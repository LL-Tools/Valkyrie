

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6537, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987;

  INV_X4 U7284 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  XNOR2_X1 U7285 ( .A(n14816), .B(n14635), .ZN(n15080) );
  NAND2_X1 U7287 ( .A1(n7847), .A2(n7846), .ZN(n14257) );
  INV_X1 U7288 ( .A(n13369), .ZN(n13031) );
  NAND2_X1 U7289 ( .A1(n9216), .A2(n9215), .ZN(n15121) );
  NAND4_X2 U7290 ( .A1(n8073), .A2(n8072), .A3(n8071), .A4(n8070), .ZN(n13979)
         );
  BUF_X2 U7291 ( .A(n10347), .Z(n9647) );
  INV_X1 U7292 ( .A(n8251), .ZN(n6855) );
  INV_X1 U7294 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n6537) );
  INV_X1 U7295 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X2 U7296 ( .A(n13743), .ZN(n13867) );
  NOR2_X1 U7297 ( .A1(n13879), .A2(n13880), .ZN(n7292) );
  AND2_X1 U7298 ( .A1(n12555), .A2(n8807), .ZN(n9321) );
  NAND2_X1 U7299 ( .A1(n9903), .A2(n7931), .ZN(n9905) );
  NAND2_X1 U7300 ( .A1(n13016), .A2(n9991), .ZN(n12862) );
  NAND3_X1 U7301 ( .A1(n9480), .A2(n9479), .A3(n10425), .ZN(n12331) );
  INV_X2 U7302 ( .A(n12331), .ZN(n9742) );
  INV_X1 U7303 ( .A(n13965), .ZN(n14119) );
  BUF_X1 U7304 ( .A(n8386), .Z(n9609) );
  AND3_X1 U7305 ( .A1(n6758), .A2(n6757), .A3(n6756), .ZN(n8222) );
  INV_X2 U7306 ( .A(n7350), .ZN(n10347) );
  INV_X1 U7307 ( .A(n15080), .ZN(n15077) );
  INV_X2 U7308 ( .A(n9321), .ZN(n10580) );
  OR2_X1 U7309 ( .A1(n9598), .A2(n9597), .ZN(n9603) );
  NAND2_X1 U7310 ( .A1(n11899), .A2(n7159), .ZN(n11900) );
  XNOR2_X1 U7311 ( .A(n9653), .B(P3_IR_REG_29__SCAN_IN), .ZN(n9663) );
  XNOR2_X1 U7312 ( .A(n8682), .B(n8680), .ZN(n13661) );
  INV_X2 U7313 ( .A(n10347), .ZN(n10425) );
  NAND2_X1 U7314 ( .A1(n9268), .A2(n9267), .ZN(n15093) );
  XNOR2_X1 U7315 ( .A(n9590), .B(n9589), .ZN(n12318) );
  XNOR2_X1 U7316 ( .A(n8886), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14676) );
  INV_X1 U7317 ( .A(n15688), .ZN(n13405) );
  OAI21_X1 U7318 ( .B1(n14072), .B2(n8461), .A(n8465), .ZN(n14046) );
  NAND4_X2 U7319 ( .A1(n8113), .A2(n8112), .A3(n8111), .A4(n8110), .ZN(n13977)
         );
  INV_X1 U7320 ( .A(n14293), .ZN(n14308) );
  BUF_X4 U7321 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n15497) );
  AND2_X1 U7322 ( .A1(n8904), .A2(n8903), .ZN(n11674) );
  INV_X1 U7323 ( .A(n15399), .ZN(n15418) );
  AOI21_X2 U7324 ( .B1(n7769), .B2(n8147), .A(n7768), .ZN(n7767) );
  OAI21_X2 U7325 ( .B1(n8436), .B2(n8435), .A(n8002), .ZN(n8553) );
  NAND4_X2 U7326 ( .A1(n8052), .A2(n8051), .A3(n8050), .A4(n8049), .ZN(n13980)
         );
  INV_X1 U7327 ( .A(n9697), .ZN(n6539) );
  OAI22_X1 U7328 ( .A1(n14069), .A2(n14068), .B1(n14413), .B2(n13866), .ZN(
        n14035) );
  NAND2_X1 U7329 ( .A1(n8048), .A2(n9647), .ZN(n6540) );
  INV_X4 U7330 ( .A(n8043), .ZN(n8102) );
  OAI21_X2 U7331 ( .B1(n6748), .B2(n6747), .A(n6744), .ZN(n12906) );
  NAND2_X4 U7332 ( .A1(n15642), .A2(n13937), .ZN(n8587) );
  XNOR2_X2 U7333 ( .A(n8806), .B(n8805), .ZN(n12556) );
  XNOR2_X2 U7334 ( .A(n8454), .B(n8453), .ZN(n8541) );
  OAI21_X2 U7335 ( .B1(n8452), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8454) );
  NAND2_X2 U7336 ( .A1(n8382), .A2(n8381), .ZN(n14345) );
  BUF_X4 U7337 ( .A(n9715), .Z(n9722) );
  AND2_X1 U7338 ( .A1(n15262), .A2(n15263), .ZN(n15270) );
  INV_X1 U7339 ( .A(n13973), .ZN(n11435) );
  INV_X1 U7340 ( .A(n11669), .ZN(n12813) );
  BUF_X2 U7341 ( .A(n8074), .Z(n9606) );
  MUX2_X1 U7342 ( .A(n10258), .B(n10257), .S(n13405), .Z(n10267) );
  AOI21_X1 U7343 ( .B1(n12481), .B2(n12523), .A(n12480), .ZN(n12515) );
  OR2_X1 U7344 ( .A1(n10260), .A2(n13540), .ZN(n10249) );
  AND3_X1 U7345 ( .A1(n6934), .A2(n6932), .A3(n6930), .ZN(n10257) );
  OR2_X1 U7346 ( .A1(n10260), .A2(n13488), .ZN(n10236) );
  XNOR2_X1 U7347 ( .A(n13323), .B(n13322), .ZN(n13453) );
  NAND2_X1 U7348 ( .A1(n13333), .A2(n10228), .ZN(n13323) );
  OAI21_X1 U7349 ( .B1(n7300), .B2(n6797), .A(n15478), .ZN(n6796) );
  MUX2_X1 U7350 ( .A(n15198), .B(n15197), .S(n15478), .Z(n15199) );
  NAND2_X1 U7351 ( .A1(n14483), .A2(n9283), .ZN(n9328) );
  INV_X1 U7352 ( .A(n12884), .ZN(n13296) );
  NAND2_X1 U7353 ( .A1(n15074), .A2(n7164), .ZN(n7300) );
  AND2_X1 U7354 ( .A1(n15090), .A2(n15091), .ZN(n7172) );
  NAND2_X1 U7355 ( .A1(n6906), .A2(n7100), .ZN(n15096) );
  AOI21_X1 U7356 ( .B1(n12820), .B2(n12819), .A(n12818), .ZN(n14069) );
  AOI211_X1 U7357 ( .C1(n14031), .C2(n14030), .A(n8582), .B(n14029), .ZN(
        n14319) );
  NAND2_X1 U7358 ( .A1(n13645), .A2(n13644), .ZN(n12893) );
  XNOR2_X1 U7359 ( .A(n12991), .B(n13324), .ZN(n13312) );
  AND2_X1 U7360 ( .A1(n7253), .A2(n7255), .ZN(n15083) );
  INV_X1 U7361 ( .A(n12817), .ZN(n12820) );
  AOI21_X1 U7362 ( .B1(n15073), .B2(n15377), .A(n15072), .ZN(n15074) );
  CLKBUF_X1 U7363 ( .A(n14125), .Z(n7128) );
  NAND2_X1 U7364 ( .A1(n10141), .A2(n10140), .ZN(n13327) );
  OAI21_X1 U7365 ( .B1(n14125), .B2(n7640), .A(n7638), .ZN(n12817) );
  AND2_X1 U7366 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  NAND2_X1 U7367 ( .A1(n7676), .A2(n6910), .ZN(n7911) );
  OAI21_X1 U7368 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(n10181) );
  NAND2_X1 U7369 ( .A1(n9601), .A2(n9600), .ZN(n14031) );
  INV_X1 U7370 ( .A(n14322), .ZN(n14040) );
  AOI21_X1 U7371 ( .B1(n6651), .B2(n7869), .A(n7866), .ZN(n7865) );
  NAND2_X1 U7372 ( .A1(n6767), .A2(n7859), .ZN(n14598) );
  NAND2_X1 U7373 ( .A1(n7273), .A2(n7815), .ZN(n14923) );
  NAND3_X1 U7374 ( .A1(n6953), .A2(n9869), .A3(n6952), .ZN(n12294) );
  OAI21_X1 U7375 ( .B1(n10023), .B2(n7718), .A(n7717), .ZN(n10136) );
  NAND2_X1 U7376 ( .A1(n9278), .A2(n9277), .ZN(n14856) );
  NAND2_X1 U7377 ( .A1(n6913), .A2(n6912), .ZN(n15024) );
  AND2_X1 U7378 ( .A1(n13862), .A2(n13963), .ZN(n12818) );
  INV_X1 U7379 ( .A(n14082), .ZN(n13862) );
  NAND2_X1 U7380 ( .A1(n9959), .A2(n9971), .ZN(n9972) );
  NAND2_X1 U7381 ( .A1(n7874), .A2(n11377), .ZN(n12018) );
  NAND2_X1 U7382 ( .A1(n9958), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9971) );
  NAND2_X1 U7383 ( .A1(n9232), .A2(n9231), .ZN(n15111) );
  OR2_X1 U7384 ( .A1(n9958), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9959) );
  NAND2_X1 U7385 ( .A1(n11379), .A2(n11378), .ZN(n11377) );
  NAND2_X1 U7386 ( .A1(n11272), .A2(n8962), .ZN(n11379) );
  NOR2_X1 U7387 ( .A1(n11890), .A2(n6588), .ZN(n7877) );
  NAND2_X1 U7388 ( .A1(n8356), .A2(n8355), .ZN(n14196) );
  NAND2_X1 U7389 ( .A1(n8335), .A2(n8334), .ZN(n14365) );
  NOR2_X2 U7390 ( .A1(n11945), .A2(n15188), .ZN(n12106) );
  NAND2_X1 U7391 ( .A1(n7597), .A2(n7594), .ZN(n7593) );
  NAND2_X1 U7392 ( .A1(n8269), .A2(n8268), .ZN(n14383) );
  OR2_X1 U7393 ( .A1(n8319), .A2(n7973), .ZN(n7597) );
  NAND2_X1 U7394 ( .A1(n8255), .A2(n8254), .ZN(n14389) );
  OAI21_X1 U7395 ( .B1(n7248), .B2(n7247), .A(n7245), .ZN(n12064) );
  NAND2_X1 U7396 ( .A1(n8212), .A2(n8211), .ZN(n14405) );
  NAND2_X1 U7397 ( .A1(n8192), .A2(n8191), .ZN(n13794) );
  NAND2_X1 U7398 ( .A1(n8968), .A2(n8967), .ZN(n12598) );
  NAND2_X1 U7399 ( .A1(n8237), .A2(n8236), .ZN(n14393) );
  NAND2_X1 U7400 ( .A1(n12372), .A2(n12371), .ZN(n12483) );
  NAND2_X1 U7401 ( .A1(n9065), .A2(n9064), .ZN(n15188) );
  AND2_X1 U7402 ( .A1(n8956), .A2(n8955), .ZN(n15440) );
  NAND2_X1 U7403 ( .A1(n8145), .A2(n8144), .ZN(n13777) );
  INV_X1 U7404 ( .A(n13726), .ZN(n13727) );
  NAND2_X1 U7405 ( .A1(n8174), .A2(n8173), .ZN(n13789) );
  NAND2_X1 U7406 ( .A1(n9048), .A2(n9047), .ZN(n12619) );
  NAND2_X1 U7407 ( .A1(n7918), .A2(n9736), .ZN(n13114) );
  NAND2_X1 U7408 ( .A1(n6850), .A2(n6849), .ZN(n13904) );
  NAND2_X2 U7409 ( .A1(n8809), .A2(n15397), .ZN(n9136) );
  NAND2_X1 U7410 ( .A1(n7190), .A2(n6597), .ZN(n13111) );
  XNOR2_X1 U7411 ( .A(n8155), .B(n8154), .ZN(n10390) );
  AND4_X1 U7412 ( .A1(n9726), .A2(n9725), .A3(n9724), .A4(n9723), .ZN(n11414)
         );
  NAND4_X1 U7413 ( .A1(n8178), .A2(n8177), .A3(n8176), .A4(n8175), .ZN(n13974)
         );
  AND2_X1 U7414 ( .A1(n8912), .A2(n6897), .ZN(n12581) );
  AND2_X1 U7415 ( .A1(n8917), .A2(n8916), .ZN(n15427) );
  NAND2_X2 U7416 ( .A1(n8853), .A2(n12719), .ZN(n8958) );
  AND2_X1 U7417 ( .A1(n6539), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9698) );
  NAND2_X1 U7418 ( .A1(n8201), .A2(n8167), .ZN(n8181) );
  XNOR2_X1 U7419 ( .A(n8116), .B(n8115), .ZN(n10392) );
  NAND4_X2 U7420 ( .A1(n8093), .A2(n8092), .A3(n8091), .A4(n8090), .ZN(n13978)
         );
  NAND4_X1 U7421 ( .A1(n8130), .A2(n8129), .A3(n8128), .A4(n8127), .ZN(n13976)
         );
  INV_X2 U7422 ( .A(n8570), .ZN(n12833) );
  INV_X4 U7423 ( .A(n8587), .ZN(n8687) );
  NAND4_X1 U7424 ( .A1(n8851), .A2(n8850), .A3(n8849), .A4(n8848), .ZN(n12041)
         );
  CLKBUF_X3 U7425 ( .A(n8068), .Z(n8721) );
  AND3_X2 U7426 ( .A1(n8874), .A2(n8873), .A3(n6605), .ZN(n15410) );
  AND2_X2 U7427 ( .A1(n12964), .A2(n9662), .ZN(n9746) );
  NAND2_X1 U7428 ( .A1(n10706), .A2(n10707), .ZN(n10705) );
  CLKBUF_X2 U7429 ( .A(n8131), .Z(n8148) );
  AND2_X2 U7430 ( .A1(n8792), .A2(n8793), .ZN(n9310) );
  NAND2_X1 U7431 ( .A1(n9629), .A2(n9628), .ZN(n10043) );
  AOI21_X1 U7432 ( .B1(n8095), .B2(n8098), .A(n8100), .ZN(n7941) );
  XNOR2_X1 U7433 ( .A(n9468), .B(n9470), .ZN(n12526) );
  MUX2_X1 U7434 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9627), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n9629) );
  INV_X2 U7435 ( .A(n7072), .ZN(n9944) );
  INV_X2 U7436 ( .A(n7916), .ZN(n9573) );
  NAND2_X2 U7437 ( .A1(n12720), .A2(n12557), .ZN(n15397) );
  OR2_X1 U7438 ( .A1(n9471), .A2(n9370), .ZN(n9473) );
  INV_X1 U7439 ( .A(n8792), .ZN(n15224) );
  NAND2_X1 U7440 ( .A1(n7680), .A2(n7677), .ZN(n15227) );
  NAND2_X2 U7441 ( .A1(n9335), .A2(n15230), .ZN(n8832) );
  AND2_X1 U7442 ( .A1(n11695), .A2(n12558), .ZN(n12719) );
  NAND2_X2 U7443 ( .A1(n10490), .A2(n13953), .ZN(n8048) );
  OR2_X1 U7444 ( .A1(n8791), .A2(n7681), .ZN(n7680) );
  NAND2_X1 U7445 ( .A1(n8759), .A2(n8760), .ZN(n15230) );
  XNOR2_X1 U7446 ( .A(n8456), .B(P2_IR_REG_21__SCAN_IN), .ZN(n13941) );
  OR2_X1 U7447 ( .A1(n8472), .A2(n8266), .ZN(n8451) );
  INV_X2 U7448 ( .A(n15221), .ZN(n15236) );
  OR2_X1 U7449 ( .A1(n9467), .A2(n7567), .ZN(n9626) );
  NOR2_X1 U7450 ( .A1(n9467), .A2(n7568), .ZN(n9471) );
  AND2_X1 U7451 ( .A1(n8789), .A2(n8756), .ZN(n8791) );
  OAI21_X1 U7452 ( .B1(n9100), .B2(n8804), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8806) );
  CLKBUF_X1 U7453 ( .A(n9650), .Z(n9654) );
  NAND2_X1 U7454 ( .A1(n6916), .A2(SI_0_), .ZN(n8053) );
  XNOR2_X1 U7455 ( .A(n7946), .B(SI_6_), .ZN(n8133) );
  CLKBUF_X1 U7456 ( .A(n8802), .Z(n8803) );
  AND3_X1 U7457 ( .A1(n9389), .A2(n7562), .A3(n9357), .ZN(n9380) );
  NOR2_X1 U7458 ( .A1(n8744), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n6890) );
  NOR2_X1 U7459 ( .A1(n8763), .A2(n8921), .ZN(n8802) );
  OR2_X1 U7460 ( .A1(n8161), .A2(n8160), .ZN(n8195) );
  AND2_X1 U7461 ( .A1(n9487), .A2(n9486), .ZN(n9389) );
  NAND4_X2 U7462 ( .A1(n14653), .A2(n8870), .A3(n8749), .A4(n8748), .ZN(n8921)
         );
  AND3_X1 U7463 ( .A1(n9360), .A2(n9359), .A3(n9358), .ZN(n9494) );
  NOR2_X1 U7464 ( .A1(n7784), .A2(n8266), .ZN(n7020) );
  AND3_X1 U7465 ( .A1(n8006), .A2(n8005), .A3(n8004), .ZN(n8351) );
  NAND2_X1 U7466 ( .A1(n6763), .A2(n8743), .ZN(n8744) );
  NAND2_X1 U7467 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n15497), .ZN(n8042) );
  AND2_X1 U7468 ( .A1(n9486), .A2(n9379), .ZN(n7561) );
  NOR2_X1 U7469 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8004) );
  NOR2_X1 U7470 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8005) );
  NOR2_X1 U7471 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6765) );
  NOR2_X1 U7472 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6763) );
  NOR2_X1 U7473 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8006) );
  NOR2_X1 U7474 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8746) );
  INV_X1 U7475 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8805) );
  NOR2_X1 U7476 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n8745) );
  INV_X1 U7477 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8483) );
  NOR2_X1 U7478 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n8751) );
  NOR2_X1 U7479 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n8750) );
  NOR2_X1 U7480 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6764) );
  INV_X1 U7481 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9365) );
  INV_X1 U7482 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9004) );
  INV_X1 U7483 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9408) );
  INV_X1 U7484 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7935) );
  INV_X1 U7485 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7295) );
  INV_X2 U7486 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8870) );
  NOR2_X2 U7487 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9487) );
  INV_X1 U7488 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9486) );
  NOR2_X1 U7489 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n9382) );
  INV_X1 U7490 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8749) );
  INV_X4 U7491 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7492 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8748) );
  NOR2_X1 U7493 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9353) );
  INV_X1 U7494 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n15697) );
  INV_X1 U7495 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9443) );
  AOI21_X2 U7496 ( .B1(n7566), .B2(n7565), .A(n7563), .ZN(n11784) );
  NAND2_X1 U7497 ( .A1(n8148), .A2(n8136), .ZN(n8116) );
  INV_X4 U7498 ( .A(n9790), .ZN(n9995) );
  NAND2_X2 U7499 ( .A1(n7101), .A2(n9288), .ZN(n8853) );
  INV_X1 U7500 ( .A(n7350), .ZN(n6541) );
  NAND2_X1 U7501 ( .A1(n6542), .A2(n10348), .ZN(n8066) );
  AOI21_X2 U7502 ( .B1(n7939), .B2(n7938), .A(n7929), .ZN(n8098) );
  INV_X2 U7503 ( .A(n13768), .ZN(n13743) );
  NAND2_X2 U7504 ( .A1(n12964), .A2(n13545), .ZN(n9697) );
  INV_X1 U7505 ( .A(n8043), .ZN(n6542) );
  INV_X1 U7506 ( .A(n9136), .ZN(n6543) );
  AND2_X4 U7507 ( .A1(n8832), .A2(n10425), .ZN(n8868) );
  NOR2_X4 U7508 ( .A1(n14257), .A2(n14372), .ZN(n14242) );
  INV_X1 U7509 ( .A(n6908), .ZN(n6907) );
  OAI21_X1 U7510 ( .B1(n6910), .B2(n6909), .A(n14850), .ZN(n6908) );
  INV_X1 U7511 ( .A(n12953), .ZN(n6909) );
  NAND2_X1 U7512 ( .A1(n13861), .A2(n7723), .ZN(n7722) );
  INV_X1 U7513 ( .A(n7963), .ZN(n7575) );
  NOR2_X1 U7514 ( .A1(n10011), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7232) );
  NOR2_X1 U7515 ( .A1(n8459), .A2(n13563), .ZN(n8565) );
  INV_X1 U7516 ( .A(n7330), .ZN(n7329) );
  OAI21_X1 U7517 ( .B1(n7331), .B2(n7335), .A(n8296), .ZN(n7330) );
  INV_X1 U7518 ( .A(n7332), .ZN(n7331) );
  NAND2_X1 U7519 ( .A1(n8048), .A2(n10425), .ZN(n8074) );
  NAND2_X1 U7520 ( .A1(n15087), .A2(n14837), .ZN(n12983) );
  AOI21_X1 U7521 ( .B1(n12751), .B2(n7812), .A(n6637), .ZN(n7811) );
  AND2_X1 U7522 ( .A1(n9663), .A2(n13545), .ZN(n9759) );
  AND2_X1 U7523 ( .A1(n10395), .A2(n10082), .ZN(n10242) );
  NAND2_X1 U7524 ( .A1(n8048), .A2(n9647), .ZN(n8043) );
  NAND2_X1 U7525 ( .A1(n8022), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8439) );
  INV_X1 U7526 ( .A(n8428), .ZN(n8022) );
  AND2_X1 U7527 ( .A1(n12839), .A2(n12821), .ZN(n14043) );
  NAND2_X1 U7528 ( .A1(n8855), .A2(n6775), .ZN(n11000) );
  OR2_X1 U7529 ( .A1(n12036), .A2(n9136), .ZN(n6775) );
  AOI22_X1 U7530 ( .A1(n8854), .A2(n12038), .B1(n8856), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n8855) );
  INV_X1 U7531 ( .A(n9310), .ZN(n9273) );
  AND4_X1 U7532 ( .A1(n12925), .A2(n12924), .A3(n12923), .A4(n12922), .ZN(
        n12926) );
  INV_X1 U7533 ( .A(n7103), .ZN(n12917) );
  NOR2_X1 U7534 ( .A1(n14885), .A2(n7675), .ZN(n7674) );
  INV_X1 U7535 ( .A(n12951), .ZN(n7675) );
  OR2_X1 U7536 ( .A1(n12600), .A2(n12599), .ZN(n11933) );
  XNOR2_X1 U7537 ( .A(n8790), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U7538 ( .A1(n15219), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U7539 ( .A1(n9264), .A2(n7075), .ZN(n14483) );
  OR2_X1 U7540 ( .A1(n9266), .A2(n9265), .ZN(n7075) );
  NAND2_X1 U7541 ( .A1(n12587), .A2(n12589), .ZN(n6989) );
  OR2_X1 U7542 ( .A1(n12681), .A2(n12680), .ZN(n12682) );
  AND2_X1 U7543 ( .A1(n7722), .A2(n13856), .ZN(n7720) );
  AOI21_X1 U7544 ( .B1(n7213), .B2(n7211), .A(n6624), .ZN(n7210) );
  INV_X1 U7545 ( .A(n10096), .ZN(n7211) );
  NAND2_X1 U7546 ( .A1(n11133), .A2(n10105), .ZN(n11050) );
  INV_X1 U7547 ( .A(n7070), .ZN(n7069) );
  OAI21_X1 U7548 ( .B1(n9928), .B2(n7071), .A(n9955), .ZN(n7070) );
  INV_X1 U7549 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U7550 ( .A1(n7058), .A2(n9755), .ZN(n7057) );
  INV_X1 U7551 ( .A(n9640), .ZN(n7058) );
  NOR2_X1 U7552 ( .A1(n6854), .A2(n13745), .ZN(n6851) );
  NAND2_X1 U7553 ( .A1(n8417), .A2(n7991), .ZN(n7995) );
  AOI21_X1 U7554 ( .B1(n7980), .B2(n8348), .A(n7979), .ZN(n7981) );
  OAI21_X1 U7555 ( .B1(n10319), .B2(n10318), .A(n10317), .ZN(n10375) );
  NAND2_X1 U7556 ( .A1(n9990), .A2(n9989), .ZN(n9991) );
  NOR2_X1 U7557 ( .A1(n13142), .A2(n6886), .ZN(n9422) );
  NOR2_X1 U7558 ( .A1(n9671), .A2(n11162), .ZN(n6886) );
  INV_X1 U7559 ( .A(n10915), .ZN(n7399) );
  OR2_X1 U7560 ( .A1(n9511), .A2(n7439), .ZN(n7434) );
  AND2_X1 U7561 ( .A1(n7436), .A2(n10482), .ZN(n7435) );
  OR2_X1 U7562 ( .A1(n13174), .A2(n7443), .ZN(n7436) );
  NAND2_X1 U7563 ( .A1(n7216), .A2(n7214), .ZN(n13308) );
  NOR2_X1 U7564 ( .A1(n13312), .A2(n7215), .ZN(n7214) );
  INV_X1 U7565 ( .A(n7217), .ZN(n7215) );
  NAND2_X1 U7566 ( .A1(n7237), .A2(n13369), .ZN(n12454) );
  OR2_X1 U7567 ( .A1(n11050), .A2(n12491), .ZN(n7207) );
  AND2_X1 U7568 ( .A1(n12497), .A2(n10108), .ZN(n7898) );
  OR2_X1 U7569 ( .A1(n13110), .A2(n11644), .ZN(n12393) );
  NAND2_X1 U7570 ( .A1(n12393), .A2(n12394), .ZN(n7213) );
  NAND2_X1 U7571 ( .A1(n11206), .A2(n11657), .ZN(n12384) );
  INV_X1 U7572 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n9732) );
  OR2_X1 U7573 ( .A1(n10178), .A2(n10201), .ZN(n12471) );
  NAND2_X1 U7574 ( .A1(n10127), .A2(n6630), .ZN(n13337) );
  NOR2_X1 U7575 ( .A1(n13351), .A2(n7195), .ZN(n7194) );
  INV_X1 U7576 ( .A(n12453), .ZN(n7195) );
  OR2_X1 U7577 ( .A1(n13521), .A2(n13022), .ZN(n12348) );
  AND2_X1 U7578 ( .A1(n10113), .A2(n7892), .ZN(n7891) );
  NAND2_X1 U7579 ( .A1(n7893), .A2(n10112), .ZN(n7892) );
  OR2_X1 U7580 ( .A1(n9483), .A2(n9475), .ZN(n9480) );
  AND2_X1 U7581 ( .A1(n9480), .A2(n9479), .ZN(n7072) );
  NOR2_X1 U7582 ( .A1(n10007), .A2(n7697), .ZN(n7696) );
  INV_X1 U7583 ( .A(n9992), .ZN(n7697) );
  AND2_X1 U7584 ( .A1(n7561), .A2(n9487), .ZN(n7560) );
  INV_X1 U7585 ( .A(n7701), .ZN(n7700) );
  OAI21_X1 U7586 ( .B1(n7703), .B2(n7702), .A(n9681), .ZN(n7701) );
  NOR2_X1 U7587 ( .A1(n11431), .A2(n7793), .ZN(n7792) );
  INV_X1 U7588 ( .A(n8619), .ZN(n7793) );
  AND2_X1 U7589 ( .A1(n13980), .A2(n8582), .ZN(n13673) );
  XNOR2_X1 U7590 ( .A(n13741), .B(n8587), .ZN(n13672) );
  OAI21_X1 U7591 ( .B1(n13865), .B2(n13864), .A(n13863), .ZN(n13878) );
  OAI21_X1 U7592 ( .B1(n7329), .B2(n6735), .A(n8315), .ZN(n6734) );
  NOR2_X1 U7593 ( .A1(n8526), .A2(n7623), .ZN(n7622) );
  INV_X1 U7594 ( .A(n7625), .ZN(n7623) );
  AOI21_X1 U7595 ( .B1(n7335), .B2(n7333), .A(n6634), .ZN(n7332) );
  INV_X1 U7596 ( .A(n6593), .ZN(n7333) );
  NAND2_X1 U7597 ( .A1(n10898), .A2(n13904), .ZN(n10897) );
  AND2_X1 U7598 ( .A1(n15610), .A2(n8498), .ZN(n8704) );
  NAND2_X1 U7599 ( .A1(n14138), .A2(n8536), .ZN(n14125) );
  AND2_X1 U7600 ( .A1(n8541), .A2(n13941), .ZN(n13747) );
  INV_X1 U7601 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7787) );
  NOR2_X1 U7602 ( .A1(n8171), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7145) );
  OR2_X1 U7603 ( .A1(n14955), .A2(n14964), .ZN(n12949) );
  OR2_X1 U7604 ( .A1(n15150), .A2(n14602), .ZN(n12767) );
  OR2_X1 U7605 ( .A1(n15171), .A2(n14541), .ZN(n12909) );
  NAND2_X1 U7606 ( .A1(n12708), .A2(n12707), .ZN(n14816) );
  NOR2_X1 U7607 ( .A1(n6578), .A2(n6723), .ZN(n7599) );
  NAND2_X1 U7608 ( .A1(n8555), .A2(n8554), .ZN(n8700) );
  OAI21_X1 U7609 ( .B1(n8553), .B2(n15772), .A(n8552), .ZN(n8555) );
  NOR2_X1 U7610 ( .A1(n7982), .A2(n7595), .ZN(n7594) );
  INV_X1 U7611 ( .A(n7975), .ZN(n7595) );
  NAND3_X1 U7612 ( .A1(n8765), .A2(n6774), .A3(n7097), .ZN(n7096) );
  INV_X1 U7613 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7097) );
  INV_X1 U7614 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9302) );
  XNOR2_X1 U7615 ( .A(n8345), .B(SI_18_), .ZN(n8344) );
  INV_X1 U7616 ( .A(n7574), .ZN(n7573) );
  OAI21_X1 U7617 ( .B1(n8249), .B2(n7575), .A(n7967), .ZN(n7574) );
  XNOR2_X1 U7618 ( .A(n7971), .B(SI_16_), .ZN(n8299) );
  NAND4_X1 U7619 ( .A1(n7296), .A2(n7295), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6785) );
  INV_X1 U7620 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7296) );
  NAND2_X1 U7621 ( .A1(n10384), .A2(n10383), .ZN(n10753) );
  OAI22_X1 U7622 ( .A1(n12098), .A2(n12097), .B1(P3_ADDR_REG_11__SCAN_IN), 
        .B2(n14766), .ZN(n15255) );
  NAND2_X1 U7623 ( .A1(n7530), .A2(n7533), .ZN(n7529) );
  INV_X1 U7624 ( .A(n13088), .ZN(n7530) );
  NAND2_X1 U7625 ( .A1(n11900), .A2(n7915), .ZN(n12237) );
  INV_X1 U7626 ( .A(n13324), .ZN(n12888) );
  INV_X1 U7627 ( .A(n13118), .ZN(n11415) );
  NAND2_X1 U7628 ( .A1(n6948), .A2(n6947), .ZN(n7566) );
  INV_X1 U7629 ( .A(n11629), .ZN(n6947) );
  NOR2_X1 U7630 ( .A1(n9924), .A2(n7541), .ZN(n7540) );
  INV_X1 U7631 ( .A(n9904), .ZN(n7541) );
  NAND2_X1 U7632 ( .A1(n10029), .A2(n10073), .ZN(n10080) );
  INV_X1 U7633 ( .A(n9759), .ZN(n10189) );
  OR2_X1 U7634 ( .A1(n9422), .A2(n9544), .ZN(n7400) );
  NAND2_X1 U7635 ( .A1(n13201), .A2(n9564), .ZN(n13203) );
  NAND2_X1 U7636 ( .A1(n9460), .A2(n13260), .ZN(n13268) );
  AND2_X1 U7637 ( .A1(n6809), .A2(n6806), .ZN(n6805) );
  INV_X1 U7638 ( .A(n13276), .ZN(n6806) );
  AND2_X1 U7639 ( .A1(n6966), .A2(n9515), .ZN(n6965) );
  NAND2_X1 U7640 ( .A1(n10229), .A2(n12469), .ZN(n13295) );
  NAND2_X1 U7641 ( .A1(n13311), .A2(n13312), .ZN(n10229) );
  NAND2_X1 U7642 ( .A1(n13366), .A2(n12509), .ZN(n10227) );
  OR2_X1 U7643 ( .A1(n13373), .A2(n13073), .ZN(n12453) );
  OR2_X1 U7644 ( .A1(n9962), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U7645 ( .A1(n11645), .A2(n11169), .ZN(n12392) );
  INV_X1 U7646 ( .A(n12353), .ZN(n7197) );
  NAND2_X1 U7647 ( .A1(n13416), .A2(n10121), .ZN(n12540) );
  OR2_X1 U7648 ( .A1(n13535), .A2(n13101), .ZN(n12353) );
  AND2_X1 U7649 ( .A1(n7740), .A2(n10118), .ZN(n7899) );
  OR2_X1 U7650 ( .A1(n13484), .A2(n13413), .ZN(n12356) );
  NAND2_X1 U7651 ( .A1(n6873), .A2(n7739), .ZN(n13422) );
  AOI21_X1 U7652 ( .B1(n7743), .B2(n7742), .A(n7740), .ZN(n7739) );
  NAND2_X1 U7653 ( .A1(n12197), .A2(n6559), .ZN(n6873) );
  NAND2_X1 U7654 ( .A1(n12197), .A2(n12501), .ZN(n7744) );
  NAND2_X1 U7655 ( .A1(n7221), .A2(n7219), .ZN(n12277) );
  AOI21_X1 U7656 ( .B1(n7222), .B2(n7223), .A(n7220), .ZN(n7219) );
  NAND2_X1 U7657 ( .A1(n10116), .A2(n7222), .ZN(n7221) );
  NAND2_X1 U7658 ( .A1(n12142), .A2(n12422), .ZN(n10116) );
  NAND2_X1 U7659 ( .A1(n7072), .A2(n9647), .ZN(n9790) );
  NAND2_X1 U7660 ( .A1(n12531), .A2(n10042), .ZN(n11358) );
  AND3_X1 U7661 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(n9662) );
  NAND2_X1 U7662 ( .A1(n12799), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9653) );
  INV_X1 U7663 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U7664 ( .A1(n9929), .A2(n9928), .ZN(n9942) );
  NAND2_X1 U7665 ( .A1(n7042), .A2(n9635), .ZN(n9728) );
  NAND2_X1 U7666 ( .A1(n9389), .A2(n9355), .ZN(n9407) );
  INV_X1 U7667 ( .A(n9389), .ZN(n9403) );
  NOR2_X1 U7668 ( .A1(n12125), .A2(n7026), .ZN(n7025) );
  INV_X1 U7669 ( .A(n8634), .ZN(n7026) );
  XNOR2_X1 U7670 ( .A(n8587), .B(n15632), .ZN(n10802) );
  NAND2_X1 U7671 ( .A1(n7806), .A2(n12894), .ZN(n7805) );
  INV_X1 U7672 ( .A(n7808), .ZN(n7806) );
  NAND2_X1 U7673 ( .A1(n12893), .A2(n7807), .ZN(n7804) );
  NOR2_X1 U7674 ( .A1(n7808), .A2(n8689), .ZN(n7807) );
  AND4_X1 U7675 ( .A1(n8166), .A2(n8165), .A3(n8164), .A4(n8163), .ZN(n11197)
         );
  AND2_X1 U7676 ( .A1(n7386), .A2(n10489), .ZN(n7378) );
  INV_X1 U7677 ( .A(n7373), .ZN(n7366) );
  AOI21_X1 U7678 ( .B1(n8722), .B2(n8721), .A(n8720), .ZN(n14047) );
  AND2_X1 U7679 ( .A1(n8573), .A2(n8572), .ZN(n14065) );
  NAND2_X1 U7680 ( .A1(n6864), .A2(n8405), .ZN(n14114) );
  AOI21_X1 U7681 ( .B1(n7622), .B2(n7621), .A(n7620), .ZN(n7619) );
  INV_X1 U7682 ( .A(n7627), .ZN(n7621) );
  INV_X1 U7683 ( .A(n13920), .ZN(n7620) );
  OAI21_X1 U7684 ( .B1(n6743), .B2(n11956), .A(n6741), .ZN(n12086) );
  NAND2_X1 U7685 ( .A1(n8458), .A2(n8457), .ZN(n14307) );
  INV_X1 U7686 ( .A(n14118), .ZN(n14304) );
  XNOR2_X1 U7687 ( .A(n14077), .B(n14046), .ZN(n14068) );
  INV_X1 U7688 ( .A(n13874), .ZN(n13875) );
  XNOR2_X1 U7689 ( .A(n13875), .B(n14047), .ZN(n13931) );
  AND2_X1 U7690 ( .A1(n8539), .A2(n10271), .ZN(n14103) );
  OAI21_X1 U7691 ( .B1(n14173), .B2(n7632), .A(n7630), .ZN(n14138) );
  INV_X1 U7692 ( .A(n7631), .ZN(n7630) );
  OAI21_X1 U7693 ( .B1(n7634), .B2(n7632), .A(n14139), .ZN(n7631) );
  INV_X2 U7694 ( .A(n8074), .ZN(n8354) );
  INV_X2 U7695 ( .A(n8048), .ZN(n8353) );
  XNOR2_X1 U7696 ( .A(n8026), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U7697 ( .A1(n8028), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8026) );
  INV_X1 U7698 ( .A(n8028), .ZN(n6746) );
  OR2_X1 U7699 ( .A1(n14500), .A2(n7870), .ZN(n7869) );
  INV_X1 U7700 ( .A(n7872), .ZN(n7870) );
  AND3_X1 U7701 ( .A1(n8859), .A2(n8858), .A3(n8857), .ZN(n11001) );
  INV_X1 U7702 ( .A(n14649), .ZN(n12812) );
  AOI21_X1 U7703 ( .B1(n7865), .B2(n7867), .A(n7863), .ZN(n7862) );
  INV_X1 U7704 ( .A(n14524), .ZN(n7863) );
  NAND2_X1 U7705 ( .A1(n14773), .A2(n6751), .ZN(n10811) );
  NOR2_X1 U7706 ( .A1(n10614), .A2(n6752), .ZN(n6751) );
  INV_X1 U7707 ( .A(n10612), .ZN(n6752) );
  OR2_X1 U7708 ( .A1(n11338), .A2(n11344), .ZN(n11440) );
  INV_X1 U7709 ( .A(n6798), .ZN(n14841) );
  AND2_X1 U7710 ( .A1(n14833), .A2(n12745), .ZN(n14853) );
  NOR2_X1 U7711 ( .A1(n14880), .A2(n6911), .ZN(n6910) );
  INV_X1 U7712 ( .A(n12952), .ZN(n6911) );
  NAND2_X1 U7713 ( .A1(n14972), .A2(n6915), .ZN(n7308) );
  AND2_X1 U7714 ( .A1(n6698), .A2(n12946), .ZN(n6915) );
  AOI21_X1 U7715 ( .B1(n7818), .B2(n7816), .A(n6646), .ZN(n7815) );
  NAND2_X1 U7716 ( .A1(n7265), .A2(n7263), .ZN(n7273) );
  AOI21_X1 U7717 ( .B1(n7822), .B2(n7821), .A(n6647), .ZN(n7820) );
  INV_X1 U7718 ( .A(n12912), .ZN(n7821) );
  OR2_X1 U7719 ( .A1(n15024), .A2(n12942), .ZN(n7689) );
  NOR2_X1 U7720 ( .A1(n12749), .A2(n7830), .ZN(n7829) );
  INV_X1 U7721 ( .A(n11837), .ZN(n7830) );
  NAND2_X1 U7722 ( .A1(n12754), .A2(n12064), .ZN(n7814) );
  INV_X2 U7723 ( .A(n8832), .ZN(n9176) );
  INV_X1 U7724 ( .A(n15397), .ZN(n15377) );
  INV_X1 U7725 ( .A(n8804), .ZN(n6889) );
  INV_X1 U7726 ( .A(n15219), .ZN(n7679) );
  INV_X1 U7727 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8756) );
  XNOR2_X1 U7728 ( .A(n10752), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n10387) );
  NAND2_X1 U7729 ( .A1(n7488), .A2(n7491), .ZN(n12103) );
  AND2_X1 U7730 ( .A1(n9377), .A2(n10047), .ZN(n9378) );
  NAND2_X1 U7731 ( .A1(n8438), .A2(n8437), .ZN(n13859) );
  NAND2_X1 U7732 ( .A1(n8445), .A2(n8444), .ZN(n13964) );
  INV_X1 U7733 ( .A(n14413), .ZN(n14077) );
  AND2_X1 U7734 ( .A1(n9284), .A2(n9285), .ZN(n7101) );
  NAND2_X2 U7735 ( .A1(n7080), .A2(n7081), .ZN(n14586) );
  AOI21_X1 U7736 ( .B1(n7880), .B2(n7882), .A(n7082), .ZN(n7081) );
  NAND2_X1 U7737 ( .A1(n14578), .A2(n7880), .ZN(n7080) );
  INV_X1 U7738 ( .A(n14588), .ZN(n7082) );
  NAND2_X1 U7739 ( .A1(n9317), .A2(n9316), .ZN(n14837) );
  NAND2_X1 U7740 ( .A1(n8799), .A2(n8798), .ZN(n14870) );
  NAND2_X1 U7741 ( .A1(n9255), .A2(n9254), .ZN(n14887) );
  OR2_X1 U7742 ( .A1(n14874), .A2(n9273), .ZN(n9255) );
  NAND2_X1 U7743 ( .A1(n9239), .A2(n9238), .ZN(n14907) );
  OR2_X1 U7744 ( .A1(n14894), .A2(n9273), .ZN(n9239) );
  NAND2_X1 U7745 ( .A1(n6860), .A2(n9474), .ZN(n6859) );
  NAND2_X1 U7746 ( .A1(n7885), .A2(n12368), .ZN(n6860) );
  AND2_X1 U7747 ( .A1(n7729), .A2(n6693), .ZN(n7283) );
  NAND2_X1 U7748 ( .A1(n13819), .A2(n13821), .ZN(n7729) );
  INV_X1 U7749 ( .A(n13822), .ZN(n7287) );
  NAND2_X1 U7750 ( .A1(n12580), .A2(n12579), .ZN(n12584) );
  AOI21_X1 U7751 ( .B1(n12640), .B2(n7429), .A(n7428), .ZN(n7427) );
  NAND2_X1 U7752 ( .A1(n12660), .A2(n12653), .ZN(n7428) );
  NOR2_X1 U7753 ( .A1(n12633), .A2(n7430), .ZN(n7429) );
  AND2_X1 U7754 ( .A1(n6993), .A2(n12668), .ZN(n6992) );
  NAND2_X1 U7755 ( .A1(n12665), .A2(n6994), .ZN(n6993) );
  INV_X1 U7756 ( .A(n12665), .ZN(n6996) );
  NAND2_X1 U7757 ( .A1(n7282), .A2(n13842), .ZN(n7280) );
  AOI21_X1 U7758 ( .B1(n7482), .B2(n7480), .A(n7479), .ZN(n12681) );
  NOR2_X1 U7759 ( .A1(n12677), .A2(n12676), .ZN(n7479) );
  AND2_X1 U7760 ( .A1(n7481), .A2(n12675), .ZN(n7480) );
  AND2_X1 U7761 ( .A1(n13427), .A2(n7220), .ZN(n6846) );
  INV_X1 U7762 ( .A(n12444), .ZN(n7137) );
  NAND2_X1 U7763 ( .A1(n12686), .A2(n12688), .ZN(n7185) );
  NOR2_X1 U7764 ( .A1(n6564), .A2(n6650), .ZN(n7009) );
  NAND2_X1 U7765 ( .A1(n12698), .A2(n7469), .ZN(n7468) );
  INV_X1 U7766 ( .A(n12697), .ZN(n7469) );
  INV_X1 U7767 ( .A(n12468), .ZN(n6837) );
  OAI21_X1 U7768 ( .B1(n6555), .B2(n6861), .A(n7181), .ZN(n7136) );
  AND2_X1 U7769 ( .A1(n13322), .A2(n12464), .ZN(n7181) );
  NAND2_X1 U7770 ( .A1(n12468), .A2(n6836), .ZN(n6835) );
  INV_X1 U7771 ( .A(n13312), .ZN(n6836) );
  NOR2_X1 U7772 ( .A1(n10969), .A2(n9504), .ZN(n9505) );
  AND2_X1 U7773 ( .A1(n10329), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9504) );
  INV_X1 U7774 ( .A(n7441), .ZN(n7439) );
  NAND2_X1 U7775 ( .A1(n13110), .A2(n11644), .ZN(n12394) );
  INV_X1 U7776 ( .A(n12409), .ZN(n7756) );
  NOR2_X1 U7777 ( .A1(n7756), .A2(n7753), .ZN(n7752) );
  INV_X1 U7778 ( .A(n12403), .ZN(n7753) );
  INV_X1 U7779 ( .A(n9941), .ZN(n7071) );
  AOI21_X1 U7780 ( .B1(n7720), .B2(n13858), .A(n6665), .ZN(n7290) );
  NOR2_X1 U7781 ( .A1(n8257), .A2(n8256), .ZN(n6791) );
  NAND2_X1 U7782 ( .A1(n7310), .A2(n12944), .ZN(n7309) );
  NAND2_X1 U7783 ( .A1(n14978), .A2(n12943), .ZN(n14995) );
  AND2_X1 U7784 ( .A1(n7579), .A2(n8406), .ZN(n7578) );
  INV_X1 U7785 ( .A(n8299), .ZN(n7090) );
  NOR2_X1 U7786 ( .A1(n7574), .A2(n7090), .ZN(n7088) );
  NAND2_X1 U7787 ( .A1(n10377), .A2(n10376), .ZN(n10382) );
  OR2_X1 U7788 ( .A1(n14714), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10761) );
  INV_X1 U7789 ( .A(n10761), .ZN(n6923) );
  INV_X1 U7790 ( .A(n10043), .ZN(n10193) );
  OAI211_X1 U7791 ( .C1(n6823), .C2(n11361), .A(n6822), .B(n6821), .ZN(n7314)
         );
  NAND2_X1 U7792 ( .A1(n6565), .A2(n6825), .ZN(n6821) );
  OR2_X1 U7793 ( .A1(n6825), .A2(n11361), .ZN(n6822) );
  NAND2_X1 U7794 ( .A1(n10337), .A2(n7389), .ZN(n7388) );
  INV_X1 U7795 ( .A(n7394), .ZN(n7389) );
  NAND2_X1 U7796 ( .A1(n7451), .A2(n6973), .ZN(n7450) );
  AND2_X1 U7797 ( .A1(n7452), .A2(n6700), .ZN(n6973) );
  AND2_X1 U7798 ( .A1(n7450), .A2(n10786), .ZN(n9507) );
  OAI21_X1 U7799 ( .B1(n6979), .B2(n6978), .A(n6977), .ZN(n9508) );
  INV_X1 U7800 ( .A(n11481), .ZN(n6978) );
  AOI21_X1 U7801 ( .B1(n11482), .B2(n11481), .A(n6982), .ZN(n6977) );
  NOR2_X1 U7802 ( .A1(n11480), .A2(n11367), .ZN(n6982) );
  NAND2_X1 U7803 ( .A1(n13188), .A2(n9437), .ZN(n9441) );
  OR2_X1 U7804 ( .A1(n7439), .A2(n13174), .ZN(n7438) );
  NAND2_X1 U7805 ( .A1(n10156), .A2(n15909), .ZN(n10171) );
  INV_X1 U7806 ( .A(n10157), .ZN(n10156) );
  NOR2_X1 U7807 ( .A1(n6544), .A2(n7202), .ZN(n7201) );
  AND2_X1 U7808 ( .A1(n9914), .A2(n7243), .ZN(n7242) );
  INV_X1 U7809 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7243) );
  INV_X1 U7810 ( .A(n9916), .ZN(n9915) );
  INV_X1 U7811 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7240) );
  INV_X1 U7812 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9845) );
  INV_X1 U7813 ( .A(n9847), .ZN(n9846) );
  NOR2_X1 U7814 ( .A1(n9794), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7235) );
  NAND2_X1 U7815 ( .A1(n6636), .A2(n10216), .ZN(n7762) );
  NAND2_X1 U7816 ( .A1(n6596), .A2(n6550), .ZN(n7742) );
  AOI21_X1 U7817 ( .B1(n7224), .B2(n7228), .A(n6635), .ZN(n7222) );
  OAI21_X1 U7818 ( .B1(n12404), .B2(n7756), .A(n12411), .ZN(n7755) );
  NOR2_X1 U7819 ( .A1(n7079), .A2(n12493), .ZN(n6875) );
  INV_X1 U7820 ( .A(n7752), .ZN(n7079) );
  NAND2_X1 U7821 ( .A1(n7752), .A2(n7078), .ZN(n7077) );
  INV_X1 U7822 ( .A(n12399), .ZN(n7078) );
  NAND2_X1 U7823 ( .A1(n9623), .A2(n10046), .ZN(n10049) );
  NOR2_X1 U7824 ( .A1(n9490), .A2(n9489), .ZN(n9495) );
  INV_X1 U7825 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7570) );
  OR2_X1 U7826 ( .A1(n9451), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n9456) );
  NAND2_X1 U7827 ( .A1(n9838), .A2(n9837), .ZN(n9859) );
  INV_X1 U7828 ( .A(n9812), .ZN(n7705) );
  INV_X1 U7829 ( .A(n9644), .ZN(n7702) );
  INV_X1 U7830 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9646) );
  AND2_X1 U7831 ( .A1(n7700), .A2(n7057), .ZN(n7054) );
  NAND2_X1 U7832 ( .A1(n7700), .A2(n6563), .ZN(n7055) );
  INV_X1 U7833 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9355) );
  INV_X1 U7834 ( .A(n8665), .ZN(n7800) );
  AOI21_X1 U7835 ( .B1(n8654), .B2(n7035), .A(n7034), .ZN(n7033) );
  INV_X1 U7836 ( .A(n13639), .ZN(n7034) );
  INV_X1 U7837 ( .A(n8645), .ZN(n7035) );
  INV_X1 U7838 ( .A(n8654), .ZN(n7036) );
  NOR2_X1 U7839 ( .A1(n13877), .A2(n6639), .ZN(n7294) );
  INV_X1 U7840 ( .A(n12906), .ZN(n8030) );
  OAI22_X1 U7841 ( .A1(n12164), .A2(n12163), .B1(n12162), .B2(n12161), .ZN(
        n13999) );
  NOR2_X1 U7842 ( .A1(n8540), .A2(n7644), .ZN(n7642) );
  INV_X1 U7843 ( .A(n7646), .ZN(n7639) );
  AOI21_X1 U7844 ( .B1(n6645), .B2(n7930), .A(n7347), .ZN(n7346) );
  INV_X1 U7845 ( .A(n13899), .ZN(n7347) );
  INV_X1 U7846 ( .A(n7904), .ZN(n7349) );
  NOR2_X1 U7847 ( .A1(n7857), .A2(n14196), .ZN(n7856) );
  INV_X1 U7848 ( .A(n7858), .ZN(n7857) );
  INV_X1 U7849 ( .A(n8298), .ZN(n6735) );
  INV_X1 U7850 ( .A(n8264), .ZN(n7336) );
  NAND2_X1 U7851 ( .A1(n8020), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8240) );
  INV_X1 U7852 ( .A(n8214), .ZN(n8020) );
  NOR2_X1 U7853 ( .A1(n15650), .A2(n13777), .ZN(n7844) );
  AND2_X1 U7854 ( .A1(n8507), .A2(n8506), .ZN(n7609) );
  OR2_X1 U7855 ( .A1(n13976), .A2(n13777), .ZN(n8506) );
  INV_X1 U7856 ( .A(n7771), .ZN(n7769) );
  INV_X1 U7857 ( .A(n11538), .ZN(n7768) );
  INV_X1 U7858 ( .A(n8147), .ZN(n7770) );
  NOR2_X1 U7859 ( .A1(n11520), .A2(n7772), .ZN(n7771) );
  INV_X1 U7860 ( .A(n8106), .ZN(n7772) );
  XNOR2_X1 U7861 ( .A(n13980), .B(n13741), .ZN(n13903) );
  NAND2_X1 U7862 ( .A1(n13744), .A2(n13745), .ZN(n12003) );
  INV_X1 U7863 ( .A(n14046), .ZN(n13866) );
  INV_X1 U7864 ( .A(n8528), .ZN(n7650) );
  OAI21_X1 U7865 ( .B1(n6853), .B2(n6854), .A(n13745), .ZN(n6849) );
  NAND2_X1 U7866 ( .A1(n6852), .A2(n6851), .ZN(n6850) );
  INV_X1 U7867 ( .A(n6853), .ZN(n6852) );
  AND2_X1 U7868 ( .A1(n8472), .A2(n8471), .ZN(n8481) );
  NOR2_X1 U7869 ( .A1(n8142), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8156) );
  INV_X1 U7870 ( .A(n12719), .ZN(n8807) );
  INV_X1 U7871 ( .A(n12704), .ZN(n7003) );
  NAND2_X1 U7872 ( .A1(n7474), .A2(n12702), .ZN(n7473) );
  AND2_X1 U7873 ( .A1(n7465), .A2(n7001), .ZN(n7000) );
  NAND2_X1 U7874 ( .A1(n12710), .A2(n7466), .ZN(n7465) );
  NAND2_X1 U7875 ( .A1(n12704), .A2(n7002), .ZN(n7001) );
  INV_X1 U7876 ( .A(n12709), .ZN(n7466) );
  INV_X1 U7877 ( .A(n15227), .ZN(n8793) );
  NAND2_X1 U7878 ( .A1(n8787), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9250) );
  INV_X1 U7879 ( .A(n9248), .ZN(n8787) );
  OR2_X1 U7880 ( .A1(n9202), .A2(n14589), .ZN(n9217) );
  NOR2_X1 U7881 ( .A1(n7823), .A2(n7269), .ZN(n7268) );
  INV_X1 U7882 ( .A(n12910), .ZN(n7269) );
  OR2_X1 U7883 ( .A1(n7912), .A2(n7909), .ZN(n7905) );
  INV_X1 U7884 ( .A(n7905), .ZN(n7671) );
  NAND2_X1 U7885 ( .A1(n12749), .A2(n7670), .ZN(n7669) );
  INV_X1 U7886 ( .A(n11834), .ZN(n7670) );
  NAND2_X1 U7887 ( .A1(n11833), .A2(n11832), .ZN(n6899) );
  INV_X1 U7888 ( .A(n14646), .ZN(n12591) );
  NAND2_X1 U7889 ( .A1(n9647), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7834) );
  INV_X1 U7890 ( .A(n9589), .ZN(n7603) );
  NAND2_X1 U7891 ( .A1(n8557), .A2(n8556), .ZN(n8559) );
  OR2_X1 U7892 ( .A1(n8700), .A2(n13551), .ZN(n8558) );
  OR2_X1 U7893 ( .A1(n7994), .A2(n7581), .ZN(n7579) );
  NAND2_X1 U7894 ( .A1(n7995), .A2(n6603), .ZN(n7580) );
  NAND2_X1 U7895 ( .A1(n7593), .A2(n7981), .ZN(n8375) );
  XNOR2_X1 U7896 ( .A(n8375), .B(SI_20_), .ZN(n8374) );
  NAND2_X1 U7897 ( .A1(n7977), .A2(SI_19_), .ZN(n8348) );
  NAND2_X1 U7898 ( .A1(n7597), .A2(n7975), .ZN(n8345) );
  AOI21_X1 U7899 ( .B1(n7573), .B2(n7575), .A(n7572), .ZN(n7571) );
  INV_X1 U7900 ( .A(n7970), .ZN(n7572) );
  OR2_X1 U7901 ( .A1(n9142), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U7902 ( .A1(n6780), .A2(n7963), .ZN(n8276) );
  OAI21_X1 U7903 ( .B1(n8234), .B2(n6779), .A(n6777), .ZN(n6780) );
  INV_X1 U7904 ( .A(n6778), .ZN(n6777) );
  OAI21_X1 U7905 ( .B1(n8233), .B2(n6779), .A(n8249), .ZN(n6778) );
  XNOR2_X1 U7906 ( .A(n8276), .B(n15956), .ZN(n8279) );
  NAND2_X1 U7907 ( .A1(n6776), .A2(n7961), .ZN(n8250) );
  NAND2_X1 U7908 ( .A1(n8234), .A2(n8233), .ZN(n6776) );
  NAND2_X1 U7909 ( .A1(n7350), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6787) );
  OAI21_X1 U7910 ( .B1(n6541), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n7614), .ZN(
        n8062) );
  NAND2_X1 U7911 ( .A1(n10347), .A2(n9633), .ZN(n7614) );
  XNOR2_X1 U7912 ( .A(n15696), .B(P1_ADDR_REG_2__SCAN_IN), .ZN(n10318) );
  OAI21_X1 U7913 ( .B1(n11762), .B2(n7495), .A(n12094), .ZN(n7494) );
  OR2_X1 U7914 ( .A1(n15312), .A2(n6652), .ZN(n7501) );
  NAND2_X1 U7915 ( .A1(n6925), .A2(n15302), .ZN(n15309) );
  NAND2_X1 U7916 ( .A1(n15301), .A2(n15300), .ZN(n6925) );
  INV_X1 U7917 ( .A(n13555), .ZN(n10046) );
  NAND2_X1 U7918 ( .A1(n7526), .A2(n7529), .ZN(n7525) );
  INV_X1 U7919 ( .A(n7531), .ZN(n7526) );
  NAND2_X1 U7920 ( .A1(n7528), .A2(n7529), .ZN(n7527) );
  INV_X1 U7921 ( .A(n12992), .ZN(n7528) );
  NAND2_X1 U7922 ( .A1(n13019), .A2(n9991), .ZN(n7559) );
  INV_X1 U7923 ( .A(n9991), .ZN(n7556) );
  NOR2_X1 U7924 ( .A1(n9768), .A2(n11814), .ZN(n7565) );
  NAND2_X1 U7925 ( .A1(n7564), .A2(n6612), .ZN(n7563) );
  NAND2_X1 U7926 ( .A1(n11784), .A2(n11785), .ZN(n11899) );
  NOR2_X1 U7927 ( .A1(n9940), .A2(n7544), .ZN(n7538) );
  AOI21_X1 U7928 ( .B1(n7534), .B2(n7537), .A(n6944), .ZN(n6943) );
  INV_X1 U7929 ( .A(n13009), .ZN(n6944) );
  NAND2_X1 U7930 ( .A1(n7552), .A2(n7551), .ZN(n7550) );
  INV_X1 U7931 ( .A(n12237), .ZN(n7552) );
  INV_X1 U7932 ( .A(n13111), .ZN(n11645) );
  OR3_X1 U7933 ( .A1(n12520), .A2(n12522), .A3(n12521), .ZN(n7189) );
  AND2_X1 U7934 ( .A1(n12344), .A2(n12345), .ZN(n7928) );
  OR2_X1 U7935 ( .A1(n12478), .A2(n12477), .ZN(n12344) );
  NAND2_X1 U7936 ( .A1(n12471), .A2(n12470), .ZN(n12884) );
  INV_X1 U7937 ( .A(n12367), .ZN(n12531) );
  NAND2_X1 U7938 ( .A1(n9679), .A2(n9678), .ZN(n9680) );
  NAND2_X1 U7939 ( .A1(n9748), .A2(n11652), .ZN(n9679) );
  AND4_X1 U7940 ( .A1(n9752), .A2(n9751), .A3(n9750), .A4(n9749), .ZN(n11632)
         );
  AND2_X1 U7941 ( .A1(n9520), .A2(n10872), .ZN(n10829) );
  NAND2_X1 U7942 ( .A1(n7314), .A2(n10836), .ZN(n9520) );
  OAI21_X1 U7943 ( .B1(n10836), .B2(n7420), .A(n9401), .ZN(n10834) );
  AND2_X1 U7944 ( .A1(n9400), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7420) );
  XNOR2_X1 U7945 ( .A(n10326), .B(n6887), .ZN(n7391) );
  OR2_X1 U7946 ( .A1(n9419), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U7947 ( .A1(n6828), .A2(n6826), .ZN(n9543) );
  AOI21_X1 U7948 ( .B1(n6829), .B2(n6831), .A(n6827), .ZN(n6826) );
  NAND2_X1 U7949 ( .A1(n9533), .A2(n6829), .ZN(n6828) );
  INV_X1 U7950 ( .A(n7400), .ZN(n10916) );
  OAI211_X1 U7951 ( .C1(n7400), .C2(n7399), .A(n9425), .B(n7398), .ZN(n9429)
         );
  NAND2_X1 U7952 ( .A1(n7403), .A2(n7396), .ZN(n7398) );
  NOR2_X1 U7953 ( .A1(n7399), .A2(n10783), .ZN(n7396) );
  NAND2_X1 U7954 ( .A1(n9430), .A2(n11466), .ZN(n11468) );
  NAND2_X1 U7955 ( .A1(n9429), .A2(n10358), .ZN(n11465) );
  NAND2_X1 U7956 ( .A1(n13163), .A2(n13162), .ZN(n13182) );
  NAND2_X1 U7957 ( .A1(n13189), .A2(n13190), .ZN(n13188) );
  NAND2_X1 U7958 ( .A1(n13203), .A2(n6811), .ZN(n6812) );
  NOR2_X1 U7959 ( .A1(n10291), .A2(n6814), .ZN(n6811) );
  NAND2_X1 U7960 ( .A1(n9512), .A2(n9566), .ZN(n10289) );
  AOI21_X1 U7961 ( .B1(n13234), .B2(n13231), .A(n13230), .ZN(n13256) );
  NAND2_X1 U7962 ( .A1(n7414), .A2(n7418), .ZN(n7415) );
  NAND2_X1 U7963 ( .A1(n13308), .A2(n7709), .ZN(n7708) );
  NAND2_X1 U7964 ( .A1(n7216), .A2(n7217), .ZN(n13309) );
  OAI21_X1 U7965 ( .B1(n7191), .B2(n7102), .A(n12460), .ZN(n13311) );
  NOR2_X1 U7966 ( .A1(n10227), .A2(n7192), .ZN(n7102) );
  NAND2_X1 U7967 ( .A1(n13341), .A2(n10134), .ZN(n13320) );
  NAND2_X1 U7968 ( .A1(n10072), .A2(n10071), .ZN(n10142) );
  AOI21_X1 U7969 ( .B1(n6870), .B2(n6872), .A(n6869), .ZN(n6868) );
  NAND2_X1 U7970 ( .A1(n12349), .A2(n12350), .ZN(n13393) );
  OR2_X1 U7971 ( .A1(n9896), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9916) );
  AND2_X1 U7972 ( .A1(n7896), .A2(n12494), .ZN(n7895) );
  INV_X1 U7973 ( .A(n7235), .ZN(n9804) );
  NAND2_X1 U7974 ( .A1(n7205), .A2(n7207), .ZN(n11058) );
  NAND2_X1 U7975 ( .A1(n11058), .A2(n7898), .ZN(n11147) );
  AOI21_X1 U7976 ( .B1(n12491), .B2(n7761), .A(n7760), .ZN(n7759) );
  NAND2_X1 U7977 ( .A1(n11126), .A2(n7073), .ZN(n7758) );
  INV_X1 U7978 ( .A(n12393), .ZN(n7760) );
  NAND2_X1 U7979 ( .A1(n7231), .A2(n9665), .ZN(n9687) );
  INV_X1 U7980 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9665) );
  INV_X1 U7981 ( .A(n9685), .ZN(n7231) );
  INV_X1 U7982 ( .A(n7213), .ZN(n12491) );
  NAND2_X1 U7983 ( .A1(n11141), .A2(n12384), .ZN(n11126) );
  INV_X1 U7984 ( .A(n11121), .ZN(n12490) );
  NAND2_X1 U7985 ( .A1(n11126), .A2(n12490), .ZN(n11128) );
  INV_X1 U7986 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9664) );
  INV_X1 U7987 ( .A(n7887), .ZN(n12487) );
  INV_X1 U7988 ( .A(n12526), .ZN(n12522) );
  INV_X1 U7989 ( .A(n10097), .ZN(n11357) );
  AND2_X1 U7990 ( .A1(n10253), .A2(n10252), .ZN(n10256) );
  NAND2_X1 U7991 ( .A1(n10043), .A2(n12526), .ZN(n10232) );
  OAI21_X1 U7992 ( .B1(n13295), .B2(n10230), .A(n12471), .ZN(n12518) );
  NAND2_X1 U7993 ( .A1(n6931), .A2(n6554), .ZN(n6930) );
  INV_X1 U7994 ( .A(n13298), .ZN(n6931) );
  NAND2_X1 U7995 ( .A1(n13298), .A2(n6935), .ZN(n6934) );
  NOR2_X1 U7996 ( .A1(n12510), .A2(n6936), .ZN(n6935) );
  NAND2_X1 U7997 ( .A1(n10179), .A2(n13398), .ZN(n6936) );
  AOI21_X1 U7998 ( .B1(n12510), .B2(n6933), .A(n10202), .ZN(n6932) );
  NOR2_X1 U7999 ( .A1(n10179), .A2(n13428), .ZN(n6933) );
  AND2_X1 U8000 ( .A1(n10185), .A2(n10184), .ZN(n10192) );
  NAND2_X1 U8001 ( .A1(n10155), .A2(n10154), .ZN(n12991) );
  NAND2_X1 U8002 ( .A1(n13549), .A2(n9742), .ZN(n10155) );
  INV_X1 U8003 ( .A(n10132), .ZN(n13338) );
  NAND2_X1 U8004 ( .A1(n12539), .A2(n6551), .ZN(n13392) );
  INV_X1 U8005 ( .A(n12349), .ZN(n6872) );
  INV_X1 U8006 ( .A(n6871), .ZN(n6870) );
  OAI21_X1 U8007 ( .B1(n12445), .B2(n6872), .A(n12350), .ZN(n6871) );
  AND2_X1 U8008 ( .A1(n12348), .A2(n12347), .ZN(n13381) );
  NAND2_X1 U8009 ( .A1(n12540), .A2(n12541), .ZN(n12539) );
  NAND2_X1 U8010 ( .A1(n13422), .A2(n7198), .ZN(n7083) );
  NOR2_X1 U8011 ( .A1(n10225), .A2(n7199), .ZN(n7198) );
  INV_X1 U8012 ( .A(n12356), .ZN(n7199) );
  AND2_X1 U8013 ( .A1(n9968), .A2(n9967), .ZN(n13414) );
  AND2_X1 U8014 ( .A1(n12353), .A2(n12357), .ZN(n13411) );
  NAND2_X1 U8015 ( .A1(n6596), .A2(n12438), .ZN(n7743) );
  INV_X1 U8016 ( .A(n7742), .ZN(n7741) );
  AND2_X1 U8017 ( .A1(n12427), .A2(n12439), .ZN(n12223) );
  NAND2_X1 U8018 ( .A1(n6874), .A2(n6632), .ZN(n12197) );
  NAND2_X1 U8019 ( .A1(n11848), .A2(n7773), .ZN(n6874) );
  AND2_X1 U8020 ( .A1(n7890), .A2(n10114), .ZN(n7889) );
  INV_X1 U8021 ( .A(n7920), .ZN(n7187) );
  AND2_X1 U8022 ( .A1(n10221), .A2(n12430), .ZN(n7773) );
  AND2_X1 U8023 ( .A1(n7920), .A2(n12430), .ZN(n12502) );
  NAND2_X1 U8024 ( .A1(n11324), .A2(n12416), .ZN(n11848) );
  NAND2_X1 U8025 ( .A1(n10111), .A2(n12499), .ZN(n11321) );
  NAND2_X1 U8026 ( .A1(n6876), .A2(n12410), .ZN(n11325) );
  NAND2_X1 U8027 ( .A1(n9387), .A2(n9386), .ZN(n10081) );
  OAI22_X1 U8028 ( .A1(n12322), .A2(n12321), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n12905), .ZN(n12796) );
  NAND2_X1 U8029 ( .A1(n7044), .A2(n10152), .ZN(n10167) );
  NAND2_X1 U8030 ( .A1(n10138), .A2(n7045), .ZN(n7044) );
  NOR2_X1 U8031 ( .A1(n7917), .A2(n7046), .ZN(n7045) );
  NOR2_X1 U8032 ( .A1(n9365), .A2(n9370), .ZN(n6958) );
  INV_X1 U8033 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9375) );
  AOI21_X1 U8034 ( .B1(n7693), .B2(n7695), .A(n7692), .ZN(n7691) );
  OAI21_X1 U8035 ( .B1(n9972), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n9971), .ZN(
        n9975) );
  NAND2_X1 U8036 ( .A1(n9975), .A2(n9974), .ZN(n9993) );
  INV_X1 U8037 ( .A(n9461), .ZN(n9463) );
  AND2_X1 U8038 ( .A1(n9941), .A2(n9927), .ZN(n9928) );
  INV_X1 U8039 ( .A(n7714), .ZN(n7713) );
  OAI21_X1 U8040 ( .B1(n9820), .B2(n7715), .A(n9858), .ZN(n7714) );
  INV_X1 U8041 ( .A(n9789), .ZN(n7065) );
  INV_X1 U8042 ( .A(n7064), .ZN(n7063) );
  OAI21_X1 U8043 ( .B1(n9787), .B2(n7065), .A(n9810), .ZN(n7064) );
  XNOR2_X1 U8044 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9810) );
  XNOR2_X1 U8045 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9787) );
  NOR2_X1 U8046 ( .A1(n9645), .A2(n7704), .ZN(n7703) );
  AND2_X1 U8047 ( .A1(n10436), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9645) );
  INV_X1 U8048 ( .A(n9642), .ZN(n7704) );
  XNOR2_X1 U8049 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9681) );
  NAND2_X1 U8050 ( .A1(n9641), .A2(n9640), .ZN(n9756) );
  INV_X1 U8051 ( .A(n9487), .ZN(n9399) );
  INV_X1 U8052 ( .A(n8602), .ZN(n7041) );
  AND2_X1 U8053 ( .A1(n10803), .A2(n8602), .ZN(n7037) );
  INV_X1 U8054 ( .A(n13976), .ZN(n13776) );
  NAND2_X1 U8055 ( .A1(n7024), .A2(n6627), .ZN(n13568) );
  AND2_X1 U8056 ( .A1(n7790), .A2(n11191), .ZN(n7023) );
  INV_X1 U8057 ( .A(n11775), .ZN(n7789) );
  AND2_X1 U8058 ( .A1(n8649), .A2(n8650), .ZN(n13629) );
  AND2_X1 U8059 ( .A1(n10695), .A2(n8588), .ZN(n7012) );
  AND2_X1 U8060 ( .A1(n8601), .A2(n8596), .ZN(n7794) );
  AND2_X1 U8061 ( .A1(n8706), .A2(n8705), .ZN(n8726) );
  INV_X1 U8062 ( .A(n8646), .ZN(n13627) );
  NAND2_X1 U8063 ( .A1(n12833), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8177) );
  NOR2_X1 U8064 ( .A1(n15501), .A2(n7357), .ZN(n15500) );
  NAND2_X1 U8065 ( .A1(n15497), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U8066 ( .A1(n7379), .A2(n7376), .ZN(n7375) );
  NAND2_X1 U8067 ( .A1(n10938), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7373) );
  INV_X1 U8068 ( .A(n10936), .ZN(n7369) );
  AOI21_X1 U8069 ( .B1(n7365), .B2(n10935), .A(n6666), .ZN(n7363) );
  AND2_X1 U8070 ( .A1(n15553), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7371) );
  AND2_X1 U8071 ( .A1(n7363), .A2(n7361), .ZN(n7360) );
  INV_X1 U8072 ( .A(n15556), .ZN(n7361) );
  NAND2_X1 U8073 ( .A1(n7125), .A2(n7124), .ZN(n14011) );
  INV_X1 U8074 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7124) );
  INV_X1 U8075 ( .A(n13996), .ZN(n7125) );
  OR2_X1 U8076 ( .A1(n14322), .A2(n14065), .ZN(n12839) );
  NAND2_X1 U8077 ( .A1(n12841), .A2(n12842), .ZN(n7778) );
  AND2_X1 U8078 ( .A1(n9592), .A2(n9591), .ZN(n13874) );
  NAND2_X1 U8079 ( .A1(n7780), .A2(n7779), .ZN(n14045) );
  NOR2_X1 U8080 ( .A1(n12830), .A2(n14042), .ZN(n7779) );
  INV_X1 U8081 ( .A(n14063), .ZN(n7780) );
  NAND2_X1 U8082 ( .A1(n6788), .A2(n12830), .ZN(n14044) );
  OR2_X1 U8083 ( .A1(n14063), .A2(n14042), .ZN(n6788) );
  NAND2_X1 U8084 ( .A1(n14036), .A2(n14040), .ZN(n14038) );
  INV_X1 U8085 ( .A(n6794), .ZN(n8426) );
  OR2_X1 U8086 ( .A1(n14161), .A2(n7636), .ZN(n7635) );
  NOR2_X2 U8087 ( .A1(n14174), .A2(n14345), .ZN(n14164) );
  OAI21_X1 U8088 ( .B1(n14215), .B2(n8330), .A(n8331), .ZN(n14201) );
  NAND2_X1 U8089 ( .A1(n7328), .A2(n7329), .ZN(n6732) );
  NOR2_X1 U8090 ( .A1(n7616), .A2(n14250), .ZN(n7615) );
  INV_X1 U8091 ( .A(n7619), .ZN(n7616) );
  NAND2_X1 U8092 ( .A1(n7626), .A2(n13574), .ZN(n7625) );
  NOR2_X1 U8093 ( .A1(n8525), .A2(n7628), .ZN(n7627) );
  INV_X1 U8094 ( .A(n12084), .ZN(n7628) );
  INV_X1 U8095 ( .A(n8248), .ZN(n7338) );
  NAND2_X1 U8096 ( .A1(n12086), .A2(n8246), .ZN(n7781) );
  NAND2_X1 U8097 ( .A1(n14286), .A2(n8523), .ZN(n12090) );
  AOI21_X1 U8098 ( .B1(n7324), .B2(n7327), .A(n7321), .ZN(n7320) );
  NAND2_X1 U8099 ( .A1(n11537), .A2(n7324), .ZN(n7322) );
  AOI21_X1 U8100 ( .B1(n13914), .B2(n7326), .A(n7325), .ZN(n7324) );
  NAND2_X1 U8101 ( .A1(n11537), .A2(n11553), .ZN(n7323) );
  OR2_X2 U8102 ( .A1(n11606), .A2(n15632), .ZN(n11604) );
  NAND2_X1 U8103 ( .A1(n8424), .A2(n8423), .ZN(n14129) );
  INV_X1 U8104 ( .A(n7635), .ZN(n7634) );
  OAI21_X1 U8105 ( .B1(n14161), .B2(n7633), .A(n8535), .ZN(n7632) );
  NAND2_X1 U8106 ( .A1(n8534), .A2(n8533), .ZN(n7633) );
  OAI22_X2 U8107 ( .A1(n14183), .A2(n8532), .B1(n14440), .B2(n14153), .ZN(
        n14173) );
  OR2_X1 U8108 ( .A1(n14228), .A2(n14227), .ZN(n14230) );
  NAND2_X1 U8109 ( .A1(n12090), .A2(n12085), .ZN(n8524) );
  XNOR2_X1 U8110 ( .A(n13747), .B(n13944), .ZN(n7782) );
  INV_X1 U8111 ( .A(n15640), .ZN(n15651) );
  AND3_X1 U8112 ( .A1(n15616), .A2(n11229), .A3(n8727), .ZN(n8546) );
  NOR2_X1 U8113 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6745) );
  AND2_X1 U8114 ( .A1(n8351), .A2(n7787), .ZN(n7785) );
  NAND2_X1 U8115 ( .A1(n7145), .A2(n8188), .ZN(n8209) );
  OR2_X1 U8116 ( .A1(n9250), .A2(n14608), .ZN(n9271) );
  NAND2_X1 U8117 ( .A1(n12171), .A2(n6631), .ZN(n14489) );
  OR2_X1 U8118 ( .A1(n9213), .A2(n9214), .ZN(n7873) );
  NAND2_X1 U8119 ( .A1(n8780), .A2(n8779), .ZN(n9010) );
  AND2_X1 U8120 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n8779) );
  INV_X1 U8121 ( .A(n8990), .ZN(n8780) );
  NAND2_X1 U8122 ( .A1(n8786), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9202) );
  INV_X1 U8123 ( .A(n9200), .ZN(n8786) );
  AND2_X1 U8124 ( .A1(n7872), .A2(n7873), .ZN(n7871) );
  INV_X1 U8125 ( .A(n11000), .ZN(n8861) );
  INV_X1 U8126 ( .A(n9061), .ZN(n7876) );
  AND2_X1 U8127 ( .A1(n6678), .A2(n8981), .ZN(n7874) );
  INV_X1 U8128 ( .A(n7861), .ZN(n7860) );
  OAI21_X1 U8129 ( .B1(n6548), .B2(n9157), .A(n14547), .ZN(n7861) );
  INV_X1 U8130 ( .A(n14856), .ZN(n14614) );
  NAND2_X1 U8131 ( .A1(n9269), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n12973) );
  INV_X1 U8132 ( .A(n9271), .ZN(n9269) );
  INV_X1 U8133 ( .A(n8931), .ZN(n9311) );
  INV_X1 U8134 ( .A(n12714), .ZN(n9203) );
  NAND2_X1 U8135 ( .A1(n10588), .A2(n6737), .ZN(n14688) );
  INV_X1 U8136 ( .A(n6738), .ZN(n6737) );
  OAI21_X1 U8137 ( .B1(n14676), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6739), .ZN(
        n6738) );
  NAND2_X1 U8138 ( .A1(n10593), .A2(n10592), .ZN(n15337) );
  AND2_X1 U8139 ( .A1(n9002), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9003) );
  OR2_X1 U8140 ( .A1(n9001), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U8141 ( .A1(n10811), .A2(n10810), .ZN(n10854) );
  NAND2_X1 U8142 ( .A1(n6753), .A2(n11440), .ZN(n11441) );
  AND2_X1 U8143 ( .A1(n11339), .A2(n6754), .ZN(n6753) );
  OR2_X1 U8144 ( .A1(n14816), .A2(n15087), .ZN(n7656) );
  NAND2_X1 U8145 ( .A1(n15068), .A2(n7655), .ZN(n7654) );
  INV_X1 U8146 ( .A(n7656), .ZN(n7655) );
  NAND2_X1 U8147 ( .A1(n14856), .A2(n15029), .ZN(n12930) );
  NOR2_X1 U8148 ( .A1(n14832), .A2(n12979), .ZN(n12955) );
  NAND2_X1 U8149 ( .A1(n14854), .A2(n6592), .ZN(n7255) );
  NAND2_X1 U8150 ( .A1(n7260), .A2(n7257), .ZN(n7256) );
  INV_X1 U8151 ( .A(n14833), .ZN(n7257) );
  INV_X1 U8152 ( .A(n14853), .ZN(n14850) );
  INV_X1 U8153 ( .A(n7161), .ZN(n9233) );
  NAND2_X1 U8154 ( .A1(n14950), .A2(n7661), .ZN(n14912) );
  NAND2_X1 U8155 ( .A1(n9198), .A2(n9197), .ZN(n14955) );
  NOR2_X2 U8156 ( .A1(n14963), .A2(n15143), .ZN(n14966) );
  NAND2_X1 U8157 ( .A1(n15028), .A2(n7268), .ZN(n7262) );
  NAND2_X1 U8158 ( .A1(n7268), .A2(n15039), .ZN(n7267) );
  NOR2_X1 U8159 ( .A1(n7688), .A2(n12747), .ZN(n7687) );
  AOI21_X1 U8160 ( .B1(n6914), .B2(n15039), .A(n6644), .ZN(n6912) );
  NAND2_X1 U8161 ( .A1(n12939), .A2(n12938), .ZN(n15057) );
  NAND2_X1 U8162 ( .A1(n9023), .A2(n9022), .ZN(n12600) );
  OAI211_X1 U8163 ( .C1(n11706), .C2(n6892), .A(n6655), .B(n6891), .ZN(n11838)
         );
  OR2_X1 U8164 ( .A1(n6892), .A2(n11705), .ZN(n6891) );
  INV_X1 U8165 ( .A(n7249), .ZN(n6892) );
  NOR2_X1 U8166 ( .A1(n12756), .A2(n7250), .ZN(n7249) );
  INV_X1 U8167 ( .A(n11707), .ZN(n7250) );
  NAND2_X1 U8168 ( .A1(n11706), .A2(n11705), .ZN(n11708) );
  AND2_X1 U8169 ( .A1(n7813), .A2(n15351), .ZN(n11680) );
  INV_X1 U8170 ( .A(n12577), .ZN(n7246) );
  INV_X1 U8171 ( .A(n15237), .ZN(n11697) );
  NAND2_X1 U8172 ( .A1(n6664), .A2(n7098), .ZN(n7177) );
  NAND2_X1 U8173 ( .A1(n7100), .A2(n7099), .ZN(n7098) );
  NAND2_X1 U8174 ( .A1(n8834), .A2(n8833), .ZN(n15150) );
  NAND2_X1 U8175 ( .A1(n9164), .A2(n9163), .ZN(n15161) );
  NAND2_X1 U8176 ( .A1(n9125), .A2(n9124), .ZN(n15171) );
  INV_X1 U8177 ( .A(n15471), .ZN(n15189) );
  AND2_X1 U8178 ( .A1(n8926), .A2(n8925), .ZN(n15434) );
  AND3_X1 U8179 ( .A1(n12790), .A2(n10573), .A3(n10572), .ZN(n11664) );
  AND2_X1 U8180 ( .A1(n10574), .A2(n11665), .ZN(n10778) );
  AND2_X1 U8181 ( .A1(n8853), .A2(n10515), .ZN(n11667) );
  INV_X1 U8182 ( .A(n8759), .ZN(n8789) );
  NAND2_X1 U8183 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n7681) );
  NOR2_X1 U8184 ( .A1(n8804), .A2(n8744), .ZN(n8764) );
  NAND2_X1 U8185 ( .A1(n7988), .A2(n7987), .ZN(n8417) );
  NAND2_X1 U8186 ( .A1(n7593), .A2(n6622), .ZN(n7988) );
  XNOR2_X1 U8187 ( .A(n9303), .B(n9302), .ZN(n10468) );
  XNOR2_X1 U8188 ( .A(n8417), .B(n8393), .ZN(n8810) );
  XNOR2_X1 U8189 ( .A(n8774), .B(P1_IR_REG_21__SCAN_IN), .ZN(n11695) );
  XNOR2_X1 U8190 ( .A(n8374), .B(n8363), .ZN(n11202) );
  AND2_X1 U8191 ( .A1(n6784), .A2(n6783), .ZN(n8221) );
  OAI21_X1 U8192 ( .B1(n8148), .B2(n8141), .A(n8139), .ZN(n7605) );
  NAND2_X1 U8193 ( .A1(n7104), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10308) );
  XNOR2_X1 U8194 ( .A(n10308), .B(n7483), .ZN(n10303) );
  XNOR2_X1 U8195 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n7483) );
  AOI21_X1 U8196 ( .B1(n15244), .B2(n15243), .A(n7906), .ZN(n10388) );
  XNOR2_X1 U8197 ( .A(n10753), .B(n10385), .ZN(n10752) );
  NAND2_X1 U8198 ( .A1(n10759), .A2(n10758), .ZN(n10764) );
  NAND2_X1 U8199 ( .A1(n11754), .A2(n11753), .ZN(n11761) );
  INV_X1 U8200 ( .A(n15258), .ZN(n7507) );
  NAND2_X1 U8201 ( .A1(n15268), .A2(n15267), .ZN(n15279) );
  XNOR2_X1 U8202 ( .A(n15309), .B(n6924), .ZN(n15311) );
  INV_X1 U8203 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U8204 ( .A1(n6926), .A2(n7501), .ZN(n7113) );
  INV_X1 U8205 ( .A(n15297), .ZN(n6926) );
  OR2_X1 U8206 ( .A1(n7501), .A2(n6553), .ZN(n7115) );
  NAND2_X1 U8207 ( .A1(n7502), .A2(n6652), .ZN(n7116) );
  INV_X1 U8208 ( .A(n7503), .ZN(n7502) );
  OAI21_X1 U8209 ( .B1(n6553), .B2(n6652), .A(n15312), .ZN(n7503) );
  NAND2_X1 U8210 ( .A1(n7522), .A2(n7529), .ZN(n12993) );
  NAND2_X1 U8211 ( .A1(n10010), .A2(n10009), .ZN(n13373) );
  AND3_X1 U8212 ( .A1(n9731), .A2(n9730), .A3(n9729), .ZN(n11395) );
  NAND2_X1 U8213 ( .A1(n11412), .A2(n6950), .ZN(n11410) );
  INV_X1 U8214 ( .A(n7514), .ZN(n6950) );
  OAI21_X1 U8215 ( .B1(n9712), .B2(n10026), .A(n11411), .ZN(n7514) );
  NAND2_X1 U8216 ( .A1(n13059), .A2(n9970), .ZN(n13018) );
  OR2_X1 U8217 ( .A1(n9969), .A2(n13414), .ZN(n9970) );
  AND2_X1 U8218 ( .A1(n9825), .A2(n9824), .ZN(n12256) );
  AND2_X1 U8219 ( .A1(n10063), .A2(n13058), .ZN(n10064) );
  OR2_X1 U8220 ( .A1(n10035), .A2(n12858), .ZN(n6956) );
  OAI21_X1 U8221 ( .B1(n7237), .B2(n13081), .A(n10094), .ZN(n10095) );
  AND2_X1 U8222 ( .A1(n10018), .A2(n10017), .ZN(n13073) );
  XNOR2_X1 U8223 ( .A(n12862), .B(n9998), .ZN(n13068) );
  OR2_X1 U8224 ( .A1(n12331), .A2(n9718), .ZN(n9721) );
  INV_X1 U8225 ( .A(n13098), .ZN(n13058) );
  NAND2_X1 U8226 ( .A1(n10068), .A2(n15681), .ZN(n13096) );
  NAND2_X1 U8227 ( .A1(n10149), .A2(n10148), .ZN(n13342) );
  NAND2_X1 U8228 ( .A1(n10034), .A2(n10033), .ZN(n13369) );
  INV_X1 U8229 ( .A(n13073), .ZN(n13385) );
  NAND2_X1 U8230 ( .A1(n10005), .A2(n10004), .ZN(n13397) );
  NAND2_X1 U8231 ( .A1(n9987), .A2(n9986), .ZN(n13384) );
  INV_X1 U8232 ( .A(n13414), .ZN(n13395) );
  NAND2_X1 U8233 ( .A1(n9953), .A2(n9952), .ZN(n13101) );
  NAND2_X1 U8234 ( .A1(n9922), .A2(n9921), .ZN(n13102) );
  NAND2_X1 U8235 ( .A1(n9883), .A2(n9882), .ZN(n13103) );
  NAND2_X1 U8236 ( .A1(n12270), .A2(n9748), .ZN(n9866) );
  INV_X1 U8237 ( .A(n12266), .ZN(n13104) );
  NAND2_X1 U8238 ( .A1(n12259), .A2(n9748), .ZN(n9830) );
  NAND2_X1 U8239 ( .A1(n12245), .A2(n9748), .ZN(n9809) );
  INV_X1 U8240 ( .A(n11414), .ZN(n13115) );
  NAND4_X1 U8241 ( .A1(n9704), .A2(n9703), .A3(n9702), .A4(n9701), .ZN(n13118)
         );
  NAND2_X1 U8242 ( .A1(n13169), .A2(n6960), .ZN(n13170) );
  INV_X1 U8243 ( .A(n6812), .ZN(n10290) );
  NAND2_X1 U8244 ( .A1(n13203), .A2(n6813), .ZN(n10292) );
  AND3_X1 U8245 ( .A1(n13269), .A2(n13268), .A3(n13267), .ZN(n13270) );
  NAND2_X1 U8246 ( .A1(n6968), .A2(n6966), .ZN(n13286) );
  NAND2_X1 U8247 ( .A1(n13279), .A2(n13280), .ZN(n7316) );
  INV_X1 U8248 ( .A(n13278), .ZN(n7317) );
  AND2_X1 U8249 ( .A1(n13275), .A2(n13276), .ZN(n7319) );
  XNOR2_X1 U8250 ( .A(n7127), .B(n7126), .ZN(n9584) );
  INV_X1 U8251 ( .A(n9576), .ZN(n7126) );
  NAND2_X1 U8252 ( .A1(n7152), .A2(n7151), .ZN(n7127) );
  OAI211_X1 U8253 ( .C1(n6965), .C2(n9575), .A(n6964), .B(n6963), .ZN(n9517)
         );
  NAND2_X1 U8254 ( .A1(n6969), .A2(n6724), .ZN(n6963) );
  INV_X1 U8255 ( .A(n13242), .ZN(n13284) );
  NAND2_X1 U8256 ( .A1(n9932), .A2(n9931), .ZN(n13484) );
  NAND2_X1 U8257 ( .A1(n11146), .A2(n12403), .ZN(n7757) );
  AND3_X1 U8258 ( .A1(n9745), .A2(n9744), .A3(n9743), .ZN(n11507) );
  AND2_X1 U8259 ( .A1(n10043), .A2(n12522), .ZN(n15679) );
  NAND2_X1 U8260 ( .A1(n9676), .A2(n9675), .ZN(n11169) );
  OR2_X1 U8261 ( .A1(n15691), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n6937) );
  INV_X1 U8262 ( .A(n10192), .ZN(n10264) );
  INV_X1 U8263 ( .A(n10178), .ZN(n13497) );
  NAND2_X1 U8264 ( .A1(n9997), .A2(n9996), .ZN(n13521) );
  NAND2_X1 U8265 ( .A1(n9946), .A2(n9945), .ZN(n13535) );
  NAND2_X1 U8266 ( .A1(n15691), .A2(n13474), .ZN(n13540) );
  OR2_X1 U8267 ( .A1(n10245), .A2(n10244), .ZN(n10246) );
  NAND2_X1 U8268 ( .A1(n8566), .A2(n8460), .ZN(n14072) );
  AND2_X1 U8269 ( .A1(n7803), .A2(n13561), .ZN(n7802) );
  AND3_X1 U8270 ( .A1(n7014), .A2(n7013), .A3(n8581), .ZN(n10562) );
  NAND2_X1 U8271 ( .A1(n8308), .A2(n8307), .ZN(n14372) );
  NAND2_X1 U8272 ( .A1(n8592), .A2(n10803), .ZN(n10809) );
  AND2_X1 U8273 ( .A1(n13711), .A2(n8582), .ZN(n13712) );
  INV_X1 U8274 ( .A(n13725), .ZN(n13693) );
  INV_X1 U8275 ( .A(n13964), .ZN(n13698) );
  NAND2_X1 U8276 ( .A1(n7804), .A2(n7805), .ZN(n13707) );
  AOI211_X1 U8277 ( .C1(n13936), .C2(n13940), .A(n13941), .B(n13935), .ZN(
        n13951) );
  NOR4_X1 U8278 ( .A1(n13933), .A2(n13932), .A3(n13931), .A4(n13930), .ZN(
        n13934) );
  OR2_X1 U8279 ( .A1(n14123), .A2(n8461), .ZN(n8433) );
  NAND2_X1 U8280 ( .A1(n10708), .A2(n7378), .ZN(n7380) );
  NAND2_X1 U8281 ( .A1(n14067), .A2(n14307), .ZN(n6839) );
  OR2_X1 U8282 ( .A1(n14063), .A2(n14062), .ZN(n14067) );
  INV_X1 U8283 ( .A(n14066), .ZN(n6842) );
  AND2_X1 U8284 ( .A1(n8018), .A2(n8017), .ZN(n14082) );
  NAND2_X1 U8285 ( .A1(n7343), .A2(n12900), .ZN(n14089) );
  XNOR2_X1 U8286 ( .A(n10272), .B(n13928), .ZN(n7344) );
  INV_X1 U8287 ( .A(n14282), .ZN(n14297) );
  NAND2_X1 U8288 ( .A1(n15615), .A2(n8716), .ZN(n14290) );
  AND2_X1 U8289 ( .A1(n8702), .A2(n8701), .ZN(n14413) );
  NAND2_X1 U8290 ( .A1(n15670), .A2(n14347), .ZN(n14401) );
  OAI211_X1 U8291 ( .C1(n9603), .C2(n7584), .A(n9607), .B(n7582), .ZN(n13872)
         );
  NAND2_X1 U8292 ( .A1(n7588), .A2(n8102), .ZN(n7584) );
  NAND2_X1 U8293 ( .A1(n9603), .A2(n7583), .ZN(n7582) );
  INV_X1 U8294 ( .A(n14031), .ZN(n14411) );
  OR2_X1 U8295 ( .A1(n14089), .A2(n7341), .ZN(n7340) );
  OR2_X1 U8296 ( .A1(n14094), .A2(n7342), .ZN(n7341) );
  AND2_X1 U8297 ( .A1(n13859), .A2(n15651), .ZN(n7342) );
  NAND2_X1 U8298 ( .A1(n7643), .A2(n7641), .ZN(n10274) );
  INV_X1 U8299 ( .A(n7644), .ZN(n7641) );
  NAND2_X1 U8300 ( .A1(n7128), .A2(n7646), .ZN(n7643) );
  NAND2_X1 U8301 ( .A1(n15659), .A2(n14347), .ZN(n14461) );
  NAND2_X1 U8302 ( .A1(n8502), .A2(n8501), .ZN(n15614) );
  NOR2_X1 U8303 ( .A1(n8008), .A2(n6659), .ZN(n6856) );
  NAND2_X1 U8304 ( .A1(n12808), .A2(n7879), .ZN(n11015) );
  AND2_X1 U8305 ( .A1(n8906), .A2(n8893), .ZN(n7879) );
  INV_X1 U8306 ( .A(n11013), .ZN(n8906) );
  INV_X1 U8307 ( .A(n9328), .ZN(n7074) );
  NAND2_X1 U8308 ( .A1(n9344), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14611) );
  NAND2_X1 U8309 ( .A1(n12173), .A2(n12172), .ZN(n12171) );
  NAND2_X1 U8310 ( .A1(n9178), .A2(n9177), .ZN(n15156) );
  INV_X1 U8311 ( .A(n14600), .ZN(n14609) );
  OR2_X1 U8312 ( .A1(n6771), .A2(n7865), .ZN(n6770) );
  INV_X1 U8313 ( .A(n14607), .ZN(n7173) );
  INV_X1 U8314 ( .A(n14619), .ZN(n14621) );
  NAND2_X1 U8315 ( .A1(n7184), .A2(n7183), .ZN(n6782) );
  OR2_X1 U8316 ( .A1(n12789), .A2(n7924), .ZN(n7184) );
  INV_X1 U8317 ( .A(n12793), .ZN(n7176) );
  OR2_X1 U8318 ( .A1(n10617), .A2(n10616), .ZN(n14805) );
  INV_X1 U8319 ( .A(n12556), .ZN(n14809) );
  NAND2_X1 U8320 ( .A1(n12717), .A2(n12716), .ZN(n15064) );
  NAND2_X1 U8321 ( .A1(n12723), .A2(n12722), .ZN(n14829) );
  OAI211_X1 U8322 ( .C1(n15075), .C2(n15060), .A(n7690), .B(n6895), .ZN(n6894)
         );
  INV_X1 U8323 ( .A(n12988), .ZN(n7690) );
  NAND2_X1 U8324 ( .A1(n15073), .A2(n12989), .ZN(n6895) );
  INV_X1 U8325 ( .A(n7177), .ZN(n15075) );
  NAND2_X1 U8326 ( .A1(n15096), .A2(n15461), .ZN(n6900) );
  NAND2_X1 U8327 ( .A1(n8762), .A2(n8761), .ZN(n14860) );
  AND2_X1 U8328 ( .A1(n12950), .A2(n7307), .ZN(n7306) );
  NAND2_X1 U8329 ( .A1(n7308), .A2(n12950), .ZN(n14911) );
  INV_X1 U8330 ( .A(n14985), .ZN(n15392) );
  NAND2_X1 U8331 ( .A1(n7258), .A2(n7165), .ZN(n7164) );
  NAND2_X1 U8332 ( .A1(n6902), .A2(n6901), .ZN(n15195) );
  AND2_X1 U8333 ( .A1(n6556), .A2(n6681), .ZN(n6901) );
  NAND2_X1 U8334 ( .A1(n15096), .A2(n6903), .ZN(n6902) );
  NOR2_X1 U8335 ( .A1(n15109), .A2(n7838), .ZN(n7837) );
  INV_X1 U8336 ( .A(n14871), .ZN(n7838) );
  OAI21_X1 U8337 ( .B1(n14864), .B2(n7828), .A(n7825), .ZN(n14868) );
  AND2_X1 U8338 ( .A1(n8756), .A2(n15732), .ZN(n7878) );
  XNOR2_X1 U8339 ( .A(n6772), .B(P1_IR_REG_22__SCAN_IN), .ZN(n15237) );
  OAI21_X1 U8340 ( .B1(n8775), .B2(n6773), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6772) );
  NAND2_X1 U8341 ( .A1(n8765), .A2(n6774), .ZN(n6773) );
  AND2_X1 U8342 ( .A1(n10373), .A2(n10372), .ZN(n15244) );
  XNOR2_X1 U8343 ( .A(n10378), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15243) );
  OR2_X1 U8344 ( .A1(n10773), .A2(n10772), .ZN(n7497) );
  NAND2_X1 U8345 ( .A1(n10773), .A2(n10772), .ZN(n7498) );
  NAND2_X1 U8346 ( .A1(n15259), .A2(n15258), .ZN(n15262) );
  NAND2_X1 U8347 ( .A1(n15251), .A2(n15250), .ZN(n7505) );
  INV_X1 U8348 ( .A(n15270), .ZN(n7511) );
  NOR2_X1 U8349 ( .A1(n15284), .A2(n7179), .ZN(n7178) );
  NAND2_X1 U8350 ( .A1(n15270), .A2(n7513), .ZN(n7106) );
  AOI21_X1 U8351 ( .B1(n7510), .B2(n7512), .A(n7509), .ZN(n7508) );
  INV_X1 U8352 ( .A(n15293), .ZN(n7166) );
  NAND2_X1 U8353 ( .A1(n15298), .A2(n15297), .ZN(n15304) );
  XNOR2_X1 U8354 ( .A(n15308), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15303) );
  INV_X1 U8355 ( .A(n15311), .ZN(n15308) );
  OAI21_X1 U8356 ( .B1(n7276), .B2(n7275), .A(n7726), .ZN(n13813) );
  NAND2_X1 U8357 ( .A1(n13809), .A2(n7727), .ZN(n7726) );
  INV_X1 U8358 ( .A(n12583), .ZN(n6988) );
  NAND2_X1 U8359 ( .A1(n6857), .A2(n12375), .ZN(n12379) );
  NAND2_X1 U8360 ( .A1(n13822), .A2(n7286), .ZN(n7285) );
  AOI21_X1 U8361 ( .B1(n12595), .B2(n12594), .A(n12592), .ZN(n12593) );
  NAND2_X1 U8362 ( .A1(n12639), .A2(n12645), .ZN(n7430) );
  NAND2_X1 U8363 ( .A1(n13831), .A2(n7732), .ZN(n7731) );
  OAI21_X1 U8364 ( .B1(n12666), .B2(n6995), .A(n6991), .ZN(n6990) );
  AND2_X1 U8365 ( .A1(n12667), .A2(n6996), .ZN(n6995) );
  AND2_X1 U8366 ( .A1(n14995), .A2(n6992), .ZN(n6991) );
  MUX2_X1 U8367 ( .A(n14942), .B(n14971), .S(n12730), .Z(n12677) );
  INV_X1 U8368 ( .A(n12685), .ZN(n7010) );
  NAND2_X1 U8369 ( .A1(n13843), .A2(n7735), .ZN(n7734) );
  NOR2_X1 U8370 ( .A1(n6642), .A2(n6545), .ZN(n7279) );
  OAI21_X1 U8371 ( .B1(n6845), .B2(n6663), .A(n6844), .ZN(n12449) );
  AND2_X1 U8372 ( .A1(n12448), .A2(n12447), .ZN(n6844) );
  AOI21_X1 U8373 ( .B1(n12443), .B2(n6846), .A(n12362), .ZN(n6845) );
  NAND2_X1 U8374 ( .A1(n15646), .A2(n13941), .ZN(n13768) );
  NAND2_X1 U8375 ( .A1(n7147), .A2(n13338), .ZN(n6861) );
  INV_X1 U8376 ( .A(n12465), .ZN(n7147) );
  AND3_X1 U8377 ( .A1(n12388), .A2(n12384), .A3(n11119), .ZN(n7208) );
  INV_X1 U8378 ( .A(n13861), .ZN(n7721) );
  NOR2_X1 U8379 ( .A1(n7291), .A2(n6546), .ZN(n7289) );
  NOR2_X1 U8380 ( .A1(n6653), .A2(n7720), .ZN(n7291) );
  INV_X1 U8381 ( .A(n8317), .ZN(n7974) );
  NOR2_X1 U8382 ( .A1(n12223), .A2(n7225), .ZN(n7224) );
  INV_X1 U8383 ( .A(n10117), .ZN(n7225) );
  INV_X1 U8384 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9361) );
  OR2_X1 U8385 ( .A1(n13872), .A2(n13959), .ZN(n13893) );
  MUX2_X1 U8386 ( .A(n13961), .B(n13875), .S(n13867), .Z(n13886) );
  MUX2_X1 U8387 ( .A(n13962), .B(n14322), .S(n13867), .Z(n13883) );
  AOI21_X1 U8388 ( .B1(n7750), .B2(n13901), .A(n7749), .ZN(n7748) );
  INV_X1 U8389 ( .A(n11955), .ZN(n7750) );
  INV_X1 U8390 ( .A(n14298), .ZN(n7749) );
  NOR2_X1 U8391 ( .A1(n12699), .A2(n12701), .ZN(n7007) );
  AND2_X1 U8392 ( .A1(n7471), .A2(n7006), .ZN(n7005) );
  NAND2_X1 U8393 ( .A1(n12699), .A2(n12701), .ZN(n7006) );
  NAND2_X1 U8394 ( .A1(n12703), .A2(n7472), .ZN(n7471) );
  INV_X1 U8395 ( .A(n12702), .ZN(n7472) );
  NAND2_X1 U8396 ( .A1(n12560), .A2(n12557), .ZN(n12733) );
  NOR2_X1 U8397 ( .A1(n9105), .A2(n9104), .ZN(n7163) );
  AND2_X1 U8398 ( .A1(n14834), .A2(n12954), .ZN(n7311) );
  NOR2_X1 U8399 ( .A1(n7813), .A2(n11678), .ZN(n7810) );
  INV_X1 U8400 ( .A(n11688), .ZN(n7812) );
  AND2_X1 U8401 ( .A1(n7603), .A2(n9593), .ZN(n7600) );
  INV_X1 U8402 ( .A(n9588), .ZN(n7602) );
  INV_X1 U8403 ( .A(n7961), .ZN(n6779) );
  AND2_X1 U8404 ( .A1(n7925), .A2(n8152), .ZN(n7945) );
  NAND2_X1 U8405 ( .A1(n7305), .A2(n7947), .ZN(n8201) );
  NAND2_X1 U8406 ( .A1(n10347), .A2(n10430), .ZN(n7182) );
  INV_X1 U8407 ( .A(n8053), .ZN(n8057) );
  OAI21_X1 U8408 ( .B1(n11755), .B2(n11756), .A(n6920), .ZN(n6919) );
  NAND2_X1 U8409 ( .A1(n11757), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n6920) );
  INV_X1 U8410 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6918) );
  INV_X1 U8411 ( .A(n13507), .ZN(n12874) );
  NAND2_X1 U8412 ( .A1(n9769), .A2(n9770), .ZN(n7564) );
  NAND2_X1 U8413 ( .A1(n6834), .A2(n6833), .ZN(n12473) );
  NAND2_X1 U8414 ( .A1(n12467), .A2(n6549), .ZN(n6834) );
  AOI21_X1 U8415 ( .B1(n6549), .B2(n6837), .A(n6661), .ZN(n6833) );
  AND3_X1 U8416 ( .A1(n7395), .A2(n7394), .A3(n13122), .ZN(n7393) );
  OAI21_X1 U8417 ( .B1(n9573), .B2(P3_REG1_REG_2__SCAN_IN), .A(n7118), .ZN(
        n9522) );
  NAND2_X1 U8418 ( .A1(n9573), .A2(n6887), .ZN(n7118) );
  NOR2_X1 U8419 ( .A1(n10964), .A2(n9412), .ZN(n9417) );
  INV_X1 U8420 ( .A(n11474), .ZN(n6819) );
  INV_X1 U8421 ( .A(n11304), .ZN(n6820) );
  OAI21_X1 U8422 ( .B1(n10920), .B2(n10919), .A(n7445), .ZN(n7448) );
  NOR2_X1 U8423 ( .A1(n7446), .A2(n6629), .ZN(n7445) );
  NOR2_X1 U8424 ( .A1(n10918), .A2(n10919), .ZN(n7446) );
  NOR2_X1 U8425 ( .A1(n7413), .A2(n13166), .ZN(n7408) );
  NOR2_X1 U8426 ( .A1(n7408), .A2(n13161), .ZN(n7407) );
  NOR2_X1 U8427 ( .A1(n7463), .A2(n13221), .ZN(n7462) );
  OAI21_X1 U8428 ( .B1(n7462), .B2(n15927), .A(n7457), .ZN(n7456) );
  NAND2_X1 U8429 ( .A1(n7463), .A2(n13221), .ZN(n7457) );
  AND2_X1 U8430 ( .A1(n6812), .A2(n6580), .ZN(n9569) );
  INV_X1 U8431 ( .A(n9568), .ZN(n7313) );
  NAND2_X1 U8432 ( .A1(n13244), .A2(n6983), .ZN(n9513) );
  OR2_X1 U8433 ( .A1(n9892), .A2(n12221), .ZN(n6983) );
  INV_X1 U8434 ( .A(n13267), .ZN(n7418) );
  NAND2_X1 U8435 ( .A1(n13337), .A2(n6939), .ZN(n7216) );
  AND2_X1 U8436 ( .A1(n10150), .A2(n10133), .ZN(n6939) );
  AOI21_X1 U8437 ( .B1(n10150), .B2(n7218), .A(n6648), .ZN(n7217) );
  INV_X1 U8438 ( .A(n10134), .ZN(n7218) );
  NAND2_X1 U8439 ( .A1(n12456), .A2(n10228), .ZN(n7192) );
  OR2_X1 U8440 ( .A1(n7192), .A2(n7194), .ZN(n7167) );
  OR2_X1 U8441 ( .A1(n10142), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n10157) );
  OR2_X1 U8442 ( .A1(n13327), .A2(n12996), .ZN(n12461) );
  INV_X1 U8443 ( .A(n7232), .ZN(n10028) );
  INV_X1 U8444 ( .A(n12347), .ZN(n6869) );
  NOR2_X1 U8445 ( .A1(n6587), .A2(n7206), .ZN(n7205) );
  NOR2_X1 U8446 ( .A1(n7213), .A2(n11121), .ZN(n7073) );
  INV_X1 U8447 ( .A(n12392), .ZN(n7761) );
  INV_X1 U8448 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n7236) );
  NAND2_X1 U8449 ( .A1(n12380), .A2(n12381), .ZN(n11064) );
  NAND2_X1 U8450 ( .A1(n12377), .A2(n12376), .ZN(n11026) );
  OR2_X1 U8451 ( .A1(n12462), .A2(n12514), .ZN(n10204) );
  INV_X1 U8452 ( .A(n7224), .ZN(n7223) );
  NAND2_X1 U8453 ( .A1(n7891), .A2(n7894), .ZN(n7890) );
  INV_X1 U8454 ( .A(n10112), .ZN(n7894) );
  INV_X1 U8455 ( .A(n12498), .ZN(n12406) );
  NAND2_X1 U8456 ( .A1(n12240), .A2(n13106), .ZN(n12408) );
  INV_X1 U8457 ( .A(n7207), .ZN(n10106) );
  NAND2_X1 U8458 ( .A1(n10105), .A2(n12489), .ZN(n7209) );
  INV_X1 U8459 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n9657) );
  INV_X1 U8460 ( .A(n10137), .ZN(n7046) );
  INV_X1 U8461 ( .A(n10019), .ZN(n7692) );
  INV_X1 U8462 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7569) );
  AOI21_X1 U8463 ( .B1(n7069), .B2(n7071), .A(n7068), .ZN(n7067) );
  INV_X1 U8464 ( .A(n9957), .ZN(n7068) );
  NAND2_X1 U8465 ( .A1(n6715), .A2(n9837), .ZN(n7715) );
  INV_X1 U8466 ( .A(n7715), .ZN(n7712) );
  INV_X1 U8467 ( .A(n9821), .ZN(n9820) );
  INV_X1 U8468 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9774) );
  AND3_X1 U8469 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .A3(P2_REG3_REG_3__SCAN_IN), .ZN(n8107) );
  NAND2_X1 U8470 ( .A1(n6705), .A2(n8695), .ZN(n7808) );
  INV_X1 U8471 ( .A(n10720), .ZN(n7376) );
  NAND2_X1 U8472 ( .A1(n7355), .A2(n7354), .ZN(n7353) );
  NAND2_X1 U8473 ( .A1(n15598), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7354) );
  NAND2_X1 U8474 ( .A1(n15593), .A2(n15594), .ZN(n7355) );
  AND2_X1 U8475 ( .A1(n14128), .A2(n6679), .ZN(n14036) );
  AND2_X1 U8476 ( .A1(n12850), .A2(n8567), .ZN(n8725) );
  NOR2_X1 U8477 ( .A1(n13862), .A2(n7853), .ZN(n7852) );
  INV_X1 U8478 ( .A(n7854), .ZN(n7853) );
  NOR2_X1 U8479 ( .A1(n13859), .A2(n14109), .ZN(n7854) );
  NOR2_X1 U8480 ( .A1(n8398), .A2(n8397), .ZN(n6794) );
  OR2_X1 U8481 ( .A1(n8384), .A2(n8383), .ZN(n8398) );
  NAND2_X1 U8482 ( .A1(n6792), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8384) );
  NOR2_X1 U8483 ( .A1(n8324), .A2(n8323), .ZN(n6793) );
  NOR2_X1 U8484 ( .A1(n14365), .A2(n14368), .ZN(n7858) );
  NAND2_X1 U8485 ( .A1(n6791), .A2(n6710), .ZN(n8309) );
  OR2_X1 U8486 ( .A1(n14383), .A2(n7849), .ZN(n7848) );
  INV_X1 U8487 ( .A(n6791), .ZN(n8290) );
  OR2_X1 U8488 ( .A1(n14389), .A2(n14393), .ZN(n7849) );
  INV_X1 U8489 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8238) );
  INV_X1 U8490 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8239) );
  OR3_X1 U8491 ( .A1(n8240), .A2(n8239), .A3(n8238), .ZN(n8257) );
  INV_X1 U8492 ( .A(n11553), .ZN(n7326) );
  INV_X1 U8493 ( .A(n11864), .ZN(n7325) );
  INV_X1 U8494 ( .A(n8516), .ZN(n7613) );
  OR2_X1 U8495 ( .A1(n8195), .A2(n8019), .ZN(n8214) );
  NAND2_X1 U8496 ( .A1(n8107), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8161) );
  INV_X1 U8497 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8160) );
  AND2_X1 U8498 ( .A1(n8504), .A2(n7610), .ZN(n11078) );
  NAND2_X1 U8499 ( .A1(n13733), .A2(n11256), .ZN(n7610) );
  AOI21_X1 U8500 ( .B1(n7748), .B2(n7751), .A(n14299), .ZN(n7746) );
  INV_X1 U8501 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8473) );
  INV_X1 U8502 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8118) );
  NAND2_X1 U8503 ( .A1(n7144), .A2(n7143), .ZN(n8117) );
  INV_X1 U8504 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7143) );
  INV_X1 U8505 ( .A(n8077), .ZN(n7144) );
  NOR2_X1 U8506 ( .A1(n9179), .A2(n8785), .ZN(n7162) );
  INV_X1 U8507 ( .A(n8818), .ZN(n8809) );
  NAND2_X1 U8508 ( .A1(n14676), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6739) );
  AND2_X1 U8509 ( .A1(n7661), .A2(n7660), .ZN(n7659) );
  INV_X1 U8510 ( .A(n15111), .ZN(n7660) );
  NOR2_X1 U8511 ( .A1(n9217), .A2(n14501), .ZN(n7161) );
  NOR2_X1 U8512 ( .A1(n15121), .A2(n7662), .ZN(n7661) );
  NAND2_X1 U8513 ( .A1(n15129), .A2(n14636), .ZN(n7103) );
  NOR2_X1 U8514 ( .A1(n7817), .A2(n7264), .ZN(n7263) );
  INV_X1 U8515 ( .A(n12914), .ZN(n7264) );
  INV_X1 U8516 ( .A(n7818), .ZN(n7817) );
  AND2_X1 U8517 ( .A1(n14947), .A2(n7819), .ZN(n7818) );
  NAND2_X1 U8518 ( .A1(n14973), .A2(n12915), .ZN(n7819) );
  INV_X1 U8519 ( .A(n12915), .ZN(n7816) );
  NAND3_X1 U8520 ( .A1(n7267), .A2(n7261), .A3(n7262), .ZN(n7265) );
  AND2_X1 U8521 ( .A1(n7820), .A2(n7310), .ZN(n7261) );
  NAND2_X1 U8522 ( .A1(n12911), .A2(n12912), .ZN(n7824) );
  NAND2_X1 U8523 ( .A1(n15001), .A2(n6802), .ZN(n14963) );
  NOR2_X1 U8524 ( .A1(n15150), .A2(n15156), .ZN(n6802) );
  INV_X1 U8525 ( .A(n12940), .ZN(n6914) );
  NAND2_X1 U8526 ( .A1(n7163), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9147) );
  INV_X1 U8527 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9146) );
  OR2_X1 U8528 ( .A1(n9147), .A2(n9146), .ZN(n9166) );
  NOR2_X1 U8529 ( .A1(n7665), .A2(n15171), .ZN(n7664) );
  NOR2_X1 U8530 ( .A1(n15175), .A2(n15183), .ZN(n7666) );
  INV_X1 U8531 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9104) );
  INV_X1 U8532 ( .A(n7163), .ZN(n9127) );
  NAND2_X1 U8533 ( .A1(n11980), .A2(n14638), .ZN(n12907) );
  NAND2_X1 U8534 ( .A1(n7160), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9049) );
  INV_X1 U8535 ( .A(n9024), .ZN(n7160) );
  INV_X1 U8536 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n15783) );
  INV_X1 U8537 ( .A(n11736), .ZN(n7831) );
  NAND2_X1 U8538 ( .A1(n8781), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9024) );
  INV_X1 U8539 ( .A(n9010), .ZN(n8781) );
  INV_X1 U8540 ( .A(n12756), .ZN(n7156) );
  NOR2_X1 U8541 ( .A1(n15077), .A2(n12987), .ZN(n7099) );
  OR2_X1 U8542 ( .A1(n15129), .A2(n14636), .ZN(n14902) );
  OAI21_X1 U8543 ( .B1(n7686), .B2(n7685), .A(n12945), .ZN(n7684) );
  INV_X1 U8544 ( .A(n12942), .ZN(n7685) );
  INV_X1 U8545 ( .A(n7687), .ZN(n7686) );
  INV_X1 U8546 ( .A(n9602), .ZN(n7591) );
  NAND2_X1 U8547 ( .A1(n7998), .A2(n7997), .ZN(n8436) );
  NAND2_X1 U8548 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  INV_X1 U8549 ( .A(n7984), .ZN(n7596) );
  INV_X1 U8550 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n15704) );
  INV_X1 U8551 ( .A(n7086), .ZN(n7085) );
  OAI21_X1 U8552 ( .B1(n7571), .B2(n7090), .A(n7972), .ZN(n7086) );
  XNOR2_X1 U8553 ( .A(n7960), .B(SI_12_), .ZN(n8233) );
  NAND2_X1 U8554 ( .A1(n7952), .A2(n7955), .ZN(n6784) );
  NAND2_X1 U8555 ( .A1(n8132), .A2(n8133), .ZN(n8149) );
  AND2_X1 U8556 ( .A1(n8085), .A2(SI_3_), .ZN(n7929) );
  INV_X1 U8557 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n10320) );
  XNOR2_X1 U8558 ( .A(n10382), .B(n10974), .ZN(n10381) );
  AOI21_X1 U8559 ( .B1(n10752), .B2(n6707), .A(n6922), .ZN(n10768) );
  OAI21_X1 U8560 ( .B1(n10754), .B2(n6923), .A(n6714), .ZN(n6922) );
  OR2_X1 U8561 ( .A1(n6919), .A2(n6918), .ZN(n11764) );
  NAND2_X1 U8562 ( .A1(n6919), .A2(n6918), .ZN(n11765) );
  OAI21_X1 U8563 ( .B1(n15279), .B2(n15278), .A(n15280), .ZN(n15289) );
  INV_X1 U8564 ( .A(n7508), .ZN(n7108) );
  NAND2_X1 U8565 ( .A1(n15291), .A2(n15290), .ZN(n15301) );
  NAND2_X1 U8566 ( .A1(n15289), .A2(n15288), .ZN(n15291) );
  NOR2_X1 U8567 ( .A1(n12881), .A2(n7532), .ZN(n7531) );
  INV_X1 U8568 ( .A(n12877), .ZN(n7532) );
  AOI21_X1 U8569 ( .B1(n7548), .B2(n9836), .A(n6719), .ZN(n7546) );
  NAND2_X1 U8570 ( .A1(n6949), .A2(n9754), .ZN(n6948) );
  NAND2_X1 U8571 ( .A1(n11390), .A2(n6945), .ZN(n6949) );
  NOR2_X1 U8572 ( .A1(n11505), .A2(n6946), .ZN(n6945) );
  INV_X1 U8573 ( .A(n9739), .ZN(n6946) );
  NOR2_X1 U8574 ( .A1(n12204), .A2(n7549), .ZN(n7548) );
  INV_X1 U8575 ( .A(n9835), .ZN(n7549) );
  INV_X1 U8576 ( .A(n13093), .ZN(n13069) );
  NAND2_X1 U8577 ( .A1(n11410), .A2(n9714), .ZN(n11400) );
  NOR2_X1 U8578 ( .A1(n10213), .A2(n10061), .ZN(n10238) );
  AND2_X1 U8579 ( .A1(n6557), .A2(n6951), .ZN(n6954) );
  NAND2_X1 U8580 ( .A1(n7548), .A2(n6955), .ZN(n6951) );
  INV_X1 U8581 ( .A(n7915), .ZN(n6955) );
  AND2_X1 U8582 ( .A1(n12343), .A2(n12342), .ZN(n12477) );
  AND3_X1 U8583 ( .A1(n9851), .A2(n9850), .A3(n9849), .ZN(n12266) );
  AND4_X1 U8584 ( .A1(n9670), .A2(n9669), .A3(n9668), .A4(n9667), .ZN(n10107)
         );
  INV_X1 U8585 ( .A(n7314), .ZN(n9519) );
  NAND2_X1 U8586 ( .A1(n10829), .A2(n11180), .ZN(n10874) );
  INV_X1 U8587 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15696) );
  NAND2_X1 U8588 ( .A1(n7392), .A2(n7391), .ZN(n7395) );
  INV_X1 U8589 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10974) );
  NAND2_X1 U8590 ( .A1(n7423), .A2(n7425), .ZN(n7422) );
  NOR2_X1 U8591 ( .A1(n7423), .A2(n11218), .ZN(n7424) );
  NAND2_X1 U8592 ( .A1(n6884), .A2(n6883), .ZN(n10964) );
  OR2_X1 U8593 ( .A1(n10965), .A2(n10966), .ZN(n6883) );
  NAND2_X1 U8594 ( .A1(n6882), .A2(n6880), .ZN(n6884) );
  INV_X1 U8595 ( .A(n7393), .ZN(n6882) );
  NAND2_X1 U8596 ( .A1(n13120), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n13119) );
  NAND2_X1 U8597 ( .A1(n6803), .A2(n10871), .ZN(n13123) );
  NAND2_X1 U8598 ( .A1(n10874), .A2(n10872), .ZN(n6803) );
  AND2_X1 U8599 ( .A1(n13151), .A2(n6974), .ZN(n10846) );
  INV_X1 U8600 ( .A(n6830), .ZN(n6829) );
  OAI21_X1 U8601 ( .B1(n10960), .B2(n6831), .A(n10842), .ZN(n6830) );
  NAND2_X1 U8602 ( .A1(n10846), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n13153) );
  NAND2_X1 U8603 ( .A1(n6975), .A2(n6972), .ZN(n7452) );
  NOR2_X1 U8604 ( .A1(n13152), .A2(n9535), .ZN(n6972) );
  NAND3_X1 U8605 ( .A1(n13151), .A2(n6660), .A3(n6974), .ZN(n7451) );
  NAND2_X1 U8606 ( .A1(n10920), .A2(n10918), .ZN(n7444) );
  NAND2_X1 U8607 ( .A1(n6816), .A2(n6815), .ZN(n11477) );
  AOI21_X1 U8608 ( .B1(n6818), .B2(n11303), .A(n11473), .ZN(n6815) );
  NAND2_X1 U8609 ( .A1(n11305), .A2(n6818), .ZN(n6816) );
  AOI21_X1 U8610 ( .B1(n9556), .B2(n6820), .A(n6819), .ZN(n6818) );
  NAND2_X1 U8611 ( .A1(n6817), .A2(n9556), .ZN(n11475) );
  NAND2_X1 U8612 ( .A1(n11305), .A2(n11304), .ZN(n6817) );
  NAND2_X1 U8613 ( .A1(n6980), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n6979) );
  INV_X1 U8614 ( .A(n7447), .ZN(n6980) );
  AND2_X1 U8615 ( .A1(n7448), .A2(n10358), .ZN(n11482) );
  NAND2_X1 U8616 ( .A1(n11468), .A2(n7408), .ZN(n7410) );
  NAND2_X1 U8617 ( .A1(n11468), .A2(n7412), .ZN(n7404) );
  NAND2_X1 U8618 ( .A1(n6885), .A2(n7405), .ZN(n13189) );
  NOR2_X1 U8619 ( .A1(n7407), .A2(n7406), .ZN(n7405) );
  NAND2_X1 U8620 ( .A1(n9430), .A2(n6608), .ZN(n6885) );
  NOR2_X1 U8621 ( .A1(n7412), .A2(n7411), .ZN(n7406) );
  OR2_X1 U8622 ( .A1(n9581), .A2(n9482), .ZN(n9516) );
  AND2_X1 U8623 ( .A1(n7442), .A2(n13207), .ZN(n7441) );
  NAND2_X1 U8624 ( .A1(n7130), .A2(n13207), .ZN(n9442) );
  NAND2_X1 U8625 ( .A1(n13182), .A2(n9562), .ZN(n13201) );
  NAND4_X1 U8626 ( .A1(n7434), .A2(n7433), .A3(n7437), .A4(n7432), .ZN(n13195)
         );
  NAND2_X1 U8627 ( .A1(n7435), .A2(n7443), .ZN(n7432) );
  AND2_X1 U8628 ( .A1(n7438), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U8629 ( .A1(n7431), .A2(n7435), .ZN(n10286) );
  XNOR2_X1 U8630 ( .A(n9569), .B(n13221), .ZN(n13217) );
  NAND2_X1 U8631 ( .A1(n10289), .A2(n7462), .ZN(n7461) );
  NAND2_X1 U8632 ( .A1(n10285), .A2(n9449), .ZN(n9453) );
  NAND2_X1 U8633 ( .A1(n6984), .A2(n13238), .ZN(n13244) );
  OAI21_X1 U8634 ( .B1(n10289), .B2(n7458), .A(n7455), .ZN(n6984) );
  NOR2_X1 U8635 ( .A1(n13221), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7458) );
  INV_X1 U8636 ( .A(n7456), .ZN(n7455) );
  NAND2_X1 U8637 ( .A1(n10289), .A2(n7464), .ZN(n7454) );
  OR2_X1 U8638 ( .A1(n7460), .A2(n7459), .ZN(n13241) );
  NAND2_X1 U8639 ( .A1(n7461), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7460) );
  INV_X1 U8640 ( .A(n13239), .ZN(n7459) );
  OR2_X1 U8641 ( .A1(n9460), .A2(n13260), .ZN(n7419) );
  NAND2_X1 U8642 ( .A1(n9513), .A2(n13260), .ZN(n13282) );
  NAND2_X1 U8643 ( .A1(n6967), .A2(n6971), .ZN(n6966) );
  INV_X1 U8644 ( .A(n13282), .ZN(n6967) );
  NAND2_X1 U8645 ( .A1(n6583), .A2(n6810), .ZN(n6809) );
  NAND2_X1 U8646 ( .A1(n6808), .A2(n6585), .ZN(n6807) );
  INV_X1 U8647 ( .A(n13255), .ZN(n6808) );
  NAND2_X1 U8648 ( .A1(n13255), .A2(n6810), .ZN(n6804) );
  NAND2_X1 U8649 ( .A1(n6969), .A2(n6584), .ZN(n6968) );
  OR2_X1 U8650 ( .A1(n10171), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n10263) );
  NAND2_X1 U8651 ( .A1(n13308), .A2(n10164), .ZN(n13297) );
  NAND2_X1 U8652 ( .A1(n7232), .A2(n10027), .ZN(n10073) );
  OAI21_X1 U8653 ( .B1(n6551), .B2(n6544), .A(n6623), .ZN(n7901) );
  NAND2_X1 U8654 ( .A1(n9979), .A2(n9978), .ZN(n9999) );
  INV_X1 U8655 ( .A(n9980), .ZN(n9979) );
  OR2_X1 U8656 ( .A1(n9999), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n10011) );
  INV_X1 U8657 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7241) );
  NAND2_X1 U8658 ( .A1(n9915), .A2(n7242), .ZN(n9947) );
  AND2_X1 U8659 ( .A1(n6577), .A2(n7239), .ZN(n7238) );
  INV_X1 U8660 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7239) );
  NAND2_X1 U8661 ( .A1(n9846), .A2(n6577), .ZN(n9895) );
  NAND2_X1 U8662 ( .A1(n9846), .A2(n9845), .ZN(n9863) );
  NAND2_X1 U8663 ( .A1(n7233), .A2(n9826), .ZN(n9847) );
  INV_X1 U8664 ( .A(n9827), .ZN(n7233) );
  NAND2_X1 U8665 ( .A1(n7235), .A2(n7234), .ZN(n9827) );
  INV_X1 U8666 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U8667 ( .A1(n11056), .A2(n12399), .ZN(n11146) );
  NAND2_X1 U8668 ( .A1(n9780), .A2(n9779), .ZN(n9794) );
  INV_X1 U8669 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9779) );
  INV_X1 U8670 ( .A(n9781), .ZN(n9780) );
  NAND2_X1 U8671 ( .A1(n7230), .A2(n7229), .ZN(n9781) );
  INV_X1 U8672 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7229) );
  INV_X1 U8673 ( .A(n9687), .ZN(n7230) );
  NAND2_X1 U8674 ( .A1(n11057), .A2(n7206), .ZN(n11056) );
  OR2_X1 U8675 ( .A1(n9762), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U8676 ( .A1(n6865), .A2(n10219), .ZN(n11139) );
  AND2_X1 U8677 ( .A1(n12388), .A2(n12384), .ZN(n12489) );
  NAND2_X1 U8678 ( .A1(n11139), .A2(n12489), .ZN(n11141) );
  NAND2_X1 U8679 ( .A1(n9732), .A2(n7236), .ZN(n9760) );
  INV_X1 U8680 ( .A(n11064), .ZN(n12486) );
  INV_X1 U8681 ( .A(n11026), .ZN(n12485) );
  NAND2_X1 U8682 ( .A1(n10216), .A2(n12368), .ZN(n11037) );
  INV_X1 U8683 ( .A(n12483), .ZN(n11036) );
  INV_X1 U8684 ( .A(n11405), .ZN(n11044) );
  NAND2_X1 U8685 ( .A1(n7887), .A2(n11411), .ZN(n10100) );
  NAND2_X1 U8686 ( .A1(n12324), .A2(n12323), .ZN(n12519) );
  AND2_X1 U8687 ( .A1(n13290), .A2(n13289), .ZN(n13489) );
  NAND2_X1 U8688 ( .A1(n7193), .A2(n12456), .ZN(n13334) );
  NAND2_X1 U8689 ( .A1(n13334), .A2(n13338), .ZN(n13333) );
  AND2_X1 U8690 ( .A1(n9902), .A2(n9901), .ZN(n12275) );
  CLKBUF_X1 U8691 ( .A(n11278), .Z(n11279) );
  AND2_X1 U8692 ( .A1(n7754), .A2(n7077), .ZN(n7076) );
  NAND2_X1 U8693 ( .A1(n6875), .A2(n11057), .ZN(n6877) );
  INV_X1 U8694 ( .A(n7755), .ZN(n7754) );
  NAND2_X1 U8695 ( .A1(n12410), .A2(n12408), .ZN(n12498) );
  OAI21_X1 U8696 ( .B1(n10181), .B2(n10180), .A(n10183), .ZN(n12322) );
  NOR2_X1 U8697 ( .A1(n9652), .A2(n6824), .ZN(n6823) );
  NOR2_X1 U8698 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6824) );
  OR2_X1 U8699 ( .A1(n9483), .A2(n15811), .ZN(n6825) );
  AND2_X1 U8700 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n11613), .ZN(n7718) );
  NAND2_X1 U8701 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7719), .ZN(n7717) );
  AOI21_X1 U8702 ( .B1(n7694), .B2(n7696), .A(n6726), .ZN(n7693) );
  INV_X1 U8703 ( .A(n9974), .ZN(n7694) );
  INV_X1 U8704 ( .A(n7696), .ZN(n7695) );
  NAND2_X1 U8705 ( .A1(n7570), .A2(n9470), .ZN(n7567) );
  AND2_X1 U8706 ( .A1(n9382), .A2(n9381), .ZN(n9383) );
  AND2_X1 U8707 ( .A1(n9906), .A2(n9888), .ZN(n9889) );
  AND2_X1 U8708 ( .A1(n9886), .A2(n9872), .ZN(n9873) );
  AND2_X1 U8709 ( .A1(n9854), .A2(n9839), .ZN(n9840) );
  AOI21_X1 U8710 ( .B1(n7063), .B2(n7065), .A(n6670), .ZN(n7061) );
  NAND2_X1 U8711 ( .A1(n7716), .A2(n9820), .ZN(n9838) );
  INV_X1 U8712 ( .A(n9822), .ZN(n7716) );
  OR2_X1 U8713 ( .A1(n9423), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9426) );
  XNOR2_X1 U8714 ( .A(n9774), .B(P1_DATAO_REG_8__SCAN_IN), .ZN(n9771) );
  NAND2_X1 U8715 ( .A1(n7056), .A2(n6621), .ZN(n9773) );
  NAND2_X1 U8716 ( .A1(n9641), .A2(n7054), .ZN(n7056) );
  AOI21_X1 U8717 ( .B1(n7700), .B2(n7702), .A(n6662), .ZN(n7698) );
  INV_X1 U8718 ( .A(n9407), .ZN(n9390) );
  OR2_X1 U8719 ( .A1(n9413), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U8720 ( .A1(n9638), .A2(n9637), .ZN(n9741) );
  XNOR2_X1 U8721 ( .A(n10349), .B(P1_DATAO_REG_2__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U8722 ( .A1(n7153), .A2(n9632), .ZN(n9716) );
  OR2_X1 U8723 ( .A1(n8439), .A2(n8024), .ZN(n8459) );
  AND2_X1 U8724 ( .A1(n7805), .A2(n6682), .ZN(n7803) );
  INV_X1 U8725 ( .A(n8660), .ZN(n7801) );
  NAND2_X1 U8726 ( .A1(n7799), .A2(n7798), .ZN(n7797) );
  INV_X1 U8727 ( .A(n8673), .ZN(n7799) );
  NOR2_X1 U8728 ( .A1(n6589), .A2(n7800), .ZN(n7798) );
  NOR2_X1 U8729 ( .A1(n6591), .A2(n7031), .ZN(n7030) );
  INV_X1 U8730 ( .A(n7033), .ZN(n7031) );
  NAND2_X1 U8731 ( .A1(n7033), .A2(n7036), .ZN(n7028) );
  NAND2_X1 U8732 ( .A1(n8021), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8324) );
  INV_X1 U8733 ( .A(n8309), .ZN(n8021) );
  INV_X1 U8734 ( .A(n6793), .ZN(n8337) );
  XNOR2_X1 U8735 ( .A(n10802), .B(n8589), .ZN(n10695) );
  NAND2_X1 U8736 ( .A1(n8618), .A2(n8617), .ZN(n11383) );
  NAND2_X1 U8737 ( .A1(n13606), .A2(n8582), .ZN(n10537) );
  AOI21_X1 U8738 ( .B1(n11385), .B2(n7792), .A(n6568), .ZN(n7790) );
  INV_X1 U8739 ( .A(n7792), .ZN(n7791) );
  INV_X1 U8740 ( .A(n8123), .ZN(n8570) );
  NAND2_X1 U8741 ( .A1(n8721), .A2(n11582), .ZN(n8111) );
  NAND2_X1 U8742 ( .A1(n8721), .A2(n10694), .ZN(n8091) );
  NAND2_X1 U8743 ( .A1(n8040), .A2(n8038), .ZN(n6854) );
  NAND2_X1 U8744 ( .A1(n8039), .A2(n8037), .ZN(n6853) );
  AND2_X1 U8745 ( .A1(n8045), .A2(n8044), .ZN(n13750) );
  AND2_X1 U8746 ( .A1(n10498), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7356) );
  INV_X1 U8747 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10519) );
  INV_X1 U8748 ( .A(n10492), .ZN(n7386) );
  NAND2_X1 U8749 ( .A1(n10743), .A2(n10744), .ZN(n10940) );
  NAND2_X1 U8750 ( .A1(n11620), .A2(n11619), .ZN(n15568) );
  INV_X1 U8751 ( .A(n8252), .ZN(n7786) );
  XNOR2_X1 U8752 ( .A(n12158), .B(n12161), .ZN(n12156) );
  XNOR2_X1 U8753 ( .A(n13999), .B(n12166), .ZN(n13997) );
  XNOR2_X1 U8754 ( .A(n7353), .B(n14001), .ZN(n14009) );
  XNOR2_X1 U8755 ( .A(n7351), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14016) );
  OAI22_X1 U8756 ( .A1(n14009), .A2(n15922), .B1(n7352), .B2(n14008), .ZN(
        n7351) );
  INV_X1 U8757 ( .A(n7353), .ZN(n7352) );
  AND2_X1 U8758 ( .A1(n8565), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8722) );
  NOR2_X1 U8759 ( .A1(n14038), .A2(n13875), .ZN(n14027) );
  AND2_X1 U8760 ( .A1(n6790), .A2(n6789), .ZN(n14063) );
  AND2_X1 U8761 ( .A1(n12828), .A2(n14068), .ZN(n6789) );
  NAND2_X1 U8762 ( .A1(n14114), .A2(n12829), .ZN(n6790) );
  AOI21_X1 U8763 ( .B1(n7642), .B2(n7639), .A(n6656), .ZN(n7638) );
  INV_X1 U8764 ( .A(n7642), .ZN(n7640) );
  AND2_X1 U8765 ( .A1(n14128), .A2(n7852), .ZN(n14074) );
  NAND2_X1 U8766 ( .A1(n14128), .A2(n7854), .ZN(n10268) );
  NAND2_X1 U8767 ( .A1(n14128), .A2(n14418), .ZN(n14105) );
  NAND2_X1 U8768 ( .A1(n6794), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U8769 ( .A1(n14114), .A2(n10270), .ZN(n14121) );
  AND2_X1 U8770 ( .A1(n14126), .A2(n14423), .ZN(n14128) );
  OAI21_X1 U8771 ( .B1(n7345), .B2(n6595), .A(n6749), .ZN(n14135) );
  INV_X1 U8772 ( .A(n6750), .ZN(n6749) );
  OAI21_X1 U8773 ( .B1(n7346), .B2(n6595), .A(n8392), .ZN(n6750) );
  INV_X1 U8774 ( .A(n8533), .ZN(n7636) );
  NOR2_X1 U8775 ( .A1(n14173), .A2(n8534), .ZN(n7637) );
  NAND2_X1 U8776 ( .A1(n14242), .A2(n6560), .ZN(n14174) );
  NAND2_X1 U8777 ( .A1(n14242), .A2(n7856), .ZN(n14193) );
  NAND2_X1 U8778 ( .A1(n6793), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8357) );
  INV_X1 U8779 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n13595) );
  NAND2_X1 U8780 ( .A1(n7348), .A2(n7904), .ZN(n14151) );
  INV_X1 U8781 ( .A(n14201), .ZN(n7348) );
  NAND2_X1 U8782 ( .A1(n6736), .A2(n8316), .ZN(n14215) );
  OAI21_X1 U8783 ( .B1(n7328), .B2(n6735), .A(n6733), .ZN(n6736) );
  INV_X1 U8784 ( .A(n6734), .ZN(n6733) );
  OAI21_X1 U8785 ( .B1(n7781), .B2(n7334), .A(n7332), .ZN(n14251) );
  NOR2_X1 U8786 ( .A1(n14259), .A2(n7848), .ZN(n7846) );
  INV_X1 U8787 ( .A(n14288), .ZN(n7847) );
  NOR2_X1 U8788 ( .A1(n14288), .A2(n14393), .ZN(n12187) );
  NAND2_X1 U8789 ( .A1(n11956), .A2(n11955), .ZN(n7747) );
  OAI21_X1 U8790 ( .B1(n11535), .B2(n8517), .A(n7611), .ZN(n11953) );
  AND2_X1 U8791 ( .A1(n7612), .A2(n8521), .ZN(n7611) );
  NAND2_X1 U8792 ( .A1(n8518), .A2(n7613), .ZN(n7612) );
  NAND2_X1 U8793 ( .A1(n11527), .A2(n7844), .ZN(n11557) );
  AOI21_X1 U8794 ( .B1(n7767), .B2(n7770), .A(n13738), .ZN(n7764) );
  NAND2_X1 U8795 ( .A1(n11527), .A2(n15641), .ZN(n11543) );
  NAND2_X1 U8796 ( .A1(n7766), .A2(n8147), .ZN(n11539) );
  NAND2_X1 U8797 ( .A1(n11596), .A2(n7771), .ZN(n7766) );
  NAND2_X1 U8798 ( .A1(n11596), .A2(n8106), .ZN(n11521) );
  NAND2_X1 U8799 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8108) );
  OR2_X1 U8800 ( .A1(n11261), .A2(n13767), .ZN(n11606) );
  NAND2_X1 U8801 ( .A1(n13903), .A2(n6731), .ZN(n12002) );
  NOR2_X1 U8802 ( .A1(n8704), .A2(n8499), .ZN(n11229) );
  NOR2_X1 U8803 ( .A1(n7586), .A2(n8043), .ZN(n7583) );
  NOR2_X1 U8804 ( .A1(n7589), .A2(n7587), .ZN(n7586) );
  INV_X1 U8805 ( .A(n7590), .ZN(n7587) );
  NAND2_X1 U8806 ( .A1(n7592), .A2(n7590), .ZN(n7588) );
  NOR2_X1 U8807 ( .A1(n14103), .A2(n7647), .ZN(n7646) );
  INV_X1 U8808 ( .A(n8538), .ZN(n7647) );
  OAI22_X1 U8809 ( .A1(n7645), .A2(n14103), .B1(n14418), .B2(n14119), .ZN(
        n7644) );
  INV_X1 U8810 ( .A(n8537), .ZN(n7645) );
  AOI21_X1 U8811 ( .B1(n14227), .B2(n6552), .A(n6633), .ZN(n7649) );
  NAND2_X1 U8812 ( .A1(n11535), .A2(n8516), .ZN(n11550) );
  AOI22_X1 U8813 ( .A1(n8354), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8353), .B2(
        n10503), .ZN(n8104) );
  AND2_X1 U8814 ( .A1(n13940), .A2(n13944), .ZN(n15646) );
  INV_X1 U8815 ( .A(n15646), .ZN(n15636) );
  NOR3_X1 U8816 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .A3(
        P2_IR_REG_19__SCAN_IN), .ZN(n8007) );
  NOR2_X1 U8817 ( .A1(n8014), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n8011) );
  NOR2_X1 U8818 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7783) );
  INV_X1 U8819 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U8820 ( .A1(n7018), .A2(n7017), .ZN(n7016) );
  INV_X1 U8821 ( .A(n7783), .ZN(n7018) );
  INV_X1 U8822 ( .A(n8014), .ZN(n7017) );
  AND2_X1 U8823 ( .A1(n8481), .A2(n8483), .ZN(n8475) );
  NAND2_X1 U8824 ( .A1(n8475), .A2(n8473), .ZN(n8479) );
  XNOR2_X1 U8825 ( .A(n8484), .B(n8483), .ZN(n11490) );
  INV_X1 U8826 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U8827 ( .A1(n6855), .A2(n7787), .ZN(n8252) );
  NOR2_X1 U8828 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6758) );
  NOR2_X1 U8829 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6757) );
  INV_X1 U8830 ( .A(n8156), .ZN(n8224) );
  OR2_X1 U8831 ( .A1(n8169), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8171) );
  INV_X1 U8832 ( .A(n7145), .ZN(n8187) );
  INV_X1 U8833 ( .A(n7162), .ZN(n8837) );
  NAND2_X1 U8834 ( .A1(n7162), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9200) );
  OR2_X1 U8835 ( .A1(n9049), .A2(n15783), .ZN(n9066) );
  NAND2_X1 U8836 ( .A1(n7868), .A2(n7869), .ZN(n7867) );
  INV_X1 U8837 ( .A(n14560), .ZN(n7868) );
  NAND2_X1 U8838 ( .A1(n11015), .A2(n8909), .ZN(n11420) );
  INV_X1 U8839 ( .A(n7881), .ZN(n7880) );
  OAI21_X1 U8840 ( .B1(n7882), .B2(n14577), .A(n9212), .ZN(n7881) );
  OAI21_X1 U8841 ( .B1(n10569), .B2(P1_D_REG_1__SCAN_IN), .A(n10555), .ZN(
        n10574) );
  NAND2_X1 U8842 ( .A1(n8778), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8990) );
  NOR2_X1 U8843 ( .A1(n9245), .A2(n9244), .ZN(n7866) );
  AOI21_X1 U8844 ( .B1(n7000), .B2(n6625), .A(n6571), .ZN(n6999) );
  NOR4_X1 U8845 ( .A1(n12780), .A2(n15077), .A3(n12772), .A4(n12771), .ZN(
        n12773) );
  OR2_X1 U8846 ( .A1(n8931), .A2(n8911), .ZN(n8912) );
  INV_X1 U8847 ( .A(n6898), .ZN(n6897) );
  OAI211_X1 U8848 ( .C1(n10591), .C2(n12714), .A(n8913), .B(n8914), .ZN(n6898)
         );
  INV_X1 U8849 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14685) );
  NAND2_X1 U8850 ( .A1(n10608), .A2(n10607), .ZN(n14771) );
  NAND2_X1 U8851 ( .A1(n8803), .A2(n15704), .ZN(n7478) );
  OR2_X1 U8852 ( .A1(n9100), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U8853 ( .A1(n10469), .A2(n8832), .ZN(n10470) );
  NAND2_X1 U8854 ( .A1(n6798), .A2(n12967), .ZN(n14817) );
  NAND2_X1 U8855 ( .A1(n12981), .A2(n12983), .ZN(n12956) );
  AND2_X1 U8856 ( .A1(n9271), .A2(n8788), .ZN(n14857) );
  AND2_X1 U8857 ( .A1(n14950), .A2(n7657), .ZN(n14875) );
  NOR2_X1 U8858 ( .A1(n14879), .A2(n7658), .ZN(n7657) );
  INV_X1 U8859 ( .A(n7659), .ZN(n7658) );
  NAND2_X1 U8860 ( .A1(n7161), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9248) );
  AND2_X1 U8861 ( .A1(n14904), .A2(n14866), .ZN(n14886) );
  NAND2_X1 U8862 ( .A1(n14904), .A2(n7827), .ZN(n14884) );
  NAND2_X1 U8863 ( .A1(n15120), .A2(n12951), .ZN(n14883) );
  NAND2_X1 U8864 ( .A1(n14950), .A2(n15129), .ZN(n14928) );
  INV_X1 U8865 ( .A(n14922), .ZN(n14926) );
  NAND2_X1 U8866 ( .A1(n14902), .A2(n7103), .ZN(n14922) );
  OR2_X1 U8867 ( .A1(n14923), .A2(n14922), .ZN(n14920) );
  NAND2_X1 U8868 ( .A1(n14972), .A2(n12946), .ZN(n14924) );
  AND2_X1 U8869 ( .A1(n14966), .A2(n15135), .ZN(n14950) );
  NAND2_X1 U8870 ( .A1(n14960), .A2(n12915), .ZN(n14940) );
  NAND2_X1 U8871 ( .A1(n6562), .A2(n14961), .ZN(n14960) );
  NAND2_X1 U8872 ( .A1(n8784), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9179) );
  INV_X1 U8873 ( .A(n9166), .ZN(n8784) );
  NOR2_X1 U8874 ( .A1(n15034), .A2(n15161), .ZN(n15001) );
  NAND2_X1 U8875 ( .A1(n15001), .A2(n15007), .ZN(n15002) );
  NAND2_X1 U8876 ( .A1(n7270), .A2(n12910), .ZN(n15014) );
  NAND2_X1 U8877 ( .A1(n7272), .A2(n7271), .ZN(n7270) );
  INV_X1 U8878 ( .A(n15028), .ZN(n7272) );
  NAND2_X1 U8879 ( .A1(n12909), .A2(n12746), .ZN(n15055) );
  NAND2_X1 U8880 ( .A1(n12106), .A2(n7664), .ZN(n15049) );
  INV_X1 U8881 ( .A(n15055), .ZN(n15045) );
  NAND2_X1 U8882 ( .A1(n12106), .A2(n7666), .ZN(n15051) );
  NAND2_X1 U8883 ( .A1(n12655), .A2(n12907), .ZN(n12765) );
  INV_X1 U8884 ( .A(n12765), .ZN(n12660) );
  NAND2_X1 U8885 ( .A1(n8782), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9085) );
  INV_X1 U8886 ( .A(n9066), .ZN(n8782) );
  NAND2_X1 U8887 ( .A1(n8783), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9105) );
  INV_X1 U8888 ( .A(n9085), .ZN(n8783) );
  AND2_X1 U8889 ( .A1(n12106), .A2(n12647), .ZN(n12107) );
  AND2_X1 U8890 ( .A1(n11991), .A2(n7669), .ZN(n7668) );
  NAND2_X1 U8891 ( .A1(n7671), .A2(n12749), .ZN(n7667) );
  OR2_X1 U8892 ( .A1(n12077), .A2(n6799), .ZN(n11945) );
  OR2_X1 U8893 ( .A1(n12600), .A2(n12619), .ZN(n6799) );
  NAND2_X1 U8894 ( .A1(n12072), .A2(n12749), .ZN(n11992) );
  NAND2_X1 U8895 ( .A1(n6801), .A2(n6800), .ZN(n12077) );
  AND2_X1 U8896 ( .A1(n12601), .A2(n7651), .ZN(n6800) );
  INV_X1 U8897 ( .A(n15362), .ZN(n6801) );
  INV_X1 U8898 ( .A(n11712), .ZN(n7651) );
  NOR2_X1 U8899 ( .A1(n11712), .A2(n15362), .ZN(n11742) );
  INV_X1 U8900 ( .A(n11682), .ZN(n7673) );
  NAND2_X1 U8901 ( .A1(n7652), .A2(n15376), .ZN(n15362) );
  AND2_X1 U8902 ( .A1(n15440), .A2(n15434), .ZN(n7652) );
  NOR2_X1 U8903 ( .A1(n15375), .A2(n14572), .ZN(n15376) );
  NAND2_X1 U8904 ( .A1(n15434), .A2(n15376), .ZN(n15361) );
  XNOR2_X1 U8905 ( .A(n11674), .B(n12812), .ZN(n12753) );
  AOI21_X1 U8906 ( .B1(n9176), .B2(n14676), .A(n7832), .ZN(n8887) );
  AND2_X1 U8907 ( .A1(n12037), .A2(n15418), .ZN(n15396) );
  INV_X1 U8908 ( .A(n14816), .ZN(n15071) );
  AOI21_X1 U8909 ( .B1(n15084), .B2(n15083), .A(n15082), .ZN(n7165) );
  NOR2_X1 U8910 ( .A1(n7259), .A2(n7252), .ZN(n7251) );
  NOR2_X1 U8911 ( .A1(n7254), .A2(n6592), .ZN(n7252) );
  OR2_X1 U8912 ( .A1(n15080), .A2(n15081), .ZN(n7259) );
  XNOR2_X1 U8913 ( .A(n14817), .B(n15071), .ZN(n15073) );
  OR2_X1 U8914 ( .A1(n15461), .A2(n15468), .ZN(n6903) );
  AOI21_X1 U8915 ( .B1(n7827), .B2(n7307), .A(n7826), .ZN(n7825) );
  INV_X1 U8916 ( .A(n14867), .ZN(n7826) );
  NAND2_X1 U8917 ( .A1(n11838), .A2(n11837), .ZN(n12074) );
  NAND2_X1 U8918 ( .A1(n10575), .A2(n9331), .ZN(n15471) );
  AND2_X1 U8919 ( .A1(n11697), .A2(n12557), .ZN(n10575) );
  NAND2_X1 U8920 ( .A1(n9605), .A2(n7591), .ZN(n7590) );
  NOR2_X1 U8921 ( .A1(n9605), .A2(n7591), .ZN(n7589) );
  INV_X1 U8922 ( .A(n9605), .ZN(n7592) );
  INV_X1 U8923 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n15732) );
  INV_X1 U8924 ( .A(n8744), .ZN(n6888) );
  AND2_X1 U8925 ( .A1(n9603), .A2(n9599), .ZN(n12805) );
  XNOR2_X1 U8926 ( .A(n9594), .B(n9593), .ZN(n12904) );
  XNOR2_X1 U8927 ( .A(n8700), .B(n8699), .ZN(n12316) );
  XNOR2_X1 U8928 ( .A(n8773), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9288) );
  OAI21_X1 U8929 ( .B1(n8772), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8773) );
  AND2_X1 U8930 ( .A1(n8771), .A2(n8772), .ZN(n9285) );
  XNOR2_X1 U8931 ( .A(n8407), .B(n8406), .ZN(n11611) );
  XNOR2_X1 U8932 ( .A(n8380), .B(n8379), .ZN(n11287) );
  INV_X1 U8933 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8742) );
  INV_X1 U8934 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8741) );
  OAI21_X1 U8935 ( .B1(n8344), .B2(n7976), .A(n8346), .ZN(n8350) );
  XNOR2_X1 U8936 ( .A(n8344), .B(n8343), .ZN(n10993) );
  NAND2_X1 U8937 ( .A1(n7089), .A2(n7571), .ZN(n8300) );
  NAND2_X1 U8938 ( .A1(n8250), .A2(n7573), .ZN(n7089) );
  AND2_X1 U8939 ( .A1(n9143), .A2(n9173), .ZN(n11802) );
  XNOR2_X1 U8940 ( .A(n7135), .B(n8281), .ZN(n10704) );
  OAI22_X1 U8941 ( .A1(n8279), .A2(n8278), .B1(n8277), .B2(SI_14_), .ZN(n7135)
         );
  XNOR2_X1 U8942 ( .A(n8181), .B(n8179), .ZN(n10441) );
  OR2_X1 U8943 ( .A1(n8953), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U8944 ( .A1(n8870), .A2(n14653), .ZN(n8900) );
  XNOR2_X1 U8945 ( .A(n8087), .B(n8086), .ZN(n10363) );
  NAND2_X1 U8946 ( .A1(n10306), .A2(n10305), .ZN(n10314) );
  NAND2_X1 U8947 ( .A1(n15242), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n7486) );
  NAND2_X1 U8948 ( .A1(n7486), .A2(n7484), .ZN(n10372) );
  NOR2_X1 U8949 ( .A1(n10321), .A2(n7485), .ZN(n7484) );
  INV_X1 U8950 ( .A(n10315), .ZN(n7485) );
  XNOR2_X1 U8951 ( .A(n10381), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U8952 ( .A1(n10751), .A2(n10750), .ZN(n10756) );
  XNOR2_X1 U8953 ( .A(n10768), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n10767) );
  NAND2_X1 U8954 ( .A1(n7112), .A2(n10774), .ZN(n7111) );
  INV_X1 U8955 ( .A(n10772), .ZN(n7112) );
  NAND2_X1 U8956 ( .A1(n6917), .A2(n11765), .ZN(n12098) );
  NAND2_X1 U8957 ( .A1(n11764), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U8958 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  NAND2_X1 U8959 ( .A1(n11762), .A2(n7495), .ZN(n7490) );
  OAI21_X1 U8960 ( .B1(n15270), .B2(n7109), .A(n7107), .ZN(n15294) );
  NOR2_X1 U8961 ( .A1(n7110), .A2(n7178), .ZN(n7109) );
  AOI22_X1 U8962 ( .A1(n7110), .A2(n7108), .B1(n7178), .B2(n7510), .ZN(n7107)
         );
  AOI21_X1 U8963 ( .B1(n7508), .B2(n7179), .A(P2_ADDR_REG_15__SCAN_IN), .ZN(
        n7110) );
  AOI21_X1 U8964 ( .B1(n15311), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n15310), .ZN(
        n15321) );
  NAND2_X1 U8965 ( .A1(n7545), .A2(n7546), .ZN(n12263) );
  NAND2_X1 U8966 ( .A1(n12237), .A2(n7548), .ZN(n7545) );
  AND2_X1 U8967 ( .A1(n11901), .A2(n11898), .ZN(n7159) );
  NAND2_X1 U8968 ( .A1(n11400), .A2(n11401), .ZN(n11399) );
  NAND2_X1 U8969 ( .A1(n6942), .A2(n7534), .ZN(n13010) );
  NAND2_X1 U8970 ( .A1(n9905), .A2(n7536), .ZN(n6942) );
  OAI21_X1 U8971 ( .B1(n9905), .B2(n7535), .A(n6943), .ZN(n13008) );
  OAI21_X1 U8972 ( .B1(n12885), .B2(n7518), .A(n7517), .ZN(n7516) );
  NAND2_X1 U8973 ( .A1(n12885), .A2(n7523), .ZN(n7517) );
  AND2_X1 U8974 ( .A1(n7523), .A2(n7527), .ZN(n7518) );
  NOR2_X1 U8975 ( .A1(n12885), .A2(n7524), .ZN(n7519) );
  NAND2_X1 U8976 ( .A1(n12885), .A2(n7521), .ZN(n7520) );
  INV_X1 U8977 ( .A(n7527), .ZN(n7521) );
  NOR2_X1 U8978 ( .A1(n9713), .A2(n9711), .ZN(n11412) );
  NAND2_X1 U8979 ( .A1(n9715), .A2(n7888), .ZN(n11409) );
  OAI211_X1 U8980 ( .C1(n12331), .C2(n10353), .A(n6928), .B(n6927), .ZN(n10097) );
  OR2_X1 U8981 ( .A1(n9790), .A2(n15702), .ZN(n6928) );
  NAND2_X1 U8982 ( .A1(n9944), .A2(n9518), .ZN(n6927) );
  OAI21_X1 U8983 ( .B1(n12961), .B2(n12331), .A(n9977), .ZN(n13024) );
  AND2_X1 U8984 ( .A1(n7555), .A2(n12873), .ZN(n7554) );
  AND2_X1 U8985 ( .A1(n12872), .A2(n12871), .ZN(n12873) );
  NAND2_X1 U8986 ( .A1(n7557), .A2(n7556), .ZN(n7555) );
  INV_X1 U8987 ( .A(n7566), .ZN(n11641) );
  INV_X1 U8988 ( .A(n6948), .ZN(n11630) );
  NAND2_X1 U8989 ( .A1(n9905), .A2(n9904), .ZN(n13048) );
  AND4_X1 U8990 ( .A1(n9766), .A2(n9765), .A3(n9764), .A4(n9763), .ZN(n11657)
         );
  NAND2_X1 U8991 ( .A1(n9748), .A2(n11635), .ZN(n9764) );
  NAND2_X1 U8992 ( .A1(n11390), .A2(n9739), .ZN(n11506) );
  AOI21_X1 U8993 ( .B1(n6943), .B2(n7535), .A(n6615), .ZN(n6941) );
  NAND2_X1 U8994 ( .A1(n7550), .A2(n9835), .ZN(n12203) );
  NAND2_X1 U8995 ( .A1(n7550), .A2(n7548), .ZN(n12206) );
  NAND3_X1 U8996 ( .A1(n13396), .A2(n10090), .A3(n10238), .ZN(n13072) );
  INV_X1 U8997 ( .A(n13096), .ZN(n13081) );
  NAND2_X1 U8998 ( .A1(n7539), .A2(n7543), .ZN(n13079) );
  NAND2_X1 U8999 ( .A1(n9905), .A2(n7540), .ZN(n7539) );
  OR2_X1 U9000 ( .A1(n12533), .A2(n10091), .ZN(n13093) );
  NOR2_X1 U9001 ( .A1(n7189), .A2(n12528), .ZN(n7051) );
  NOR2_X1 U9002 ( .A1(n12518), .A2(n12517), .ZN(n12528) );
  OAI21_X1 U9003 ( .B1(n12520), .B2(n12521), .A(n6572), .ZN(n7188) );
  NOR2_X1 U9004 ( .A1(n7053), .A2(n12884), .ZN(n7052) );
  INV_X1 U9005 ( .A(n12477), .ZN(n13290) );
  NAND2_X1 U9006 ( .A1(n10163), .A2(n10162), .ZN(n13324) );
  NAND2_X1 U9007 ( .A1(n10079), .A2(n10078), .ZN(n13353) );
  NAND2_X1 U9008 ( .A1(n11907), .A2(n9748), .ZN(n9797) );
  NAND4_X1 U9009 ( .A1(n9691), .A2(n9690), .A3(n9689), .A4(n9688), .ZN(n13110)
         );
  NAND2_X1 U9010 ( .A1(n9748), .A2(n11648), .ZN(n9689) );
  NOR2_X1 U9011 ( .A1(n9680), .A2(n7919), .ZN(n7190) );
  INV_X1 U9012 ( .A(n11657), .ZN(n13112) );
  NAND2_X1 U9013 ( .A1(n9759), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9736) );
  CLKBUF_X1 U9014 ( .A(n13117), .Z(n7138) );
  AND2_X1 U9015 ( .A1(n9521), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11180) );
  OAI21_X1 U9016 ( .B1(n9573), .B2(P3_REG1_REG_0__SCAN_IN), .A(n7168), .ZN(
        n9521) );
  NAND2_X1 U9017 ( .A1(n9573), .A2(n11174), .ZN(n7168) );
  AOI21_X1 U9018 ( .B1(n9518), .B2(n11172), .A(n9499), .ZN(n10828) );
  INV_X1 U9019 ( .A(n7391), .ZN(n10870) );
  NAND2_X1 U9020 ( .A1(n9533), .A2(n10960), .ZN(n10961) );
  AOI21_X1 U9021 ( .B1(n13140), .B2(n13138), .A(n13139), .ZN(n13142) );
  INV_X1 U9022 ( .A(n7403), .ZN(n7402) );
  XNOR2_X1 U9023 ( .A(n9424), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10924) );
  NAND2_X1 U9024 ( .A1(n9548), .A2(n10791), .ZN(n10913) );
  OR2_X1 U9025 ( .A1(n9429), .A2(n10358), .ZN(n7134) );
  OR2_X1 U9026 ( .A1(n11299), .A2(n11300), .ZN(n11470) );
  NAND2_X1 U9027 ( .A1(n7409), .A2(n7410), .ZN(n13160) );
  NOR2_X1 U9028 ( .A1(n13175), .A2(n11371), .ZN(n6959) );
  INV_X1 U9029 ( .A(n9380), .ZN(n9434) );
  NAND2_X1 U9030 ( .A1(n10286), .A2(n7440), .ZN(n13197) );
  NAND2_X1 U9031 ( .A1(n13176), .A2(n7441), .ZN(n7440) );
  XNOR2_X1 U9032 ( .A(n9453), .B(n9876), .ZN(n13214) );
  NAND2_X1 U9033 ( .A1(n7710), .A2(n7707), .ZN(n13449) );
  AOI21_X1 U9034 ( .B1(n13450), .B2(n13368), .A(n6878), .ZN(n7710) );
  INV_X1 U9035 ( .A(n13314), .ZN(n6878) );
  XNOR2_X1 U9036 ( .A(n13311), .B(n13312), .ZN(n13450) );
  NAND2_X1 U9037 ( .A1(n7133), .A2(n7131), .ZN(n13452) );
  NAND2_X1 U9038 ( .A1(n13453), .A2(n13368), .ZN(n7133) );
  INV_X1 U9039 ( .A(n7132), .ZN(n7131) );
  OAI21_X1 U9040 ( .B1(n13326), .B2(n13428), .A(n13325), .ZN(n7132) );
  NAND2_X1 U9041 ( .A1(n10227), .A2(n12453), .ZN(n13349) );
  NAND2_X1 U9042 ( .A1(n7200), .A2(n12445), .ZN(n13391) );
  AND2_X1 U9043 ( .A1(n12539), .A2(n10122), .ZN(n13394) );
  NAND2_X1 U9044 ( .A1(n12277), .A2(n10118), .ZN(n13426) );
  AND2_X1 U9045 ( .A1(n9913), .A2(n9912), .ZN(n13051) );
  NAND2_X1 U9046 ( .A1(n11147), .A2(n10109), .ZN(n11249) );
  NAND2_X1 U9047 ( .A1(n11049), .A2(n12491), .ZN(n11048) );
  NAND2_X1 U9048 ( .A1(n11128), .A2(n12392), .ZN(n11049) );
  OR2_X1 U9049 ( .A1(n10262), .A2(n10261), .ZN(n13403) );
  OR2_X1 U9050 ( .A1(n11358), .A2(n10067), .ZN(n15681) );
  XNOR2_X1 U9051 ( .A(n11351), .B(n7887), .ZN(n11354) );
  INV_X1 U9052 ( .A(n13403), .ZN(n13438) );
  INV_X1 U9053 ( .A(n13482), .ZN(n13469) );
  INV_X1 U9054 ( .A(n12519), .ZN(n13494) );
  INV_X1 U9055 ( .A(n12991), .ZN(n13501) );
  AND2_X1 U9056 ( .A1(n13344), .A2(n13343), .ZN(n13506) );
  NAND2_X1 U9057 ( .A1(n13392), .A2(n10123), .ZN(n13383) );
  OR2_X1 U9058 ( .A1(n7200), .A2(n6872), .ZN(n6867) );
  INV_X1 U9059 ( .A(n13024), .ZN(n13528) );
  NAND2_X1 U9060 ( .A1(n13424), .A2(n10119), .ZN(n13412) );
  NAND2_X1 U9061 ( .A1(n13422), .A2(n12356), .ZN(n13408) );
  INV_X1 U9062 ( .A(n7737), .ZN(n13423) );
  AOI21_X1 U9063 ( .B1(n7744), .B2(n7738), .A(n7741), .ZN(n7737) );
  INV_X1 U9064 ( .A(n7743), .ZN(n7738) );
  INV_X1 U9065 ( .A(n13051), .ZN(n12288) );
  NAND2_X1 U9066 ( .A1(n9894), .A2(n9893), .ZN(n13042) );
  NAND2_X1 U9067 ( .A1(n10116), .A2(n7227), .ZN(n7226) );
  NAND2_X1 U9068 ( .A1(n9878), .A2(n9877), .ZN(n12302) );
  NAND2_X1 U9069 ( .A1(n7774), .A2(n12430), .ZN(n12141) );
  OR2_X1 U9070 ( .A1(n11848), .A2(n7187), .ZN(n7774) );
  AND2_X1 U9071 ( .A1(n9844), .A2(n9843), .ZN(n12420) );
  NAND2_X1 U9072 ( .A1(n11321), .A2(n10112), .ZN(n11849) );
  INV_X1 U9073 ( .A(n12256), .ZN(n11498) );
  AND2_X1 U9074 ( .A1(n10081), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10395) );
  INV_X1 U9075 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9651) );
  INV_X1 U9076 ( .A(n9662), .ZN(n13545) );
  XNOR2_X1 U9077 ( .A(n10167), .B(n10153), .ZN(n13549) );
  NAND2_X1 U9078 ( .A1(n6825), .A2(n6823), .ZN(n7916) );
  NAND2_X1 U9079 ( .A1(n6957), .A2(n9369), .ZN(n13555) );
  OAI21_X1 U9080 ( .B1(n9374), .B2(P3_IR_REG_25__SCAN_IN), .A(n6958), .ZN(
        n6957) );
  NOR2_X1 U9081 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n9368) );
  INV_X1 U9082 ( .A(SI_26_), .ZN(n15772) );
  XNOR2_X1 U9083 ( .A(n9376), .B(n9375), .ZN(n13559) );
  NAND2_X1 U9084 ( .A1(n9372), .A2(n9370), .ZN(n9371) );
  XNOR2_X1 U9085 ( .A(n10023), .B(n7169), .ZN(n12181) );
  XNOR2_X1 U9086 ( .A(n7719), .B(n11613), .ZN(n7169) );
  INV_X1 U9087 ( .A(SI_23_), .ZN(n11731) );
  XNOR2_X1 U9088 ( .A(n9472), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12367) );
  OAI21_X1 U9089 ( .B1(n9628), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U9090 ( .A1(n9993), .A2(n9992), .ZN(n10008) );
  INV_X1 U9091 ( .A(SI_21_), .ZN(n12960) );
  NAND2_X1 U9092 ( .A1(n9976), .A2(n9993), .ZN(n12961) );
  OR2_X1 U9093 ( .A1(n9975), .A2(n9974), .ZN(n9976) );
  INV_X1 U9094 ( .A(SI_19_), .ZN(n10798) );
  NAND2_X1 U9095 ( .A1(n9942), .A2(n9941), .ZN(n9956) );
  INV_X1 U9096 ( .A(SI_16_), .ZN(n15925) );
  INV_X1 U9097 ( .A(SI_14_), .ZN(n15956) );
  INV_X1 U9098 ( .A(SI_12_), .ZN(n10438) );
  INV_X1 U9099 ( .A(SI_11_), .ZN(n15810) );
  NAND2_X1 U9100 ( .A1(n7706), .A2(n9812), .ZN(n9816) );
  OAI21_X1 U9101 ( .B1(n9788), .B2(n7065), .A(n7063), .ZN(n7706) );
  INV_X1 U9102 ( .A(SI_10_), .ZN(n10366) );
  NAND2_X1 U9103 ( .A1(n7062), .A2(n9789), .ZN(n9811) );
  NAND2_X1 U9104 ( .A1(n9788), .A2(n9787), .ZN(n7062) );
  XNOR2_X1 U9105 ( .A(n9395), .B(n15697), .ZN(n10367) );
  NAND2_X1 U9106 ( .A1(n7699), .A2(n9644), .ZN(n9682) );
  NAND2_X1 U9107 ( .A1(n9643), .A2(n7703), .ZN(n7699) );
  NAND2_X1 U9108 ( .A1(n9643), .A2(n9642), .ZN(n9674) );
  XNOR2_X1 U9109 ( .A(n9409), .B(n9408), .ZN(n10329) );
  NAND2_X1 U9110 ( .A1(n9405), .A2(n9407), .ZN(n10337) );
  NAND2_X1 U9111 ( .A1(n9398), .A2(n9403), .ZN(n10326) );
  MUX2_X1 U9112 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9397), .S(
        P3_IR_REG_2__SCAN_IN), .Z(n9398) );
  NAND2_X1 U9113 ( .A1(n7475), .A2(n9399), .ZN(n10836) );
  INV_X1 U9114 ( .A(n7476), .ZN(n7475) );
  NAND2_X1 U9115 ( .A1(n7040), .A2(n7038), .ZN(n10983) );
  INV_X1 U9116 ( .A(n7039), .ZN(n7038) );
  OAI21_X1 U9117 ( .B1(n7794), .B2(n7041), .A(n10979), .ZN(n7039) );
  NAND2_X2 U9118 ( .A1(n8159), .A2(n8158), .ZN(n15650) );
  AND2_X1 U9119 ( .A1(n7024), .A2(n6600), .ZN(n13569) );
  NAND2_X1 U9120 ( .A1(n11383), .A2(n8619), .ZN(n11432) );
  NAND2_X1 U9121 ( .A1(n7795), .A2(n8665), .ZN(n13613) );
  NAND2_X1 U9122 ( .A1(n13638), .A2(n6589), .ZN(n7795) );
  OR2_X1 U9123 ( .A1(n8048), .A2(n7840), .ZN(n7841) );
  NAND2_X1 U9124 ( .A1(n7029), .A2(n7027), .ZN(n13619) );
  AND2_X1 U9125 ( .A1(n7796), .A2(n6699), .ZN(n7027) );
  NAND2_X1 U9126 ( .A1(n13626), .A2(n7030), .ZN(n7029) );
  AND2_X1 U9127 ( .A1(n8672), .A2(n7797), .ZN(n7796) );
  NAND2_X1 U9128 ( .A1(n13626), .A2(n8645), .ZN(n7032) );
  NAND3_X1 U9129 ( .A1(n8686), .A2(n8685), .A3(n8684), .ZN(n13645) );
  INV_X1 U9130 ( .A(n13717), .ZN(n13701) );
  NAND2_X1 U9131 ( .A1(n12131), .A2(n8634), .ZN(n12126) );
  NAND2_X1 U9132 ( .A1(n8396), .A2(n8395), .ZN(n14145) );
  NAND2_X1 U9133 ( .A1(n8228), .A2(n8227), .ZN(n14399) );
  NAND2_X1 U9134 ( .A1(n13638), .A2(n8660), .ZN(n13690) );
  NAND2_X1 U9135 ( .A1(n10809), .A2(n7794), .ZN(n10981) );
  NAND2_X1 U9136 ( .A1(n10809), .A2(n8596), .ZN(n10888) );
  NAND2_X1 U9137 ( .A1(n7606), .A2(n8102), .ZN(n8145) );
  AND2_X1 U9138 ( .A1(n8717), .A2(n14290), .ZN(n13725) );
  NAND2_X1 U9139 ( .A1(n8466), .A2(n10483), .ZN(n14116) );
  INV_X1 U9140 ( .A(n14064), .ZN(n13963) );
  NAND2_X1 U9141 ( .A1(n8415), .A2(n8414), .ZN(n13965) );
  OR2_X1 U9142 ( .A1(n14107), .A2(n8461), .ZN(n8415) );
  NAND2_X1 U9143 ( .A1(n8404), .A2(n8403), .ZN(n13967) );
  INV_X1 U9144 ( .A(n11197), .ZN(n13975) );
  OR2_X1 U9145 ( .A1(n6854), .A2(n6853), .ZN(n13981) );
  NAND2_X1 U9146 ( .A1(n15517), .A2(n15516), .ZN(n15515) );
  NAND2_X1 U9147 ( .A1(n7383), .A2(n10489), .ZN(n10529) );
  OR2_X1 U9148 ( .A1(n10708), .A2(n10526), .ZN(n7383) );
  NAND2_X1 U9149 ( .A1(n7382), .A2(n7386), .ZN(n7381) );
  INV_X1 U9150 ( .A(n7384), .ZN(n7382) );
  AOI21_X1 U9151 ( .B1(n10489), .B2(n10526), .A(n7385), .ZN(n7384) );
  INV_X1 U9152 ( .A(n10493), .ZN(n7385) );
  NAND2_X1 U9153 ( .A1(n10508), .A2(n10509), .ZN(n10729) );
  AND2_X1 U9154 ( .A1(n7380), .A2(n7377), .ZN(n10719) );
  NAND2_X1 U9155 ( .A1(n7367), .A2(n7373), .ZN(n15544) );
  NAND2_X1 U9156 ( .A1(n7369), .A2(n7368), .ZN(n7367) );
  NAND2_X1 U9157 ( .A1(n7362), .A2(n7363), .ZN(n15555) );
  AND2_X1 U9158 ( .A1(n7362), .A2(n7360), .ZN(n15554) );
  NAND2_X1 U9159 ( .A1(n10936), .A2(n7365), .ZN(n7362) );
  AND2_X1 U9160 ( .A1(n15540), .A2(n10942), .ZN(n15560) );
  INV_X1 U9161 ( .A(n7370), .ZN(n11107) );
  AOI21_X1 U9162 ( .B1(n7360), .B2(n7364), .A(n7371), .ZN(n7358) );
  INV_X1 U9163 ( .A(n7360), .ZN(n7359) );
  OR2_X1 U9164 ( .A1(n15568), .A2(n15567), .ZN(n15569) );
  NOR2_X1 U9165 ( .A1(n15571), .A2(n6703), .ZN(n12164) );
  AND2_X1 U9166 ( .A1(n15498), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15595) );
  NAND2_X1 U9167 ( .A1(n14010), .A2(n13994), .ZN(n13996) );
  INV_X1 U9168 ( .A(n15579), .ZN(n15603) );
  NAND2_X1 U9169 ( .A1(n8452), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U9170 ( .A1(n12843), .A2(n7777), .ZN(n12854) );
  AOI21_X1 U9171 ( .B1(n14045), .B2(n6601), .A(n7778), .ZN(n7777) );
  OAI21_X1 U9172 ( .B1(n8467), .B2(n14217), .A(n13704), .ZN(n14085) );
  NAND2_X1 U9173 ( .A1(n6732), .A2(n8298), .ZN(n14226) );
  NAND2_X1 U9174 ( .A1(n7617), .A2(n7619), .ZN(n14249) );
  NAND2_X1 U9175 ( .A1(n7624), .A2(n7625), .ZN(n14278) );
  NAND2_X1 U9176 ( .A1(n8524), .A2(n7627), .ZN(n7624) );
  NAND2_X1 U9177 ( .A1(n7337), .A2(n8264), .ZN(n14266) );
  NAND2_X1 U9178 ( .A1(n7781), .A2(n6593), .ZN(n7337) );
  NAND2_X1 U9179 ( .A1(n7781), .A2(n8248), .ZN(n12184) );
  NOR2_X1 U9180 ( .A1(n12854), .A2(n7775), .ZN(n12846) );
  OR2_X1 U9181 ( .A1(n12853), .A2(n7776), .ZN(n7775) );
  AND2_X1 U9182 ( .A1(n13875), .A2(n15651), .ZN(n7776) );
  XOR2_X1 U9183 ( .A(n13931), .B(n12822), .Z(n12857) );
  AOI21_X1 U9184 ( .B1(n14035), .B2(n12830), .A(n7908), .ZN(n12822) );
  NOR2_X1 U9185 ( .A1(n14325), .A2(n14324), .ZN(n14326) );
  OR2_X1 U9186 ( .A1(n14323), .A2(n7907), .ZN(n14324) );
  NAND2_X1 U9187 ( .A1(n6839), .A2(n6838), .ZN(n14415) );
  AND2_X1 U9188 ( .A1(n14328), .A2(n6842), .ZN(n6838) );
  NOR2_X1 U9189 ( .A1(n14085), .A2(n8470), .ZN(n8547) );
  NAND2_X1 U9190 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  NAND2_X1 U9191 ( .A1(n13862), .A2(n15651), .ZN(n8468) );
  INV_X1 U9192 ( .A(n14084), .ZN(n8469) );
  AOI21_X1 U9193 ( .B1(n7128), .B2(n8538), .A(n8537), .ZN(n14104) );
  INV_X1 U9194 ( .A(n14129), .ZN(n14423) );
  INV_X1 U9195 ( .A(n14145), .ZN(n14428) );
  INV_X1 U9196 ( .A(n7629), .ZN(n14140) );
  AOI21_X1 U9197 ( .B1(n14173), .B2(n7634), .A(n7632), .ZN(n7629) );
  NAND2_X1 U9198 ( .A1(n14230), .A2(n8528), .ZN(n14213) );
  NAND2_X1 U9199 ( .A1(n8524), .A2(n12084), .ZN(n12183) );
  AND2_X1 U9200 ( .A1(n8730), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15615) );
  INV_X1 U9201 ( .A(n8029), .ZN(n12807) );
  INV_X1 U9202 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12905) );
  NAND2_X1 U9203 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), 
        .ZN(n6747) );
  NOR2_X1 U9204 ( .A1(n6746), .A2(n6745), .ZN(n6744) );
  INV_X1 U9205 ( .A(n8027), .ZN(n6748) );
  INV_X1 U9206 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14479) );
  XNOR2_X1 U9207 ( .A(n8474), .B(P2_IR_REG_26__SCAN_IN), .ZN(n14476) );
  OAI21_X1 U9208 ( .B1(n8479), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8474) );
  INV_X1 U9209 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11770) );
  INV_X1 U9210 ( .A(n14017), .ZN(n11528) );
  INV_X1 U9211 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10701) );
  INV_X1 U9212 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10565) );
  INV_X1 U9213 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10736) );
  INV_X1 U9214 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10477) );
  INV_X1 U9215 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10452) );
  XNOR2_X1 U9216 ( .A(n8210), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15553) );
  INV_X1 U9217 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10436) );
  INV_X1 U9218 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10430) );
  INV_X1 U9219 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9633) );
  INV_X1 U9220 ( .A(n15030), .ZN(n14541) );
  NAND2_X1 U9221 ( .A1(n12171), .A2(n9099), .ZN(n14491) );
  AND2_X1 U9222 ( .A1(n8817), .A2(n8816), .ZN(n14944) );
  NAND2_X1 U9223 ( .A1(n14586), .A2(n7873), .ZN(n14499) );
  NAND2_X1 U9224 ( .A1(n12808), .A2(n8893), .ZN(n11014) );
  NAND2_X1 U9225 ( .A1(n11377), .A2(n8981), .ZN(n11886) );
  NAND2_X1 U9226 ( .A1(n10998), .A2(n8862), .ZN(n11008) );
  INV_X1 U9227 ( .A(n14637), .ZN(n14942) );
  OR2_X1 U9228 ( .A1(n14584), .A2(n7882), .ZN(n14515) );
  NOR2_X1 U9229 ( .A1(n14584), .A2(n7883), .ZN(n14516) );
  NAND2_X1 U9230 ( .A1(n7094), .A2(n9062), .ZN(n12029) );
  NAND2_X1 U9231 ( .A1(n12029), .A2(n12028), .ZN(n12027) );
  OAI21_X1 U9232 ( .B1(n14586), .B2(n7867), .A(n7865), .ZN(n14523) );
  OAI21_X1 U9233 ( .B1(n14535), .B2(n6548), .A(n7860), .ZN(n14550) );
  NAND2_X1 U9234 ( .A1(n7864), .A2(n7869), .ZN(n14559) );
  NAND2_X1 U9235 ( .A1(n14586), .A2(n7871), .ZN(n7864) );
  AND2_X1 U9236 ( .A1(n14578), .A2(n14577), .ZN(n14584) );
  NAND2_X1 U9237 ( .A1(n8821), .A2(n8820), .ZN(n15143) );
  NAND2_X1 U9238 ( .A1(n6766), .A2(n7091), .ZN(n12173) );
  INV_X1 U9239 ( .A(n7092), .ZN(n7091) );
  OAI21_X1 U9240 ( .B1(n9062), .B2(n7093), .A(n9080), .ZN(n7092) );
  AND2_X1 U9241 ( .A1(n14571), .A2(n15031), .ZN(n14591) );
  OAI21_X1 U9242 ( .B1(n14578), .B2(n7882), .A(n7880), .ZN(n14587) );
  INV_X1 U9243 ( .A(n7877), .ZN(n12017) );
  NAND2_X1 U9244 ( .A1(n6762), .A2(n8882), .ZN(n12809) );
  AOI21_X1 U9245 ( .B1(n7860), .B2(n6548), .A(n6611), .ZN(n7859) );
  NAND2_X1 U9246 ( .A1(n14535), .A2(n7860), .ZN(n6767) );
  INV_X1 U9247 ( .A(n8909), .ZN(n6769) );
  NAND2_X1 U9248 ( .A1(n11271), .A2(n11273), .ZN(n11272) );
  INV_X1 U9249 ( .A(n14611), .ZN(n14630) );
  INV_X1 U9250 ( .A(n14617), .ZN(n14633) );
  NAND2_X1 U9251 ( .A1(n9342), .A2(n9341), .ZN(n14635) );
  OR2_X1 U9252 ( .A1(n14844), .A2(n9273), .ZN(n9278) );
  NAND2_X1 U9253 ( .A1(n9224), .A2(n9223), .ZN(n14930) );
  INV_X1 U9254 ( .A(n14944), .ZN(n14636) );
  NAND2_X1 U9255 ( .A1(n9208), .A2(n9207), .ZN(n14964) );
  INV_X1 U9256 ( .A(n12581), .ZN(n14648) );
  NAND4_X1 U9257 ( .A1(n8899), .A2(n8898), .A3(n8897), .A4(n8896), .ZN(n14649)
         );
  CLKBUF_X2 U9258 ( .A(P1_U4016), .Z(n14666) );
  INV_X1 U9259 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7104) );
  NAND2_X1 U9260 ( .A1(n14688), .A2(n14687), .ZN(n10589) );
  NAND2_X1 U9261 ( .A1(n10599), .A2(n10598), .ZN(n14732) );
  NAND2_X1 U9262 ( .A1(n10603), .A2(n10602), .ZN(n14755) );
  AND2_X1 U9263 ( .A1(n9006), .A2(n9020), .ZN(n10663) );
  NAND2_X1 U9264 ( .A1(n14773), .A2(n10612), .ZN(n10615) );
  OR2_X1 U9265 ( .A1(n10854), .A2(n10812), .ZN(n10856) );
  NAND2_X1 U9266 ( .A1(n11440), .A2(n11339), .ZN(n11340) );
  NAND2_X1 U9267 ( .A1(n11441), .A2(n11440), .ZN(n11444) );
  NAND2_X1 U9268 ( .A1(n7142), .A2(n7141), .ZN(n11799) );
  INV_X1 U9269 ( .A(n11443), .ZN(n7141) );
  INV_X1 U9270 ( .A(n11444), .ZN(n7142) );
  XNOR2_X1 U9271 ( .A(n14799), .B(n14787), .ZN(n14797) );
  AND2_X1 U9272 ( .A1(n10650), .A2(n15230), .ZN(n15332) );
  NAND2_X1 U9273 ( .A1(n14819), .A2(n15377), .ZN(n15065) );
  OAI21_X1 U9274 ( .B1(n14841), .B2(n7654), .A(n14818), .ZN(n7653) );
  NOR2_X1 U9275 ( .A1(n14841), .A2(n7656), .ZN(n14826) );
  OR2_X1 U9276 ( .A1(n14841), .A2(n7654), .ZN(n14825) );
  NAND2_X1 U9277 ( .A1(n7255), .A2(n7256), .ZN(n14836) );
  NAND2_X1 U9278 ( .A1(n6667), .A2(n7260), .ZN(n6906) );
  NAND2_X1 U9279 ( .A1(n7911), .A2(n12953), .ZN(n14851) );
  NAND2_X1 U9280 ( .A1(n6671), .A2(n14880), .ZN(n15105) );
  NAND2_X1 U9281 ( .A1(n7266), .A2(n7267), .ZN(n14982) );
  AND2_X1 U9282 ( .A1(n7262), .A2(n7820), .ZN(n7266) );
  NAND2_X1 U9283 ( .A1(n7689), .A2(n7687), .ZN(n14979) );
  NAND2_X1 U9284 ( .A1(n15057), .A2(n12940), .ZN(n15040) );
  NAND2_X1 U9285 ( .A1(n11708), .A2(n7249), .ZN(n11737) );
  NAND2_X1 U9286 ( .A1(n11708), .A2(n11707), .ZN(n11735) );
  NAND2_X1 U9287 ( .A1(n11683), .A2(n11682), .ZN(n11704) );
  NAND2_X1 U9288 ( .A1(n7814), .A2(n11688), .ZN(n15353) );
  OR2_X1 U9289 ( .A1(n15405), .A2(n11698), .ZN(n15394) );
  NAND2_X1 U9290 ( .A1(n11667), .A2(n11666), .ZN(n14985) );
  INV_X1 U9291 ( .A(n15060), .ZN(n15381) );
  INV_X1 U9292 ( .A(n15394), .ZN(n14954) );
  OR2_X1 U9293 ( .A1(n15126), .A2(n15125), .ZN(n15203) );
  NAND2_X1 U9294 ( .A1(n11667), .A2(n10569), .ZN(n15407) );
  OAI211_X1 U9295 ( .C1(n9603), .C2(n7592), .A(n7590), .B(n7585), .ZN(n12715)
         );
  NAND2_X1 U9296 ( .A1(n9603), .A2(n7589), .ZN(n7585) );
  NOR2_X1 U9297 ( .A1(n7679), .A2(n7678), .ZN(n7677) );
  NOR2_X1 U9298 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n7678) );
  NAND2_X1 U9299 ( .A1(n8759), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6795) );
  INV_X1 U9300 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11774) );
  INV_X1 U9301 ( .A(n9284), .ZN(n11772) );
  INV_X1 U9302 ( .A(n9285), .ZN(n11612) );
  XNOR2_X1 U9303 ( .A(n8422), .B(n8421), .ZN(n11494) );
  XNOR2_X1 U9304 ( .A(n7084), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15238) );
  NAND2_X1 U9305 ( .A1(n8810), .A2(n10425), .ZN(n7084) );
  INV_X1 U9306 ( .A(n11695), .ZN(n12557) );
  INV_X1 U9307 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11203) );
  INV_X1 U9308 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11158) );
  INV_X1 U9309 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10994) );
  INV_X1 U9310 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10558) );
  INV_X1 U9311 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n15737) );
  INV_X1 U9312 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10656) );
  INV_X1 U9313 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10465) );
  INV_X1 U9314 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n15797) );
  INV_X1 U9315 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10448) );
  INV_X1 U9316 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10457) );
  INV_X1 U9317 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10371) );
  INV_X1 U9318 ( .A(n7606), .ZN(n10437) );
  XNOR2_X1 U9319 ( .A(n8871), .B(n8870), .ZN(n14656) );
  XNOR2_X1 U9320 ( .A(n10303), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n15240) );
  XNOR2_X1 U9321 ( .A(n10314), .B(n10312), .ZN(n15242) );
  NAND2_X1 U9322 ( .A1(n6602), .A2(n7150), .ZN(n10373) );
  NAND2_X1 U9323 ( .A1(n7487), .A2(n10386), .ZN(n7105) );
  NAND3_X1 U9324 ( .A1(n7105), .A2(n10750), .A3(n10389), .ZN(n10751) );
  NAND2_X1 U9325 ( .A1(n10388), .A2(n10387), .ZN(n10750) );
  XNOR2_X1 U9326 ( .A(n10756), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n15246) );
  NAND2_X1 U9327 ( .A1(n6921), .A2(n10754), .ZN(n10762) );
  NAND2_X1 U9328 ( .A1(n10752), .A2(n14700), .ZN(n6921) );
  XNOR2_X1 U9329 ( .A(n10764), .B(n10760), .ZN(n15248) );
  XNOR2_X1 U9330 ( .A(n11750), .B(n11751), .ZN(n11749) );
  XNOR2_X1 U9331 ( .A(n11761), .B(n11759), .ZN(n15249) );
  NAND2_X1 U9332 ( .A1(n11762), .A2(n11763), .ZN(n7496) );
  NAND2_X1 U9333 ( .A1(n15249), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n11763) );
  INV_X1 U9334 ( .A(n7490), .ZN(n7493) );
  OAI211_X1 U9335 ( .C1(n12101), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n15252), .B(
        n6569), .ZN(n15261) );
  NAND2_X1 U9336 ( .A1(n12102), .A2(n15250), .ZN(n7506) );
  AND2_X1 U9337 ( .A1(n7116), .A2(n7115), .ZN(n7500) );
  NOR2_X1 U9338 ( .A1(n15313), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15317) );
  OAI21_X1 U9339 ( .B1(n6567), .B2(n6657), .A(n7158), .ZN(P3_U3169) );
  INV_X1 U9340 ( .A(n10095), .ZN(n7158) );
  OR4_X1 U9341 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        P3_U3196) );
  OAI21_X1 U9342 ( .B1(n13274), .B2(n7319), .A(n13248), .ZN(n7318) );
  OAI21_X1 U9343 ( .B1(n13270), .B2(n13271), .A(n13209), .ZN(n7315) );
  AOI21_X1 U9344 ( .B1(n9584), .B2(n13248), .A(n9583), .ZN(n9585) );
  INV_X1 U9345 ( .A(n7121), .ZN(n7120) );
  OAI22_X1 U9346 ( .A1(n13497), .A2(n13482), .B1(n13486), .B2(n13448), .ZN(
        n7121) );
  NAND2_X1 U9347 ( .A1(n6938), .A2(n6937), .ZN(n10250) );
  INV_X1 U9348 ( .A(n7123), .ZN(n7122) );
  OAI22_X1 U9349 ( .A1(n13497), .A2(n13536), .B1(n15691), .B2(n13496), .ZN(
        n7123) );
  INV_X1 U9350 ( .A(n8740), .ZN(n7148) );
  AOI211_X1 U9351 ( .C1(n13707), .C2(n13711), .A(n13706), .B(n13705), .ZN(
        n13708) );
  AND2_X1 U9352 ( .A1(n6839), .A2(n6842), .ZN(n14329) );
  MUX2_X1 U9353 ( .A(n14315), .B(n14314), .S(n15670), .Z(n14316) );
  MUX2_X1 U9354 ( .A(n14320), .B(n14409), .S(n15670), .Z(n14321) );
  OR2_X1 U9355 ( .A1(n14097), .A2(n14401), .ZN(n10275) );
  OAI21_X1 U9356 ( .B1(n7340), .B2(n15667), .A(n6755), .ZN(n10276) );
  NAND2_X1 U9357 ( .A1(n15667), .A2(n10273), .ZN(n6755) );
  MUX2_X1 U9358 ( .A(n9617), .B(n14314), .S(n15659), .Z(n9620) );
  MUX2_X1 U9359 ( .A(n15873), .B(n14409), .S(n15659), .Z(n14410) );
  NAND2_X1 U9360 ( .A1(n6843), .A2(n6840), .ZN(P2_U3494) );
  AOI21_X1 U9361 ( .B1(n14415), .B2(n15659), .A(n6841), .ZN(n6840) );
  INV_X1 U9362 ( .A(n14416), .ZN(n6843) );
  NOR2_X1 U9363 ( .A1(n15659), .A2(n15895), .ZN(n6841) );
  OR2_X1 U9364 ( .A1(n14097), .A2(n14461), .ZN(n10278) );
  OAI21_X1 U9365 ( .B1(n7340), .B2(n15657), .A(n7339), .ZN(n10279) );
  NAND2_X1 U9366 ( .A1(n15657), .A2(n10277), .ZN(n7339) );
  NAND2_X1 U9367 ( .A1(n7074), .A2(n7910), .ZN(n7154) );
  XNOR2_X1 U9368 ( .A(n14606), .B(n7173), .ZN(n14620) );
  NAND2_X1 U9369 ( .A1(n6781), .A2(n12792), .ZN(P1_U3242) );
  OAI21_X1 U9370 ( .B1(n12788), .B2(n6782), .A(n7176), .ZN(n6781) );
  NAND2_X1 U9371 ( .A1(n6896), .A2(n6893), .ZN(P1_U3356) );
  OR2_X1 U9372 ( .A1(n12990), .A2(n14938), .ZN(n6896) );
  INV_X1 U9373 ( .A(n6894), .ZN(n6893) );
  OAI211_X1 U9374 ( .C1(n7304), .C2(n7301), .A(n7302), .B(n7299), .ZN(P1_U3557) );
  OR2_X1 U9375 ( .A1(n15492), .A2(n7303), .ZN(n7302) );
  NAND2_X1 U9376 ( .A1(n7300), .A2(n15492), .ZN(n7299) );
  INV_X1 U9377 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7303) );
  INV_X1 U9378 ( .A(n7836), .ZN(n7835) );
  OAI21_X1 U9379 ( .B1(n7837), .B2(n7301), .A(n7839), .ZN(n7836) );
  OR2_X1 U9380 ( .A1(n15492), .A2(n15110), .ZN(n7839) );
  NAND2_X1 U9381 ( .A1(n6796), .A2(n7274), .ZN(P1_U3525) );
  NAND2_X1 U9382 ( .A1(n15477), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7274) );
  INV_X1 U9383 ( .A(n7304), .ZN(n6797) );
  NAND2_X1 U9384 ( .A1(n7171), .A2(n7170), .ZN(P1_U3524) );
  NAND2_X1 U9385 ( .A1(n15477), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7170) );
  NAND2_X1 U9386 ( .A1(n15477), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6904) );
  NAND2_X1 U9387 ( .A1(n15195), .A2(n15478), .ZN(n6905) );
  NAND2_X1 U9388 ( .A1(n7497), .A2(n7498), .ZN(n10775) );
  NAND2_X1 U9389 ( .A1(n15270), .A2(n15271), .ZN(n15275) );
  NAND2_X1 U9390 ( .A1(n7511), .A2(n15272), .ZN(n15276) );
  OAI21_X1 U9391 ( .B1(n15270), .B2(n7179), .A(n7508), .ZN(n15286) );
  NAND2_X1 U9392 ( .A1(n7106), .A2(n7178), .ZN(n15287) );
  NAND2_X1 U9393 ( .A1(n15304), .A2(n15303), .ZN(n15306) );
  INV_X1 U9394 ( .A(n13901), .ZN(n7751) );
  OR2_X1 U9395 ( .A1(n10125), .A2(n7902), .ZN(n6544) );
  NAND2_X1 U9396 ( .A1(n7928), .A2(n12346), .ZN(n12520) );
  INV_X1 U9397 ( .A(n13254), .ZN(n6969) );
  AND2_X1 U9398 ( .A1(n13841), .A2(n7281), .ZN(n6545) );
  AND2_X1 U9399 ( .A1(n13853), .A2(n7725), .ZN(n6546) );
  AND2_X1 U9400 ( .A1(n7844), .A2(n7843), .ZN(n6547) );
  INV_X1 U9401 ( .A(n13914), .ZN(n7327) );
  AND2_X1 U9402 ( .A1(n9452), .A2(n9456), .ZN(n9876) );
  AND2_X2 U9403 ( .A1(n12971), .A2(n14985), .ZN(n15405) );
  INV_X4 U9404 ( .A(n14239), .ZN(n8582) );
  INV_X4 U9405 ( .A(n8958), .ZN(n8854) );
  CLKBUF_X3 U9406 ( .A(n13743), .Z(n13855) );
  INV_X1 U9407 ( .A(n11705), .ZN(n12748) );
  NAND2_X1 U9408 ( .A1(n9161), .A2(n14546), .ZN(n6548) );
  AND2_X1 U9409 ( .A1(n13296), .A2(n6835), .ZN(n6549) );
  OAI21_X1 U9410 ( .B1(n13626), .B2(n7036), .A(n7033), .ZN(n13638) );
  INV_X1 U9411 ( .A(n12751), .ZN(n7813) );
  INV_X1 U9412 ( .A(n7535), .ZN(n7534) );
  NOR2_X1 U9413 ( .A1(n7538), .A2(n7903), .ZN(n7535) );
  NAND2_X1 U9414 ( .A1(n14517), .A2(n7884), .ZN(n7882) );
  NAND2_X1 U9415 ( .A1(n12223), .A2(n12358), .ZN(n6550) );
  AND2_X1 U9416 ( .A1(n13393), .A2(n10122), .ZN(n6551) );
  XNOR2_X1 U9417 ( .A(n14614), .B(n15093), .ZN(n14834) );
  INV_X1 U9418 ( .A(n14834), .ZN(n7260) );
  NOR2_X1 U9419 ( .A1(n13900), .A2(n7650), .ZN(n6552) );
  OR2_X1 U9420 ( .A1(n15303), .A2(n7504), .ZN(n6553) );
  NAND2_X1 U9421 ( .A1(n15238), .A2(n8832), .ZN(n15129) );
  INV_X1 U9422 ( .A(n15129), .ZN(n7662) );
  AND2_X1 U9423 ( .A1(n12510), .A2(n13398), .ZN(n6554) );
  XNOR2_X1 U9424 ( .A(n9433), .B(n9432), .ZN(n13166) );
  INV_X1 U9425 ( .A(n12493), .ZN(n7206) );
  AND4_X1 U9426 ( .A1(n12451), .A2(n12452), .A3(n12509), .A4(n7139), .ZN(n6555) );
  NAND2_X1 U9427 ( .A1(n9103), .A2(n9102), .ZN(n15175) );
  AND2_X1 U9428 ( .A1(n14839), .A2(n14838), .ZN(n6556) );
  INV_X1 U9429 ( .A(n10935), .ZN(n7368) );
  INV_X1 U9430 ( .A(n13810), .ZN(n7727) );
  AND2_X1 U9431 ( .A1(n7546), .A2(n7553), .ZN(n6557) );
  AND2_X1 U9432 ( .A1(n10772), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6558) );
  INV_X1 U9433 ( .A(n12505), .ZN(n7220) );
  INV_X1 U9434 ( .A(n9836), .ZN(n7551) );
  AND2_X1 U9435 ( .A1(n7742), .A2(n12501), .ZN(n6559) );
  AND2_X1 U9436 ( .A1(n7856), .A2(n7855), .ZN(n6560) );
  INV_X1 U9437 ( .A(n13152), .ZN(n7453) );
  AND4_X1 U9438 ( .A1(n13338), .A2(n12509), .A3(n7139), .A4(n12508), .ZN(n6561) );
  INV_X1 U9439 ( .A(n7228), .ZN(n7227) );
  AND2_X1 U9440 ( .A1(n7265), .A2(n12914), .ZN(n6562) );
  NAND2_X1 U9441 ( .A1(n15271), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7512) );
  INV_X1 U9442 ( .A(n7512), .ZN(n7179) );
  AND2_X1 U9443 ( .A1(n7057), .A2(n7059), .ZN(n6563) );
  NOR2_X1 U9444 ( .A1(n12686), .A2(n12688), .ZN(n6564) );
  AND2_X1 U9445 ( .A1(n6823), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U9446 ( .A1(n12502), .A2(n12418), .ZN(n6566) );
  NOR2_X1 U9447 ( .A1(n13002), .A2(n6956), .ZN(n6567) );
  NOR2_X1 U9448 ( .A1(n8621), .A2(n8620), .ZN(n6568) );
  AND2_X1 U9449 ( .A1(n7507), .A2(n7506), .ZN(n6569) );
  AND3_X1 U9450 ( .A1(n6888), .A2(n7878), .A3(n7244), .ZN(n6570) );
  AND2_X1 U9451 ( .A1(n7467), .A2(n12709), .ZN(n6571) );
  INV_X1 U9452 ( .A(n13854), .ZN(n7725) );
  AND2_X1 U9453 ( .A1(n12524), .A2(n12522), .ZN(n6572) );
  AND2_X1 U9454 ( .A1(n12529), .A2(n12530), .ZN(n6573) );
  NOR2_X1 U9455 ( .A1(n12598), .A2(n14645), .ZN(n6574) );
  NOR2_X1 U9456 ( .A1(n7007), .A2(n6686), .ZN(n6575) );
  OR2_X1 U9457 ( .A1(n7727), .A2(n13809), .ZN(n6576) );
  INV_X1 U9458 ( .A(n12706), .ZN(n7002) );
  INV_X1 U9459 ( .A(n13902), .ZN(n7321) );
  AND2_X1 U9460 ( .A1(n9845), .A2(n7240), .ZN(n6577) );
  AND2_X1 U9461 ( .A1(n9593), .A2(n7602), .ZN(n6578) );
  OR2_X1 U9462 ( .A1(n13166), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6579) );
  OR2_X1 U9463 ( .A1(n7313), .A2(n7312), .ZN(n6580) );
  AND2_X1 U9464 ( .A1(n11058), .A2(n10108), .ZN(n6581) );
  AND2_X1 U9465 ( .A1(n7410), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6582) );
  AND2_X1 U9466 ( .A1(n9571), .A2(n13260), .ZN(n6583) );
  NOR2_X1 U9467 ( .A1(n10916), .A2(n7401), .ZN(n10782) );
  INV_X1 U9468 ( .A(n13789), .ZN(n7843) );
  NOR2_X1 U9469 ( .A1(n15543), .A2(n7366), .ZN(n7365) );
  INV_X1 U9470 ( .A(n14389), .ZN(n7626) );
  AND2_X1 U9471 ( .A1(n6971), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n6584) );
  INV_X1 U9472 ( .A(n10919), .ZN(n7449) );
  NOR2_X1 U9473 ( .A1(n6583), .A2(n6810), .ZN(n6585) );
  NAND2_X1 U9474 ( .A1(n10518), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7464) );
  INV_X1 U9475 ( .A(n7464), .ZN(n7463) );
  INV_X1 U9476 ( .A(n13146), .ZN(n6827) );
  AND2_X1 U9477 ( .A1(n7418), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6586) );
  NAND2_X1 U9478 ( .A1(n9961), .A2(n9960), .ZN(n13057) );
  INV_X1 U9479 ( .A(n9474), .ZN(n12462) );
  INV_X1 U9480 ( .A(n10836), .ZN(n9518) );
  NAND2_X1 U9481 ( .A1(n7212), .A2(n7210), .ZN(n6587) );
  NAND2_X1 U9482 ( .A1(n7604), .A2(n8140), .ZN(n7606) );
  NAND2_X1 U9483 ( .A1(n7454), .A2(n13221), .ZN(n13239) );
  INV_X1 U9484 ( .A(n14910), .ZN(n7307) );
  INV_X1 U9485 ( .A(n9715), .ZN(n10026) );
  OAI211_X2 U9486 ( .C1(n10048), .C2(n10060), .A(n9630), .B(n10232), .ZN(n9715) );
  NOR2_X1 U9487 ( .A1(n9035), .A2(n9034), .ZN(n6588) );
  OAI211_X1 U9488 ( .C1(n14586), .C2(n6771), .A(n9262), .B(n6770), .ZN(n14606)
         );
  NAND2_X1 U9489 ( .A1(n14489), .A2(n9119), .ZN(n14535) );
  XNOR2_X1 U9490 ( .A(n13057), .B(n13414), .ZN(n12541) );
  INV_X1 U9491 ( .A(n12541), .ZN(n7202) );
  NAND2_X1 U9492 ( .A1(n10170), .A2(n10169), .ZN(n10178) );
  NAND2_X1 U9493 ( .A1(n7747), .A2(n13901), .ZN(n11954) );
  NAND2_X1 U9494 ( .A1(n7322), .A2(n7320), .ZN(n11956) );
  NOR2_X1 U9495 ( .A1(n13689), .A2(n7801), .ZN(n6589) );
  OR2_X1 U9496 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6590) );
  OR2_X1 U9497 ( .A1(n8673), .A2(n7800), .ZN(n6591) );
  AND2_X1 U9498 ( .A1(n7260), .A2(n14853), .ZN(n6592) );
  NOR2_X1 U9499 ( .A1(n8263), .A2(n7338), .ZN(n6593) );
  INV_X1 U9500 ( .A(n10228), .ZN(n7745) );
  NAND2_X1 U9501 ( .A1(n13507), .A2(n13094), .ZN(n10228) );
  AND2_X1 U9502 ( .A1(n15797), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6594) );
  AND2_X1 U9503 ( .A1(n14345), .A2(n13664), .ZN(n6595) );
  NAND2_X1 U9504 ( .A1(n9756), .A2(n9755), .ZN(n9643) );
  XNOR2_X1 U9505 ( .A(n15434), .B(n11687), .ZN(n12754) );
  XNOR2_X1 U9506 ( .A(n15427), .B(n12581), .ZN(n15367) );
  AND2_X1 U9507 ( .A1(n14242), .A2(n14222), .ZN(n14204) );
  AND2_X1 U9508 ( .A1(n11235), .A2(n8541), .ZN(n14239) );
  NAND2_X1 U9509 ( .A1(n8409), .A2(n8408), .ZN(n14109) );
  OR2_X1 U9510 ( .A1(n10224), .A2(n10223), .ZN(n6596) );
  NAND2_X1 U9511 ( .A1(n12338), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n6597) );
  AND2_X1 U9512 ( .A1(n14950), .A2(n7659), .ZN(n6598) );
  NAND2_X1 U9513 ( .A1(n13360), .A2(n13369), .ZN(n6599) );
  NAND2_X1 U9514 ( .A1(n9008), .A2(n9007), .ZN(n12603) );
  XNOR2_X1 U9515 ( .A(n9473), .B(P3_IR_REG_21__SCAN_IN), .ZN(n9625) );
  INV_X1 U9516 ( .A(n15039), .ZN(n7271) );
  NAND2_X1 U9517 ( .A1(n8638), .A2(n8637), .ZN(n6600) );
  INV_X1 U9518 ( .A(n8947), .ZN(n8812) );
  AND3_X1 U9519 ( .A1(n12840), .A2(n14307), .A3(n12839), .ZN(n6601) );
  NAND2_X1 U9520 ( .A1(n10127), .A2(n10126), .ZN(n13350) );
  NAND2_X1 U9521 ( .A1(n7226), .A2(n10117), .ZN(n12219) );
  NAND2_X1 U9522 ( .A1(n6867), .A2(n6870), .ZN(n13380) );
  AND2_X1 U9523 ( .A1(n10323), .A2(n10372), .ZN(n6602) );
  AND2_X1 U9524 ( .A1(n7994), .A2(n7581), .ZN(n6603) );
  NOR3_X1 U9525 ( .A1(n14204), .A2(n14219), .A3(n8582), .ZN(n6604) );
  XNOR2_X1 U9526 ( .A(n9396), .B(P3_IR_REG_6__SCAN_IN), .ZN(n9671) );
  INV_X1 U9527 ( .A(n12499), .ZN(n7893) );
  INV_X1 U9528 ( .A(n14880), .ZN(n7140) );
  INV_X1 U9529 ( .A(n14981), .ZN(n7310) );
  OR2_X1 U9530 ( .A1(n8832), .A2(n14656), .ZN(n6605) );
  AOI21_X1 U9531 ( .B1(n12893), .B2(n8694), .A(n12894), .ZN(n12898) );
  AND3_X1 U9532 ( .A1(n7560), .A2(n7562), .A3(n9357), .ZN(n9438) );
  NOR2_X1 U9533 ( .A1(n15500), .A2(n7356), .ZN(n6606) );
  INV_X1 U9534 ( .A(n13823), .ZN(n7286) );
  INV_X1 U9535 ( .A(n13832), .ZN(n7732) );
  INV_X1 U9536 ( .A(n13844), .ZN(n7735) );
  INV_X1 U9537 ( .A(n10786), .ZN(n9544) );
  AND2_X1 U9538 ( .A1(n7672), .A2(n11705), .ZN(n6607) );
  NAND2_X1 U9539 ( .A1(n7032), .A2(n8654), .ZN(n13637) );
  AND2_X1 U9540 ( .A1(n6579), .A2(n11466), .ZN(n6608) );
  AND2_X1 U9541 ( .A1(n8029), .A2(n8030), .ZN(n8068) );
  AND2_X1 U9542 ( .A1(n14572), .A2(n12581), .ZN(n6609) );
  OR2_X1 U9543 ( .A1(n12714), .A2(n10587), .ZN(n6610) );
  AND2_X1 U9544 ( .A1(n9171), .A2(n9172), .ZN(n6611) );
  NAND2_X1 U9545 ( .A1(n9247), .A2(n9246), .ZN(n14879) );
  INV_X1 U9546 ( .A(n15284), .ZN(n7509) );
  OR2_X1 U9547 ( .A1(n9693), .A2(n10107), .ZN(n6612) );
  AND2_X1 U9548 ( .A1(n14399), .A2(n11434), .ZN(n6613) );
  AND3_X1 U9549 ( .A1(n8577), .A2(n10537), .A3(n13602), .ZN(n6614) );
  NAND2_X1 U9550 ( .A1(n9083), .A2(n9082), .ZN(n15183) );
  AND2_X1 U9551 ( .A1(n9954), .A2(n13101), .ZN(n6615) );
  OR2_X1 U9552 ( .A1(n8775), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n6616) );
  INV_X1 U9553 ( .A(n13777), .ZN(n15641) );
  OR2_X1 U9554 ( .A1(n15304), .A2(n15303), .ZN(n6617) );
  AND2_X1 U9555 ( .A1(n7683), .A2(n7682), .ZN(n6618) );
  AND2_X1 U9556 ( .A1(n13239), .A2(n7461), .ZN(n6619) );
  INV_X1 U9557 ( .A(n7413), .ZN(n7412) );
  AND2_X1 U9558 ( .A1(n14872), .A2(n14871), .ZN(n6620) );
  AND2_X1 U9559 ( .A1(n7698), .A2(n7055), .ZN(n6621) );
  AND2_X1 U9560 ( .A1(n7596), .A2(n7981), .ZN(n6622) );
  OR2_X1 U9561 ( .A1(n10124), .A2(n13022), .ZN(n6623) );
  AND2_X1 U9562 ( .A1(n13110), .A2(n11094), .ZN(n6624) );
  INV_X1 U9563 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9372) );
  INV_X1 U9564 ( .A(n7524), .ZN(n7523) );
  OAI22_X1 U9565 ( .A1(n12992), .A2(n7525), .B1(n13324), .B2(n12883), .ZN(
        n7524) );
  AND2_X1 U9566 ( .A1(n12706), .A2(n7003), .ZN(n6625) );
  OR2_X1 U9567 ( .A1(n7637), .A2(n7635), .ZN(n6626) );
  INV_X1 U9568 ( .A(n14368), .ZN(n14222) );
  NAND2_X1 U9569 ( .A1(n8322), .A2(n8321), .ZN(n14368) );
  AND2_X1 U9570 ( .A1(n13570), .A2(n6600), .ZN(n6627) );
  AND2_X1 U9571 ( .A1(n12426), .A2(n12438), .ZN(n12501) );
  INV_X1 U9572 ( .A(n12501), .ZN(n7736) );
  NAND2_X1 U9573 ( .A1(n12302), .A2(n13103), .ZN(n6628) );
  AND2_X1 U9574 ( .A1(n10362), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6629) );
  INV_X1 U9575 ( .A(n7537), .ZN(n7536) );
  NAND2_X1 U9576 ( .A1(n7542), .A2(n7540), .ZN(n7537) );
  AND2_X1 U9577 ( .A1(n6599), .A2(n10126), .ZN(n6630) );
  AND2_X1 U9578 ( .A1(n9116), .A2(n9099), .ZN(n6631) );
  AND2_X1 U9579 ( .A1(n7095), .A2(n12431), .ZN(n6632) );
  INV_X1 U9580 ( .A(n13860), .ZN(n7723) );
  INV_X1 U9581 ( .A(n7365), .ZN(n7364) );
  NOR2_X1 U9582 ( .A1(n14368), .A2(n14231), .ZN(n6633) );
  INV_X1 U9583 ( .A(n7544), .ZN(n7543) );
  AND2_X1 U9584 ( .A1(n14383), .A2(n8274), .ZN(n6634) );
  AND2_X1 U9585 ( .A1(n13042), .A2(n13049), .ZN(n6635) );
  NAND2_X1 U9586 ( .A1(n15272), .A2(n15274), .ZN(n7513) );
  INV_X1 U9587 ( .A(n7513), .ZN(n7510) );
  NAND2_X1 U9588 ( .A1(n12277), .A2(n7899), .ZN(n13424) );
  INV_X1 U9589 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8743) );
  INV_X1 U9590 ( .A(n7884), .ZN(n7883) );
  AND2_X1 U9591 ( .A1(n12371), .A2(n12368), .ZN(n6636) );
  AND2_X1 U9592 ( .A1(n12590), .A2(n12591), .ZN(n6637) );
  AND2_X1 U9593 ( .A1(n9189), .A2(n9190), .ZN(n6638) );
  AND2_X1 U9594 ( .A1(n13881), .A2(n13882), .ZN(n6639) );
  NAND2_X1 U9595 ( .A1(n8943), .A2(n11421), .ZN(n6640) );
  NAND2_X1 U9596 ( .A1(n10724), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6641) );
  NOR2_X1 U9597 ( .A1(n13843), .A2(n7735), .ZN(n6642) );
  NAND2_X1 U9598 ( .A1(n15093), .A2(n14614), .ZN(n6643) );
  INV_X1 U9599 ( .A(n7823), .ZN(n7822) );
  NOR2_X1 U9600 ( .A1(n15166), .A2(n15016), .ZN(n6644) );
  OR2_X1 U9601 ( .A1(n14152), .A2(n7349), .ZN(n6645) );
  NOR2_X1 U9602 ( .A1(n14955), .A2(n14580), .ZN(n6646) );
  NOR2_X1 U9603 ( .A1(n15156), .A2(n12913), .ZN(n6647) );
  INV_X1 U9604 ( .A(n7335), .ZN(n7334) );
  NOR2_X1 U9605 ( .A1(n8275), .A2(n7336), .ZN(n7335) );
  AND2_X1 U9606 ( .A1(n13327), .A2(n13342), .ZN(n6648) );
  INV_X1 U9607 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7936) );
  OR2_X1 U9608 ( .A1(n12595), .A2(n12594), .ZN(n6649) );
  AND2_X1 U9609 ( .A1(n7010), .A2(n7011), .ZN(n6650) );
  INV_X1 U9610 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10678) );
  NOR2_X1 U9611 ( .A1(n14560), .A2(n7871), .ZN(n6651) );
  INV_X1 U9612 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10428) );
  NOR2_X1 U9613 ( .A1(n13494), .A2(n13290), .ZN(n12521) );
  INV_X1 U9614 ( .A(n10849), .ZN(n9535) );
  AND2_X1 U9615 ( .A1(n15303), .A2(n7504), .ZN(n6652) );
  AND2_X1 U9616 ( .A1(n7722), .A2(n13858), .ZN(n6653) );
  INV_X1 U9617 ( .A(n7903), .ZN(n7542) );
  OR2_X1 U9618 ( .A1(n9467), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n6654) );
  AND2_X1 U9619 ( .A1(n12356), .A2(n12355), .ZN(n13427) );
  INV_X1 U9620 ( .A(n13427), .ZN(n7740) );
  NOR2_X1 U9621 ( .A1(n11832), .A2(n7831), .ZN(n6655) );
  NOR2_X1 U9622 ( .A1(n13859), .A2(n13964), .ZN(n6656) );
  INV_X1 U9623 ( .A(n7828), .ZN(n7827) );
  NAND2_X1 U9624 ( .A1(n14866), .A2(n14885), .ZN(n7828) );
  NAND2_X1 U9625 ( .A1(n10065), .A2(n10064), .ZN(n6657) );
  OR3_X1 U9626 ( .A1(n14841), .A2(n14818), .A3(n7654), .ZN(n6658) );
  OR2_X1 U9627 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6659) );
  AND2_X1 U9628 ( .A1(n7453), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n6660) );
  AND2_X1 U9629 ( .A1(n12472), .A2(n12471), .ZN(n6661) );
  AND3_X1 U9630 ( .A1(n9494), .A2(n9363), .A3(n9362), .ZN(n9367) );
  INV_X1 U9631 ( .A(n8937), .ZN(n8938) );
  OAI21_X1 U9632 ( .B1(n11419), .B2(n14567), .A(n11422), .ZN(n8937) );
  INV_X1 U9633 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6774) );
  AND2_X1 U9634 ( .A1(n9646), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6662) );
  OR2_X1 U9635 ( .A1(n12541), .A2(n7137), .ZN(n6663) );
  AND2_X1 U9636 ( .A1(n14164), .A2(n14428), .ZN(n14126) );
  AND2_X1 U9637 ( .A1(n14849), .A2(n7311), .ZN(n14832) );
  INV_X1 U9638 ( .A(n14832), .ZN(n7100) );
  AND2_X1 U9639 ( .A1(n12986), .A2(n12985), .ZN(n6664) );
  AND2_X1 U9640 ( .A1(n7721), .A2(n13860), .ZN(n6665) );
  AND2_X1 U9641 ( .A1(n15539), .A2(n7372), .ZN(n6666) );
  NAND2_X1 U9642 ( .A1(n14849), .A2(n12954), .ZN(n6667) );
  NOR3_X1 U9643 ( .A1(n12768), .A2(n14996), .A3(n14981), .ZN(n6668) );
  INV_X1 U9644 ( .A(n6792), .ZN(n8367) );
  NOR2_X1 U9645 ( .A1(n8357), .A2(n13595), .ZN(n6792) );
  AND2_X1 U9646 ( .A1(n10425), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6669) );
  OR2_X1 U9647 ( .A1(n6594), .A2(n7705), .ZN(n6670) );
  NAND2_X1 U9648 ( .A1(n12456), .A2(n12454), .ZN(n13351) );
  INV_X1 U9649 ( .A(n13351), .ZN(n7139) );
  NAND2_X1 U9650 ( .A1(n7676), .A2(n12952), .ZN(n6671) );
  INV_X1 U9651 ( .A(n12028), .ZN(n7093) );
  INV_X1 U9652 ( .A(n12587), .ZN(n7477) );
  INV_X1 U9653 ( .A(n7379), .ZN(n7377) );
  NAND2_X1 U9654 ( .A1(n7381), .A2(n6641), .ZN(n7379) );
  INV_X1 U9655 ( .A(n12710), .ZN(n7467) );
  INV_X1 U9656 ( .A(n12698), .ZN(n7470) );
  INV_X1 U9657 ( .A(n12703), .ZN(n7474) );
  INV_X1 U9658 ( .A(n13841), .ZN(n7282) );
  NOR2_X1 U9659 ( .A1(n15317), .A2(n15316), .ZN(n6672) );
  INV_X1 U9660 ( .A(n13842), .ZN(n7281) );
  NAND2_X1 U9661 ( .A1(n8887), .A2(n8888), .ZN(n15399) );
  AND3_X1 U9662 ( .A1(n13287), .A2(n7317), .A3(n7316), .ZN(n6673) );
  AND2_X1 U9663 ( .A1(n13450), .A2(n13465), .ZN(n6674) );
  OR2_X1 U9664 ( .A1(n9569), .A2(n9876), .ZN(n6675) );
  AND2_X1 U9665 ( .A1(n13898), .A2(n13876), .ZN(n6676) );
  AND2_X1 U9666 ( .A1(n12528), .A2(n6572), .ZN(n6677) );
  NOR2_X1 U9667 ( .A1(n11885), .A2(n6588), .ZN(n6678) );
  AND2_X1 U9668 ( .A1(n7852), .A2(n14413), .ZN(n6679) );
  AND2_X1 U9669 ( .A1(n12978), .A2(n7311), .ZN(n6680) );
  AND2_X1 U9670 ( .A1(n15095), .A2(n15094), .ZN(n6681) );
  NAND2_X1 U9671 ( .A1(n8697), .A2(n8696), .ZN(n6682) );
  AND2_X1 U9672 ( .A1(n12884), .A2(n10164), .ZN(n6683) );
  OR2_X1 U9673 ( .A1(n7637), .A2(n7636), .ZN(n6684) );
  AND2_X1 U9674 ( .A1(n8515), .A2(n8514), .ZN(n6685) );
  NOR2_X1 U9675 ( .A1(n8184), .A2(n7948), .ZN(n8202) );
  AND2_X1 U9676 ( .A1(n7470), .A2(n12697), .ZN(n6686) );
  AND2_X1 U9677 ( .A1(n10120), .A2(n10119), .ZN(n6687) );
  AND2_X1 U9678 ( .A1(n12407), .A2(n12405), .ZN(n6688) );
  INV_X1 U9679 ( .A(n12667), .ZN(n6994) );
  AND2_X1 U9680 ( .A1(n6988), .A2(n12579), .ZN(n6689) );
  OR2_X1 U9681 ( .A1(n13821), .A2(n13819), .ZN(n6690) );
  OR2_X1 U9682 ( .A1(n7725), .A2(n13853), .ZN(n6691) );
  AND2_X1 U9683 ( .A1(n15704), .A2(n8743), .ZN(n6692) );
  NAND2_X1 U9684 ( .A1(n13823), .A2(n7287), .ZN(n6693) );
  AND2_X1 U9685 ( .A1(n12461), .A2(n12460), .ZN(n13322) );
  AND2_X1 U9686 ( .A1(n7378), .A2(n7376), .ZN(n6694) );
  OR2_X1 U9687 ( .A1(n7011), .A2(n7010), .ZN(n6695) );
  INV_X1 U9688 ( .A(n10109), .ZN(n7897) );
  NAND2_X1 U9689 ( .A1(n12406), .A2(n6688), .ZN(n6696) );
  OR2_X1 U9690 ( .A1(n13831), .A2(n7732), .ZN(n6697) );
  INV_X1 U9691 ( .A(n13794), .ZN(n12061) );
  NOR2_X1 U9692 ( .A1(n14926), .A2(n12948), .ZN(n6698) );
  OR2_X1 U9693 ( .A1(n6591), .A2(n7028), .ZN(n6699) );
  OR2_X1 U9694 ( .A1(n9671), .A2(n9539), .ZN(n6700) );
  INV_X1 U9695 ( .A(n7548), .ZN(n7547) );
  INV_X1 U9696 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n15811) );
  INV_X1 U9697 ( .A(n7254), .ZN(n7253) );
  NAND2_X1 U9698 ( .A1(n7256), .A2(n6643), .ZN(n7254) );
  INV_X1 U9699 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8012) );
  INV_X1 U9700 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7244) );
  INV_X1 U9701 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9379) );
  INV_X1 U9702 ( .A(n7558), .ZN(n7557) );
  NAND2_X1 U9703 ( .A1(n12861), .A2(n7559), .ZN(n7558) );
  NAND2_X1 U9704 ( .A1(n12588), .A2(n7477), .ZN(n6701) );
  INV_X1 U9705 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10432) );
  AND2_X2 U9706 ( .A1(n12724), .A2(n12561), .ZN(n12571) );
  NAND2_X1 U9707 ( .A1(n10025), .A2(n10024), .ZN(n13360) );
  INV_X1 U9708 ( .A(n13360), .ZN(n7237) );
  NAND2_X1 U9709 ( .A1(n7404), .A2(n13166), .ZN(n7409) );
  INV_X1 U9710 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n6887) );
  AND2_X1 U9711 ( .A1(n13944), .A2(n11289), .ZN(n11235) );
  NAND2_X1 U9712 ( .A1(n8365), .A2(n8364), .ZN(n14353) );
  INV_X1 U9713 ( .A(n14353), .ZN(n7855) );
  NAND2_X1 U9714 ( .A1(n10130), .A2(n10129), .ZN(n13507) );
  AND3_X1 U9715 ( .A1(n11527), .A2(n6547), .A3(n12061), .ZN(n11872) );
  NOR2_X1 U9716 ( .A1(n14288), .A2(n7849), .ZN(n12188) );
  NAND2_X1 U9717 ( .A1(n7765), .A2(n7764), .ZN(n11537) );
  INV_X1 U9718 ( .A(n15150), .ZN(n7119) );
  AND2_X1 U9719 ( .A1(n14242), .A2(n7858), .ZN(n6702) );
  XNOR2_X1 U9720 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9755) );
  INV_X1 U9721 ( .A(n9755), .ZN(n7059) );
  INV_X1 U9722 ( .A(n7443), .ZN(n7442) );
  NOR2_X1 U9723 ( .A1(n13187), .A2(n11487), .ZN(n7443) );
  NAND2_X1 U9724 ( .A1(n7323), .A2(n13914), .ZN(n11552) );
  AND2_X1 U9725 ( .A1(n15566), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U9726 ( .A1(n6929), .A2(n7889), .ZN(n12142) );
  NAND2_X1 U9727 ( .A1(n7757), .A2(n12404), .ZN(n11247) );
  OR2_X1 U9728 ( .A1(n13501), .A2(n13482), .ZN(n6704) );
  NOR2_X1 U9729 ( .A1(n6979), .A2(n11482), .ZN(n11311) );
  XOR2_X1 U9730 ( .A(n8697), .B(n8696), .Z(n6705) );
  NOR2_X1 U9731 ( .A1(n8775), .A2(n7096), .ZN(n9300) );
  OAI21_X1 U9732 ( .B1(n10049), .B2(P3_D_REG_0__SCAN_IN), .A(n9624), .ZN(
        n10048) );
  OAI21_X1 U9733 ( .B1(n8937), .B2(n11015), .A(n6768), .ZN(n11271) );
  INV_X1 U9734 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9446) );
  OR2_X1 U9735 ( .A1(n13501), .A2(n13536), .ZN(n6706) );
  NAND2_X1 U9736 ( .A1(n9463), .A2(n9462), .ZN(n9467) );
  AND2_X1 U9737 ( .A1(n10761), .A2(n14700), .ZN(n6707) );
  INV_X1 U9738 ( .A(n7022), .ZN(n8618) );
  NAND2_X1 U9739 ( .A1(n8611), .A2(n11191), .ZN(n7022) );
  AND2_X1 U9740 ( .A1(n11737), .A2(n11736), .ZN(n6708) );
  AND2_X1 U9741 ( .A1(n7209), .A2(n10096), .ZN(n6709) );
  INV_X1 U9742 ( .A(n7851), .ZN(n14270) );
  NOR2_X1 U9743 ( .A1(n14288), .A2(n7848), .ZN(n7851) );
  AND2_X1 U9744 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n6710) );
  AND2_X1 U9745 ( .A1(n6582), .A2(n7409), .ZN(n6711) );
  AND2_X1 U9746 ( .A1(n9508), .A2(n13166), .ZN(n13175) );
  AND2_X1 U9747 ( .A1(n7774), .A2(n7773), .ZN(n6712) );
  INV_X1 U9748 ( .A(n6814), .ZN(n6813) );
  NOR2_X1 U9749 ( .A1(n9565), .A2(n10482), .ZN(n6814) );
  NAND2_X1 U9750 ( .A1(n8511), .A2(n8510), .ZN(n6713) );
  NAND2_X1 U9751 ( .A1(n14714), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U9752 ( .A1(n10465), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6715) );
  NOR2_X1 U9753 ( .A1(n6587), .A2(n10106), .ZN(n6716) );
  AND2_X1 U9754 ( .A1(n9442), .A2(n10282), .ZN(n6717) );
  AND2_X1 U9755 ( .A1(n7242), .A2(n7241), .ZN(n6718) );
  NAND2_X1 U9756 ( .A1(n7782), .A2(n11528), .ZN(n15642) );
  NAND2_X1 U9757 ( .A1(n8287), .A2(n8286), .ZN(n14259) );
  INV_X1 U9758 ( .A(n14259), .ZN(n7850) );
  NAND2_X1 U9759 ( .A1(n7403), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7401) );
  AND2_X2 U9760 ( .A1(n10247), .A2(n10246), .ZN(n15693) );
  INV_X2 U9761 ( .A(n15657), .ZN(n15659) );
  INV_X2 U9762 ( .A(n15667), .ZN(n15670) );
  AND2_X2 U9763 ( .A1(n11664), .A2(n10778), .ZN(n15478) );
  AND2_X1 U9764 ( .A1(n9852), .A2(n13104), .ZN(n6719) );
  INV_X1 U9765 ( .A(n10518), .ZN(n7312) );
  AND2_X2 U9766 ( .A1(n10214), .A2(n10252), .ZN(n13486) );
  INV_X1 U9767 ( .A(n13486), .ZN(n13478) );
  NAND2_X1 U9768 ( .A1(n10042), .A2(n10193), .ZN(n10060) );
  INV_X1 U9769 ( .A(n13428), .ZN(n13398) );
  NAND2_X1 U9770 ( .A1(n6877), .A2(n7076), .ZN(n11277) );
  NAND2_X1 U9771 ( .A1(n9145), .A2(n9144), .ZN(n15166) );
  INV_X1 U9772 ( .A(n15166), .ZN(n7663) );
  INV_X1 U9773 ( .A(n13207), .ZN(n10482) );
  AND2_X2 U9774 ( .A1(n10779), .A2(n10778), .ZN(n15492) );
  INV_X1 U9775 ( .A(n15492), .ZN(n7301) );
  INV_X1 U9776 ( .A(n10970), .ZN(n7423) );
  INV_X1 U9777 ( .A(n14307), .ZN(n14217) );
  AND2_X1 U9778 ( .A1(n6976), .A2(n11481), .ZN(n6720) );
  NAND2_X1 U9779 ( .A1(n7422), .A2(n7421), .ZN(n10969) );
  AND2_X1 U9780 ( .A1(n7397), .A2(n10915), .ZN(n6721) );
  OR2_X1 U9781 ( .A1(n10916), .A2(n7402), .ZN(n6722) );
  AND2_X1 U9782 ( .A1(n9595), .A2(n15965), .ZN(n6723) );
  AND2_X1 U9783 ( .A1(n6584), .A2(n6970), .ZN(n6724) );
  NAND2_X1 U9784 ( .A1(n7444), .A2(n7449), .ZN(n6725) );
  INV_X1 U9785 ( .A(n13281), .ZN(n6971) );
  NAND2_X1 U9786 ( .A1(n11527), .A2(n6547), .ZN(n7845) );
  AND2_X1 U9787 ( .A1(n11365), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6726) );
  AND2_X1 U9788 ( .A1(n7380), .A2(n7381), .ZN(n6727) );
  AND2_X1 U9789 ( .A1(n11415), .A2(n10930), .ZN(n12365) );
  INV_X1 U9790 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7719) );
  INV_X1 U9791 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7372) );
  INV_X1 U9792 ( .A(n9575), .ZN(n6970) );
  INV_X1 U9793 ( .A(n10841), .ZN(n6831) );
  AND2_X1 U9794 ( .A1(n12794), .A2(n12326), .ZN(n6728) );
  AND2_X1 U9795 ( .A1(n7105), .A2(n10750), .ZN(n6729) );
  INV_X1 U9796 ( .A(n10498), .ZN(n7840) );
  INV_X1 U9797 ( .A(SI_24_), .ZN(n7581) );
  INV_X1 U9798 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7504) );
  INV_X1 U9799 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7298) );
  NAND2_X1 U9800 ( .A1(n10186), .A2(n9748), .ZN(n12343) );
  AOI21_X1 U9801 ( .B1(n13303), .B2(n9748), .A(n10177), .ZN(n10201) );
  NAND2_X1 U9802 ( .A1(n13315), .A2(n9748), .ZN(n10163) );
  NAND2_X1 U9803 ( .A1(n13328), .A2(n9748), .ZN(n10149) );
  NAND2_X1 U9804 ( .A1(n13346), .A2(n9748), .ZN(n10079) );
  NAND2_X1 U9805 ( .A1(n13374), .A2(n9748), .ZN(n10018) );
  NAND2_X1 U9806 ( .A1(n13388), .A2(n9748), .ZN(n10005) );
  NAND2_X1 U9807 ( .A1(n10080), .A2(n9748), .ZN(n10034) );
  NAND2_X1 U9808 ( .A1(n13064), .A2(n9748), .ZN(n9968) );
  NAND2_X1 U9809 ( .A1(n13401), .A2(n9748), .ZN(n9987) );
  NAND2_X1 U9810 ( .A1(n13409), .A2(n9748), .ZN(n9953) );
  NAND2_X1 U9811 ( .A1(n13434), .A2(n9748), .ZN(n9939) );
  NAND2_X1 U9812 ( .A1(n12297), .A2(n9748), .ZN(n9883) );
  NAND2_X1 U9813 ( .A1(n13041), .A2(n9748), .ZN(n9902) );
  NAND2_X1 U9814 ( .A1(n13054), .A2(n9748), .ZN(n9922) );
  NAND2_X1 U9815 ( .A1(n12211), .A2(n9748), .ZN(n9851) );
  AND2_X2 U9816 ( .A1(n12721), .A2(n9335), .ZN(n15031) );
  AND2_X1 U9817 ( .A1(n15237), .A2(n11695), .ZN(n12721) );
  NAND2_X1 U9818 ( .A1(n6730), .A2(n14800), .ZN(n14802) );
  NAND2_X1 U9819 ( .A1(n14797), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U9820 ( .A1(n14778), .A2(n14777), .ZN(n14799) );
  NAND2_X1 U9821 ( .A1(n12002), .A2(n8067), .ZN(n11255) );
  NAND2_X1 U9822 ( .A1(n12003), .A2(n10897), .ZN(n6731) );
  NAND2_X1 U9823 ( .A1(n6740), .A2(n7746), .ZN(n14301) );
  NAND2_X1 U9824 ( .A1(n11956), .A2(n7748), .ZN(n6740) );
  AOI21_X1 U9825 ( .B1(n7746), .B2(n6742), .A(n6613), .ZN(n6741) );
  INV_X1 U9826 ( .A(n7748), .ZN(n6742) );
  INV_X1 U9827 ( .A(n7746), .ZN(n6743) );
  NAND2_X1 U9828 ( .A1(n14135), .A2(n13924), .ZN(n6864) );
  INV_X1 U9829 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6754) );
  INV_X1 U9830 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6756) );
  NOR2_X1 U9831 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6761) );
  NOR2_X1 U9832 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n6760) );
  NOR2_X2 U9833 ( .A1(n8251), .A2(n8008), .ZN(n8013) );
  NAND2_X2 U9834 ( .A1(n6759), .A2(n8222), .ZN(n8251) );
  AND4_X2 U9835 ( .A1(n8063), .A2(n6761), .A3(n6760), .A4(n8075), .ZN(n6759)
         );
  NOR2_X2 U9836 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8063) );
  OAI21_X1 U9837 ( .B1(n11008), .B2(n11009), .A(n6762), .ZN(n11010) );
  NAND2_X1 U9838 ( .A1(n11008), .A2(n11009), .ZN(n6762) );
  NAND4_X1 U9839 ( .A1(n6765), .A2(n6764), .A3(n8741), .A4(n8742), .ZN(n8804)
         );
  NAND3_X1 U9840 ( .A1(n7875), .A2(n12028), .A3(n12018), .ZN(n6766) );
  AOI21_X2 U9841 ( .B1(n14598), .B2(n14599), .A(n6638), .ZN(n14509) );
  AOI21_X1 U9842 ( .B1(n8938), .B2(n6769), .A(n6640), .ZN(n6768) );
  INV_X1 U9843 ( .A(n7862), .ZN(n6771) );
  INV_X2 U9844 ( .A(n9136), .ZN(n9318) );
  NAND3_X1 U9845 ( .A1(n6784), .A2(n8220), .A3(n6783), .ZN(n7959) );
  NAND4_X1 U9846 ( .A1(n7305), .A2(n7955), .A3(n8202), .A4(n7947), .ZN(n6783)
         );
  NAND2_X2 U9847 ( .A1(n6786), .A2(n6785), .ZN(n7350) );
  NAND4_X1 U9848 ( .A1(n7297), .A2(n7298), .A3(n7935), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n6786) );
  OAI21_X1 U9849 ( .B1(n7350), .B2(n10432), .A(n6787), .ZN(n8085) );
  XNOR2_X2 U9850 ( .A(n6795), .B(n8756), .ZN(n9335) );
  NAND4_X1 U9851 ( .A1(n8754), .A2(n6889), .A3(n6890), .A4(n8755), .ZN(n8759)
         );
  NOR2_X2 U9852 ( .A1(n14855), .A2(n15093), .ZN(n6798) );
  NAND3_X1 U9853 ( .A1(n6807), .A2(n6809), .A3(n6804), .ZN(n13275) );
  NAND3_X1 U9854 ( .A1(n6807), .A2(n6805), .A3(n6804), .ZN(n7152) );
  NOR2_X1 U9855 ( .A1(n13255), .A2(n6583), .ZN(n9572) );
  INV_X1 U9856 ( .A(n13280), .ZN(n6810) );
  OAI21_X1 U9857 ( .B1(n9533), .B2(n6831), .A(n6829), .ZN(n10843) );
  OR2_X1 U9858 ( .A1(n12467), .A2(n6837), .ZN(n6832) );
  NAND2_X1 U9859 ( .A1(n6832), .A2(n6549), .ZN(n12474) );
  NAND4_X1 U9860 ( .A1(n12415), .A2(n12402), .A3(n12401), .A4(n12400), .ZN(
        n6847) );
  NAND2_X1 U9861 ( .A1(n6848), .A2(n6847), .ZN(n12424) );
  AOI21_X1 U9862 ( .B1(n12415), .B2(n6696), .A(n6566), .ZN(n6848) );
  NAND2_X1 U9863 ( .A1(n9481), .A2(n7072), .ZN(n9581) );
  AND2_X2 U9864 ( .A1(n8013), .A2(n8011), .ZN(n8015) );
  NAND3_X1 U9865 ( .A1(n8011), .A2(n6856), .A3(n6855), .ZN(n8028) );
  NAND3_X1 U9866 ( .A1(n6859), .A2(n12370), .A3(n6858), .ZN(n6857) );
  OR2_X1 U9867 ( .A1(n12363), .A2(n9474), .ZN(n6858) );
  NAND2_X1 U9868 ( .A1(n6862), .A2(n12530), .ZN(n7049) );
  OAI21_X1 U9869 ( .B1(n12515), .B2(n12482), .A(n6863), .ZN(n6862) );
  NAND2_X1 U9870 ( .A1(n12515), .A2(n12514), .ZN(n6863) );
  NAND3_X1 U9871 ( .A1(n7762), .A2(n7922), .A3(n7763), .ZN(n6865) );
  NAND2_X1 U9872 ( .A1(n6866), .A2(n6868), .ZN(n10226) );
  NAND2_X1 U9873 ( .A1(n7200), .A2(n6870), .ZN(n6866) );
  NAND2_X1 U9874 ( .A1(n11277), .A2(n12406), .ZN(n6876) );
  NAND2_X1 U9875 ( .A1(n9742), .A2(n10344), .ZN(n9709) );
  NAND2_X1 U9876 ( .A1(n6879), .A2(n9567), .ZN(n10285) );
  NAND2_X1 U9877 ( .A1(n13208), .A2(n10282), .ZN(n6879) );
  NOR2_X1 U9878 ( .A1(n7393), .A2(n9406), .ZN(n13120) );
  NOR2_X1 U9879 ( .A1(n6881), .A2(n9406), .ZN(n6880) );
  OR2_X1 U9880 ( .A1(n10966), .A2(n9525), .ZN(n6881) );
  NAND3_X1 U9881 ( .A1(n7419), .A2(n6586), .A3(n13268), .ZN(n7416) );
  NAND4_X1 U9882 ( .A1(n6570), .A2(n8755), .A3(n6889), .A4(n8754), .ZN(n15219)
         );
  NOR2_X2 U9883 ( .A1(n8921), .A2(n8753), .ZN(n8754) );
  NAND2_X2 U9884 ( .A1(n11838), .A2(n7829), .ZN(n11973) );
  OAI21_X2 U9885 ( .B1(n14923), .B2(n12927), .A(n12926), .ZN(n14854) );
  NAND2_X1 U9886 ( .A1(n6899), .A2(n11834), .ZN(n12072) );
  OAI22_X2 U9887 ( .A1(n6899), .A2(n7667), .B1(n7668), .B2(n7905), .ZN(n12105)
         );
  AND2_X1 U9888 ( .A1(n6900), .A2(n6556), .ZN(n15097) );
  NAND2_X1 U9889 ( .A1(n6905), .A2(n6904), .ZN(P1_U3523) );
  OAI21_X2 U9890 ( .B1(n7676), .B2(n6909), .A(n6907), .ZN(n14849) );
  NAND3_X1 U9891 ( .A1(n12939), .A2(n12938), .A3(n15039), .ZN(n6913) );
  NAND2_X2 U9892 ( .A1(n7308), .A2(n7306), .ZN(n15120) );
  MUX2_X1 U9893 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n7350), .Z(n6916) );
  NAND3_X1 U9894 ( .A1(n7114), .A2(n7500), .A3(n7499), .ZN(n15313) );
  NAND2_X1 U9895 ( .A1(n10111), .A2(n7891), .ZN(n6929) );
  NAND4_X1 U9896 ( .A1(n6934), .A2(n6932), .A3(n15691), .A4(n6930), .ZN(n6938)
         );
  NAND2_X1 U9897 ( .A1(n13424), .A2(n6687), .ZN(n13416) );
  NAND3_X1 U9898 ( .A1(n7207), .A2(n10109), .A3(n7205), .ZN(n7204) );
  NAND2_X1 U9899 ( .A1(n13337), .A2(n10133), .ZN(n13341) );
  NAND2_X1 U9900 ( .A1(n9905), .A2(n6943), .ZN(n6940) );
  NAND2_X1 U9901 ( .A1(n6940), .A2(n6941), .ZN(n13061) );
  INV_X1 U9902 ( .A(n6949), .ZN(n11504) );
  NAND3_X1 U9903 ( .A1(n6557), .A2(n7547), .A3(n6951), .ZN(n6952) );
  NAND2_X1 U9904 ( .A1(n11900), .A2(n6954), .ZN(n6953) );
  AOI21_X2 U9905 ( .B1(n13068), .B2(n13022), .A(n10006), .ZN(n13002) );
  NAND2_X1 U9906 ( .A1(n9367), .A2(n9380), .ZN(n9387) );
  NAND2_X1 U9907 ( .A1(n6959), .A2(n6962), .ZN(n13169) );
  NAND2_X1 U9908 ( .A1(n9509), .A2(n7411), .ZN(n6962) );
  NAND2_X1 U9909 ( .A1(n9510), .A2(n6962), .ZN(n6961) );
  NAND2_X1 U9910 ( .A1(n6961), .A2(n11371), .ZN(n6960) );
  NAND3_X1 U9911 ( .A1(n6968), .A2(n6965), .A3(n9575), .ZN(n6964) );
  OR2_X1 U9912 ( .A1(n13254), .A2(n12285), .ZN(n13283) );
  NAND2_X1 U9913 ( .A1(n9505), .A2(n9535), .ZN(n6974) );
  NAND2_X1 U9914 ( .A1(n6975), .A2(n10849), .ZN(n13151) );
  INV_X1 U9915 ( .A(n9505), .ZN(n6975) );
  INV_X1 U9916 ( .A(n11482), .ZN(n6981) );
  NAND2_X1 U9917 ( .A1(n6979), .A2(n6981), .ZN(n6976) );
  NOR2_X1 U9918 ( .A1(n7447), .A2(n11482), .ZN(n11310) );
  NAND2_X1 U9919 ( .A1(n12580), .A2(n6689), .ZN(n6987) );
  NAND2_X1 U9920 ( .A1(n6985), .A2(n6989), .ZN(n12595) );
  NAND3_X1 U9921 ( .A1(n12585), .A2(n6701), .A3(n6986), .ZN(n6985) );
  NAND2_X1 U9922 ( .A1(n6987), .A2(n12582), .ZN(n6986) );
  NAND2_X1 U9923 ( .A1(n7923), .A2(n6990), .ZN(n7482) );
  NAND2_X1 U9924 ( .A1(n12733), .A2(n12558), .ZN(n12724) );
  NAND2_X1 U9925 ( .A1(n12555), .A2(n6997), .ZN(n12560) );
  OR2_X1 U9926 ( .A1(n15237), .A2(n12556), .ZN(n6997) );
  NAND2_X1 U9927 ( .A1(n12705), .A2(n7000), .ZN(n6998) );
  NAND2_X1 U9928 ( .A1(n6998), .A2(n6999), .ZN(n12789) );
  NAND2_X1 U9929 ( .A1(n7004), .A2(n7005), .ZN(n7175) );
  NAND2_X1 U9930 ( .A1(n7174), .A2(n6575), .ZN(n7004) );
  NAND2_X1 U9931 ( .A1(n7008), .A2(n7009), .ZN(n7186) );
  NAND3_X1 U9932 ( .A1(n12682), .A2(n12683), .A3(n6695), .ZN(n7008) );
  INV_X1 U9933 ( .A(n12684), .ZN(n7011) );
  NAND2_X1 U9934 ( .A1(n10688), .A2(n7012), .ZN(n10689) );
  NAND2_X1 U9935 ( .A1(n10562), .A2(n10561), .ZN(n10688) );
  NAND2_X1 U9936 ( .A1(n8578), .A2(n6614), .ZN(n7013) );
  NAND3_X1 U9937 ( .A1(n8576), .A2(n8578), .A3(n13678), .ZN(n7014) );
  OR3_X2 U9938 ( .A1(n8015), .A2(n8266), .A3(n8012), .ZN(n7015) );
  NAND3_X2 U9939 ( .A1(n8027), .A2(n7015), .A3(n6590), .ZN(n10490) );
  NAND2_X1 U9940 ( .A1(n8015), .A2(n8012), .ZN(n8027) );
  OAI22_X2 U9941 ( .A1(n7016), .A2(n8455), .B1(n7783), .B2(n7020), .ZN(n7019)
         );
  NAND2_X2 U9942 ( .A1(n8016), .A2(n7019), .ZN(n13953) );
  NAND2_X1 U9943 ( .A1(n8611), .A2(n7023), .ZN(n7021) );
  NAND2_X1 U9944 ( .A1(n7021), .A2(n7788), .ZN(n8626) );
  NAND2_X1 U9945 ( .A1(n12131), .A2(n7025), .ZN(n7024) );
  NAND2_X1 U9946 ( .A1(n8592), .A2(n7037), .ZN(n7040) );
  NAND2_X1 U9947 ( .A1(n9728), .A2(n9636), .ZN(n9638) );
  NAND2_X1 U9948 ( .A1(n9716), .A2(n9634), .ZN(n7042) );
  NAND2_X1 U9949 ( .A1(n7043), .A2(n7691), .ZN(n10022) );
  NAND2_X1 U9950 ( .A1(n9975), .A2(n7693), .ZN(n7043) );
  NAND2_X1 U9951 ( .A1(n10138), .A2(n10137), .ZN(n10151) );
  NAND2_X1 U9952 ( .A1(n12513), .A2(n12530), .ZN(n7047) );
  NAND4_X1 U9953 ( .A1(n7049), .A2(n7048), .A3(n7047), .A4(n12534), .ZN(
        P3_U3296) );
  NAND3_X1 U9954 ( .A1(n7050), .A2(n6573), .A3(n7188), .ZN(n7048) );
  NOR2_X1 U9955 ( .A1(n6677), .A2(n7051), .ZN(n7050) );
  NAND4_X1 U9956 ( .A1(n12511), .A2(n12510), .A3(n7928), .A4(n7052), .ZN(n7146) );
  NAND3_X1 U9957 ( .A1(n6561), .A2(n13322), .A3(n13312), .ZN(n7053) );
  NAND2_X1 U9958 ( .A1(n9788), .A2(n7063), .ZN(n7060) );
  NAND2_X1 U9959 ( .A1(n7060), .A2(n7061), .ZN(n9818) );
  NAND2_X1 U9960 ( .A1(n9929), .A2(n7069), .ZN(n7066) );
  NAND2_X1 U9961 ( .A1(n7066), .A2(n7067), .ZN(n9958) );
  NAND2_X1 U9962 ( .A1(n7083), .A2(n7196), .ZN(n7200) );
  NAND2_X1 U9963 ( .A1(n7083), .A2(n12353), .ZN(n12538) );
  NAND2_X1 U9964 ( .A1(n12809), .A2(n12810), .ZN(n12808) );
  AND2_X1 U9965 ( .A1(n8881), .A2(n8882), .ZN(n11009) );
  NAND2_X1 U9966 ( .A1(n8250), .A2(n7088), .ZN(n7087) );
  NAND2_X1 U9967 ( .A1(n7087), .A2(n7085), .ZN(n8319) );
  NAND2_X1 U9968 ( .A1(n7875), .A2(n12018), .ZN(n7094) );
  NAND2_X1 U9969 ( .A1(n7773), .A2(n7187), .ZN(n7095) );
  NAND2_X1 U9970 ( .A1(n9300), .A2(n9302), .ZN(n8769) );
  MUX2_X1 U9971 ( .A(n10436), .B(n10371), .S(n7350), .Z(n7946) );
  OAI21_X1 U9972 ( .B1(n14815), .B2(n7104), .A(n10476), .ZN(P1_U3243) );
  INV_X1 U9973 ( .A(n15294), .ZN(n7117) );
  AOI21_X1 U9974 ( .B1(n10773), .B2(n7111), .A(n6558), .ZN(n11750) );
  NAND3_X1 U9975 ( .A1(n7497), .A2(n7498), .A3(n10774), .ZN(n11020) );
  NAND2_X1 U9976 ( .A1(n15298), .A2(n7113), .ZN(n7114) );
  INV_X1 U9977 ( .A(n12103), .ZN(n12101) );
  NAND3_X1 U9978 ( .A1(n7488), .A2(n7491), .A3(n12100), .ZN(n15251) );
  NAND2_X1 U9979 ( .A1(n11025), .A2(n11024), .ZN(n11755) );
  NAND2_X1 U9980 ( .A1(n7117), .A2(n7166), .ZN(n15296) );
  NAND2_X1 U9981 ( .A1(n11477), .A2(n9559), .ZN(n13163) );
  OAI211_X1 U9982 ( .C1(n13338), .C2(n7745), .A(n7167), .B(n12461), .ZN(n7191)
         );
  INV_X1 U9983 ( .A(n7666), .ZN(n7665) );
  NAND3_X1 U9984 ( .A1(n7664), .A2(n7663), .A3(n12106), .ZN(n15034) );
  OAI21_X1 U9985 ( .B1(n13495), .B2(n13478), .A(n7120), .ZN(P3_U3487) );
  OAI21_X1 U9986 ( .B1(n13495), .B2(n15693), .A(n7122), .ZN(P3_U3455) );
  NAND2_X1 U9987 ( .A1(n15246), .A2(n15245), .ZN(n10759) );
  NAND2_X1 U9988 ( .A1(n13602), .A2(n10537), .ZN(n13600) );
  NAND2_X1 U9989 ( .A1(n7492), .A2(n7495), .ZN(n7491) );
  NAND2_X2 U9990 ( .A1(n15560), .A2(n15559), .ZN(n15558) );
  XNOR2_X2 U9991 ( .A(n8064), .B(P2_IR_REG_2__SCAN_IN), .ZN(n12536) );
  NAND2_X1 U9992 ( .A1(n9552), .A2(n10911), .ZN(n11305) );
  NAND2_X1 U9993 ( .A1(n9543), .A2(n13147), .ZN(n10789) );
  OAI21_X2 U9994 ( .B1(n9192), .B2(n9191), .A(n14507), .ZN(n14578) );
  NAND2_X1 U9995 ( .A1(n7129), .A2(n7914), .ZN(P2_U3192) );
  NAND2_X1 U9996 ( .A1(n7149), .A2(n7148), .ZN(n7129) );
  NAND2_X1 U9997 ( .A1(n8105), .A2(n13908), .ZN(n11596) );
  NAND2_X1 U9998 ( .A1(n7344), .A2(n14307), .ZN(n7343) );
  NAND3_X1 U9999 ( .A1(n9442), .A2(n10282), .A3(P3_REG2_REG_13__SCAN_IN), .ZN(
        n13208) );
  INV_X1 U10000 ( .A(n9441), .ZN(n7130) );
  NAND2_X1 U10001 ( .A1(n11465), .A2(n7134), .ZN(n11299) );
  INV_X1 U10002 ( .A(n13252), .ZN(n7417) );
  NAND3_X1 U10003 ( .A1(n12663), .A2(n12661), .A3(n12662), .ZN(n7426) );
  NAND2_X1 U10004 ( .A1(n7136), .A2(n12466), .ZN(n12467) );
  NAND2_X1 U10005 ( .A1(n11681), .A2(n11680), .ZN(n11683) );
  NAND2_X1 U10006 ( .A1(n7177), .A2(n15476), .ZN(n7304) );
  NAND2_X1 U10007 ( .A1(n12105), .A2(n11993), .ZN(n11995) );
  NAND2_X1 U10008 ( .A1(n11734), .A2(n11733), .ZN(n11833) );
  NAND3_X1 U10009 ( .A1(n15085), .A2(n15086), .A3(n15476), .ZN(n15092) );
  NAND2_X1 U10010 ( .A1(n7617), .A2(n7615), .ZN(n14247) );
  XNOR2_X1 U10011 ( .A(n7146), .B(n12526), .ZN(n12512) );
  NAND2_X2 U10012 ( .A1(n8564), .A2(n8563), .ZN(n14322) );
  NAND2_X1 U10013 ( .A1(n15296), .A2(n15592), .ZN(n15298) );
  NAND2_X1 U10014 ( .A1(n7486), .A2(n10315), .ZN(n10322) );
  NAND2_X1 U10015 ( .A1(n7618), .A2(n7622), .ZN(n7617) );
  NAND4_X1 U10016 ( .A1(n7609), .A2(n8509), .A3(n11078), .A4(n8508), .ZN(n7608) );
  NAND2_X1 U10017 ( .A1(n11953), .A2(n7751), .ZN(n11952) );
  OAI21_X1 U10018 ( .B1(n13560), .B2(n13695), .A(n8711), .ZN(n7149) );
  INV_X1 U10019 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7150) );
  INV_X1 U10020 ( .A(n9485), .ZN(n7562) );
  INV_X1 U10021 ( .A(n7152), .ZN(n13274) );
  NAND2_X1 U10022 ( .A1(n9572), .A2(n13280), .ZN(n7151) );
  NAND2_X1 U10023 ( .A1(n13215), .A2(n6675), .ZN(n13234) );
  NAND2_X1 U10024 ( .A1(n9631), .A2(n9700), .ZN(n7153) );
  NAND2_X1 U10025 ( .A1(n12540), .A2(n7201), .ZN(n7203) );
  INV_X1 U10026 ( .A(n10123), .ZN(n7902) );
  NAND2_X1 U10027 ( .A1(n10227), .A2(n7194), .ZN(n7193) );
  NAND3_X1 U10028 ( .A1(n6676), .A2(n7294), .A3(n13878), .ZN(n7293) );
  NAND3_X1 U10029 ( .A1(n7154), .A2(n9352), .A3(n9351), .ZN(P1_U3220) );
  NOR2_X1 U10030 ( .A1(n7877), .A2(n7876), .ZN(n7875) );
  NAND2_X1 U10031 ( .A1(n12813), .A2(n12039), .ZN(n12566) );
  NAND2_X1 U10032 ( .A1(n11676), .A2(n11675), .ZN(n15374) );
  NAND2_X1 U10033 ( .A1(n7157), .A2(n7155), .ZN(n11734) );
  NOR2_X1 U10034 ( .A1(n7156), .A2(n6607), .ZN(n7155) );
  NAND2_X1 U10035 ( .A1(n11683), .A2(n7672), .ZN(n7157) );
  NAND2_X1 U10036 ( .A1(n9818), .A2(n9817), .ZN(n9822) );
  INV_X1 U10037 ( .A(n10098), .ZN(n13117) );
  NAND2_X1 U10038 ( .A1(n13365), .A2(n13367), .ZN(n10127) );
  NAND2_X1 U10039 ( .A1(n13451), .A2(n6704), .ZN(P3_U3486) );
  NAND2_X1 U10040 ( .A1(n13500), .A2(n6706), .ZN(P3_U3454) );
  NAND2_X1 U10041 ( .A1(n10228), .A2(n10131), .ZN(n10132) );
  NAND2_X1 U10042 ( .A1(n13217), .A2(n13216), .ZN(n13215) );
  NAND2_X1 U10043 ( .A1(n7203), .A2(n7900), .ZN(n13365) );
  NAND2_X1 U10044 ( .A1(n9422), .A2(n9544), .ZN(n7403) );
  NAND2_X1 U10045 ( .A1(n7417), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13269) );
  NAND2_X1 U10046 ( .A1(n7390), .A2(n7388), .ZN(n9406) );
  NAND2_X1 U10047 ( .A1(n15120), .A2(n7674), .ZN(n7676) );
  NAND2_X1 U10048 ( .A1(n15194), .A2(n15478), .ZN(n7171) );
  NAND2_X1 U10049 ( .A1(n15092), .A2(n7172), .ZN(n15194) );
  NAND2_X1 U10050 ( .A1(n12796), .A2(n6728), .ZN(n12333) );
  NAND2_X2 U10051 ( .A1(n8089), .A2(n8088), .ZN(n13767) );
  NAND3_X1 U10052 ( .A1(n12696), .A2(n12695), .A3(n7468), .ZN(n7174) );
  NAND2_X1 U10053 ( .A1(n7175), .A2(n7473), .ZN(n12705) );
  OAI21_X1 U10054 ( .B1(n7427), .B2(n7426), .A(n12664), .ZN(n12666) );
  NAND3_X1 U10055 ( .A1(n15024), .A2(n7309), .A3(n7687), .ZN(n7683) );
  NAND2_X1 U10056 ( .A1(n15374), .A2(n7247), .ZN(n15350) );
  NAND3_X1 U10057 ( .A1(n10237), .A2(n10235), .A3(n10236), .ZN(P3_U3488) );
  NAND3_X1 U10058 ( .A1(n10250), .A2(n10248), .A3(n10249), .ZN(P3_U3456) );
  NAND2_X1 U10059 ( .A1(n7601), .A2(n9588), .ZN(n9594) );
  NAND2_X2 U10060 ( .A1(n13568), .A2(n8644), .ZN(n13626) );
  INV_X1 U10061 ( .A(n7901), .ZN(n7900) );
  AND2_X4 U10062 ( .A1(n9663), .A2(n9662), .ZN(n9748) );
  NAND2_X1 U10063 ( .A1(n9476), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9483) );
  AOI21_X1 U10064 ( .B1(n12748), .B2(n7673), .A(n6574), .ZN(n7672) );
  NAND2_X1 U10065 ( .A1(n7941), .A2(n7180), .ZN(n8131) );
  NAND3_X1 U10066 ( .A1(n8080), .A2(n8079), .A3(n8098), .ZN(n7180) );
  NAND2_X1 U10067 ( .A1(n7934), .A2(n11995), .ZN(n12939) );
  NAND2_X2 U10068 ( .A1(n8104), .A2(n8103), .ZN(n15632) );
  NAND2_X1 U10069 ( .A1(n13619), .A2(n8677), .ZN(n8682) );
  XNOR2_X1 U10070 ( .A(n10136), .B(n10128), .ZN(n13556) );
  NAND3_X1 U10071 ( .A1(n10267), .A2(n10265), .A3(n10266), .ZN(P3_U3204) );
  NAND2_X1 U10072 ( .A1(n9910), .A2(n9909), .ZN(n9926) );
  NAND2_X1 U10073 ( .A1(n9907), .A2(n9906), .ZN(n9910) );
  NAND2_X1 U10074 ( .A1(n7186), .A2(n7185), .ZN(n12691) );
  OAI21_X2 U10075 ( .B1(n10347), .B2(P2_DATAO_REG_4__SCAN_IN), .A(n7182), .ZN(
        n7942) );
  NAND2_X1 U10076 ( .A1(n12789), .A2(n12743), .ZN(n7183) );
  NAND2_X1 U10077 ( .A1(n12677), .A2(n12676), .ZN(n7481) );
  NAND2_X1 U10078 ( .A1(n11656), .A2(n13111), .ZN(n12390) );
  INV_X2 U10079 ( .A(n9663), .ZN(n12964) );
  NOR2_X1 U10080 ( .A1(n12541), .A2(n7197), .ZN(n7196) );
  NAND2_X1 U10081 ( .A1(n7895), .A2(n7204), .ZN(n11248) );
  NAND2_X1 U10082 ( .A1(n11248), .A2(n10110), .ZN(n11280) );
  NAND3_X1 U10083 ( .A1(n7208), .A2(n7213), .A3(n11121), .ZN(n7212) );
  OAI21_X1 U10084 ( .B1(n10116), .B2(n7223), .A(n7222), .ZN(n12273) );
  NAND2_X1 U10085 ( .A1(n10116), .A2(n10115), .ZN(n12195) );
  NAND2_X1 U10086 ( .A1(n10115), .A2(n6628), .ZN(n7228) );
  NAND3_X1 U10087 ( .A1(n9732), .A2(n7236), .A3(n9664), .ZN(n9762) );
  NAND2_X1 U10088 ( .A1(n9846), .A2(n7238), .ZN(n9896) );
  NAND2_X1 U10089 ( .A1(n9915), .A2(n6718), .ZN(n9962) );
  NAND2_X1 U10090 ( .A1(n9915), .A2(n9914), .ZN(n9933) );
  NAND3_X1 U10091 ( .A1(n8754), .A2(n8755), .A3(n8764), .ZN(n8757) );
  NAND2_X1 U10092 ( .A1(n7248), .A2(n12577), .ZN(n15368) );
  AOI21_X1 U10093 ( .B1(n15367), .B2(n7246), .A(n6609), .ZN(n7245) );
  INV_X1 U10094 ( .A(n15367), .ZN(n7247) );
  NAND2_X1 U10095 ( .A1(n11722), .A2(n12753), .ZN(n7248) );
  NAND2_X1 U10096 ( .A1(n14854), .A2(n14853), .ZN(n14852) );
  OAI21_X1 U10097 ( .B1(n14854), .B2(n7254), .A(n7251), .ZN(n7258) );
  OAI21_X1 U10098 ( .B1(n13807), .B2(n13808), .A(n6576), .ZN(n7275) );
  AOI21_X1 U10099 ( .B1(n13807), .B2(n13808), .A(n7277), .ZN(n7276) );
  INV_X1 U10100 ( .A(n13806), .ZN(n7277) );
  NAND3_X1 U10101 ( .A1(n13840), .A2(n13839), .A3(n7280), .ZN(n7278) );
  NAND2_X1 U10102 ( .A1(n7278), .A2(n7279), .ZN(n7733) );
  NAND2_X1 U10103 ( .A1(n7728), .A2(n7283), .ZN(n7284) );
  NAND2_X1 U10104 ( .A1(n7284), .A2(n7285), .ZN(n13827) );
  NAND2_X1 U10105 ( .A1(n7724), .A2(n7289), .ZN(n7288) );
  NAND2_X1 U10106 ( .A1(n7288), .A2(n7290), .ZN(n13865) );
  OAI21_X2 U10107 ( .B1(n7293), .B2(n7292), .A(n13897), .ZN(n13949) );
  INV_X2 U10108 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7297) );
  NAND2_X1 U10109 ( .A1(n8131), .A2(n7945), .ZN(n7305) );
  NAND3_X1 U10110 ( .A1(n7682), .A2(n7683), .A3(n14973), .ZN(n14972) );
  NAND2_X1 U10111 ( .A1(n7684), .A2(n7309), .ZN(n7682) );
  NAND2_X1 U10112 ( .A1(n14849), .A2(n6680), .ZN(n12986) );
  NAND3_X1 U10113 ( .A1(n9380), .A2(n9367), .A3(n9366), .ZN(n9476) );
  NAND3_X1 U10114 ( .A1(n7318), .A2(n6673), .A3(n7315), .ZN(P3_U3200) );
  OAI211_X4 U10115 ( .C1(n6540), .C2(n10429), .A(n7841), .B(n7842), .ZN(n13745) );
  NAND2_X1 U10116 ( .A1(n7781), .A2(n7332), .ZN(n7328) );
  NAND2_X1 U10117 ( .A1(n14201), .A2(n7930), .ZN(n7345) );
  XNOR2_X1 U10118 ( .A(n8053), .B(n8041), .ZN(n8869) );
  XNOR2_X1 U10119 ( .A(n8054), .B(SI_1_), .ZN(n8041) );
  MUX2_X1 U10120 ( .A(n10428), .B(n10368), .S(n7350), .Z(n8054) );
  MUX2_X1 U10121 ( .A(n15952), .B(P2_REG1_REG_1__SCAN_IN), .S(n10498), .Z(
        n15501) );
  XNOR2_X2 U10122 ( .A(n8042), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10498) );
  OAI21_X1 U10123 ( .B1(n10936), .B2(n7359), .A(n7358), .ZN(n7370) );
  NAND2_X1 U10124 ( .A1(n7374), .A2(n7375), .ZN(n10738) );
  NAND2_X1 U10125 ( .A1(n10708), .A2(n6694), .ZN(n7374) );
  OAI21_X1 U10126 ( .B1(P3_IR_REG_31__SCAN_IN), .B2(P3_IR_REG_1__SCAN_IN), .A(
        n7387), .ZN(n7476) );
  NAND3_X1 U10127 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), 
        .A3(P3_IR_REG_0__SCAN_IN), .ZN(n7387) );
  NAND3_X1 U10128 ( .A1(n7392), .A2(n10337), .A3(n7391), .ZN(n7390) );
  INV_X1 U10129 ( .A(n7395), .ZN(n10868) );
  INV_X1 U10130 ( .A(n10869), .ZN(n7392) );
  NAND2_X1 U10131 ( .A1(n10326), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7394) );
  NAND2_X1 U10132 ( .A1(n7400), .A2(n7401), .ZN(n7397) );
  INV_X1 U10133 ( .A(n13166), .ZN(n7411) );
  NOR2_X1 U10134 ( .A1(n11480), .A2(n15928), .ZN(n7413) );
  NAND3_X1 U10135 ( .A1(n7416), .A2(n9466), .A3(n7415), .ZN(n9469) );
  INV_X1 U10136 ( .A(n13268), .ZN(n7414) );
  NAND2_X1 U10137 ( .A1(n7419), .A2(n13268), .ZN(n13252) );
  NAND2_X1 U10138 ( .A1(n7415), .A2(n7416), .ZN(n13271) );
  NAND4_X1 U10139 ( .A1(n9503), .A2(n10970), .A3(n7425), .A4(
        P3_REG1_REG_3__SCAN_IN), .ZN(n7421) );
  NAND2_X1 U10140 ( .A1(n7424), .A2(n9503), .ZN(n13131) );
  AND2_X1 U10141 ( .A1(n9503), .A2(n10970), .ZN(n13132) );
  INV_X1 U10142 ( .A(n10971), .ZN(n7425) );
  OR2_X1 U10143 ( .A1(n9511), .A2(n7443), .ZN(n7431) );
  NAND2_X1 U10144 ( .A1(n9511), .A2(n7435), .ZN(n7433) );
  NAND2_X1 U10145 ( .A1(n9511), .A2(n13174), .ZN(n13176) );
  MUX2_X1 U10146 ( .A(n15418), .B(n12570), .S(n12571), .Z(n12572) );
  NOR2_X1 U10147 ( .A1(n7448), .A2(n10358), .ZN(n7447) );
  NAND2_X1 U10148 ( .A1(n7452), .A2(n7451), .ZN(n13155) );
  INV_X1 U10149 ( .A(n7450), .ZN(n9506) );
  NAND2_X1 U10150 ( .A1(n12691), .A2(n12692), .ZN(n12690) );
  NAND2_X1 U10151 ( .A1(n8803), .A2(n6692), .ZN(n9100) );
  NAND2_X1 U10152 ( .A1(n7478), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9063) );
  AND2_X1 U10153 ( .A1(n9046), .A2(n7478), .ZN(n14768) );
  INV_X1 U10154 ( .A(n10388), .ZN(n7487) );
  NAND2_X1 U10155 ( .A1(n7493), .A2(n11763), .ZN(n12096) );
  NAND2_X1 U10156 ( .A1(n7489), .A2(n11763), .ZN(n7488) );
  NAND2_X1 U10157 ( .A1(n7494), .A2(n7490), .ZN(n7489) );
  INV_X1 U10158 ( .A(n7494), .ZN(n7492) );
  INV_X1 U10159 ( .A(n11767), .ZN(n7495) );
  NAND2_X1 U10160 ( .A1(n7496), .A2(n11767), .ZN(n12095) );
  OAI21_X1 U10161 ( .B1(n15304), .B2(n6652), .A(n7502), .ZN(n15315) );
  NAND2_X1 U10162 ( .A1(n15304), .A2(n7502), .ZN(n7499) );
  NAND2_X1 U10163 ( .A1(n7505), .A2(n15252), .ZN(n15259) );
  NAND2_X1 U10164 ( .A1(n12878), .A2(n7519), .ZN(n7515) );
  OAI211_X1 U10165 ( .C1(n12878), .C2(n7520), .A(n7515), .B(n7516), .ZN(n12892) );
  NAND2_X1 U10166 ( .A1(n12878), .A2(n7531), .ZN(n7522) );
  NAND2_X1 U10167 ( .A1(n12878), .A2(n12877), .ZN(n13087) );
  INV_X1 U10168 ( .A(n12881), .ZN(n7533) );
  NOR2_X1 U10169 ( .A1(n9923), .A2(n13430), .ZN(n7544) );
  INV_X1 U10170 ( .A(n12262), .ZN(n7553) );
  OAI21_X1 U10171 ( .B1(n13018), .B2(n7558), .A(n7554), .ZN(n13027) );
  OR2_X2 U10172 ( .A1(n13018), .A2(n13019), .ZN(n13016) );
  NAND4_X1 U10173 ( .A1(n7562), .A2(n9357), .A3(n7560), .A4(n9383), .ZN(n9461)
         );
  NAND3_X1 U10174 ( .A1(n9470), .A2(n7570), .A3(n7569), .ZN(n7568) );
  NAND2_X1 U10175 ( .A1(n9364), .A2(n9372), .ZN(n9374) );
  INV_X1 U10176 ( .A(n7995), .ZN(n7576) );
  NAND2_X1 U10177 ( .A1(n7576), .A2(SI_24_), .ZN(n7577) );
  NAND3_X1 U10178 ( .A1(n7577), .A2(n7578), .A3(n7580), .ZN(n7998) );
  NAND3_X1 U10179 ( .A1(n7580), .A2(n7579), .A3(n7577), .ZN(n8407) );
  NAND2_X1 U10180 ( .A1(n7598), .A2(n7599), .ZN(n9598) );
  NAND3_X1 U10181 ( .A1(n8559), .A2(n7600), .A3(n8558), .ZN(n7598) );
  NAND2_X1 U10182 ( .A1(n8559), .A2(n8558), .ZN(n9590) );
  NAND3_X1 U10183 ( .A1(n8559), .A2(n8558), .A3(n7603), .ZN(n7601) );
  INV_X1 U10184 ( .A(n7605), .ZN(n7604) );
  NAND2_X1 U10185 ( .A1(n7606), .A2(n8868), .ZN(n8956) );
  NAND3_X1 U10186 ( .A1(n7608), .A2(n7607), .A3(n6685), .ZN(n11536) );
  NAND3_X1 U10187 ( .A1(n11078), .A2(n7609), .A3(n6713), .ZN(n7607) );
  INV_X1 U10188 ( .A(n8524), .ZN(n7618) );
  NAND2_X1 U10189 ( .A1(n14228), .A2(n6552), .ZN(n7648) );
  NAND2_X1 U10190 ( .A1(n7648), .A2(n7649), .ZN(n14199) );
  OR2_X1 U10191 ( .A1(n8872), .A2(n10368), .ZN(n8873) );
  NAND2_X2 U10192 ( .A1(n8832), .A2(n9647), .ZN(n8872) );
  NAND2_X1 U10193 ( .A1(n6658), .A2(n7653), .ZN(n14819) );
  OAI21_X1 U10194 ( .B1(n11683), .B2(n11705), .A(n7672), .ZN(n11732) );
  MUX2_X1 U10195 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15239), .S(n8832), .Z(n12038)
         );
  NAND2_X1 U10196 ( .A1(n7689), .A2(n12941), .ZN(n14994) );
  INV_X1 U10197 ( .A(n12943), .ZN(n7688) );
  OAI21_X1 U10198 ( .B1(n9975), .B2(n7695), .A(n7693), .ZN(n10020) );
  NOR2_X1 U10199 ( .A1(n13449), .A2(n6674), .ZN(n13498) );
  NAND2_X1 U10200 ( .A1(n7708), .A2(n13398), .ZN(n7707) );
  NAND2_X1 U10201 ( .A1(n13309), .A2(n13312), .ZN(n7709) );
  NAND2_X1 U10202 ( .A1(n9822), .A2(n7712), .ZN(n7711) );
  NAND2_X1 U10203 ( .A1(n7711), .A2(n7713), .ZN(n9871) );
  NAND3_X1 U10204 ( .A1(n13852), .A2(n13851), .A3(n6691), .ZN(n7724) );
  NAND3_X1 U10205 ( .A1(n13818), .A2(n13817), .A3(n6690), .ZN(n7728) );
  NAND2_X1 U10206 ( .A1(n7730), .A2(n7731), .ZN(n13835) );
  NAND3_X1 U10207 ( .A1(n13830), .A2(n6697), .A3(n13829), .ZN(n7730) );
  NAND2_X1 U10208 ( .A1(n7733), .A2(n7734), .ZN(n13847) );
  NAND2_X1 U10209 ( .A1(n7744), .A2(n12438), .ZN(n12222) );
  NAND2_X1 U10210 ( .A1(n7758), .A2(n7759), .ZN(n11057) );
  NAND2_X1 U10211 ( .A1(n12483), .A2(n12371), .ZN(n7763) );
  NAND2_X1 U10212 ( .A1(n11039), .A2(n12371), .ZN(n11027) );
  NAND2_X1 U10213 ( .A1(n11037), .A2(n11036), .ZN(n11039) );
  NAND2_X1 U10214 ( .A1(n11596), .A2(n7767), .ZN(n7765) );
  NAND2_X1 U10215 ( .A1(n6855), .A2(n7785), .ZN(n8452) );
  NAND2_X1 U10216 ( .A1(n7786), .A2(n8265), .ZN(n8282) );
  OAI21_X1 U10217 ( .B1(n8618), .B2(n7791), .A(n7790), .ZN(n11776) );
  AOI21_X1 U10218 ( .B1(n7790), .B2(n7791), .A(n7789), .ZN(n7788) );
  NAND2_X1 U10219 ( .A1(n7804), .A2(n7802), .ZN(n13560) );
  AND2_X1 U10220 ( .A1(n7804), .A2(n7803), .ZN(n13562) );
  NAND2_X1 U10221 ( .A1(n12064), .A2(n7810), .ZN(n7809) );
  NAND2_X1 U10222 ( .A1(n7809), .A2(n7811), .ZN(n11706) );
  OAI21_X1 U10223 ( .B1(n15014), .B2(n12911), .A(n12912), .ZN(n14997) );
  NAND2_X1 U10224 ( .A1(n14995), .A2(n7824), .ZN(n7823) );
  NAND2_X1 U10225 ( .A1(n14864), .A2(n14910), .ZN(n14904) );
  INV_X1 U10226 ( .A(n8832), .ZN(n7833) );
  NOR2_X1 U10227 ( .A1(n7833), .A2(n7834), .ZN(n7832) );
  INV_X2 U10228 ( .A(n8872), .ZN(n9175) );
  AND2_X1 U10229 ( .A1(n14872), .A2(n7837), .ZN(n15197) );
  OAI21_X1 U10230 ( .B1(n14872), .B2(n7301), .A(n7835), .ZN(P1_U3553) );
  NAND2_X1 U10231 ( .A1(n8048), .A2(n6669), .ZN(n7842) );
  INV_X1 U10232 ( .A(n7845), .ZN(n11871) );
  NAND2_X1 U10233 ( .A1(n9230), .A2(n9229), .ZN(n7872) );
  NAND2_X1 U10234 ( .A1(n9195), .A2(n9196), .ZN(n7884) );
  NAND2_X1 U10235 ( .A1(n12363), .A2(n12368), .ZN(n7887) );
  NAND2_X1 U10236 ( .A1(n12366), .A2(n12487), .ZN(n7885) );
  XNOR2_X1 U10237 ( .A(n7886), .B(n12487), .ZN(n15678) );
  INV_X1 U10238 ( .A(n12365), .ZN(n7886) );
  NOR2_X1 U10239 ( .A1(n12365), .A2(n12487), .ZN(n7888) );
  OR2_X1 U10240 ( .A1(n7898), .A2(n7897), .ZN(n7896) );
  NAND2_X1 U10241 ( .A1(n6683), .A2(n13308), .ZN(n13298) );
  NAND2_X1 U10242 ( .A1(n8531), .A2(n8530), .ZN(n14183) );
  XNOR2_X1 U10243 ( .A(n8553), .B(n8003), .ZN(n14477) );
  NAND2_X1 U10244 ( .A1(n10541), .A2(n13756), .ZN(n11233) );
  OR2_X1 U10245 ( .A1(n15156), .A2(n15015), .ZN(n14978) );
  AND2_X1 U10246 ( .A1(n14151), .A2(n14150), .ZN(n14185) );
  NAND2_X1 U10247 ( .A1(n11686), .A2(n11685), .ZN(n11722) );
  XNOR2_X1 U10248 ( .A(n15083), .B(n12928), .ZN(n12932) );
  INV_X1 U10249 ( .A(n12832), .ZN(n9613) );
  INV_X1 U10250 ( .A(n12520), .ZN(n12523) );
  OR2_X1 U10251 ( .A1(n14128), .A2(n14127), .ZN(n14336) );
  AND2_X4 U10252 ( .A1(n15224), .A2(n8793), .ZN(n8947) );
  OR2_X1 U10253 ( .A1(n8958), .A2(n12036), .ZN(n8858) );
  NAND2_X1 U10254 ( .A1(n9310), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8867) );
  NAND2_X1 U10255 ( .A1(n14509), .A2(n14508), .ZN(n14507) );
  XNOR2_X2 U10256 ( .A(n13977), .B(n13726), .ZN(n13907) );
  NAND2_X4 U10257 ( .A1(n8122), .A2(n8121), .ZN(n13726) );
  OAI211_X4 U10258 ( .C1(n9606), .C2(n9633), .A(n8066), .B(n8065), .ZN(n13741)
         );
  AND2_X2 U10259 ( .A1(n10262), .A2(n15681), .ZN(n15688) );
  AND2_X1 U10260 ( .A1(n13077), .A2(n13413), .ZN(n7903) );
  OR2_X1 U10261 ( .A1(n14365), .A2(n8529), .ZN(n7904) );
  INV_X1 U10262 ( .A(n14088), .ZN(n8543) );
  AND2_X1 U10263 ( .A1(n10577), .A2(n10576), .ZN(n15355) );
  AND2_X1 U10264 ( .A1(n10379), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7906) );
  AND2_X1 U10265 ( .A1(n14322), .A2(n15651), .ZN(n7907) );
  AND2_X1 U10266 ( .A1(n14322), .A2(n13962), .ZN(n7908) );
  NOR2_X1 U10267 ( .A1(n11990), .A2(n11989), .ZN(n7909) );
  AND2_X1 U10268 ( .A1(n9329), .A2(n14621), .ZN(n7910) );
  NOR2_X1 U10269 ( .A1(n11987), .A2(n11932), .ZN(n7912) );
  AND3_X1 U10270 ( .A1(n6676), .A2(n13890), .A3(n13885), .ZN(n7913) );
  AND2_X1 U10271 ( .A1(n8739), .A2(n8738), .ZN(n7914) );
  OR2_X1 U10272 ( .A1(n9803), .A2(n12242), .ZN(n7915) );
  INV_X1 U10273 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9370) );
  AND2_X1 U10274 ( .A1(n15233), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7917) );
  AND3_X1 U10275 ( .A1(n9735), .A2(n9734), .A3(n9733), .ZN(n7918) );
  AND2_X1 U10276 ( .A1(n9759), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U10277 ( .A1(n10220), .A2(n12266), .ZN(n7920) );
  AND2_X2 U10278 ( .A1(n9474), .A2(n10088), .ZN(n13396) );
  OR2_X1 U10279 ( .A1(n14047), .A2(n14118), .ZN(n7921) );
  INV_X1 U10280 ( .A(n10329), .ZN(n9411) );
  INV_X1 U10281 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9410) );
  INV_X1 U10282 ( .A(n14043), .ZN(n12830) );
  AND2_X1 U10283 ( .A1(n12377), .A2(n12380), .ZN(n7922) );
  INV_X1 U10284 ( .A(n14459), .ZN(n9618) );
  INV_X1 U10285 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8266) );
  INV_X1 U10286 ( .A(n9476), .ZN(n9478) );
  AND3_X1 U10287 ( .A1(n12674), .A2(n12673), .A3(n12914), .ZN(n7923) );
  OR2_X1 U10288 ( .A1(n12774), .A2(n12775), .ZN(n7924) );
  AND2_X1 U10289 ( .A1(n8134), .A2(n8136), .ZN(n7925) );
  AND3_X1 U10290 ( .A1(n8740), .A2(n8713), .A3(n13711), .ZN(n7926) );
  INV_X1 U10291 ( .A(n12956), .ZN(n12928) );
  AND2_X1 U10292 ( .A1(n9655), .A2(n9657), .ZN(n7927) );
  INV_X1 U10293 ( .A(n13101), .ZN(n13432) );
  INV_X1 U10294 ( .A(n12422), .ZN(n10221) );
  INV_X1 U10295 ( .A(n13872), .ZN(n14317) );
  AND2_X1 U10296 ( .A1(n8372), .A2(n14154), .ZN(n7930) );
  OR2_X1 U10297 ( .A1(n13035), .A2(n12275), .ZN(n7931) );
  AND2_X1 U10298 ( .A1(n8182), .A2(n8167), .ZN(n7932) );
  NOR2_X1 U10299 ( .A1(n11971), .A2(n11970), .ZN(n7933) );
  AND2_X1 U10300 ( .A1(n12765), .A2(n11994), .ZN(n7934) );
  AND2_X1 U10301 ( .A1(n13732), .A2(n13731), .ZN(n13774) );
  AND2_X1 U10302 ( .A1(n13914), .A2(n13785), .ZN(n13786) );
  INV_X1 U10303 ( .A(n12687), .ZN(n12688) );
  NAND2_X1 U10304 ( .A1(n12694), .A2(n12693), .ZN(n12695) );
  NOR2_X1 U10305 ( .A1(n12863), .A2(n13022), .ZN(n12859) );
  NAND2_X1 U10306 ( .A1(n11026), .A2(n11064), .ZN(n10104) );
  AND2_X1 U10307 ( .A1(n15811), .A2(n9486), .ZN(n9488) );
  OAI21_X1 U10308 ( .B1(n14536), .B2(n14534), .A(n9158), .ZN(n9156) );
  NOR2_X1 U10309 ( .A1(n12041), .A2(n11693), .ZN(n12562) );
  NOR2_X1 U10310 ( .A1(n12860), .A2(n12859), .ZN(n12861) );
  NAND2_X1 U10311 ( .A1(n13117), .A2(n11357), .ZN(n12363) );
  NAND3_X1 U10312 ( .A1(n9408), .A2(n9356), .A3(n9355), .ZN(n9492) );
  INV_X1 U10313 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9462) );
  INV_X1 U10314 ( .A(n13384), .ZN(n9989) );
  NOR2_X1 U10315 ( .A1(n9411), .A2(n9410), .ZN(n9412) );
  OAI21_X1 U10316 ( .B1(n13582), .B2(n13966), .A(n13579), .ZN(n8678) );
  NAND2_X1 U10317 ( .A1(n13895), .A2(n13894), .ZN(n13896) );
  INV_X1 U10318 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8075) );
  INV_X1 U10319 ( .A(n12984), .ZN(n12985) );
  AOI21_X1 U10320 ( .B1(n11973), .B2(n11972), .A(n7933), .ZN(n12110) );
  AND2_X1 U10321 ( .A1(n8853), .A2(n9333), .ZN(n9343) );
  AND2_X1 U10322 ( .A1(n9834), .A2(n12248), .ZN(n9835) );
  INV_X1 U10323 ( .A(n9746), .ZN(n10176) );
  INV_X1 U10324 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n9826) );
  AND2_X1 U10325 ( .A1(n12516), .A2(n12346), .ZN(n12510) );
  INV_X1 U10326 ( .A(n13411), .ZN(n10120) );
  INV_X1 U10327 ( .A(n9387), .ZN(n9364) );
  INV_X1 U10328 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9391) );
  OAI21_X1 U10329 ( .B1(n14040), .B2(n13725), .A(n8736), .ZN(n8737) );
  INV_X1 U10330 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8323) );
  NOR2_X1 U10331 ( .A1(n7913), .A2(n13896), .ZN(n13897) );
  AND2_X1 U10332 ( .A1(n8025), .A2(n8459), .ZN(n14080) );
  INV_X1 U10333 ( .A(n13903), .ZN(n12004) );
  INV_X1 U10334 ( .A(n10541), .ZN(n11232) );
  OR2_X1 U10335 ( .A1(n8301), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8303) );
  NAND2_X1 U10336 ( .A1(n9210), .A2(n9211), .ZN(n9212) );
  AND2_X1 U10337 ( .A1(n14571), .A2(n15029), .ZN(n14600) );
  OR2_X1 U10338 ( .A1(n11452), .A2(n11453), .ZN(n11804) );
  XNOR2_X1 U10339 ( .A(n14650), .B(n15399), .ZN(n15386) );
  NAND2_X1 U10340 ( .A1(n8553), .A2(n15772), .ZN(n8554) );
  INV_X1 U10341 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8765) );
  INV_X1 U10342 ( .A(n13342), .ZN(n12996) );
  INV_X1 U10343 ( .A(n13397), .ZN(n13022) );
  INV_X1 U10344 ( .A(n13103), .ZN(n13039) );
  OR2_X1 U10345 ( .A1(n9738), .A2(n11403), .ZN(n9739) );
  INV_X1 U10346 ( .A(n13114), .ZN(n11403) );
  INV_X1 U10347 ( .A(n13353), .ZN(n13094) );
  NOR2_X1 U10348 ( .A1(n10232), .A2(n10070), .ZN(n10090) );
  AND2_X1 U10349 ( .A1(n9939), .A2(n9938), .ZN(n13413) );
  NAND2_X1 U10350 ( .A1(n10845), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n13140) );
  INV_X1 U10351 ( .A(n13102), .ZN(n13430) );
  AND2_X1 U10352 ( .A1(n10213), .A2(n10212), .ZN(n10252) );
  AND2_X1 U10353 ( .A1(n10207), .A2(n12525), .ZN(n13428) );
  AND2_X1 U10354 ( .A1(n10234), .A2(n10233), .ZN(n13313) );
  NAND2_X1 U10355 ( .A1(n9652), .A2(n7927), .ZN(n9661) );
  NOR2_X1 U10356 ( .A1(n9478), .A2(n9368), .ZN(n9369) );
  AND2_X1 U10357 ( .A1(n9992), .A2(n9973), .ZN(n9974) );
  AND2_X1 U10358 ( .A1(n9925), .A2(n9908), .ZN(n9909) );
  NAND2_X1 U10359 ( .A1(n9390), .A2(n9408), .ZN(n9413) );
  INV_X1 U10360 ( .A(n8737), .ZN(n8738) );
  INV_X1 U10361 ( .A(n10887), .ZN(n8601) );
  OR2_X1 U10362 ( .A1(n13703), .A2(n14116), .ZN(n13587) );
  INV_X1 U10363 ( .A(n13966), .ZN(n13665) );
  INV_X1 U10364 ( .A(n13970), .ZN(n14153) );
  INV_X1 U10365 ( .A(n13977), .ZN(n11597) );
  AND2_X1 U10366 ( .A1(n13959), .A2(n9616), .ZN(n14318) );
  INV_X1 U10367 ( .A(n14269), .ZN(n13574) );
  INV_X1 U10368 ( .A(n14591), .ZN(n14613) );
  INV_X1 U10369 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14714) );
  OR2_X1 U10370 ( .A1(n10672), .A2(n10671), .ZN(n14762) );
  OR2_X1 U10371 ( .A1(n10859), .A2(n10860), .ZN(n10861) );
  INV_X1 U10372 ( .A(n15064), .ZN(n14818) );
  NAND2_X1 U10373 ( .A1(n14635), .A2(n15031), .ZN(n12929) );
  INV_X1 U10374 ( .A(n15031), .ZN(n14943) );
  OR2_X1 U10375 ( .A1(n9334), .A2(n10567), .ZN(n10777) );
  AND2_X1 U10376 ( .A1(n11697), .A2(n12558), .ZN(n12720) );
  INV_X1 U10377 ( .A(n12758), .ZN(n11989) );
  NAND2_X1 U10378 ( .A1(n15377), .A2(n14809), .ZN(n11665) );
  XNOR2_X1 U10379 ( .A(n8350), .B(n8349), .ZN(n8831) );
  XNOR2_X1 U10380 ( .A(n7962), .B(SI_13_), .ZN(n8249) );
  INV_X1 U10381 ( .A(n12102), .ZN(n12100) );
  INV_X1 U10382 ( .A(n13072), .ZN(n13089) );
  INV_X1 U10383 ( .A(n12275), .ZN(n13049) );
  AND2_X1 U10384 ( .A1(n9581), .A2(n9580), .ZN(n15694) );
  AND2_X1 U10385 ( .A1(n9579), .A2(n9578), .ZN(n13261) );
  INV_X1 U10386 ( .A(n13261), .ZN(n13279) );
  AND2_X1 U10387 ( .A1(P3_U3897), .A2(n13548), .ZN(n13248) );
  INV_X1 U10388 ( .A(n15681), .ZN(n15675) );
  AND2_X1 U10389 ( .A1(n11283), .A2(n11282), .ZN(n11372) );
  NAND2_X1 U10390 ( .A1(n12431), .A2(n12425), .ZN(n12422) );
  INV_X1 U10391 ( .A(n13536), .ZN(n13520) );
  NAND2_X1 U10392 ( .A1(n13313), .A2(n11359), .ZN(n13474) );
  INV_X1 U10393 ( .A(n10048), .ZN(n10341) );
  OAI211_X1 U10394 ( .C1(n9373), .C2(n9372), .A(n9374), .B(n9371), .ZN(n9621)
         );
  AND2_X1 U10395 ( .A1(n9957), .A2(n9943), .ZN(n9955) );
  AND2_X1 U10396 ( .A1(n8726), .A2(n8708), .ZN(n13711) );
  INV_X1 U10397 ( .A(n13944), .ZN(n13954) );
  AND2_X1 U10398 ( .A1(n8036), .A2(n8035), .ZN(n14064) );
  INV_X1 U10399 ( .A(n8721), .ZN(n8461) );
  NAND2_X2 U10400 ( .A1(n13750), .A2(n8046), .ZN(n10541) );
  AND2_X1 U10401 ( .A1(n10491), .A2(n13953), .ZN(n15596) );
  OR2_X1 U10402 ( .A1(n10486), .A2(n10485), .ZN(n10495) );
  NAND2_X1 U10403 ( .A1(n14050), .A2(n14049), .ZN(n14325) );
  INV_X1 U10404 ( .A(n14275), .ZN(n14295) );
  INV_X1 U10405 ( .A(n14116), .ZN(n14302) );
  NAND2_X2 U10406 ( .A1(n11230), .A2(n14290), .ZN(n14293) );
  INV_X1 U10407 ( .A(n15614), .ZN(n8705) );
  INV_X1 U10408 ( .A(n14461), .ZN(n8549) );
  AND2_X1 U10409 ( .A1(n15642), .A2(n15636), .ZN(n15655) );
  AND2_X1 U10410 ( .A1(n8486), .A2(n14476), .ZN(n15610) );
  AND2_X1 U10411 ( .A1(n10281), .A2(n11490), .ZN(n8730) );
  NOR2_X1 U10412 ( .A1(n10777), .A2(n10574), .ZN(n14571) );
  NOR2_X2 U10413 ( .A1(n11923), .A2(n15471), .ZN(n14617) );
  OR2_X1 U10414 ( .A1(n12973), .A2(n9336), .ZN(n9342) );
  INV_X1 U10415 ( .A(n14804), .ZN(n15340) );
  INV_X1 U10416 ( .A(n14805), .ZN(n15338) );
  NAND2_X1 U10417 ( .A1(n12930), .A2(n12929), .ZN(n12931) );
  INV_X1 U10418 ( .A(n15405), .ZN(n15005) );
  INV_X1 U10419 ( .A(n10777), .ZN(n10779) );
  INV_X1 U10420 ( .A(n14829), .ZN(n15068) );
  INV_X1 U10421 ( .A(n15476), .ZN(n15456) );
  NAND2_X1 U10422 ( .A1(n15447), .A2(n15446), .ZN(n15476) );
  NAND2_X1 U10423 ( .A1(n9288), .A2(n9287), .ZN(n10569) );
  INV_X1 U10424 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U10425 ( .A1(n10062), .A2(n10242), .ZN(n13098) );
  INV_X1 U10426 ( .A(n13248), .ZN(n13277) );
  OR2_X1 U10427 ( .A1(n9516), .A2(n9573), .ZN(n13242) );
  NAND2_X1 U10428 ( .A1(n9577), .A2(n9498), .ZN(n13288) );
  NAND2_X1 U10429 ( .A1(n13405), .A2(n10259), .ZN(n13441) );
  INV_X1 U10430 ( .A(n11395), .ZN(n11220) );
  OR2_X1 U10431 ( .A1(n13478), .A2(n11358), .ZN(n13482) );
  AND2_X1 U10432 ( .A1(n11323), .A2(n11322), .ZN(n11500) );
  INV_X2 U10433 ( .A(n15693), .ZN(n15691) );
  OR2_X1 U10434 ( .A1(n15693), .A2(n11358), .ZN(n13536) );
  INV_X1 U10435 ( .A(SI_13_), .ZN(n10480) );
  INV_X1 U10436 ( .A(n10924), .ZN(n10362) );
  INV_X1 U10437 ( .A(n14109), .ZN(n14418) );
  INV_X1 U10438 ( .A(n13711), .ZN(n13695) );
  NAND2_X1 U10439 ( .A1(n10539), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13717) );
  INV_X1 U10440 ( .A(n14065), .ZN(n13962) );
  NAND2_X1 U10441 ( .A1(n8433), .A2(n8432), .ZN(n13966) );
  INV_X1 U10442 ( .A(n15595), .ZN(n15584) );
  INV_X1 U10443 ( .A(n15596), .ZN(n15586) );
  OR2_X1 U10444 ( .A1(n10495), .A2(P2_U3088), .ZN(n15609) );
  NAND2_X1 U10445 ( .A1(n14293), .A2(n11529), .ZN(n14275) );
  NAND2_X1 U10446 ( .A1(n14293), .A2(n11515), .ZN(n14279) );
  NAND2_X1 U10447 ( .A1(n15670), .A2(n15651), .ZN(n14400) );
  NAND2_X1 U10448 ( .A1(n8546), .A2(n8705), .ZN(n15667) );
  NAND2_X1 U10449 ( .A1(n8543), .A2(n8549), .ZN(n8550) );
  NAND2_X1 U10450 ( .A1(n15659), .A2(n15651), .ZN(n14459) );
  NAND2_X1 U10451 ( .A1(n8546), .A2(n15614), .ZN(n15657) );
  INV_X1 U10452 ( .A(n15612), .ZN(n15611) );
  NOR2_X1 U10453 ( .A1(n15617), .A2(n15610), .ZN(n15612) );
  INV_X1 U10454 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11316) );
  INV_X1 U10455 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10461) );
  INV_X1 U10456 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10434) );
  NAND3_X1 U10457 ( .A1(n11663), .A2(n9307), .A3(n9306), .ZN(n14619) );
  OR2_X1 U10458 ( .A1(n10617), .A2(n14664), .ZN(n14804) );
  OR2_X1 U10459 ( .A1(n12971), .A2(n14809), .ZN(n14935) );
  OR2_X1 U10460 ( .A1(n15405), .A2(n11668), .ZN(n15060) );
  INV_X1 U10461 ( .A(n15478), .ZN(n15477) );
  INV_X1 U10462 ( .A(n15407), .ZN(n15406) );
  AND2_X1 U10463 ( .A1(n10468), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10515) );
  INV_X1 U10464 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12319) );
  INV_X1 U10465 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10687) );
  INV_X1 U10466 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10459) );
  AND2_X1 U10467 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10486), .ZN(P2_U3947) );
  NOR2_X1 U10468 ( .A1(n8853), .A2(n10554), .ZN(P1_U4016) );
  INV_X1 U10469 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8503) );
  INV_X1 U10470 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10349) );
  INV_X1 U10471 ( .A(n8062), .ZN(n8081) );
  INV_X1 U10472 ( .A(n8085), .ZN(n7937) );
  INV_X1 U10473 ( .A(SI_3_), .ZN(n10335) );
  NAND2_X1 U10474 ( .A1(n7937), .A2(n10335), .ZN(n7938) );
  OAI21_X1 U10475 ( .B1(n8081), .B2(SI_2_), .A(n7938), .ZN(n8095) );
  INV_X1 U10476 ( .A(SI_2_), .ZN(n10324) );
  NOR2_X1 U10477 ( .A1(n8062), .A2(n10324), .ZN(n7939) );
  INV_X1 U10478 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10352) );
  XNOR2_X1 U10479 ( .A(n7942), .B(SI_4_), .ZN(n7940) );
  INV_X1 U10480 ( .A(n7940), .ZN(n8100) );
  INV_X1 U10481 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U10482 ( .A1(n8041), .A2(n8057), .ZN(n8080) );
  INV_X1 U10483 ( .A(n8054), .ZN(n8058) );
  NAND2_X1 U10484 ( .A1(n8058), .A2(SI_1_), .ZN(n8079) );
  MUX2_X1 U10485 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10347), .Z(n8114) );
  NAND2_X1 U10486 ( .A1(n8114), .A2(SI_5_), .ZN(n8134) );
  INV_X1 U10487 ( .A(n7942), .ZN(n7943) );
  NAND2_X1 U10488 ( .A1(n7943), .A2(SI_4_), .ZN(n8136) );
  INV_X1 U10489 ( .A(n7946), .ZN(n7944) );
  NAND2_X1 U10490 ( .A1(n7944), .A2(SI_6_), .ZN(n8152) );
  NOR2_X1 U10491 ( .A1(n8114), .A2(SI_5_), .ZN(n8137) );
  INV_X1 U10492 ( .A(n8137), .ZN(n8132) );
  MUX2_X1 U10493 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6541), .Z(n7949) );
  XNOR2_X1 U10494 ( .A(n7949), .B(SI_7_), .ZN(n8154) );
  AOI21_X1 U10495 ( .B1(n8149), .B2(n8152), .A(n8154), .ZN(n7947) );
  MUX2_X1 U10496 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10347), .Z(n7950) );
  XNOR2_X1 U10497 ( .A(n7950), .B(SI_9_), .ZN(n8184) );
  MUX2_X1 U10498 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10347), .Z(n8168) );
  NOR2_X1 U10499 ( .A1(n8168), .A2(SI_8_), .ZN(n7948) );
  INV_X1 U10500 ( .A(n8202), .ZN(n7953) );
  NAND2_X1 U10501 ( .A1(n8168), .A2(SI_8_), .ZN(n8182) );
  NAND2_X1 U10502 ( .A1(n7949), .A2(SI_7_), .ZN(n8167) );
  NAND2_X1 U10503 ( .A1(n7950), .A2(SI_9_), .ZN(n8204) );
  MUX2_X1 U10504 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10347), .Z(n8206) );
  NAND2_X1 U10505 ( .A1(n8206), .A2(SI_10_), .ZN(n7951) );
  OAI211_X1 U10506 ( .C1(n7953), .C2(n7932), .A(n8204), .B(n7951), .ZN(n7952)
         );
  INV_X1 U10507 ( .A(n8206), .ZN(n7954) );
  NAND2_X1 U10508 ( .A1(n7954), .A2(n10366), .ZN(n7955) );
  MUX2_X1 U10509 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10347), .Z(n7956) );
  XNOR2_X1 U10510 ( .A(n7956), .B(n15810), .ZN(n8220) );
  INV_X1 U10511 ( .A(n7956), .ZN(n7957) );
  NAND2_X1 U10512 ( .A1(n7957), .A2(n15810), .ZN(n7958) );
  NAND2_X1 U10513 ( .A1(n7959), .A2(n7958), .ZN(n8234) );
  MUX2_X1 U10514 ( .A(n10459), .B(n10461), .S(n9647), .Z(n7960) );
  NAND2_X1 U10515 ( .A1(n7960), .A2(n10438), .ZN(n7961) );
  MUX2_X1 U10516 ( .A(n10465), .B(n10477), .S(n6541), .Z(n7962) );
  NAND2_X1 U10517 ( .A1(n7962), .A2(n10480), .ZN(n7963) );
  MUX2_X1 U10518 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6541), .Z(n8278) );
  INV_X1 U10519 ( .A(n8278), .ZN(n7965) );
  MUX2_X1 U10520 ( .A(n15737), .B(n10736), .S(n10347), .Z(n8280) );
  INV_X1 U10521 ( .A(n8280), .ZN(n7964) );
  NAND2_X1 U10522 ( .A1(n7964), .A2(SI_15_), .ZN(n7968) );
  OAI21_X1 U10523 ( .B1(n7965), .B2(n15956), .A(n7968), .ZN(n7966) );
  INV_X1 U10524 ( .A(n7966), .ZN(n7967) );
  NOR2_X1 U10525 ( .A1(n8278), .A2(SI_14_), .ZN(n7969) );
  INV_X1 U10526 ( .A(SI_15_), .ZN(n10536) );
  AOI22_X1 U10527 ( .A1(n7969), .A2(n7968), .B1(n10536), .B2(n8280), .ZN(n7970) );
  MUX2_X1 U10528 ( .A(n10558), .B(n10565), .S(n9647), .Z(n7971) );
  NAND2_X1 U10529 ( .A1(n7971), .A2(n15925), .ZN(n7972) );
  MUX2_X1 U10530 ( .A(n10687), .B(n10701), .S(n9647), .Z(n8317) );
  NOR2_X1 U10531 ( .A1(n7974), .A2(SI_17_), .ZN(n7973) );
  NAND2_X1 U10532 ( .A1(n7974), .A2(SI_17_), .ZN(n7975) );
  INV_X1 U10533 ( .A(SI_18_), .ZN(n10735) );
  MUX2_X1 U10534 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9647), .Z(n8343) );
  INV_X1 U10535 ( .A(n8343), .ZN(n7976) );
  MUX2_X1 U10536 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9647), .Z(n7977) );
  OAI21_X1 U10537 ( .B1(n10735), .B2(n7976), .A(n8348), .ZN(n7982) );
  NOR2_X1 U10538 ( .A1(n8343), .A2(SI_18_), .ZN(n7980) );
  INV_X1 U10539 ( .A(n7977), .ZN(n7978) );
  NAND2_X1 U10540 ( .A1(n7978), .A2(n10798), .ZN(n8347) );
  INV_X1 U10541 ( .A(n8347), .ZN(n7979) );
  MUX2_X1 U10542 ( .A(n11203), .B(n11316), .S(n9647), .Z(n8363) );
  INV_X1 U10543 ( .A(n8363), .ZN(n8373) );
  MUX2_X1 U10544 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9647), .Z(n8378) );
  INV_X1 U10545 ( .A(n8378), .ZN(n7983) );
  NAND2_X1 U10546 ( .A1(n7983), .A2(n12960), .ZN(n7985) );
  OAI21_X1 U10547 ( .B1(SI_20_), .B2(n8373), .A(n7985), .ZN(n7984) );
  INV_X1 U10548 ( .A(SI_20_), .ZN(n11183) );
  NOR2_X1 U10549 ( .A1(n8363), .A2(n11183), .ZN(n7986) );
  AOI22_X1 U10550 ( .A1(n7986), .A2(n7985), .B1(n8378), .B2(SI_21_), .ZN(n7987) );
  MUX2_X1 U10551 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9647), .Z(n8416) );
  MUX2_X1 U10552 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9647), .Z(n8420) );
  INV_X1 U10553 ( .A(n8420), .ZN(n7989) );
  NAND2_X1 U10554 ( .A1(n7989), .A2(n11731), .ZN(n7992) );
  OAI21_X1 U10555 ( .B1(SI_22_), .B2(n8416), .A(n7992), .ZN(n7990) );
  INV_X1 U10556 ( .A(n7990), .ZN(n7991) );
  INV_X1 U10557 ( .A(n8416), .ZN(n8394) );
  INV_X1 U10558 ( .A(SI_22_), .ZN(n8393) );
  NOR2_X1 U10559 ( .A1(n8394), .A2(n8393), .ZN(n7993) );
  AOI22_X1 U10560 ( .A1(n7993), .A2(n7992), .B1(n8420), .B2(SI_23_), .ZN(n7994) );
  MUX2_X1 U10561 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9647), .Z(n8406) );
  NAND2_X1 U10562 ( .A1(n7996), .A2(SI_24_), .ZN(n7997) );
  MUX2_X1 U10563 ( .A(n11774), .B(n11770), .S(n9647), .Z(n7999) );
  INV_X1 U10564 ( .A(SI_25_), .ZN(n13558) );
  NAND2_X1 U10565 ( .A1(n7999), .A2(n13558), .ZN(n8002) );
  INV_X1 U10566 ( .A(n7999), .ZN(n8000) );
  NAND2_X1 U10567 ( .A1(n8000), .A2(SI_25_), .ZN(n8001) );
  NAND2_X1 U10568 ( .A1(n8002), .A2(n8001), .ZN(n8435) );
  INV_X1 U10569 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15233) );
  MUX2_X1 U10570 ( .A(n15233), .B(n14479), .S(n9647), .Z(n8552) );
  XNOR2_X1 U10571 ( .A(n8552), .B(SI_26_), .ZN(n8003) );
  NAND2_X1 U10572 ( .A1(n8351), .A2(n8007), .ZN(n8008) );
  NOR2_X1 U10573 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8010) );
  NOR2_X1 U10574 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n8009) );
  NAND4_X1 U10575 ( .A1(n8010), .A2(n8009), .A3(n8483), .A4(n8473), .ZN(n8014)
         );
  INV_X1 U10576 ( .A(n8013), .ZN(n8455) );
  INV_X1 U10577 ( .A(n8015), .ZN(n8016) );
  NAND2_X1 U10578 ( .A1(n14477), .A2(n8102), .ZN(n8018) );
  OR2_X1 U10579 ( .A1(n9606), .A2(n14479), .ZN(n8017) );
  NAND2_X1 U10580 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n8019) );
  INV_X1 U10581 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8383) );
  INV_X1 U10582 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8397) );
  INV_X1 U10583 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n15875) );
  INV_X1 U10584 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8023) );
  OAI21_X1 U10585 ( .B1(n8439), .B2(n15875), .A(n8023), .ZN(n8025) );
  NAND2_X1 U10586 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n8024) );
  NAND2_X1 U10587 ( .A1(n14080), .A2(n8721), .ZN(n8036) );
  AND2_X4 U10588 ( .A1(n8029), .A2(n12906), .ZN(n12832) );
  INV_X1 U10589 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8033) );
  AND2_X2 U10590 ( .A1(n12807), .A2(n12906), .ZN(n8386) );
  NAND2_X1 U10591 ( .A1(n9609), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8032) );
  AND2_X2 U10592 ( .A1(n12807), .A2(n8030), .ZN(n8123) );
  NAND2_X1 U10593 ( .A1(n12833), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8031) );
  OAI211_X1 U10594 ( .C1(n9613), .C2(n8033), .A(n8032), .B(n8031), .ZN(n8034)
         );
  INV_X1 U10595 ( .A(n8034), .ZN(n8035) );
  OR2_X1 U10596 ( .A1(n13862), .A2(n14064), .ZN(n12826) );
  NAND2_X1 U10597 ( .A1(n13862), .A2(n14064), .ZN(n14057) );
  NAND2_X1 U10598 ( .A1(n12826), .A2(n14057), .ZN(n13927) );
  NAND2_X1 U10599 ( .A1(n8386), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8040) );
  NAND2_X1 U10600 ( .A1(n12832), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8039) );
  NAND2_X1 U10601 ( .A1(n8068), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U10602 ( .A1(n8123), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8037) );
  INV_X1 U10603 ( .A(n8869), .ZN(n10429) );
  NAND2_X1 U10604 ( .A1(n12832), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U10605 ( .A1(n8123), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8044) );
  NAND2_X1 U10606 ( .A1(n8386), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n13749) );
  NAND2_X1 U10607 ( .A1(n8068), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n13748) );
  AND2_X1 U10608 ( .A1(n13749), .A2(n13748), .ZN(n8046) );
  INV_X1 U10609 ( .A(SI_0_), .ZN(n10346) );
  NOR2_X1 U10610 ( .A1(n10425), .A2(n10346), .ZN(n8047) );
  INV_X1 U10611 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10547) );
  XNOR2_X1 U10612 ( .A(n8047), .B(n10547), .ZN(n14481) );
  MUX2_X1 U10613 ( .A(n15497), .B(n14481), .S(n8048), .Z(n13756) );
  AND2_X1 U10614 ( .A1(n11232), .A2(n13756), .ZN(n10898) );
  INV_X1 U10615 ( .A(n13981), .ZN(n13744) );
  NAND2_X1 U10616 ( .A1(n12832), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8052) );
  NAND2_X1 U10617 ( .A1(n8123), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8051) );
  NAND2_X1 U10618 ( .A1(n8068), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8050) );
  NAND2_X1 U10619 ( .A1(n8386), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8049) );
  NAND3_X1 U10620 ( .A1(n8079), .A2(SI_2_), .A3(n8053), .ZN(n8061) );
  INV_X1 U10621 ( .A(SI_1_), .ZN(n15702) );
  OAI21_X1 U10622 ( .B1(SI_2_), .B2(n15702), .A(n8058), .ZN(n8056) );
  OAI21_X1 U10623 ( .B1(SI_1_), .B2(n10324), .A(n8054), .ZN(n8055) );
  NAND2_X1 U10624 ( .A1(n8056), .A2(n8055), .ZN(n8060) );
  OAI211_X1 U10625 ( .C1(SI_1_), .C2(n8058), .A(n8057), .B(n10324), .ZN(n8059)
         );
  NAND3_X1 U10626 ( .A1(n8061), .A2(n8060), .A3(n8059), .ZN(n8082) );
  XNOR2_X1 U10627 ( .A(n8082), .B(n8062), .ZN(n10348) );
  OR2_X1 U10628 ( .A1(n8063), .A2(n8266), .ZN(n8064) );
  NAND2_X1 U10629 ( .A1(n8353), .A2(n12536), .ZN(n8065) );
  INV_X1 U10630 ( .A(n13980), .ZN(n11257) );
  NAND2_X1 U10631 ( .A1(n11257), .A2(n13741), .ZN(n8067) );
  NAND2_X1 U10632 ( .A1(n12832), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10633 ( .A1(n8123), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8072) );
  INV_X1 U10634 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U10635 ( .A1(n8721), .A2(n8069), .ZN(n8071) );
  NAND2_X1 U10636 ( .A1(n8386), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8070) );
  NAND2_X1 U10637 ( .A1(n8063), .A2(n8075), .ZN(n8077) );
  NAND2_X1 U10638 ( .A1(n8077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8076) );
  MUX2_X1 U10639 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8076), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8078) );
  AND2_X1 U10640 ( .A1(n8078), .A2(n8117), .ZN(n10501) );
  AOI22_X1 U10641 ( .A1(n8354), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8353), .B2(
        n10501), .ZN(n8089) );
  NAND2_X1 U10642 ( .A1(n8080), .A2(n8079), .ZN(n8097) );
  NAND2_X1 U10643 ( .A1(n8097), .A2(SI_2_), .ZN(n8084) );
  NAND2_X1 U10644 ( .A1(n8082), .A2(n8081), .ZN(n8083) );
  NAND2_X1 U10645 ( .A1(n8084), .A2(n8083), .ZN(n8087) );
  XNOR2_X1 U10646 ( .A(n8085), .B(SI_3_), .ZN(n8086) );
  NAND2_X1 U10647 ( .A1(n10363), .A2(n8102), .ZN(n8088) );
  XNOR2_X1 U10648 ( .A(n13979), .B(n13767), .ZN(n13910) );
  NAND2_X1 U10649 ( .A1(n11255), .A2(n13910), .ZN(n11594) );
  INV_X1 U10650 ( .A(n13979), .ZN(n11598) );
  NAND2_X1 U10651 ( .A1(n11598), .A2(n13767), .ZN(n11592) );
  NAND2_X1 U10652 ( .A1(n11594), .A2(n11592), .ZN(n8105) );
  NAND2_X1 U10653 ( .A1(n12832), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U10654 ( .A1(n8123), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8092) );
  OAI21_X1 U10655 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8108), .ZN(n11607) );
  INV_X1 U10656 ( .A(n11607), .ZN(n10694) );
  NAND2_X1 U10657 ( .A1(n8386), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8090) );
  NAND2_X1 U10658 ( .A1(n8117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8094) );
  XNOR2_X1 U10659 ( .A(n8094), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10503) );
  INV_X1 U10660 ( .A(n8095), .ZN(n8096) );
  NAND2_X1 U10661 ( .A1(n8097), .A2(n8096), .ZN(n8099) );
  NAND2_X1 U10662 ( .A1(n8099), .A2(n8098), .ZN(n8101) );
  XNOR2_X1 U10663 ( .A(n8101), .B(n8100), .ZN(n10350) );
  NAND2_X1 U10664 ( .A1(n10350), .A2(n8102), .ZN(n8103) );
  XNOR2_X1 U10665 ( .A(n13978), .B(n15632), .ZN(n13908) );
  INV_X1 U10666 ( .A(n13978), .ZN(n11256) );
  NAND2_X1 U10667 ( .A1(n11256), .A2(n15632), .ZN(n8106) );
  NAND2_X1 U10668 ( .A1(n12832), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10669 ( .A1(n8123), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8112) );
  INV_X1 U10670 ( .A(n8107), .ZN(n8125) );
  NAND2_X1 U10671 ( .A1(n8108), .A2(n10519), .ZN(n8109) );
  AND2_X1 U10672 ( .A1(n8125), .A2(n8109), .ZN(n11582) );
  NAND2_X1 U10673 ( .A1(n8386), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8110) );
  XNOR2_X1 U10674 ( .A(n8114), .B(SI_5_), .ZN(n8115) );
  NAND2_X1 U10675 ( .A1(n10392), .A2(n8102), .ZN(n8122) );
  INV_X1 U10676 ( .A(n8117), .ZN(n8119) );
  NAND2_X1 U10677 ( .A1(n8119), .A2(n8118), .ZN(n8142) );
  NAND2_X1 U10678 ( .A1(n8142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8120) );
  XNOR2_X1 U10679 ( .A(n8120), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U10680 ( .A1(n8354), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8353), .B2(
        n10525), .ZN(n8121) );
  AND2_X1 U10681 ( .A1(n11597), .A2(n13726), .ZN(n11520) );
  NAND2_X1 U10682 ( .A1(n12832), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8130) );
  NAND2_X1 U10683 ( .A1(n8123), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8129) );
  INV_X1 U10684 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8124) );
  NAND2_X1 U10685 ( .A1(n8125), .A2(n8124), .ZN(n8126) );
  AND2_X1 U10686 ( .A1(n8161), .A2(n8126), .ZN(n10886) );
  NAND2_X1 U10687 ( .A1(n8721), .A2(n10886), .ZN(n8128) );
  NAND2_X1 U10688 ( .A1(n8386), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8127) );
  INV_X1 U10689 ( .A(n8133), .ZN(n8135) );
  NAND2_X1 U10690 ( .A1(n8135), .A2(n8132), .ZN(n8141) );
  NAND3_X1 U10691 ( .A1(n8148), .A2(n7925), .A3(n8133), .ZN(n8140) );
  OAI211_X1 U10692 ( .C1(n8137), .C2(n8136), .A(n8135), .B(n8134), .ZN(n8138)
         );
  NAND2_X1 U10693 ( .A1(n8138), .A2(n8149), .ZN(n8139) );
  NAND2_X1 U10694 ( .A1(n8224), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8143) );
  XNOR2_X1 U10695 ( .A(n8143), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U10696 ( .A1(n8354), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8353), .B2(
        n10724), .ZN(n8144) );
  XNOR2_X1 U10697 ( .A(n13976), .B(n13777), .ZN(n13732) );
  NAND2_X1 U10698 ( .A1(n13727), .A2(n13977), .ZN(n8146) );
  AND2_X1 U10699 ( .A1(n13732), .A2(n8146), .ZN(n8147) );
  NAND2_X1 U10700 ( .A1(n13776), .A2(n13777), .ZN(n11538) );
  NAND2_X1 U10701 ( .A1(n8148), .A2(n7925), .ZN(n8151) );
  INV_X1 U10702 ( .A(n8149), .ZN(n8150) );
  NAND2_X1 U10703 ( .A1(n8151), .A2(n8150), .ZN(n8153) );
  NAND2_X1 U10704 ( .A1(n8153), .A2(n8152), .ZN(n8155) );
  NAND2_X1 U10705 ( .A1(n10390), .A2(n8102), .ZN(n8159) );
  NAND2_X1 U10706 ( .A1(n8156), .A2(n6756), .ZN(n8169) );
  NAND2_X1 U10707 ( .A1(n8169), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8157) );
  XNOR2_X1 U10708 ( .A(n8157), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U10709 ( .A1(n8354), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8353), .B2(
        n10740), .ZN(n8158) );
  NAND2_X1 U10710 ( .A1(n12832), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10711 ( .A1(n12833), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10712 ( .A1(n8161), .A2(n8160), .ZN(n8162) );
  AND2_X1 U10713 ( .A1(n8195), .A2(n8162), .ZN(n10988) );
  NAND2_X1 U10714 ( .A1(n8721), .A2(n10988), .ZN(n8164) );
  NAND2_X1 U10715 ( .A1(n8386), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8163) );
  XNOR2_X1 U10716 ( .A(n15650), .B(n11197), .ZN(n13738) );
  INV_X1 U10717 ( .A(n13738), .ZN(n13909) );
  NAND2_X1 U10718 ( .A1(n15650), .A2(n11197), .ZN(n11553) );
  XNOR2_X1 U10719 ( .A(n8168), .B(SI_8_), .ZN(n8179) );
  NAND2_X1 U10720 ( .A1(n10441), .A2(n8102), .ZN(n8174) );
  NAND2_X1 U10721 ( .A1(n8171), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8170) );
  MUX2_X1 U10722 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8170), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8172) );
  NAND2_X1 U10723 ( .A1(n8172), .A2(n8187), .ZN(n10934) );
  INV_X1 U10724 ( .A(n10934), .ZN(n10938) );
  AOI22_X1 U10725 ( .A1(n8354), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10938), 
        .B2(n8353), .ZN(n8173) );
  NAND2_X1 U10726 ( .A1(n12832), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8178) );
  XNOR2_X1 U10727 ( .A(n8195), .B(P2_REG3_REG_8__SCAN_IN), .ZN(n11196) );
  NAND2_X1 U10728 ( .A1(n8721), .A2(n11196), .ZN(n8176) );
  NAND2_X1 U10729 ( .A1(n9609), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8175) );
  XNOR2_X1 U10730 ( .A(n13789), .B(n13974), .ZN(n13914) );
  INV_X1 U10731 ( .A(n13974), .ZN(n10987) );
  NAND2_X1 U10732 ( .A1(n13789), .A2(n10987), .ZN(n11864) );
  INV_X1 U10733 ( .A(n8179), .ZN(n8180) );
  NAND2_X1 U10734 ( .A1(n8181), .A2(n8180), .ZN(n8183) );
  NAND2_X1 U10735 ( .A1(n8183), .A2(n8182), .ZN(n8185) );
  XNOR2_X1 U10736 ( .A(n8185), .B(n8184), .ZN(n10454) );
  NAND2_X1 U10737 ( .A1(n10454), .A2(n8102), .ZN(n8192) );
  NAND2_X1 U10738 ( .A1(n8187), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8186) );
  MUX2_X1 U10739 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8186), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8189) );
  INV_X1 U10740 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U10741 ( .A1(n8189), .A2(n8209), .ZN(n15539) );
  INV_X1 U10742 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10455) );
  OAI22_X1 U10743 ( .A1(n15539), .A2(n8048), .B1(n9606), .B2(n10455), .ZN(
        n8190) );
  INV_X1 U10744 ( .A(n8190), .ZN(n8191) );
  NAND2_X1 U10745 ( .A1(n12833), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10746 ( .A1(n9609), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8199) );
  INV_X1 U10747 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8194) );
  INV_X1 U10748 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8193) );
  OAI21_X1 U10749 ( .B1(n8195), .B2(n8194), .A(n8193), .ZN(n8196) );
  AND2_X1 U10750 ( .A1(n8214), .A2(n8196), .ZN(n11874) );
  NAND2_X1 U10751 ( .A1(n8721), .A2(n11874), .ZN(n8198) );
  NAND2_X1 U10752 ( .A1(n12832), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8197) );
  NAND4_X1 U10753 ( .A1(n8200), .A2(n8199), .A3(n8198), .A4(n8197), .ZN(n13973) );
  XNOR2_X1 U10754 ( .A(n13794), .B(n13973), .ZN(n13902) );
  NAND2_X1 U10755 ( .A1(n13794), .A2(n11435), .ZN(n11955) );
  NAND2_X1 U10756 ( .A1(n8201), .A2(n7932), .ZN(n8203) );
  NAND2_X1 U10757 ( .A1(n8203), .A2(n8202), .ZN(n8205) );
  NAND2_X1 U10758 ( .A1(n8205), .A2(n8204), .ZN(n8208) );
  XNOR2_X1 U10759 ( .A(n8206), .B(SI_10_), .ZN(n8207) );
  XNOR2_X1 U10760 ( .A(n8208), .B(n8207), .ZN(n10447) );
  NAND2_X1 U10761 ( .A1(n10447), .A2(n8102), .ZN(n8212) );
  NAND2_X1 U10762 ( .A1(n8209), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8210) );
  AOI22_X1 U10763 ( .A1(n15553), .A2(n8353), .B1(n8354), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U10764 ( .A1(n12832), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8219) );
  NAND2_X1 U10765 ( .A1(n12833), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8218) );
  INV_X1 U10766 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U10767 ( .A1(n8214), .A2(n8213), .ZN(n8215) );
  AND2_X1 U10768 ( .A1(n8240), .A2(n8215), .ZN(n11433) );
  NAND2_X1 U10769 ( .A1(n8721), .A2(n11433), .ZN(n8217) );
  NAND2_X1 U10770 ( .A1(n9609), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8216) );
  NAND4_X1 U10771 ( .A1(n8219), .A2(n8218), .A3(n8217), .A4(n8216), .ZN(n14303) );
  XNOR2_X1 U10772 ( .A(n14405), .B(n14303), .ZN(n13901) );
  INV_X1 U10773 ( .A(n14303), .ZN(n11778) );
  NAND2_X1 U10774 ( .A1(n14405), .A2(n11778), .ZN(n14298) );
  XNOR2_X1 U10775 ( .A(n8221), .B(n8220), .ZN(n10444) );
  NAND2_X1 U10776 ( .A1(n10444), .A2(n8102), .ZN(n8228) );
  INV_X1 U10777 ( .A(n8222), .ZN(n8223) );
  OAI21_X1 U10778 ( .B1(n8224), .B2(n8223), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8225) );
  MUX2_X1 U10779 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8225), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n8226) );
  NAND2_X1 U10780 ( .A1(n8226), .A2(n8251), .ZN(n11105) );
  INV_X1 U10781 ( .A(n11105), .ZN(n10943) );
  AOI22_X1 U10782 ( .A1(n8354), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8353), 
        .B2(n10943), .ZN(n8227) );
  NAND2_X1 U10783 ( .A1(n12832), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8232) );
  NAND2_X1 U10784 ( .A1(n12833), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8231) );
  XNOR2_X1 U10785 ( .A(n8240), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n11777) );
  NAND2_X1 U10786 ( .A1(n8721), .A2(n11777), .ZN(n8230) );
  NAND2_X1 U10787 ( .A1(n8386), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8229) );
  NAND4_X1 U10788 ( .A1(n8232), .A2(n8231), .A3(n8230), .A4(n8229), .ZN(n13972) );
  XNOR2_X1 U10789 ( .A(n14399), .B(n13972), .ZN(n13913) );
  INV_X1 U10790 ( .A(n13972), .ZN(n11434) );
  XNOR2_X1 U10791 ( .A(n8234), .B(n8233), .ZN(n10458) );
  NAND2_X1 U10792 ( .A1(n10458), .A2(n8102), .ZN(n8237) );
  NAND2_X1 U10793 ( .A1(n8251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8235) );
  XNOR2_X1 U10794 ( .A(n8235), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U10795 ( .A1(n8354), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8353), 
        .B2(n11618), .ZN(n8236) );
  NAND2_X1 U10796 ( .A1(n12832), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U10797 ( .A1(n12833), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8244) );
  OAI21_X1 U10798 ( .B1(n8240), .B2(n8239), .A(n8238), .ZN(n8241) );
  AND2_X1 U10799 ( .A1(n8241), .A2(n8257), .ZN(n12135) );
  NAND2_X1 U10800 ( .A1(n8721), .A2(n12135), .ZN(n8243) );
  NAND2_X1 U10801 ( .A1(n9609), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8242) );
  NAND4_X1 U10802 ( .A1(n8245), .A2(n8244), .A3(n8243), .A4(n8242), .ZN(n14305) );
  INV_X1 U10803 ( .A(n14305), .ZN(n8247) );
  OR2_X1 U10804 ( .A1(n14393), .A2(n8247), .ZN(n8246) );
  NAND2_X1 U10805 ( .A1(n14393), .A2(n8247), .ZN(n8248) );
  XNOR2_X1 U10806 ( .A(n8250), .B(n8249), .ZN(n10464) );
  NAND2_X1 U10807 ( .A1(n10464), .A2(n8102), .ZN(n8255) );
  NAND2_X1 U10808 ( .A1(n8252), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8253) );
  XNOR2_X1 U10809 ( .A(n8253), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15566) );
  AOI22_X1 U10810 ( .A1(n8354), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8353), 
        .B2(n15566), .ZN(n8254) );
  NAND2_X1 U10811 ( .A1(n12832), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U10812 ( .A1(n12833), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8261) );
  INV_X1 U10813 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U10814 ( .A1(n8257), .A2(n8256), .ZN(n8258) );
  AND2_X1 U10815 ( .A1(n8290), .A2(n8258), .ZN(n12190) );
  NAND2_X1 U10816 ( .A1(n8721), .A2(n12190), .ZN(n8260) );
  NAND2_X1 U10817 ( .A1(n9609), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8259) );
  NAND4_X1 U10818 ( .A1(n8262), .A2(n8261), .A3(n8260), .A4(n8259), .ZN(n14269) );
  AND2_X1 U10819 ( .A1(n14389), .A2(n13574), .ZN(n8263) );
  OR2_X1 U10820 ( .A1(n14389), .A2(n13574), .ZN(n8264) );
  XNOR2_X1 U10821 ( .A(n8279), .B(n8278), .ZN(n10655) );
  NAND2_X1 U10822 ( .A1(n10655), .A2(n8102), .ZN(n8269) );
  INV_X1 U10823 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U10824 ( .A1(n8282), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8267) );
  XNOR2_X1 U10825 ( .A(n8267), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U10826 ( .A1(n8354), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8353), 
        .B2(n12157), .ZN(n8268) );
  NAND2_X1 U10827 ( .A1(n12832), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8273) );
  NAND2_X1 U10828 ( .A1(n12833), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8272) );
  XNOR2_X1 U10829 ( .A(n8290), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n14273) );
  NAND2_X1 U10830 ( .A1(n8721), .A2(n14273), .ZN(n8271) );
  NAND2_X1 U10831 ( .A1(n8386), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8270) );
  NAND4_X1 U10832 ( .A1(n8273), .A2(n8272), .A3(n8271), .A4(n8270), .ZN(n14254) );
  INV_X1 U10833 ( .A(n14254), .ZN(n8274) );
  NOR2_X1 U10834 ( .A1(n14383), .A2(n8274), .ZN(n8275) );
  INV_X1 U10835 ( .A(n8276), .ZN(n8277) );
  XNOR2_X1 U10836 ( .A(n8280), .B(SI_15_), .ZN(n8281) );
  NAND2_X1 U10837 ( .A1(n10704), .A2(n8102), .ZN(n8287) );
  INV_X1 U10838 ( .A(n8282), .ZN(n8284) );
  INV_X1 U10839 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10840 ( .A1(n8284), .A2(n8283), .ZN(n8301) );
  NAND2_X1 U10841 ( .A1(n8301), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8285) );
  XNOR2_X1 U10842 ( .A(n8285), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13998) );
  AOI22_X1 U10843 ( .A1(n8354), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8353), 
        .B2(n13998), .ZN(n8286) );
  NAND2_X1 U10844 ( .A1(n12832), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U10845 ( .A1(n12833), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8294) );
  INV_X1 U10846 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8289) );
  INV_X1 U10847 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8288) );
  OAI21_X1 U10848 ( .B1(n8290), .B2(n8289), .A(n8288), .ZN(n8291) );
  AND2_X1 U10849 ( .A1(n8291), .A2(n8309), .ZN(n14260) );
  NAND2_X1 U10850 ( .A1(n8721), .A2(n14260), .ZN(n8293) );
  NAND2_X1 U10851 ( .A1(n9609), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8292) );
  NAND4_X1 U10852 ( .A1(n8295), .A2(n8294), .A3(n8293), .A4(n8292), .ZN(n14268) );
  INV_X1 U10853 ( .A(n14268), .ZN(n8297) );
  OR2_X1 U10854 ( .A1(n14259), .A2(n8297), .ZN(n8296) );
  NAND2_X1 U10855 ( .A1(n14259), .A2(n8297), .ZN(n8298) );
  XNOR2_X1 U10856 ( .A(n8300), .B(n8299), .ZN(n10557) );
  NAND2_X1 U10857 ( .A1(n10557), .A2(n8102), .ZN(n8308) );
  NAND2_X1 U10858 ( .A1(n8303), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8302) );
  MUX2_X1 U10859 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8302), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8306) );
  INV_X1 U10860 ( .A(n8303), .ZN(n8305) );
  INV_X1 U10861 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8304) );
  NAND2_X1 U10862 ( .A1(n8305), .A2(n8304), .ZN(n8332) );
  NAND2_X1 U10863 ( .A1(n8306), .A2(n8332), .ZN(n15585) );
  INV_X1 U10864 ( .A(n15585), .ZN(n13988) );
  AOI22_X1 U10865 ( .A1(n8354), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n13988), 
        .B2(n8353), .ZN(n8307) );
  NAND2_X1 U10866 ( .A1(n12833), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U10867 ( .A1(n9609), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8313) );
  INV_X1 U10868 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n15826) );
  NAND2_X1 U10869 ( .A1(n8309), .A2(n15826), .ZN(n8310) );
  AND2_X1 U10870 ( .A1(n8324), .A2(n8310), .ZN(n14235) );
  NAND2_X1 U10871 ( .A1(n8721), .A2(n14235), .ZN(n8312) );
  NAND2_X1 U10872 ( .A1(n12832), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8311) );
  NAND4_X1 U10873 ( .A1(n8314), .A2(n8313), .A3(n8312), .A4(n8311), .ZN(n14253) );
  INV_X1 U10874 ( .A(n14253), .ZN(n13719) );
  OR2_X1 U10875 ( .A1(n14372), .A2(n13719), .ZN(n8315) );
  NAND2_X1 U10876 ( .A1(n14372), .A2(n13719), .ZN(n8316) );
  XNOR2_X1 U10877 ( .A(n8317), .B(SI_17_), .ZN(n8318) );
  XNOR2_X1 U10878 ( .A(n8319), .B(n8318), .ZN(n10686) );
  NAND2_X1 U10879 ( .A1(n10686), .A2(n8102), .ZN(n8322) );
  NAND2_X1 U10880 ( .A1(n8332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8320) );
  XNOR2_X1 U10881 ( .A(n8320), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15598) );
  AOI22_X1 U10882 ( .A1(n8353), .A2(n15598), .B1(n8354), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10883 ( .A1(n8324), .A2(n8323), .ZN(n8325) );
  AND2_X1 U10884 ( .A1(n8337), .A2(n8325), .ZN(n14220) );
  NAND2_X1 U10885 ( .A1(n14220), .A2(n8721), .ZN(n8329) );
  NAND2_X1 U10886 ( .A1(n12833), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U10887 ( .A1(n12832), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U10888 ( .A1(n8386), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8326) );
  NAND4_X1 U10889 ( .A1(n8329), .A2(n8328), .A3(n8327), .A4(n8326), .ZN(n14231) );
  INV_X1 U10890 ( .A(n14231), .ZN(n13633) );
  AND2_X1 U10891 ( .A1(n14368), .A2(n13633), .ZN(n8330) );
  OR2_X1 U10892 ( .A1(n14368), .A2(n13633), .ZN(n8331) );
  NAND2_X1 U10893 ( .A1(n10993), .A2(n8102), .ZN(n8335) );
  OAI21_X1 U10894 ( .B1(n8332), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8333) );
  XNOR2_X1 U10895 ( .A(n8333), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14001) );
  AOI22_X1 U10896 ( .A1(n14001), .A2(n8353), .B1(n8354), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8334) );
  INV_X1 U10897 ( .A(n8386), .ZN(n12836) );
  INV_X1 U10898 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14442) );
  INV_X1 U10899 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U10900 ( .A1(n8337), .A2(n8336), .ZN(n8338) );
  NAND2_X1 U10901 ( .A1(n8357), .A2(n8338), .ZN(n14206) );
  OR2_X1 U10902 ( .A1(n14206), .A2(n8461), .ZN(n8342) );
  NAND2_X1 U10903 ( .A1(n12833), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U10904 ( .A1(n12832), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8339) );
  AND2_X1 U10905 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  OAI211_X1 U10906 ( .C1(n12836), .C2(n14442), .A(n8342), .B(n8341), .ZN(
        n13971) );
  INV_X1 U10907 ( .A(n13971), .ZN(n8529) );
  NAND2_X1 U10908 ( .A1(n8345), .A2(SI_18_), .ZN(n8346) );
  NAND2_X1 U10909 ( .A1(n8348), .A2(n8347), .ZN(n8349) );
  NAND2_X1 U10910 ( .A1(n8831), .A2(n8102), .ZN(n8356) );
  XNOR2_X2 U10911 ( .A(n8352), .B(P2_IR_REG_19__SCAN_IN), .ZN(n14017) );
  AOI22_X1 U10912 ( .A1(n8354), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n14017), 
        .B2(n8353), .ZN(n8355) );
  NAND2_X1 U10913 ( .A1(n8357), .A2(n13595), .ZN(n8358) );
  NAND2_X1 U10914 ( .A1(n8367), .A2(n8358), .ZN(n14191) );
  AOI22_X1 U10915 ( .A1(n12832), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n12833), 
        .B2(P2_REG1_REG_19__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10916 ( .A1(n9609), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8359) );
  OAI211_X1 U10917 ( .C1(n14191), .C2(n8461), .A(n8360), .B(n8359), .ZN(n13970) );
  NOR2_X1 U10918 ( .A1(n14196), .A2(n14153), .ZN(n14152) );
  NAND2_X1 U10919 ( .A1(n14365), .A2(n8529), .ZN(n14150) );
  NAND2_X1 U10920 ( .A1(n14150), .A2(n13970), .ZN(n8362) );
  INV_X1 U10921 ( .A(n14150), .ZN(n8361) );
  AOI22_X1 U10922 ( .A1(n14196), .A2(n8362), .B1(n8361), .B2(n14153), .ZN(
        n8372) );
  NAND2_X1 U10923 ( .A1(n11202), .A2(n8102), .ZN(n8365) );
  OR2_X1 U10924 ( .A1(n9606), .A2(n11316), .ZN(n8364) );
  INV_X1 U10925 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8371) );
  INV_X1 U10926 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U10927 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  NAND2_X1 U10928 ( .A1(n8384), .A2(n8368), .ZN(n14176) );
  OR2_X1 U10929 ( .A1(n14176), .A2(n8461), .ZN(n8370) );
  AOI22_X1 U10930 ( .A1(n12832), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n12833), 
        .B2(P2_REG1_REG_20__SCAN_IN), .ZN(n8369) );
  OAI211_X1 U10931 ( .C1(n12836), .C2(n8371), .A(n8370), .B(n8369), .ZN(n13969) );
  INV_X1 U10932 ( .A(n13969), .ZN(n13620) );
  NAND2_X1 U10933 ( .A1(n14353), .A2(n13620), .ZN(n14154) );
  OR2_X1 U10934 ( .A1(n14353), .A2(n13620), .ZN(n13899) );
  NAND2_X1 U10935 ( .A1(n8374), .A2(n8373), .ZN(n8377) );
  OR2_X1 U10936 ( .A1(n8375), .A2(n11183), .ZN(n8376) );
  NAND2_X1 U10937 ( .A1(n8377), .A2(n8376), .ZN(n8380) );
  XNOR2_X1 U10938 ( .A(n8378), .B(SI_21_), .ZN(n8379) );
  NAND2_X1 U10939 ( .A1(n11287), .A2(n8102), .ZN(n8382) );
  INV_X1 U10940 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11288) );
  OR2_X1 U10941 ( .A1(n9606), .A2(n11288), .ZN(n8381) );
  NAND2_X1 U10942 ( .A1(n8384), .A2(n8383), .ZN(n8385) );
  NAND2_X1 U10943 ( .A1(n8398), .A2(n8385), .ZN(n14158) );
  OR2_X1 U10944 ( .A1(n14158), .A2(n8461), .ZN(n8391) );
  INV_X1 U10945 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n14159) );
  NAND2_X1 U10946 ( .A1(n8386), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10947 ( .A1(n12833), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8387) );
  OAI211_X1 U10948 ( .C1(n9613), .C2(n14159), .A(n8388), .B(n8387), .ZN(n8389)
         );
  INV_X1 U10949 ( .A(n8389), .ZN(n8390) );
  NAND2_X1 U10950 ( .A1(n8391), .A2(n8390), .ZN(n13968) );
  INV_X1 U10951 ( .A(n13968), .ZN(n13664) );
  OR2_X1 U10952 ( .A1(n14345), .A2(n13664), .ZN(n8392) );
  XNOR2_X1 U10953 ( .A(n8810), .B(n8394), .ZN(n11363) );
  NAND2_X1 U10954 ( .A1(n11363), .A2(n8102), .ZN(n8396) );
  INV_X1 U10955 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11365) );
  OR2_X1 U10956 ( .A1(n9606), .A2(n11365), .ZN(n8395) );
  NAND2_X1 U10957 ( .A1(n8398), .A2(n8397), .ZN(n8399) );
  AND2_X1 U10958 ( .A1(n8426), .A2(n8399), .ZN(n13663) );
  NAND2_X1 U10959 ( .A1(n13663), .A2(n8721), .ZN(n8404) );
  INV_X1 U10960 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n14142) );
  NAND2_X1 U10961 ( .A1(n9609), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10962 ( .A1(n12833), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8400) );
  OAI211_X1 U10963 ( .C1(n9613), .C2(n14142), .A(n8401), .B(n8400), .ZN(n8402)
         );
  INV_X1 U10964 ( .A(n8402), .ZN(n8403) );
  XNOR2_X1 U10965 ( .A(n14145), .B(n13967), .ZN(n13924) );
  INV_X1 U10966 ( .A(n13967), .ZN(n14117) );
  OR2_X1 U10967 ( .A1(n14145), .A2(n14117), .ZN(n8405) );
  NAND2_X1 U10968 ( .A1(n11611), .A2(n8102), .ZN(n8409) );
  INV_X1 U10969 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11613) );
  OR2_X1 U10970 ( .A1(n9606), .A2(n11613), .ZN(n8408) );
  INV_X1 U10971 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13646) );
  NAND2_X1 U10972 ( .A1(n8428), .A2(n13646), .ZN(n8410) );
  NAND2_X1 U10973 ( .A1(n8439), .A2(n8410), .ZN(n14107) );
  INV_X1 U10974 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14106) );
  NAND2_X1 U10975 ( .A1(n9609), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8412) );
  NAND2_X1 U10976 ( .A1(n12833), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8411) );
  OAI211_X1 U10977 ( .C1(n9613), .C2(n14106), .A(n8412), .B(n8411), .ZN(n8413)
         );
  INV_X1 U10978 ( .A(n8413), .ZN(n8414) );
  NAND2_X1 U10979 ( .A1(n14109), .A2(n14119), .ZN(n10271) );
  NAND2_X1 U10980 ( .A1(n8810), .A2(n8416), .ZN(n8419) );
  NAND2_X1 U10981 ( .A1(n8417), .A2(SI_22_), .ZN(n8418) );
  NAND2_X1 U10982 ( .A1(n8419), .A2(n8418), .ZN(n8422) );
  XNOR2_X1 U10983 ( .A(n8420), .B(SI_23_), .ZN(n8421) );
  NAND2_X1 U10984 ( .A1(n11494), .A2(n8102), .ZN(n8424) );
  INV_X1 U10985 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11493) );
  OR2_X1 U10986 ( .A1(n9606), .A2(n11493), .ZN(n8423) );
  INV_X1 U10987 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10988 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  NAND2_X1 U10989 ( .A1(n8428), .A2(n8427), .ZN(n14123) );
  INV_X1 U10990 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n15711) );
  NAND2_X1 U10991 ( .A1(n12832), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U10992 ( .A1(n9609), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8429) );
  OAI211_X1 U10993 ( .C1(n8570), .C2(n15711), .A(n8430), .B(n8429), .ZN(n8431)
         );
  INV_X1 U10994 ( .A(n8431), .ZN(n8432) );
  NAND2_X1 U10995 ( .A1(n14129), .A2(n13665), .ZN(n8434) );
  AND2_X1 U10996 ( .A1(n10271), .A2(n8434), .ZN(n12823) );
  XNOR2_X1 U10997 ( .A(n8436), .B(n8435), .ZN(n11769) );
  NAND2_X1 U10998 ( .A1(n11769), .A2(n8102), .ZN(n8438) );
  OR2_X1 U10999 ( .A1(n9606), .A2(n11770), .ZN(n8437) );
  XNOR2_X1 U11000 ( .A(n8439), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14090) );
  NAND2_X1 U11001 ( .A1(n14090), .A2(n8721), .ZN(n8445) );
  INV_X1 U11002 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U11003 ( .A1(n12833), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U11004 ( .A1(n9609), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8440) );
  OAI211_X1 U11005 ( .C1(n8442), .C2(n9613), .A(n8441), .B(n8440), .ZN(n8443)
         );
  INV_X1 U11006 ( .A(n8443), .ZN(n8444) );
  XNOR2_X1 U11007 ( .A(n13859), .B(n13964), .ZN(n13928) );
  OR2_X1 U11008 ( .A1(n14109), .A2(n14119), .ZN(n8539) );
  OR2_X1 U11009 ( .A1(n14129), .A2(n13665), .ZN(n14098) );
  NAND2_X1 U11010 ( .A1(n8539), .A2(n14098), .ZN(n8446) );
  NAND2_X1 U11011 ( .A1(n8446), .A2(n10271), .ZN(n8447) );
  NAND2_X1 U11012 ( .A1(n13928), .A2(n8447), .ZN(n12825) );
  AOI21_X1 U11013 ( .B1(n14114), .B2(n12823), .A(n12825), .ZN(n8449) );
  NAND2_X1 U11014 ( .A1(n13859), .A2(n13698), .ZN(n12824) );
  INV_X1 U11015 ( .A(n12824), .ZN(n8448) );
  NOR2_X1 U11016 ( .A1(n8449), .A2(n8448), .ZN(n8450) );
  XOR2_X1 U11017 ( .A(n13927), .B(n8450), .Z(n8467) );
  NOR2_X2 U11018 ( .A1(n8455), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n8472) );
  XNOR2_X2 U11019 ( .A(n8451), .B(n8471), .ZN(n13944) );
  NAND2_X1 U11020 ( .A1(n13954), .A2(n14017), .ZN(n8458) );
  INV_X1 U11021 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U11022 ( .A1(n8455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8456) );
  INV_X1 U11023 ( .A(n13941), .ZN(n11289) );
  OR2_X1 U11024 ( .A1(n8541), .A2(n11289), .ZN(n8457) );
  INV_X1 U11025 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13563) );
  INV_X1 U11026 ( .A(n8565), .ZN(n8566) );
  NAND2_X1 U11027 ( .A1(n8459), .A2(n13563), .ZN(n8460) );
  INV_X1 U11028 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n15895) );
  NAND2_X1 U11029 ( .A1(n12832), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U11030 ( .A1(n12833), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8462) );
  OAI211_X1 U11031 ( .C1(n15895), .C2(n12836), .A(n8463), .B(n8462), .ZN(n8464) );
  INV_X1 U11032 ( .A(n8464), .ZN(n8465) );
  AND2_X1 U11033 ( .A1(n13954), .A2(n13941), .ZN(n10483) );
  NAND2_X1 U11034 ( .A1(n10483), .A2(n10490), .ZN(n14118) );
  INV_X1 U11035 ( .A(n10490), .ZN(n8466) );
  AOI22_X1 U11036 ( .A1(n14046), .A2(n14304), .B1(n14302), .B2(n13964), .ZN(
        n13704) );
  NOR2_X1 U11037 ( .A1(n13745), .A2(n13756), .ZN(n12011) );
  INV_X1 U11038 ( .A(n13741), .ZN(n15626) );
  NAND2_X1 U11039 ( .A1(n12011), .A2(n15626), .ZN(n11261) );
  NOR2_X4 U11040 ( .A1(n11604), .A2(n13726), .ZN(n11527) );
  INV_X1 U11041 ( .A(n14405), .ZN(n11964) );
  NAND2_X1 U11042 ( .A1(n11872), .A2(n11964), .ZN(n14287) );
  OR2_X2 U11043 ( .A1(n14287), .A2(n14399), .ZN(n14288) );
  INV_X1 U11044 ( .A(n14383), .ZN(n14276) );
  INV_X1 U11045 ( .A(n14365), .ZN(n14209) );
  AOI211_X1 U11046 ( .C1(n13862), .C2(n10268), .A(n14074), .B(n8582), .ZN(
        n14084) );
  NAND2_X1 U11047 ( .A1(n8541), .A2(n11528), .ZN(n13952) );
  NAND2_X1 U11048 ( .A1(n13952), .A2(n11235), .ZN(n15640) );
  INV_X1 U11049 ( .A(n8475), .ZN(n8476) );
  NAND2_X1 U11050 ( .A1(n8476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8477) );
  MUX2_X1 U11051 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8477), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8478) );
  NAND2_X1 U11052 ( .A1(n8478), .A2(n8479), .ZN(n11615) );
  INV_X1 U11053 ( .A(n11615), .ZN(n8500) );
  NAND2_X1 U11054 ( .A1(n8479), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8480) );
  XNOR2_X1 U11055 ( .A(n8480), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8487) );
  NAND3_X1 U11056 ( .A1(n14476), .A2(n8500), .A3(n8487), .ZN(n10281) );
  INV_X1 U11057 ( .A(n8481), .ZN(n8482) );
  NAND2_X1 U11058 ( .A1(n8482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8484) );
  INV_X1 U11059 ( .A(n8487), .ZN(n11771) );
  XNOR2_X1 U11060 ( .A(n11615), .B(P2_B_REG_SCAN_IN), .ZN(n8485) );
  NAND2_X1 U11061 ( .A1(n11771), .A2(n8485), .ZN(n8486) );
  INV_X1 U11062 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15618) );
  NAND2_X1 U11063 ( .A1(n15610), .A2(n15618), .ZN(n8489) );
  OR2_X1 U11064 ( .A1(n14476), .A2(n8487), .ZN(n8488) );
  NAND2_X1 U11065 ( .A1(n8489), .A2(n8488), .ZN(n11227) );
  AND2_X1 U11066 ( .A1(n15615), .A2(n11227), .ZN(n15616) );
  NOR4_X1 U11067 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8497) );
  INV_X1 U11068 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15923) );
  INV_X1 U11069 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15894) );
  INV_X1 U11070 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15842) );
  INV_X1 U11071 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15853) );
  NAND4_X1 U11072 ( .A1(n15923), .A2(n15894), .A3(n15842), .A4(n15853), .ZN(
        n15709) );
  NOR4_X1 U11073 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8493) );
  NOR4_X1 U11074 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n8492) );
  NOR4_X1 U11075 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n8491) );
  NOR4_X1 U11076 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n8490) );
  NAND4_X1 U11077 ( .A1(n8493), .A2(n8492), .A3(n8491), .A4(n8490), .ZN(n8494)
         );
  NOR4_X1 U11078 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n15709), .A4(n8494), .ZN(n8496) );
  NOR4_X1 U11079 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8495) );
  NAND3_X1 U11080 ( .A1(n8497), .A2(n8496), .A3(n8495), .ZN(n8498) );
  NAND2_X1 U11081 ( .A1(n13952), .A2(n10483), .ZN(n8729) );
  INV_X1 U11082 ( .A(n8729), .ZN(n8499) );
  AND2_X2 U11083 ( .A1(n8541), .A2(n14017), .ZN(n13940) );
  NAND2_X1 U11084 ( .A1(n13940), .A2(n11235), .ZN(n8727) );
  INV_X1 U11085 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15613) );
  NAND2_X1 U11086 ( .A1(n15610), .A2(n15613), .ZN(n8502) );
  OR2_X1 U11087 ( .A1(n8500), .A2(n14476), .ZN(n8501) );
  MUX2_X1 U11088 ( .A(n8503), .B(n8547), .S(n15670), .Z(n8545) );
  NOR2_X1 U11089 ( .A1(n13981), .A2(n13745), .ZN(n11074) );
  NOR2_X1 U11090 ( .A1(n13980), .A2(n13741), .ZN(n11077) );
  AOI21_X1 U11091 ( .B1(n12004), .B2(n11074), .A(n11077), .ZN(n8509) );
  NOR2_X1 U11092 ( .A1(n13979), .A2(n13767), .ZN(n11589) );
  NAND2_X1 U11093 ( .A1(n13978), .A2(n15632), .ZN(n8511) );
  NAND2_X1 U11094 ( .A1(n11589), .A2(n8511), .ZN(n8504) );
  INV_X1 U11095 ( .A(n15632), .ZN(n13733) );
  INV_X1 U11096 ( .A(n11233), .ZN(n13606) );
  OR2_X1 U11097 ( .A1(n13904), .A2(n13606), .ZN(n11076) );
  INV_X1 U11098 ( .A(n11076), .ZN(n8505) );
  NAND2_X1 U11099 ( .A1(n8505), .A2(n12004), .ZN(n8508) );
  NAND2_X1 U11100 ( .A1(n11597), .A2(n13727), .ZN(n8507) );
  NAND2_X1 U11101 ( .A1(n13979), .A2(n13767), .ZN(n8510) );
  NAND2_X1 U11102 ( .A1(n13977), .A2(n13726), .ZN(n8512) );
  NAND2_X1 U11103 ( .A1(n13776), .A2(n8512), .ZN(n8513) );
  NAND2_X1 U11104 ( .A1(n8513), .A2(n13777), .ZN(n8515) );
  NAND3_X1 U11105 ( .A1(n13977), .A2(n13976), .A3(n13726), .ZN(n8514) );
  NAND2_X1 U11106 ( .A1(n11536), .A2(n13738), .ZN(n11535) );
  NAND2_X1 U11107 ( .A1(n13975), .A2(n15650), .ZN(n8516) );
  OAI22_X1 U11108 ( .A1(n13794), .A2(n13973), .B1(n13789), .B2(n13974), .ZN(
        n8517) );
  INV_X1 U11109 ( .A(n8517), .ZN(n8518) );
  NAND2_X1 U11110 ( .A1(n13789), .A2(n13974), .ZN(n11861) );
  NAND2_X1 U11111 ( .A1(n11861), .A2(n11435), .ZN(n8520) );
  AND2_X1 U11112 ( .A1(n13974), .A2(n13973), .ZN(n8519) );
  AOI22_X1 U11113 ( .A1(n8520), .A2(n13794), .B1(n8519), .B2(n13789), .ZN(
        n8521) );
  NAND2_X1 U11114 ( .A1(n14405), .A2(n14303), .ZN(n8522) );
  NAND2_X1 U11115 ( .A1(n11952), .A2(n8522), .ZN(n14284) );
  INV_X1 U11116 ( .A(n13913), .ZN(n14299) );
  NAND2_X1 U11117 ( .A1(n14284), .A2(n14299), .ZN(n14286) );
  NAND2_X1 U11118 ( .A1(n14399), .A2(n13972), .ZN(n8523) );
  OR2_X1 U11119 ( .A1(n14393), .A2(n14305), .ZN(n12085) );
  NAND2_X1 U11120 ( .A1(n14393), .A2(n14305), .ZN(n12084) );
  AND2_X1 U11121 ( .A1(n14389), .A2(n14269), .ZN(n8525) );
  OR2_X1 U11122 ( .A1(n14383), .A2(n14254), .ZN(n13921) );
  INV_X1 U11123 ( .A(n13921), .ZN(n8526) );
  NAND2_X1 U11124 ( .A1(n14383), .A2(n14254), .ZN(n13920) );
  XNOR2_X1 U11125 ( .A(n14259), .B(n14268), .ZN(n14250) );
  OR2_X1 U11126 ( .A1(n14259), .A2(n14268), .ZN(n8527) );
  NAND2_X1 U11127 ( .A1(n14247), .A2(n8527), .ZN(n14228) );
  XNOR2_X1 U11128 ( .A(n14372), .B(n14253), .ZN(n14227) );
  NAND2_X1 U11129 ( .A1(n14372), .A2(n14253), .ZN(n8528) );
  AND2_X1 U11130 ( .A1(n14368), .A2(n14231), .ZN(n13900) );
  XNOR2_X1 U11131 ( .A(n14365), .B(n8529), .ZN(n14200) );
  NAND2_X1 U11132 ( .A1(n14199), .A2(n14200), .ZN(n8531) );
  OR2_X1 U11133 ( .A1(n14365), .A2(n13971), .ZN(n8530) );
  NOR2_X1 U11134 ( .A1(n14196), .A2(n13970), .ZN(n8532) );
  INV_X1 U11135 ( .A(n14196), .ZN(n14440) );
  AND2_X1 U11136 ( .A1(n14353), .A2(n13969), .ZN(n8534) );
  OR2_X1 U11137 ( .A1(n14353), .A2(n13969), .ZN(n8533) );
  XNOR2_X1 U11138 ( .A(n14345), .B(n13968), .ZN(n14161) );
  NAND2_X1 U11139 ( .A1(n14345), .A2(n13968), .ZN(n8535) );
  INV_X1 U11140 ( .A(n13924), .ZN(n14139) );
  NAND2_X1 U11141 ( .A1(n14145), .A2(n13967), .ZN(n8536) );
  OR2_X1 U11142 ( .A1(n14129), .A2(n13966), .ZN(n8538) );
  AND2_X1 U11143 ( .A1(n14129), .A2(n13966), .ZN(n8537) );
  INV_X1 U11144 ( .A(n13859), .ZN(n14092) );
  NOR2_X1 U11145 ( .A1(n14092), .A2(n13698), .ZN(n8540) );
  XOR2_X1 U11146 ( .A(n12817), .B(n13927), .Z(n14088) );
  INV_X1 U11147 ( .A(n15655), .ZN(n14347) );
  INV_X1 U11148 ( .A(n14401), .ZN(n8542) );
  NAND2_X1 U11149 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  NAND2_X1 U11150 ( .A1(n8545), .A2(n8544), .ZN(P2_U3525) );
  INV_X1 U11151 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8548) );
  MUX2_X1 U11152 ( .A(n8548), .B(n8547), .S(n15659), .Z(n8551) );
  NAND2_X1 U11153 ( .A1(n8551), .A2(n8550), .ZN(P2_U3493) );
  INV_X1 U11154 ( .A(SI_27_), .ZN(n13551) );
  NAND2_X1 U11155 ( .A1(n8700), .A2(n13551), .ZN(n8557) );
  INV_X1 U11156 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15229) );
  INV_X1 U11157 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12317) );
  MUX2_X1 U11158 ( .A(n15229), .B(n12317), .S(n9647), .Z(n8698) );
  INV_X1 U11159 ( .A(n8698), .ZN(n8556) );
  INV_X1 U11160 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10182) );
  MUX2_X1 U11161 ( .A(n10182), .B(n12319), .S(n10425), .Z(n8560) );
  NAND2_X1 U11162 ( .A1(n8560), .A2(n15944), .ZN(n9588) );
  INV_X1 U11163 ( .A(n8560), .ZN(n8561) );
  NAND2_X1 U11164 ( .A1(n8561), .A2(SI_28_), .ZN(n8562) );
  NAND2_X1 U11165 ( .A1(n9588), .A2(n8562), .ZN(n9589) );
  NAND2_X1 U11166 ( .A1(n12318), .A2(n8102), .ZN(n8564) );
  OR2_X1 U11167 ( .A1(n9606), .A2(n10182), .ZN(n8563) );
  INV_X1 U11168 ( .A(n8722), .ZN(n12850) );
  INV_X1 U11169 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11170 ( .A1(n8566), .A2(n8733), .ZN(n8567) );
  NAND2_X1 U11171 ( .A1(n8725), .A2(n8721), .ZN(n8573) );
  INV_X1 U11172 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n15950) );
  NAND2_X1 U11173 ( .A1(n12832), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U11174 ( .A1(n9609), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8568) );
  OAI211_X1 U11175 ( .C1(n8570), .C2(n15950), .A(n8569), .B(n8568), .ZN(n8571)
         );
  INV_X1 U11176 ( .A(n8571), .ZN(n8572) );
  NOR2_X1 U11177 ( .A1(n14065), .A2(n14239), .ZN(n8574) );
  INV_X1 U11178 ( .A(n13747), .ZN(n13937) );
  XNOR2_X1 U11179 ( .A(n8574), .B(n8587), .ZN(n8575) );
  XNOR2_X1 U11180 ( .A(n14040), .B(n8575), .ZN(n8740) );
  OR2_X1 U11181 ( .A1(n13756), .A2(n8587), .ZN(n13602) );
  AND2_X1 U11182 ( .A1(n13981), .A2(n8582), .ZN(n13679) );
  NAND2_X1 U11183 ( .A1(n13600), .A2(n13679), .ZN(n8576) );
  XNOR2_X1 U11184 ( .A(n8687), .B(n13745), .ZN(n13678) );
  NAND2_X1 U11185 ( .A1(n13673), .A2(n13672), .ZN(n8578) );
  INV_X1 U11186 ( .A(n13679), .ZN(n8577) );
  INV_X1 U11187 ( .A(n13672), .ZN(n8580) );
  INV_X1 U11188 ( .A(n13673), .ZN(n8579) );
  NAND2_X1 U11189 ( .A1(n8580), .A2(n8579), .ZN(n8581) );
  AND2_X1 U11190 ( .A1(n13979), .A2(n8582), .ZN(n8584) );
  XNOR2_X1 U11191 ( .A(n13767), .B(n8587), .ZN(n8583) );
  NAND2_X1 U11192 ( .A1(n8584), .A2(n8583), .ZN(n8588) );
  INV_X1 U11193 ( .A(n8583), .ZN(n10696) );
  INV_X1 U11194 ( .A(n8584), .ZN(n8585) );
  NAND2_X1 U11195 ( .A1(n10696), .A2(n8585), .ZN(n8586) );
  AND2_X1 U11196 ( .A1(n8586), .A2(n8588), .ZN(n10561) );
  NAND2_X1 U11197 ( .A1(n13978), .A2(n8582), .ZN(n8589) );
  INV_X1 U11198 ( .A(n10802), .ZN(n8590) );
  NAND2_X1 U11199 ( .A1(n8590), .A2(n8589), .ZN(n8591) );
  NAND2_X1 U11200 ( .A1(n10689), .A2(n8591), .ZN(n8592) );
  XNOR2_X1 U11201 ( .A(n13726), .B(n8587), .ZN(n8593) );
  NAND2_X1 U11202 ( .A1(n13977), .A2(n8582), .ZN(n8594) );
  XNOR2_X1 U11203 ( .A(n8593), .B(n8594), .ZN(n10803) );
  INV_X1 U11204 ( .A(n8593), .ZN(n8595) );
  NAND2_X1 U11205 ( .A1(n8595), .A2(n8594), .ZN(n8596) );
  XNOR2_X1 U11206 ( .A(n13777), .B(n8587), .ZN(n8597) );
  AND2_X1 U11207 ( .A1(n13976), .A2(n8582), .ZN(n8598) );
  NAND2_X1 U11208 ( .A1(n8597), .A2(n8598), .ZN(n8602) );
  INV_X1 U11209 ( .A(n8597), .ZN(n10982) );
  INV_X1 U11210 ( .A(n8598), .ZN(n8599) );
  NAND2_X1 U11211 ( .A1(n10982), .A2(n8599), .ZN(n8600) );
  NAND2_X1 U11212 ( .A1(n8602), .A2(n8600), .ZN(n10887) );
  XNOR2_X1 U11213 ( .A(n15650), .B(n8687), .ZN(n8603) );
  NOR2_X1 U11214 ( .A1(n11197), .A2(n14239), .ZN(n8604) );
  XNOR2_X1 U11215 ( .A(n8603), .B(n8604), .ZN(n10979) );
  INV_X1 U11216 ( .A(n8603), .ZN(n8605) );
  NAND2_X1 U11217 ( .A1(n8605), .A2(n8604), .ZN(n8606) );
  NAND2_X1 U11218 ( .A1(n10983), .A2(n8606), .ZN(n11193) );
  XNOR2_X1 U11219 ( .A(n13789), .B(n8687), .ZN(n8607) );
  NAND2_X1 U11220 ( .A1(n13974), .A2(n8582), .ZN(n8608) );
  NAND2_X1 U11221 ( .A1(n8607), .A2(n8608), .ZN(n11192) );
  NAND2_X1 U11222 ( .A1(n11193), .A2(n11192), .ZN(n8611) );
  INV_X1 U11223 ( .A(n8607), .ZN(n8610) );
  INV_X1 U11224 ( .A(n8608), .ZN(n8609) );
  NAND2_X1 U11225 ( .A1(n8610), .A2(n8609), .ZN(n11191) );
  XNOR2_X1 U11226 ( .A(n13794), .B(n8687), .ZN(n8612) );
  NAND2_X1 U11227 ( .A1(n13973), .A2(n8582), .ZN(n8613) );
  NAND2_X1 U11228 ( .A1(n8612), .A2(n8613), .ZN(n8619) );
  INV_X1 U11229 ( .A(n8612), .ZN(n8615) );
  INV_X1 U11230 ( .A(n8613), .ZN(n8614) );
  NAND2_X1 U11231 ( .A1(n8615), .A2(n8614), .ZN(n8616) );
  NAND2_X1 U11232 ( .A1(n8619), .A2(n8616), .ZN(n11385) );
  INV_X1 U11233 ( .A(n11385), .ZN(n8617) );
  XNOR2_X1 U11234 ( .A(n14405), .B(n8687), .ZN(n8621) );
  NAND2_X1 U11235 ( .A1(n14303), .A2(n8582), .ZN(n8620) );
  XNOR2_X1 U11236 ( .A(n8621), .B(n8620), .ZN(n11431) );
  XNOR2_X1 U11237 ( .A(n14399), .B(n8587), .ZN(n8624) );
  NAND2_X1 U11238 ( .A1(n13972), .A2(n8582), .ZN(n8622) );
  XNOR2_X1 U11239 ( .A(n8624), .B(n8622), .ZN(n11775) );
  INV_X1 U11240 ( .A(n8622), .ZN(n8623) );
  NAND2_X1 U11241 ( .A1(n8624), .A2(n8623), .ZN(n8625) );
  NAND2_X1 U11242 ( .A1(n8626), .A2(n8625), .ZN(n12133) );
  INV_X1 U11243 ( .A(n12133), .ZN(n8633) );
  XNOR2_X1 U11244 ( .A(n14393), .B(n8687), .ZN(n8627) );
  NAND2_X1 U11245 ( .A1(n14305), .A2(n8582), .ZN(n8628) );
  NAND2_X1 U11246 ( .A1(n8627), .A2(n8628), .ZN(n8634) );
  INV_X1 U11247 ( .A(n8627), .ZN(n8630) );
  INV_X1 U11248 ( .A(n8628), .ZN(n8629) );
  NAND2_X1 U11249 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  NAND2_X1 U11250 ( .A1(n8634), .A2(n8631), .ZN(n12134) );
  INV_X1 U11251 ( .A(n12134), .ZN(n8632) );
  NAND2_X1 U11252 ( .A1(n8633), .A2(n8632), .ZN(n12131) );
  XNOR2_X1 U11253 ( .A(n14389), .B(n8687), .ZN(n8635) );
  NAND2_X1 U11254 ( .A1(n14269), .A2(n8582), .ZN(n8636) );
  XNOR2_X1 U11255 ( .A(n8635), .B(n8636), .ZN(n12125) );
  INV_X1 U11256 ( .A(n8635), .ZN(n8638) );
  INV_X1 U11257 ( .A(n8636), .ZN(n8637) );
  XNOR2_X1 U11258 ( .A(n14383), .B(n8687), .ZN(n8639) );
  NAND2_X1 U11259 ( .A1(n14254), .A2(n8582), .ZN(n8640) );
  NAND2_X1 U11260 ( .A1(n8639), .A2(n8640), .ZN(n8644) );
  INV_X1 U11261 ( .A(n8639), .ZN(n8642) );
  INV_X1 U11262 ( .A(n8640), .ZN(n8641) );
  NAND2_X1 U11263 ( .A1(n8642), .A2(n8641), .ZN(n8643) );
  AND2_X1 U11264 ( .A1(n8644), .A2(n8643), .ZN(n13570) );
  XNOR2_X1 U11265 ( .A(n14259), .B(n8587), .ZN(n8646) );
  AND2_X1 U11266 ( .A1(n14268), .A2(n8582), .ZN(n8647) );
  XNOR2_X1 U11267 ( .A(n14372), .B(n8587), .ZN(n8649) );
  AND2_X1 U11268 ( .A1(n14253), .A2(n8582), .ZN(n8650) );
  AOI21_X1 U11269 ( .B1(n8646), .B2(n8647), .A(n13629), .ZN(n8645) );
  INV_X1 U11270 ( .A(n13629), .ZN(n8648) );
  INV_X1 U11271 ( .A(n8647), .ZN(n13710) );
  AND2_X1 U11272 ( .A1(n8648), .A2(n13710), .ZN(n8653) );
  INV_X1 U11273 ( .A(n8649), .ZN(n8652) );
  INV_X1 U11274 ( .A(n8650), .ZN(n8651) );
  AND2_X1 U11275 ( .A1(n8652), .A2(n8651), .ZN(n13628) );
  AOI21_X1 U11276 ( .B1(n13627), .B2(n8653), .A(n13628), .ZN(n8654) );
  XNOR2_X1 U11277 ( .A(n14368), .B(n8687), .ZN(n8655) );
  NAND2_X1 U11278 ( .A1(n14231), .A2(n8582), .ZN(n8656) );
  NAND2_X1 U11279 ( .A1(n8655), .A2(n8656), .ZN(n8660) );
  INV_X1 U11280 ( .A(n8655), .ZN(n8658) );
  INV_X1 U11281 ( .A(n8656), .ZN(n8657) );
  NAND2_X1 U11282 ( .A1(n8658), .A2(n8657), .ZN(n8659) );
  AND2_X1 U11283 ( .A1(n8660), .A2(n8659), .ZN(n13639) );
  XNOR2_X1 U11284 ( .A(n14365), .B(n8687), .ZN(n8661) );
  NAND2_X1 U11285 ( .A1(n13971), .A2(n8582), .ZN(n8662) );
  XNOR2_X1 U11286 ( .A(n8661), .B(n8662), .ZN(n13689) );
  INV_X1 U11287 ( .A(n8661), .ZN(n8664) );
  INV_X1 U11288 ( .A(n8662), .ZN(n8663) );
  NAND2_X1 U11289 ( .A1(n8664), .A2(n8663), .ZN(n8665) );
  XNOR2_X1 U11290 ( .A(n14353), .B(n8587), .ZN(n13615) );
  AND2_X1 U11291 ( .A1(n13969), .A2(n8582), .ZN(n8669) );
  NAND2_X1 U11292 ( .A1(n13615), .A2(n8669), .ZN(n8668) );
  XNOR2_X1 U11293 ( .A(n14196), .B(n8687), .ZN(n8667) );
  INV_X1 U11294 ( .A(n8667), .ZN(n13612) );
  NAND2_X1 U11295 ( .A1(n13970), .A2(n8582), .ZN(n13616) );
  INV_X1 U11296 ( .A(n13616), .ZN(n8666) );
  NAND2_X1 U11297 ( .A1(n13612), .A2(n8666), .ZN(n13592) );
  NAND2_X1 U11298 ( .A1(n8668), .A2(n13592), .ZN(n8673) );
  XNOR2_X1 U11299 ( .A(n14345), .B(n8587), .ZN(n8676) );
  NAND2_X1 U11300 ( .A1(n13968), .A2(n8582), .ZN(n8674) );
  XNOR2_X1 U11301 ( .A(n8676), .B(n8674), .ZN(n13617) );
  AND2_X1 U11302 ( .A1(n8667), .A2(n13616), .ZN(n13593) );
  NAND2_X1 U11303 ( .A1(n8668), .A2(n13593), .ZN(n8671) );
  INV_X1 U11304 ( .A(n13615), .ZN(n8670) );
  INV_X1 U11305 ( .A(n8669), .ZN(n13614) );
  NAND2_X1 U11306 ( .A1(n8670), .A2(n13614), .ZN(n13618) );
  AND3_X1 U11307 ( .A1(n13617), .A2(n8671), .A3(n13618), .ZN(n8672) );
  INV_X1 U11308 ( .A(n8674), .ZN(n8675) );
  NAND2_X1 U11309 ( .A1(n8676), .A2(n8675), .ZN(n8677) );
  XNOR2_X1 U11310 ( .A(n14145), .B(n8687), .ZN(n8680) );
  XNOR2_X1 U11311 ( .A(n14129), .B(n8587), .ZN(n13582) );
  AND2_X1 U11312 ( .A1(n13967), .A2(n8582), .ZN(n13579) );
  INV_X1 U11313 ( .A(n8678), .ZN(n8679) );
  NAND2_X1 U11314 ( .A1(n13661), .A2(n8679), .ZN(n8686) );
  AND2_X1 U11315 ( .A1(n13966), .A2(n8582), .ZN(n8683) );
  INV_X1 U11316 ( .A(n8680), .ZN(n8681) );
  AND2_X1 U11317 ( .A1(n8682), .A2(n8681), .ZN(n13580) );
  OAI21_X1 U11318 ( .B1(n8683), .B2(n13582), .A(n13580), .ZN(n8685) );
  INV_X1 U11319 ( .A(n8683), .ZN(n13585) );
  NAND2_X1 U11320 ( .A1(n13582), .A2(n8683), .ZN(n8684) );
  XNOR2_X1 U11321 ( .A(n14109), .B(n8687), .ZN(n12895) );
  NAND2_X1 U11322 ( .A1(n13965), .A2(n8582), .ZN(n8688) );
  NOR2_X1 U11323 ( .A1(n12895), .A2(n8688), .ZN(n8689) );
  AOI21_X1 U11324 ( .B1(n12895), .B2(n8688), .A(n8689), .ZN(n13644) );
  INV_X1 U11325 ( .A(n8689), .ZN(n8694) );
  XNOR2_X1 U11326 ( .A(n13859), .B(n8587), .ZN(n8690) );
  AND2_X1 U11327 ( .A1(n13964), .A2(n8582), .ZN(n8691) );
  NAND2_X1 U11328 ( .A1(n8690), .A2(n8691), .ZN(n8695) );
  INV_X1 U11329 ( .A(n8690), .ZN(n13699) );
  INV_X1 U11330 ( .A(n8691), .ZN(n8692) );
  NAND2_X1 U11331 ( .A1(n13699), .A2(n8692), .ZN(n8693) );
  NAND2_X1 U11332 ( .A1(n8695), .A2(n8693), .ZN(n12894) );
  XNOR2_X1 U11333 ( .A(n14082), .B(n8587), .ZN(n8697) );
  NAND2_X1 U11334 ( .A1(n13963), .A2(n8582), .ZN(n8696) );
  XNOR2_X1 U11335 ( .A(n8698), .B(SI_27_), .ZN(n8699) );
  NAND2_X1 U11336 ( .A1(n12316), .A2(n8102), .ZN(n8702) );
  OR2_X1 U11337 ( .A1(n9606), .A2(n12317), .ZN(n8701) );
  XNOR2_X1 U11338 ( .A(n14413), .B(n8587), .ZN(n8709) );
  NAND2_X1 U11339 ( .A1(n14046), .A2(n8582), .ZN(n8703) );
  NOR2_X1 U11340 ( .A1(n8709), .A2(n8703), .ZN(n8712) );
  AOI21_X1 U11341 ( .B1(n8709), .B2(n8703), .A(n8712), .ZN(n13561) );
  NOR2_X1 U11342 ( .A1(n11227), .A2(n8704), .ZN(n8706) );
  INV_X1 U11343 ( .A(n10483), .ZN(n8707) );
  AND3_X1 U11344 ( .A1(n15615), .A2(n8707), .A3(n15640), .ZN(n8708) );
  INV_X1 U11345 ( .A(n8709), .ZN(n8710) );
  NAND3_X1 U11346 ( .A1(n8710), .A2(n13712), .A3(n14046), .ZN(n8711) );
  INV_X1 U11347 ( .A(n8712), .ZN(n8713) );
  NAND2_X1 U11348 ( .A1(n13560), .A2(n7926), .ZN(n8739) );
  INV_X1 U11349 ( .A(n11235), .ZN(n8714) );
  NOR2_X1 U11350 ( .A1(n8714), .A2(n8541), .ZN(n11529) );
  AND2_X1 U11351 ( .A1(n15615), .A2(n11529), .ZN(n8715) );
  NAND2_X1 U11352 ( .A1(n8726), .A2(n8715), .ZN(n8717) );
  INV_X1 U11353 ( .A(n8727), .ZN(n8716) );
  INV_X1 U11354 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n12849) );
  NAND2_X1 U11355 ( .A1(n9609), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11356 ( .A1(n12833), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8718) );
  OAI211_X1 U11357 ( .C1(n9613), .C2(n12849), .A(n8719), .B(n8718), .ZN(n8720)
         );
  INV_X1 U11358 ( .A(n13952), .ZN(n8723) );
  AND2_X1 U11359 ( .A1(n15615), .A2(n8723), .ZN(n8724) );
  NAND2_X1 U11360 ( .A1(n8726), .A2(n8724), .ZN(n13703) );
  OR2_X1 U11361 ( .A1(n13703), .A2(n14118), .ZN(n13718) );
  INV_X1 U11362 ( .A(n8725), .ZN(n14051) );
  INV_X1 U11363 ( .A(n8726), .ZN(n8728) );
  NAND2_X1 U11364 ( .A1(n8728), .A2(n8727), .ZN(n8732) );
  AND2_X1 U11365 ( .A1(n8730), .A2(n8729), .ZN(n8731) );
  NAND2_X1 U11366 ( .A1(n8732), .A2(n8731), .ZN(n10539) );
  OAI22_X1 U11367 ( .A1(n14047), .A2(n13718), .B1(n14051), .B2(n13717), .ZN(
        n8735) );
  OAI22_X1 U11368 ( .A1(n13866), .A2(n13587), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8733), .ZN(n8734) );
  NOR2_X1 U11369 ( .A1(n8735), .A2(n8734), .ZN(n8736) );
  NOR2_X1 U11370 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n8747) );
  NAND4_X1 U11371 ( .A1(n8747), .A2(n8746), .A3(n8745), .A4(n9004), .ZN(n8763)
         );
  INV_X1 U11372 ( .A(n8763), .ZN(n8755) );
  INV_X2 U11373 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14653) );
  NOR2_X1 U11374 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8752) );
  NAND4_X1 U11375 ( .A1(n8752), .A2(n8751), .A3(n8750), .A4(n6774), .ZN(n8753)
         );
  NAND2_X1 U11376 ( .A1(n8757), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8758) );
  MUX2_X1 U11377 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8758), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n8760) );
  NAND2_X1 U11378 ( .A1(n14477), .A2(n8868), .ZN(n8762) );
  OR2_X1 U11379 ( .A1(n8872), .A2(n15233), .ZN(n8761) );
  NAND2_X1 U11380 ( .A1(n8802), .A2(n8764), .ZN(n8775) );
  INV_X1 U11381 ( .A(n8769), .ZN(n8767) );
  INV_X1 U11382 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U11383 ( .A1(n8767), .A2(n8766), .ZN(n8772) );
  NAND2_X1 U11384 ( .A1(n8772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8768) );
  XNOR2_X1 U11385 ( .A(n8768), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U11386 ( .A1(n8769), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8770) );
  MUX2_X1 U11387 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8770), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8771) );
  NAND2_X1 U11388 ( .A1(n6616), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U11389 ( .A1(n8775), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8776) );
  MUX2_X1 U11390 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8776), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8777) );
  NAND2_X1 U11391 ( .A1(n8777), .A2(n6616), .ZN(n12558) );
  NAND2_X2 U11392 ( .A1(n8853), .A2(n8807), .ZN(n8818) );
  INV_X2 U11393 ( .A(n8818), .ZN(n9323) );
  NAND2_X1 U11394 ( .A1(n14860), .A2(n9323), .ZN(n8801) );
  NAND3_X1 U11395 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8945) );
  INV_X1 U11396 ( .A(n8945), .ZN(n8778) );
  NAND2_X1 U11397 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n8785) );
  INV_X1 U11398 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14589) );
  INV_X1 U11399 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14501) );
  INV_X1 U11400 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14608) );
  NAND2_X1 U11401 ( .A1(n9250), .A2(n14608), .ZN(n8788) );
  NAND2_X1 U11402 ( .A1(n14857), .A2(n9310), .ZN(n8799) );
  NAND2_X2 U11403 ( .A1(n8792), .A2(n15227), .ZN(n12714) );
  INV_X1 U11404 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8796) );
  NAND2_X2 U11405 ( .A1(n15224), .A2(n15227), .ZN(n8931) );
  NAND2_X1 U11406 ( .A1(n9311), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11407 ( .A1(n8947), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8794) );
  OAI211_X1 U11408 ( .C1(n12714), .C2(n8796), .A(n8795), .B(n8794), .ZN(n8797)
         );
  INV_X1 U11409 ( .A(n8797), .ZN(n8798) );
  NAND2_X1 U11410 ( .A1(n14870), .A2(n8854), .ZN(n8800) );
  NAND2_X1 U11411 ( .A1(n8801), .A2(n8800), .ZN(n8808) );
  NAND2_X1 U11412 ( .A1(n15237), .A2(n12556), .ZN(n12555) );
  XNOR2_X1 U11413 ( .A(n8808), .B(n10580), .ZN(n9266) );
  AOI22_X1 U11414 ( .A1(n14860), .A2(n8854), .B1(n9318), .B2(n14870), .ZN(
        n9263) );
  INV_X1 U11415 ( .A(n9263), .ZN(n9265) );
  NAND2_X1 U11416 ( .A1(n9202), .A2(n14589), .ZN(n8811) );
  NAND2_X1 U11417 ( .A1(n9217), .A2(n8811), .ZN(n14931) );
  OR2_X1 U11418 ( .A1(n14931), .A2(n9273), .ZN(n8817) );
  INV_X1 U11419 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14929) );
  NAND2_X1 U11420 ( .A1(n9311), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8814) );
  NAND2_X1 U11421 ( .A1(n8947), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8813) );
  OAI211_X1 U11422 ( .C1(n14929), .C2(n12714), .A(n8814), .B(n8813), .ZN(n8815) );
  INV_X1 U11423 ( .A(n8815), .ZN(n8816) );
  OAI22_X1 U11424 ( .A1(n15129), .A2(n8958), .B1(n14944), .B2(n9136), .ZN(
        n9214) );
  OAI22_X1 U11425 ( .A1(n15129), .A2(n8818), .B1(n14944), .B2(n8958), .ZN(
        n8819) );
  XNOR2_X1 U11426 ( .A(n8819), .B(n10580), .ZN(n9213) );
  NAND2_X1 U11427 ( .A1(n11202), .A2(n8868), .ZN(n8821) );
  OR2_X1 U11428 ( .A1(n8872), .A2(n11203), .ZN(n8820) );
  INV_X1 U11429 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14579) );
  NAND2_X1 U11430 ( .A1(n8837), .A2(n14579), .ZN(n8822) );
  NAND2_X1 U11431 ( .A1(n9200), .A2(n8822), .ZN(n14968) );
  OR2_X1 U11432 ( .A1(n14968), .A2(n9273), .ZN(n8828) );
  INV_X1 U11433 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U11434 ( .A1(n8947), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U11435 ( .A1(n9311), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8823) );
  OAI211_X1 U11436 ( .C1(n12714), .C2(n8825), .A(n8824), .B(n8823), .ZN(n8826)
         );
  INV_X1 U11437 ( .A(n8826), .ZN(n8827) );
  NAND2_X1 U11438 ( .A1(n8828), .A2(n8827), .ZN(n14637) );
  AND2_X1 U11439 ( .A1(n14637), .A2(n9318), .ZN(n8829) );
  AOI21_X1 U11440 ( .B1(n15143), .B2(n8854), .A(n8829), .ZN(n9194) );
  INV_X1 U11441 ( .A(n9194), .ZN(n9196) );
  AOI22_X1 U11442 ( .A1(n15143), .A2(n9323), .B1(n8854), .B2(n14637), .ZN(
        n8830) );
  XNOR2_X1 U11443 ( .A(n8830), .B(n10580), .ZN(n9193) );
  INV_X1 U11444 ( .A(n9193), .ZN(n9195) );
  NAND2_X1 U11445 ( .A1(n8831), .A2(n8868), .ZN(n8834) );
  AOI22_X1 U11446 ( .A1(n9175), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14809), 
        .B2(n9176), .ZN(n8833) );
  INV_X1 U11447 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8836) );
  INV_X1 U11448 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8835) );
  OAI21_X1 U11449 ( .B1(n9179), .B2(n8836), .A(n8835), .ZN(n8838) );
  NAND2_X1 U11450 ( .A1(n8838), .A2(n8837), .ZN(n14986) );
  OR2_X1 U11451 ( .A1(n14986), .A2(n9273), .ZN(n8843) );
  INV_X1 U11452 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14801) );
  NAND2_X1 U11453 ( .A1(n8947), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8840) );
  NAND2_X1 U11454 ( .A1(n9311), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8839) );
  OAI211_X1 U11455 ( .C1(n12714), .C2(n14801), .A(n8840), .B(n8839), .ZN(n8841) );
  INV_X1 U11456 ( .A(n8841), .ZN(n8842) );
  NAND2_X1 U11457 ( .A1(n8843), .A2(n8842), .ZN(n14993) );
  AND2_X1 U11458 ( .A1(n14993), .A2(n9318), .ZN(n8844) );
  AOI21_X1 U11459 ( .B1(n15150), .B2(n8854), .A(n8844), .ZN(n9192) );
  AOI22_X1 U11460 ( .A1(n15150), .A2(n9323), .B1(n8854), .B2(n14993), .ZN(
        n8845) );
  XNOR2_X1 U11461 ( .A(n8845), .B(n10580), .ZN(n9191) );
  NAND2_X1 U11462 ( .A1(n9310), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U11463 ( .A1(n8947), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8850) );
  INV_X1 U11464 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n8846) );
  OR2_X1 U11465 ( .A1(n8931), .A2(n8846), .ZN(n8849) );
  INV_X1 U11466 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8847) );
  OR2_X1 U11467 ( .A1(n12714), .A2(n8847), .ZN(n8848) );
  INV_X1 U11468 ( .A(n12041), .ZN(n12036) );
  NAND2_X1 U11469 ( .A1(n10425), .A2(SI_0_), .ZN(n8852) );
  XNOR2_X1 U11470 ( .A(n8852), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15239) );
  INV_X1 U11471 ( .A(n8853), .ZN(n8856) );
  NAND2_X1 U11472 ( .A1(n9323), .A2(n12038), .ZN(n8859) );
  NAND2_X1 U11473 ( .A1(n8856), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8857) );
  INV_X1 U11474 ( .A(n11001), .ZN(n8860) );
  NAND2_X1 U11475 ( .A1(n8861), .A2(n8860), .ZN(n10998) );
  NAND2_X1 U11476 ( .A1(n11001), .A2(n10580), .ZN(n8862) );
  NAND2_X1 U11477 ( .A1(n8947), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8866) );
  INV_X1 U11478 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8863) );
  OR2_X1 U11479 ( .A1(n8931), .A2(n8863), .ZN(n8865) );
  INV_X1 U11480 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10586) );
  OR2_X1 U11481 ( .A1(n12714), .A2(n10586), .ZN(n8864) );
  NAND4_X2 U11482 ( .A1(n8867), .A2(n8866), .A3(n8865), .A4(n8864), .ZN(n11669) );
  NAND2_X1 U11483 ( .A1(n8868), .A2(n8869), .ZN(n8874) );
  NAND2_X1 U11484 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8871) );
  OAI22_X1 U11485 ( .A1(n12813), .A2(n8958), .B1(n8818), .B2(n15410), .ZN(
        n8875) );
  XNOR2_X1 U11486 ( .A(n8875), .B(n9321), .ZN(n8880) );
  INV_X1 U11487 ( .A(n8880), .ZN(n8878) );
  NOR2_X1 U11488 ( .A1(n8958), .A2(n15410), .ZN(n8876) );
  AOI21_X1 U11489 ( .B1(n6543), .B2(n11669), .A(n8876), .ZN(n8879) );
  INV_X1 U11490 ( .A(n8879), .ZN(n8877) );
  NAND2_X1 U11491 ( .A1(n8878), .A2(n8877), .ZN(n8881) );
  NAND2_X1 U11492 ( .A1(n8880), .A2(n8879), .ZN(n8882) );
  NAND2_X1 U11493 ( .A1(n9310), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8885) );
  NAND2_X1 U11494 ( .A1(n8947), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8884) );
  INV_X1 U11495 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15703) );
  OR2_X1 U11496 ( .A1(n8931), .A2(n15703), .ZN(n8883) );
  INV_X1 U11497 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10587) );
  NAND4_X1 U11498 ( .A1(n8885), .A2(n8884), .A3(n8883), .A4(n6610), .ZN(n14650) );
  INV_X1 U11499 ( .A(n14650), .ZN(n12570) );
  NAND2_X1 U11500 ( .A1(n10348), .A2(n8868), .ZN(n8888) );
  NAND2_X1 U11501 ( .A1(n8900), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8886) );
  OAI22_X1 U11502 ( .A1(n12570), .A2(n8958), .B1(n8818), .B2(n15418), .ZN(
        n8889) );
  XNOR2_X1 U11503 ( .A(n8889), .B(n9321), .ZN(n8892) );
  OAI22_X1 U11504 ( .A1(n9136), .A2(n12570), .B1(n15418), .B2(n8958), .ZN(
        n8890) );
  XNOR2_X1 U11505 ( .A(n8892), .B(n8890), .ZN(n12810) );
  INV_X1 U11506 ( .A(n8890), .ZN(n8891) );
  NAND2_X1 U11507 ( .A1(n8892), .A2(n8891), .ZN(n8893) );
  INV_X1 U11508 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U11509 ( .A1(n9310), .A2(n8894), .ZN(n8899) );
  NAND2_X1 U11510 ( .A1(n8947), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8898) );
  INV_X1 U11511 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10585) );
  OR2_X1 U11512 ( .A1(n12714), .A2(n10585), .ZN(n8897) );
  INV_X1 U11513 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8895) );
  OR2_X1 U11514 ( .A1(n8931), .A2(n8895), .ZN(n8896) );
  NAND2_X1 U11515 ( .A1(n10363), .A2(n8868), .ZN(n8904) );
  OAI21_X1 U11516 ( .B1(n8900), .B2(P1_IR_REG_2__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8901) );
  MUX2_X1 U11517 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8901), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8902) );
  AND2_X1 U11518 ( .A1(n8902), .A2(n8921), .ZN(n14691) );
  AOI22_X1 U11519 ( .A1(n9175), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n9176), .B2(
        n14691), .ZN(n8903) );
  OAI22_X1 U11520 ( .A1(n12812), .A2(n8958), .B1(n8818), .B2(n11674), .ZN(
        n8905) );
  XNOR2_X1 U11521 ( .A(n8905), .B(n10580), .ZN(n8908) );
  OAI22_X1 U11522 ( .A1(n9136), .A2(n12812), .B1(n11674), .B2(n8958), .ZN(
        n8907) );
  XNOR2_X1 U11523 ( .A(n8908), .B(n8907), .ZN(n11013) );
  NAND2_X1 U11524 ( .A1(n8908), .A2(n8907), .ZN(n8909) );
  NAND2_X1 U11525 ( .A1(n8947), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8914) );
  INV_X1 U11526 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8910) );
  XNOR2_X1 U11527 ( .A(n8910), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n15371) );
  NAND2_X1 U11528 ( .A1(n9310), .A2(n15371), .ZN(n8913) );
  INV_X1 U11529 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8911) );
  INV_X1 U11530 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10591) );
  NAND2_X1 U11531 ( .A1(n9318), .A2(n14648), .ZN(n8919) );
  NAND2_X1 U11532 ( .A1(n10350), .A2(n8868), .ZN(n8917) );
  NAND2_X1 U11533 ( .A1(n8921), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8915) );
  XNOR2_X1 U11534 ( .A(n8915), .B(P1_IR_REG_4__SCAN_IN), .ZN(n15339) );
  AOI22_X1 U11535 ( .A1(n9175), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9176), .B2(
        n15339), .ZN(n8916) );
  INV_X1 U11536 ( .A(n15427), .ZN(n14572) );
  NAND2_X1 U11537 ( .A1(n8854), .A2(n14572), .ZN(n8918) );
  NAND2_X1 U11538 ( .A1(n8919), .A2(n8918), .ZN(n11419) );
  OAI22_X1 U11539 ( .A1(n12581), .A2(n8958), .B1(n8818), .B2(n15427), .ZN(
        n8920) );
  XNOR2_X1 U11540 ( .A(n8920), .B(n10580), .ZN(n14567) );
  NAND2_X1 U11541 ( .A1(n10392), .A2(n8868), .ZN(n8926) );
  INV_X1 U11542 ( .A(n8921), .ZN(n8923) );
  INV_X1 U11543 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U11544 ( .A1(n8923), .A2(n8922), .ZN(n8953) );
  NAND2_X1 U11545 ( .A1(n8953), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8924) );
  XNOR2_X1 U11546 ( .A(n8924), .B(P1_IR_REG_5__SCAN_IN), .ZN(n14706) );
  AOI22_X1 U11547 ( .A1(n9175), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9176), .B2(
        n14706), .ZN(n8925) );
  INV_X1 U11548 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U11549 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n8927) );
  NAND2_X1 U11550 ( .A1(n8928), .A2(n8927), .ZN(n8929) );
  AND2_X1 U11551 ( .A1(n8945), .A2(n8929), .ZN(n12065) );
  NAND2_X1 U11552 ( .A1(n9310), .A2(n12065), .ZN(n8935) );
  NAND2_X1 U11553 ( .A1(n8947), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8934) );
  INV_X1 U11554 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10594) );
  OR2_X1 U11555 ( .A1(n12714), .A2(n10594), .ZN(n8933) );
  INV_X1 U11556 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n8930) );
  OR2_X1 U11557 ( .A1(n8931), .A2(n8930), .ZN(n8932) );
  NAND4_X1 U11558 ( .A1(n8935), .A2(n8934), .A3(n8933), .A4(n8932), .ZN(n14647) );
  INV_X1 U11559 ( .A(n14647), .ZN(n11687) );
  OAI22_X1 U11560 ( .A1(n15434), .A2(n8818), .B1(n8958), .B2(n11687), .ZN(
        n8936) );
  XNOR2_X1 U11561 ( .A(n8936), .B(n9321), .ZN(n8939) );
  INV_X1 U11562 ( .A(n15434), .ZN(n12586) );
  AOI22_X1 U11563 ( .A1(n9318), .A2(n14647), .B1(n8854), .B2(n12586), .ZN(
        n8940) );
  NAND2_X1 U11564 ( .A1(n8939), .A2(n8940), .ZN(n11422) );
  NAND3_X1 U11565 ( .A1(n11422), .A2(n14567), .A3(n11419), .ZN(n8943) );
  INV_X1 U11566 ( .A(n8939), .ZN(n8942) );
  INV_X1 U11567 ( .A(n8940), .ZN(n8941) );
  NAND2_X1 U11568 ( .A1(n8942), .A2(n8941), .ZN(n11421) );
  INV_X1 U11569 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U11570 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  AND2_X1 U11571 ( .A1(n8990), .A2(n8946), .ZN(n15358) );
  NAND2_X1 U11572 ( .A1(n9310), .A2(n15358), .ZN(n8952) );
  NAND2_X1 U11573 ( .A1(n8947), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8951) );
  INV_X1 U11574 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10597) );
  OR2_X1 U11575 ( .A1(n12714), .A2(n10597), .ZN(n8950) );
  INV_X1 U11576 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8948) );
  OR2_X1 U11577 ( .A1(n8931), .A2(n8948), .ZN(n8949) );
  NAND4_X1 U11578 ( .A1(n8952), .A2(n8951), .A3(n8950), .A4(n8949), .ZN(n14646) );
  NAND2_X1 U11579 ( .A1(n8963), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8954) );
  XNOR2_X1 U11580 ( .A(n8954), .B(P1_IR_REG_6__SCAN_IN), .ZN(n14716) );
  AOI22_X1 U11581 ( .A1(n9175), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9176), .B2(
        n14716), .ZN(n8955) );
  OAI22_X1 U11582 ( .A1(n12591), .A2(n8958), .B1(n8818), .B2(n15440), .ZN(
        n8957) );
  XNOR2_X1 U11583 ( .A(n8957), .B(n9321), .ZN(n8959) );
  OAI22_X1 U11584 ( .A1(n9136), .A2(n12591), .B1(n15440), .B2(n8958), .ZN(
        n8960) );
  XNOR2_X1 U11585 ( .A(n8959), .B(n8960), .ZN(n11273) );
  INV_X1 U11586 ( .A(n8959), .ZN(n8961) );
  NAND2_X1 U11587 ( .A1(n8961), .A2(n8960), .ZN(n8962) );
  NAND2_X1 U11588 ( .A1(n10390), .A2(n8868), .ZN(n8968) );
  INV_X1 U11589 ( .A(n8963), .ZN(n8965) );
  INV_X1 U11590 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8964) );
  NAND2_X1 U11591 ( .A1(n8965), .A2(n8964), .ZN(n8982) );
  NAND2_X1 U11592 ( .A1(n8982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8966) );
  XNOR2_X1 U11593 ( .A(n8966), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14734) );
  AOI22_X1 U11594 ( .A1(n9175), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9176), .B2(
        n14734), .ZN(n8967) );
  NAND2_X1 U11595 ( .A1(n12598), .A2(n9323), .ZN(n8975) );
  XNOR2_X1 U11596 ( .A(n8990), .B(P1_REG3_REG_7__SCAN_IN), .ZN(n11699) );
  NAND2_X1 U11597 ( .A1(n9310), .A2(n11699), .ZN(n8973) );
  NAND2_X1 U11598 ( .A1(n8947), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8972) );
  INV_X1 U11599 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11692) );
  OR2_X1 U11600 ( .A1(n12714), .A2(n11692), .ZN(n8971) );
  INV_X1 U11601 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8969) );
  OR2_X1 U11602 ( .A1(n8931), .A2(n8969), .ZN(n8970) );
  NAND4_X1 U11603 ( .A1(n8973), .A2(n8972), .A3(n8971), .A4(n8970), .ZN(n14645) );
  NAND2_X1 U11604 ( .A1(n8854), .A2(n14645), .ZN(n8974) );
  NAND2_X1 U11605 ( .A1(n8975), .A2(n8974), .ZN(n8976) );
  XNOR2_X1 U11606 ( .A(n8976), .B(n9321), .ZN(n8978) );
  INV_X1 U11607 ( .A(n14645), .ZN(n12597) );
  NAND2_X1 U11608 ( .A1(n12598), .A2(n8854), .ZN(n8977) );
  OAI21_X1 U11609 ( .B1(n9136), .B2(n12597), .A(n8977), .ZN(n8979) );
  XNOR2_X1 U11610 ( .A(n8978), .B(n8979), .ZN(n11378) );
  INV_X1 U11611 ( .A(n8978), .ZN(n8980) );
  NAND2_X1 U11612 ( .A1(n8980), .A2(n8979), .ZN(n8981) );
  NAND2_X1 U11613 ( .A1(n10441), .A2(n8868), .ZN(n8987) );
  INV_X1 U11614 ( .A(n8982), .ZN(n8984) );
  INV_X1 U11615 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U11616 ( .A1(n8984), .A2(n8983), .ZN(n9001) );
  NAND2_X1 U11617 ( .A1(n9001), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8985) );
  XNOR2_X1 U11618 ( .A(n8985), .B(P1_IR_REG_8__SCAN_IN), .ZN(n14750) );
  AOI22_X1 U11619 ( .A1(n9175), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9176), .B2(
        n14750), .ZN(n8986) );
  NAND2_X1 U11620 ( .A1(n8987), .A2(n8986), .ZN(n12607) );
  NAND2_X1 U11621 ( .A1(n12607), .A2(n9323), .ZN(n8998) );
  INV_X1 U11622 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8989) );
  INV_X1 U11623 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8988) );
  OAI21_X1 U11624 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(n8991) );
  AND2_X1 U11625 ( .A1(n9010), .A2(n8991), .ZN(n11829) );
  NAND2_X1 U11626 ( .A1(n9310), .A2(n11829), .ZN(n8996) );
  NAND2_X1 U11627 ( .A1(n8947), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8995) );
  INV_X1 U11628 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11711) );
  OR2_X1 U11629 ( .A1(n12714), .A2(n11711), .ZN(n8994) );
  INV_X1 U11630 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8992) );
  OR2_X1 U11631 ( .A1(n8931), .A2(n8992), .ZN(n8993) );
  NAND4_X1 U11632 ( .A1(n8996), .A2(n8995), .A3(n8994), .A4(n8993), .ZN(n14644) );
  NAND2_X1 U11633 ( .A1(n8854), .A2(n14644), .ZN(n8997) );
  NAND2_X1 U11634 ( .A1(n8998), .A2(n8997), .ZN(n8999) );
  XNOR2_X1 U11635 ( .A(n8999), .B(n10580), .ZN(n9040) );
  INV_X1 U11636 ( .A(n14644), .ZN(n12606) );
  NAND2_X1 U11637 ( .A1(n12607), .A2(n8854), .ZN(n9000) );
  OAI21_X1 U11638 ( .B1(n9136), .B2(n12606), .A(n9000), .ZN(n9039) );
  XNOR2_X1 U11639 ( .A(n9040), .B(n9039), .ZN(n11825) );
  NAND2_X1 U11640 ( .A1(n10454), .A2(n8868), .ZN(n9008) );
  NAND2_X1 U11641 ( .A1(n9003), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9006) );
  INV_X1 U11642 ( .A(n9003), .ZN(n9005) );
  NAND2_X1 U11643 ( .A1(n9005), .A2(n9004), .ZN(n9020) );
  AOI22_X1 U11644 ( .A1(n9175), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10663), 
        .B2(n9176), .ZN(n9007) );
  NAND2_X1 U11645 ( .A1(n12603), .A2(n9323), .ZN(n9018) );
  INV_X1 U11646 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U11647 ( .A1(n9010), .A2(n9009), .ZN(n9011) );
  AND2_X1 U11648 ( .A1(n9024), .A2(n9011), .ZN(n11918) );
  NAND2_X1 U11649 ( .A1(n9310), .A2(n11918), .ZN(n9016) );
  NAND2_X1 U11650 ( .A1(n8947), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9015) );
  INV_X1 U11651 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11741) );
  OR2_X1 U11652 ( .A1(n12714), .A2(n11741), .ZN(n9014) );
  INV_X1 U11653 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9012) );
  OR2_X1 U11654 ( .A1(n8931), .A2(n9012), .ZN(n9013) );
  NAND4_X1 U11655 ( .A1(n9016), .A2(n9015), .A3(n9014), .A4(n9013), .ZN(n14643) );
  NAND2_X1 U11656 ( .A1(n8854), .A2(n14643), .ZN(n9017) );
  NAND2_X1 U11657 ( .A1(n9018), .A2(n9017), .ZN(n9019) );
  XNOR2_X1 U11658 ( .A(n9019), .B(n10580), .ZN(n9036) );
  AOI22_X1 U11659 ( .A1(n12603), .A2(n8854), .B1(n9318), .B2(n14643), .ZN(
        n9037) );
  XNOR2_X1 U11660 ( .A(n9036), .B(n9037), .ZN(n11917) );
  INV_X1 U11661 ( .A(n11917), .ZN(n9041) );
  OR2_X1 U11662 ( .A1(n11825), .A2(n9041), .ZN(n11885) );
  NAND2_X1 U11663 ( .A1(n10447), .A2(n8868), .ZN(n9023) );
  NAND2_X1 U11664 ( .A1(n9020), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9021) );
  XNOR2_X1 U11665 ( .A(n9021), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U11666 ( .A1(n10673), .A2(n9176), .B1(n9175), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U11667 ( .A1(n12600), .A2(n9323), .ZN(n9032) );
  NAND2_X1 U11668 ( .A1(n9024), .A2(n10678), .ZN(n9025) );
  AND2_X1 U11669 ( .A1(n9049), .A2(n9025), .ZN(n11893) );
  NAND2_X1 U11670 ( .A1(n9310), .A2(n11893), .ZN(n9030) );
  NAND2_X1 U11671 ( .A1(n8947), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9029) );
  INV_X1 U11672 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10606) );
  OR2_X1 U11673 ( .A1(n12714), .A2(n10606), .ZN(n9028) );
  INV_X1 U11674 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9026) );
  OR2_X1 U11675 ( .A1(n8931), .A2(n9026), .ZN(n9027) );
  NAND4_X1 U11676 ( .A1(n9030), .A2(n9029), .A3(n9028), .A4(n9027), .ZN(n14642) );
  NAND2_X1 U11677 ( .A1(n8854), .A2(n14642), .ZN(n9031) );
  NAND2_X1 U11678 ( .A1(n9032), .A2(n9031), .ZN(n9033) );
  XNOR2_X1 U11679 ( .A(n9033), .B(n9321), .ZN(n9035) );
  AOI22_X1 U11680 ( .A1(n12600), .A2(n8854), .B1(n9318), .B2(n14642), .ZN(
        n9034) );
  XNOR2_X1 U11681 ( .A(n9035), .B(n9034), .ZN(n11888) );
  INV_X1 U11682 ( .A(n11888), .ZN(n9043) );
  INV_X1 U11683 ( .A(n9036), .ZN(n9038) );
  NAND2_X1 U11684 ( .A1(n9038), .A2(n9037), .ZN(n9042) );
  OR2_X1 U11685 ( .A1(n9040), .A2(n9039), .ZN(n11911) );
  OR2_X1 U11686 ( .A1(n9041), .A2(n11911), .ZN(n11913) );
  AND2_X1 U11687 ( .A1(n9042), .A2(n11913), .ZN(n11887) );
  AND2_X1 U11688 ( .A1(n11887), .A2(n9043), .ZN(n11890) );
  NAND2_X1 U11689 ( .A1(n10444), .A2(n8868), .ZN(n9048) );
  INV_X1 U11690 ( .A(n8803), .ZN(n9044) );
  NAND2_X1 U11691 ( .A1(n9044), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9045) );
  MUX2_X1 U11692 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9045), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n9046) );
  AOI22_X1 U11693 ( .A1(n9175), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9176), 
        .B2(n14768), .ZN(n9047) );
  NAND2_X1 U11694 ( .A1(n12619), .A2(n9323), .ZN(n9057) );
  NAND2_X1 U11695 ( .A1(n9049), .A2(n15783), .ZN(n9050) );
  AND2_X1 U11696 ( .A1(n9066), .A2(n9050), .ZN(n12117) );
  NAND2_X1 U11697 ( .A1(n9310), .A2(n12117), .ZN(n9055) );
  NAND2_X1 U11698 ( .A1(n8947), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9054) );
  INV_X1 U11699 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10609) );
  OR2_X1 U11700 ( .A1(n12714), .A2(n10609), .ZN(n9053) );
  INV_X1 U11701 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9051) );
  OR2_X1 U11702 ( .A1(n8931), .A2(n9051), .ZN(n9052) );
  NAND4_X1 U11703 ( .A1(n9055), .A2(n9054), .A3(n9053), .A4(n9052), .ZN(n14641) );
  NAND2_X1 U11704 ( .A1(n8854), .A2(n14641), .ZN(n9056) );
  NAND2_X1 U11705 ( .A1(n9057), .A2(n9056), .ZN(n9058) );
  XNOR2_X1 U11706 ( .A(n9058), .B(n9321), .ZN(n9060) );
  AOI22_X1 U11707 ( .A1(n12619), .A2(n8854), .B1(n9318), .B2(n14641), .ZN(
        n9059) );
  NAND2_X1 U11708 ( .A1(n9060), .A2(n9059), .ZN(n9061) );
  XNOR2_X1 U11709 ( .A(n9060), .B(n9059), .ZN(n12021) );
  NAND2_X1 U11710 ( .A1(n9061), .A2(n12021), .ZN(n9062) );
  NAND2_X1 U11711 ( .A1(n10458), .A2(n8868), .ZN(n9065) );
  XNOR2_X1 U11712 ( .A(n9063), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U11713 ( .A1(n9175), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9176), 
        .B2(n10815), .ZN(n9064) );
  NAND2_X1 U11714 ( .A1(n15188), .A2(n9323), .ZN(n9074) );
  INV_X1 U11715 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n12030) );
  NAND2_X1 U11716 ( .A1(n9066), .A2(n12030), .ZN(n9067) );
  AND2_X1 U11717 ( .A1(n9085), .A2(n9067), .ZN(n12033) );
  NAND2_X1 U11718 ( .A1(n9310), .A2(n12033), .ZN(n9072) );
  NAND2_X1 U11719 ( .A1(n8947), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9071) );
  INV_X1 U11720 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11944) );
  OR2_X1 U11721 ( .A1(n12714), .A2(n11944), .ZN(n9070) );
  INV_X1 U11722 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9068) );
  OR2_X1 U11723 ( .A1(n8931), .A2(n9068), .ZN(n9069) );
  NAND4_X1 U11724 ( .A1(n9072), .A2(n9071), .A3(n9070), .A4(n9069), .ZN(n14640) );
  NAND2_X1 U11725 ( .A1(n8854), .A2(n14640), .ZN(n9073) );
  NAND2_X1 U11726 ( .A1(n9074), .A2(n9073), .ZN(n9075) );
  XNOR2_X1 U11727 ( .A(n9075), .B(n10580), .ZN(n9079) );
  INV_X1 U11728 ( .A(n14640), .ZN(n12638) );
  NOR2_X1 U11729 ( .A1(n9136), .A2(n12638), .ZN(n9076) );
  AOI21_X1 U11730 ( .B1(n15188), .B2(n8854), .A(n9076), .ZN(n9077) );
  XNOR2_X1 U11731 ( .A(n9079), .B(n9077), .ZN(n12028) );
  INV_X1 U11732 ( .A(n9077), .ZN(n9078) );
  NAND2_X1 U11733 ( .A1(n9079), .A2(n9078), .ZN(n9080) );
  NAND2_X1 U11734 ( .A1(n10464), .A2(n8868), .ZN(n9083) );
  NAND2_X1 U11735 ( .A1(n9100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9081) );
  XNOR2_X1 U11736 ( .A(n9081), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U11737 ( .A1(n9175), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9176), 
        .B2(n10855), .ZN(n9082) );
  NAND2_X1 U11738 ( .A1(n15183), .A2(n9323), .ZN(n9093) );
  INV_X1 U11739 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U11740 ( .A1(n9085), .A2(n9084), .ZN(n9086) );
  AND2_X1 U11741 ( .A1(n9105), .A2(n9086), .ZN(n12175) );
  NAND2_X1 U11742 ( .A1(n9310), .A2(n12175), .ZN(n9091) );
  NAND2_X1 U11743 ( .A1(n8947), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9090) );
  INV_X1 U11744 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12114) );
  OR2_X1 U11745 ( .A1(n12714), .A2(n12114), .ZN(n9089) );
  INV_X1 U11746 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9087) );
  OR2_X1 U11747 ( .A1(n8931), .A2(n9087), .ZN(n9088) );
  NAND4_X1 U11748 ( .A1(n9091), .A2(n9090), .A3(n9089), .A4(n9088), .ZN(n14639) );
  NAND2_X1 U11749 ( .A1(n8854), .A2(n14639), .ZN(n9092) );
  NAND2_X1 U11750 ( .A1(n9093), .A2(n9092), .ZN(n9094) );
  XNOR2_X1 U11751 ( .A(n9094), .B(n10580), .ZN(n9098) );
  INV_X1 U11752 ( .A(n14639), .ZN(n11974) );
  NOR2_X1 U11753 ( .A1(n9136), .A2(n11974), .ZN(n9095) );
  AOI21_X1 U11754 ( .B1(n15183), .B2(n8854), .A(n9095), .ZN(n9096) );
  XNOR2_X1 U11755 ( .A(n9098), .B(n9096), .ZN(n12172) );
  INV_X1 U11756 ( .A(n9096), .ZN(n9097) );
  NAND2_X1 U11757 ( .A1(n9098), .A2(n9097), .ZN(n9099) );
  NAND2_X1 U11758 ( .A1(n10655), .A2(n8868), .ZN(n9103) );
  NAND2_X1 U11759 ( .A1(n9120), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9101) );
  XNOR2_X1 U11760 ( .A(n9101), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U11761 ( .A1(n9175), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9176), 
        .B2(n11335), .ZN(n9102) );
  NAND2_X1 U11762 ( .A1(n15175), .A2(n9323), .ZN(n9113) );
  NAND2_X1 U11763 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  AND2_X1 U11764 ( .A1(n9127), .A2(n9106), .ZN(n14493) );
  NAND2_X1 U11765 ( .A1(n9310), .A2(n14493), .ZN(n9111) );
  NAND2_X1 U11766 ( .A1(n8947), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9110) );
  INV_X1 U11767 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10814) );
  OR2_X1 U11768 ( .A1(n12714), .A2(n10814), .ZN(n9109) );
  INV_X1 U11769 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9107) );
  OR2_X1 U11770 ( .A1(n8931), .A2(n9107), .ZN(n9108) );
  NAND4_X1 U11771 ( .A1(n9111), .A2(n9110), .A3(n9109), .A4(n9108), .ZN(n14638) );
  NAND2_X1 U11772 ( .A1(n8854), .A2(n14638), .ZN(n9112) );
  NAND2_X1 U11773 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  XNOR2_X1 U11774 ( .A(n9114), .B(n9321), .ZN(n9118) );
  INV_X1 U11775 ( .A(n14638), .ZN(n11976) );
  NOR2_X1 U11776 ( .A1(n9136), .A2(n11976), .ZN(n9115) );
  AOI21_X1 U11777 ( .B1(n15175), .B2(n8854), .A(n9115), .ZN(n9117) );
  XNOR2_X1 U11778 ( .A(n9118), .B(n9117), .ZN(n14492) );
  INV_X1 U11779 ( .A(n14492), .ZN(n9116) );
  NAND2_X1 U11780 ( .A1(n9118), .A2(n9117), .ZN(n9119) );
  NAND2_X1 U11781 ( .A1(n10704), .A2(n8868), .ZN(n9125) );
  INV_X1 U11782 ( .A(n9120), .ZN(n9122) );
  INV_X1 U11783 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U11784 ( .A1(n9122), .A2(n9121), .ZN(n9138) );
  NAND2_X1 U11785 ( .A1(n9138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9123) );
  XNOR2_X1 U11786 ( .A(n9123), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U11787 ( .A1(n11344), .A2(n9176), .B1(n9175), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U11788 ( .A1(n15171), .A2(n9323), .ZN(n9134) );
  INV_X1 U11789 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U11790 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  NAND2_X1 U11791 ( .A1(n9147), .A2(n9128), .ZN(n14625) );
  OR2_X1 U11792 ( .A1(n14625), .A2(n9273), .ZN(n9132) );
  NAND2_X1 U11793 ( .A1(n9203), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9131) );
  NAND2_X1 U11794 ( .A1(n9311), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9130) );
  NAND2_X1 U11795 ( .A1(n8947), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9129) );
  NAND4_X1 U11796 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n15030) );
  NAND2_X1 U11797 ( .A1(n8854), .A2(n15030), .ZN(n9133) );
  NAND2_X1 U11798 ( .A1(n9134), .A2(n9133), .ZN(n9135) );
  XNOR2_X1 U11799 ( .A(n9135), .B(n9321), .ZN(n14536) );
  NOR2_X1 U11800 ( .A1(n9136), .A2(n14541), .ZN(n9137) );
  AOI21_X1 U11801 ( .B1(n15171), .B2(n8854), .A(n9137), .ZN(n14534) );
  NAND2_X1 U11802 ( .A1(n10557), .A2(n8868), .ZN(n9145) );
  INV_X1 U11803 ( .A(n9138), .ZN(n9140) );
  INV_X1 U11804 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U11805 ( .A1(n9140), .A2(n9139), .ZN(n9142) );
  NAND2_X1 U11806 ( .A1(n9142), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9141) );
  MUX2_X1 U11807 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9141), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9143) );
  AOI22_X1 U11808 ( .A1(n11802), .A2(n9176), .B1(n9175), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U11809 ( .A1(n15166), .A2(n9323), .ZN(n9152) );
  NAND2_X1 U11810 ( .A1(n9147), .A2(n9146), .ZN(n9148) );
  NAND2_X1 U11811 ( .A1(n9166), .A2(n9148), .ZN(n15036) );
  AOI22_X1 U11812 ( .A1(n9203), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9311), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U11813 ( .A1(n8947), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9149) );
  OAI211_X1 U11814 ( .C1(n15036), .C2(n9273), .A(n9150), .B(n9149), .ZN(n15016) );
  NAND2_X1 U11815 ( .A1(n8854), .A2(n15016), .ZN(n9151) );
  NAND2_X1 U11816 ( .A1(n9152), .A2(n9151), .ZN(n9153) );
  XNOR2_X1 U11817 ( .A(n9153), .B(n10580), .ZN(n14533) );
  NAND2_X1 U11818 ( .A1(n15166), .A2(n8854), .ZN(n9155) );
  NAND2_X1 U11819 ( .A1(n9318), .A2(n15016), .ZN(n9154) );
  NAND2_X1 U11820 ( .A1(n9155), .A2(n9154), .ZN(n14532) );
  NAND2_X1 U11821 ( .A1(n14533), .A2(n14532), .ZN(n9158) );
  INV_X1 U11822 ( .A(n9156), .ZN(n9157) );
  NAND3_X1 U11823 ( .A1(n14536), .A2(n14534), .A3(n9158), .ZN(n9161) );
  INV_X1 U11824 ( .A(n14533), .ZN(n9160) );
  INV_X1 U11825 ( .A(n14532), .ZN(n9159) );
  NAND2_X1 U11826 ( .A1(n9160), .A2(n9159), .ZN(n14546) );
  NAND2_X1 U11827 ( .A1(n10686), .A2(n8868), .ZN(n9164) );
  NAND2_X1 U11828 ( .A1(n9173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9162) );
  XNOR2_X1 U11829 ( .A(n9162), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14781) );
  AOI22_X1 U11830 ( .A1(n14781), .A2(n9176), .B1(n9175), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n9163) );
  INV_X1 U11831 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11801) );
  INV_X1 U11832 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9165) );
  NAND2_X1 U11833 ( .A1(n9166), .A2(n9165), .ZN(n9167) );
  NAND2_X1 U11834 ( .A1(n9179), .A2(n9167), .ZN(n15019) );
  OR2_X1 U11835 ( .A1(n15019), .A2(n9273), .ZN(n9169) );
  AOI22_X1 U11836 ( .A1(n9203), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9311), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n9168) );
  OAI211_X1 U11837 ( .C1(n8812), .C2(n11801), .A(n9169), .B(n9168), .ZN(n15032) );
  AOI22_X1 U11838 ( .A1(n15161), .A2(n8854), .B1(n9318), .B2(n15032), .ZN(
        n9172) );
  AOI22_X1 U11839 ( .A1(n15161), .A2(n9323), .B1(n8854), .B2(n15032), .ZN(
        n9170) );
  XNOR2_X1 U11840 ( .A(n9170), .B(n10580), .ZN(n9171) );
  XOR2_X1 U11841 ( .A(n9172), .B(n9171), .Z(n14547) );
  NAND2_X1 U11842 ( .A1(n10993), .A2(n8868), .ZN(n9178) );
  OAI21_X1 U11843 ( .B1(n9173), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9174) );
  XNOR2_X1 U11844 ( .A(n9174), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14798) );
  AOI22_X1 U11845 ( .A1(n14798), .A2(n9176), .B1(n9175), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U11846 ( .A1(n15156), .A2(n9323), .ZN(n9186) );
  XNOR2_X1 U11847 ( .A(n9179), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n15000) );
  NAND2_X1 U11848 ( .A1(n15000), .A2(n9310), .ZN(n9184) );
  INV_X1 U11849 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n15723) );
  NAND2_X1 U11850 ( .A1(n9203), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9181) );
  NAND2_X1 U11851 ( .A1(n8947), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9180) );
  OAI211_X1 U11852 ( .C1(n8931), .C2(n15723), .A(n9181), .B(n9180), .ZN(n9182)
         );
  INV_X1 U11853 ( .A(n9182), .ZN(n9183) );
  NAND2_X1 U11854 ( .A1(n9184), .A2(n9183), .ZN(n15015) );
  NAND2_X1 U11855 ( .A1(n15015), .A2(n8854), .ZN(n9185) );
  NAND2_X1 U11856 ( .A1(n9186), .A2(n9185), .ZN(n9187) );
  XNOR2_X1 U11857 ( .A(n9187), .B(n10580), .ZN(n9188) );
  AOI22_X1 U11858 ( .A1(n15156), .A2(n8854), .B1(n9318), .B2(n15015), .ZN(
        n9190) );
  XNOR2_X1 U11859 ( .A(n9188), .B(n9190), .ZN(n14599) );
  INV_X1 U11860 ( .A(n9188), .ZN(n9189) );
  XOR2_X1 U11861 ( .A(n9192), .B(n9191), .Z(n14508) );
  XOR2_X1 U11862 ( .A(n9194), .B(n9193), .Z(n14577) );
  NAND2_X1 U11863 ( .A1(n11287), .A2(n8868), .ZN(n9198) );
  INV_X1 U11864 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11291) );
  OR2_X1 U11865 ( .A1(n8872), .A2(n11291), .ZN(n9197) );
  INV_X1 U11866 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U11867 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  NAND2_X1 U11868 ( .A1(n9202), .A2(n9201), .ZN(n14952) );
  OR2_X1 U11869 ( .A1(n14952), .A2(n9273), .ZN(n9208) );
  INV_X1 U11870 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15718) );
  NAND2_X1 U11871 ( .A1(n9203), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11872 ( .A1(n8947), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9204) );
  OAI211_X1 U11873 ( .C1(n8931), .C2(n15718), .A(n9205), .B(n9204), .ZN(n9206)
         );
  INV_X1 U11874 ( .A(n9206), .ZN(n9207) );
  AOI22_X1 U11875 ( .A1(n14955), .A2(n8854), .B1(n9318), .B2(n14964), .ZN(
        n9211) );
  AOI22_X1 U11876 ( .A1(n14955), .A2(n9323), .B1(n8854), .B2(n14964), .ZN(
        n9209) );
  XNOR2_X1 U11877 ( .A(n9209), .B(n10580), .ZN(n9210) );
  XOR2_X1 U11878 ( .A(n9211), .B(n9210), .Z(n14517) );
  XOR2_X1 U11879 ( .A(n9214), .B(n9213), .Z(n14588) );
  NAND2_X1 U11880 ( .A1(n11494), .A2(n8868), .ZN(n9216) );
  INV_X1 U11881 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11496) );
  OR2_X1 U11882 ( .A1(n8872), .A2(n11496), .ZN(n9215) );
  NAND2_X1 U11883 ( .A1(n15121), .A2(n9323), .ZN(n9226) );
  NAND2_X1 U11884 ( .A1(n9217), .A2(n14501), .ZN(n9218) );
  AND2_X1 U11885 ( .A1(n9233), .A2(n9218), .ZN(n14914) );
  NAND2_X1 U11886 ( .A1(n14914), .A2(n9310), .ZN(n9224) );
  INV_X1 U11887 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11888 ( .A1(n8947), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11889 ( .A1(n9311), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9219) );
  OAI211_X1 U11890 ( .C1(n12714), .C2(n9221), .A(n9220), .B(n9219), .ZN(n9222)
         );
  INV_X1 U11891 ( .A(n9222), .ZN(n9223) );
  NAND2_X1 U11892 ( .A1(n14930), .A2(n8854), .ZN(n9225) );
  NAND2_X1 U11893 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  XNOR2_X1 U11894 ( .A(n9227), .B(n10580), .ZN(n9228) );
  AOI22_X1 U11895 ( .A1(n15121), .A2(n8854), .B1(n9318), .B2(n14930), .ZN(
        n9229) );
  XNOR2_X1 U11896 ( .A(n9228), .B(n9229), .ZN(n14500) );
  INV_X1 U11897 ( .A(n9228), .ZN(n9230) );
  NAND2_X1 U11898 ( .A1(n11611), .A2(n8868), .ZN(n9232) );
  OR2_X1 U11899 ( .A1(n8872), .A2(n7719), .ZN(n9231) );
  INV_X1 U11900 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14561) );
  NAND2_X1 U11901 ( .A1(n9233), .A2(n14561), .ZN(n9234) );
  NAND2_X1 U11902 ( .A1(n9248), .A2(n9234), .ZN(n14894) );
  INV_X1 U11903 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14895) );
  NAND2_X1 U11904 ( .A1(n8947), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U11905 ( .A1(n9311), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9235) );
  OAI211_X1 U11906 ( .C1(n12714), .C2(n14895), .A(n9236), .B(n9235), .ZN(n9237) );
  INV_X1 U11907 ( .A(n9237), .ZN(n9238) );
  AOI22_X1 U11908 ( .A1(n15111), .A2(n8854), .B1(n9318), .B2(n14907), .ZN(
        n9243) );
  NAND2_X1 U11909 ( .A1(n15111), .A2(n9323), .ZN(n9241) );
  NAND2_X1 U11910 ( .A1(n14907), .A2(n8854), .ZN(n9240) );
  NAND2_X1 U11911 ( .A1(n9241), .A2(n9240), .ZN(n9242) );
  XNOR2_X1 U11912 ( .A(n9242), .B(n10580), .ZN(n9245) );
  XOR2_X1 U11913 ( .A(n9243), .B(n9245), .Z(n14560) );
  INV_X1 U11914 ( .A(n9243), .ZN(n9244) );
  NAND2_X1 U11915 ( .A1(n11769), .A2(n8868), .ZN(n9247) );
  OR2_X1 U11916 ( .A1(n8872), .A2(n11774), .ZN(n9246) );
  NAND2_X1 U11917 ( .A1(n14879), .A2(n9323), .ZN(n9257) );
  INV_X1 U11918 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14525) );
  NAND2_X1 U11919 ( .A1(n9248), .A2(n14525), .ZN(n9249) );
  NAND2_X1 U11920 ( .A1(n9250), .A2(n9249), .ZN(n14874) );
  INV_X1 U11921 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14873) );
  NAND2_X1 U11922 ( .A1(n9311), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11923 ( .A1(n8947), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9251) );
  OAI211_X1 U11924 ( .C1(n14873), .C2(n12714), .A(n9252), .B(n9251), .ZN(n9253) );
  INV_X1 U11925 ( .A(n9253), .ZN(n9254) );
  NAND2_X1 U11926 ( .A1(n14887), .A2(n8854), .ZN(n9256) );
  NAND2_X1 U11927 ( .A1(n9257), .A2(n9256), .ZN(n9258) );
  XNOR2_X1 U11928 ( .A(n9258), .B(n10580), .ZN(n9259) );
  AOI22_X1 U11929 ( .A1(n14879), .A2(n8854), .B1(n9318), .B2(n14887), .ZN(
        n9260) );
  XNOR2_X1 U11930 ( .A(n9259), .B(n9260), .ZN(n14524) );
  INV_X1 U11931 ( .A(n9259), .ZN(n9261) );
  NAND2_X1 U11932 ( .A1(n9261), .A2(n9260), .ZN(n9262) );
  XNOR2_X1 U11933 ( .A(n9266), .B(n9263), .ZN(n14607) );
  NAND2_X1 U11934 ( .A1(n14606), .A2(n14607), .ZN(n9264) );
  NAND2_X1 U11935 ( .A1(n12316), .A2(n8868), .ZN(n9268) );
  OR2_X1 U11936 ( .A1(n8872), .A2(n15229), .ZN(n9267) );
  NAND2_X1 U11937 ( .A1(n15093), .A2(n9323), .ZN(n9280) );
  INV_X1 U11938 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U11939 ( .A1(n9271), .A2(n9270), .ZN(n9272) );
  NAND2_X1 U11940 ( .A1(n12973), .A2(n9272), .ZN(n14844) );
  INV_X1 U11941 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14843) );
  NAND2_X1 U11942 ( .A1(n8947), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U11943 ( .A1(n9311), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9274) );
  OAI211_X1 U11944 ( .C1(n12714), .C2(n14843), .A(n9275), .B(n9274), .ZN(n9276) );
  INV_X1 U11945 ( .A(n9276), .ZN(n9277) );
  NAND2_X1 U11946 ( .A1(n14856), .A2(n8854), .ZN(n9279) );
  NAND2_X1 U11947 ( .A1(n9280), .A2(n9279), .ZN(n9281) );
  XNOR2_X1 U11948 ( .A(n9281), .B(n9321), .ZN(n9327) );
  AND2_X1 U11949 ( .A1(n14856), .A2(n9318), .ZN(n9282) );
  AOI21_X1 U11950 ( .B1(n15093), .B2(n8854), .A(n9282), .ZN(n9326) );
  XNOR2_X1 U11951 ( .A(n9327), .B(n9326), .ZN(n14482) );
  INV_X1 U11952 ( .A(n14482), .ZN(n9283) );
  NAND2_X1 U11953 ( .A1(n11772), .A2(P1_B_REG_SCAN_IN), .ZN(n9286) );
  MUX2_X1 U11954 ( .A(P1_B_REG_SCAN_IN), .B(n9286), .S(n11612), .Z(n9287) );
  INV_X1 U11955 ( .A(n9288), .ZN(n15234) );
  NAND2_X1 U11956 ( .A1(n15234), .A2(n11772), .ZN(n10555) );
  INV_X1 U11957 ( .A(n10574), .ZN(n11663) );
  NOR4_X1 U11958 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9292) );
  NOR4_X1 U11959 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9291) );
  NOR4_X1 U11960 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9290) );
  NOR4_X1 U11961 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9289) );
  AND4_X1 U11962 ( .A1(n9292), .A2(n9291), .A3(n9290), .A4(n9289), .ZN(n9298)
         );
  INV_X1 U11963 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15964) );
  INV_X1 U11964 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15760) );
  NAND2_X1 U11965 ( .A1(n15964), .A2(n15760), .ZN(n15710) );
  INV_X1 U11966 ( .A(n15710), .ZN(n9296) );
  NOR4_X1 U11967 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n9295) );
  NOR4_X1 U11968 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9294) );
  NOR4_X1 U11969 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9293) );
  AND4_X1 U11970 ( .A1(n9296), .A2(n9295), .A3(n9294), .A4(n9293), .ZN(n9297)
         );
  NAND2_X1 U11971 ( .A1(n9298), .A2(n9297), .ZN(n10570) );
  INV_X1 U11972 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n15985) );
  NOR2_X1 U11973 ( .A1(n10570), .A2(n15985), .ZN(n9299) );
  NAND2_X1 U11974 ( .A1(n15234), .A2(n11612), .ZN(n10568) );
  OAI21_X1 U11975 ( .B1(n10569), .B2(n9299), .A(n10568), .ZN(n9334) );
  INV_X1 U11976 ( .A(n9334), .ZN(n9307) );
  INV_X1 U11977 ( .A(n9300), .ZN(n9301) );
  NAND2_X1 U11978 ( .A1(n9301), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9303) );
  INV_X1 U11979 ( .A(n11667), .ZN(n10467) );
  NAND2_X1 U11980 ( .A1(n12556), .A2(n12558), .ZN(n9331) );
  INV_X1 U11981 ( .A(n12721), .ZN(n9304) );
  NAND2_X1 U11982 ( .A1(n15471), .A2(n9304), .ZN(n9305) );
  NOR2_X1 U11983 ( .A1(n10467), .A2(n9305), .ZN(n9306) );
  NAND2_X1 U11984 ( .A1(n12318), .A2(n8868), .ZN(n9309) );
  OR2_X1 U11985 ( .A1(n8872), .A2(n12319), .ZN(n9308) );
  NAND2_X2 U11986 ( .A1(n9309), .A2(n9308), .ZN(n15087) );
  NAND2_X1 U11987 ( .A1(n15087), .A2(n8854), .ZN(n9320) );
  XNOR2_X1 U11988 ( .A(n12973), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n12934) );
  NAND2_X1 U11989 ( .A1(n12934), .A2(n9310), .ZN(n9317) );
  INV_X1 U11990 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U11991 ( .A1(n8947), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U11992 ( .A1(n9311), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9312) );
  OAI211_X1 U11993 ( .C1(n12714), .C2(n9314), .A(n9313), .B(n9312), .ZN(n9315)
         );
  INV_X1 U11994 ( .A(n9315), .ZN(n9316) );
  NAND2_X1 U11995 ( .A1(n14837), .A2(n9318), .ZN(n9319) );
  NAND2_X1 U11996 ( .A1(n9320), .A2(n9319), .ZN(n9322) );
  XNOR2_X1 U11997 ( .A(n9322), .B(n9321), .ZN(n9325) );
  AOI22_X1 U11998 ( .A1(n15087), .A2(n9323), .B1(n8854), .B2(n14837), .ZN(
        n9324) );
  XNOR2_X1 U11999 ( .A(n9325), .B(n9324), .ZN(n9348) );
  NAND2_X1 U12000 ( .A1(n9327), .A2(n9326), .ZN(n9347) );
  NAND4_X1 U12001 ( .A1(n9328), .A2(n14621), .A3(n9348), .A4(n9347), .ZN(n9352) );
  INV_X1 U12002 ( .A(n9348), .ZN(n9329) );
  OR2_X1 U12003 ( .A1(n10574), .A2(n9334), .ZN(n9330) );
  NAND2_X1 U12004 ( .A1(n9330), .A2(n11665), .ZN(n11002) );
  NAND2_X1 U12005 ( .A1(n11002), .A2(n11667), .ZN(n11923) );
  NAND2_X1 U12006 ( .A1(n12721), .A2(n9331), .ZN(n9332) );
  AND2_X1 U12007 ( .A1(n9332), .A2(n10468), .ZN(n9333) );
  NAND2_X1 U12008 ( .A1(n9343), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10567) );
  INV_X1 U12009 ( .A(n9335), .ZN(n14664) );
  AND2_X2 U12010 ( .A1(n12721), .A2(n14664), .ZN(n15029) );
  NAND2_X1 U12011 ( .A1(n9310), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9336) );
  INV_X1 U12012 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U12013 ( .A1(n8947), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9338) );
  INV_X1 U12014 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n15830) );
  OR2_X1 U12015 ( .A1(n8931), .A2(n15830), .ZN(n9337) );
  OAI211_X1 U12016 ( .C1(n12714), .C2(n9339), .A(n9338), .B(n9337), .ZN(n9340)
         );
  INV_X1 U12017 ( .A(n9340), .ZN(n9341) );
  AOI22_X1 U12018 ( .A1(n14635), .A2(n14591), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(n6537), .ZN(n9346) );
  NAND2_X1 U12019 ( .A1(n11002), .A2(n9343), .ZN(n9344) );
  NAND2_X1 U12020 ( .A1(n12934), .A2(n14630), .ZN(n9345) );
  OAI211_X1 U12021 ( .C1(n14614), .C2(n14609), .A(n9346), .B(n9345), .ZN(n9350) );
  NOR3_X1 U12022 ( .A1(n9348), .A2(n14619), .A3(n9347), .ZN(n9349) );
  AOI211_X1 U12023 ( .C1(n14617), .C2(n15087), .A(n9350), .B(n9349), .ZN(n9351) );
  NOR2_X1 U12024 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n9354) );
  NAND4_X1 U12025 ( .A1(n9354), .A2(n9353), .A3(n15697), .A4(n9391), .ZN(n9485) );
  INV_X1 U12026 ( .A(n9492), .ZN(n9357) );
  NOR2_X1 U12027 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), 
        .ZN(n9360) );
  NOR2_X1 U12028 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), 
        .ZN(n9359) );
  NOR2_X1 U12029 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n9358) );
  NAND3_X1 U12030 ( .A1(n9443), .A2(n9446), .A3(n9379), .ZN(n9489) );
  INV_X1 U12031 ( .A(n9489), .ZN(n9363) );
  NAND2_X1 U12032 ( .A1(n9382), .A2(n9361), .ZN(n9484) );
  INV_X1 U12033 ( .A(n9484), .ZN(n9362) );
  NAND3_X1 U12034 ( .A1(n9372), .A2(n9365), .A3(n9375), .ZN(n9491) );
  INV_X1 U12035 ( .A(n9491), .ZN(n9366) );
  NAND2_X1 U12036 ( .A1(n9387), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9373) );
  INV_X1 U12037 ( .A(n9621), .ZN(n9377) );
  NAND2_X1 U12038 ( .A1(n9374), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9376) );
  INV_X1 U12039 ( .A(n13559), .ZN(n10047) );
  NAND2_X1 U12040 ( .A1(n10046), .A2(n9378), .ZN(n10082) );
  INV_X1 U12041 ( .A(n10082), .ZN(n9388) );
  NOR2_X1 U12042 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), 
        .ZN(n9381) );
  INV_X1 U12043 ( .A(n9494), .ZN(n9384) );
  OAI21_X1 U12044 ( .B1(n9461), .B2(n9384), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9385) );
  MUX2_X1 U12045 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9385), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n9386) );
  AND2_X2 U12046 ( .A1(n9388), .A2(n10395), .ZN(P3_U3897) );
  INV_X1 U12047 ( .A(n9415), .ZN(n9392) );
  NAND2_X1 U12048 ( .A1(n9392), .A2(n9391), .ZN(n9419) );
  INV_X1 U12049 ( .A(n9426), .ZN(n9394) );
  INV_X1 U12050 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9393) );
  NAND2_X1 U12051 ( .A1(n9394), .A2(n9393), .ZN(n9431) );
  NAND2_X1 U12052 ( .A1(n9431), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9395) );
  INV_X1 U12053 ( .A(n10367), .ZN(n11480) );
  INV_X1 U12054 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n15928) );
  NAND2_X1 U12055 ( .A1(n9415), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9396) );
  INV_X1 U12056 ( .A(n9671), .ZN(n13143) );
  NAND2_X1 U12057 ( .A1(n9399), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9397) );
  INV_X1 U12058 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9400) );
  NAND2_X1 U12059 ( .A1(n9487), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9401) );
  INV_X1 U12060 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15687) );
  NOR2_X1 U12061 ( .A1(n10834), .A2(n15687), .ZN(n10833) );
  INV_X1 U12062 ( .A(n9401), .ZN(n9402) );
  NOR2_X1 U12063 ( .A1(n10833), .A2(n9402), .ZN(n10869) );
  NAND2_X1 U12064 ( .A1(n9403), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9404) );
  MUX2_X1 U12065 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9404), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n9405) );
  INV_X1 U12066 ( .A(n10337), .ZN(n13122) );
  INV_X1 U12067 ( .A(n9406), .ZN(n10965) );
  NAND2_X1 U12068 ( .A1(n9407), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9409) );
  XNOR2_X1 U12069 ( .A(n10329), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n10966) );
  NAND2_X1 U12070 ( .A1(n9413), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9414) );
  MUX2_X1 U12071 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9414), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n9416) );
  NAND2_X1 U12072 ( .A1(n9416), .A2(n9415), .ZN(n10849) );
  NOR2_X1 U12073 ( .A1(n9417), .A2(n9535), .ZN(n9418) );
  AOI21_X1 U12074 ( .B1(n9417), .B2(n9535), .A(n9418), .ZN(n10845) );
  INV_X1 U12075 ( .A(n9418), .ZN(n13138) );
  INV_X1 U12076 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11162) );
  XNOR2_X1 U12077 ( .A(n9671), .B(n11162), .ZN(n13139) );
  NAND2_X1 U12078 ( .A1(n9419), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9421) );
  INV_X1 U12079 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9420) );
  XNOR2_X1 U12080 ( .A(n9421), .B(n9420), .ZN(n10786) );
  NAND2_X1 U12081 ( .A1(n9423), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9424) );
  XNOR2_X1 U12082 ( .A(n10924), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n10915) );
  NAND2_X1 U12083 ( .A1(n10362), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U12084 ( .A1(n9426), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9427) );
  MUX2_X1 U12085 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9427), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n9428) );
  NAND2_X1 U12086 ( .A1(n9428), .A2(n9431), .ZN(n10358) );
  INV_X1 U12087 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11300) );
  NAND2_X1 U12088 ( .A1(n11470), .A2(n11465), .ZN(n9430) );
  XNOR2_X1 U12089 ( .A(n10367), .B(n15928), .ZN(n11466) );
  OAI21_X1 U12090 ( .B1(n9431), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9433) );
  INV_X1 U12091 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9432) );
  INV_X1 U12092 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n13161) );
  NAND2_X1 U12093 ( .A1(n9434), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9435) );
  XNOR2_X1 U12094 ( .A(n9435), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13187) );
  INV_X1 U12095 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11499) );
  NOR2_X1 U12096 ( .A1(n13187), .A2(n11499), .ZN(n9436) );
  AOI21_X1 U12097 ( .B1(n13187), .B2(n11499), .A(n9436), .ZN(n13190) );
  INV_X1 U12098 ( .A(n9436), .ZN(n9437) );
  INV_X1 U12099 ( .A(n9438), .ZN(n9439) );
  NAND2_X1 U12100 ( .A1(n9439), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9440) );
  XNOR2_X1 U12101 ( .A(n9440), .B(P3_IR_REG_13__SCAN_IN), .ZN(n13207) );
  NAND2_X1 U12102 ( .A1(n9441), .A2(n10482), .ZN(n10282) );
  NAND2_X1 U12103 ( .A1(n9438), .A2(n9443), .ZN(n9445) );
  NAND2_X1 U12104 ( .A1(n9445), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9444) );
  MUX2_X1 U12105 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9444), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n9448) );
  INV_X1 U12106 ( .A(n9445), .ZN(n9447) );
  NAND2_X1 U12107 ( .A1(n9447), .A2(n9446), .ZN(n9451) );
  NAND2_X1 U12108 ( .A1(n9448), .A2(n9451), .ZN(n10518) );
  INV_X1 U12109 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12144) );
  XNOR2_X1 U12110 ( .A(n10518), .B(n12144), .ZN(n9567) );
  NAND2_X1 U12111 ( .A1(n10518), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9449) );
  NAND2_X1 U12112 ( .A1(n9451), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9450) );
  MUX2_X1 U12113 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9450), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n9452) );
  NAND2_X1 U12114 ( .A1(n13214), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9455) );
  INV_X1 U12115 ( .A(n9876), .ZN(n13221) );
  NAND2_X1 U12116 ( .A1(n9453), .A2(n13221), .ZN(n9454) );
  NAND2_X1 U12117 ( .A1(n9455), .A2(n9454), .ZN(n13227) );
  NAND2_X1 U12118 ( .A1(n9456), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9457) );
  XNOR2_X1 U12119 ( .A(n9457), .B(P3_IR_REG_16__SCAN_IN), .ZN(n9892) );
  XNOR2_X1 U12120 ( .A(n9892), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13228) );
  NAND2_X1 U12121 ( .A1(n13227), .A2(n13228), .ZN(n13226) );
  INV_X1 U12122 ( .A(n9892), .ZN(n13237) );
  NAND2_X1 U12123 ( .A1(n13237), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9458) );
  NAND2_X1 U12124 ( .A1(n13226), .A2(n9458), .ZN(n9460) );
  NAND2_X1 U12125 ( .A1(n9461), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9459) );
  XNOR2_X1 U12126 ( .A(n9459), .B(P3_IR_REG_17__SCAN_IN), .ZN(n10551) );
  INV_X1 U12127 ( .A(n10551), .ZN(n13260) );
  INV_X1 U12128 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U12129 ( .A1(n9467), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9464) );
  XNOR2_X1 U12130 ( .A(n9464), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13280) );
  INV_X1 U12131 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13436) );
  OR2_X1 U12132 ( .A1(n13280), .A2(n13436), .ZN(n9466) );
  NAND2_X1 U12133 ( .A1(n13280), .A2(n13436), .ZN(n9465) );
  NAND2_X1 U12134 ( .A1(n9466), .A2(n9465), .ZN(n13267) );
  NAND2_X1 U12135 ( .A1(n6654), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9468) );
  XNOR2_X1 U12136 ( .A(n12526), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n9574) );
  XNOR2_X1 U12137 ( .A(n9469), .B(n9574), .ZN(n9587) );
  INV_X1 U12138 ( .A(n9471), .ZN(n9628) );
  AND2_X2 U12139 ( .A1(n12367), .A2(n9625), .ZN(n9474) );
  NAND2_X1 U12140 ( .A1(n9474), .A2(n10081), .ZN(n9481) );
  NAND2_X1 U12141 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), 
        .ZN(n9475) );
  NOR2_X1 U12142 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), 
        .ZN(n9477) );
  OAI21_X1 U12143 ( .B1(n9478), .B2(n9370), .A(n9477), .ZN(n9479) );
  INV_X1 U12144 ( .A(n10242), .ZN(n10070) );
  NOR2_X1 U12145 ( .A1(n10081), .A2(P3_U3151), .ZN(n12530) );
  INV_X1 U12146 ( .A(n12530), .ZN(n12535) );
  NAND2_X1 U12147 ( .A1(n10070), .A2(n12535), .ZN(n9580) );
  INV_X1 U12148 ( .A(n9580), .ZN(n9482) );
  INV_X1 U12149 ( .A(n9516), .ZN(n9577) );
  NOR2_X1 U12150 ( .A1(n9485), .A2(n9484), .ZN(n9496) );
  NAND2_X1 U12151 ( .A1(n9488), .A2(n9487), .ZN(n9490) );
  NOR2_X1 U12152 ( .A1(n9492), .A2(n9491), .ZN(n9493) );
  NAND4_X1 U12153 ( .A1(n9495), .A2(n9496), .A3(n9494), .A4(n9493), .ZN(n9650)
         );
  NAND2_X1 U12154 ( .A1(n9654), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9497) );
  XNOR2_X1 U12155 ( .A(n9497), .B(P3_IR_REG_28__SCAN_IN), .ZN(n10198) );
  NAND2_X1 U12156 ( .A1(n9573), .A2(n10198), .ZN(n10069) );
  INV_X1 U12157 ( .A(n10069), .ZN(n9498) );
  INV_X1 U12158 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12221) );
  INV_X1 U12159 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12147) );
  INV_X1 U12160 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11487) );
  INV_X1 U12161 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11367) );
  NAND2_X1 U12162 ( .A1(n9400), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11172) );
  NOR2_X1 U12163 ( .A1(n11172), .A2(P3_IR_REG_1__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U12164 ( .A1(n10828), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10827) );
  INV_X1 U12165 ( .A(n9499), .ZN(n9500) );
  NAND2_X1 U12166 ( .A1(n10827), .A2(n9500), .ZN(n10880) );
  INV_X1 U12167 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n11046) );
  XNOR2_X1 U12168 ( .A(n10326), .B(n11046), .ZN(n10881) );
  NAND2_X1 U12169 ( .A1(n10880), .A2(n10881), .ZN(n10879) );
  NAND2_X1 U12170 ( .A1(n10326), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U12171 ( .A1(n10879), .A2(n9501), .ZN(n9502) );
  OR2_X1 U12172 ( .A1(n9502), .A2(n10337), .ZN(n9503) );
  NAND2_X1 U12173 ( .A1(n9502), .A2(n10337), .ZN(n10970) );
  XNOR2_X1 U12174 ( .A(n10329), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n10971) );
  INV_X1 U12175 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9539) );
  XNOR2_X1 U12176 ( .A(n9671), .B(n9539), .ZN(n13152) );
  AOI21_X1 U12177 ( .B1(n9506), .B2(n9544), .A(n9507), .ZN(n10784) );
  NAND2_X1 U12178 ( .A1(n10784), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n10920) );
  INV_X1 U12179 ( .A(n9507), .ZN(n10918) );
  INV_X1 U12180 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11101) );
  XNOR2_X1 U12181 ( .A(n10924), .B(n11101), .ZN(n10919) );
  INV_X1 U12182 ( .A(n10358), .ZN(n11309) );
  XNOR2_X1 U12183 ( .A(n10367), .B(n11367), .ZN(n11481) );
  INV_X1 U12184 ( .A(n9508), .ZN(n9509) );
  INV_X1 U12185 ( .A(n13175), .ZN(n9510) );
  NAND2_X1 U12186 ( .A1(n13169), .A2(n9510), .ZN(n9511) );
  XNOR2_X1 U12187 ( .A(n13187), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n13174) );
  INV_X1 U12188 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15738) );
  NAND2_X1 U12189 ( .A1(n13195), .A2(n10286), .ZN(n9512) );
  XNOR2_X1 U12190 ( .A(n10518), .B(n12147), .ZN(n9566) );
  INV_X1 U12191 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n15927) );
  XNOR2_X1 U12192 ( .A(n9892), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13238) );
  OAI21_X1 U12193 ( .B1(n9513), .B2(n13260), .A(n13282), .ZN(n13254) );
  INV_X1 U12194 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12285) );
  INV_X1 U12195 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n15759) );
  OR2_X1 U12196 ( .A1(n13280), .A2(n15759), .ZN(n9515) );
  NAND2_X1 U12197 ( .A1(n13280), .A2(n15759), .ZN(n9514) );
  NAND2_X1 U12198 ( .A1(n9515), .A2(n9514), .ZN(n13281) );
  XNOR2_X1 U12199 ( .A(n12526), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U12200 ( .A1(n9517), .A2(n13284), .ZN(n9586) );
  MUX2_X1 U12201 ( .A(P3_REG1_REG_17__SCAN_IN), .B(P3_REG2_REG_17__SCAN_IN), 
        .S(n9573), .Z(n9571) );
  MUX2_X1 U12202 ( .A(P3_REG1_REG_14__SCAN_IN), .B(P3_REG2_REG_14__SCAN_IN), 
        .S(n9573), .Z(n9568) );
  MUX2_X1 U12203 ( .A(P3_REG1_REG_13__SCAN_IN), .B(P3_REG2_REG_13__SCAN_IN), 
        .S(n9573), .Z(n9565) );
  INV_X1 U12204 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11361) );
  NAND2_X1 U12205 ( .A1(n9519), .A2(n9518), .ZN(n10872) );
  INV_X1 U12206 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10956) );
  INV_X1 U12207 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11174) );
  INV_X1 U12208 ( .A(n10326), .ZN(n10878) );
  NAND2_X1 U12209 ( .A1(n9522), .A2(n10878), .ZN(n13124) );
  INV_X1 U12210 ( .A(n9522), .ZN(n9523) );
  NAND2_X1 U12211 ( .A1(n9523), .A2(n10326), .ZN(n9524) );
  AND2_X1 U12212 ( .A1(n13124), .A2(n9524), .ZN(n10871) );
  NAND2_X1 U12213 ( .A1(n13123), .A2(n13124), .ZN(n9529) );
  INV_X1 U12214 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11218) );
  INV_X1 U12215 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9525) );
  MUX2_X1 U12216 ( .A(n11218), .B(n9525), .S(n9573), .Z(n9526) );
  NAND2_X1 U12217 ( .A1(n9526), .A2(n13122), .ZN(n10958) );
  INV_X1 U12218 ( .A(n9526), .ZN(n9527) );
  NAND2_X1 U12219 ( .A1(n9527), .A2(n10337), .ZN(n9528) );
  AND2_X1 U12220 ( .A1(n10958), .A2(n9528), .ZN(n13125) );
  NAND2_X1 U12221 ( .A1(n9529), .A2(n13125), .ZN(n13128) );
  NAND2_X1 U12222 ( .A1(n13128), .A2(n10958), .ZN(n9533) );
  INV_X1 U12223 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11244) );
  MUX2_X1 U12224 ( .A(n11244), .B(n9410), .S(n9573), .Z(n9530) );
  NAND2_X1 U12225 ( .A1(n9530), .A2(n9411), .ZN(n10841) );
  INV_X1 U12226 ( .A(n9530), .ZN(n9531) );
  NAND2_X1 U12227 ( .A1(n9531), .A2(n10329), .ZN(n9532) );
  AND2_X1 U12228 ( .A1(n10841), .A2(n9532), .ZN(n10960) );
  INV_X1 U12229 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9534) );
  INV_X1 U12230 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11186) );
  MUX2_X1 U12231 ( .A(n9534), .B(n11186), .S(n9573), .Z(n9536) );
  NAND2_X1 U12232 ( .A1(n9536), .A2(n9535), .ZN(n13146) );
  INV_X1 U12233 ( .A(n9536), .ZN(n9537) );
  NAND2_X1 U12234 ( .A1(n9537), .A2(n10849), .ZN(n9538) );
  AND2_X1 U12235 ( .A1(n13146), .A2(n9538), .ZN(n10842) );
  MUX2_X1 U12236 ( .A(n9539), .B(n11162), .S(n9573), .Z(n9540) );
  NAND2_X1 U12237 ( .A1(n9540), .A2(n9671), .ZN(n10790) );
  INV_X1 U12238 ( .A(n9540), .ZN(n9541) );
  NAND2_X1 U12239 ( .A1(n9541), .A2(n13143), .ZN(n9542) );
  AND2_X1 U12240 ( .A1(n10790), .A2(n9542), .ZN(n13147) );
  NAND2_X1 U12241 ( .A1(n10789), .A2(n10790), .ZN(n9548) );
  INV_X1 U12242 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11215) );
  INV_X1 U12243 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10783) );
  MUX2_X1 U12244 ( .A(n11215), .B(n10783), .S(n9573), .Z(n9545) );
  NAND2_X1 U12245 ( .A1(n9545), .A2(n9544), .ZN(n10909) );
  INV_X1 U12246 ( .A(n9545), .ZN(n9546) );
  NAND2_X1 U12247 ( .A1(n9546), .A2(n10786), .ZN(n9547) );
  AND2_X1 U12248 ( .A1(n10909), .A2(n9547), .ZN(n10791) );
  NAND2_X1 U12249 ( .A1(n10913), .A2(n10909), .ZN(n9552) );
  INV_X1 U12250 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11088) );
  MUX2_X1 U12251 ( .A(n11101), .B(n11088), .S(n9573), .Z(n9549) );
  NAND2_X1 U12252 ( .A1(n9549), .A2(n10924), .ZN(n11304) );
  INV_X1 U12253 ( .A(n9549), .ZN(n9550) );
  NAND2_X1 U12254 ( .A1(n9550), .A2(n10362), .ZN(n9551) );
  AND2_X1 U12255 ( .A1(n11304), .A2(n9551), .ZN(n10911) );
  INV_X1 U12256 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11241) );
  MUX2_X1 U12257 ( .A(n11241), .B(n11300), .S(n9573), .Z(n9553) );
  NAND2_X1 U12258 ( .A1(n11309), .A2(n9553), .ZN(n11474) );
  INV_X1 U12259 ( .A(n9553), .ZN(n9554) );
  NAND2_X1 U12260 ( .A1(n10358), .A2(n9554), .ZN(n9555) );
  NAND2_X1 U12261 ( .A1(n11474), .A2(n9555), .ZN(n11303) );
  INV_X1 U12262 ( .A(n11303), .ZN(n9556) );
  MUX2_X1 U12263 ( .A(P3_REG1_REG_10__SCAN_IN), .B(P3_REG2_REG_10__SCAN_IN), 
        .S(n9573), .Z(n9557) );
  OR2_X1 U12264 ( .A1(n9557), .A2(n10367), .ZN(n9559) );
  NAND2_X1 U12265 ( .A1(n10367), .A2(n9557), .ZN(n9558) );
  NAND2_X1 U12266 ( .A1(n9559), .A2(n9558), .ZN(n11473) );
  INV_X1 U12267 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11371) );
  MUX2_X1 U12268 ( .A(n11371), .B(n13161), .S(n9573), .Z(n9560) );
  XNOR2_X1 U12269 ( .A(n13166), .B(n9560), .ZN(n13162) );
  INV_X1 U12270 ( .A(n9560), .ZN(n9561) );
  OR2_X1 U12271 ( .A1(n13166), .A2(n9561), .ZN(n13181) );
  MUX2_X1 U12272 ( .A(P3_REG1_REG_12__SCAN_IN), .B(P3_REG2_REG_12__SCAN_IN), 
        .S(n9573), .Z(n9563) );
  XNOR2_X1 U12273 ( .A(n9563), .B(n13187), .ZN(n13180) );
  AND2_X1 U12274 ( .A1(n13181), .A2(n13180), .ZN(n9562) );
  XNOR2_X1 U12275 ( .A(n9565), .B(n13207), .ZN(n13199) );
  INV_X1 U12276 ( .A(n13187), .ZN(n10440) );
  NAND2_X1 U12277 ( .A1(n9563), .A2(n10440), .ZN(n13200) );
  AND2_X1 U12278 ( .A1(n13199), .A2(n13200), .ZN(n9564) );
  INV_X1 U12279 ( .A(n9566), .ZN(n10287) );
  INV_X1 U12280 ( .A(n9567), .ZN(n10283) );
  MUX2_X1 U12281 ( .A(n10287), .B(n10283), .S(n9573), .Z(n10291) );
  MUX2_X1 U12282 ( .A(P3_REG1_REG_15__SCAN_IN), .B(P3_REG2_REG_15__SCAN_IN), 
        .S(n9573), .Z(n13216) );
  INV_X1 U12283 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12231) );
  MUX2_X1 U12284 ( .A(n12221), .B(n12231), .S(n9573), .Z(n9570) );
  NAND2_X1 U12285 ( .A1(n9570), .A2(n9892), .ZN(n13231) );
  NOR2_X1 U12286 ( .A1(n9570), .A2(n9892), .ZN(n13230) );
  XOR2_X1 U12287 ( .A(n10551), .B(n9571), .Z(n13257) );
  NOR2_X1 U12288 ( .A1(n13256), .A2(n13257), .ZN(n13255) );
  MUX2_X1 U12289 ( .A(P3_REG1_REG_18__SCAN_IN), .B(P3_REG2_REG_18__SCAN_IN), 
        .S(n9573), .Z(n13276) );
  MUX2_X1 U12290 ( .A(n9575), .B(n9574), .S(n9573), .Z(n9576) );
  INV_X1 U12291 ( .A(n10198), .ZN(n13548) );
  NAND2_X1 U12292 ( .A1(n9577), .A2(n13548), .ZN(n9579) );
  NAND2_X1 U12293 ( .A1(P3_U3897), .A2(n10198), .ZN(n9578) );
  NAND2_X1 U12294 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13011)
         );
  NAND2_X1 U12295 ( .A1(n15694), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n9582) );
  OAI211_X1 U12296 ( .C1(n13261), .C2(n12526), .A(n13011), .B(n9582), .ZN(
        n9583) );
  OAI211_X1 U12297 ( .C1(n9587), .C2(n13288), .A(n9586), .B(n9585), .ZN(
        P3_U3201) );
  INV_X1 U12298 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9617) );
  INV_X1 U12299 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15226) );
  MUX2_X1 U12300 ( .A(n12905), .B(n15226), .S(n10425), .Z(n9595) );
  XNOR2_X1 U12301 ( .A(n9595), .B(SI_29_), .ZN(n9593) );
  NAND2_X1 U12302 ( .A1(n12904), .A2(n8102), .ZN(n9592) );
  OR2_X1 U12303 ( .A1(n9606), .A2(n12905), .ZN(n9591) );
  INV_X1 U12304 ( .A(SI_29_), .ZN(n15965) );
  MUX2_X1 U12305 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n10425), .Z(n9596) );
  NAND2_X1 U12306 ( .A1(n9596), .A2(SI_30_), .ZN(n9602) );
  OAI21_X1 U12307 ( .B1(SI_30_), .B2(n9596), .A(n9602), .ZN(n9597) );
  NAND2_X1 U12308 ( .A1(n9598), .A2(n9597), .ZN(n9599) );
  NAND2_X1 U12309 ( .A1(n12805), .A2(n8102), .ZN(n9601) );
  INV_X1 U12310 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12806) );
  OR2_X1 U12311 ( .A1(n9606), .A2(n12806), .ZN(n9600) );
  NAND2_X1 U12312 ( .A1(n14027), .A2(n14411), .ZN(n14028) );
  MUX2_X1 U12313 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n10425), .Z(n9604) );
  XNOR2_X1 U12314 ( .A(n9604), .B(SI_31_), .ZN(n9605) );
  INV_X1 U12315 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14467) );
  OR2_X1 U12316 ( .A1(n9606), .A2(n14467), .ZN(n9607) );
  XNOR2_X1 U12317 ( .A(n14028), .B(n13872), .ZN(n9608) );
  NOR2_X2 U12318 ( .A1(n9608), .A2(n8582), .ZN(n14023) );
  INV_X1 U12319 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9612) );
  NAND2_X1 U12320 ( .A1(n12833), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U12321 ( .A1(n9609), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9610) );
  OAI211_X1 U12322 ( .C1(n9613), .C2(n9612), .A(n9611), .B(n9610), .ZN(n13959)
         );
  INV_X1 U12323 ( .A(P2_B_REG_SCAN_IN), .ZN(n9614) );
  NOR2_X1 U12324 ( .A1(n13953), .A2(n9614), .ZN(n9615) );
  OR2_X1 U12325 ( .A1(n14118), .A2(n9615), .ZN(n12837) );
  INV_X1 U12326 ( .A(n12837), .ZN(n9616) );
  NOR2_X1 U12327 ( .A1(n14023), .A2(n14318), .ZN(n14314) );
  NAND2_X1 U12328 ( .A1(n13872), .A2(n9618), .ZN(n9619) );
  NAND2_X1 U12329 ( .A1(n9620), .A2(n9619), .ZN(P2_U3498) );
  XNOR2_X1 U12330 ( .A(n9621), .B(P3_B_REG_SCAN_IN), .ZN(n9622) );
  NAND2_X1 U12331 ( .A1(n9622), .A2(n13559), .ZN(n9623) );
  NAND2_X1 U12332 ( .A1(n13555), .A2(n9621), .ZN(n9624) );
  INV_X1 U12333 ( .A(n9625), .ZN(n10042) );
  NAND2_X1 U12334 ( .A1(n9626), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9627) );
  NAND2_X1 U12335 ( .A1(n10043), .A2(n9625), .ZN(n9630) );
  NAND2_X1 U12336 ( .A1(n10547), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9707) );
  INV_X1 U12337 ( .A(n9707), .ZN(n9631) );
  XNOR2_X1 U12338 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9700) );
  NAND2_X1 U12339 ( .A1(n10428), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9632) );
  INV_X1 U12340 ( .A(n9717), .ZN(n9634) );
  NAND2_X1 U12341 ( .A1(n9633), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9635) );
  XNOR2_X1 U12342 ( .A(n10432), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n9727) );
  INV_X1 U12343 ( .A(n9727), .ZN(n9636) );
  NAND2_X1 U12344 ( .A1(n10432), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9637) );
  XNOR2_X1 U12345 ( .A(n10430), .B(P2_DATAO_REG_4__SCAN_IN), .ZN(n9740) );
  INV_X1 U12346 ( .A(n9740), .ZN(n9639) );
  NAND2_X1 U12347 ( .A1(n9741), .A2(n9639), .ZN(n9641) );
  NAND2_X1 U12348 ( .A1(n10430), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12349 ( .A1(n10434), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U12350 ( .A1(n10371), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9644) );
  XNOR2_X1 U12351 ( .A(n9773), .B(n9771), .ZN(n10359) );
  NAND2_X1 U12352 ( .A1(n10359), .A2(n9742), .ZN(n9649) );
  AOI22_X1 U12353 ( .A1(n10924), .A2(n9944), .B1(n9995), .B2(SI_8_), .ZN(n9648) );
  NAND2_X1 U12354 ( .A1(n9649), .A2(n9648), .ZN(n11819) );
  XNOR2_X1 U12355 ( .A(n9722), .B(n11819), .ZN(n9693) );
  INV_X1 U12356 ( .A(n9650), .ZN(n9652) );
  NAND2_X1 U12357 ( .A1(n9652), .A2(n9651), .ZN(n12799) );
  NOR2_X1 U12358 ( .A1(P3_IR_REG_29__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), 
        .ZN(n9655) );
  NAND3_X1 U12359 ( .A1(n9654), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_IR_REG_30__SCAN_IN), .ZN(n9660) );
  INV_X1 U12360 ( .A(n9655), .ZN(n9658) );
  XNOR2_X1 U12361 ( .A(P3_IR_REG_31__SCAN_IN), .B(P3_IR_REG_30__SCAN_IN), .ZN(
        n9656) );
  OAI21_X1 U12362 ( .B1(n9658), .B2(n9657), .A(n9656), .ZN(n9659) );
  NAND2_X1 U12363 ( .A1(n9746), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9670) );
  INV_X2 U12364 ( .A(n10189), .ZN(n12337) );
  NAND2_X1 U12365 ( .A1(n12337), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9669) );
  NAND2_X1 U12366 ( .A1(n9687), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U12367 ( .A1(n9781), .A2(n9666), .ZN(n11820) );
  NAND2_X1 U12368 ( .A1(n9748), .A2(n11820), .ZN(n9668) );
  INV_X4 U12369 ( .A(n9697), .ZN(n12338) );
  NAND2_X1 U12370 ( .A1(n12338), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9667) );
  XNOR2_X1 U12371 ( .A(n9693), .B(n10107), .ZN(n11814) );
  AND2_X1 U12372 ( .A1(n9944), .A2(n9671), .ZN(n9672) );
  AOI21_X1 U12373 ( .B1(n9995), .B2(SI_6_), .A(n9672), .ZN(n9676) );
  XNOR2_X1 U12374 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9673) );
  XNOR2_X1 U12375 ( .A(n9674), .B(n9673), .ZN(n10330) );
  NAND2_X1 U12376 ( .A1(n10330), .A2(n9742), .ZN(n9675) );
  INV_X1 U12377 ( .A(n11169), .ZN(n11656) );
  XNOR2_X1 U12378 ( .A(n9722), .B(n11656), .ZN(n11642) );
  NAND2_X1 U12379 ( .A1(n9762), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9677) );
  NAND2_X1 U12380 ( .A1(n9685), .A2(n9677), .ZN(n11652) );
  NAND2_X1 U12381 ( .A1(n9746), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9678) );
  NAND2_X1 U12382 ( .A1(n11642), .A2(n13111), .ZN(n11643) );
  XNOR2_X1 U12383 ( .A(n9682), .B(n9681), .ZN(n10354) );
  NAND2_X1 U12384 ( .A1(n10354), .A2(n9742), .ZN(n9684) );
  INV_X1 U12385 ( .A(SI_7_), .ZN(n10355) );
  AOI22_X1 U12386 ( .A1(n9995), .A2(n10355), .B1(n10786), .B2(n9944), .ZN(
        n9683) );
  NAND2_X1 U12387 ( .A1(n9684), .A2(n9683), .ZN(n11644) );
  NAND2_X1 U12388 ( .A1(n9746), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9691) );
  NAND2_X1 U12389 ( .A1(n9759), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9690) );
  NAND2_X1 U12390 ( .A1(n9685), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U12391 ( .A1(n9687), .A2(n9686), .ZN(n11648) );
  NAND2_X1 U12392 ( .A1(n12338), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9688) );
  XNOR2_X1 U12393 ( .A(n9722), .B(n12491), .ZN(n11811) );
  OAI21_X1 U12394 ( .B1(n11814), .B2(n11643), .A(n11811), .ZN(n9770) );
  INV_X1 U12395 ( .A(n13110), .ZN(n11817) );
  INV_X1 U12396 ( .A(n11811), .ZN(n9692) );
  OAI21_X1 U12397 ( .B1(n11814), .B2(n11817), .A(n9692), .ZN(n9769) );
  NAND2_X1 U12398 ( .A1(n9759), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9696) );
  NAND2_X1 U12399 ( .A1(n9748), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9695) );
  NAND2_X1 U12400 ( .A1(n9746), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9694) );
  NAND3_X1 U12401 ( .A1(n9696), .A2(n9695), .A3(n9694), .ZN(n9699) );
  NOR2_X2 U12402 ( .A1(n9699), .A2(n9698), .ZN(n10098) );
  XNOR2_X1 U12403 ( .A(n9700), .B(n9707), .ZN(n10353) );
  NAND2_X1 U12404 ( .A1(n12338), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U12405 ( .A1(n9746), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9703) );
  NAND2_X1 U12406 ( .A1(n9759), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9702) );
  NAND2_X1 U12407 ( .A1(n9748), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9701) );
  INV_X1 U12408 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9705) );
  NAND2_X1 U12409 ( .A1(n9705), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U12410 ( .A1(n9707), .A2(n9706), .ZN(n10344) );
  NAND2_X1 U12411 ( .A1(n9944), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9708) );
  OAI211_X1 U12412 ( .C1(n9790), .C2(n10346), .A(n9709), .B(n9708), .ZN(n10930) );
  NAND2_X1 U12413 ( .A1(n12363), .A2(n12365), .ZN(n10216) );
  INV_X1 U12414 ( .A(n10216), .ZN(n9712) );
  XNOR2_X1 U12415 ( .A(n9715), .B(n11357), .ZN(n9710) );
  NOR2_X1 U12416 ( .A1(n9710), .A2(n7138), .ZN(n9713) );
  NOR3_X1 U12417 ( .A1(n9715), .A2(n10098), .A3(n11357), .ZN(n9711) );
  NAND2_X1 U12418 ( .A1(n10930), .A2(n13118), .ZN(n11411) );
  INV_X1 U12419 ( .A(n9713), .ZN(n9714) );
  XNOR2_X1 U12420 ( .A(n9716), .B(n9717), .ZN(n10325) );
  INV_X1 U12421 ( .A(n10325), .ZN(n9718) );
  NAND2_X1 U12422 ( .A1(n9995), .A2(n10324), .ZN(n9720) );
  NAND2_X1 U12423 ( .A1(n9944), .A2(n10326), .ZN(n9719) );
  AND3_X1 U12424 ( .A1(n9721), .A2(n9720), .A3(n9719), .ZN(n11405) );
  XNOR2_X1 U12425 ( .A(n9722), .B(n11405), .ZN(n9737) );
  NAND2_X1 U12426 ( .A1(n12338), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U12427 ( .A1(n9759), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U12428 ( .A1(n9746), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9724) );
  NAND2_X1 U12429 ( .A1(n9748), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9723) );
  XNOR2_X1 U12430 ( .A(n9737), .B(n13115), .ZN(n11401) );
  XNOR2_X1 U12431 ( .A(n9728), .B(n9727), .ZN(n10336) );
  NAND2_X1 U12432 ( .A1(n9742), .A2(n10336), .ZN(n9731) );
  NAND2_X1 U12433 ( .A1(n9995), .A2(n10335), .ZN(n9730) );
  NAND2_X1 U12434 ( .A1(n9944), .A2(n10337), .ZN(n9729) );
  XNOR2_X1 U12435 ( .A(n9722), .B(n11395), .ZN(n9738) );
  NAND2_X1 U12436 ( .A1(n9748), .A2(n9732), .ZN(n9735) );
  NAND2_X1 U12437 ( .A1(n12338), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9734) );
  NAND2_X1 U12438 ( .A1(n9746), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9733) );
  XNOR2_X1 U12439 ( .A(n9738), .B(n13114), .ZN(n11391) );
  NAND2_X1 U12440 ( .A1(n9737), .A2(n11414), .ZN(n11392) );
  NAND3_X1 U12441 ( .A1(n11399), .A2(n11391), .A3(n11392), .ZN(n11390) );
  XNOR2_X1 U12442 ( .A(n9741), .B(n9740), .ZN(n10328) );
  NAND2_X1 U12443 ( .A1(n9742), .A2(n10328), .ZN(n9745) );
  INV_X1 U12444 ( .A(SI_4_), .ZN(n10327) );
  NAND2_X1 U12445 ( .A1(n9995), .A2(n10327), .ZN(n9744) );
  NAND2_X1 U12446 ( .A1(n9944), .A2(n10329), .ZN(n9743) );
  XNOR2_X1 U12447 ( .A(n9715), .B(n11507), .ZN(n9753) );
  NAND2_X1 U12448 ( .A1(n9746), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U12449 ( .A1(n9759), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9751) );
  NAND2_X1 U12450 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9747) );
  NAND2_X1 U12451 ( .A1(n9760), .A2(n9747), .ZN(n11511) );
  NAND2_X1 U12452 ( .A1(n9748), .A2(n11511), .ZN(n9750) );
  NAND2_X1 U12453 ( .A1(n12338), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U12454 ( .A1(n9753), .A2(n11632), .ZN(n9754) );
  OAI21_X1 U12455 ( .B1(n9753), .B2(n11632), .A(n9754), .ZN(n11505) );
  XNOR2_X1 U12456 ( .A(n9756), .B(n7059), .ZN(n10334) );
  NAND2_X1 U12457 ( .A1(n9742), .A2(n10334), .ZN(n9758) );
  NAND2_X1 U12458 ( .A1(n9944), .A2(n10849), .ZN(n9757) );
  OAI211_X1 U12459 ( .C1(n9790), .C2(SI_5_), .A(n9758), .B(n9757), .ZN(n11631)
         );
  INV_X1 U12460 ( .A(n11631), .ZN(n11206) );
  XNOR2_X1 U12461 ( .A(n9715), .B(n11206), .ZN(n9767) );
  NAND2_X1 U12462 ( .A1(n9746), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9766) );
  NAND2_X1 U12463 ( .A1(n9759), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9765) );
  NAND2_X1 U12464 ( .A1(n9760), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U12465 ( .A1(n9762), .A2(n9761), .ZN(n11635) );
  NAND2_X1 U12466 ( .A1(n12338), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9763) );
  XNOR2_X1 U12467 ( .A(n9767), .B(n11657), .ZN(n11629) );
  NAND2_X1 U12468 ( .A1(n9767), .A2(n11657), .ZN(n11639) );
  OAI211_X1 U12469 ( .C1(n11642), .C2(n13111), .A(n11639), .B(n11811), .ZN(
        n9768) );
  INV_X1 U12470 ( .A(n9771), .ZN(n9772) );
  NAND2_X1 U12471 ( .A1(n9773), .A2(n9772), .ZN(n9776) );
  NAND2_X1 U12472 ( .A1(n9774), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U12473 ( .A1(n9776), .A2(n9775), .ZN(n9788) );
  XNOR2_X1 U12474 ( .A(n9788), .B(n9787), .ZN(n10356) );
  NAND2_X1 U12475 ( .A1(n10356), .A2(n9742), .ZN(n9778) );
  INV_X1 U12476 ( .A(SI_9_), .ZN(n10357) );
  AOI22_X1 U12477 ( .A1(n10358), .A2(n9944), .B1(n9995), .B2(n10357), .ZN(
        n9777) );
  NAND2_X1 U12478 ( .A1(n9778), .A2(n9777), .ZN(n11793) );
  XNOR2_X1 U12479 ( .A(n9722), .B(n11793), .ZN(n9800) );
  NAND2_X1 U12480 ( .A1(n9746), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9786) );
  NAND2_X1 U12481 ( .A1(n12337), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9785) );
  NAND2_X1 U12482 ( .A1(n9781), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9782) );
  NAND2_X1 U12483 ( .A1(n9794), .A2(n9782), .ZN(n11790) );
  NAND2_X1 U12484 ( .A1(n9748), .A2(n11790), .ZN(n9784) );
  NAND2_X1 U12485 ( .A1(n12338), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9783) );
  NAND4_X1 U12486 ( .A1(n9786), .A2(n9785), .A3(n9784), .A4(n9783), .ZN(n13108) );
  INV_X1 U12487 ( .A(n13108), .ZN(n11905) );
  XNOR2_X1 U12488 ( .A(n9800), .B(n11905), .ZN(n11785) );
  NAND2_X1 U12489 ( .A1(n10457), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9789) );
  XNOR2_X1 U12490 ( .A(n9811), .B(n9810), .ZN(n10365) );
  NAND2_X1 U12491 ( .A1(n10365), .A2(n9742), .ZN(n9793) );
  NOR2_X1 U12492 ( .A1(n9790), .A2(SI_10_), .ZN(n9791) );
  AOI21_X1 U12493 ( .B1(n10367), .B2(n9944), .A(n9791), .ZN(n9792) );
  NAND2_X1 U12494 ( .A1(n9793), .A2(n9792), .ZN(n11910) );
  XNOR2_X1 U12495 ( .A(n11910), .B(n9722), .ZN(n9802) );
  NAND2_X1 U12496 ( .A1(n9746), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U12497 ( .A1(n12337), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U12498 ( .A1(n9794), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9795) );
  NAND2_X1 U12499 ( .A1(n9804), .A2(n9795), .ZN(n11907) );
  NAND2_X1 U12500 ( .A1(n12338), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9796) );
  NAND4_X1 U12501 ( .A1(n9799), .A2(n9798), .A3(n9797), .A4(n9796), .ZN(n13107) );
  INV_X1 U12502 ( .A(n13107), .ZN(n12242) );
  XNOR2_X1 U12503 ( .A(n9802), .B(n12242), .ZN(n11901) );
  INV_X1 U12504 ( .A(n9800), .ZN(n9801) );
  NAND2_X1 U12505 ( .A1(n9801), .A2(n11905), .ZN(n11898) );
  INV_X1 U12506 ( .A(n9802), .ZN(n9803) );
  NAND2_X1 U12507 ( .A1(n9804), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U12508 ( .A1(n9827), .A2(n9805), .ZN(n12245) );
  NAND2_X1 U12509 ( .A1(n9746), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9808) );
  NAND2_X1 U12510 ( .A1(n12337), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U12511 ( .A1(n12338), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9806) );
  NAND4_X1 U12512 ( .A1(n9809), .A2(n9808), .A3(n9807), .A4(n9806), .ZN(n13106) );
  INV_X1 U12513 ( .A(n13106), .ZN(n12255) );
  NAND2_X1 U12514 ( .A1(n10448), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9812) );
  XNOR2_X1 U12515 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9813) );
  XNOR2_X1 U12516 ( .A(n9816), .B(n9813), .ZN(n10369) );
  NAND2_X1 U12517 ( .A1(n10369), .A2(n9742), .ZN(n9815) );
  AOI22_X1 U12518 ( .A1(n13166), .A2(n9944), .B1(n9995), .B2(n15810), .ZN(
        n9814) );
  NAND2_X1 U12519 ( .A1(n9815), .A2(n9814), .ZN(n12240) );
  XNOR2_X1 U12520 ( .A(n12240), .B(n10026), .ZN(n12235) );
  NAND2_X1 U12521 ( .A1(n10452), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U12522 ( .A1(n10459), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U12523 ( .A1(n10461), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U12524 ( .A1(n9837), .A2(n9819), .ZN(n9821) );
  NAND2_X1 U12525 ( .A1(n9822), .A2(n9821), .ZN(n9823) );
  NAND2_X1 U12526 ( .A1(n9838), .A2(n9823), .ZN(n10439) );
  OR2_X1 U12527 ( .A1(n10439), .A2(n12331), .ZN(n9825) );
  AOI22_X1 U12528 ( .A1(n9995), .A2(SI_12_), .B1(n13187), .B2(n9944), .ZN(
        n9824) );
  XNOR2_X1 U12529 ( .A(n12256), .B(n9715), .ZN(n9832) );
  INV_X1 U12530 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U12531 ( .A1(n9827), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9828) );
  NAND2_X1 U12532 ( .A1(n9847), .A2(n9828), .ZN(n12259) );
  AOI22_X1 U12533 ( .A1(n9746), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n12337), 
        .B2(P3_REG1_REG_12__SCAN_IN), .ZN(n9829) );
  OAI211_X1 U12534 ( .C1(n9697), .C2(n9831), .A(n9830), .B(n9829), .ZN(n13105)
         );
  NAND2_X1 U12535 ( .A1(n9832), .A2(n13105), .ZN(n12249) );
  OAI21_X1 U12536 ( .B1(n12255), .B2(n12235), .A(n12249), .ZN(n9836) );
  NAND3_X1 U12537 ( .A1(n12249), .A2(n12255), .A3(n12235), .ZN(n9834) );
  INV_X1 U12538 ( .A(n9832), .ZN(n9833) );
  INV_X1 U12539 ( .A(n13105), .ZN(n12209) );
  NAND2_X1 U12540 ( .A1(n9833), .A2(n12209), .ZN(n12248) );
  NAND2_X1 U12541 ( .A1(n9859), .A2(n10465), .ZN(n9854) );
  OR2_X1 U12542 ( .A1(n9859), .A2(n10465), .ZN(n9839) );
  NAND2_X1 U12543 ( .A1(n9840), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9855) );
  INV_X1 U12544 ( .A(n9840), .ZN(n9841) );
  NAND2_X1 U12545 ( .A1(n9841), .A2(n10477), .ZN(n9842) );
  NAND2_X1 U12546 ( .A1(n9855), .A2(n9842), .ZN(n10481) );
  OR2_X1 U12547 ( .A1(n10481), .A2(n12331), .ZN(n9844) );
  AOI22_X1 U12548 ( .A1(n9995), .A2(SI_13_), .B1(n13207), .B2(n9944), .ZN(
        n9843) );
  XNOR2_X1 U12549 ( .A(n12420), .B(n9722), .ZN(n9852) );
  NAND2_X1 U12550 ( .A1(n9847), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U12551 ( .A1(n9863), .A2(n9848), .ZN(n12211) );
  AOI22_X1 U12552 ( .A1(n9746), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n12337), 
        .B2(P3_REG1_REG_13__SCAN_IN), .ZN(n9850) );
  NAND2_X1 U12553 ( .A1(n12338), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9849) );
  NOR2_X1 U12554 ( .A1(n9852), .A2(n13104), .ZN(n12204) );
  NAND2_X1 U12555 ( .A1(n10656), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9870) );
  INV_X1 U12556 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10684) );
  NAND2_X1 U12557 ( .A1(n10684), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9853) );
  NAND2_X1 U12558 ( .A1(n9870), .A2(n9853), .ZN(n9857) );
  NAND3_X1 U12559 ( .A1(n9855), .A2(n9857), .A3(n9854), .ZN(n9860) );
  AND2_X1 U12560 ( .A1(n10477), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n9856) );
  NOR2_X1 U12561 ( .A1(n9857), .A2(n9856), .ZN(n9858) );
  NAND2_X1 U12562 ( .A1(n9860), .A2(n9871), .ZN(n10517) );
  NAND2_X1 U12563 ( .A1(n10517), .A2(n9742), .ZN(n9862) );
  AOI22_X1 U12564 ( .A1(n9995), .A2(n15956), .B1(n10518), .B2(n9944), .ZN(
        n9861) );
  NAND2_X1 U12565 ( .A1(n9862), .A2(n9861), .ZN(n12267) );
  XNOR2_X1 U12566 ( .A(n12267), .B(n9722), .ZN(n9867) );
  INV_X1 U12567 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U12568 ( .A1(n9863), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9864) );
  NAND2_X1 U12569 ( .A1(n9895), .A2(n9864), .ZN(n12270) );
  AOI22_X1 U12570 ( .A1(n9746), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n12337), 
        .B2(P3_REG1_REG_14__SCAN_IN), .ZN(n9865) );
  OAI211_X1 U12571 ( .C1(n9697), .C2(n12151), .A(n9866), .B(n9865), .ZN(n12207) );
  XNOR2_X1 U12572 ( .A(n9867), .B(n12207), .ZN(n12262) );
  INV_X1 U12573 ( .A(n9867), .ZN(n9868) );
  INV_X1 U12574 ( .A(n12207), .ZN(n12300) );
  NAND2_X1 U12575 ( .A1(n9868), .A2(n12300), .ZN(n9869) );
  NAND2_X1 U12576 ( .A1(n9871), .A2(n9870), .ZN(n9874) );
  NAND2_X1 U12577 ( .A1(n15737), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9886) );
  NAND2_X1 U12578 ( .A1(n10736), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U12579 ( .A1(n9874), .A2(n9873), .ZN(n9887) );
  OR2_X1 U12580 ( .A1(n9874), .A2(n9873), .ZN(n9875) );
  AND2_X1 U12581 ( .A1(n9887), .A2(n9875), .ZN(n10534) );
  NAND2_X1 U12582 ( .A1(n10534), .A2(n9742), .ZN(n9878) );
  AOI22_X1 U12583 ( .A1(n9876), .A2(n9944), .B1(n9995), .B2(SI_15_), .ZN(n9877) );
  XNOR2_X1 U12584 ( .A(n12302), .B(n10026), .ZN(n12295) );
  XNOR2_X1 U12585 ( .A(n9895), .B(P3_REG3_REG_15__SCAN_IN), .ZN(n12297) );
  INV_X1 U12586 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15758) );
  NAND2_X1 U12587 ( .A1(n12337), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U12588 ( .A1(n12338), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9879) );
  OAI211_X1 U12589 ( .C1(n15758), .C2(n10176), .A(n9880), .B(n9879), .ZN(n9881) );
  INV_X1 U12590 ( .A(n9881), .ZN(n9882) );
  NOR2_X1 U12591 ( .A1(n12295), .A2(n13103), .ZN(n9885) );
  INV_X1 U12592 ( .A(n12295), .ZN(n9884) );
  OAI22_X1 U12593 ( .A1(n12294), .A2(n9885), .B1(n13039), .B2(n9884), .ZN(
        n13037) );
  INV_X1 U12594 ( .A(n13037), .ZN(n9903) );
  NAND2_X1 U12595 ( .A1(n9887), .A2(n9886), .ZN(n9890) );
  NAND2_X1 U12596 ( .A1(n10558), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9906) );
  NAND2_X1 U12597 ( .A1(n10565), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9888) );
  NAND2_X1 U12598 ( .A1(n9890), .A2(n9889), .ZN(n9907) );
  OR2_X1 U12599 ( .A1(n9890), .A2(n9889), .ZN(n9891) );
  AND2_X1 U12600 ( .A1(n9907), .A2(n9891), .ZN(n10548) );
  NAND2_X1 U12601 ( .A1(n10548), .A2(n9742), .ZN(n9894) );
  AOI22_X1 U12602 ( .A1(n9892), .A2(n9944), .B1(SI_16_), .B2(n9995), .ZN(n9893) );
  XNOR2_X1 U12603 ( .A(n13042), .B(n9715), .ZN(n13035) );
  NAND2_X1 U12604 ( .A1(n9896), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U12605 ( .A1(n9916), .A2(n9897), .ZN(n13041) );
  NAND2_X1 U12606 ( .A1(n12337), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9899) );
  NAND2_X1 U12607 ( .A1(n12338), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9898) );
  OAI211_X1 U12608 ( .C1(n12231), .C2(n10176), .A(n9899), .B(n9898), .ZN(n9900) );
  INV_X1 U12609 ( .A(n9900), .ZN(n9901) );
  NAND2_X1 U12610 ( .A1(n13035), .A2(n12275), .ZN(n9904) );
  NAND2_X1 U12611 ( .A1(n10687), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U12612 ( .A1(n10701), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9908) );
  OR2_X1 U12613 ( .A1(n9910), .A2(n9909), .ZN(n9911) );
  NAND2_X1 U12614 ( .A1(n9926), .A2(n9911), .ZN(n10553) );
  OR2_X1 U12615 ( .A1(n10553), .A2(n12331), .ZN(n9913) );
  AOI22_X1 U12616 ( .A1(n9995), .A2(SI_17_), .B1(n10551), .B2(n9944), .ZN(
        n9912) );
  XNOR2_X1 U12617 ( .A(n13051), .B(n9715), .ZN(n13046) );
  INV_X1 U12618 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9914) );
  NAND2_X1 U12619 ( .A1(n9916), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U12620 ( .A1(n9933), .A2(n9917), .ZN(n13054) );
  NAND2_X1 U12621 ( .A1(n12338), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U12622 ( .A1(n12337), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9918) );
  OAI211_X1 U12623 ( .C1(n10176), .C2(n13253), .A(n9919), .B(n9918), .ZN(n9920) );
  INV_X1 U12624 ( .A(n9920), .ZN(n9921) );
  NOR2_X1 U12625 ( .A1(n13046), .A2(n13102), .ZN(n9924) );
  INV_X1 U12626 ( .A(n13046), .ZN(n9923) );
  NAND2_X1 U12627 ( .A1(n9926), .A2(n9925), .ZN(n9929) );
  NAND2_X1 U12628 ( .A1(n10994), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9941) );
  INV_X1 U12629 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10997) );
  NAND2_X1 U12630 ( .A1(n10997), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9927) );
  OR2_X1 U12631 ( .A1(n9929), .A2(n9928), .ZN(n9930) );
  NAND2_X1 U12632 ( .A1(n9942), .A2(n9930), .ZN(n10734) );
  OR2_X1 U12633 ( .A1(n10734), .A2(n12331), .ZN(n9932) );
  AOI22_X1 U12634 ( .A1(n13280), .A2(n9944), .B1(n9995), .B2(SI_18_), .ZN(
        n9931) );
  XNOR2_X1 U12635 ( .A(n13484), .B(n9722), .ZN(n13077) );
  NAND2_X1 U12636 ( .A1(n9933), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U12637 ( .A1(n9947), .A2(n9934), .ZN(n13434) );
  NAND2_X1 U12638 ( .A1(n9746), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U12639 ( .A1(n12338), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9935) );
  OAI211_X1 U12640 ( .C1(n10189), .C2(n15759), .A(n9936), .B(n9935), .ZN(n9937) );
  INV_X1 U12641 ( .A(n9937), .ZN(n9938) );
  NOR2_X1 U12642 ( .A1(n13077), .A2(n13413), .ZN(n9940) );
  NAND2_X1 U12643 ( .A1(n11158), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9957) );
  INV_X1 U12644 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U12645 ( .A1(n11159), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9943) );
  XNOR2_X1 U12646 ( .A(n9956), .B(n9955), .ZN(n10799) );
  NAND2_X1 U12647 ( .A1(n10799), .A2(n9742), .ZN(n9946) );
  AOI22_X1 U12648 ( .A1(n12526), .A2(n9944), .B1(n9995), .B2(n10798), .ZN(
        n9945) );
  XNOR2_X1 U12649 ( .A(n13535), .B(n9715), .ZN(n9954) );
  NAND2_X1 U12650 ( .A1(n9947), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12651 ( .A1(n9962), .A2(n9948), .ZN(n13409) );
  INV_X1 U12652 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13418) );
  NAND2_X1 U12653 ( .A1(n6539), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12654 ( .A1(n12337), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9949) );
  OAI211_X1 U12655 ( .C1(n10176), .C2(n13418), .A(n9950), .B(n9949), .ZN(n9951) );
  INV_X1 U12656 ( .A(n9951), .ZN(n9952) );
  XNOR2_X1 U12657 ( .A(n9954), .B(n13432), .ZN(n13009) );
  XNOR2_X1 U12658 ( .A(n9972), .B(n11203), .ZN(n11182) );
  NAND2_X1 U12659 ( .A1(n11182), .A2(n9742), .ZN(n9961) );
  NAND2_X1 U12660 ( .A1(n9995), .A2(SI_20_), .ZN(n9960) );
  XNOR2_X1 U12661 ( .A(n13057), .B(n9715), .ZN(n9969) );
  NAND2_X1 U12662 ( .A1(n9962), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9963) );
  NAND2_X1 U12663 ( .A1(n9980), .A2(n9963), .ZN(n13064) );
  INV_X1 U12664 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12550) );
  NAND2_X1 U12665 ( .A1(n12338), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U12666 ( .A1(n12337), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9964) );
  OAI211_X1 U12667 ( .C1(n10176), .C2(n12550), .A(n9965), .B(n9964), .ZN(n9966) );
  INV_X1 U12668 ( .A(n9966), .ZN(n9967) );
  XNOR2_X1 U12669 ( .A(n9969), .B(n13395), .ZN(n13060) );
  NAND2_X1 U12670 ( .A1(n13061), .A2(n13060), .ZN(n13059) );
  NAND2_X1 U12671 ( .A1(n11291), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9992) );
  NAND2_X1 U12672 ( .A1(n11288), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U12673 ( .A1(n9995), .A2(SI_21_), .ZN(n9977) );
  XNOR2_X1 U12674 ( .A(n13528), .B(n9715), .ZN(n9988) );
  INV_X1 U12675 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9978) );
  NAND2_X1 U12676 ( .A1(n9980), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U12677 ( .A1(n9999), .A2(n9981), .ZN(n13401) );
  INV_X1 U12678 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U12679 ( .A1(n12337), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9983) );
  NAND2_X1 U12680 ( .A1(n12338), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9982) );
  OAI211_X1 U12681 ( .C1(n9984), .C2(n10176), .A(n9983), .B(n9982), .ZN(n9985)
         );
  INV_X1 U12682 ( .A(n9985), .ZN(n9986) );
  XNOR2_X1 U12683 ( .A(n9988), .B(n13384), .ZN(n13019) );
  INV_X1 U12684 ( .A(n9988), .ZN(n9990) );
  INV_X1 U12685 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9994) );
  XNOR2_X1 U12686 ( .A(n9994), .B(P1_DATAO_REG_22__SCAN_IN), .ZN(n10007) );
  XNOR2_X1 U12687 ( .A(n10008), .B(n10007), .ZN(n11348) );
  NAND2_X1 U12688 ( .A1(n11348), .A2(n9742), .ZN(n9997) );
  NAND2_X1 U12689 ( .A1(n9995), .A2(SI_22_), .ZN(n9996) );
  XNOR2_X1 U12690 ( .A(n13521), .B(n9722), .ZN(n12863) );
  INV_X1 U12691 ( .A(n12863), .ZN(n9998) );
  NAND2_X1 U12692 ( .A1(n9999), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n10000) );
  NAND2_X1 U12693 ( .A1(n10011), .A2(n10000), .ZN(n13388) );
  INV_X1 U12694 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U12695 ( .A1(n12338), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U12696 ( .A1(n12337), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n10001) );
  OAI211_X1 U12697 ( .C1(n10176), .C2(n13387), .A(n10002), .B(n10001), .ZN(
        n10003) );
  INV_X1 U12698 ( .A(n10003), .ZN(n10004) );
  AND2_X1 U12699 ( .A1(n12862), .A2(n12863), .ZN(n10006) );
  XNOR2_X1 U12700 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n10019) );
  XNOR2_X1 U12701 ( .A(n10020), .B(n10019), .ZN(n11729) );
  NAND2_X1 U12702 ( .A1(n11729), .A2(n9742), .ZN(n10010) );
  NAND2_X1 U12703 ( .A1(n9995), .A2(SI_23_), .ZN(n10009) );
  XNOR2_X1 U12704 ( .A(n13373), .B(n10026), .ZN(n13000) );
  NAND2_X1 U12705 ( .A1(n10011), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U12706 ( .A1(n10028), .A2(n10012), .ZN(n13374) );
  INV_X1 U12707 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U12708 ( .A1(n12338), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U12709 ( .A1(n12337), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n10013) );
  OAI211_X1 U12710 ( .C1(n10176), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10016) );
  INV_X1 U12711 ( .A(n10016), .ZN(n10017) );
  AND2_X1 U12712 ( .A1(n13000), .A2(n13385), .ZN(n12858) );
  NAND2_X1 U12713 ( .A1(n11493), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n10021) );
  NAND2_X1 U12714 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  NAND2_X1 U12715 ( .A1(n12181), .A2(n9742), .ZN(n10025) );
  NAND2_X1 U12716 ( .A1(n9995), .A2(SI_24_), .ZN(n10024) );
  XNOR2_X1 U12717 ( .A(n13360), .B(n10026), .ZN(n12865) );
  INV_X1 U12718 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U12719 ( .A1(n10028), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n10029) );
  INV_X1 U12720 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13357) );
  NAND2_X1 U12721 ( .A1(n6539), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U12722 ( .A1(n12337), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n10030) );
  OAI211_X1 U12723 ( .C1(n10176), .C2(n13357), .A(n10031), .B(n10030), .ZN(
        n10032) );
  INV_X1 U12724 ( .A(n10032), .ZN(n10033) );
  XNOR2_X1 U12725 ( .A(n12865), .B(n13031), .ZN(n10035) );
  INV_X1 U12726 ( .A(n13000), .ZN(n12867) );
  NAND2_X1 U12727 ( .A1(n12867), .A2(n13073), .ZN(n12866) );
  NAND3_X1 U12728 ( .A1(n13002), .A2(n12866), .A3(n10035), .ZN(n10065) );
  NOR2_X1 U12729 ( .A1(n13369), .A2(n13385), .ZN(n12868) );
  INV_X1 U12730 ( .A(n12868), .ZN(n10037) );
  AOI21_X1 U12731 ( .B1(n13369), .B2(n13385), .A(n12867), .ZN(n10036) );
  AOI21_X1 U12732 ( .B1(n12867), .B2(n10037), .A(n10036), .ZN(n10041) );
  AOI21_X1 U12733 ( .B1(n13031), .B2(n13385), .A(n12867), .ZN(n10039) );
  AOI21_X1 U12734 ( .B1(n13073), .B2(n13369), .A(n13000), .ZN(n10038) );
  OAI21_X1 U12735 ( .B1(n10039), .B2(n10038), .A(n12865), .ZN(n10040) );
  OAI21_X1 U12736 ( .B1(n10041), .B2(n12865), .A(n10040), .ZN(n10063) );
  NAND2_X1 U12737 ( .A1(n10042), .A2(n10043), .ZN(n10205) );
  XNOR2_X1 U12738 ( .A(n12367), .B(n10205), .ZN(n10045) );
  NAND2_X1 U12739 ( .A1(n10042), .A2(n12526), .ZN(n10044) );
  NAND2_X1 U12740 ( .A1(n10045), .A2(n10044), .ZN(n10239) );
  NAND2_X1 U12741 ( .A1(n10239), .A2(n11358), .ZN(n10928) );
  OAI22_X1 U12742 ( .A1(n10049), .A2(P3_D_REG_1__SCAN_IN), .B1(n10047), .B2(
        n10046), .ZN(n10208) );
  INV_X1 U12743 ( .A(n10208), .ZN(n10338) );
  INV_X1 U12744 ( .A(n10049), .ZN(n10397) );
  NOR4_X1 U12745 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n10058) );
  INV_X1 U12746 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n15907) );
  INV_X1 U12747 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n15790) );
  INV_X1 U12748 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15843) );
  INV_X1 U12749 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n15840) );
  NAND4_X1 U12750 ( .A1(n15907), .A2(n15790), .A3(n15843), .A4(n15840), .ZN(
        n10055) );
  NOR4_X1 U12751 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n10053) );
  NOR4_X1 U12752 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n10052) );
  NOR4_X1 U12753 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n10051) );
  NOR4_X1 U12754 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n10050) );
  NAND4_X1 U12755 ( .A1(n10053), .A2(n10052), .A3(n10051), .A4(n10050), .ZN(
        n10054) );
  NOR4_X1 U12756 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        n10055), .A4(n10054), .ZN(n10057) );
  NOR4_X1 U12757 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n10056) );
  NAND3_X1 U12758 ( .A1(n10058), .A2(n10057), .A3(n10056), .ZN(n10059) );
  NAND2_X1 U12759 ( .A1(n10397), .A2(n10059), .ZN(n10211) );
  NAND3_X1 U12760 ( .A1(n10338), .A2(n10341), .A3(n10211), .ZN(n10244) );
  NAND2_X1 U12761 ( .A1(n12367), .A2(n12522), .ZN(n10207) );
  OR2_X1 U12762 ( .A1(n10207), .A2(n10060), .ZN(n10241) );
  NAND2_X1 U12763 ( .A1(n10208), .A2(n10048), .ZN(n10213) );
  INV_X1 U12764 ( .A(n10211), .ZN(n10061) );
  INV_X1 U12765 ( .A(n10238), .ZN(n10091) );
  OAI22_X1 U12766 ( .A1(n10928), .A2(n10244), .B1(n10241), .B2(n10091), .ZN(
        n10062) );
  INV_X1 U12767 ( .A(n10244), .ZN(n10066) );
  INV_X1 U12768 ( .A(n11358), .ZN(n13485) );
  NAND3_X1 U12769 ( .A1(n10066), .A2(n10242), .A3(n13485), .ZN(n10068) );
  NAND2_X1 U12770 ( .A1(n15679), .A2(n10242), .ZN(n10067) );
  NAND2_X1 U12771 ( .A1(n10069), .A2(n7072), .ZN(n10088) );
  INV_X1 U12772 ( .A(n10073), .ZN(n10072) );
  INV_X1 U12773 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U12774 ( .A1(n10073), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U12775 ( .A1(n10142), .A2(n10074), .ZN(n13346) );
  INV_X1 U12776 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n13345) );
  NAND2_X1 U12777 ( .A1(n6539), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U12778 ( .A1(n12337), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n10075) );
  OAI211_X1 U12779 ( .C1(n10176), .C2(n13345), .A(n10076), .B(n10075), .ZN(
        n10077) );
  INV_X1 U12780 ( .A(n10077), .ZN(n10078) );
  INV_X1 U12781 ( .A(n10080), .ZN(n13358) );
  INV_X1 U12782 ( .A(n10232), .ZN(n12514) );
  AND3_X1 U12783 ( .A1(n10204), .A2(n10082), .A3(n10081), .ZN(n10084) );
  NAND2_X1 U12784 ( .A1(n10239), .A2(n10244), .ZN(n10083) );
  OAI211_X1 U12785 ( .C1(n10238), .C2(n10241), .A(n10084), .B(n10083), .ZN(
        n10085) );
  NAND2_X1 U12786 ( .A1(n10085), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10087) );
  NAND2_X1 U12787 ( .A1(n9474), .A2(n10090), .ZN(n10245) );
  OR2_X1 U12788 ( .A1(n10245), .A2(n10238), .ZN(n10086) );
  NAND2_X2 U12789 ( .A1(n10087), .A2(n10086), .ZN(n13090) );
  INV_X1 U12790 ( .A(n13090), .ZN(n11661) );
  INV_X1 U12791 ( .A(n10088), .ZN(n10089) );
  AND2_X2 U12792 ( .A1(n9474), .A2(n10089), .ZN(n13352) );
  NAND2_X1 U12793 ( .A1(n13352), .A2(n10090), .ZN(n12533) );
  AOI22_X1 U12794 ( .A1(n13385), .A2(n13069), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10092) );
  OAI21_X1 U12795 ( .B1(n13358), .B2(n11661), .A(n10092), .ZN(n10093) );
  AOI21_X1 U12796 ( .B1(n13089), .B2(n13353), .A(n10093), .ZN(n10094) );
  INV_X1 U12797 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10215) );
  NAND2_X1 U12798 ( .A1(n11631), .A2(n13112), .ZN(n12388) );
  NAND2_X1 U12799 ( .A1(n12392), .A2(n12390), .ZN(n11121) );
  NAND2_X1 U12800 ( .A1(n11657), .A2(n11631), .ZN(n11119) );
  NAND2_X1 U12801 ( .A1(n11169), .A2(n13111), .ZN(n10096) );
  INV_X1 U12802 ( .A(n11644), .ZN(n11094) );
  AND2_X1 U12803 ( .A1(n11121), .A2(n11119), .ZN(n10105) );
  NAND2_X1 U12804 ( .A1(n10098), .A2(n10097), .ZN(n12368) );
  NAND2_X1 U12805 ( .A1(n10098), .A2(n11357), .ZN(n10099) );
  NAND2_X1 U12806 ( .A1(n10100), .A2(n10099), .ZN(n11040) );
  NAND2_X1 U12807 ( .A1(n11044), .A2(n13115), .ZN(n12372) );
  NAND2_X1 U12808 ( .A1(n11414), .A2(n11405), .ZN(n12371) );
  NAND2_X1 U12809 ( .A1(n11040), .A2(n12483), .ZN(n10102) );
  NAND2_X1 U12810 ( .A1(n11414), .A2(n11044), .ZN(n10101) );
  NAND2_X1 U12811 ( .A1(n10102), .A2(n10101), .ZN(n11028) );
  NAND2_X1 U12812 ( .A1(n11220), .A2(n13114), .ZN(n12377) );
  NAND2_X1 U12813 ( .A1(n11403), .A2(n11395), .ZN(n12376) );
  INV_X1 U12814 ( .A(n11507), .ZN(n11246) );
  INV_X1 U12815 ( .A(n11632), .ZN(n13113) );
  NAND2_X1 U12816 ( .A1(n11246), .A2(n13113), .ZN(n12380) );
  NAND2_X1 U12817 ( .A1(n11632), .A2(n11507), .ZN(n12381) );
  AND2_X1 U12818 ( .A1(n11395), .A2(n13114), .ZN(n11066) );
  AOI22_X1 U12819 ( .A1(n11064), .A2(n11066), .B1(n11507), .B2(n13113), .ZN(
        n10103) );
  OAI21_X2 U12820 ( .B1(n11028), .B2(n10104), .A(n10103), .ZN(n11133) );
  OR2_X1 U12821 ( .A1(n11819), .A2(n10107), .ZN(n12398) );
  NAND2_X1 U12822 ( .A1(n11819), .A2(n10107), .ZN(n12399) );
  NAND2_X1 U12823 ( .A1(n12398), .A2(n12399), .ZN(n12493) );
  INV_X1 U12824 ( .A(n10107), .ZN(n13109) );
  OR2_X1 U12825 ( .A1(n11819), .A2(n13109), .ZN(n10108) );
  XNOR2_X1 U12826 ( .A(n11793), .B(n13108), .ZN(n12497) );
  OR2_X1 U12827 ( .A1(n11793), .A2(n11905), .ZN(n10109) );
  OR2_X1 U12828 ( .A1(n11910), .A2(n13107), .ZN(n12411) );
  NAND2_X1 U12829 ( .A1(n11910), .A2(n13107), .ZN(n12409) );
  NAND2_X1 U12830 ( .A1(n12411), .A2(n12409), .ZN(n12494) );
  OR2_X1 U12831 ( .A1(n11910), .A2(n12242), .ZN(n10110) );
  OR2_X1 U12832 ( .A1(n12240), .A2(n13106), .ZN(n12410) );
  NAND2_X1 U12833 ( .A1(n11280), .A2(n12498), .ZN(n11278) );
  OR2_X1 U12834 ( .A1(n12240), .A2(n12255), .ZN(n11319) );
  NAND2_X1 U12835 ( .A1(n11278), .A2(n11319), .ZN(n10111) );
  NAND2_X1 U12836 ( .A1(n12256), .A2(n13105), .ZN(n12417) );
  NAND2_X1 U12837 ( .A1(n11498), .A2(n12209), .ZN(n12416) );
  NAND2_X1 U12838 ( .A1(n12417), .A2(n12416), .ZN(n12499) );
  NAND2_X1 U12839 ( .A1(n11498), .A2(n13105), .ZN(n10112) );
  NAND2_X1 U12840 ( .A1(n12420), .A2(n12266), .ZN(n10113) );
  INV_X1 U12841 ( .A(n12420), .ZN(n10220) );
  NAND2_X1 U12842 ( .A1(n10220), .A2(n13104), .ZN(n10114) );
  OR2_X1 U12843 ( .A1(n12267), .A2(n12207), .ZN(n12431) );
  NAND2_X1 U12844 ( .A1(n12267), .A2(n12207), .ZN(n12425) );
  OR2_X1 U12845 ( .A1(n12267), .A2(n12300), .ZN(n10115) );
  INV_X1 U12846 ( .A(n12302), .ZN(n10222) );
  NAND2_X1 U12847 ( .A1(n10222), .A2(n13039), .ZN(n10117) );
  OR2_X1 U12848 ( .A1(n13042), .A2(n12275), .ZN(n12427) );
  NAND2_X1 U12849 ( .A1(n13042), .A2(n12275), .ZN(n12439) );
  NAND2_X1 U12850 ( .A1(n13051), .A2(n13102), .ZN(n12358) );
  NAND2_X1 U12851 ( .A1(n12288), .A2(n13430), .ZN(n12351) );
  NAND2_X1 U12852 ( .A1(n12358), .A2(n12351), .ZN(n12505) );
  NAND2_X1 U12853 ( .A1(n12288), .A2(n13102), .ZN(n10118) );
  NAND2_X1 U12854 ( .A1(n13484), .A2(n13413), .ZN(n12355) );
  INV_X1 U12855 ( .A(n13484), .ZN(n13082) );
  NAND2_X1 U12856 ( .A1(n13082), .A2(n13413), .ZN(n10119) );
  NAND2_X1 U12857 ( .A1(n13535), .A2(n13101), .ZN(n12357) );
  OR2_X1 U12858 ( .A1(n13535), .A2(n13432), .ZN(n10121) );
  NAND2_X1 U12859 ( .A1(n13057), .A2(n13395), .ZN(n10122) );
  NAND2_X1 U12860 ( .A1(n13528), .A2(n13384), .ZN(n12350) );
  NAND2_X1 U12861 ( .A1(n13024), .A2(n9989), .ZN(n12349) );
  NAND2_X1 U12862 ( .A1(n13528), .A2(n9989), .ZN(n10123) );
  NOR2_X1 U12863 ( .A1(n13521), .A2(n13397), .ZN(n10125) );
  INV_X1 U12864 ( .A(n13521), .ZN(n10124) );
  NAND2_X1 U12865 ( .A1(n13373), .A2(n13073), .ZN(n12457) );
  NAND2_X1 U12866 ( .A1(n12453), .A2(n12457), .ZN(n13367) );
  NAND2_X1 U12867 ( .A1(n13373), .A2(n13385), .ZN(n10126) );
  XNOR2_X1 U12868 ( .A(n11770), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n10128) );
  NAND2_X1 U12869 ( .A1(n13556), .A2(n9742), .ZN(n10130) );
  NAND2_X1 U12870 ( .A1(n9995), .A2(SI_25_), .ZN(n10129) );
  NAND2_X1 U12871 ( .A1(n12874), .A2(n13353), .ZN(n10131) );
  OR2_X1 U12872 ( .A1(n13360), .A2(n13369), .ZN(n13336) );
  AND2_X1 U12873 ( .A1(n10132), .A2(n13336), .ZN(n10133) );
  NAND2_X1 U12874 ( .A1(n13507), .A2(n13353), .ZN(n10134) );
  NAND2_X1 U12875 ( .A1(n11770), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n10135) );
  NAND2_X1 U12876 ( .A1(n10136), .A2(n10135), .ZN(n10138) );
  NAND2_X1 U12877 ( .A1(n11774), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n10137) );
  XNOR2_X1 U12878 ( .A(n14479), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n10139) );
  XNOR2_X1 U12879 ( .A(n10151), .B(n10139), .ZN(n13553) );
  NAND2_X1 U12880 ( .A1(n13553), .A2(n9742), .ZN(n10141) );
  NAND2_X1 U12881 ( .A1(n9995), .A2(SI_26_), .ZN(n10140) );
  NAND2_X1 U12882 ( .A1(n10142), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n10143) );
  NAND2_X1 U12883 ( .A1(n10157), .A2(n10143), .ZN(n13328) );
  INV_X1 U12884 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n10146) );
  NAND2_X1 U12885 ( .A1(n12337), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U12886 ( .A1(n12338), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n10144) );
  OAI211_X1 U12887 ( .C1(n10176), .C2(n10146), .A(n10145), .B(n10144), .ZN(
        n10147) );
  INV_X1 U12888 ( .A(n10147), .ZN(n10148) );
  OR2_X1 U12889 ( .A1(n13327), .A2(n13342), .ZN(n10150) );
  NAND2_X1 U12890 ( .A1(n14479), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n10152) );
  XNOR2_X1 U12891 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n10153) );
  NAND2_X1 U12892 ( .A1(n9995), .A2(SI_27_), .ZN(n10154) );
  INV_X1 U12893 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15909) );
  NAND2_X1 U12894 ( .A1(n10157), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U12895 ( .A1(n10171), .A2(n10158), .ZN(n13315) );
  INV_X1 U12896 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n15829) );
  NAND2_X1 U12897 ( .A1(n9746), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U12898 ( .A1(n12338), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n10159) );
  OAI211_X1 U12899 ( .C1(n10189), .C2(n15829), .A(n10160), .B(n10159), .ZN(
        n10161) );
  INV_X1 U12900 ( .A(n10161), .ZN(n10162) );
  OR2_X1 U12901 ( .A1(n12991), .A2(n13324), .ZN(n10164) );
  AND2_X1 U12902 ( .A1(n12317), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n10166) );
  NAND2_X1 U12903 ( .A1(n15229), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n10165) );
  XNOR2_X1 U12904 ( .A(n10182), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n10168) );
  XNOR2_X1 U12905 ( .A(n10181), .B(n10168), .ZN(n13546) );
  NAND2_X1 U12906 ( .A1(n13546), .A2(n9742), .ZN(n10170) );
  NAND2_X1 U12907 ( .A1(n9995), .A2(SI_28_), .ZN(n10169) );
  NAND2_X1 U12908 ( .A1(n10171), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U12909 ( .A1(n10263), .A2(n10172), .ZN(n13303) );
  INV_X1 U12910 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U12911 ( .A1(n6539), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n10174) );
  NAND2_X1 U12912 ( .A1(n12337), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n10173) );
  OAI211_X1 U12913 ( .C1(n10176), .C2(n10175), .A(n10174), .B(n10173), .ZN(
        n10177) );
  NAND2_X1 U12914 ( .A1(n10178), .A2(n10201), .ZN(n12470) );
  INV_X1 U12915 ( .A(n10201), .ZN(n13310) );
  NAND2_X1 U12916 ( .A1(n10178), .A2(n13310), .ZN(n10179) );
  AND2_X1 U12917 ( .A1(n12319), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10180) );
  NAND2_X1 U12918 ( .A1(n10182), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n10183) );
  XNOR2_X1 U12919 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12320) );
  XNOR2_X1 U12920 ( .A(n12322), .B(n12320), .ZN(n12963) );
  NAND2_X1 U12921 ( .A1(n12963), .A2(n9742), .ZN(n10185) );
  NAND2_X1 U12922 ( .A1(n9995), .A2(SI_29_), .ZN(n10184) );
  INV_X1 U12923 ( .A(n10263), .ZN(n10186) );
  NAND2_X1 U12924 ( .A1(n9746), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n10188) );
  NAND2_X1 U12925 ( .A1(n12338), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10187) );
  OAI211_X1 U12926 ( .C1(n10215), .C2(n10189), .A(n10188), .B(n10187), .ZN(
        n10190) );
  INV_X1 U12927 ( .A(n10190), .ZN(n10191) );
  NAND2_X1 U12928 ( .A1(n12343), .A2(n10191), .ZN(n13300) );
  NAND2_X1 U12929 ( .A1(n10192), .A2(n13300), .ZN(n12516) );
  INV_X1 U12930 ( .A(n13300), .ZN(n12886) );
  NAND2_X1 U12931 ( .A1(n10264), .A2(n12886), .ZN(n12346) );
  NAND2_X1 U12932 ( .A1(n9625), .A2(n10193), .ZN(n12525) );
  INV_X1 U12933 ( .A(n13352), .ZN(n13431) );
  NAND2_X1 U12934 ( .A1(n12338), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n10196) );
  NAND2_X1 U12935 ( .A1(n9746), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n10195) );
  NAND2_X1 U12936 ( .A1(n12337), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n10194) );
  AND3_X1 U12937 ( .A1(n10196), .A2(n10195), .A3(n10194), .ZN(n10197) );
  NAND2_X1 U12938 ( .A1(n12343), .A2(n10197), .ZN(n13100) );
  NAND2_X1 U12939 ( .A1(n10198), .A2(P3_B_REG_SCAN_IN), .ZN(n10199) );
  AND2_X1 U12940 ( .A1(n13396), .A2(n10199), .ZN(n13289) );
  NAND2_X1 U12941 ( .A1(n13100), .A2(n13289), .ZN(n10200) );
  OAI21_X1 U12942 ( .B1(n10201), .B2(n13431), .A(n10200), .ZN(n10202) );
  NOR2_X1 U12943 ( .A1(n10043), .A2(n12522), .ZN(n10203) );
  NAND2_X1 U12944 ( .A1(n12367), .A2(n10203), .ZN(n10233) );
  NAND2_X1 U12945 ( .A1(n12462), .A2(n10233), .ZN(n10251) );
  NAND2_X1 U12946 ( .A1(n10204), .A2(n10251), .ZN(n10254) );
  NAND2_X1 U12947 ( .A1(n12531), .A2(n10205), .ZN(n10206) );
  NAND3_X1 U12948 ( .A1(n10207), .A2(n10206), .A3(n10232), .ZN(n10209) );
  NAND3_X1 U12949 ( .A1(n10209), .A2(n12462), .A3(n10208), .ZN(n10210) );
  OAI21_X1 U12950 ( .B1(n10254), .B2(n10341), .A(n10210), .ZN(n10214) );
  AND2_X1 U12951 ( .A1(n10211), .A2(n10242), .ZN(n10212) );
  MUX2_X1 U12952 ( .A(n10215), .B(n10257), .S(n13486), .Z(n10237) );
  INV_X1 U12953 ( .A(n12510), .ZN(n10231) );
  INV_X1 U12954 ( .A(n12380), .ZN(n10217) );
  OAI21_X1 U12955 ( .B1(n12376), .B2(n10217), .A(n12381), .ZN(n10218) );
  INV_X1 U12956 ( .A(n10218), .ZN(n10219) );
  NAND2_X1 U12957 ( .A1(n11793), .A2(n13108), .ZN(n12403) );
  OR2_X1 U12958 ( .A1(n11793), .A2(n13108), .ZN(n12404) );
  NAND2_X1 U12959 ( .A1(n11325), .A2(n7893), .ZN(n11324) );
  NAND2_X1 U12960 ( .A1(n12420), .A2(n13104), .ZN(n12430) );
  NAND2_X1 U12961 ( .A1(n10222), .A2(n13103), .ZN(n12426) );
  NAND2_X1 U12962 ( .A1(n12302), .A2(n13039), .ZN(n12438) );
  INV_X1 U12963 ( .A(n12358), .ZN(n10224) );
  AND2_X1 U12964 ( .A1(n12439), .A2(n12351), .ZN(n10223) );
  INV_X1 U12965 ( .A(n12357), .ZN(n10225) );
  OR2_X1 U12966 ( .A1(n13057), .A2(n13414), .ZN(n12445) );
  NAND2_X1 U12967 ( .A1(n13521), .A2(n13022), .ZN(n12347) );
  NAND2_X1 U12968 ( .A1(n10226), .A2(n12348), .ZN(n13366) );
  INV_X1 U12969 ( .A(n13367), .ZN(n12509) );
  NAND2_X1 U12970 ( .A1(n13360), .A2(n13031), .ZN(n12456) );
  NAND2_X1 U12971 ( .A1(n13327), .A2(n12996), .ZN(n12460) );
  NAND2_X1 U12972 ( .A1(n12991), .A2(n12888), .ZN(n12469) );
  INV_X1 U12973 ( .A(n12470), .ZN(n10230) );
  XOR2_X1 U12974 ( .A(n10231), .B(n12518), .Z(n10260) );
  OR2_X1 U12975 ( .A1(n10928), .A2(n10232), .ZN(n10234) );
  NAND2_X1 U12976 ( .A1(n12531), .A2(n15679), .ZN(n11359) );
  NAND2_X1 U12977 ( .A1(n13474), .A2(n13486), .ZN(n13488) );
  NAND2_X1 U12978 ( .A1(n10264), .A2(n13469), .ZN(n10235) );
  NAND2_X1 U12979 ( .A1(n10239), .A2(n10238), .ZN(n10240) );
  OAI21_X1 U12980 ( .B1(n10241), .B2(n10244), .A(n10240), .ZN(n10243) );
  NAND2_X1 U12981 ( .A1(n10243), .A2(n10242), .ZN(n10247) );
  NAND2_X1 U12982 ( .A1(n10264), .A2(n13520), .ZN(n10248) );
  INV_X1 U12983 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U12984 ( .A1(n10251), .A2(n10338), .ZN(n10253) );
  NAND2_X1 U12985 ( .A1(n10254), .A2(n10341), .ZN(n10255) );
  NAND2_X1 U12986 ( .A1(n10256), .A2(n10255), .ZN(n10262) );
  NAND2_X1 U12987 ( .A1(n15679), .A2(n9625), .ZN(n15677) );
  NAND2_X1 U12988 ( .A1(n13313), .A2(n15677), .ZN(n10259) );
  OR2_X1 U12989 ( .A1(n10260), .A2(n13441), .ZN(n10266) );
  OR2_X1 U12990 ( .A1(n11358), .A2(n15679), .ZN(n10261) );
  NOR2_X1 U12991 ( .A1(n10263), .A2(n15681), .ZN(n13291) );
  AOI21_X1 U12992 ( .B1(n10264), .B2(n13438), .A(n13291), .ZN(n10265) );
  INV_X1 U12993 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10273) );
  INV_X1 U12994 ( .A(n10268), .ZN(n10269) );
  AOI211_X1 U12995 ( .C1(n13859), .C2(n14105), .A(n10269), .B(n8582), .ZN(
        n14094) );
  XNOR2_X1 U12996 ( .A(n14129), .B(n13665), .ZN(n14124) );
  INV_X1 U12997 ( .A(n14124), .ZN(n10270) );
  NAND3_X1 U12998 ( .A1(n14121), .A2(n14103), .A3(n14098), .ZN(n14099) );
  NAND2_X1 U12999 ( .A1(n14099), .A2(n10271), .ZN(n10272) );
  AOI22_X1 U13000 ( .A1(n13963), .A2(n14304), .B1(n14302), .B2(n13965), .ZN(
        n12900) );
  XOR2_X1 U13001 ( .A(n13928), .B(n10274), .Z(n14097) );
  NAND2_X1 U13002 ( .A1(n10276), .A2(n10275), .ZN(P2_U3524) );
  INV_X1 U13003 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10277) );
  NAND2_X1 U13004 ( .A1(n10279), .A2(n10278), .ZN(P2_U3492) );
  INV_X1 U13005 ( .A(n11490), .ZN(n10280) );
  NOR2_X1 U13006 ( .A1(n10281), .A2(n10280), .ZN(n10486) );
  INV_X1 U13007 ( .A(n10515), .ZN(n10554) );
  NAND3_X1 U13008 ( .A1(n13208), .A2(n10283), .A3(n10282), .ZN(n10284) );
  AOI21_X1 U13009 ( .B1(n10285), .B2(n10284), .A(n13288), .ZN(n10297) );
  NAND3_X1 U13010 ( .A1(n13195), .A2(n10287), .A3(n10286), .ZN(n10288) );
  AOI21_X1 U13011 ( .B1(n10289), .B2(n10288), .A(n13242), .ZN(n10296) );
  AOI211_X1 U13012 ( .C1(n10292), .C2(n10291), .A(n13277), .B(n10290), .ZN(
        n10295) );
  NAND2_X1 U13013 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12264)
         );
  NAND2_X1 U13014 ( .A1(n15694), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n10293) );
  OAI211_X1 U13015 ( .C1(n13261), .C2(n10518), .A(n12264), .B(n10293), .ZN(
        n10294) );
  INV_X1 U13016 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U13017 ( .A1(n10298), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n10299) );
  NAND2_X1 U13018 ( .A1(n10308), .A2(n10299), .ZN(n10300) );
  INV_X1 U13019 ( .A(n10300), .ZN(n10302) );
  INV_X1 U13020 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10301) );
  AND2_X1 U13021 ( .A1(n10300), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n15241) );
  AOI21_X1 U13022 ( .B1(n10302), .B2(n10301), .A(n15241), .ZN(SUB_1596_U53) );
  NAND2_X1 U13023 ( .A1(n15240), .A2(n15241), .ZN(n10306) );
  INV_X1 U13024 ( .A(n10303), .ZN(n10304) );
  NAND2_X1 U13025 ( .A1(n10304), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10305) );
  INV_X1 U13026 ( .A(n10318), .ZN(n10311) );
  INV_X1 U13027 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n15695) );
  NAND2_X1 U13028 ( .A1(n15695), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U13029 ( .A1(n10308), .A2(n10307), .ZN(n10310) );
  INV_X1 U13030 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10832) );
  NAND2_X1 U13031 ( .A1(n10832), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n10309) );
  NAND2_X1 U13032 ( .A1(n10310), .A2(n10309), .ZN(n10319) );
  XNOR2_X1 U13033 ( .A(n10319), .B(n10311), .ZN(n10312) );
  INV_X1 U13034 ( .A(n10312), .ZN(n10313) );
  NAND2_X1 U13035 ( .A1(n10314), .A2(n10313), .ZN(n10315) );
  INV_X1 U13036 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10316) );
  NAND2_X1 U13037 ( .A1(n10316), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10317) );
  XNOR2_X1 U13038 ( .A(n10375), .B(n10320), .ZN(n10374) );
  XNOR2_X1 U13039 ( .A(n10374), .B(n14685), .ZN(n10321) );
  NAND2_X1 U13040 ( .A1(n10322), .A2(n10321), .ZN(n10323) );
  OAI21_X1 U13041 ( .B1(n6602), .B2(n7150), .A(n10373), .ZN(SUB_1596_U60) );
  AND2_X1 U13042 ( .A1(n10425), .A2(P3_U3151), .ZN(n11728) );
  INV_X2 U13043 ( .A(n11728), .ZN(n12962) );
  NOR2_X1 U13044 ( .A1(n10425), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12800) );
  INV_X2 U13045 ( .A(n12800), .ZN(n13550) );
  OAI222_X1 U13046 ( .A1(n10326), .A2(P3_U3151), .B1(n12962), .B2(n10325), 
        .C1(n10324), .C2(n13550), .ZN(P3_U3293) );
  OAI222_X1 U13047 ( .A1(n10329), .A2(P3_U3151), .B1(n12962), .B2(n10328), 
        .C1(n10327), .C2(n13550), .ZN(P3_U3291) );
  INV_X1 U13048 ( .A(n10330), .ZN(n10332) );
  INV_X1 U13049 ( .A(SI_6_), .ZN(n10331) );
  OAI222_X1 U13050 ( .A1(n13143), .A2(P3_U3151), .B1(n12962), .B2(n10332), 
        .C1(n10331), .C2(n13550), .ZN(P3_U3289) );
  INV_X1 U13051 ( .A(SI_5_), .ZN(n10333) );
  OAI222_X1 U13052 ( .A1(n10849), .A2(P3_U3151), .B1(n12962), .B2(n10334), 
        .C1(n10333), .C2(n13550), .ZN(P3_U3290) );
  OAI222_X1 U13053 ( .A1(n10337), .A2(P3_U3151), .B1(n12962), .B2(n10336), 
        .C1(n10335), .C2(n13550), .ZN(P3_U3292) );
  INV_X1 U13054 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U13055 ( .A1(n10338), .A2(n10395), .ZN(n10339) );
  OAI21_X1 U13056 ( .B1(n10395), .B2(n10340), .A(n10339), .ZN(P3_U3377) );
  INV_X1 U13057 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10343) );
  NAND2_X1 U13058 ( .A1(n10341), .A2(n10395), .ZN(n10342) );
  OAI21_X1 U13059 ( .B1(n10395), .B2(n10343), .A(n10342), .ZN(P3_U3376) );
  AOI22_X1 U13060 ( .A1(n11728), .A2(n10344), .B1(P3_IR_REG_0__SCAN_IN), .B2(
        P3_STATE_REG_SCAN_IN), .ZN(n10345) );
  OAI21_X1 U13061 ( .B1(n13550), .B2(n10346), .A(n10345), .ZN(P3_U3295) );
  AND2_X1 U13062 ( .A1(n9647), .A2(P1_U3086), .ZN(n10442) );
  INV_X2 U13063 ( .A(n10442), .ZN(n15232) );
  NOR2_X1 U13064 ( .A1(n9647), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15221) );
  INV_X1 U13065 ( .A(n10348), .ZN(n12537) );
  INV_X1 U13066 ( .A(n14676), .ZN(n14674) );
  OAI222_X1 U13067 ( .A1(n15232), .A2(n10349), .B1(n15236), .B2(n12537), .C1(
        P1_U3086), .C2(n14674), .ZN(P1_U3353) );
  INV_X1 U13068 ( .A(n10350), .ZN(n10431) );
  INV_X1 U13069 ( .A(n15339), .ZN(n10351) );
  OAI222_X1 U13070 ( .A1(n15232), .A2(n10352), .B1(n15236), .B2(n10431), .C1(
        n6537), .C2(n10351), .ZN(P1_U3351) );
  OAI222_X1 U13071 ( .A1(n12962), .A2(n10353), .B1(n13550), .B2(n15702), .C1(
        P3_U3151), .C2(n10836), .ZN(P3_U3294) );
  OAI222_X1 U13072 ( .A1(P3_U3151), .A2(n10786), .B1(n13550), .B2(n10355), 
        .C1(n12962), .C2(n10354), .ZN(P3_U3288) );
  OAI222_X1 U13073 ( .A1(P3_U3151), .A2(n10358), .B1(n13550), .B2(n10357), 
        .C1(n12962), .C2(n10356), .ZN(P3_U3286) );
  INV_X1 U13074 ( .A(SI_8_), .ZN(n10361) );
  INV_X1 U13075 ( .A(n10359), .ZN(n10360) );
  OAI222_X1 U13076 ( .A1(P3_U3151), .A2(n10362), .B1(n13550), .B2(n10361), 
        .C1(n12962), .C2(n10360), .ZN(P3_U3287) );
  INV_X1 U13077 ( .A(n10363), .ZN(n10433) );
  INV_X1 U13078 ( .A(n14691), .ZN(n10364) );
  OAI222_X1 U13079 ( .A1(n15232), .A2(n7936), .B1(n15236), .B2(n10433), .C1(
        P1_U3086), .C2(n10364), .ZN(P1_U3352) );
  OAI222_X1 U13080 ( .A1(P3_U3151), .A2(n10367), .B1(n13550), .B2(n10366), 
        .C1(n12962), .C2(n10365), .ZN(P3_U3285) );
  OAI222_X1 U13081 ( .A1(n15236), .A2(n10429), .B1(n14656), .B2(n6537), .C1(
        n10368), .C2(n15232), .ZN(P1_U3354) );
  OAI222_X1 U13082 ( .A1(n13166), .A2(P3_U3151), .B1(n12962), .B2(n10369), 
        .C1(n13550), .C2(n15810), .ZN(P3_U3284) );
  INV_X1 U13083 ( .A(n14716), .ZN(n10370) );
  OAI222_X1 U13084 ( .A1(n15232), .A2(n10371), .B1(n15236), .B2(n10437), .C1(
        n6537), .C2(n10370), .ZN(P1_U3349) );
  NAND2_X1 U13085 ( .A1(n10374), .A2(n14685), .ZN(n10377) );
  NAND2_X1 U13086 ( .A1(n10375), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10376) );
  INV_X1 U13087 ( .A(n10378), .ZN(n10379) );
  INV_X1 U13088 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10380) );
  NAND2_X1 U13089 ( .A1(n10381), .A2(n10380), .ZN(n10384) );
  NAND2_X1 U13090 ( .A1(n10382), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10383) );
  INV_X1 U13091 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n10385) );
  INV_X1 U13092 ( .A(n10387), .ZN(n10386) );
  INV_X1 U13093 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10389) );
  OAI21_X1 U13094 ( .B1(n6729), .B2(n10389), .A(n10751), .ZN(SUB_1596_U58) );
  INV_X1 U13095 ( .A(n10390), .ZN(n10427) );
  AOI22_X1 U13096 ( .A1(n14734), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10442), .ZN(n10391) );
  OAI21_X1 U13097 ( .B1(n10427), .B2(n15236), .A(n10391), .ZN(P1_U3348) );
  INV_X1 U13098 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10394) );
  INV_X1 U13099 ( .A(n10392), .ZN(n10435) );
  INV_X1 U13100 ( .A(n14706), .ZN(n10393) );
  OAI222_X1 U13101 ( .A1(n15232), .A2(n10394), .B1(n15236), .B2(n10435), .C1(
        P1_U3086), .C2(n10393), .ZN(P1_U3350) );
  INV_X1 U13102 ( .A(n10395), .ZN(n10396) );
  NOR2_X1 U13103 ( .A1(n10397), .A2(n10396), .ZN(n10399) );
  CLKBUF_X1 U13104 ( .A(n10399), .Z(n10423) );
  NOR2_X1 U13105 ( .A1(n10423), .A2(n15843), .ZN(P3_U3253) );
  NOR2_X1 U13106 ( .A1(n10423), .A2(n15790), .ZN(P3_U3256) );
  INV_X1 U13107 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10398) );
  NOR2_X1 U13108 ( .A1(n10423), .A2(n10398), .ZN(P3_U3257) );
  INV_X1 U13109 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n15859) );
  NOR2_X1 U13110 ( .A1(n10423), .A2(n15859), .ZN(P3_U3234) );
  INV_X1 U13111 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10400) );
  NOR2_X1 U13112 ( .A1(n10399), .A2(n10400), .ZN(P3_U3262) );
  INV_X1 U13113 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10401) );
  NOR2_X1 U13114 ( .A1(n10423), .A2(n10401), .ZN(P3_U3252) );
  INV_X1 U13115 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10402) );
  NOR2_X1 U13116 ( .A1(n10423), .A2(n10402), .ZN(P3_U3254) );
  INV_X1 U13117 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10403) );
  NOR2_X1 U13118 ( .A1(n10399), .A2(n10403), .ZN(P3_U3242) );
  INV_X1 U13119 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10404) );
  NOR2_X1 U13120 ( .A1(n10399), .A2(n10404), .ZN(P3_U3243) );
  INV_X1 U13121 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10405) );
  NOR2_X1 U13122 ( .A1(n10399), .A2(n10405), .ZN(P3_U3244) );
  INV_X1 U13123 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10406) );
  NOR2_X1 U13124 ( .A1(n10399), .A2(n10406), .ZN(P3_U3258) );
  INV_X1 U13125 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10407) );
  NOR2_X1 U13126 ( .A1(n10423), .A2(n10407), .ZN(P3_U3259) );
  INV_X1 U13127 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10408) );
  NOR2_X1 U13128 ( .A1(n10399), .A2(n10408), .ZN(P3_U3240) );
  INV_X1 U13129 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10409) );
  NOR2_X1 U13130 ( .A1(n10399), .A2(n10409), .ZN(P3_U3241) );
  INV_X1 U13131 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10410) );
  NOR2_X1 U13132 ( .A1(n10399), .A2(n10410), .ZN(P3_U3235) );
  INV_X1 U13133 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10411) );
  NOR2_X1 U13134 ( .A1(n10399), .A2(n10411), .ZN(P3_U3245) );
  NOR2_X1 U13135 ( .A1(n10423), .A2(n15907), .ZN(P3_U3246) );
  INV_X1 U13136 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10412) );
  NOR2_X1 U13137 ( .A1(n10399), .A2(n10412), .ZN(P3_U3260) );
  INV_X1 U13138 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10413) );
  NOR2_X1 U13139 ( .A1(n10423), .A2(n10413), .ZN(P3_U3261) );
  INV_X1 U13140 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10414) );
  NOR2_X1 U13141 ( .A1(n10423), .A2(n10414), .ZN(P3_U3247) );
  INV_X1 U13142 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10415) );
  NOR2_X1 U13143 ( .A1(n10423), .A2(n10415), .ZN(P3_U3263) );
  NOR2_X1 U13144 ( .A1(n10423), .A2(n15840), .ZN(P3_U3250) );
  INV_X1 U13145 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10416) );
  NOR2_X1 U13146 ( .A1(n10423), .A2(n10416), .ZN(P3_U3255) );
  INV_X1 U13147 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10417) );
  NOR2_X1 U13148 ( .A1(n10423), .A2(n10417), .ZN(P3_U3249) );
  INV_X1 U13149 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10418) );
  NOR2_X1 U13150 ( .A1(n10399), .A2(n10418), .ZN(P3_U3238) );
  INV_X1 U13151 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10419) );
  NOR2_X1 U13152 ( .A1(n10423), .A2(n10419), .ZN(P3_U3251) );
  INV_X1 U13153 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10420) );
  NOR2_X1 U13154 ( .A1(n10423), .A2(n10420), .ZN(P3_U3239) );
  INV_X1 U13155 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10421) );
  NOR2_X1 U13156 ( .A1(n10423), .A2(n10421), .ZN(P3_U3236) );
  INV_X1 U13157 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10422) );
  NOR2_X1 U13158 ( .A1(n10423), .A2(n10422), .ZN(P3_U3248) );
  INV_X1 U13159 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10424) );
  NOR2_X1 U13160 ( .A1(n10423), .A2(n10424), .ZN(P3_U3237) );
  INV_X1 U13161 ( .A(n10740), .ZN(n10733) );
  NOR2_X1 U13162 ( .A1(n10425), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14470) );
  INV_X2 U13163 ( .A(n14470), .ZN(n10996) );
  INV_X1 U13164 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10426) );
  NAND2_X1 U13165 ( .A1(n10425), .A2(P2_U3088), .ZN(n11492) );
  OAI222_X1 U13166 ( .A1(n10733), .A2(P2_U3088), .B1(n10996), .B2(n10427), 
        .C1(n10426), .C2(n11492), .ZN(P2_U3320) );
  INV_X1 U13167 ( .A(n11492), .ZN(n14473) );
  INV_X1 U13168 ( .A(n14473), .ZN(n14478) );
  OAI222_X1 U13169 ( .A1(P2_U3088), .A2(n7840), .B1(n10996), .B2(n10429), .C1(
        n10428), .C2(n14478), .ZN(P2_U3326) );
  INV_X1 U13170 ( .A(n10503), .ZN(n10718) );
  OAI222_X1 U13171 ( .A1(n10718), .A2(P2_U3088), .B1(n10996), .B2(n10431), 
        .C1(n10430), .C2(n14478), .ZN(P2_U3323) );
  INV_X1 U13172 ( .A(n10501), .ZN(n15525) );
  OAI222_X1 U13173 ( .A1(n15525), .A2(P2_U3088), .B1(n10996), .B2(n10433), 
        .C1(n10432), .C2(n14478), .ZN(P2_U3324) );
  INV_X1 U13174 ( .A(n10525), .ZN(n10533) );
  OAI222_X1 U13175 ( .A1(n10533), .A2(P2_U3088), .B1(n10996), .B2(n10435), 
        .C1(n10434), .C2(n14478), .ZN(P2_U3322) );
  INV_X1 U13176 ( .A(n10724), .ZN(n10514) );
  OAI222_X1 U13177 ( .A1(n10514), .A2(P2_U3088), .B1(n10996), .B2(n10437), 
        .C1(n10436), .C2(n14478), .ZN(P2_U3321) );
  OAI222_X1 U13178 ( .A1(P3_U3151), .A2(n10440), .B1(n12962), .B2(n10439), 
        .C1(n10438), .C2(n13550), .ZN(P3_U3283) );
  INV_X1 U13179 ( .A(n10441), .ZN(n10446) );
  AOI22_X1 U13180 ( .A1(n14750), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10442), .ZN(n10443) );
  OAI21_X1 U13181 ( .B1(n10446), .B2(n15236), .A(n10443), .ZN(P1_U3347) );
  INV_X1 U13182 ( .A(n10444), .ZN(n10453) );
  INV_X1 U13183 ( .A(n14768), .ZN(n10644) );
  OAI222_X1 U13184 ( .A1(n15236), .A2(n10453), .B1(n10644), .B2(P1_U3086), 
        .C1(n15797), .C2(n15232), .ZN(P1_U3344) );
  INV_X1 U13185 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10445) );
  OAI222_X1 U13186 ( .A1(n10934), .A2(P2_U3088), .B1(n10996), .B2(n10446), 
        .C1(n10445), .C2(n11492), .ZN(P2_U3319) );
  INV_X1 U13187 ( .A(n10447), .ZN(n10450) );
  INV_X1 U13188 ( .A(n10673), .ZN(n10681) );
  OAI222_X1 U13189 ( .A1(n15232), .A2(n10448), .B1(n15236), .B2(n10450), .C1(
        n6537), .C2(n10681), .ZN(P1_U3345) );
  INV_X1 U13190 ( .A(n15553), .ZN(n10451) );
  INV_X1 U13191 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10449) );
  OAI222_X1 U13192 ( .A1(n10451), .A2(P2_U3088), .B1(n10996), .B2(n10450), 
        .C1(n10449), .C2(n11492), .ZN(P2_U3317) );
  OAI222_X1 U13193 ( .A1(P2_U3088), .A2(n11105), .B1(n10996), .B2(n10453), 
        .C1(n10452), .C2(n11492), .ZN(P2_U3316) );
  INV_X1 U13194 ( .A(n10454), .ZN(n10456) );
  OAI222_X1 U13195 ( .A1(n15539), .A2(P2_U3088), .B1(n10996), .B2(n10456), 
        .C1(n10455), .C2(n11492), .ZN(P2_U3318) );
  INV_X1 U13196 ( .A(n10663), .ZN(n10641) );
  OAI222_X1 U13197 ( .A1(n15232), .A2(n10457), .B1(n15236), .B2(n10456), .C1(
        P1_U3086), .C2(n10641), .ZN(P1_U3346) );
  INV_X1 U13198 ( .A(n10458), .ZN(n10462) );
  INV_X1 U13199 ( .A(n10815), .ZN(n10618) );
  OAI222_X1 U13200 ( .A1(n15236), .A2(n10462), .B1(n10618), .B2(P1_U3086), 
        .C1(n10459), .C2(n15232), .ZN(P1_U3343) );
  INV_X1 U13201 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n15795) );
  NAND2_X1 U13202 ( .A1(n12207), .A2(P3_U3897), .ZN(n10460) );
  OAI21_X1 U13203 ( .B1(P3_U3897), .B2(n15795), .A(n10460), .ZN(P3_U3505) );
  INV_X1 U13204 ( .A(n11618), .ZN(n10463) );
  OAI222_X1 U13205 ( .A1(P2_U3088), .A2(n10463), .B1(n10996), .B2(n10462), 
        .C1(n10461), .C2(n11492), .ZN(P2_U3315) );
  INV_X1 U13206 ( .A(n10464), .ZN(n10478) );
  INV_X1 U13207 ( .A(n10855), .ZN(n10867) );
  OAI222_X1 U13208 ( .A1(n15236), .A2(n10478), .B1(n10867), .B2(n6537), .C1(
        n10465), .C2(n15232), .ZN(P1_U3342) );
  INV_X1 U13209 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n15821) );
  NAND2_X1 U13210 ( .A1(n13049), .A2(P3_U3897), .ZN(n10466) );
  OAI21_X1 U13211 ( .B1(P3_U3897), .B2(n15821), .A(n10466), .ZN(P3_U3507) );
  OR2_X1 U13212 ( .A1(n10468), .A2(n6537), .ZN(n12793) );
  NAND2_X1 U13213 ( .A1(n10467), .A2(n12793), .ZN(n10472) );
  NAND2_X1 U13214 ( .A1(n10468), .A2(n12721), .ZN(n10469) );
  AND2_X1 U13215 ( .A1(n10472), .A2(n10470), .ZN(n15342) );
  INV_X1 U13216 ( .A(n15342), .ZN(n14815) );
  INV_X1 U13217 ( .A(n10470), .ZN(n10471) );
  NAND2_X1 U13218 ( .A1(n10472), .A2(n10471), .ZN(n10617) );
  INV_X1 U13219 ( .A(n10617), .ZN(n10650) );
  INV_X1 U13220 ( .A(n15230), .ZN(n12969) );
  NAND2_X1 U13221 ( .A1(n12969), .A2(n8847), .ZN(n10473) );
  AND2_X1 U13222 ( .A1(n14664), .A2(n10473), .ZN(n14668) );
  OAI21_X1 U13223 ( .B1(n12969), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14668), .ZN(
        n10474) );
  XNOR2_X1 U13224 ( .A(n10474), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13225 ( .A1(n10650), .A2(n10475), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n6537), .ZN(n10476) );
  INV_X1 U13226 ( .A(n15566), .ZN(n10479) );
  OAI222_X1 U13227 ( .A1(P2_U3088), .A2(n10479), .B1(n10996), .B2(n10478), 
        .C1(n10477), .C2(n11492), .ZN(P2_U3314) );
  OAI222_X1 U13228 ( .A1(P3_U3151), .A2(n10482), .B1(n12962), .B2(n10481), 
        .C1(n10480), .C2(n13550), .ZN(P3_U3282) );
  NOR2_X1 U13229 ( .A1(n15342), .A2(n14666), .ZN(P1_U3085) );
  NAND2_X1 U13230 ( .A1(n10483), .A2(n11490), .ZN(n10484) );
  AND2_X1 U13231 ( .A1(n8048), .A2(n10484), .ZN(n10485) );
  AND2_X1 U13232 ( .A1(n10495), .A2(n10490), .ZN(n15498) );
  INV_X1 U13233 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n15952) );
  INV_X1 U13234 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10487) );
  INV_X1 U13235 ( .A(n15497), .ZN(n15502) );
  INV_X1 U13236 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n15661) );
  MUX2_X1 U13237 ( .A(n15661), .B(P2_REG1_REG_2__SCAN_IN), .S(n12536), .Z(
        n15519) );
  NOR2_X1 U13238 ( .A1(n6606), .A2(n15519), .ZN(n15518) );
  AOI21_X1 U13239 ( .B1(n12536), .B2(P2_REG1_REG_2__SCAN_IN), .A(n15518), .ZN(
        n15529) );
  INV_X1 U13240 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11264) );
  MUX2_X1 U13241 ( .A(n11264), .B(P2_REG1_REG_3__SCAN_IN), .S(n10501), .Z(
        n15530) );
  NOR2_X1 U13242 ( .A1(n15529), .A2(n15530), .ZN(n15528) );
  AOI21_X1 U13243 ( .B1(n10501), .B2(P2_REG1_REG_3__SCAN_IN), .A(n15528), .ZN(
        n10709) );
  INV_X1 U13244 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15663) );
  MUX2_X1 U13245 ( .A(n15663), .B(P2_REG1_REG_4__SCAN_IN), .S(n10503), .Z(
        n10710) );
  NOR2_X1 U13246 ( .A1(n10709), .A2(n10710), .ZN(n10708) );
  NOR2_X1 U13247 ( .A1(n10718), .A2(n15663), .ZN(n10526) );
  INV_X1 U13248 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10488) );
  MUX2_X1 U13249 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10488), .S(n10525), .Z(
        n10489) );
  NAND2_X1 U13250 ( .A1(n10525), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10493) );
  INV_X1 U13251 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15665) );
  MUX2_X1 U13252 ( .A(n15665), .B(P2_REG1_REG_6__SCAN_IN), .S(n10724), .Z(
        n10492) );
  NOR2_X1 U13253 ( .A1(n10490), .A2(P2_U3088), .ZN(n14472) );
  NAND2_X1 U13254 ( .A1(n10495), .A2(n14472), .ZN(n10507) );
  INV_X1 U13255 ( .A(n10507), .ZN(n10491) );
  NAND3_X1 U13256 ( .A1(n10529), .A2(n10493), .A3(n10492), .ZN(n10494) );
  NAND3_X1 U13257 ( .A1(n6727), .A2(n15596), .A3(n10494), .ZN(n10513) );
  INV_X1 U13258 ( .A(n15609), .ZN(n15527) );
  NAND2_X1 U13259 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10890) );
  INV_X1 U13260 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11526) );
  MUX2_X1 U13261 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11526), .S(n10724), .Z(
        n10509) );
  INV_X1 U13262 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10496) );
  MUX2_X1 U13263 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10496), .S(n12536), .Z(
        n15517) );
  INV_X1 U13264 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10497) );
  MUX2_X1 U13265 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10497), .S(n10498), .Z(
        n15506) );
  AND2_X1 U13266 ( .A1(n15497), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n15507) );
  NAND2_X1 U13267 ( .A1(n15506), .A2(n15507), .ZN(n15505) );
  NAND2_X1 U13268 ( .A1(n10498), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10499) );
  NAND2_X1 U13269 ( .A1(n15505), .A2(n10499), .ZN(n15516) );
  NAND2_X1 U13270 ( .A1(n12536), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10500) );
  NAND2_X1 U13271 ( .A1(n15515), .A2(n10500), .ZN(n15533) );
  INV_X1 U13272 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11565) );
  MUX2_X1 U13273 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11565), .S(n10501), .Z(
        n15534) );
  NAND2_X1 U13274 ( .A1(n15533), .A2(n15534), .ZN(n15532) );
  NAND2_X1 U13275 ( .A1(n10501), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10502) );
  NAND2_X1 U13276 ( .A1(n15532), .A2(n10502), .ZN(n10706) );
  INV_X1 U13277 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11603) );
  MUX2_X1 U13278 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11603), .S(n10503), .Z(
        n10707) );
  NAND2_X1 U13279 ( .A1(n10503), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U13280 ( .A1(n10705), .A2(n10521), .ZN(n10505) );
  INV_X1 U13281 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11581) );
  MUX2_X1 U13282 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11581), .S(n10525), .Z(
        n10504) );
  NAND2_X1 U13283 ( .A1(n10505), .A2(n10504), .ZN(n10523) );
  NAND2_X1 U13284 ( .A1(n10525), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U13285 ( .A1(n10523), .A2(n10506), .ZN(n10508) );
  OR2_X1 U13286 ( .A1(n10507), .A2(n13953), .ZN(n15579) );
  OAI211_X1 U13287 ( .C1(n10509), .C2(n10508), .A(n15603), .B(n10729), .ZN(
        n10510) );
  NAND2_X1 U13288 ( .A1(n10890), .A2(n10510), .ZN(n10511) );
  AOI21_X1 U13289 ( .B1(n15527), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n10511), .ZN(
        n10512) );
  OAI211_X1 U13290 ( .C1(n15584), .C2(n10514), .A(n10513), .B(n10512), .ZN(
        P2_U3220) );
  INV_X1 U13291 ( .A(n10568), .ZN(n10516) );
  AOI22_X1 U13292 ( .A1(n15407), .A2(n15985), .B1(n10516), .B2(n10515), .ZN(
        P1_U3445) );
  OAI222_X1 U13293 ( .A1(P3_U3151), .A2(n10518), .B1(n13550), .B2(n15956), 
        .C1(n12962), .C2(n10517), .ZN(P3_U3281) );
  NOR2_X1 U13294 ( .A1(n10519), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10800) );
  MUX2_X1 U13295 ( .A(n11581), .B(P2_REG2_REG_5__SCAN_IN), .S(n10525), .Z(
        n10520) );
  NAND3_X1 U13296 ( .A1(n10705), .A2(n10521), .A3(n10520), .ZN(n10522) );
  AND3_X1 U13297 ( .A1(n15603), .A2(n10523), .A3(n10522), .ZN(n10524) );
  AOI211_X1 U13298 ( .C1(n15527), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n10800), .B(
        n10524), .ZN(n10532) );
  MUX2_X1 U13299 ( .A(n10488), .B(P2_REG1_REG_5__SCAN_IN), .S(n10525), .Z(
        n10528) );
  INV_X1 U13300 ( .A(n10526), .ZN(n10527) );
  NAND2_X1 U13301 ( .A1(n10528), .A2(n10527), .ZN(n10530) );
  OAI211_X1 U13302 ( .C1(n10708), .C2(n10530), .A(n10529), .B(n15596), .ZN(
        n10531) );
  OAI211_X1 U13303 ( .C1(n15584), .C2(n10533), .A(n10532), .B(n10531), .ZN(
        P2_U3219) );
  INV_X1 U13304 ( .A(n10534), .ZN(n10535) );
  OAI222_X1 U13305 ( .A1(P3_U3151), .A2(n13221), .B1(n13550), .B2(n10536), 
        .C1(n12962), .C2(n10535), .ZN(P3_U3280) );
  INV_X1 U13306 ( .A(n10537), .ZN(n10538) );
  OAI21_X1 U13307 ( .B1(n13695), .B2(n10538), .A(n13725), .ZN(n10540) );
  OR2_X1 U13308 ( .A1(n10539), .A2(P2_U3088), .ZN(n13676) );
  AOI22_X1 U13309 ( .A1(n10540), .A2(n13756), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13676), .ZN(n10543) );
  NAND3_X1 U13310 ( .A1(n13712), .A2(n10541), .A3(n11233), .ZN(n10542) );
  OAI211_X1 U13311 ( .C1(n13744), .C2(n13718), .A(n10543), .B(n10542), .ZN(
        P2_U3204) );
  INV_X1 U13312 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n15798) );
  INV_X1 U13313 ( .A(n13413), .ZN(n10544) );
  NAND2_X1 U13314 ( .A1(n10544), .A2(P3_U3897), .ZN(n10545) );
  OAI21_X1 U13315 ( .B1(P3_U3897), .B2(n15798), .A(n10545), .ZN(P3_U3509) );
  NAND2_X1 U13316 ( .A1(n14666), .A2(n12041), .ZN(n10546) );
  OAI21_X1 U13317 ( .B1(n14666), .B2(n10547), .A(n10546), .ZN(P1_U3560) );
  INV_X1 U13318 ( .A(n10548), .ZN(n10549) );
  OAI222_X1 U13319 ( .A1(P3_U3151), .A2(n13237), .B1(n12962), .B2(n10549), 
        .C1(n15925), .C2(n13550), .ZN(P3_U3279) );
  OAI22_X1 U13320 ( .A1(n10551), .A2(P3_U3151), .B1(SI_17_), .B2(n13550), .ZN(
        n10552) );
  AOI21_X1 U13321 ( .B1(n10553), .B2(n11728), .A(n10552), .ZN(P3_U3278) );
  OAI22_X1 U13322 ( .A1(n15406), .A2(P1_D_REG_1__SCAN_IN), .B1(n10555), .B2(
        n10554), .ZN(n10556) );
  INV_X1 U13323 ( .A(n10556), .ZN(P1_U3446) );
  INV_X1 U13324 ( .A(n10557), .ZN(n10566) );
  INV_X1 U13325 ( .A(n11802), .ZN(n11459) );
  OAI222_X1 U13326 ( .A1(n15236), .A2(n10566), .B1(n11459), .B2(P1_U3086), 
        .C1(n10558), .C2(n15232), .ZN(P1_U3339) );
  INV_X1 U13327 ( .A(n13587), .ZN(n13722) );
  AOI22_X1 U13328 ( .A1(n13717), .A2(n8069), .B1(P2_STATE_REG_SCAN_IN), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n10560) );
  INV_X1 U13329 ( .A(n13767), .ZN(n13769) );
  OAI22_X1 U13330 ( .A1(n13769), .A2(n13725), .B1(n13718), .B2(n11256), .ZN(
        n10559) );
  AOI211_X1 U13331 ( .C1(n13722), .C2(n13980), .A(n10560), .B(n10559), .ZN(
        n10564) );
  OAI211_X1 U13332 ( .C1(n10562), .C2(n10561), .A(n10688), .B(n13711), .ZN(
        n10563) );
  NAND2_X1 U13333 ( .A1(n10564), .A2(n10563), .ZN(P2_U3190) );
  OAI222_X1 U13334 ( .A1(P2_U3088), .A2(n15585), .B1(n10996), .B2(n10566), 
        .C1(n10565), .C2(n14478), .ZN(P2_U3311) );
  INV_X1 U13335 ( .A(n10567), .ZN(n12790) );
  OAI21_X1 U13336 ( .B1(n10569), .B2(P1_D_REG_0__SCAN_IN), .A(n10568), .ZN(
        n10573) );
  INV_X1 U13337 ( .A(n10569), .ZN(n10571) );
  NAND2_X1 U13338 ( .A1(n10571), .A2(n10570), .ZN(n10572) );
  INV_X1 U13339 ( .A(n12038), .ZN(n11693) );
  INV_X1 U13340 ( .A(n10575), .ZN(n10583) );
  NAND2_X1 U13341 ( .A1(n14809), .A2(n15237), .ZN(n10577) );
  INV_X1 U13342 ( .A(n12558), .ZN(n12559) );
  NAND2_X1 U13343 ( .A1(n11695), .A2(n12559), .ZN(n10576) );
  INV_X1 U13344 ( .A(n12555), .ZN(n10578) );
  NAND2_X1 U13345 ( .A1(n10578), .A2(n12719), .ZN(n10579) );
  NAND2_X1 U13346 ( .A1(n10580), .A2(n10579), .ZN(n11668) );
  OR2_X1 U13347 ( .A1(n11668), .A2(n14809), .ZN(n15447) );
  NAND2_X1 U13348 ( .A1(n12720), .A2(n14809), .ZN(n15446) );
  NAND2_X1 U13349 ( .A1(n12041), .A2(n12038), .ZN(n12050) );
  OAI21_X1 U13350 ( .B1(n12041), .B2(n12038), .A(n12050), .ZN(n12750) );
  INV_X1 U13351 ( .A(n12750), .ZN(n10581) );
  OAI21_X1 U13352 ( .B1(n15389), .B2(n15476), .A(n10581), .ZN(n10582) );
  NAND2_X1 U13353 ( .A1(n11669), .A2(n15031), .ZN(n11880) );
  OAI211_X1 U13354 ( .C1(n11693), .C2(n10583), .A(n10582), .B(n11880), .ZN(
        n10780) );
  NAND2_X1 U13355 ( .A1(n15478), .A2(n10780), .ZN(n10584) );
  OAI21_X1 U13356 ( .B1(n15478), .B2(n8846), .A(n10584), .ZN(P1_U3459) );
  MUX2_X1 U13357 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10585), .S(n14691), .Z(
        n10590) );
  MUX2_X1 U13358 ( .A(n10586), .B(P1_REG2_REG_1__SCAN_IN), .S(n14656), .Z(
        n14651) );
  AND2_X1 U13359 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14663) );
  NAND2_X1 U13360 ( .A1(n14651), .A2(n14663), .ZN(n14670) );
  OR2_X1 U13361 ( .A1(n14656), .A2(n10586), .ZN(n14669) );
  NAND2_X1 U13362 ( .A1(n14670), .A2(n14669), .ZN(n10588) );
  NAND2_X1 U13363 ( .A1(n14676), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14687) );
  NAND2_X1 U13364 ( .A1(n10590), .A2(n10589), .ZN(n15335) );
  NAND2_X1 U13365 ( .A1(n14691), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n15334) );
  NAND2_X1 U13366 ( .A1(n15335), .A2(n15334), .ZN(n10593) );
  MUX2_X1 U13367 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10591), .S(n15339), .Z(
        n10592) );
  NAND2_X1 U13368 ( .A1(n15339), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14708) );
  NAND2_X1 U13369 ( .A1(n15337), .A2(n14708), .ZN(n10596) );
  MUX2_X1 U13370 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10594), .S(n14706), .Z(
        n10595) );
  NAND2_X1 U13371 ( .A1(n10596), .A2(n10595), .ZN(n14719) );
  NAND2_X1 U13372 ( .A1(n14706), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14718) );
  NAND2_X1 U13373 ( .A1(n14719), .A2(n14718), .ZN(n10599) );
  MUX2_X1 U13374 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10597), .S(n14716), .Z(
        n10598) );
  NAND2_X1 U13375 ( .A1(n14716), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14731) );
  NAND2_X1 U13376 ( .A1(n14732), .A2(n14731), .ZN(n10601) );
  MUX2_X1 U13377 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11692), .S(n14734), .Z(
        n10600) );
  NAND2_X1 U13378 ( .A1(n10601), .A2(n10600), .ZN(n14753) );
  NAND2_X1 U13379 ( .A1(n14734), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n14752) );
  NAND2_X1 U13380 ( .A1(n14753), .A2(n14752), .ZN(n10603) );
  MUX2_X1 U13381 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11711), .S(n14750), .Z(
        n10602) );
  NAND2_X1 U13382 ( .A1(n14750), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U13383 ( .A1(n14755), .A2(n10665), .ZN(n10605) );
  MUX2_X1 U13384 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11741), .S(n10663), .Z(
        n10604) );
  NAND2_X1 U13385 ( .A1(n10605), .A2(n10604), .ZN(n10676) );
  NAND2_X1 U13386 ( .A1(n10663), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10675) );
  NAND2_X1 U13387 ( .A1(n10676), .A2(n10675), .ZN(n10608) );
  MUX2_X1 U13388 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10606), .S(n10673), .Z(
        n10607) );
  NAND2_X1 U13389 ( .A1(n10673), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n14770) );
  NAND2_X1 U13390 ( .A1(n14771), .A2(n14770), .ZN(n10611) );
  MUX2_X1 U13391 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10609), .S(n14768), .Z(
        n10610) );
  NAND2_X1 U13392 ( .A1(n10611), .A2(n10610), .ZN(n14773) );
  NAND2_X1 U13393 ( .A1(n14768), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10612) );
  MUX2_X1 U13394 ( .A(n11944), .B(P1_REG2_REG_12__SCAN_IN), .S(n10815), .Z(
        n10614) );
  INV_X1 U13395 ( .A(n10811), .ZN(n10613) );
  AOI21_X1 U13396 ( .B1(n10615), .B2(n10614), .A(n10613), .ZN(n10654) );
  OR2_X1 U13397 ( .A1(n9335), .A2(n15230), .ZN(n10616) );
  NOR2_X1 U13398 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12030), .ZN(n10620) );
  NOR2_X1 U13399 ( .A1(n14804), .A2(n10618), .ZN(n10619) );
  AOI211_X1 U13400 ( .C1(n15342), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n10620), 
        .B(n10619), .ZN(n10653) );
  INV_X1 U13401 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10621) );
  XNOR2_X1 U13402 ( .A(n10815), .B(n10621), .ZN(n10649) );
  INV_X1 U13403 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10622) );
  MUX2_X1 U13404 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10622), .S(n14691), .Z(
        n10630) );
  INV_X1 U13405 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10623) );
  MUX2_X1 U13406 ( .A(n10623), .B(P1_REG1_REG_1__SCAN_IN), .S(n14656), .Z(
        n10625) );
  AND2_X1 U13407 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10624) );
  NAND2_X1 U13408 ( .A1(n10625), .A2(n10624), .ZN(n14678) );
  OR2_X1 U13409 ( .A1(n14656), .A2(n10623), .ZN(n14677) );
  NAND2_X1 U13410 ( .A1(n14678), .A2(n14677), .ZN(n10628) );
  INV_X1 U13411 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10626) );
  MUX2_X1 U13412 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10626), .S(n14676), .Z(
        n10627) );
  NAND2_X1 U13413 ( .A1(n10628), .A2(n10627), .ZN(n14693) );
  NAND2_X1 U13414 ( .A1(n14676), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14692) );
  NAND2_X1 U13415 ( .A1(n14693), .A2(n14692), .ZN(n10629) );
  NAND2_X1 U13416 ( .A1(n10630), .A2(n10629), .ZN(n15329) );
  NAND2_X1 U13417 ( .A1(n14691), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n15328) );
  NAND2_X1 U13418 ( .A1(n15329), .A2(n15328), .ZN(n10633) );
  INV_X1 U13419 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10631) );
  MUX2_X1 U13420 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10631), .S(n15339), .Z(
        n10632) );
  NAND2_X1 U13421 ( .A1(n10633), .A2(n10632), .ZN(n15331) );
  NAND2_X1 U13422 ( .A1(n15339), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10634) );
  AND2_X1 U13423 ( .A1(n15331), .A2(n10634), .ZN(n14704) );
  INV_X1 U13424 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15483) );
  MUX2_X1 U13425 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n15483), .S(n14706), .Z(
        n14703) );
  NAND2_X1 U13426 ( .A1(n14704), .A2(n14703), .ZN(n14702) );
  OR2_X1 U13427 ( .A1(n14706), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10635) );
  NAND2_X1 U13428 ( .A1(n14702), .A2(n10635), .ZN(n14722) );
  INV_X1 U13429 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15756) );
  MUX2_X1 U13430 ( .A(n15756), .B(P1_REG1_REG_6__SCAN_IN), .S(n14716), .Z(
        n14721) );
  OR2_X1 U13431 ( .A1(n14722), .A2(n14721), .ZN(n14737) );
  NAND2_X1 U13432 ( .A1(n14716), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n14736) );
  NAND2_X1 U13433 ( .A1(n14737), .A2(n14736), .ZN(n10638) );
  INV_X1 U13434 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10636) );
  MUX2_X1 U13435 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10636), .S(n14734), .Z(
        n10637) );
  NAND2_X1 U13436 ( .A1(n10638), .A2(n10637), .ZN(n14739) );
  NAND2_X1 U13437 ( .A1(n14734), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10639) );
  AND2_X1 U13438 ( .A1(n14739), .A2(n10639), .ZN(n14748) );
  INV_X1 U13439 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n15487) );
  MUX2_X1 U13440 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n15487), .S(n14750), .Z(
        n14747) );
  NAND2_X1 U13441 ( .A1(n14748), .A2(n14747), .ZN(n14746) );
  OR2_X1 U13442 ( .A1(n14750), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10658) );
  NAND2_X1 U13443 ( .A1(n14746), .A2(n10658), .ZN(n10640) );
  INV_X1 U13444 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15489) );
  MUX2_X1 U13445 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15489), .S(n10663), .Z(
        n10657) );
  NAND2_X1 U13446 ( .A1(n10640), .A2(n10657), .ZN(n10661) );
  NAND2_X1 U13447 ( .A1(n10641), .A2(n15489), .ZN(n10642) );
  NAND2_X1 U13448 ( .A1(n10661), .A2(n10642), .ZN(n10672) );
  INV_X1 U13449 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15943) );
  MUX2_X1 U13450 ( .A(n15943), .B(P1_REG1_REG_10__SCAN_IN), .S(n10673), .Z(
        n10671) );
  NAND2_X1 U13451 ( .A1(n10673), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n14761) );
  INV_X1 U13452 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10643) );
  NAND2_X1 U13453 ( .A1(n10644), .A2(n10643), .ZN(n10647) );
  NAND2_X1 U13454 ( .A1(n14768), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10645) );
  AND2_X1 U13455 ( .A1(n10647), .A2(n10645), .ZN(n14760) );
  AND2_X1 U13456 ( .A1(n14761), .A2(n14760), .ZN(n10646) );
  NAND2_X1 U13457 ( .A1(n14762), .A2(n10646), .ZN(n14759) );
  NAND2_X1 U13458 ( .A1(n14759), .A2(n10647), .ZN(n10648) );
  NAND2_X1 U13459 ( .A1(n10648), .A2(n10649), .ZN(n10817) );
  OAI21_X1 U13460 ( .B1(n10649), .B2(n10648), .A(n10817), .ZN(n10651) );
  NAND2_X1 U13461 ( .A1(n10651), .A2(n15332), .ZN(n10652) );
  OAI211_X1 U13462 ( .C1(n10654), .C2(n14805), .A(n10653), .B(n10652), .ZN(
        P1_U3255) );
  INV_X1 U13463 ( .A(n10655), .ZN(n10685) );
  INV_X1 U13464 ( .A(n11335), .ZN(n11329) );
  OAI222_X1 U13465 ( .A1(n15236), .A2(n10685), .B1(n11329), .B2(n6537), .C1(
        n10656), .C2(n15232), .ZN(P1_U3341) );
  INV_X1 U13466 ( .A(n10657), .ZN(n10659) );
  NAND3_X1 U13467 ( .A1(n14746), .A2(n10659), .A3(n10658), .ZN(n10660) );
  AND2_X1 U13468 ( .A1(n10661), .A2(n10660), .ZN(n10669) );
  INV_X1 U13469 ( .A(n15332), .ZN(n11347) );
  AND2_X1 U13470 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n11919) );
  INV_X1 U13471 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n11757) );
  NOR2_X1 U13472 ( .A1(n14815), .A2(n11757), .ZN(n10662) );
  AOI211_X1 U13473 ( .C1(n15340), .C2(n10663), .A(n11919), .B(n10662), .ZN(
        n10668) );
  MUX2_X1 U13474 ( .A(n11741), .B(P1_REG2_REG_9__SCAN_IN), .S(n10663), .Z(
        n10664) );
  NAND3_X1 U13475 ( .A1(n14755), .A2(n10665), .A3(n10664), .ZN(n10666) );
  NAND3_X1 U13476 ( .A1(n15338), .A2(n10676), .A3(n10666), .ZN(n10667) );
  OAI211_X1 U13477 ( .C1(n10669), .C2(n11347), .A(n10668), .B(n10667), .ZN(
        P1_U3252) );
  INV_X1 U13478 ( .A(n14762), .ZN(n10670) );
  AOI211_X1 U13479 ( .C1(n10672), .C2(n10671), .A(n11347), .B(n10670), .ZN(
        n10683) );
  MUX2_X1 U13480 ( .A(n10606), .B(P1_REG2_REG_10__SCAN_IN), .S(n10673), .Z(
        n10674) );
  NAND3_X1 U13481 ( .A1(n10676), .A2(n10675), .A3(n10674), .ZN(n10677) );
  NAND3_X1 U13482 ( .A1(n15338), .A2(n14771), .A3(n10677), .ZN(n10680) );
  NOR2_X1 U13483 ( .A1(n10678), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11895) );
  AOI21_X1 U13484 ( .B1(n15342), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11895), 
        .ZN(n10679) );
  OAI211_X1 U13485 ( .C1(n14804), .C2(n10681), .A(n10680), .B(n10679), .ZN(
        n10682) );
  OR2_X1 U13486 ( .A1(n10683), .A2(n10682), .ZN(P1_U3253) );
  INV_X1 U13487 ( .A(n12157), .ZN(n12161) );
  OAI222_X1 U13488 ( .A1(P2_U3088), .A2(n12161), .B1(n10996), .B2(n10685), 
        .C1(n10684), .C2(n14478), .ZN(P2_U3313) );
  INV_X1 U13489 ( .A(n10686), .ZN(n10702) );
  INV_X1 U13490 ( .A(n14781), .ZN(n11810) );
  OAI222_X1 U13491 ( .A1(n15236), .A2(n10702), .B1(n11810), .B2(n6537), .C1(
        n10687), .C2(n15232), .ZN(P1_U3338) );
  INV_X1 U13492 ( .A(n10688), .ZN(n10691) );
  INV_X1 U13493 ( .A(n10695), .ZN(n10690) );
  INV_X1 U13494 ( .A(n10689), .ZN(n10805) );
  AOI21_X1 U13495 ( .B1(n10691), .B2(n10690), .A(n10805), .ZN(n10700) );
  INV_X1 U13496 ( .A(n13718), .ZN(n13675) );
  NAND2_X1 U13497 ( .A1(n13675), .A2(n13977), .ZN(n10692) );
  NAND2_X1 U13498 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10714) );
  OAI211_X1 U13499 ( .C1(n13733), .C2(n13725), .A(n10692), .B(n10714), .ZN(
        n10693) );
  AOI21_X1 U13500 ( .B1(n10694), .B2(n13701), .A(n10693), .ZN(n10699) );
  INV_X1 U13501 ( .A(n13712), .ZN(n13697) );
  NOR3_X1 U13502 ( .A1(n13697), .A2(n10696), .A3(n10695), .ZN(n10697) );
  OAI21_X1 U13503 ( .B1(n10697), .B2(n13722), .A(n13979), .ZN(n10698) );
  OAI211_X1 U13504 ( .C1(n10700), .C2(n13695), .A(n10699), .B(n10698), .ZN(
        P2_U3202) );
  INV_X1 U13505 ( .A(n15598), .ZN(n10703) );
  OAI222_X1 U13506 ( .A1(P2_U3088), .A2(n10703), .B1(n10996), .B2(n10702), 
        .C1(n10701), .C2(n14478), .ZN(P2_U3310) );
  INV_X1 U13507 ( .A(n10704), .ZN(n10737) );
  INV_X1 U13508 ( .A(n11344), .ZN(n11448) );
  OAI222_X1 U13509 ( .A1(n15236), .A2(n10737), .B1(n11448), .B2(P1_U3086), 
        .C1(n15737), .C2(n15232), .ZN(P1_U3340) );
  OAI211_X1 U13510 ( .C1(n10707), .C2(n10706), .A(n15603), .B(n10705), .ZN(
        n10713) );
  AOI211_X1 U13511 ( .C1(n10710), .C2(n10709), .A(n10708), .B(n15586), .ZN(
        n10711) );
  INV_X1 U13512 ( .A(n10711), .ZN(n10712) );
  NAND2_X1 U13513 ( .A1(n10713), .A2(n10712), .ZN(n10716) );
  INV_X1 U13514 ( .A(n10714), .ZN(n10715) );
  AOI211_X1 U13515 ( .C1(n15527), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n10716), .B(
        n10715), .ZN(n10717) );
  OAI21_X1 U13516 ( .B1(n15584), .B2(n10718), .A(n10717), .ZN(P2_U3218) );
  NAND2_X1 U13517 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n10986) );
  INV_X1 U13518 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15668) );
  MUX2_X1 U13519 ( .A(n15668), .B(P2_REG1_REG_7__SCAN_IN), .S(n10740), .Z(
        n10720) );
  AOI211_X1 U13520 ( .C1(n10720), .C2(n10719), .A(n10738), .B(n15586), .ZN(
        n10721) );
  INV_X1 U13521 ( .A(n10721), .ZN(n10722) );
  NAND2_X1 U13522 ( .A1(n10986), .A2(n10722), .ZN(n10723) );
  AOI21_X1 U13523 ( .B1(n15527), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n10723), .ZN(
        n10732) );
  NAND2_X1 U13524 ( .A1(n10724), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10728) );
  NAND2_X1 U13525 ( .A1(n10729), .A2(n10728), .ZN(n10726) );
  INV_X1 U13526 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11542) );
  MUX2_X1 U13527 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11542), .S(n10740), .Z(
        n10725) );
  NAND2_X1 U13528 ( .A1(n10726), .A2(n10725), .ZN(n10742) );
  MUX2_X1 U13529 ( .A(n11542), .B(P2_REG2_REG_7__SCAN_IN), .S(n10740), .Z(
        n10727) );
  NAND3_X1 U13530 ( .A1(n10729), .A2(n10728), .A3(n10727), .ZN(n10730) );
  NAND3_X1 U13531 ( .A1(n15603), .A2(n10742), .A3(n10730), .ZN(n10731) );
  OAI211_X1 U13532 ( .C1(n15584), .C2(n10733), .A(n10732), .B(n10731), .ZN(
        P2_U3221) );
  OAI222_X1 U13533 ( .A1(P3_U3151), .A2(n6810), .B1(n13550), .B2(n10735), .C1(
        n12962), .C2(n10734), .ZN(P3_U3277) );
  INV_X1 U13534 ( .A(n13998), .ZN(n12166) );
  OAI222_X1 U13535 ( .A1(P2_U3088), .A2(n12166), .B1(n10996), .B2(n10737), 
        .C1(n10736), .C2(n14478), .ZN(P2_U3312) );
  AOI21_X1 U13536 ( .B1(n10740), .B2(P2_REG1_REG_7__SCAN_IN), .A(n10738), .ZN(
        n10936) );
  INV_X1 U13537 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10933) );
  XNOR2_X1 U13538 ( .A(n10934), .B(n10933), .ZN(n10935) );
  XOR2_X1 U13539 ( .A(n10936), .B(n10935), .Z(n10739) );
  NAND2_X1 U13540 ( .A1(n15596), .A2(n10739), .ZN(n10746) );
  INV_X1 U13541 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11556) );
  MUX2_X1 U13542 ( .A(n11556), .B(P2_REG2_REG_8__SCAN_IN), .S(n10934), .Z(
        n10744) );
  NAND2_X1 U13543 ( .A1(n10740), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10741) );
  NAND2_X1 U13544 ( .A1(n10742), .A2(n10741), .ZN(n10743) );
  OAI211_X1 U13545 ( .C1(n10744), .C2(n10743), .A(n15603), .B(n10940), .ZN(
        n10745) );
  NAND2_X1 U13546 ( .A1(n10746), .A2(n10745), .ZN(n10748) );
  NAND2_X1 U13547 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11195) );
  INV_X1 U13548 ( .A(n11195), .ZN(n10747) );
  AOI211_X1 U13549 ( .C1(n15527), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10748), .B(
        n10747), .ZN(n10749) );
  OAI21_X1 U13550 ( .B1(n15584), .B2(n10934), .A(n10749), .ZN(P2_U3222) );
  INV_X1 U13551 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14700) );
  NAND2_X1 U13552 ( .A1(n10753), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10754) );
  XNOR2_X1 U13553 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n10755) );
  XNOR2_X1 U13554 ( .A(n10762), .B(n10755), .ZN(n15245) );
  INV_X1 U13555 ( .A(n10756), .ZN(n10757) );
  NAND2_X1 U13556 ( .A1(n10757), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10758) );
  INV_X1 U13557 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10760) );
  INV_X1 U13558 ( .A(n10767), .ZN(n10763) );
  XNOR2_X1 U13559 ( .A(n10763), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15247) );
  NAND2_X1 U13560 ( .A1(n15248), .A2(n15247), .ZN(n10766) );
  NAND2_X1 U13561 ( .A1(n10764), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10765) );
  NAND2_X1 U13562 ( .A1(n10766), .A2(n10765), .ZN(n10773) );
  NAND2_X1 U13563 ( .A1(n10767), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10770) );
  INV_X1 U13564 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15897) );
  NAND2_X1 U13565 ( .A1(n10768), .A2(n15897), .ZN(n10769) );
  NAND2_X1 U13566 ( .A1(n10770), .A2(n10769), .ZN(n11022) );
  XNOR2_X1 U13567 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n11021) );
  INV_X1 U13568 ( .A(n11021), .ZN(n10771) );
  XNOR2_X1 U13569 ( .A(n11022), .B(n10771), .ZN(n10772) );
  NAND2_X1 U13570 ( .A1(n10775), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U13571 ( .A1(n11020), .A2(n10776), .ZN(SUB_1596_U55) );
  INV_X1 U13572 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14654) );
  NAND2_X1 U13573 ( .A1(n15492), .A2(n10780), .ZN(n10781) );
  OAI21_X1 U13574 ( .B1(n15492), .B2(n14654), .A(n10781), .ZN(P1_U3528) );
  AOI21_X1 U13575 ( .B1(n10783), .B2(n6722), .A(n10782), .ZN(n10797) );
  OAI21_X1 U13576 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10784), .A(n10920), .ZN(
        n10788) );
  AND2_X1 U13577 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11647) );
  AOI21_X1 U13578 ( .B1(n15694), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11647), .ZN(
        n10785) );
  OAI21_X1 U13579 ( .B1(n13261), .B2(n10786), .A(n10785), .ZN(n10787) );
  AOI21_X1 U13580 ( .B1(n10788), .B2(n13284), .A(n10787), .ZN(n10796) );
  INV_X1 U13581 ( .A(n10789), .ZN(n13149) );
  INV_X1 U13582 ( .A(n10790), .ZN(n10792) );
  NOR3_X1 U13583 ( .A1(n13149), .A2(n10792), .A3(n10791), .ZN(n10794) );
  INV_X1 U13584 ( .A(n10913), .ZN(n10793) );
  OAI21_X1 U13585 ( .B1(n10794), .B2(n10793), .A(n13248), .ZN(n10795) );
  OAI211_X1 U13586 ( .C1(n10797), .C2(n13288), .A(n10796), .B(n10795), .ZN(
        P3_U3189) );
  OAI222_X1 U13587 ( .A1(P3_U3151), .A2(n12526), .B1(n12962), .B2(n10799), 
        .C1(n10798), .C2(n13550), .ZN(P3_U3276) );
  INV_X1 U13588 ( .A(n13703), .ZN(n13666) );
  OAI22_X1 U13589 ( .A1(n11256), .A2(n14116), .B1(n13776), .B2(n14118), .ZN(
        n11079) );
  AOI21_X1 U13590 ( .B1(n13666), .B2(n11079), .A(n10800), .ZN(n10801) );
  OAI21_X1 U13591 ( .B1(n13727), .B2(n13725), .A(n10801), .ZN(n10807) );
  AOI22_X1 U13592 ( .A1(n13712), .A2(n13978), .B1(n13711), .B2(n10802), .ZN(
        n10804) );
  NOR3_X1 U13593 ( .A1(n10805), .A2(n10804), .A3(n10803), .ZN(n10806) );
  AOI211_X1 U13594 ( .C1(n13701), .C2(n11582), .A(n10807), .B(n10806), .ZN(
        n10808) );
  OAI21_X1 U13595 ( .B1(n13695), .B2(n10809), .A(n10808), .ZN(P2_U3199) );
  OR2_X1 U13596 ( .A1(n10815), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10810) );
  MUX2_X1 U13597 ( .A(n12114), .B(P1_REG2_REG_13__SCAN_IN), .S(n10855), .Z(
        n10812) );
  NAND2_X1 U13598 ( .A1(n10855), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10813) );
  NAND2_X1 U13599 ( .A1(n10856), .A2(n10813), .ZN(n11334) );
  XNOR2_X1 U13600 ( .A(n11335), .B(n10814), .ZN(n11333) );
  XNOR2_X1 U13601 ( .A(n11334), .B(n11333), .ZN(n10826) );
  OR2_X1 U13602 ( .A1(n10815), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10816) );
  NAND2_X1 U13603 ( .A1(n10817), .A2(n10816), .ZN(n10859) );
  XNOR2_X1 U13604 ( .A(n10855), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10860) );
  INV_X1 U13605 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11328) );
  XNOR2_X1 U13606 ( .A(n11335), .B(n11328), .ZN(n10819) );
  NAND2_X1 U13607 ( .A1(n10855), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10820) );
  AND2_X1 U13608 ( .A1(n10819), .A2(n10820), .ZN(n10818) );
  NAND2_X1 U13609 ( .A1(n10861), .A2(n10818), .ZN(n11331) );
  INV_X1 U13610 ( .A(n11331), .ZN(n10822) );
  AOI21_X1 U13611 ( .B1(n10861), .B2(n10820), .A(n10819), .ZN(n10821) );
  OAI21_X1 U13612 ( .B1(n10822), .B2(n10821), .A(n15332), .ZN(n10825) );
  INV_X1 U13613 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15277) );
  NAND2_X1 U13614 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14494)
         );
  OAI21_X1 U13615 ( .B1(n14815), .B2(n15277), .A(n14494), .ZN(n10823) );
  AOI21_X1 U13616 ( .B1(n11335), .B2(n15340), .A(n10823), .ZN(n10824) );
  OAI211_X1 U13617 ( .C1(n10826), .C2(n14805), .A(n10825), .B(n10824), .ZN(
        P1_U3257) );
  OAI21_X1 U13618 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n10828), .A(n10827), .ZN(
        n10839) );
  INV_X1 U13619 ( .A(n15694), .ZN(n13273) );
  OAI21_X1 U13620 ( .B1(n10829), .B2(n11180), .A(n10874), .ZN(n10830) );
  AOI22_X1 U13621 ( .A1(n10830), .A2(n13248), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10831) );
  OAI21_X1 U13622 ( .B1(n13273), .B2(n10832), .A(n10831), .ZN(n10838) );
  AOI21_X1 U13623 ( .B1(n15687), .B2(n10834), .A(n10833), .ZN(n10835) );
  OAI22_X1 U13624 ( .A1(n13261), .A2(n10836), .B1(n10835), .B2(n13288), .ZN(
        n10837) );
  AOI211_X1 U13625 ( .C1(n13284), .C2(n10839), .A(n10838), .B(n10837), .ZN(
        n10840) );
  INV_X1 U13626 ( .A(n10840), .ZN(P3_U3183) );
  NOR2_X1 U13627 ( .A1(n10842), .A2(n6831), .ZN(n10844) );
  INV_X1 U13628 ( .A(n10843), .ZN(n13148) );
  AOI21_X1 U13629 ( .B1(n10844), .B2(n10961), .A(n13148), .ZN(n10853) );
  OAI21_X1 U13630 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n10845), .A(n13140), .ZN(
        n10848) );
  INV_X1 U13631 ( .A(n13288), .ZN(n13209) );
  OAI21_X1 U13632 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n10846), .A(n13153), .ZN(
        n10847) );
  AOI22_X1 U13633 ( .A1(n10848), .A2(n13209), .B1(n13284), .B2(n10847), .ZN(
        n10852) );
  AND2_X1 U13634 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11634) );
  NOR2_X1 U13635 ( .A1(n13261), .A2(n10849), .ZN(n10850) );
  AOI211_X1 U13636 ( .C1(n15694), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n11634), .B(
        n10850), .ZN(n10851) );
  OAI211_X1 U13637 ( .C1(n10853), .C2(n13277), .A(n10852), .B(n10851), .ZN(
        P3_U3187) );
  INV_X1 U13638 ( .A(n10854), .ZN(n10858) );
  MUX2_X1 U13639 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n12114), .S(n10855), .Z(
        n10857) );
  OAI211_X1 U13640 ( .C1(n10858), .C2(n10857), .A(n15338), .B(n10856), .ZN(
        n10866) );
  NAND2_X1 U13641 ( .A1(n6537), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12174) );
  AOI21_X1 U13642 ( .B1(n10860), .B2(n10859), .A(n11347), .ZN(n10862) );
  NAND2_X1 U13643 ( .A1(n10862), .A2(n10861), .ZN(n10863) );
  NAND2_X1 U13644 ( .A1(n12174), .A2(n10863), .ZN(n10864) );
  AOI21_X1 U13645 ( .B1(n15342), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10864), 
        .ZN(n10865) );
  OAI211_X1 U13646 ( .C1(n14804), .C2(n10867), .A(n10866), .B(n10865), .ZN(
        P1_U3256) );
  AOI21_X1 U13647 ( .B1(n10870), .B2(n10869), .A(n10868), .ZN(n10885) );
  INV_X1 U13648 ( .A(n10871), .ZN(n10873) );
  NAND3_X1 U13649 ( .A1(n10874), .A2(n10873), .A3(n10872), .ZN(n10875) );
  AOI21_X1 U13650 ( .B1(n13123), .B2(n10875), .A(n13277), .ZN(n10877) );
  INV_X1 U13651 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11408) );
  OAI22_X1 U13652 ( .A1(n13273), .A2(n15696), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11408), .ZN(n10876) );
  AOI211_X1 U13653 ( .C1(n10878), .C2(n13279), .A(n10877), .B(n10876), .ZN(
        n10884) );
  OAI21_X1 U13654 ( .B1(n10881), .B2(n10880), .A(n10879), .ZN(n10882) );
  NAND2_X1 U13655 ( .A1(n13284), .A2(n10882), .ZN(n10883) );
  OAI211_X1 U13656 ( .C1(n10885), .C2(n13288), .A(n10884), .B(n10883), .ZN(
        P3_U3184) );
  INV_X1 U13657 ( .A(n10886), .ZN(n11530) );
  AOI21_X1 U13658 ( .B1(n10888), .B2(n10887), .A(n13695), .ZN(n10889) );
  NAND2_X1 U13659 ( .A1(n10889), .A2(n10981), .ZN(n10893) );
  AOI22_X1 U13660 ( .A1(n13975), .A2(n14304), .B1(n14302), .B2(n13977), .ZN(
        n11524) );
  OAI21_X1 U13661 ( .B1(n13703), .B2(n11524), .A(n10890), .ZN(n10891) );
  AOI21_X1 U13662 ( .B1(n13693), .B2(n13777), .A(n10891), .ZN(n10892) );
  OAI211_X1 U13663 ( .C1(n13717), .C2(n11530), .A(n10893), .B(n10892), .ZN(
        P2_U3211) );
  NAND2_X1 U13664 ( .A1(n13606), .A2(n13904), .ZN(n10894) );
  NAND2_X1 U13665 ( .A1(n11076), .A2(n10894), .ZN(n12306) );
  NAND2_X1 U13666 ( .A1(n13745), .A2(n13756), .ZN(n10895) );
  NAND2_X1 U13667 ( .A1(n10895), .A2(n14239), .ZN(n10896) );
  NOR2_X1 U13668 ( .A1(n12011), .A2(n10896), .ZN(n12308) );
  INV_X1 U13669 ( .A(n15642), .ZN(n11601) );
  NAND2_X1 U13670 ( .A1(n12306), .A2(n11601), .ZN(n10902) );
  OAI21_X1 U13671 ( .B1(n10898), .B2(n13904), .A(n10897), .ZN(n10899) );
  NAND2_X1 U13672 ( .A1(n10899), .A2(n14307), .ZN(n10901) );
  AOI22_X1 U13673 ( .A1(n10541), .A2(n14302), .B1(n14304), .B2(n13980), .ZN(
        n10900) );
  NAND3_X1 U13674 ( .A1(n10902), .A2(n10901), .A3(n10900), .ZN(n12305) );
  AOI211_X1 U13675 ( .C1(n15646), .C2(n12306), .A(n12308), .B(n12305), .ZN(
        n10908) );
  INV_X1 U13676 ( .A(n13745), .ZN(n13742) );
  OAI22_X1 U13677 ( .A1(n14400), .A2(n13742), .B1(n15670), .B2(n15952), .ZN(
        n10903) );
  INV_X1 U13678 ( .A(n10903), .ZN(n10904) );
  OAI21_X1 U13679 ( .B1(n10908), .B2(n15667), .A(n10904), .ZN(P2_U3500) );
  INV_X1 U13680 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10905) );
  OAI22_X1 U13681 ( .A1(n14459), .A2(n13742), .B1(n15659), .B2(n10905), .ZN(
        n10906) );
  INV_X1 U13682 ( .A(n10906), .ZN(n10907) );
  OAI21_X1 U13683 ( .B1(n10908), .B2(n15657), .A(n10907), .ZN(P2_U3433) );
  INV_X1 U13684 ( .A(n10909), .ZN(n10910) );
  NOR2_X1 U13685 ( .A1(n10911), .A2(n10910), .ZN(n10914) );
  INV_X1 U13686 ( .A(n11305), .ZN(n10912) );
  AOI21_X1 U13687 ( .B1(n10914), .B2(n10913), .A(n10912), .ZN(n10927) );
  NOR3_X1 U13688 ( .A1(n10782), .A2(n10916), .A3(n10915), .ZN(n10917) );
  OAI21_X1 U13689 ( .B1(n6721), .B2(n10917), .A(n13209), .ZN(n10926) );
  INV_X1 U13690 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U13691 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11815) );
  OAI21_X1 U13692 ( .B1(n13273), .B2(n11023), .A(n11815), .ZN(n10923) );
  NAND3_X1 U13693 ( .A1(n10920), .A2(n10919), .A3(n10918), .ZN(n10921) );
  AOI21_X1 U13694 ( .B1(n6725), .B2(n10921), .A(n13242), .ZN(n10922) );
  AOI211_X1 U13695 ( .C1(n10924), .C2(n13279), .A(n10923), .B(n10922), .ZN(
        n10925) );
  OAI211_X1 U13696 ( .C1(n10927), .C2(n13277), .A(n10926), .B(n10925), .ZN(
        P3_U3190) );
  NAND2_X1 U13697 ( .A1(n10928), .A2(n13428), .ZN(n10929) );
  INV_X1 U13698 ( .A(n10930), .ZN(n11460) );
  AND2_X1 U13699 ( .A1(n11460), .A2(n13118), .ZN(n12364) );
  OR2_X1 U13700 ( .A1(n12364), .A2(n12365), .ZN(n12484) );
  AOI22_X1 U13701 ( .A1(n10929), .A2(n12484), .B1(n13396), .B2(n7138), .ZN(
        n10955) );
  MUX2_X1 U13702 ( .A(n10955), .B(n11174), .S(n15688), .Z(n10932) );
  AOI22_X1 U13703 ( .A1(n13438), .A2(n10930), .B1(n15675), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10931) );
  NAND2_X1 U13704 ( .A1(n10932), .A2(n10931), .ZN(P3_U3233) );
  XOR2_X1 U13705 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n15539), .Z(n15543) );
  INV_X1 U13706 ( .A(n15539), .ZN(n15546) );
  XNOR2_X1 U13707 ( .A(n15553), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n15556) );
  XNOR2_X1 U13708 ( .A(n10943), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n11106) );
  XNOR2_X1 U13709 ( .A(n11107), .B(n11106), .ZN(n10952) );
  AND2_X1 U13710 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11780) );
  INV_X1 U13711 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n12094) );
  NOR2_X1 U13712 ( .A1(n15609), .A2(n12094), .ZN(n10937) );
  AOI211_X1 U13713 ( .C1(n15595), .C2(n10943), .A(n11780), .B(n10937), .ZN(
        n10951) );
  INV_X1 U13714 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11870) );
  MUX2_X1 U13715 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11870), .S(n15539), .Z(
        n10941) );
  NAND2_X1 U13716 ( .A1(n10938), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10939) );
  NAND2_X1 U13717 ( .A1(n10940), .A2(n10939), .ZN(n15538) );
  OR2_X2 U13718 ( .A1(n10941), .A2(n15538), .ZN(n15540) );
  NAND2_X1 U13719 ( .A1(n15539), .A2(n11870), .ZN(n10942) );
  INV_X1 U13720 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11960) );
  MUX2_X1 U13721 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n11960), .S(n15553), .Z(
        n15559) );
  NAND2_X1 U13722 ( .A1(n15553), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10947) );
  NAND2_X1 U13723 ( .A1(n10943), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10944) );
  INV_X1 U13724 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n14292) );
  NAND2_X1 U13725 ( .A1(n11105), .A2(n14292), .ZN(n11111) );
  AND2_X1 U13726 ( .A1(n10944), .A2(n11111), .ZN(n10946) );
  AND2_X1 U13727 ( .A1(n10947), .A2(n10946), .ZN(n10945) );
  NAND2_X1 U13728 ( .A1(n15558), .A2(n10945), .ZN(n11113) );
  INV_X1 U13729 ( .A(n11113), .ZN(n10949) );
  AOI21_X1 U13730 ( .B1(n15558), .B2(n10947), .A(n10946), .ZN(n10948) );
  OAI21_X1 U13731 ( .B1(n10949), .B2(n10948), .A(n15603), .ZN(n10950) );
  OAI211_X1 U13732 ( .C1(n10952), .C2(n15586), .A(n10951), .B(n10950), .ZN(
        P2_U3225) );
  INV_X1 U13733 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10953) );
  MUX2_X1 U13734 ( .A(n10955), .B(n10953), .S(n15693), .Z(n10954) );
  OAI21_X1 U13735 ( .B1(n11460), .B2(n13536), .A(n10954), .ZN(P3_U3390) );
  MUX2_X1 U13736 ( .A(n10956), .B(n10955), .S(n13486), .Z(n10957) );
  OAI21_X1 U13737 ( .B1(n11460), .B2(n13482), .A(n10957), .ZN(P3_U3459) );
  INV_X1 U13738 ( .A(n10958), .ZN(n10959) );
  NOR2_X1 U13739 ( .A1(n10960), .A2(n10959), .ZN(n10963) );
  INV_X1 U13740 ( .A(n10961), .ZN(n10962) );
  AOI21_X1 U13741 ( .B1(n10963), .B2(n13128), .A(n10962), .ZN(n10978) );
  INV_X1 U13742 ( .A(n10964), .ZN(n10968) );
  NAND3_X1 U13743 ( .A1(n13119), .A2(n10966), .A3(n10965), .ZN(n10967) );
  AOI21_X1 U13744 ( .B1(n10968), .B2(n10967), .A(n13288), .ZN(n10976) );
  AND3_X1 U13745 ( .A1(n13131), .A2(n10971), .A3(n10970), .ZN(n10972) );
  OAI21_X1 U13746 ( .B1(n10969), .B2(n10972), .A(n13284), .ZN(n10973) );
  NAND2_X1 U13747 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11508) );
  OAI211_X1 U13748 ( .C1(n13273), .C2(n10974), .A(n10973), .B(n11508), .ZN(
        n10975) );
  AOI211_X1 U13749 ( .C1(n9411), .C2(n13279), .A(n10976), .B(n10975), .ZN(
        n10977) );
  OAI21_X1 U13750 ( .B1(n10978), .B2(n13277), .A(n10977), .ZN(P3_U3186) );
  INV_X1 U13751 ( .A(n10979), .ZN(n10980) );
  AOI21_X1 U13752 ( .B1(n10981), .B2(n10980), .A(n13695), .ZN(n10985) );
  NOR3_X1 U13753 ( .A1(n13697), .A2(n13776), .A3(n10982), .ZN(n10984) );
  OAI21_X1 U13754 ( .B1(n10985), .B2(n10984), .A(n10983), .ZN(n10992) );
  OAI21_X1 U13755 ( .B1(n13718), .B2(n10987), .A(n10986), .ZN(n10990) );
  INV_X1 U13756 ( .A(n10988), .ZN(n11545) );
  OAI22_X1 U13757 ( .A1(n13776), .A2(n13587), .B1(n13717), .B2(n11545), .ZN(
        n10989) );
  AOI211_X1 U13758 ( .C1(n15650), .C2(n13693), .A(n10990), .B(n10989), .ZN(
        n10991) );
  NAND2_X1 U13759 ( .A1(n10992), .A2(n10991), .ZN(P2_U3185) );
  INV_X1 U13760 ( .A(n10993), .ZN(n10995) );
  INV_X1 U13761 ( .A(n14798), .ZN(n14787) );
  OAI222_X1 U13762 ( .A1(n15232), .A2(n10994), .B1(n15236), .B2(n10995), .C1(
        n6537), .C2(n14787), .ZN(P1_U3337) );
  INV_X1 U13763 ( .A(n14001), .ZN(n14008) );
  OAI222_X1 U13764 ( .A1(n11492), .A2(n10997), .B1(n10996), .B2(n10995), .C1(
        n14008), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13765 ( .A(n10998), .ZN(n10999) );
  AOI21_X1 U13766 ( .B1(n11001), .B2(n11000), .A(n10999), .ZN(n14662) );
  NAND2_X1 U13767 ( .A1(n11002), .A2(n12790), .ZN(n12814) );
  NAND2_X1 U13768 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n12814), .ZN(n11003) );
  OAI21_X1 U13769 ( .B1(n14662), .B2(n14619), .A(n11003), .ZN(n11004) );
  AOI21_X1 U13770 ( .B1(n14591), .B2(n11669), .A(n11004), .ZN(n11005) );
  OAI21_X1 U13771 ( .B1(n11693), .B2(n14633), .A(n11005), .ZN(P1_U3232) );
  NOR2_X1 U13772 ( .A1(n12570), .A2(n14943), .ZN(n12045) );
  INV_X1 U13773 ( .A(n12045), .ZN(n11006) );
  INV_X1 U13774 ( .A(n14571), .ZN(n14628) );
  OAI22_X1 U13775 ( .A1(n14609), .A2(n12036), .B1(n11006), .B2(n14628), .ZN(
        n11007) );
  AOI21_X1 U13776 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n12814), .A(n11007), .ZN(
        n11012) );
  NAND2_X1 U13777 ( .A1(n11010), .A2(n14621), .ZN(n11011) );
  OAI211_X1 U13778 ( .C1(n15410), .C2(n14633), .A(n11012), .B(n11011), .ZN(
        P1_U3222) );
  AOI21_X1 U13779 ( .B1(n11014), .B2(n11013), .A(n14619), .ZN(n11016) );
  NAND2_X1 U13780 ( .A1(n11016), .A2(n11015), .ZN(n11019) );
  AOI22_X1 U13781 ( .A1(n15031), .A2(n14648), .B1(n14650), .B2(n15029), .ZN(
        n11724) );
  NAND2_X1 U13782 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14684) );
  OAI21_X1 U13783 ( .B1(n14628), .B2(n11724), .A(n14684), .ZN(n11017) );
  AOI21_X1 U13784 ( .B1(n14630), .B2(n8894), .A(n11017), .ZN(n11018) );
  OAI211_X1 U13785 ( .C1(n11674), .C2(n14633), .A(n11019), .B(n11018), .ZN(
        P1_U3218) );
  NAND2_X1 U13786 ( .A1(n11022), .A2(n11021), .ZN(n11025) );
  NAND2_X1 U13787 ( .A1(n11023), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n11024) );
  XNOR2_X1 U13788 ( .A(n11757), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n11756) );
  XNOR2_X1 U13789 ( .A(n11755), .B(n11756), .ZN(n11751) );
  INV_X1 U13790 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15781) );
  XNOR2_X1 U13791 ( .A(n11749), .B(n15781), .ZN(SUB_1596_U54) );
  NAND2_X1 U13792 ( .A1(n11027), .A2(n12485), .ZN(n11063) );
  OAI21_X1 U13793 ( .B1(n11027), .B2(n12485), .A(n11063), .ZN(n11211) );
  NOR2_X1 U13794 ( .A1(n11028), .A2(n12485), .ZN(n11067) );
  NAND2_X1 U13795 ( .A1(n11028), .A2(n12485), .ZN(n11029) );
  NAND2_X1 U13796 ( .A1(n11029), .A2(n13398), .ZN(n11030) );
  OR2_X1 U13797 ( .A1(n11067), .A2(n11030), .ZN(n11032) );
  AOI22_X1 U13798 ( .A1(n13396), .A2(n13113), .B1(n13352), .B2(n13115), .ZN(
        n11031) );
  NAND2_X1 U13799 ( .A1(n11032), .A2(n11031), .ZN(n11208) );
  AOI21_X1 U13800 ( .B1(n13474), .B2(n11211), .A(n11208), .ZN(n11217) );
  INV_X1 U13801 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n11033) );
  OAI22_X1 U13802 ( .A1(n11220), .A2(n13536), .B1(n15691), .B2(n11033), .ZN(
        n11034) );
  INV_X1 U13803 ( .A(n11034), .ZN(n11035) );
  OAI21_X1 U13804 ( .B1(n15693), .B2(n11217), .A(n11035), .ZN(P3_U3399) );
  OR2_X1 U13805 ( .A1(n11037), .A2(n11036), .ZN(n11038) );
  AND2_X1 U13806 ( .A1(n11039), .A2(n11038), .ZN(n15672) );
  AOI22_X1 U13807 ( .A1(n13396), .A2(n13114), .B1(n13352), .B2(n7138), .ZN(
        n11043) );
  XNOR2_X1 U13808 ( .A(n12483), .B(n11040), .ZN(n11041) );
  NAND2_X1 U13809 ( .A1(n13398), .A2(n11041), .ZN(n11042) );
  OAI211_X1 U13810 ( .C1(n13313), .C2(n15672), .A(n11043), .B(n11042), .ZN(
        n15674) );
  OR2_X1 U13811 ( .A1(n11358), .A2(n11044), .ZN(n15671) );
  OAI21_X1 U13812 ( .B1(n15672), .B2(n11359), .A(n15671), .ZN(n11045) );
  NOR2_X1 U13813 ( .A1(n15674), .A2(n11045), .ZN(n15692) );
  MUX2_X1 U13814 ( .A(n11046), .B(n15692), .S(n13486), .Z(n11047) );
  INV_X1 U13815 ( .A(n11047), .ZN(P3_U3461) );
  OAI21_X1 U13816 ( .B1(n11049), .B2(n12491), .A(n11048), .ZN(n11093) );
  NAND2_X1 U13817 ( .A1(n11050), .A2(n6709), .ZN(n11051) );
  XNOR2_X1 U13818 ( .A(n11051), .B(n12491), .ZN(n11052) );
  NAND2_X1 U13819 ( .A1(n11052), .A2(n13398), .ZN(n11054) );
  AOI22_X1 U13820 ( .A1(n13352), .A2(n13111), .B1(n13396), .B2(n13109), .ZN(
        n11053) );
  NAND2_X1 U13821 ( .A1(n11054), .A2(n11053), .ZN(n11095) );
  AOI21_X1 U13822 ( .B1(n11093), .B2(n13474), .A(n11095), .ZN(n11214) );
  AOI22_X1 U13823 ( .A1(n13520), .A2(n11094), .B1(P3_REG0_REG_7__SCAN_IN), 
        .B2(n15693), .ZN(n11055) );
  OAI21_X1 U13824 ( .B1(n11214), .B2(n15693), .A(n11055), .ZN(P3_U3411) );
  OAI21_X1 U13825 ( .B1(n11057), .B2(n7206), .A(n11056), .ZN(n11086) );
  OAI21_X1 U13826 ( .B1(n6716), .B2(n12493), .A(n11058), .ZN(n11059) );
  NAND2_X1 U13827 ( .A1(n11059), .A2(n13398), .ZN(n11061) );
  AOI22_X1 U13828 ( .A1(n13352), .A2(n13110), .B1(n13396), .B2(n13108), .ZN(
        n11060) );
  NAND2_X1 U13829 ( .A1(n11061), .A2(n11060), .ZN(n11087) );
  AOI21_X1 U13830 ( .B1(n11086), .B2(n13474), .A(n11087), .ZN(n11100) );
  AOI22_X1 U13831 ( .A1(n13520), .A2(n11819), .B1(P3_REG0_REG_8__SCAN_IN), 
        .B2(n15693), .ZN(n11062) );
  OAI21_X1 U13832 ( .B1(n11100), .B2(n15693), .A(n11062), .ZN(P3_U3414) );
  NAND2_X1 U13833 ( .A1(n11063), .A2(n12376), .ZN(n11065) );
  XNOR2_X1 U13834 ( .A(n11065), .B(n12486), .ZN(n11221) );
  NOR2_X1 U13835 ( .A1(n11067), .A2(n11066), .ZN(n11068) );
  XNOR2_X1 U13836 ( .A(n11068), .B(n12486), .ZN(n11070) );
  AOI22_X1 U13837 ( .A1(n13396), .A2(n13112), .B1(n13352), .B2(n13114), .ZN(
        n11069) );
  OAI21_X1 U13838 ( .B1(n11070), .B2(n13428), .A(n11069), .ZN(n11222) );
  AOI21_X1 U13839 ( .B1(n11221), .B2(n13474), .A(n11222), .ZN(n11243) );
  INV_X1 U13840 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n11071) );
  OAI22_X1 U13841 ( .A1(n11246), .A2(n13536), .B1(n15691), .B2(n11071), .ZN(
        n11072) );
  INV_X1 U13842 ( .A(n11072), .ZN(n11073) );
  OAI21_X1 U13843 ( .B1(n11243), .B2(n15693), .A(n11073), .ZN(P3_U3402) );
  INV_X1 U13844 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11083) );
  INV_X1 U13845 ( .A(n11074), .ZN(n11075) );
  NAND2_X1 U13846 ( .A1(n11076), .A2(n11075), .ZN(n11999) );
  AND2_X1 U13847 ( .A1(n11999), .A2(n12004), .ZN(n12001) );
  NOR2_X1 U13848 ( .A1(n12001), .A2(n11077), .ZN(n11254) );
  OAI21_X1 U13849 ( .B1(n11254), .B2(n6713), .A(n11078), .ZN(n11518) );
  XNOR2_X1 U13850 ( .A(n11518), .B(n13907), .ZN(n11588) );
  XNOR2_X1 U13851 ( .A(n11521), .B(n13907), .ZN(n11080) );
  AOI21_X1 U13852 ( .B1(n11080), .B2(n14307), .A(n11079), .ZN(n11580) );
  AOI211_X1 U13853 ( .C1(n13726), .C2(n11604), .A(n8582), .B(n11527), .ZN(
        n11585) );
  AOI21_X1 U13854 ( .B1(n15651), .B2(n13726), .A(n11585), .ZN(n11081) );
  OAI211_X1 U13855 ( .C1(n11588), .C2(n15655), .A(n11580), .B(n11081), .ZN(
        n11084) );
  NAND2_X1 U13856 ( .A1(n11084), .A2(n15659), .ZN(n11082) );
  OAI21_X1 U13857 ( .B1(n15659), .B2(n11083), .A(n11082), .ZN(P2_U3445) );
  NAND2_X1 U13858 ( .A1(n11084), .A2(n15670), .ZN(n11085) );
  OAI21_X1 U13859 ( .B1(n15670), .B2(n10488), .A(n11085), .ZN(P2_U3504) );
  INV_X1 U13860 ( .A(n11086), .ZN(n11092) );
  AOI22_X1 U13861 ( .A1(n13438), .A2(n11819), .B1(n15675), .B2(n11820), .ZN(
        n11091) );
  INV_X1 U13862 ( .A(n11087), .ZN(n11089) );
  MUX2_X1 U13863 ( .A(n11089), .B(n11088), .S(n15688), .Z(n11090) );
  OAI211_X1 U13864 ( .C1(n11092), .C2(n13441), .A(n11091), .B(n11090), .ZN(
        P3_U3225) );
  INV_X1 U13865 ( .A(n11093), .ZN(n11099) );
  AOI22_X1 U13866 ( .A1(n13438), .A2(n11094), .B1(n15675), .B2(n11648), .ZN(
        n11098) );
  MUX2_X1 U13867 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n11095), .S(n13405), .Z(
        n11096) );
  INV_X1 U13868 ( .A(n11096), .ZN(n11097) );
  OAI211_X1 U13869 ( .C1(n11099), .C2(n13441), .A(n11098), .B(n11097), .ZN(
        P3_U3226) );
  INV_X1 U13870 ( .A(n11819), .ZN(n11103) );
  MUX2_X1 U13871 ( .A(n11101), .B(n11100), .S(n13486), .Z(n11102) );
  OAI21_X1 U13872 ( .B1(n11103), .B2(n13482), .A(n11102), .ZN(P3_U3467) );
  XNOR2_X1 U13873 ( .A(n11618), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n11616) );
  INV_X1 U13874 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11104) );
  OAI22_X1 U13875 ( .A1(n11107), .A2(n11106), .B1(n11105), .B2(n11104), .ZN(
        n11617) );
  XOR2_X1 U13876 ( .A(n11616), .B(n11617), .Z(n11118) );
  INV_X1 U13877 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15250) );
  NAND2_X1 U13878 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n12136)
         );
  OAI21_X1 U13879 ( .B1(n15609), .B2(n15250), .A(n12136), .ZN(n11116) );
  NAND2_X1 U13880 ( .A1(n11113), .A2(n11111), .ZN(n11109) );
  INV_X1 U13881 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11108) );
  MUX2_X1 U13882 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11108), .S(n11618), .Z(
        n11110) );
  NAND2_X1 U13883 ( .A1(n11109), .A2(n11110), .ZN(n11620) );
  INV_X1 U13884 ( .A(n11110), .ZN(n11112) );
  NAND3_X1 U13885 ( .A1(n11113), .A2(n11112), .A3(n11111), .ZN(n11114) );
  AOI21_X1 U13886 ( .B1(n11620), .B2(n11114), .A(n15579), .ZN(n11115) );
  AOI211_X1 U13887 ( .C1(n15595), .C2(n11618), .A(n11116), .B(n11115), .ZN(
        n11117) );
  OAI21_X1 U13888 ( .B1(n11118), .B2(n15586), .A(n11117), .ZN(P2_U3226) );
  OR2_X1 U13889 ( .A1(n11133), .A2(n12489), .ZN(n11135) );
  NAND2_X1 U13890 ( .A1(n11135), .A2(n11119), .ZN(n11120) );
  XNOR2_X1 U13891 ( .A(n11121), .B(n11120), .ZN(n11125) );
  NAND2_X1 U13892 ( .A1(n13396), .A2(n13110), .ZN(n11123) );
  NAND2_X1 U13893 ( .A1(n13352), .A2(n13112), .ZN(n11122) );
  NAND2_X1 U13894 ( .A1(n11123), .A2(n11122), .ZN(n11124) );
  AOI21_X1 U13895 ( .B1(n11125), .B2(n13398), .A(n11124), .ZN(n11163) );
  OR2_X1 U13896 ( .A1(n11126), .A2(n12490), .ZN(n11127) );
  NAND2_X1 U13897 ( .A1(n11128), .A2(n11127), .ZN(n11161) );
  NAND2_X1 U13898 ( .A1(n11161), .A2(n13474), .ZN(n11129) );
  NAND2_X1 U13899 ( .A1(n11163), .A2(n11129), .ZN(n11167) );
  INV_X1 U13900 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11130) );
  OAI22_X1 U13901 ( .A1(n11656), .A2(n13536), .B1(n15691), .B2(n11130), .ZN(
        n11131) );
  AOI21_X1 U13902 ( .B1(n11167), .B2(n15691), .A(n11131), .ZN(n11132) );
  INV_X1 U13903 ( .A(n11132), .ZN(P3_U3408) );
  NAND2_X1 U13904 ( .A1(n11133), .A2(n12489), .ZN(n11134) );
  NAND2_X1 U13905 ( .A1(n11135), .A2(n11134), .ZN(n11136) );
  NAND2_X1 U13906 ( .A1(n11136), .A2(n13398), .ZN(n11138) );
  AOI22_X1 U13907 ( .A1(n13396), .A2(n13111), .B1(n13352), .B2(n13113), .ZN(
        n11137) );
  AND2_X1 U13908 ( .A1(n11138), .A2(n11137), .ZN(n11187) );
  OR2_X1 U13909 ( .A1(n11139), .A2(n12489), .ZN(n11140) );
  NAND2_X1 U13910 ( .A1(n11141), .A2(n11140), .ZN(n11185) );
  NAND2_X1 U13911 ( .A1(n13474), .A2(n11185), .ZN(n11142) );
  NAND2_X1 U13912 ( .A1(n11187), .A2(n11142), .ZN(n11204) );
  INV_X1 U13913 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11143) );
  OAI22_X1 U13914 ( .A1(n11631), .A2(n13536), .B1(n15691), .B2(n11143), .ZN(
        n11144) );
  AOI21_X1 U13915 ( .B1(n15691), .B2(n11204), .A(n11144), .ZN(n11145) );
  INV_X1 U13916 ( .A(n11145), .ZN(P3_U3405) );
  INV_X1 U13917 ( .A(n11359), .ZN(n13465) );
  XNOR2_X1 U13918 ( .A(n11146), .B(n12497), .ZN(n11157) );
  INV_X1 U13919 ( .A(n11157), .ZN(n11150) );
  AOI22_X1 U13920 ( .A1(n13352), .A2(n13109), .B1(n13396), .B2(n13107), .ZN(
        n11149) );
  OAI211_X1 U13921 ( .C1(n6581), .C2(n12497), .A(n11147), .B(n13398), .ZN(
        n11148) );
  OAI211_X1 U13922 ( .C1(n11157), .C2(n13313), .A(n11149), .B(n11148), .ZN(
        n11152) );
  AOI21_X1 U13923 ( .B1(n13465), .B2(n11150), .A(n11152), .ZN(n11240) );
  INV_X1 U13924 ( .A(n11793), .ZN(n11154) );
  AOI22_X1 U13925 ( .A1(n13520), .A2(n11154), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n15693), .ZN(n11151) );
  OAI21_X1 U13926 ( .B1(n11240), .B2(n15693), .A(n11151), .ZN(P3_U3417) );
  NOR2_X1 U13927 ( .A1(n15688), .A2(n15677), .ZN(n13377) );
  INV_X1 U13928 ( .A(n13377), .ZN(n13363) );
  INV_X1 U13929 ( .A(n11152), .ZN(n11153) );
  MUX2_X1 U13930 ( .A(n11300), .B(n11153), .S(n13405), .Z(n11156) );
  AOI22_X1 U13931 ( .A1(n13438), .A2(n11154), .B1(n15675), .B2(n11790), .ZN(
        n11155) );
  OAI211_X1 U13932 ( .C1(n11157), .C2(n13363), .A(n11156), .B(n11155), .ZN(
        P3_U3224) );
  INV_X1 U13933 ( .A(n8831), .ZN(n11160) );
  OAI222_X1 U13934 ( .A1(n15232), .A2(n11158), .B1(n15236), .B2(n11160), .C1(
        P1_U3086), .C2(n12556), .ZN(P1_U3336) );
  OAI222_X1 U13935 ( .A1(n11528), .A2(P2_U3088), .B1(n10996), .B2(n11160), 
        .C1(n11159), .C2(n14478), .ZN(P2_U3308) );
  INV_X1 U13936 ( .A(n11161), .ZN(n11166) );
  MUX2_X1 U13937 ( .A(n11163), .B(n11162), .S(n15688), .Z(n11165) );
  AOI22_X1 U13938 ( .A1(n13438), .A2(n11169), .B1(n15675), .B2(n11652), .ZN(
        n11164) );
  OAI211_X1 U13939 ( .C1(n11166), .C2(n13441), .A(n11165), .B(n11164), .ZN(
        P3_U3227) );
  MUX2_X1 U13940 ( .A(n11167), .B(P3_REG1_REG_6__SCAN_IN), .S(n13478), .Z(
        n11168) );
  AOI21_X1 U13941 ( .B1(n13469), .B2(n11169), .A(n11168), .ZN(n11170) );
  INV_X1 U13942 ( .A(n11170), .ZN(P3_U3465) );
  NAND3_X1 U13943 ( .A1(n13288), .A2(n13242), .A3(n13277), .ZN(n11179) );
  AOI21_X1 U13944 ( .B1(n13248), .B2(n7916), .A(n13284), .ZN(n11173) );
  AOI22_X1 U13945 ( .A1(n15694), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11171) );
  OAI21_X1 U13946 ( .B1(n11173), .B2(n11172), .A(n11171), .ZN(n11178) );
  AOI21_X1 U13947 ( .B1(n9573), .B2(n13248), .A(n13209), .ZN(n11175) );
  NOR2_X1 U13948 ( .A1(n11175), .A2(n11174), .ZN(n11176) );
  MUX2_X1 U13949 ( .A(n13279), .B(n11176), .S(n9400), .Z(n11177) );
  AOI211_X1 U13950 ( .C1(n11180), .C2(n11179), .A(n11178), .B(n11177), .ZN(
        n11181) );
  INV_X1 U13951 ( .A(n11181), .ZN(P3_U3182) );
  INV_X1 U13952 ( .A(n11182), .ZN(n11184) );
  OAI222_X1 U13953 ( .A1(P3_U3151), .A2(n10043), .B1(n12962), .B2(n11184), 
        .C1(n11183), .C2(n13550), .ZN(P3_U3275) );
  INV_X1 U13954 ( .A(n11185), .ZN(n11190) );
  MUX2_X1 U13955 ( .A(n11187), .B(n11186), .S(n15688), .Z(n11189) );
  AOI22_X1 U13956 ( .A1(n13438), .A2(n11206), .B1(n15675), .B2(n11635), .ZN(
        n11188) );
  OAI211_X1 U13957 ( .C1(n11190), .C2(n13441), .A(n11189), .B(n11188), .ZN(
        P3_U3228) );
  NAND2_X1 U13958 ( .A1(n11192), .A2(n11191), .ZN(n11194) );
  XOR2_X1 U13959 ( .A(n11194), .B(n11193), .Z(n11201) );
  OAI21_X1 U13960 ( .B1(n13718), .B2(n11435), .A(n11195), .ZN(n11199) );
  INV_X1 U13961 ( .A(n11196), .ZN(n11559) );
  OAI22_X1 U13962 ( .A1(n11197), .A2(n13587), .B1(n13717), .B2(n11559), .ZN(
        n11198) );
  AOI211_X1 U13963 ( .C1(n13789), .C2(n13693), .A(n11199), .B(n11198), .ZN(
        n11200) );
  OAI21_X1 U13964 ( .B1(n11201), .B2(n13695), .A(n11200), .ZN(P2_U3193) );
  INV_X1 U13965 ( .A(n11202), .ZN(n11317) );
  OAI222_X1 U13966 ( .A1(n15236), .A2(n11317), .B1(n12558), .B2(n6537), .C1(
        n11203), .C2(n15232), .ZN(P1_U3335) );
  MUX2_X1 U13967 ( .A(P3_REG1_REG_5__SCAN_IN), .B(n11204), .S(n13486), .Z(
        n11205) );
  AOI21_X1 U13968 ( .B1(n13469), .B2(n11206), .A(n11205), .ZN(n11207) );
  INV_X1 U13969 ( .A(n11207), .ZN(P3_U3464) );
  INV_X1 U13970 ( .A(n13441), .ZN(n11212) );
  MUX2_X1 U13971 ( .A(n11208), .B(P3_REG2_REG_3__SCAN_IN), .S(n15688), .Z(
        n11210) );
  OAI22_X1 U13972 ( .A1(n13403), .A2(n11220), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15681), .ZN(n11209) );
  AOI211_X1 U13973 ( .C1(n11212), .C2(n11211), .A(n11210), .B(n11209), .ZN(
        n11213) );
  INV_X1 U13974 ( .A(n11213), .ZN(P3_U3230) );
  MUX2_X1 U13975 ( .A(n11215), .B(n11214), .S(n13486), .Z(n11216) );
  OAI21_X1 U13976 ( .B1(n13482), .B2(n11644), .A(n11216), .ZN(P3_U3466) );
  MUX2_X1 U13977 ( .A(n11218), .B(n11217), .S(n13486), .Z(n11219) );
  OAI21_X1 U13978 ( .B1(n13482), .B2(n11220), .A(n11219), .ZN(P3_U3462) );
  INV_X1 U13979 ( .A(n11221), .ZN(n11226) );
  INV_X1 U13980 ( .A(n11222), .ZN(n11223) );
  MUX2_X1 U13981 ( .A(n9410), .B(n11223), .S(n13405), .Z(n11225) );
  AOI22_X1 U13982 ( .A1(n13438), .A2(n11507), .B1(n15675), .B2(n11511), .ZN(
        n11224) );
  OAI211_X1 U13983 ( .C1(n13441), .C2(n11226), .A(n11225), .B(n11224), .ZN(
        P3_U3229) );
  INV_X1 U13984 ( .A(n11227), .ZN(n11228) );
  NAND4_X1 U13985 ( .A1(n11229), .A2(n15615), .A3(n11228), .A4(n15614), .ZN(
        n11230) );
  NAND2_X1 U13986 ( .A1(n13940), .A2(n13941), .ZN(n11514) );
  INV_X1 U13987 ( .A(n11514), .ZN(n11231) );
  NAND2_X1 U13988 ( .A1(n14293), .A2(n11231), .ZN(n14265) );
  INV_X1 U13989 ( .A(n13756), .ZN(n13757) );
  NAND2_X1 U13990 ( .A1(n11232), .A2(n13757), .ZN(n11234) );
  NAND2_X1 U13991 ( .A1(n11234), .A2(n11233), .ZN(n15621) );
  NAND2_X1 U13992 ( .A1(n13756), .A2(n11235), .ZN(n15619) );
  AOI21_X1 U13993 ( .B1(n14217), .B2(n15642), .A(n15621), .ZN(n11236) );
  AOI21_X1 U13994 ( .B1(n14304), .B2(n13981), .A(n11236), .ZN(n15620) );
  OAI21_X1 U13995 ( .B1(n13940), .B2(n15619), .A(n15620), .ZN(n11237) );
  NAND2_X1 U13996 ( .A1(n11237), .A2(n14293), .ZN(n11239) );
  INV_X1 U13997 ( .A(n14290), .ZN(n14272) );
  AOI22_X1 U13998 ( .A1(n14308), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n14272), .ZN(n11238) );
  OAI211_X1 U13999 ( .C1(n14265), .C2(n15621), .A(n11239), .B(n11238), .ZN(
        P2_U3265) );
  MUX2_X1 U14000 ( .A(n11241), .B(n11240), .S(n13486), .Z(n11242) );
  OAI21_X1 U14001 ( .B1(n13482), .B2(n11793), .A(n11242), .ZN(P3_U3468) );
  MUX2_X1 U14002 ( .A(n11244), .B(n11243), .S(n13486), .Z(n11245) );
  OAI21_X1 U14003 ( .B1(n13482), .B2(n11246), .A(n11245), .ZN(P3_U3463) );
  XNOR2_X1 U14004 ( .A(n11247), .B(n12494), .ZN(n11297) );
  INV_X1 U14005 ( .A(n11297), .ZN(n11252) );
  AOI22_X1 U14006 ( .A1(n13352), .A2(n13108), .B1(n13396), .B2(n13106), .ZN(
        n11251) );
  OAI211_X1 U14007 ( .C1(n11249), .C2(n12494), .A(n11248), .B(n13398), .ZN(
        n11250) );
  OAI211_X1 U14008 ( .C1(n11297), .C2(n13313), .A(n11251), .B(n11250), .ZN(
        n11292) );
  AOI21_X1 U14009 ( .B1(n13465), .B2(n11252), .A(n11292), .ZN(n11366) );
  INV_X1 U14010 ( .A(n11910), .ZN(n11294) );
  AOI22_X1 U14011 ( .A1(n13520), .A2(n11294), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n15693), .ZN(n11253) );
  OAI21_X1 U14012 ( .B1(n11366), .B2(n15693), .A(n11253), .ZN(P3_U3420) );
  NOR2_X1 U14013 ( .A1(n11254), .A2(n13910), .ZN(n11590) );
  AOI21_X1 U14014 ( .B1(n11254), .B2(n13910), .A(n11590), .ZN(n11570) );
  OAI21_X1 U14015 ( .B1(n11255), .B2(n13910), .A(n11594), .ZN(n11260) );
  OAI22_X1 U14016 ( .A1(n11257), .A2(n14116), .B1(n11256), .B2(n14118), .ZN(
        n11259) );
  NOR2_X1 U14017 ( .A1(n11570), .A2(n15642), .ZN(n11258) );
  AOI211_X1 U14018 ( .C1(n14307), .C2(n11260), .A(n11259), .B(n11258), .ZN(
        n11564) );
  AOI21_X1 U14019 ( .B1(n11261), .B2(n13767), .A(n8582), .ZN(n11262) );
  AND2_X1 U14020 ( .A1(n11262), .A2(n11606), .ZN(n11567) );
  INV_X1 U14021 ( .A(n11567), .ZN(n11263) );
  OAI211_X1 U14022 ( .C1(n11570), .C2(n15636), .A(n11564), .B(n11263), .ZN(
        n11269) );
  OAI22_X1 U14023 ( .A1(n14400), .A2(n13769), .B1(n15670), .B2(n11264), .ZN(
        n11265) );
  AOI21_X1 U14024 ( .B1(n11269), .B2(n15670), .A(n11265), .ZN(n11266) );
  INV_X1 U14025 ( .A(n11266), .ZN(P2_U3502) );
  INV_X1 U14026 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11267) );
  OAI22_X1 U14027 ( .A1(n14459), .A2(n13769), .B1(n15659), .B2(n11267), .ZN(
        n11268) );
  AOI21_X1 U14028 ( .B1(n11269), .B2(n15659), .A(n11268), .ZN(n11270) );
  INV_X1 U14029 ( .A(n11270), .ZN(P2_U3439) );
  OAI211_X1 U14030 ( .C1(n11271), .C2(n11273), .A(n11272), .B(n14621), .ZN(
        n11276) );
  AOI22_X1 U14031 ( .A1(n15031), .A2(n14645), .B1(n14647), .B2(n15029), .ZN(
        n15354) );
  NAND2_X1 U14032 ( .A1(n6537), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14713) );
  OAI21_X1 U14033 ( .B1(n14628), .B2(n15354), .A(n14713), .ZN(n11274) );
  AOI21_X1 U14034 ( .B1(n15358), .B2(n14630), .A(n11274), .ZN(n11275) );
  OAI211_X1 U14035 ( .C1(n15440), .C2(n14633), .A(n11276), .B(n11275), .ZN(
        P1_U3239) );
  XNOR2_X1 U14036 ( .A(n11277), .B(n12498), .ZN(n11376) );
  OR2_X1 U14037 ( .A1(n11280), .A2(n12498), .ZN(n11281) );
  NAND3_X1 U14038 ( .A1(n11279), .A2(n11281), .A3(n13398), .ZN(n11283) );
  AOI22_X1 U14039 ( .A1(n13352), .A2(n13107), .B1(n13396), .B2(n13105), .ZN(
        n11282) );
  INV_X1 U14040 ( .A(n11372), .ZN(n11284) );
  NAND2_X1 U14041 ( .A1(n11284), .A2(n15691), .ZN(n11286) );
  INV_X1 U14042 ( .A(n12240), .ZN(n11373) );
  AOI22_X1 U14043 ( .A1(n13520), .A2(n11373), .B1(P3_REG0_REG_11__SCAN_IN), 
        .B2(n15693), .ZN(n11285) );
  OAI211_X1 U14044 ( .C1(n11376), .C2(n13540), .A(n11286), .B(n11285), .ZN(
        P3_U3423) );
  INV_X1 U14045 ( .A(n11287), .ZN(n11290) );
  OAI222_X1 U14046 ( .A1(n11289), .A2(P2_U3088), .B1(n10996), .B2(n11290), 
        .C1(n11288), .C2(n14478), .ZN(P2_U3306) );
  OAI222_X1 U14047 ( .A1(n15232), .A2(n11291), .B1(n15236), .B2(n11290), .C1(
        n6537), .C2(n12557), .ZN(P1_U3334) );
  INV_X1 U14048 ( .A(n11292), .ZN(n11293) );
  MUX2_X1 U14049 ( .A(n15928), .B(n11293), .S(n13405), .Z(n11296) );
  AOI22_X1 U14050 ( .A1(n13438), .A2(n11294), .B1(n15675), .B2(n11907), .ZN(
        n11295) );
  OAI211_X1 U14051 ( .C1(n11297), .C2(n13363), .A(n11296), .B(n11295), .ZN(
        P3_U3223) );
  INV_X1 U14052 ( .A(n11470), .ZN(n11298) );
  AOI21_X1 U14053 ( .B1(n11300), .B2(n11299), .A(n11298), .ZN(n11315) );
  INV_X1 U14054 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n11302) );
  AND2_X1 U14055 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11787) );
  INV_X1 U14056 ( .A(n11787), .ZN(n11301) );
  OAI21_X1 U14057 ( .B1(n13273), .B2(n11302), .A(n11301), .ZN(n11308) );
  NAND3_X1 U14058 ( .A1(n11305), .A2(n11304), .A3(n11303), .ZN(n11306) );
  AOI21_X1 U14059 ( .B1(n11475), .B2(n11306), .A(n13277), .ZN(n11307) );
  AOI211_X1 U14060 ( .C1(n11309), .C2(n13279), .A(n11308), .B(n11307), .ZN(
        n11314) );
  NOR2_X1 U14061 ( .A1(n11310), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n11312) );
  OAI21_X1 U14062 ( .B1(n11312), .B2(n11311), .A(n13284), .ZN(n11313) );
  OAI211_X1 U14063 ( .C1(n11315), .C2(n13288), .A(n11314), .B(n11313), .ZN(
        P3_U3191) );
  OAI222_X1 U14064 ( .A1(P2_U3088), .A2(n8541), .B1(n10996), .B2(n11317), .C1(
        n11316), .C2(n14478), .ZN(P2_U3307) );
  INV_X1 U14065 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n15827) );
  NAND2_X1 U14066 ( .A1(n13353), .A2(P3_U3897), .ZN(n11318) );
  OAI21_X1 U14067 ( .B1(P3_U3897), .B2(n15827), .A(n11318), .ZN(P3_U3516) );
  NAND3_X1 U14068 ( .A1(n11279), .A2(n7893), .A3(n11319), .ZN(n11320) );
  NAND3_X1 U14069 ( .A1(n11321), .A2(n13398), .A3(n11320), .ZN(n11323) );
  AOI22_X1 U14070 ( .A1(n13396), .A2(n13104), .B1(n13352), .B2(n13106), .ZN(
        n11322) );
  OAI21_X1 U14071 ( .B1(n11325), .B2(n7893), .A(n11324), .ZN(n11497) );
  INV_X1 U14072 ( .A(n13540), .ZN(n13529) );
  NAND2_X1 U14073 ( .A1(n11497), .A2(n13529), .ZN(n11327) );
  AOI22_X1 U14074 ( .A1(n13520), .A2(n11498), .B1(P3_REG0_REG_12__SCAN_IN), 
        .B2(n15693), .ZN(n11326) );
  OAI211_X1 U14075 ( .C1(n15693), .C2(n11500), .A(n11327), .B(n11326), .ZN(
        P3_U3426) );
  NAND2_X1 U14076 ( .A1(n11329), .A2(n11328), .ZN(n11330) );
  NAND2_X1 U14077 ( .A1(n11331), .A2(n11330), .ZN(n11449) );
  XNOR2_X1 U14078 ( .A(n11449), .B(n11344), .ZN(n11447) );
  XNOR2_X1 U14079 ( .A(n11447), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n11346) );
  INV_X1 U14080 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U14081 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14627)
         );
  OAI21_X1 U14082 ( .B1(n14815), .B2(n11332), .A(n14627), .ZN(n11343) );
  NAND2_X1 U14083 ( .A1(n11334), .A2(n11333), .ZN(n11337) );
  NAND2_X1 U14084 ( .A1(n11335), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11336) );
  NAND2_X1 U14085 ( .A1(n11337), .A2(n11336), .ZN(n11338) );
  NAND2_X1 U14086 ( .A1(n11338), .A2(n11344), .ZN(n11339) );
  NAND2_X1 U14087 ( .A1(n11340), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11341) );
  AOI21_X1 U14088 ( .B1(n11441), .B2(n11341), .A(n14805), .ZN(n11342) );
  AOI211_X1 U14089 ( .C1(n15340), .C2(n11344), .A(n11343), .B(n11342), .ZN(
        n11345) );
  OAI21_X1 U14090 ( .B1(n11347), .B2(n11346), .A(n11345), .ZN(P1_U3258) );
  INV_X1 U14091 ( .A(n11348), .ZN(n11350) );
  OAI22_X1 U14092 ( .A1(n12367), .A2(P3_U3151), .B1(SI_22_), .B2(n13550), .ZN(
        n11349) );
  AOI21_X1 U14093 ( .B1(n11350), .B2(n11728), .A(n11349), .ZN(P3_U3273) );
  INV_X1 U14094 ( .A(n11411), .ZN(n11351) );
  NAND2_X1 U14095 ( .A1(n13352), .A2(n13118), .ZN(n11353) );
  NAND2_X1 U14096 ( .A1(n13396), .A2(n13115), .ZN(n11352) );
  OAI211_X1 U14097 ( .C1(n13428), .C2(n11354), .A(n11353), .B(n11352), .ZN(
        n11355) );
  INV_X1 U14098 ( .A(n11355), .ZN(n11356) );
  OAI21_X1 U14099 ( .B1(n13313), .B2(n15678), .A(n11356), .ZN(n15685) );
  OR2_X1 U14100 ( .A1(n11358), .A2(n11357), .ZN(n15680) );
  OAI21_X1 U14101 ( .B1(n15678), .B2(n11359), .A(n15680), .ZN(n11360) );
  NOR2_X1 U14102 ( .A1(n15685), .A2(n11360), .ZN(n15689) );
  MUX2_X1 U14103 ( .A(n11361), .B(n15689), .S(n13486), .Z(n11362) );
  INV_X1 U14104 ( .A(n11362), .ZN(P3_U3460) );
  INV_X1 U14105 ( .A(n11363), .ZN(n11364) );
  OAI222_X1 U14106 ( .A1(n11492), .A2(n11365), .B1(n10996), .B2(n11364), .C1(
        P2_U3088), .C2(n13944), .ZN(P2_U3305) );
  MUX2_X1 U14107 ( .A(n11367), .B(n11366), .S(n13486), .Z(n11368) );
  OAI21_X1 U14108 ( .B1(n13482), .B2(n11910), .A(n11368), .ZN(P3_U3469) );
  MUX2_X1 U14109 ( .A(n11372), .B(n13161), .S(n15688), .Z(n11370) );
  AOI22_X1 U14110 ( .A1(n13438), .A2(n11373), .B1(n15675), .B2(n12245), .ZN(
        n11369) );
  OAI211_X1 U14111 ( .C1(n11376), .C2(n13441), .A(n11370), .B(n11369), .ZN(
        P3_U3222) );
  MUX2_X1 U14112 ( .A(n11372), .B(n11371), .S(n13478), .Z(n11375) );
  NAND2_X1 U14113 ( .A1(n13469), .A2(n11373), .ZN(n11374) );
  OAI211_X1 U14114 ( .C1(n13488), .C2(n11376), .A(n11375), .B(n11374), .ZN(
        P3_U3470) );
  NAND2_X1 U14115 ( .A1(n12598), .A2(n15189), .ZN(n15448) );
  OAI211_X1 U14116 ( .C1(n11379), .C2(n11378), .A(n11377), .B(n14621), .ZN(
        n11382) );
  AOI22_X1 U14117 ( .A1(n15029), .A2(n14646), .B1(n14644), .B2(n15031), .ZN(
        n11689) );
  NAND2_X1 U14118 ( .A1(n6537), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14727) );
  OAI21_X1 U14119 ( .B1(n14628), .B2(n11689), .A(n14727), .ZN(n11380) );
  AOI21_X1 U14120 ( .B1(n11699), .B2(n14630), .A(n11380), .ZN(n11381) );
  OAI211_X1 U14121 ( .C1(n11923), .C2(n15448), .A(n11382), .B(n11381), .ZN(
        P1_U3213) );
  INV_X1 U14122 ( .A(n11383), .ZN(n11384) );
  AOI21_X1 U14123 ( .B1(n11385), .B2(n7022), .A(n11384), .ZN(n11389) );
  AOI22_X1 U14124 ( .A1(n13722), .A2(n13974), .B1(n13701), .B2(n11874), .ZN(
        n11386) );
  NAND2_X1 U14125 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n15548) );
  OAI211_X1 U14126 ( .C1(n11778), .C2(n13718), .A(n11386), .B(n15548), .ZN(
        n11387) );
  AOI21_X1 U14127 ( .B1(n13794), .B2(n13693), .A(n11387), .ZN(n11388) );
  OAI21_X1 U14128 ( .B1(n11389), .B2(n13695), .A(n11388), .ZN(P2_U3203) );
  NAND2_X1 U14129 ( .A1(n11390), .A2(n13058), .ZN(n11398) );
  AOI21_X1 U14130 ( .B1(n11399), .B2(n11392), .A(n11391), .ZN(n11397) );
  OAI22_X1 U14131 ( .A1(n13093), .A2(n11414), .B1(n13072), .B2(n11632), .ZN(
        n11394) );
  MUX2_X1 U14132 ( .A(n13090), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n11393) );
  AOI211_X1 U14133 ( .C1(n11395), .C2(n13096), .A(n11394), .B(n11393), .ZN(
        n11396) );
  OAI21_X1 U14134 ( .B1(n11398), .B2(n11397), .A(n11396), .ZN(P3_U3158) );
  NOR2_X1 U14135 ( .A1(n13090), .A2(P3_U3151), .ZN(n11464) );
  OAI21_X1 U14136 ( .B1(n11401), .B2(n11400), .A(n11399), .ZN(n11402) );
  NAND2_X1 U14137 ( .A1(n11402), .A2(n13058), .ZN(n11407) );
  OAI22_X1 U14138 ( .A1(n13093), .A2(n10098), .B1(n13072), .B2(n11403), .ZN(
        n11404) );
  AOI21_X1 U14139 ( .B1(n11405), .B2(n13096), .A(n11404), .ZN(n11406) );
  OAI211_X1 U14140 ( .C1(n11464), .C2(n11408), .A(n11407), .B(n11406), .ZN(
        P3_U3177) );
  INV_X1 U14141 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15682) );
  OAI211_X1 U14142 ( .C1(n11412), .C2(n11411), .A(n11410), .B(n11409), .ZN(
        n11413) );
  NAND2_X1 U14143 ( .A1(n11413), .A2(n13058), .ZN(n11418) );
  OAI22_X1 U14144 ( .A1(n13093), .A2(n11415), .B1(n13072), .B2(n11414), .ZN(
        n11416) );
  AOI21_X1 U14145 ( .B1(n10097), .B2(n13096), .A(n11416), .ZN(n11417) );
  OAI211_X1 U14146 ( .C1(n11464), .C2(n15682), .A(n11418), .B(n11417), .ZN(
        P3_U3162) );
  XOR2_X1 U14147 ( .A(n11420), .B(n11419), .Z(n14566) );
  AOI22_X1 U14148 ( .A1(n14566), .A2(n14567), .B1(n11420), .B2(n11419), .ZN(
        n11424) );
  NAND2_X1 U14149 ( .A1(n11422), .A2(n11421), .ZN(n11423) );
  XNOR2_X1 U14150 ( .A(n11424), .B(n11423), .ZN(n11430) );
  NAND2_X1 U14151 ( .A1(n14648), .A2(n15029), .ZN(n11426) );
  NAND2_X1 U14152 ( .A1(n14646), .A2(n15031), .ZN(n11425) );
  AND2_X1 U14153 ( .A1(n11426), .A2(n11425), .ZN(n15432) );
  NAND2_X1 U14154 ( .A1(n14630), .A2(n12065), .ZN(n11427) );
  NAND2_X1 U14155 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14699) );
  OAI211_X1 U14156 ( .C1(n15432), .C2(n14628), .A(n11427), .B(n14699), .ZN(
        n11428) );
  AOI21_X1 U14157 ( .B1(n14617), .B2(n12586), .A(n11428), .ZN(n11429) );
  OAI21_X1 U14158 ( .B1(n11430), .B2(n14619), .A(n11429), .ZN(P1_U3227) );
  XNOR2_X1 U14159 ( .A(n11432), .B(n11431), .ZN(n11439) );
  INV_X1 U14160 ( .A(n11433), .ZN(n11963) );
  NAND2_X1 U14161 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n15550)
         );
  OAI22_X1 U14162 ( .A1(n11435), .A2(n14116), .B1(n11434), .B2(n14118), .ZN(
        n11958) );
  NAND2_X1 U14163 ( .A1(n13666), .A2(n11958), .ZN(n11436) );
  OAI211_X1 U14164 ( .C1(n13717), .C2(n11963), .A(n15550), .B(n11436), .ZN(
        n11437) );
  AOI21_X1 U14165 ( .B1(n14405), .B2(n13693), .A(n11437), .ZN(n11438) );
  OAI21_X1 U14166 ( .B1(n11439), .B2(n13695), .A(n11438), .ZN(P2_U3189) );
  INV_X1 U14167 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11442) );
  MUX2_X1 U14168 ( .A(n11442), .B(P1_REG2_REG_16__SCAN_IN), .S(n11802), .Z(
        n11443) );
  AOI21_X1 U14169 ( .B1(n11444), .B2(n11443), .A(n14805), .ZN(n11445) );
  NAND2_X1 U14170 ( .A1(n11445), .A2(n11799), .ZN(n11458) );
  NAND2_X1 U14171 ( .A1(n6537), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14539) );
  INV_X1 U14172 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11446) );
  NAND2_X1 U14173 ( .A1(n11447), .A2(n11446), .ZN(n11451) );
  NAND2_X1 U14174 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  NAND2_X1 U14175 ( .A1(n11451), .A2(n11450), .ZN(n11452) );
  XNOR2_X1 U14176 ( .A(n11802), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U14177 ( .A1(n11453), .A2(n11452), .ZN(n11454) );
  NAND3_X1 U14178 ( .A1(n15332), .A2(n11804), .A3(n11454), .ZN(n11455) );
  NAND2_X1 U14179 ( .A1(n14539), .A2(n11455), .ZN(n11456) );
  AOI21_X1 U14180 ( .B1(n15342), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11456), 
        .ZN(n11457) );
  OAI211_X1 U14181 ( .C1(n14804), .C2(n11459), .A(n11458), .B(n11457), .ZN(
        P1_U3259) );
  INV_X1 U14182 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11463) );
  OAI22_X1 U14183 ( .A1(n13081), .A2(n11460), .B1(n13072), .B2(n10098), .ZN(
        n11461) );
  AOI21_X1 U14184 ( .B1(n13058), .B2(n12484), .A(n11461), .ZN(n11462) );
  OAI21_X1 U14185 ( .B1(n11464), .B2(n11463), .A(n11462), .ZN(P3_U3172) );
  INV_X1 U14186 ( .A(n11465), .ZN(n11467) );
  NOR2_X1 U14187 ( .A1(n11467), .A2(n11466), .ZN(n11471) );
  INV_X1 U14188 ( .A(n11468), .ZN(n11469) );
  AOI21_X1 U14189 ( .B1(n11471), .B2(n11470), .A(n11469), .ZN(n11486) );
  INV_X1 U14190 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11472) );
  NAND2_X1 U14191 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11903)
         );
  OAI21_X1 U14192 ( .B1(n13273), .B2(n11472), .A(n11903), .ZN(n11479) );
  NAND3_X1 U14193 ( .A1(n11475), .A2(n11474), .A3(n11473), .ZN(n11476) );
  AOI21_X1 U14194 ( .B1(n11477), .B2(n11476), .A(n13277), .ZN(n11478) );
  AOI211_X1 U14195 ( .C1(n11480), .C2(n13279), .A(n11479), .B(n11478), .ZN(
        n11485) );
  NOR3_X1 U14196 ( .A1(n11311), .A2(n11482), .A3(n11481), .ZN(n11483) );
  OAI21_X1 U14197 ( .B1(n6720), .B2(n11483), .A(n13284), .ZN(n11484) );
  OAI211_X1 U14198 ( .C1(n11486), .C2(n13288), .A(n11485), .B(n11484), .ZN(
        P3_U3192) );
  INV_X1 U14199 ( .A(n13488), .ZN(n13477) );
  AOI22_X1 U14200 ( .A1(n11497), .A2(n13477), .B1(n13469), .B2(n11498), .ZN(
        n11489) );
  MUX2_X1 U14201 ( .A(n11500), .B(n11487), .S(n13478), .Z(n11488) );
  NAND2_X1 U14202 ( .A1(n11489), .A2(n11488), .ZN(P3_U3471) );
  NAND2_X1 U14203 ( .A1(n11494), .A2(n14470), .ZN(n11491) );
  OR2_X1 U14204 ( .A1(n11490), .A2(P2_U3088), .ZN(n13957) );
  OAI211_X1 U14205 ( .C1(n11493), .C2(n11492), .A(n11491), .B(n13957), .ZN(
        P2_U3304) );
  NAND2_X1 U14206 ( .A1(n11494), .A2(n15221), .ZN(n11495) );
  OAI211_X1 U14207 ( .C1(n11496), .C2(n15232), .A(n11495), .B(n12793), .ZN(
        P1_U3332) );
  INV_X1 U14208 ( .A(n11497), .ZN(n11503) );
  AOI22_X1 U14209 ( .A1(n11498), .A2(n13438), .B1(n15675), .B2(n12259), .ZN(
        n11502) );
  MUX2_X1 U14210 ( .A(n11500), .B(n11499), .S(n15688), .Z(n11501) );
  OAI211_X1 U14211 ( .C1(n11503), .C2(n13441), .A(n11502), .B(n11501), .ZN(
        P3_U3221) );
  AOI21_X1 U14212 ( .B1(n11506), .B2(n11505), .A(n11504), .ZN(n11513) );
  AOI22_X1 U14213 ( .A1(n13069), .A2(n13114), .B1(n11507), .B2(n13096), .ZN(
        n11509) );
  OAI211_X1 U14214 ( .C1(n11657), .C2(n13072), .A(n11509), .B(n11508), .ZN(
        n11510) );
  AOI21_X1 U14215 ( .B1(n11511), .B2(n13090), .A(n11510), .ZN(n11512) );
  OAI21_X1 U14216 ( .B1(n11513), .B2(n13098), .A(n11512), .ZN(P3_U3170) );
  NAND2_X1 U14217 ( .A1(n15642), .A2(n11514), .ZN(n11515) );
  INV_X1 U14218 ( .A(n11518), .ZN(n11516) );
  AOI21_X1 U14219 ( .B1(n11516), .B2(n13977), .A(n13726), .ZN(n11517) );
  AOI21_X1 U14220 ( .B1(n11597), .B2(n11518), .A(n11517), .ZN(n11519) );
  INV_X1 U14221 ( .A(n13732), .ZN(n13905) );
  XNOR2_X1 U14222 ( .A(n11519), .B(n13905), .ZN(n15643) );
  INV_X1 U14223 ( .A(n11539), .ZN(n11523) );
  AOI211_X1 U14224 ( .C1(n11521), .C2(n13907), .A(n11520), .B(n13732), .ZN(
        n11522) );
  OAI21_X1 U14225 ( .B1(n11523), .B2(n11522), .A(n14307), .ZN(n11525) );
  AND2_X1 U14226 ( .A1(n11525), .A2(n11524), .ZN(n15639) );
  MUX2_X1 U14227 ( .A(n11526), .B(n15639), .S(n14293), .Z(n11534) );
  OAI211_X1 U14228 ( .C1(n11527), .C2(n15641), .A(n11543), .B(n14239), .ZN(
        n15638) );
  INV_X1 U14229 ( .A(n15638), .ZN(n11532) );
  AND2_X2 U14230 ( .A1(n14293), .A2(n11528), .ZN(n14282) );
  OAI22_X1 U14231 ( .A1(n14275), .A2(n15641), .B1(n14290), .B2(n11530), .ZN(
        n11531) );
  AOI21_X1 U14232 ( .B1(n11532), .B2(n14282), .A(n11531), .ZN(n11533) );
  OAI211_X1 U14233 ( .C1(n14279), .C2(n15643), .A(n11534), .B(n11533), .ZN(
        P2_U3259) );
  OAI21_X1 U14234 ( .B1(n11536), .B2(n13738), .A(n11535), .ZN(n15654) );
  NAND3_X1 U14235 ( .A1(n11539), .A2(n13738), .A3(n11538), .ZN(n11540) );
  NAND2_X1 U14236 ( .A1(n11537), .A2(n11540), .ZN(n11541) );
  AOI222_X1 U14237 ( .A1(n14307), .A2(n11541), .B1(n13974), .B2(n14304), .C1(
        n13976), .C2(n14302), .ZN(n15653) );
  MUX2_X1 U14238 ( .A(n11542), .B(n15653), .S(n14293), .Z(n11549) );
  AOI21_X1 U14239 ( .B1(n11543), .B2(n15650), .A(n8582), .ZN(n11544) );
  AND2_X1 U14240 ( .A1(n11544), .A2(n11557), .ZN(n15649) );
  INV_X1 U14241 ( .A(n15650), .ZN(n11546) );
  OAI22_X1 U14242 ( .A1(n14275), .A2(n11546), .B1(n11545), .B2(n14290), .ZN(
        n11547) );
  AOI21_X1 U14243 ( .B1(n15649), .B2(n14282), .A(n11547), .ZN(n11548) );
  OAI211_X1 U14244 ( .C1(n14279), .C2(n15654), .A(n11549), .B(n11548), .ZN(
        P2_U3258) );
  NAND2_X1 U14245 ( .A1(n11550), .A2(n7327), .ZN(n11862) );
  OR2_X1 U14246 ( .A1(n11550), .A2(n7327), .ZN(n11551) );
  NAND2_X1 U14247 ( .A1(n11862), .A2(n11551), .ZN(n11579) );
  NAND3_X1 U14248 ( .A1(n11537), .A2(n7327), .A3(n11553), .ZN(n11554) );
  NAND2_X1 U14249 ( .A1(n11552), .A2(n11554), .ZN(n11555) );
  AOI222_X1 U14250 ( .A1(n14307), .A2(n11555), .B1(n13973), .B2(n14304), .C1(
        n13975), .C2(n14302), .ZN(n11572) );
  MUX2_X1 U14251 ( .A(n11556), .B(n11572), .S(n14293), .Z(n11563) );
  INV_X1 U14252 ( .A(n11557), .ZN(n11558) );
  OAI211_X1 U14253 ( .C1(n7843), .C2(n11558), .A(n7845), .B(n14239), .ZN(
        n11571) );
  INV_X1 U14254 ( .A(n11571), .ZN(n11561) );
  OAI22_X1 U14255 ( .A1(n14275), .A2(n7843), .B1(n14290), .B2(n11559), .ZN(
        n11560) );
  AOI21_X1 U14256 ( .B1(n11561), .B2(n14282), .A(n11560), .ZN(n11562) );
  OAI211_X1 U14257 ( .C1(n14279), .C2(n11579), .A(n11563), .B(n11562), .ZN(
        P2_U3257) );
  MUX2_X1 U14258 ( .A(n11565), .B(n11564), .S(n14293), .Z(n11569) );
  OAI22_X1 U14259 ( .A1(n14275), .A2(n13769), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14290), .ZN(n11566) );
  AOI21_X1 U14260 ( .B1(n14282), .B2(n11567), .A(n11566), .ZN(n11568) );
  OAI211_X1 U14261 ( .C1(n11570), .C2(n14265), .A(n11569), .B(n11568), .ZN(
        P2_U3262) );
  NAND2_X1 U14262 ( .A1(n11572), .A2(n11571), .ZN(n11575) );
  NAND2_X1 U14263 ( .A1(n11575), .A2(n15659), .ZN(n11574) );
  AOI22_X1 U14264 ( .A1(n9618), .A2(n13789), .B1(P2_REG0_REG_8__SCAN_IN), .B2(
        n15657), .ZN(n11573) );
  OAI211_X1 U14265 ( .C1(n11579), .C2(n14461), .A(n11574), .B(n11573), .ZN(
        P2_U3454) );
  NAND2_X1 U14266 ( .A1(n11575), .A2(n15670), .ZN(n11578) );
  INV_X1 U14267 ( .A(n14400), .ZN(n11576) );
  AOI22_X1 U14268 ( .A1(n11576), .A2(n13789), .B1(P2_REG1_REG_8__SCAN_IN), 
        .B2(n15667), .ZN(n11577) );
  OAI211_X1 U14269 ( .C1(n11579), .C2(n14401), .A(n11578), .B(n11577), .ZN(
        P2_U3507) );
  MUX2_X1 U14270 ( .A(n11581), .B(n11580), .S(n14293), .Z(n11587) );
  INV_X1 U14271 ( .A(n11582), .ZN(n11583) );
  OAI22_X1 U14272 ( .A1(n14275), .A2(n13727), .B1(n14290), .B2(n11583), .ZN(
        n11584) );
  AOI21_X1 U14273 ( .B1(n11585), .B2(n14282), .A(n11584), .ZN(n11586) );
  OAI211_X1 U14274 ( .C1(n14279), .C2(n11588), .A(n11587), .B(n11586), .ZN(
        P2_U3260) );
  NOR2_X1 U14275 ( .A1(n11590), .A2(n11589), .ZN(n11591) );
  XNOR2_X1 U14276 ( .A(n11591), .B(n13908), .ZN(n11602) );
  INV_X1 U14277 ( .A(n11602), .ZN(n15635) );
  INV_X1 U14278 ( .A(n13908), .ZN(n11593) );
  NAND3_X1 U14279 ( .A1(n11594), .A2(n11593), .A3(n11592), .ZN(n11595) );
  AOI21_X1 U14280 ( .B1(n11596), .B2(n11595), .A(n14217), .ZN(n11600) );
  OAI22_X1 U14281 ( .A1(n11598), .A2(n14116), .B1(n11597), .B2(n14118), .ZN(
        n11599) );
  AOI211_X1 U14282 ( .C1(n11602), .C2(n11601), .A(n11600), .B(n11599), .ZN(
        n15634) );
  MUX2_X1 U14283 ( .A(n11603), .B(n15634), .S(n14293), .Z(n11610) );
  INV_X1 U14284 ( .A(n11604), .ZN(n11605) );
  AOI211_X1 U14285 ( .C1(n15632), .C2(n11606), .A(n8582), .B(n11605), .ZN(
        n15631) );
  OAI22_X1 U14286 ( .A1(n14275), .A2(n13733), .B1(n11607), .B2(n14290), .ZN(
        n11608) );
  AOI21_X1 U14287 ( .B1(n15631), .B2(n14282), .A(n11608), .ZN(n11609) );
  OAI211_X1 U14288 ( .C1(n15635), .C2(n14265), .A(n11610), .B(n11609), .ZN(
        P2_U3261) );
  INV_X1 U14289 ( .A(n11611), .ZN(n11614) );
  OAI222_X1 U14290 ( .A1(n15232), .A2(n7719), .B1(n15236), .B2(n11614), .C1(
        n11612), .C2(n6537), .ZN(P1_U3331) );
  OAI222_X1 U14291 ( .A1(n11615), .A2(P2_U3088), .B1(n10996), .B2(n11614), 
        .C1(n11613), .C2(n14478), .ZN(P2_U3303) );
  OAI22_X1 U14292 ( .A1(n11617), .A2(n11616), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n11618), .ZN(n15572) );
  XNOR2_X1 U14293 ( .A(n15566), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n15573) );
  NOR2_X1 U14294 ( .A1(n15572), .A2(n15573), .ZN(n15571) );
  XNOR2_X1 U14295 ( .A(n12157), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n12163) );
  XNOR2_X1 U14296 ( .A(n12164), .B(n12163), .ZN(n11628) );
  NAND2_X1 U14297 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n13572)
         );
  OR2_X1 U14298 ( .A1(n11618), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11619) );
  INV_X1 U14299 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11621) );
  MUX2_X1 U14300 ( .A(n11621), .B(P2_REG2_REG_13__SCAN_IN), .S(n15566), .Z(
        n15567) );
  NAND2_X1 U14301 ( .A1(n15566), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11622) );
  NAND2_X1 U14302 ( .A1(n15569), .A2(n11622), .ZN(n12158) );
  XOR2_X1 U14303 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n12156), .Z(n11623) );
  NAND2_X1 U14304 ( .A1(n15603), .A2(n11623), .ZN(n11624) );
  NAND2_X1 U14305 ( .A1(n13572), .A2(n11624), .ZN(n11626) );
  INV_X1 U14306 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15274) );
  NOR2_X1 U14307 ( .A1(n15609), .A2(n15274), .ZN(n11625) );
  AOI211_X1 U14308 ( .C1(n15595), .C2(n12157), .A(n11626), .B(n11625), .ZN(
        n11627) );
  OAI21_X1 U14309 ( .B1(n11628), .B2(n15586), .A(n11627), .ZN(P2_U3228) );
  AOI21_X1 U14310 ( .B1(n11630), .B2(n11629), .A(n11641), .ZN(n11638) );
  OAI22_X1 U14311 ( .A1(n11632), .A2(n13093), .B1(n13081), .B2(n11631), .ZN(
        n11633) );
  AOI211_X1 U14312 ( .C1(n13089), .C2(n13111), .A(n11634), .B(n11633), .ZN(
        n11637) );
  NAND2_X1 U14313 ( .A1(n13090), .A2(n11635), .ZN(n11636) );
  OAI211_X1 U14314 ( .C1(n11638), .C2(n13098), .A(n11637), .B(n11636), .ZN(
        P3_U3167) );
  INV_X1 U14315 ( .A(n11639), .ZN(n11640) );
  NOR2_X1 U14316 ( .A1(n11641), .A2(n11640), .ZN(n11655) );
  XNOR2_X1 U14317 ( .A(n11642), .B(n11645), .ZN(n11654) );
  NAND2_X1 U14318 ( .A1(n11655), .A2(n11654), .ZN(n11653) );
  NAND2_X1 U14319 ( .A1(n11653), .A2(n11643), .ZN(n11812) );
  XNOR2_X1 U14320 ( .A(n11812), .B(n11811), .ZN(n11651) );
  OAI22_X1 U14321 ( .A1(n11645), .A2(n13093), .B1(n13081), .B2(n11644), .ZN(
        n11646) );
  AOI211_X1 U14322 ( .C1(n13089), .C2(n13109), .A(n11647), .B(n11646), .ZN(
        n11650) );
  NAND2_X1 U14323 ( .A1(n13090), .A2(n11648), .ZN(n11649) );
  OAI211_X1 U14324 ( .C1(n11651), .C2(n13098), .A(n11650), .B(n11649), .ZN(
        P3_U3153) );
  INV_X1 U14325 ( .A(n11652), .ZN(n11662) );
  OAI211_X1 U14326 ( .C1(n11655), .C2(n11654), .A(n11653), .B(n13058), .ZN(
        n11660) );
  AND2_X1 U14327 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n13145) );
  OAI22_X1 U14328 ( .A1(n11657), .A2(n13093), .B1(n13081), .B2(n11656), .ZN(
        n11658) );
  AOI211_X1 U14329 ( .C1(n13089), .C2(n13110), .A(n13145), .B(n11658), .ZN(
        n11659) );
  OAI211_X1 U14330 ( .C1(n11662), .C2(n11661), .A(n11660), .B(n11659), .ZN(
        P3_U3179) );
  NAND2_X1 U14331 ( .A1(n11664), .A2(n11663), .ZN(n12971) );
  INV_X1 U14332 ( .A(n11665), .ZN(n11666) );
  INV_X1 U14333 ( .A(n15410), .ZN(n12039) );
  NAND2_X1 U14334 ( .A1(n11669), .A2(n15410), .ZN(n12565) );
  NAND2_X1 U14335 ( .A1(n12566), .A2(n12565), .ZN(n12049) );
  NAND2_X1 U14336 ( .A1(n12049), .A2(n12050), .ZN(n11671) );
  NAND2_X1 U14337 ( .A1(n12813), .A2(n15410), .ZN(n11670) );
  NAND2_X1 U14338 ( .A1(n11671), .A2(n11670), .ZN(n15385) );
  INV_X1 U14339 ( .A(n15386), .ZN(n15384) );
  NAND2_X1 U14340 ( .A1(n15385), .A2(n15384), .ZN(n11673) );
  NAND2_X1 U14341 ( .A1(n12570), .A2(n15418), .ZN(n11672) );
  NAND2_X1 U14342 ( .A1(n11673), .A2(n11672), .ZN(n11718) );
  INV_X1 U14343 ( .A(n12753), .ZN(n11723) );
  NAND2_X1 U14344 ( .A1(n11718), .A2(n11723), .ZN(n11676) );
  NAND2_X1 U14345 ( .A1(n12812), .A2(n11674), .ZN(n11675) );
  NAND2_X1 U14346 ( .A1(n12581), .A2(n15427), .ZN(n12062) );
  NAND2_X1 U14347 ( .A1(n15434), .A2(n11687), .ZN(n11677) );
  AND2_X1 U14348 ( .A1(n12062), .A2(n11677), .ZN(n15349) );
  NAND2_X1 U14349 ( .A1(n15350), .A2(n15349), .ZN(n11681) );
  XNOR2_X1 U14350 ( .A(n15440), .B(n12591), .ZN(n12751) );
  INV_X1 U14351 ( .A(n11677), .ZN(n11679) );
  INV_X1 U14352 ( .A(n12754), .ZN(n11678) );
  OR2_X1 U14353 ( .A1(n11679), .A2(n11678), .ZN(n15351) );
  NAND2_X1 U14354 ( .A1(n15440), .A2(n12591), .ZN(n11682) );
  XNOR2_X1 U14355 ( .A(n12598), .B(n14645), .ZN(n11705) );
  XNOR2_X1 U14356 ( .A(n11704), .B(n11705), .ZN(n15445) );
  NAND2_X1 U14357 ( .A1(n12562), .A2(n12565), .ZN(n11684) );
  NAND2_X1 U14358 ( .A1(n11684), .A2(n12566), .ZN(n15387) );
  NAND2_X1 U14359 ( .A1(n15386), .A2(n15387), .ZN(n11686) );
  NAND2_X1 U14360 ( .A1(n12570), .A2(n15399), .ZN(n11685) );
  INV_X1 U14361 ( .A(n11674), .ZN(n11721) );
  NAND2_X1 U14362 ( .A1(n11721), .A2(n12812), .ZN(n12577) );
  NAND2_X1 U14363 ( .A1(n12586), .A2(n11687), .ZN(n11688) );
  INV_X1 U14364 ( .A(n15440), .ZN(n12590) );
  XNOR2_X1 U14365 ( .A(n11706), .B(n12748), .ZN(n11690) );
  OAI21_X1 U14366 ( .B1(n11690), .B2(n15355), .A(n11689), .ZN(n15451) );
  INV_X1 U14367 ( .A(n15451), .ZN(n11691) );
  MUX2_X1 U14368 ( .A(n11692), .B(n11691), .S(n15005), .Z(n11703) );
  INV_X1 U14369 ( .A(n14935), .ZN(n15400) );
  AND2_X1 U14370 ( .A1(n15410), .A2(n11693), .ZN(n12037) );
  NAND2_X1 U14371 ( .A1(n15396), .A2(n11674), .ZN(n15375) );
  XNOR2_X1 U14372 ( .A(n15362), .B(n12598), .ZN(n11694) );
  NOR2_X1 U14373 ( .A1(n11694), .A2(n15397), .ZN(n15449) );
  OR2_X1 U14374 ( .A1(n11695), .A2(n12558), .ZN(n12786) );
  INV_X1 U14375 ( .A(n12786), .ZN(n11696) );
  NAND2_X1 U14376 ( .A1(n11697), .A2(n11696), .ZN(n11698) );
  INV_X1 U14377 ( .A(n12598), .ZN(n12596) );
  INV_X1 U14378 ( .A(n11699), .ZN(n11700) );
  OAI22_X1 U14379 ( .A1(n15394), .A2(n12596), .B1(n11700), .B2(n14985), .ZN(
        n11701) );
  AOI21_X1 U14380 ( .B1(n15400), .B2(n15449), .A(n11701), .ZN(n11702) );
  OAI211_X1 U14381 ( .C1(n15060), .C2(n15445), .A(n11703), .B(n11702), .ZN(
        P1_U3286) );
  XNOR2_X1 U14382 ( .A(n12607), .B(n12606), .ZN(n12756) );
  XOR2_X1 U14383 ( .A(n11732), .B(n12756), .Z(n15457) );
  NAND2_X1 U14384 ( .A1(n12598), .A2(n12597), .ZN(n11707) );
  XOR2_X1 U14385 ( .A(n12756), .B(n11735), .Z(n11710) );
  INV_X2 U14386 ( .A(n15355), .ZN(n15389) );
  AOI22_X1 U14387 ( .A1(n15029), .A2(n14645), .B1(n14643), .B2(n15031), .ZN(
        n11826) );
  INV_X1 U14388 ( .A(n11826), .ZN(n11709) );
  AOI21_X1 U14389 ( .B1(n11710), .B2(n15389), .A(n11709), .ZN(n15458) );
  MUX2_X1 U14390 ( .A(n11711), .B(n15458), .S(n15005), .Z(n11717) );
  OR2_X1 U14391 ( .A1(n15362), .A2(n12598), .ZN(n11713) );
  OR2_X1 U14392 ( .A1(n12607), .A2(n12598), .ZN(n11712) );
  AOI211_X1 U14393 ( .C1(n12607), .C2(n11713), .A(n15397), .B(n11742), .ZN(
        n15453) );
  INV_X1 U14394 ( .A(n12607), .ZN(n12605) );
  INV_X1 U14395 ( .A(n11829), .ZN(n11714) );
  OAI22_X1 U14396 ( .A1(n15394), .A2(n12605), .B1(n11714), .B2(n14985), .ZN(
        n11715) );
  AOI21_X1 U14397 ( .B1(n15453), .B2(n15400), .A(n11715), .ZN(n11716) );
  OAI211_X1 U14398 ( .C1(n15060), .C2(n15457), .A(n11717), .B(n11716), .ZN(
        P1_U3285) );
  XNOR2_X1 U14399 ( .A(n11718), .B(n12753), .ZN(n15421) );
  OAI211_X1 U14400 ( .C1(n15396), .C2(n11674), .A(n15377), .B(n15375), .ZN(
        n15422) );
  AOI22_X1 U14401 ( .A1(n15405), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n15392), 
        .B2(n8894), .ZN(n11719) );
  OAI21_X1 U14402 ( .B1(n14935), .B2(n15422), .A(n11719), .ZN(n11720) );
  AOI21_X1 U14403 ( .B1(n14954), .B2(n11721), .A(n11720), .ZN(n11727) );
  XNOR2_X1 U14404 ( .A(n11723), .B(n11722), .ZN(n11725) );
  OAI21_X1 U14405 ( .B1(n11725), .B2(n15355), .A(n11724), .ZN(n15424) );
  NAND2_X1 U14406 ( .A1(n15005), .A2(n15424), .ZN(n11726) );
  OAI211_X1 U14407 ( .C1(n15060), .C2(n15421), .A(n11727), .B(n11726), .ZN(
        P1_U3290) );
  NAND2_X1 U14408 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  OAI211_X1 U14409 ( .C1(n11731), .C2(n13550), .A(n11730), .B(n12535), .ZN(
        P3_U3272) );
  OR2_X1 U14410 ( .A1(n12607), .A2(n14644), .ZN(n11733) );
  INV_X1 U14411 ( .A(n14643), .ZN(n12602) );
  XNOR2_X1 U14412 ( .A(n12603), .B(n12602), .ZN(n11832) );
  XNOR2_X1 U14413 ( .A(n11833), .B(n11832), .ZN(n15467) );
  INV_X1 U14414 ( .A(n15467), .ZN(n11748) );
  OR2_X1 U14415 ( .A1(n12607), .A2(n12606), .ZN(n11736) );
  INV_X1 U14416 ( .A(n11832), .ZN(n12761) );
  OAI21_X1 U14417 ( .B1(n6708), .B2(n12761), .A(n11838), .ZN(n11740) );
  NAND2_X1 U14418 ( .A1(n14642), .A2(n15031), .ZN(n11739) );
  NAND2_X1 U14419 ( .A1(n14644), .A2(n15029), .ZN(n11738) );
  NAND2_X1 U14420 ( .A1(n11739), .A2(n11738), .ZN(n11920) );
  AOI21_X1 U14421 ( .B1(n11740), .B2(n15389), .A(n11920), .ZN(n15465) );
  MUX2_X1 U14422 ( .A(n11741), .B(n15465), .S(n15005), .Z(n11747) );
  INV_X1 U14423 ( .A(n12603), .ZN(n12601) );
  OAI211_X1 U14424 ( .C1(n11742), .C2(n12601), .A(n12077), .B(n15377), .ZN(
        n15463) );
  INV_X1 U14425 ( .A(n15463), .ZN(n11745) );
  INV_X1 U14426 ( .A(n11918), .ZN(n11743) );
  OAI22_X1 U14427 ( .A1(n15394), .A2(n12601), .B1(n14985), .B2(n11743), .ZN(
        n11744) );
  AOI21_X1 U14428 ( .B1(n11745), .B2(n15400), .A(n11744), .ZN(n11746) );
  OAI211_X1 U14429 ( .C1(n15060), .C2(n11748), .A(n11747), .B(n11746), .ZN(
        P1_U3284) );
  NAND2_X1 U14430 ( .A1(n11749), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11754) );
  INV_X1 U14431 ( .A(n11750), .ZN(n11752) );
  NAND2_X1 U14432 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  NAND2_X1 U14433 ( .A1(n11765), .A2(n11764), .ZN(n11758) );
  XNOR2_X1 U14434 ( .A(n11758), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n11759) );
  INV_X1 U14435 ( .A(n11759), .ZN(n11760) );
  INV_X1 U14436 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14766) );
  XNOR2_X1 U14437 ( .A(n14766), .B(P3_ADDR_REG_11__SCAN_IN), .ZN(n12097) );
  INV_X1 U14438 ( .A(n12097), .ZN(n11766) );
  XNOR2_X1 U14439 ( .A(n12098), .B(n11766), .ZN(n11767) );
  NAND2_X1 U14440 ( .A1(n12096), .A2(n12095), .ZN(n11768) );
  XNOR2_X1 U14441 ( .A(n11768), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  INV_X1 U14442 ( .A(n11769), .ZN(n11773) );
  OAI222_X1 U14443 ( .A1(n11771), .A2(P2_U3088), .B1(n10996), .B2(n11773), 
        .C1(n11770), .C2(n14478), .ZN(P2_U3302) );
  OAI222_X1 U14444 ( .A1(n15232), .A2(n11774), .B1(n15236), .B2(n11773), .C1(
        n11772), .C2(P1_U3086), .ZN(P1_U3330) );
  XNOR2_X1 U14445 ( .A(n11776), .B(n11775), .ZN(n11783) );
  INV_X1 U14446 ( .A(n11777), .ZN(n14291) );
  OAI22_X1 U14447 ( .A1(n11778), .A2(n13587), .B1(n13717), .B2(n14291), .ZN(
        n11779) );
  AOI211_X1 U14448 ( .C1(n13675), .C2(n14305), .A(n11780), .B(n11779), .ZN(
        n11782) );
  NAND2_X1 U14449 ( .A1(n13693), .A2(n14399), .ZN(n11781) );
  OAI211_X1 U14450 ( .C1(n11783), .C2(n13695), .A(n11782), .B(n11781), .ZN(
        P2_U3208) );
  OAI21_X1 U14451 ( .B1(n11785), .B2(n11784), .A(n11899), .ZN(n11786) );
  NAND2_X1 U14452 ( .A1(n11786), .A2(n13058), .ZN(n11792) );
  AOI21_X1 U14453 ( .B1(n13069), .B2(n13109), .A(n11787), .ZN(n11788) );
  OAI21_X1 U14454 ( .B1(n12242), .B2(n13072), .A(n11788), .ZN(n11789) );
  AOI21_X1 U14455 ( .B1(n11790), .B2(n13090), .A(n11789), .ZN(n11791) );
  OAI211_X1 U14456 ( .C1(n13081), .C2(n11793), .A(n11792), .B(n11791), .ZN(
        P3_U3171) );
  NAND2_X1 U14457 ( .A1(n11802), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11798) );
  NAND2_X1 U14458 ( .A1(n11799), .A2(n11798), .ZN(n11796) );
  INV_X1 U14459 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11794) );
  MUX2_X1 U14460 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n11794), .S(n14781), .Z(
        n11795) );
  NAND2_X1 U14461 ( .A1(n11796), .A2(n11795), .ZN(n14778) );
  MUX2_X1 U14462 ( .A(n11794), .B(P1_REG2_REG_17__SCAN_IN), .S(n14781), .Z(
        n11797) );
  NAND3_X1 U14463 ( .A1(n11799), .A2(n11798), .A3(n11797), .ZN(n11800) );
  NAND3_X1 U14464 ( .A1(n14778), .A2(n15338), .A3(n11800), .ZN(n11809) );
  NAND2_X1 U14465 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14553)
         );
  XNOR2_X1 U14466 ( .A(n14781), .B(n11801), .ZN(n14779) );
  NAND2_X1 U14467 ( .A1(n11802), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11803) );
  NAND2_X1 U14468 ( .A1(n11804), .A2(n11803), .ZN(n14780) );
  XOR2_X1 U14469 ( .A(n14779), .B(n14780), .Z(n11805) );
  NAND2_X1 U14470 ( .A1(n15332), .A2(n11805), .ZN(n11806) );
  NAND2_X1 U14471 ( .A1(n14553), .A2(n11806), .ZN(n11807) );
  AOI21_X1 U14472 ( .B1(n15342), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11807), 
        .ZN(n11808) );
  OAI211_X1 U14473 ( .C1(n14804), .C2(n11810), .A(n11809), .B(n11808), .ZN(
        P1_U3260) );
  MUX2_X1 U14474 ( .A(n13110), .B(n11812), .S(n11811), .Z(n11813) );
  XOR2_X1 U14475 ( .A(n11814), .B(n11813), .Z(n11823) );
  NAND2_X1 U14476 ( .A1(n13089), .A2(n13108), .ZN(n11816) );
  OAI211_X1 U14477 ( .C1(n11817), .C2(n13093), .A(n11816), .B(n11815), .ZN(
        n11818) );
  AOI21_X1 U14478 ( .B1(n11819), .B2(n13096), .A(n11818), .ZN(n11822) );
  NAND2_X1 U14479 ( .A1(n13090), .A2(n11820), .ZN(n11821) );
  OAI211_X1 U14480 ( .C1(n11823), .C2(n13098), .A(n11822), .B(n11821), .ZN(
        P3_U3161) );
  OR2_X1 U14481 ( .A1(n11886), .A2(n11825), .ZN(n11912) );
  INV_X1 U14482 ( .A(n11912), .ZN(n11824) );
  AOI21_X1 U14483 ( .B1(n11825), .B2(n11886), .A(n11824), .ZN(n11831) );
  NAND2_X1 U14484 ( .A1(n12607), .A2(n15189), .ZN(n15455) );
  NOR2_X1 U14485 ( .A1(n11923), .A2(n15455), .ZN(n11828) );
  NAND2_X1 U14486 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n14743) );
  OAI21_X1 U14487 ( .B1(n14628), .B2(n11826), .A(n14743), .ZN(n11827) );
  AOI211_X1 U14488 ( .C1(n14630), .C2(n11829), .A(n11828), .B(n11827), .ZN(
        n11830) );
  OAI21_X1 U14489 ( .B1(n11831), .B2(n14619), .A(n11830), .ZN(P1_U3221) );
  OR2_X1 U14490 ( .A1(n12603), .A2(n14643), .ZN(n11834) );
  INV_X1 U14491 ( .A(n14642), .ZN(n12599) );
  NAND2_X1 U14492 ( .A1(n12600), .A2(n12599), .ZN(n11835) );
  NAND2_X1 U14493 ( .A1(n11933), .A2(n11835), .ZN(n12749) );
  OR2_X1 U14494 ( .A1(n12600), .A2(n14642), .ZN(n11985) );
  NAND2_X1 U14495 ( .A1(n11992), .A2(n11985), .ZN(n11927) );
  XNOR2_X1 U14496 ( .A(n12619), .B(n14641), .ZN(n12758) );
  XNOR2_X1 U14497 ( .A(n11927), .B(n11989), .ZN(n12123) );
  INV_X1 U14498 ( .A(n12619), .ZN(n12617) );
  OAI21_X1 U14499 ( .B1(n12077), .B2(n12600), .A(n12619), .ZN(n11836) );
  NAND3_X1 U14500 ( .A1(n11836), .A2(n15377), .A3(n11945), .ZN(n12119) );
  OAI21_X1 U14501 ( .B1(n12617), .B2(n15471), .A(n12119), .ZN(n11844) );
  NAND2_X1 U14502 ( .A1(n12603), .A2(n12602), .ZN(n11837) );
  NAND2_X1 U14503 ( .A1(n11973), .A2(n11933), .ZN(n11839) );
  NAND2_X1 U14504 ( .A1(n11839), .A2(n12758), .ZN(n11930) );
  NAND3_X1 U14505 ( .A1(n11973), .A2(n11989), .A3(n11933), .ZN(n11840) );
  NAND3_X1 U14506 ( .A1(n11930), .A2(n15389), .A3(n11840), .ZN(n11843) );
  NAND2_X1 U14507 ( .A1(n14640), .A2(n15031), .ZN(n11842) );
  NAND2_X1 U14508 ( .A1(n14642), .A2(n15029), .ZN(n11841) );
  AND2_X1 U14509 ( .A1(n11842), .A2(n11841), .ZN(n12023) );
  NAND2_X1 U14510 ( .A1(n11843), .A2(n12023), .ZN(n12120) );
  AOI211_X1 U14511 ( .C1(n12123), .C2(n15476), .A(n11844), .B(n12120), .ZN(
        n11847) );
  NAND2_X1 U14512 ( .A1(n7301), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11845) );
  OAI21_X1 U14513 ( .B1(n11847), .B2(n7301), .A(n11845), .ZN(P1_U3539) );
  NAND2_X1 U14514 ( .A1(n15477), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11846) );
  OAI21_X1 U14515 ( .B1(n11847), .B2(n15477), .A(n11846), .ZN(P1_U3492) );
  XOR2_X1 U14516 ( .A(n11848), .B(n12502), .Z(n11860) );
  XOR2_X1 U14517 ( .A(n11849), .B(n12502), .Z(n11850) );
  INV_X1 U14518 ( .A(n13396), .ZN(n13433) );
  OAI222_X1 U14519 ( .A1(n11850), .A2(n13428), .B1(n13433), .B2(n12300), .C1(
        n13431), .C2(n12209), .ZN(n11858) );
  OAI22_X1 U14520 ( .A1(n12420), .A2(n13482), .B1(n13486), .B2(n15738), .ZN(
        n11851) );
  AOI21_X1 U14521 ( .B1(n11858), .B2(n13486), .A(n11851), .ZN(n11852) );
  OAI21_X1 U14522 ( .B1(n13488), .B2(n11860), .A(n11852), .ZN(P3_U3472) );
  AOI22_X1 U14523 ( .A1(n15688), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15675), 
        .B2(n12211), .ZN(n11853) );
  OAI21_X1 U14524 ( .B1(n12420), .B2(n13403), .A(n11853), .ZN(n11854) );
  AOI21_X1 U14525 ( .B1(n11858), .B2(n13405), .A(n11854), .ZN(n11855) );
  OAI21_X1 U14526 ( .B1(n13441), .B2(n11860), .A(n11855), .ZN(P3_U3220) );
  INV_X1 U14527 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n11856) );
  OAI22_X1 U14528 ( .A1(n12420), .A2(n13536), .B1(n11856), .B2(n15691), .ZN(
        n11857) );
  AOI21_X1 U14529 ( .B1(n11858), .B2(n15691), .A(n11857), .ZN(n11859) );
  OAI21_X1 U14530 ( .B1(n13540), .B2(n11860), .A(n11859), .ZN(P3_U3429) );
  NAND2_X1 U14531 ( .A1(n11862), .A2(n11861), .ZN(n11863) );
  XNOR2_X1 U14532 ( .A(n11863), .B(n7321), .ZN(n12054) );
  INV_X1 U14533 ( .A(n11956), .ZN(n11866) );
  AND3_X1 U14534 ( .A1(n11552), .A2(n7321), .A3(n11864), .ZN(n11865) );
  OAI21_X1 U14535 ( .B1(n11866), .B2(n11865), .A(n14307), .ZN(n11868) );
  AOI22_X1 U14536 ( .A1(n14302), .A2(n13974), .B1(n14303), .B2(n14304), .ZN(
        n11867) );
  OAI211_X1 U14537 ( .C1(n12054), .C2(n15642), .A(n11868), .B(n11867), .ZN(
        n12055) );
  INV_X1 U14538 ( .A(n12055), .ZN(n11869) );
  MUX2_X1 U14539 ( .A(n11870), .B(n11869), .S(n14293), .Z(n11878) );
  OAI21_X1 U14540 ( .B1(n11871), .B2(n12061), .A(n14239), .ZN(n11873) );
  NOR2_X1 U14541 ( .A1(n11873), .A2(n11872), .ZN(n12056) );
  INV_X1 U14542 ( .A(n11874), .ZN(n11875) );
  OAI22_X1 U14543 ( .A1(n14275), .A2(n12061), .B1(n14290), .B2(n11875), .ZN(
        n11876) );
  AOI21_X1 U14544 ( .B1(n12056), .B2(n14282), .A(n11876), .ZN(n11877) );
  OAI211_X1 U14545 ( .C1(n12054), .C2(n14265), .A(n11878), .B(n11877), .ZN(
        P2_U3256) );
  NAND2_X1 U14546 ( .A1(n15005), .A2(n15389), .ZN(n14938) );
  INV_X1 U14547 ( .A(n14938), .ZN(n14983) );
  NOR2_X1 U14548 ( .A1(n14983), .A2(n15381), .ZN(n11884) );
  INV_X1 U14549 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11879) );
  OAI22_X1 U14550 ( .A1(n15405), .A2(n11880), .B1(n11879), .B2(n14985), .ZN(
        n11881) );
  AOI21_X1 U14551 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n15405), .A(n11881), .ZN(
        n11883) );
  NOR2_X1 U14552 ( .A1(n14935), .A2(n15397), .ZN(n12989) );
  OAI21_X1 U14553 ( .B1(n14954), .B2(n12989), .A(n12038), .ZN(n11882) );
  OAI211_X1 U14554 ( .C1(n11884), .C2(n12750), .A(n11883), .B(n11882), .ZN(
        P1_U3293) );
  INV_X1 U14555 ( .A(n12600), .ZN(n15472) );
  OR2_X1 U14556 ( .A1(n11886), .A2(n11885), .ZN(n11914) );
  NAND2_X1 U14557 ( .A1(n11914), .A2(n11887), .ZN(n11889) );
  AOI21_X1 U14558 ( .B1(n11889), .B2(n11888), .A(n14619), .ZN(n11892) );
  NAND2_X1 U14559 ( .A1(n11914), .A2(n11890), .ZN(n11891) );
  NAND2_X1 U14560 ( .A1(n11892), .A2(n11891), .ZN(n11897) );
  INV_X1 U14561 ( .A(n11893), .ZN(n12076) );
  OAI22_X1 U14562 ( .A1(n14609), .A2(n12602), .B1(n12076), .B2(n14611), .ZN(
        n11894) );
  AOI211_X1 U14563 ( .C1(n14591), .C2(n14641), .A(n11895), .B(n11894), .ZN(
        n11896) );
  OAI211_X1 U14564 ( .C1(n15472), .C2(n14633), .A(n11897), .B(n11896), .ZN(
        P1_U3217) );
  AND2_X1 U14565 ( .A1(n11899), .A2(n11898), .ZN(n11902) );
  OAI211_X1 U14566 ( .C1(n11902), .C2(n11901), .A(n13058), .B(n11900), .ZN(
        n11909) );
  NAND2_X1 U14567 ( .A1(n13089), .A2(n13106), .ZN(n11904) );
  OAI211_X1 U14568 ( .C1(n11905), .C2(n13093), .A(n11904), .B(n11903), .ZN(
        n11906) );
  AOI21_X1 U14569 ( .B1(n11907), .B2(n13090), .A(n11906), .ZN(n11908) );
  OAI211_X1 U14570 ( .C1(n13081), .C2(n11910), .A(n11909), .B(n11908), .ZN(
        P3_U3157) );
  NAND2_X1 U14571 ( .A1(n11912), .A2(n11911), .ZN(n11916) );
  AND2_X1 U14572 ( .A1(n11914), .A2(n11913), .ZN(n11915) );
  OAI21_X1 U14573 ( .B1(n11917), .B2(n11916), .A(n11915), .ZN(n11925) );
  NAND2_X1 U14574 ( .A1(n12603), .A2(n15189), .ZN(n15464) );
  NAND2_X1 U14575 ( .A1(n14630), .A2(n11918), .ZN(n11922) );
  AOI21_X1 U14576 ( .B1(n14571), .B2(n11920), .A(n11919), .ZN(n11921) );
  OAI211_X1 U14577 ( .C1(n15464), .C2(n11923), .A(n11922), .B(n11921), .ZN(
        n11924) );
  AOI21_X1 U14578 ( .B1(n11925), .B2(n14621), .A(n11924), .ZN(n11926) );
  INV_X1 U14579 ( .A(n11926), .ZN(P1_U3231) );
  NAND2_X1 U14580 ( .A1(n11927), .A2(n11989), .ZN(n11928) );
  OR2_X1 U14581 ( .A1(n12619), .A2(n14641), .ZN(n11984) );
  NAND2_X1 U14582 ( .A1(n11928), .A2(n11984), .ZN(n11929) );
  XNOR2_X1 U14583 ( .A(n15188), .B(n14640), .ZN(n12762) );
  XNOR2_X1 U14584 ( .A(n11929), .B(n12762), .ZN(n15191) );
  INV_X1 U14585 ( .A(n14641), .ZN(n12618) );
  OR2_X1 U14586 ( .A1(n12619), .A2(n12618), .ZN(n11931) );
  NAND2_X1 U14587 ( .A1(n11930), .A2(n11931), .ZN(n11939) );
  INV_X1 U14588 ( .A(n12762), .ZN(n11932) );
  OR2_X1 U14589 ( .A1(n11932), .A2(n11931), .ZN(n11934) );
  AND2_X1 U14590 ( .A1(n11933), .A2(n11934), .ZN(n11968) );
  NAND2_X1 U14591 ( .A1(n11973), .A2(n11968), .ZN(n11937) );
  INV_X1 U14592 ( .A(n11934), .ZN(n11936) );
  AND2_X1 U14593 ( .A1(n12758), .A2(n12762), .ZN(n11935) );
  OR2_X1 U14594 ( .A1(n11936), .A2(n11935), .ZN(n11970) );
  NAND2_X1 U14595 ( .A1(n11937), .A2(n11970), .ZN(n11938) );
  OAI211_X1 U14596 ( .C1(n12762), .C2(n11939), .A(n11938), .B(n15389), .ZN(
        n11942) );
  NAND2_X1 U14597 ( .A1(n14639), .A2(n15031), .ZN(n11941) );
  NAND2_X1 U14598 ( .A1(n14641), .A2(n15029), .ZN(n11940) );
  AND2_X1 U14599 ( .A1(n11941), .A2(n11940), .ZN(n12031) );
  NAND2_X1 U14600 ( .A1(n11942), .A2(n12031), .ZN(n15186) );
  INV_X1 U14601 ( .A(n15186), .ZN(n11943) );
  MUX2_X1 U14602 ( .A(n11944), .B(n11943), .S(n15005), .Z(n11951) );
  NAND2_X1 U14603 ( .A1(n11945), .A2(n15188), .ZN(n11946) );
  NAND2_X1 U14604 ( .A1(n11946), .A2(n15377), .ZN(n11947) );
  NOR2_X1 U14605 ( .A1(n12106), .A2(n11947), .ZN(n15187) );
  INV_X1 U14606 ( .A(n15188), .ZN(n12637) );
  INV_X1 U14607 ( .A(n12033), .ZN(n11948) );
  OAI22_X1 U14608 ( .A1(n15394), .A2(n12637), .B1(n11948), .B2(n14985), .ZN(
        n11949) );
  AOI21_X1 U14609 ( .B1(n15187), .B2(n15400), .A(n11949), .ZN(n11950) );
  OAI211_X1 U14610 ( .C1(n15060), .C2(n15191), .A(n11951), .B(n11950), .ZN(
        P1_U3281) );
  OAI21_X1 U14611 ( .B1(n7751), .B2(n11953), .A(n11952), .ZN(n14408) );
  NAND3_X1 U14612 ( .A1(n11956), .A2(n7751), .A3(n11955), .ZN(n11957) );
  AOI21_X1 U14613 ( .B1(n11954), .B2(n11957), .A(n14217), .ZN(n11959) );
  NOR2_X1 U14614 ( .A1(n11959), .A2(n11958), .ZN(n14407) );
  MUX2_X1 U14615 ( .A(n11960), .B(n14407), .S(n14293), .Z(n11967) );
  INV_X1 U14616 ( .A(n11872), .ZN(n11962) );
  INV_X1 U14617 ( .A(n14287), .ZN(n11961) );
  AOI211_X1 U14618 ( .C1(n14405), .C2(n11962), .A(n8582), .B(n11961), .ZN(
        n14404) );
  OAI22_X1 U14619 ( .A1(n14275), .A2(n11964), .B1(n14290), .B2(n11963), .ZN(
        n11965) );
  AOI21_X1 U14620 ( .B1(n14404), .B2(n14282), .A(n11965), .ZN(n11966) );
  OAI211_X1 U14621 ( .C1(n14279), .C2(n14408), .A(n11967), .B(n11966), .ZN(
        P2_U3255) );
  OR2_X1 U14622 ( .A1(n15188), .A2(n12638), .ZN(n11969) );
  AND2_X1 U14623 ( .A1(n11968), .A2(n11969), .ZN(n11972) );
  INV_X1 U14624 ( .A(n11969), .ZN(n11971) );
  XNOR2_X1 U14625 ( .A(n15183), .B(n14639), .ZN(n12763) );
  NAND2_X1 U14626 ( .A1(n12110), .A2(n12763), .ZN(n12109) );
  OR2_X1 U14627 ( .A1(n15183), .A2(n11974), .ZN(n11975) );
  NAND2_X1 U14628 ( .A1(n12109), .A2(n11975), .ZN(n11977) );
  NAND2_X1 U14629 ( .A1(n15175), .A2(n11976), .ZN(n12655) );
  NAND2_X1 U14630 ( .A1(n11977), .A2(n12660), .ZN(n12908) );
  OAI211_X1 U14631 ( .C1(n11977), .C2(n12660), .A(n12908), .B(n15389), .ZN(
        n11979) );
  AOI22_X1 U14632 ( .A1(n15030), .A2(n15031), .B1(n15029), .B2(n14639), .ZN(
        n11978) );
  AND2_X1 U14633 ( .A1(n11979), .A2(n11978), .ZN(n15180) );
  INV_X1 U14634 ( .A(n15183), .ZN(n12647) );
  INV_X1 U14635 ( .A(n15175), .ZN(n11980) );
  OAI211_X1 U14636 ( .C1(n12107), .C2(n11980), .A(n15377), .B(n15051), .ZN(
        n15177) );
  AOI22_X1 U14637 ( .A1(n15405), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n14493), 
        .B2(n15392), .ZN(n11982) );
  NAND2_X1 U14638 ( .A1(n15175), .A2(n14954), .ZN(n11981) );
  OAI211_X1 U14639 ( .C1(n15177), .C2(n14935), .A(n11982), .B(n11981), .ZN(
        n11983) );
  INV_X1 U14640 ( .A(n11983), .ZN(n11998) );
  OR2_X1 U14641 ( .A1(n15188), .A2(n14640), .ZN(n11986) );
  AND2_X1 U14642 ( .A1(n11984), .A2(n11986), .ZN(n11988) );
  AND2_X1 U14643 ( .A1(n11985), .A2(n11988), .ZN(n11991) );
  INV_X1 U14644 ( .A(n11986), .ZN(n11987) );
  INV_X1 U14645 ( .A(n11988), .ZN(n11990) );
  INV_X1 U14646 ( .A(n12763), .ZN(n11993) );
  OR2_X1 U14647 ( .A1(n15183), .A2(n14639), .ZN(n11994) );
  NAND2_X1 U14648 ( .A1(n11995), .A2(n11994), .ZN(n11996) );
  NAND2_X1 U14649 ( .A1(n11996), .A2(n12660), .ZN(n15176) );
  NAND3_X1 U14650 ( .A1(n12939), .A2(n15176), .A3(n15381), .ZN(n11997) );
  OAI211_X1 U14651 ( .C1(n15180), .C2(n15405), .A(n11998), .B(n11997), .ZN(
        P1_U3279) );
  NOR2_X1 U14652 ( .A1(n11999), .A2(n12004), .ZN(n12000) );
  NOR2_X1 U14653 ( .A1(n12001), .A2(n12000), .ZN(n15624) );
  AOI22_X1 U14654 ( .A1(n14302), .A2(n13981), .B1(n13979), .B2(n14304), .ZN(
        n12008) );
  INV_X1 U14655 ( .A(n12002), .ZN(n12006) );
  AND3_X1 U14656 ( .A1(n10897), .A2(n12004), .A3(n12003), .ZN(n12005) );
  OAI21_X1 U14657 ( .B1(n12006), .B2(n12005), .A(n14307), .ZN(n12007) );
  OAI211_X1 U14658 ( .C1(n15624), .C2(n15642), .A(n12008), .B(n12007), .ZN(
        n15627) );
  INV_X1 U14659 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n12009) );
  OAI22_X1 U14660 ( .A1(n14293), .A2(n10496), .B1(n12009), .B2(n14290), .ZN(
        n12010) );
  AOI21_X1 U14661 ( .B1(n14295), .B2(n13741), .A(n12010), .ZN(n12014) );
  OAI211_X1 U14662 ( .C1(n12011), .C2(n15626), .A(n11261), .B(n14239), .ZN(
        n15625) );
  INV_X1 U14663 ( .A(n15625), .ZN(n12012) );
  NAND2_X1 U14664 ( .A1(n14282), .A2(n12012), .ZN(n12013) );
  OAI211_X1 U14665 ( .C1(n15624), .C2(n14265), .A(n12014), .B(n12013), .ZN(
        n12015) );
  AOI21_X1 U14666 ( .B1(n15627), .B2(n14293), .A(n12015), .ZN(n12016) );
  INV_X1 U14667 ( .A(n12016), .ZN(P2_U3263) );
  AND2_X1 U14668 ( .A1(n12018), .A2(n12017), .ZN(n12020) );
  NOR2_X1 U14669 ( .A1(n12020), .A2(n12021), .ZN(n12019) );
  AOI21_X1 U14670 ( .B1(n12021), .B2(n12020), .A(n12019), .ZN(n12026) );
  NAND2_X1 U14671 ( .A1(n14630), .A2(n12117), .ZN(n12022) );
  NAND2_X1 U14672 ( .A1(n6537), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n14765) );
  OAI211_X1 U14673 ( .C1(n12023), .C2(n14628), .A(n12022), .B(n14765), .ZN(
        n12024) );
  AOI21_X1 U14674 ( .B1(n14617), .B2(n12619), .A(n12024), .ZN(n12025) );
  OAI21_X1 U14675 ( .B1(n12026), .B2(n14619), .A(n12025), .ZN(P1_U3236) );
  OAI211_X1 U14676 ( .C1(n12029), .C2(n12028), .A(n12027), .B(n14621), .ZN(
        n12035) );
  OAI22_X1 U14677 ( .A1(n14628), .A2(n12031), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12030), .ZN(n12032) );
  AOI21_X1 U14678 ( .B1(n12033), .B2(n14630), .A(n12032), .ZN(n12034) );
  OAI211_X1 U14679 ( .C1(n12637), .C2(n14633), .A(n12035), .B(n12034), .ZN(
        P1_U3224) );
  INV_X1 U14680 ( .A(n15029), .ZN(n14941) );
  OAI21_X1 U14681 ( .B1(n12049), .B2(n12036), .A(n15389), .ZN(n12044) );
  INV_X1 U14682 ( .A(n12037), .ZN(n15398) );
  NAND2_X1 U14683 ( .A1(n12039), .A2(n12038), .ZN(n12040) );
  NAND2_X1 U14684 ( .A1(n15398), .A2(n12040), .ZN(n12047) );
  XNOR2_X1 U14685 ( .A(n12047), .B(n11669), .ZN(n12042) );
  AOI21_X1 U14686 ( .B1(n12042), .B2(n15389), .A(n12041), .ZN(n12043) );
  AOI21_X1 U14687 ( .B1(n14941), .B2(n12044), .A(n12043), .ZN(n12046) );
  NOR2_X1 U14688 ( .A1(n12046), .A2(n12045), .ZN(n15411) );
  OR2_X1 U14689 ( .A1(n12047), .A2(n15397), .ZN(n15409) );
  INV_X1 U14690 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n12048) );
  OAI22_X1 U14691 ( .A1(n14935), .A2(n15409), .B1(n12048), .B2(n14985), .ZN(
        n12052) );
  INV_X1 U14692 ( .A(n12049), .ZN(n12752) );
  XNOR2_X1 U14693 ( .A(n12752), .B(n12050), .ZN(n15408) );
  OAI22_X1 U14694 ( .A1(n15410), .A2(n15394), .B1(n15060), .B2(n15408), .ZN(
        n12051) );
  AOI211_X1 U14695 ( .C1(n15405), .C2(P1_REG2_REG_1__SCAN_IN), .A(n12052), .B(
        n12051), .ZN(n12053) );
  OAI21_X1 U14696 ( .B1(n15405), .B2(n15411), .A(n12053), .ZN(P1_U3292) );
  INV_X1 U14697 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15782) );
  INV_X1 U14698 ( .A(n12054), .ZN(n12057) );
  AOI211_X1 U14699 ( .C1(n15646), .C2(n12057), .A(n12056), .B(n12055), .ZN(
        n12059) );
  MUX2_X1 U14700 ( .A(n15782), .B(n12059), .S(n15659), .Z(n12058) );
  OAI21_X1 U14701 ( .B1(n12061), .B2(n14459), .A(n12058), .ZN(P2_U3457) );
  MUX2_X1 U14702 ( .A(n7372), .B(n12059), .S(n15670), .Z(n12060) );
  OAI21_X1 U14703 ( .B1(n12061), .B2(n14400), .A(n12060), .ZN(P2_U3508) );
  NAND2_X1 U14704 ( .A1(n15350), .A2(n12062), .ZN(n12063) );
  XNOR2_X1 U14705 ( .A(n12063), .B(n12754), .ZN(n15435) );
  XNOR2_X1 U14706 ( .A(n12064), .B(n12754), .ZN(n15438) );
  OR2_X1 U14707 ( .A1(n15405), .A2(n14809), .ZN(n14962) );
  OAI211_X1 U14708 ( .C1(n15376), .C2(n15434), .A(n15377), .B(n15361), .ZN(
        n15433) );
  INV_X1 U14709 ( .A(n15432), .ZN(n12066) );
  AOI22_X1 U14710 ( .A1(n15005), .A2(n12066), .B1(n12065), .B2(n15392), .ZN(
        n12067) );
  OAI21_X1 U14711 ( .B1(n10594), .B2(n15005), .A(n12067), .ZN(n12068) );
  AOI21_X1 U14712 ( .B1(n14954), .B2(n12586), .A(n12068), .ZN(n12069) );
  OAI21_X1 U14713 ( .B1(n14962), .B2(n15433), .A(n12069), .ZN(n12070) );
  AOI21_X1 U14714 ( .B1(n14983), .B2(n15438), .A(n12070), .ZN(n12071) );
  OAI21_X1 U14715 ( .B1(n15060), .B2(n15435), .A(n12071), .ZN(P1_U3288) );
  XNOR2_X1 U14716 ( .A(n12072), .B(n12749), .ZN(n15475) );
  INV_X1 U14717 ( .A(n15475), .ZN(n12083) );
  INV_X1 U14718 ( .A(n11973), .ZN(n12073) );
  AOI211_X1 U14719 ( .C1(n12749), .C2(n12074), .A(n15355), .B(n12073), .ZN(
        n15473) );
  INV_X1 U14720 ( .A(n15473), .ZN(n12075) );
  NAND2_X1 U14721 ( .A1(n14643), .A2(n15029), .ZN(n15469) );
  OAI211_X1 U14722 ( .C1(n14985), .C2(n12076), .A(n12075), .B(n15469), .ZN(
        n12081) );
  XNOR2_X1 U14723 ( .A(n12077), .B(n15472), .ZN(n12078) );
  AOI22_X1 U14724 ( .A1(n12078), .A2(n15377), .B1(n15031), .B2(n14641), .ZN(
        n15470) );
  NOR2_X1 U14725 ( .A1(n15470), .A2(n14935), .ZN(n12080) );
  OAI22_X1 U14726 ( .A1(n15472), .A2(n15394), .B1(n15005), .B2(n10606), .ZN(
        n12079) );
  AOI211_X1 U14727 ( .C1(n12081), .C2(n15005), .A(n12080), .B(n12079), .ZN(
        n12082) );
  OAI21_X1 U14728 ( .B1(n12083), .B2(n15060), .A(n12082), .ZN(P1_U3283) );
  NAND2_X1 U14729 ( .A1(n12085), .A2(n12084), .ZN(n13915) );
  XNOR2_X1 U14730 ( .A(n12086), .B(n13915), .ZN(n12087) );
  AOI222_X1 U14731 ( .A1(n14307), .A2(n12087), .B1(n14269), .B2(n14304), .C1(
        n13972), .C2(n14302), .ZN(n14395) );
  AOI211_X1 U14732 ( .C1(n14393), .C2(n14288), .A(n8582), .B(n12187), .ZN(
        n14392) );
  INV_X1 U14733 ( .A(n14393), .ZN(n12089) );
  AOI22_X1 U14734 ( .A1(n14308), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12135), 
        .B2(n14272), .ZN(n12088) );
  OAI21_X1 U14735 ( .B1(n12089), .B2(n14275), .A(n12088), .ZN(n12092) );
  XOR2_X1 U14736 ( .A(n12090), .B(n13915), .Z(n14396) );
  NOR2_X1 U14737 ( .A1(n14396), .A2(n14279), .ZN(n12091) );
  AOI211_X1 U14738 ( .C1(n14392), .C2(n14282), .A(n12092), .B(n12091), .ZN(
        n12093) );
  OAI21_X1 U14739 ( .B1(n14395), .B2(n14308), .A(n12093), .ZN(P2_U3253) );
  XNOR2_X1 U14740 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n12099) );
  XNOR2_X1 U14741 ( .A(n15255), .B(n12099), .ZN(n12102) );
  NAND2_X1 U14742 ( .A1(n12103), .A2(n12102), .ZN(n15252) );
  NAND2_X1 U14743 ( .A1(n15251), .A2(n15252), .ZN(n12104) );
  XNOR2_X1 U14744 ( .A(n12104), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  XNOR2_X1 U14745 ( .A(n12105), .B(n12763), .ZN(n15185) );
  INV_X1 U14746 ( .A(n12106), .ZN(n12108) );
  AOI211_X1 U14747 ( .C1(n15183), .C2(n12108), .A(n15397), .B(n12107), .ZN(
        n15182) );
  OAI211_X1 U14748 ( .C1(n12110), .C2(n12763), .A(n12109), .B(n15389), .ZN(
        n12112) );
  AOI22_X1 U14749 ( .A1(n15029), .A2(n14640), .B1(n14638), .B2(n15031), .ZN(
        n12111) );
  NAND2_X1 U14750 ( .A1(n12112), .A2(n12111), .ZN(n15181) );
  AOI21_X1 U14751 ( .B1(n15182), .B2(n12556), .A(n15181), .ZN(n12113) );
  MUX2_X1 U14752 ( .A(n12114), .B(n12113), .S(n15005), .Z(n12116) );
  AOI22_X1 U14753 ( .A1(n14954), .A2(n15183), .B1(n12175), .B2(n15392), .ZN(
        n12115) );
  OAI211_X1 U14754 ( .C1(n15185), .C2(n15060), .A(n12116), .B(n12115), .ZN(
        P1_U3280) );
  AOI22_X1 U14755 ( .A1(n14954), .A2(n12619), .B1(n15392), .B2(n12117), .ZN(
        n12118) );
  OAI21_X1 U14756 ( .B1(n12119), .B2(n14935), .A(n12118), .ZN(n12122) );
  MUX2_X1 U14757 ( .A(n12120), .B(P1_REG2_REG_11__SCAN_IN), .S(n15405), .Z(
        n12121) );
  AOI211_X1 U14758 ( .C1(n15381), .C2(n12123), .A(n12122), .B(n12121), .ZN(
        n12124) );
  INV_X1 U14759 ( .A(n12124), .ZN(P1_U3282) );
  XNOR2_X1 U14760 ( .A(n12126), .B(n12125), .ZN(n12130) );
  AOI22_X1 U14761 ( .A1(n14302), .A2(n14305), .B1(n14254), .B2(n14304), .ZN(
        n12185) );
  NAND2_X1 U14762 ( .A1(n13701), .A2(n12190), .ZN(n12127) );
  NAND2_X1 U14763 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n15564)
         );
  OAI211_X1 U14764 ( .C1(n12185), .C2(n13703), .A(n12127), .B(n15564), .ZN(
        n12128) );
  AOI21_X1 U14765 ( .B1(n14389), .B2(n13693), .A(n12128), .ZN(n12129) );
  OAI21_X1 U14766 ( .B1(n12130), .B2(n13695), .A(n12129), .ZN(P2_U3206) );
  INV_X1 U14767 ( .A(n12131), .ZN(n12132) );
  AOI21_X1 U14768 ( .B1(n12134), .B2(n12133), .A(n12132), .ZN(n12140) );
  AOI22_X1 U14769 ( .A1(n13722), .A2(n13972), .B1(n13701), .B2(n12135), .ZN(
        n12137) );
  OAI211_X1 U14770 ( .C1(n13574), .C2(n13718), .A(n12137), .B(n12136), .ZN(
        n12138) );
  AOI21_X1 U14771 ( .B1(n14393), .B2(n13693), .A(n12138), .ZN(n12139) );
  OAI21_X1 U14772 ( .B1(n12140), .B2(n13695), .A(n12139), .ZN(P2_U3196) );
  AOI21_X1 U14773 ( .B1(n12422), .B2(n12141), .A(n6712), .ZN(n12155) );
  XNOR2_X1 U14774 ( .A(n12142), .B(n10221), .ZN(n12143) );
  AOI222_X1 U14775 ( .A1(n13104), .A2(n13352), .B1(n13398), .B2(n12143), .C1(
        n13103), .C2(n13396), .ZN(n12150) );
  MUX2_X1 U14776 ( .A(n12144), .B(n12150), .S(n13405), .Z(n12146) );
  INV_X1 U14777 ( .A(n12267), .ZN(n12152) );
  AOI22_X1 U14778 ( .A1(n12152), .A2(n13438), .B1(n15675), .B2(n12270), .ZN(
        n12145) );
  OAI211_X1 U14779 ( .C1(n12155), .C2(n13441), .A(n12146), .B(n12145), .ZN(
        P3_U3219) );
  MUX2_X1 U14780 ( .A(n12147), .B(n12150), .S(n13486), .Z(n12149) );
  NAND2_X1 U14781 ( .A1(n12152), .A2(n13469), .ZN(n12148) );
  OAI211_X1 U14782 ( .C1(n12155), .C2(n13488), .A(n12149), .B(n12148), .ZN(
        P3_U3473) );
  MUX2_X1 U14783 ( .A(n12151), .B(n12150), .S(n15691), .Z(n12154) );
  NAND2_X1 U14784 ( .A1(n12152), .A2(n13520), .ZN(n12153) );
  OAI211_X1 U14785 ( .C1(n12155), .C2(n13540), .A(n12154), .B(n12153), .ZN(
        P3_U3432) );
  NAND2_X1 U14786 ( .A1(n12156), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n12160) );
  NAND2_X1 U14787 ( .A1(n12158), .A2(n12157), .ZN(n12159) );
  NAND2_X1 U14788 ( .A1(n12160), .A2(n12159), .ZN(n13984) );
  XNOR2_X1 U14789 ( .A(n13984), .B(n12166), .ZN(n13983) );
  XNOR2_X1 U14790 ( .A(n13983), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n12170) );
  INV_X1 U14791 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12162) );
  INV_X1 U14792 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14380) );
  XNOR2_X1 U14793 ( .A(n13997), .B(n14380), .ZN(n12168) );
  AND2_X1 U14794 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n13721) );
  AOI21_X1 U14795 ( .B1(n15527), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n13721), 
        .ZN(n12165) );
  OAI21_X1 U14796 ( .B1(n15584), .B2(n12166), .A(n12165), .ZN(n12167) );
  AOI21_X1 U14797 ( .B1(n12168), .B2(n15596), .A(n12167), .ZN(n12169) );
  OAI21_X1 U14798 ( .B1(n12170), .B2(n15579), .A(n12169), .ZN(P2_U3229) );
  OAI211_X1 U14799 ( .C1(n12173), .C2(n12172), .A(n12171), .B(n14621), .ZN(
        n12180) );
  INV_X1 U14800 ( .A(n12174), .ZN(n12178) );
  INV_X1 U14801 ( .A(n12175), .ZN(n12176) );
  OAI22_X1 U14802 ( .A1(n14609), .A2(n12638), .B1(n12176), .B2(n14611), .ZN(
        n12177) );
  AOI211_X1 U14803 ( .C1(n14591), .C2(n14638), .A(n12178), .B(n12177), .ZN(
        n12179) );
  OAI211_X1 U14804 ( .C1(n12647), .C2(n14633), .A(n12180), .B(n12179), .ZN(
        P1_U3234) );
  INV_X1 U14805 ( .A(n12181), .ZN(n12182) );
  OAI222_X1 U14806 ( .A1(n9621), .A2(P3_U3151), .B1(n12962), .B2(n12182), .C1(
        n7581), .C2(n13550), .ZN(P3_U3271) );
  XNOR2_X1 U14807 ( .A(n14389), .B(n13574), .ZN(n13919) );
  XNOR2_X1 U14808 ( .A(n12183), .B(n13919), .ZN(n14456) );
  XNOR2_X1 U14809 ( .A(n12184), .B(n13919), .ZN(n12186) );
  OAI21_X1 U14810 ( .B1(n12186), .B2(n14217), .A(n12185), .ZN(n14387) );
  NAND2_X1 U14811 ( .A1(n14387), .A2(n14293), .ZN(n12194) );
  INV_X1 U14812 ( .A(n12187), .ZN(n12189) );
  AOI211_X1 U14813 ( .C1(n14389), .C2(n12189), .A(n12188), .B(n8582), .ZN(
        n14388) );
  AOI22_X1 U14814 ( .A1(n14308), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12190), 
        .B2(n14272), .ZN(n12191) );
  OAI21_X1 U14815 ( .B1(n7626), .B2(n14275), .A(n12191), .ZN(n12192) );
  AOI21_X1 U14816 ( .B1(n14388), .B2(n14282), .A(n12192), .ZN(n12193) );
  OAI211_X1 U14817 ( .C1(n14456), .C2(n14279), .A(n12194), .B(n12193), .ZN(
        P2_U3252) );
  XNOR2_X1 U14818 ( .A(n12195), .B(n12501), .ZN(n12196) );
  AOI222_X1 U14819 ( .A1(n12207), .A2(n13352), .B1(n13398), .B2(n12196), .C1(
        n13049), .C2(n13396), .ZN(n12215) );
  MUX2_X1 U14820 ( .A(n15927), .B(n12215), .S(n13486), .Z(n12199) );
  XNOR2_X1 U14821 ( .A(n12197), .B(n12501), .ZN(n12214) );
  AOI22_X1 U14822 ( .A1(n12214), .A2(n13477), .B1(n13469), .B2(n12302), .ZN(
        n12198) );
  NAND2_X1 U14823 ( .A1(n12199), .A2(n12198), .ZN(P3_U3474) );
  INV_X1 U14824 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12200) );
  MUX2_X1 U14825 ( .A(n12200), .B(n12215), .S(n15691), .Z(n12202) );
  AOI22_X1 U14826 ( .A1(n12214), .A2(n13529), .B1(n13520), .B2(n12302), .ZN(
        n12201) );
  NAND2_X1 U14827 ( .A1(n12202), .A2(n12201), .ZN(P3_U3435) );
  OAI21_X1 U14828 ( .B1(n6719), .B2(n12204), .A(n12203), .ZN(n12205) );
  OAI211_X1 U14829 ( .C1(n12206), .C2(n6719), .A(n13058), .B(n12205), .ZN(
        n12213) );
  NAND2_X1 U14830 ( .A1(n13089), .A2(n12207), .ZN(n12208) );
  NAND2_X1 U14831 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13198)
         );
  OAI211_X1 U14832 ( .C1(n12209), .C2(n13093), .A(n12208), .B(n13198), .ZN(
        n12210) );
  AOI21_X1 U14833 ( .B1(n12211), .B2(n13090), .A(n12210), .ZN(n12212) );
  OAI211_X1 U14834 ( .C1(n12420), .C2(n13081), .A(n12213), .B(n12212), .ZN(
        P3_U3174) );
  INV_X1 U14835 ( .A(n12214), .ZN(n12218) );
  MUX2_X1 U14836 ( .A(n15758), .B(n12215), .S(n13405), .Z(n12217) );
  AOI22_X1 U14837 ( .A1(n12302), .A2(n13438), .B1(n12297), .B2(n15675), .ZN(
        n12216) );
  OAI211_X1 U14838 ( .C1(n12218), .C2(n13441), .A(n12217), .B(n12216), .ZN(
        P3_U3218) );
  INV_X1 U14839 ( .A(n12223), .ZN(n12504) );
  XNOR2_X1 U14840 ( .A(n12219), .B(n12504), .ZN(n12220) );
  AOI222_X1 U14841 ( .A1(n12220), .A2(n13398), .B1(n13102), .B2(n13396), .C1(
        n13103), .C2(n13352), .ZN(n12230) );
  MUX2_X1 U14842 ( .A(n12221), .B(n12230), .S(n13486), .Z(n12225) );
  NAND2_X1 U14843 ( .A1(n12222), .A2(n12223), .ZN(n12279) );
  OAI21_X1 U14844 ( .B1(n12222), .B2(n12223), .A(n12279), .ZN(n12229) );
  AOI22_X1 U14845 ( .A1(n12229), .A2(n13477), .B1(n13469), .B2(n13042), .ZN(
        n12224) );
  NAND2_X1 U14846 ( .A1(n12225), .A2(n12224), .ZN(P3_U3475) );
  INV_X1 U14847 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12226) );
  MUX2_X1 U14848 ( .A(n12226), .B(n12230), .S(n15691), .Z(n12228) );
  AOI22_X1 U14849 ( .A1(n12229), .A2(n13529), .B1(n13520), .B2(n13042), .ZN(
        n12227) );
  NAND2_X1 U14850 ( .A1(n12228), .A2(n12227), .ZN(P3_U3438) );
  INV_X1 U14851 ( .A(n12229), .ZN(n12234) );
  MUX2_X1 U14852 ( .A(n12231), .B(n12230), .S(n13405), .Z(n12233) );
  AOI22_X1 U14853 ( .A1(n13042), .A2(n13438), .B1(n15675), .B2(n13041), .ZN(
        n12232) );
  OAI211_X1 U14854 ( .C1(n12234), .C2(n13441), .A(n12233), .B(n12232), .ZN(
        P3_U3217) );
  INV_X1 U14855 ( .A(n12235), .ZN(n12236) );
  NOR2_X1 U14856 ( .A1(n12237), .A2(n12236), .ZN(n12250) );
  INV_X1 U14857 ( .A(n12250), .ZN(n12238) );
  NAND2_X1 U14858 ( .A1(n12237), .A2(n12236), .ZN(n12251) );
  NAND2_X1 U14859 ( .A1(n12238), .A2(n12251), .ZN(n12239) );
  XNOR2_X1 U14860 ( .A(n12239), .B(n12255), .ZN(n12247) );
  NOR2_X1 U14861 ( .A1(n12240), .A2(n13081), .ZN(n12244) );
  NAND2_X1 U14862 ( .A1(n13089), .A2(n13105), .ZN(n12241) );
  NAND2_X1 U14863 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n13165)
         );
  OAI211_X1 U14864 ( .C1(n12242), .C2(n13093), .A(n12241), .B(n13165), .ZN(
        n12243) );
  AOI211_X1 U14865 ( .C1(n12245), .C2(n13090), .A(n12244), .B(n12243), .ZN(
        n12246) );
  OAI21_X1 U14866 ( .B1(n12247), .B2(n13098), .A(n12246), .ZN(P3_U3176) );
  NAND2_X1 U14867 ( .A1(n12249), .A2(n12248), .ZN(n12253) );
  AOI21_X1 U14868 ( .B1(n12255), .B2(n12251), .A(n12250), .ZN(n12252) );
  XOR2_X1 U14869 ( .A(n12253), .B(n12252), .Z(n12261) );
  NAND2_X1 U14870 ( .A1(n13089), .A2(n13104), .ZN(n12254) );
  NAND2_X1 U14871 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13179)
         );
  OAI211_X1 U14872 ( .C1(n12255), .C2(n13093), .A(n12254), .B(n13179), .ZN(
        n12258) );
  NOR2_X1 U14873 ( .A1(n12256), .A2(n13081), .ZN(n12257) );
  AOI211_X1 U14874 ( .C1(n12259), .C2(n13090), .A(n12258), .B(n12257), .ZN(
        n12260) );
  OAI21_X1 U14875 ( .B1(n12261), .B2(n13098), .A(n12260), .ZN(P3_U3164) );
  XOR2_X1 U14876 ( .A(n12263), .B(n12262), .Z(n12272) );
  NAND2_X1 U14877 ( .A1(n13089), .A2(n13103), .ZN(n12265) );
  OAI211_X1 U14878 ( .C1(n12266), .C2(n13093), .A(n12265), .B(n12264), .ZN(
        n12269) );
  NOR2_X1 U14879 ( .A1(n12267), .A2(n13081), .ZN(n12268) );
  AOI211_X1 U14880 ( .C1(n12270), .C2(n13090), .A(n12269), .B(n12268), .ZN(
        n12271) );
  OAI21_X1 U14881 ( .B1(n12272), .B2(n13098), .A(n12271), .ZN(P3_U3155) );
  INV_X1 U14882 ( .A(n12273), .ZN(n12274) );
  AOI21_X1 U14883 ( .B1(n12274), .B2(n7220), .A(n13428), .ZN(n12278) );
  OAI22_X1 U14884 ( .A1(n13413), .A2(n13433), .B1(n12275), .B2(n13431), .ZN(
        n12276) );
  AOI21_X1 U14885 ( .B1(n12278), .B2(n12277), .A(n12276), .ZN(n12290) );
  MUX2_X1 U14886 ( .A(n13253), .B(n12290), .S(n13405), .Z(n12284) );
  NAND2_X1 U14887 ( .A1(n12279), .A2(n12439), .ZN(n12280) );
  XNOR2_X1 U14888 ( .A(n12280), .B(n7220), .ZN(n12289) );
  INV_X1 U14889 ( .A(n13054), .ZN(n12281) );
  OAI22_X1 U14890 ( .A1(n13051), .A2(n13403), .B1(n12281), .B2(n15681), .ZN(
        n12282) );
  AOI21_X1 U14891 ( .B1(n12289), .B2(n11212), .A(n12282), .ZN(n12283) );
  NAND2_X1 U14892 ( .A1(n12284), .A2(n12283), .ZN(P3_U3216) );
  AOI22_X1 U14893 ( .A1(n12289), .A2(n13477), .B1(n13469), .B2(n12288), .ZN(
        n12287) );
  MUX2_X1 U14894 ( .A(n12285), .B(n12290), .S(n13486), .Z(n12286) );
  NAND2_X1 U14895 ( .A1(n12287), .A2(n12286), .ZN(P3_U3476) );
  AOI22_X1 U14896 ( .A1(n12289), .A2(n13529), .B1(n13520), .B2(n12288), .ZN(
        n12293) );
  INV_X1 U14897 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12291) );
  MUX2_X1 U14898 ( .A(n12291), .B(n12290), .S(n15691), .Z(n12292) );
  NAND2_X1 U14899 ( .A1(n12293), .A2(n12292), .ZN(P3_U3441) );
  XNOR2_X1 U14900 ( .A(n12295), .B(n13103), .ZN(n12296) );
  XNOR2_X1 U14901 ( .A(n12294), .B(n12296), .ZN(n12304) );
  NAND2_X1 U14902 ( .A1(n13090), .A2(n12297), .ZN(n12299) );
  AND2_X1 U14903 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13218) );
  AOI21_X1 U14904 ( .B1(n13089), .B2(n13049), .A(n13218), .ZN(n12298) );
  OAI211_X1 U14905 ( .C1(n12300), .C2(n13093), .A(n12299), .B(n12298), .ZN(
        n12301) );
  AOI21_X1 U14906 ( .B1(n12302), .B2(n13096), .A(n12301), .ZN(n12303) );
  OAI21_X1 U14907 ( .B1(n12304), .B2(n13098), .A(n12303), .ZN(P3_U3181) );
  MUX2_X1 U14908 ( .A(n12305), .B(P2_REG2_REG_1__SCAN_IN), .S(n14308), .Z(
        n12315) );
  INV_X1 U14909 ( .A(n14265), .ZN(n12307) );
  NAND2_X1 U14910 ( .A1(n12307), .A2(n12306), .ZN(n12313) );
  NAND2_X1 U14911 ( .A1(n14282), .A2(n12308), .ZN(n12312) );
  INV_X1 U14912 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n12309) );
  OR2_X1 U14913 ( .A1(n14290), .A2(n12309), .ZN(n12311) );
  OR2_X1 U14914 ( .A1(n14275), .A2(n13742), .ZN(n12310) );
  NAND4_X1 U14915 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12314) );
  OR2_X1 U14916 ( .A1(n12315), .A2(n12314), .ZN(P2_U3264) );
  INV_X1 U14917 ( .A(n12316), .ZN(n15231) );
  OAI222_X1 U14918 ( .A1(P2_U3088), .A2(n13953), .B1(n10996), .B2(n15231), 
        .C1(n12317), .C2(n14478), .ZN(P2_U3300) );
  INV_X1 U14919 ( .A(n12318), .ZN(n14475) );
  OAI222_X1 U14920 ( .A1(n15232), .A2(n12319), .B1(n15236), .B2(n14475), .C1(
        P1_U3086), .C2(n9335), .ZN(P1_U3327) );
  INV_X1 U14921 ( .A(n12320), .ZN(n12321) );
  XNOR2_X1 U14922 ( .A(n12806), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n12795) );
  XNOR2_X1 U14923 ( .A(n12796), .B(n12795), .ZN(n13542) );
  NAND2_X1 U14924 ( .A1(n13542), .A2(n9742), .ZN(n12324) );
  NAND2_X1 U14925 ( .A1(n9995), .A2(SI_30_), .ZN(n12323) );
  INV_X1 U14926 ( .A(n13100), .ZN(n12476) );
  NAND2_X1 U14927 ( .A1(n12519), .A2(n12476), .ZN(n12345) );
  XNOR2_X1 U14928 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12326) );
  INV_X1 U14929 ( .A(n12326), .ZN(n12797) );
  INV_X1 U14930 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15223) );
  NAND2_X1 U14931 ( .A1(n15223), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U14932 ( .A1(n12797), .A2(n12325), .ZN(n12334) );
  NAND2_X1 U14933 ( .A1(n12806), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12794) );
  OAI21_X1 U14934 ( .B1(n12326), .B2(n15223), .A(n12806), .ZN(n12329) );
  NAND2_X1 U14935 ( .A1(n12326), .A2(n15223), .ZN(n12327) );
  NAND2_X1 U14936 ( .A1(n12327), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12328) );
  AND2_X1 U14937 ( .A1(n12329), .A2(n12328), .ZN(n12330) );
  NOR2_X1 U14938 ( .A1(n12331), .A2(n12330), .ZN(n12332) );
  OAI211_X1 U14939 ( .C1(n12796), .C2(n12334), .A(n12333), .B(n12332), .ZN(
        n12336) );
  NAND2_X1 U14940 ( .A1(n9995), .A2(SI_31_), .ZN(n12335) );
  NAND2_X1 U14941 ( .A1(n12336), .A2(n12335), .ZN(n12478) );
  NAND2_X1 U14942 ( .A1(n9746), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12341) );
  NAND2_X1 U14943 ( .A1(n12337), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U14944 ( .A1(n6539), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12339) );
  AND3_X1 U14945 ( .A1(n12341), .A2(n12340), .A3(n12339), .ZN(n12342) );
  MUX2_X1 U14946 ( .A(n12461), .B(n12460), .S(n9474), .Z(n12466) );
  MUX2_X1 U14947 ( .A(n12347), .B(n12348), .S(n9474), .Z(n12452) );
  MUX2_X1 U14948 ( .A(n12350), .B(n12349), .S(n9474), .Z(n12450) );
  INV_X1 U14949 ( .A(n13393), .ZN(n12448) );
  MUX2_X1 U14950 ( .A(n12357), .B(n12353), .S(n9474), .Z(n12444) );
  INV_X1 U14951 ( .A(n12351), .ZN(n12352) );
  NAND2_X1 U14952 ( .A1(n13427), .A2(n12352), .ZN(n12354) );
  NAND3_X1 U14953 ( .A1(n12354), .A2(n12353), .A3(n12355), .ZN(n12361) );
  INV_X1 U14954 ( .A(n12355), .ZN(n12359) );
  OAI211_X1 U14955 ( .C1(n12359), .C2(n12358), .A(n12357), .B(n12356), .ZN(
        n12360) );
  MUX2_X1 U14956 ( .A(n12361), .B(n12360), .S(n9474), .Z(n12362) );
  INV_X1 U14957 ( .A(n12364), .ZN(n12366) );
  OAI22_X1 U14958 ( .A1(n12367), .A2(n12366), .B1(n12365), .B2(n9625), .ZN(
        n12369) );
  AOI21_X1 U14959 ( .B1(n12369), .B2(n12368), .A(n12483), .ZN(n12370) );
  AND2_X1 U14960 ( .A1(n12376), .A2(n12371), .ZN(n12374) );
  AND2_X1 U14961 ( .A1(n12377), .A2(n12372), .ZN(n12373) );
  MUX2_X1 U14962 ( .A(n12374), .B(n12373), .S(n9474), .Z(n12375) );
  MUX2_X1 U14963 ( .A(n12377), .B(n12376), .S(n9474), .Z(n12378) );
  NAND3_X1 U14964 ( .A1(n12379), .A2(n12486), .A3(n12378), .ZN(n12383) );
  MUX2_X1 U14965 ( .A(n12381), .B(n12380), .S(n9474), .Z(n12382) );
  NAND3_X1 U14966 ( .A1(n12383), .A2(n12489), .A3(n12382), .ZN(n12387) );
  NAND2_X1 U14967 ( .A1(n12392), .A2(n12384), .ZN(n12385) );
  NAND2_X1 U14968 ( .A1(n9474), .A2(n12385), .ZN(n12386) );
  NAND2_X1 U14969 ( .A1(n12387), .A2(n12386), .ZN(n12391) );
  NAND2_X1 U14970 ( .A1(n12390), .A2(n12388), .ZN(n12389) );
  AOI22_X1 U14971 ( .A1(n12391), .A2(n12390), .B1(n12462), .B2(n12389), .ZN(
        n12397) );
  OAI21_X1 U14972 ( .B1(n9474), .B2(n12392), .A(n12491), .ZN(n12396) );
  MUX2_X1 U14973 ( .A(n12394), .B(n12393), .S(n9474), .Z(n12395) );
  OAI211_X1 U14974 ( .C1(n12397), .C2(n12396), .A(n7206), .B(n12395), .ZN(
        n12402) );
  INV_X1 U14975 ( .A(n12497), .ZN(n12401) );
  MUX2_X1 U14976 ( .A(n12399), .B(n12398), .S(n9474), .Z(n12400) );
  INV_X1 U14977 ( .A(n12494), .ZN(n12407) );
  MUX2_X1 U14978 ( .A(n12404), .B(n12403), .S(n12462), .Z(n12405) );
  OAI211_X1 U14979 ( .C1(n12498), .C2(n12409), .A(n12417), .B(n12408), .ZN(
        n12413) );
  OAI211_X1 U14980 ( .C1(n12498), .C2(n12411), .A(n12416), .B(n12410), .ZN(
        n12412) );
  MUX2_X1 U14981 ( .A(n12413), .B(n12412), .S(n12462), .Z(n12414) );
  INV_X1 U14982 ( .A(n12414), .ZN(n12415) );
  MUX2_X1 U14983 ( .A(n12417), .B(n12416), .S(n9474), .Z(n12418) );
  OR2_X1 U14984 ( .A1(n9474), .A2(n13104), .ZN(n12419) );
  NOR2_X1 U14985 ( .A1(n12420), .A2(n12419), .ZN(n12421) );
  NOR2_X1 U14986 ( .A1(n12422), .A2(n12421), .ZN(n12423) );
  NAND2_X1 U14987 ( .A1(n12424), .A2(n12423), .ZN(n12433) );
  AOI21_X1 U14988 ( .B1(n12433), .B2(n12425), .A(n7736), .ZN(n12429) );
  NAND2_X1 U14989 ( .A1(n12427), .A2(n12426), .ZN(n12428) );
  OAI21_X1 U14990 ( .B1(n12429), .B2(n12428), .A(n12462), .ZN(n12437) );
  INV_X1 U14991 ( .A(n12430), .ZN(n12432) );
  OAI22_X1 U14992 ( .A1(n12433), .A2(n12432), .B1(n12431), .B2(n12462), .ZN(
        n12434) );
  NAND2_X1 U14993 ( .A1(n12434), .A2(n12501), .ZN(n12436) );
  INV_X1 U14994 ( .A(n12439), .ZN(n12435) );
  AOI21_X1 U14995 ( .B1(n12437), .B2(n12436), .A(n12435), .ZN(n12442) );
  AOI21_X1 U14996 ( .B1(n12439), .B2(n12438), .A(n12462), .ZN(n12441) );
  NAND2_X1 U14997 ( .A1(n13049), .A2(n9474), .ZN(n12440) );
  OAI22_X1 U14998 ( .A1(n12442), .A2(n12441), .B1(n13042), .B2(n12440), .ZN(
        n12443) );
  NAND2_X1 U14999 ( .A1(n13057), .A2(n13414), .ZN(n12446) );
  MUX2_X1 U15000 ( .A(n12446), .B(n12445), .S(n9474), .Z(n12447) );
  NAND3_X1 U15001 ( .A1(n13381), .A2(n12450), .A3(n12449), .ZN(n12451) );
  NAND2_X1 U15002 ( .A1(n12454), .A2(n12453), .ZN(n12455) );
  AND2_X1 U15003 ( .A1(n12455), .A2(n12456), .ZN(n12459) );
  OAI21_X1 U15004 ( .B1(n13351), .B2(n12457), .A(n12456), .ZN(n12458) );
  MUX2_X1 U15005 ( .A(n12459), .B(n12458), .S(n9474), .Z(n12465) );
  MUX2_X1 U15006 ( .A(n12462), .B(n13353), .S(n12874), .Z(n12463) );
  OAI21_X1 U15007 ( .B1(n13094), .B2(n9474), .A(n12463), .ZN(n12464) );
  OR3_X1 U15008 ( .A1(n12991), .A2(n12888), .A3(n9474), .ZN(n12468) );
  NAND3_X1 U15009 ( .A1(n12470), .A2(n9474), .A3(n12469), .ZN(n12472) );
  OAI211_X1 U15010 ( .C1(n12474), .C2(n9474), .A(n12473), .B(n12516), .ZN(
        n12481) );
  NAND2_X1 U15011 ( .A1(n12478), .A2(n12477), .ZN(n12475) );
  OAI21_X1 U15012 ( .B1(n12519), .B2(n12476), .A(n12475), .ZN(n12479) );
  INV_X1 U15013 ( .A(n12479), .ZN(n12511) );
  NAND2_X1 U15014 ( .A1(n12479), .A2(n12478), .ZN(n12524) );
  OAI21_X1 U15015 ( .B1(n12511), .B2(n13290), .A(n12524), .ZN(n12480) );
  INV_X1 U15016 ( .A(n15679), .ZN(n12482) );
  INV_X1 U15017 ( .A(n13322), .ZN(n13321) );
  INV_X1 U15018 ( .A(n13381), .ZN(n13382) );
  NOR2_X1 U15019 ( .A1(n12484), .A2(n12483), .ZN(n12488) );
  AND4_X1 U15020 ( .A1(n12488), .A2(n12487), .A3(n12486), .A4(n12485), .ZN(
        n12492) );
  NAND4_X1 U15021 ( .A1(n12492), .A2(n12491), .A3(n12490), .A4(n12489), .ZN(
        n12495) );
  OR3_X1 U15022 ( .A1(n12495), .A2(n12494), .A3(n12493), .ZN(n12496) );
  NOR4_X1 U15023 ( .A1(n12499), .A2(n12498), .A3(n12497), .A4(n12496), .ZN(
        n12500) );
  NAND4_X1 U15024 ( .A1(n10221), .A2(n12502), .A3(n12501), .A4(n12500), .ZN(
        n12503) );
  NOR4_X1 U15025 ( .A1(n7740), .A2(n12505), .A3(n12504), .A4(n12503), .ZN(
        n12506) );
  NAND2_X1 U15026 ( .A1(n12506), .A2(n13411), .ZN(n12507) );
  NOR4_X1 U15027 ( .A1(n13382), .A2(n13393), .A3(n12541), .A4(n12507), .ZN(
        n12508) );
  NOR2_X1 U15028 ( .A1(n12512), .A2(n10060), .ZN(n12513) );
  INV_X1 U15029 ( .A(n12516), .ZN(n12517) );
  INV_X1 U15030 ( .A(n12524), .ZN(n12527) );
  AOI21_X1 U15031 ( .B1(n12527), .B2(n12526), .A(n12525), .ZN(n12529) );
  NAND2_X1 U15032 ( .A1(n12531), .A2(n12530), .ZN(n12532) );
  OAI211_X1 U15033 ( .C1(n12533), .C2(n13548), .A(P3_B_REG_SCAN_IN), .B(n12532), .ZN(n12534) );
  INV_X1 U15034 ( .A(n12536), .ZN(n15512) );
  OAI222_X1 U15035 ( .A1(n15512), .A2(P2_U3088), .B1(n10996), .B2(n12537), 
        .C1(n9633), .C2(n14478), .ZN(P2_U3325) );
  XNOR2_X1 U15036 ( .A(n12538), .B(n12541), .ZN(n12554) );
  OAI211_X1 U15037 ( .C1(n12541), .C2(n12540), .A(n12539), .B(n13398), .ZN(
        n12543) );
  AOI22_X1 U15038 ( .A1(n13384), .A2(n13396), .B1(n13352), .B2(n13101), .ZN(
        n12542) );
  AND2_X1 U15039 ( .A1(n12543), .A2(n12542), .ZN(n12551) );
  INV_X1 U15040 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12544) );
  MUX2_X1 U15041 ( .A(n12551), .B(n12544), .S(n15693), .Z(n12546) );
  NAND2_X1 U15042 ( .A1(n13057), .A2(n13520), .ZN(n12545) );
  OAI211_X1 U15043 ( .C1(n12554), .C2(n13540), .A(n12546), .B(n12545), .ZN(
        P3_U3447) );
  INV_X1 U15044 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12547) );
  MUX2_X1 U15045 ( .A(n12547), .B(n12551), .S(n13486), .Z(n12549) );
  NAND2_X1 U15046 ( .A1(n13057), .A2(n13469), .ZN(n12548) );
  OAI211_X1 U15047 ( .C1(n12554), .C2(n13488), .A(n12549), .B(n12548), .ZN(
        P3_U3479) );
  MUX2_X1 U15048 ( .A(n12551), .B(n12550), .S(n15688), .Z(n12553) );
  AOI22_X1 U15049 ( .A1(n13057), .A2(n13438), .B1(n15675), .B2(n13064), .ZN(
        n12552) );
  OAI211_X1 U15050 ( .C1(n12554), .C2(n13441), .A(n12553), .B(n12552), .ZN(
        P3_U3213) );
  NAND2_X1 U15051 ( .A1(n12560), .A2(n12559), .ZN(n12561) );
  XNOR2_X1 U15052 ( .A(n12562), .B(n12571), .ZN(n12564) );
  NAND2_X1 U15053 ( .A1(n12750), .A2(n12719), .ZN(n12563) );
  NAND3_X1 U15054 ( .A1(n12752), .A2(n12564), .A3(n12563), .ZN(n12568) );
  INV_X4 U15055 ( .A(n12571), .ZN(n12730) );
  MUX2_X1 U15056 ( .A(n12566), .B(n12565), .S(n12730), .Z(n12567) );
  NAND2_X1 U15057 ( .A1(n12568), .A2(n12567), .ZN(n12574) );
  NAND2_X1 U15058 ( .A1(n12571), .A2(n15399), .ZN(n12569) );
  NAND2_X1 U15059 ( .A1(n12570), .A2(n12569), .ZN(n12573) );
  OAI21_X1 U15060 ( .B1(n12574), .B2(n12573), .A(n12572), .ZN(n12576) );
  NAND3_X1 U15061 ( .A1(n12574), .A2(n15399), .A3(n12573), .ZN(n12575) );
  NAND3_X1 U15062 ( .A1(n12576), .A2(n12575), .A3(n12753), .ZN(n12580) );
  NAND2_X1 U15063 ( .A1(n11674), .A2(n14649), .ZN(n12578) );
  MUX2_X1 U15064 ( .A(n12578), .B(n12577), .S(n12730), .Z(n12579) );
  MUX2_X1 U15065 ( .A(n12581), .B(n15427), .S(n12571), .Z(n12583) );
  MUX2_X1 U15066 ( .A(n14648), .B(n14572), .S(n12730), .Z(n12582) );
  NAND2_X1 U15067 ( .A1(n12584), .A2(n12583), .ZN(n12585) );
  MUX2_X1 U15068 ( .A(n12586), .B(n14647), .S(n12571), .Z(n12588) );
  MUX2_X1 U15069 ( .A(n12586), .B(n14647), .S(n12730), .Z(n12587) );
  INV_X1 U15070 ( .A(n12588), .ZN(n12589) );
  MUX2_X1 U15071 ( .A(n12590), .B(n14646), .S(n12730), .Z(n12594) );
  MUX2_X1 U15072 ( .A(n15440), .B(n12591), .S(n12571), .Z(n12592) );
  INV_X1 U15073 ( .A(n12593), .ZN(n12611) );
  MUX2_X1 U15074 ( .A(n12597), .B(n12596), .S(n12730), .Z(n12635) );
  MUX2_X1 U15075 ( .A(n14645), .B(n12598), .S(n12571), .Z(n12634) );
  MUX2_X1 U15076 ( .A(n12599), .B(n15472), .S(n12571), .Z(n12621) );
  MUX2_X1 U15077 ( .A(n14642), .B(n12600), .S(n12730), .Z(n12620) );
  NAND2_X1 U15078 ( .A1(n12621), .A2(n12620), .ZN(n12628) );
  MUX2_X1 U15079 ( .A(n12602), .B(n12601), .S(n12571), .Z(n12625) );
  MUX2_X1 U15080 ( .A(n14643), .B(n12603), .S(n12730), .Z(n12624) );
  NAND2_X1 U15081 ( .A1(n12625), .A2(n12624), .ZN(n12604) );
  AND2_X1 U15082 ( .A1(n12628), .A2(n12604), .ZN(n12612) );
  MUX2_X1 U15083 ( .A(n12606), .B(n12605), .S(n12571), .Z(n12614) );
  MUX2_X1 U15084 ( .A(n14644), .B(n12607), .S(n12730), .Z(n12613) );
  NAND2_X1 U15085 ( .A1(n12614), .A2(n12613), .ZN(n12608) );
  AND2_X1 U15086 ( .A1(n12612), .A2(n12608), .ZN(n12636) );
  OAI21_X1 U15087 ( .B1(n12635), .B2(n12634), .A(n12636), .ZN(n12609) );
  INV_X1 U15088 ( .A(n12609), .ZN(n12610) );
  NAND3_X1 U15089 ( .A1(n12611), .A2(n6649), .A3(n12610), .ZN(n12640) );
  INV_X1 U15090 ( .A(n12612), .ZN(n12632) );
  INV_X1 U15091 ( .A(n12613), .ZN(n12616) );
  INV_X1 U15092 ( .A(n12614), .ZN(n12615) );
  NAND2_X1 U15093 ( .A1(n12616), .A2(n12615), .ZN(n12631) );
  MUX2_X1 U15094 ( .A(n12618), .B(n12617), .S(n12730), .Z(n12642) );
  MUX2_X1 U15095 ( .A(n14641), .B(n12619), .S(n12571), .Z(n12641) );
  INV_X1 U15096 ( .A(n12620), .ZN(n12623) );
  INV_X1 U15097 ( .A(n12621), .ZN(n12622) );
  AOI22_X1 U15098 ( .A1(n12642), .A2(n12641), .B1(n12623), .B2(n12622), .ZN(
        n12630) );
  INV_X1 U15099 ( .A(n12624), .ZN(n12627) );
  INV_X1 U15100 ( .A(n12625), .ZN(n12626) );
  NAND3_X1 U15101 ( .A1(n12628), .A2(n12627), .A3(n12626), .ZN(n12629) );
  OAI211_X1 U15102 ( .C1(n12632), .C2(n12631), .A(n12630), .B(n12629), .ZN(
        n12633) );
  NAND3_X1 U15103 ( .A1(n12636), .A2(n12635), .A3(n12634), .ZN(n12639) );
  MUX2_X1 U15104 ( .A(n12638), .B(n12637), .S(n12730), .Z(n12651) );
  MUX2_X1 U15105 ( .A(n14640), .B(n15188), .S(n12571), .Z(n12650) );
  NAND2_X1 U15106 ( .A1(n12651), .A2(n12650), .ZN(n12645) );
  INV_X1 U15107 ( .A(n12641), .ZN(n12644) );
  INV_X1 U15108 ( .A(n12642), .ZN(n12643) );
  NAND3_X1 U15109 ( .A1(n12645), .A2(n12644), .A3(n12643), .ZN(n12649) );
  MUX2_X1 U15110 ( .A(n14639), .B(n15183), .S(n12730), .Z(n12657) );
  NAND2_X1 U15111 ( .A1(n14639), .A2(n12730), .ZN(n12646) );
  OAI211_X1 U15112 ( .C1(n12647), .C2(n12730), .A(n12657), .B(n12646), .ZN(
        n12648) );
  OAI211_X1 U15113 ( .C1(n12651), .C2(n12650), .A(n12649), .B(n12648), .ZN(
        n12652) );
  INV_X1 U15114 ( .A(n12652), .ZN(n12653) );
  NAND2_X1 U15115 ( .A1(n12909), .A2(n12907), .ZN(n12654) );
  NAND2_X1 U15116 ( .A1(n12654), .A2(n12730), .ZN(n12663) );
  NAND2_X1 U15117 ( .A1(n15171), .A2(n14541), .ZN(n12746) );
  NAND2_X1 U15118 ( .A1(n12746), .A2(n12655), .ZN(n12656) );
  NAND2_X1 U15119 ( .A1(n12656), .A2(n12571), .ZN(n12662) );
  INV_X1 U15120 ( .A(n12657), .ZN(n12659) );
  MUX2_X1 U15121 ( .A(n14639), .B(n15183), .S(n12571), .Z(n12658) );
  NAND3_X1 U15122 ( .A1(n12660), .A2(n12659), .A3(n12658), .ZN(n12661) );
  MUX2_X1 U15123 ( .A(n12746), .B(n12909), .S(n12571), .Z(n12664) );
  MUX2_X1 U15124 ( .A(n15016), .B(n15166), .S(n12730), .Z(n12667) );
  MUX2_X1 U15125 ( .A(n15016), .B(n15166), .S(n12571), .Z(n12665) );
  NAND2_X1 U15126 ( .A1(n15156), .A2(n15015), .ZN(n12943) );
  MUX2_X1 U15127 ( .A(n15032), .B(n15161), .S(n12571), .Z(n12671) );
  NAND2_X1 U15128 ( .A1(n15161), .A2(n15032), .ZN(n12941) );
  NAND2_X1 U15129 ( .A1(n12671), .A2(n12941), .ZN(n12668) );
  INV_X1 U15130 ( .A(n14993), .ZN(n14602) );
  OAI21_X1 U15131 ( .B1(n15015), .B2(n12730), .A(n12943), .ZN(n12669) );
  NAND2_X1 U15132 ( .A1(n12767), .A2(n12669), .ZN(n12670) );
  OAI21_X1 U15133 ( .B1(n12571), .B2(n15156), .A(n12670), .ZN(n12674) );
  NOR2_X1 U15134 ( .A1(n15161), .A2(n15032), .ZN(n12942) );
  NOR2_X1 U15135 ( .A1(n12671), .A2(n12942), .ZN(n12672) );
  NAND2_X1 U15136 ( .A1(n14995), .A2(n12672), .ZN(n12673) );
  NAND2_X1 U15137 ( .A1(n15150), .A2(n14602), .ZN(n12914) );
  MUX2_X1 U15138 ( .A(n12914), .B(n12767), .S(n12730), .Z(n12675) );
  INV_X1 U15139 ( .A(n15143), .ZN(n14971) );
  MUX2_X1 U15140 ( .A(n14637), .B(n15143), .S(n12571), .Z(n12676) );
  MUX2_X1 U15141 ( .A(n14964), .B(n14955), .S(n12571), .Z(n12680) );
  NAND2_X1 U15142 ( .A1(n12681), .A2(n12680), .ZN(n12679) );
  MUX2_X1 U15143 ( .A(n14964), .B(n14955), .S(n12730), .Z(n12678) );
  NAND2_X1 U15144 ( .A1(n12679), .A2(n12678), .ZN(n12683) );
  MUX2_X1 U15145 ( .A(n14636), .B(n7662), .S(n12730), .Z(n12685) );
  MUX2_X1 U15146 ( .A(n14944), .B(n15129), .S(n12571), .Z(n12684) );
  MUX2_X1 U15147 ( .A(n14930), .B(n15121), .S(n12571), .Z(n12687) );
  MUX2_X1 U15148 ( .A(n14930), .B(n15121), .S(n12730), .Z(n12686) );
  MUX2_X1 U15149 ( .A(n14907), .B(n15111), .S(n12730), .Z(n12692) );
  MUX2_X1 U15150 ( .A(n14907), .B(n15111), .S(n12571), .Z(n12689) );
  NAND2_X1 U15151 ( .A1(n12690), .A2(n12689), .ZN(n12696) );
  INV_X1 U15152 ( .A(n12691), .ZN(n12694) );
  INV_X1 U15153 ( .A(n12692), .ZN(n12693) );
  MUX2_X1 U15154 ( .A(n14887), .B(n14879), .S(n12571), .Z(n12698) );
  MUX2_X1 U15155 ( .A(n14887), .B(n14879), .S(n12730), .Z(n12697) );
  MUX2_X1 U15156 ( .A(n14870), .B(n14860), .S(n12730), .Z(n12700) );
  MUX2_X1 U15157 ( .A(n14870), .B(n14860), .S(n12571), .Z(n12699) );
  INV_X1 U15158 ( .A(n12700), .ZN(n12701) );
  MUX2_X1 U15159 ( .A(n14856), .B(n15093), .S(n12571), .Z(n12703) );
  MUX2_X1 U15160 ( .A(n14856), .B(n15093), .S(n12730), .Z(n12702) );
  MUX2_X1 U15161 ( .A(n14837), .B(n15087), .S(n12730), .Z(n12706) );
  MUX2_X1 U15162 ( .A(n15087), .B(n14837), .S(n12730), .Z(n12704) );
  NAND2_X1 U15163 ( .A1(n12904), .A2(n8868), .ZN(n12708) );
  OR2_X1 U15164 ( .A1(n8872), .A2(n15226), .ZN(n12707) );
  MUX2_X1 U15165 ( .A(n14635), .B(n14816), .S(n12571), .Z(n12710) );
  MUX2_X1 U15166 ( .A(n14635), .B(n14816), .S(n12730), .Z(n12709) );
  INV_X1 U15167 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14820) );
  NAND2_X1 U15168 ( .A1(n8947), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12713) );
  INV_X1 U15169 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n12711) );
  OR2_X1 U15170 ( .A1(n8931), .A2(n12711), .ZN(n12712) );
  OAI211_X1 U15171 ( .C1(n12714), .C2(n14820), .A(n12713), .B(n12712), .ZN(
        n14822) );
  NAND2_X1 U15172 ( .A1(n12715), .A2(n8868), .ZN(n12717) );
  INV_X1 U15173 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15217) );
  OR2_X1 U15174 ( .A1(n8872), .A2(n15217), .ZN(n12716) );
  MUX2_X1 U15175 ( .A(n14822), .B(n12571), .S(n15064), .Z(n12718) );
  NAND2_X1 U15176 ( .A1(n12571), .A2(n14822), .ZN(n12732) );
  NAND2_X1 U15177 ( .A1(n12718), .A2(n12732), .ZN(n12781) );
  NAND2_X1 U15178 ( .A1(n14809), .A2(n12719), .ZN(n14840) );
  OAI21_X1 U15179 ( .B1(n12721), .B2(n12720), .A(n14840), .ZN(n12783) );
  AND2_X1 U15180 ( .A1(n12783), .A2(n12786), .ZN(n12779) );
  NAND2_X1 U15181 ( .A1(n12781), .A2(n12779), .ZN(n12774) );
  NAND2_X1 U15182 ( .A1(n12805), .A2(n8868), .ZN(n12723) );
  OR2_X1 U15183 ( .A1(n8872), .A2(n15223), .ZN(n12722) );
  INV_X1 U15184 ( .A(n12724), .ZN(n12728) );
  INV_X1 U15185 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n12727) );
  NAND2_X1 U15186 ( .A1(n8947), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n12726) );
  INV_X1 U15187 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15858) );
  OR2_X1 U15188 ( .A1(n8931), .A2(n15858), .ZN(n12725) );
  OAI211_X1 U15189 ( .C1(n12714), .C2(n12727), .A(n12726), .B(n12725), .ZN(
        n14634) );
  OAI21_X1 U15190 ( .B1(n14822), .B2(n12728), .A(n14634), .ZN(n12729) );
  INV_X1 U15191 ( .A(n12729), .ZN(n12731) );
  MUX2_X1 U15192 ( .A(n14829), .B(n12731), .S(n12730), .Z(n12738) );
  INV_X1 U15193 ( .A(n14634), .ZN(n12744) );
  AOI21_X1 U15194 ( .B1(n12733), .B2(n12732), .A(n12744), .ZN(n12734) );
  AOI21_X1 U15195 ( .B1(n14829), .B2(n12730), .A(n12734), .ZN(n12739) );
  NOR2_X1 U15196 ( .A1(n12738), .A2(n12739), .ZN(n12775) );
  INV_X1 U15197 ( .A(n14822), .ZN(n12735) );
  XNOR2_X1 U15198 ( .A(n15064), .B(n12735), .ZN(n12780) );
  INV_X1 U15199 ( .A(n12780), .ZN(n12737) );
  INV_X1 U15200 ( .A(n12783), .ZN(n12736) );
  AND2_X1 U15201 ( .A1(n12737), .A2(n12736), .ZN(n12776) );
  INV_X1 U15202 ( .A(n12776), .ZN(n12742) );
  INV_X1 U15203 ( .A(n12738), .ZN(n12741) );
  INV_X1 U15204 ( .A(n12739), .ZN(n12740) );
  NOR2_X1 U15205 ( .A1(n12741), .A2(n12740), .ZN(n12777) );
  NOR2_X1 U15206 ( .A1(n12742), .A2(n12777), .ZN(n12743) );
  XNOR2_X1 U15207 ( .A(n14829), .B(n12744), .ZN(n12772) );
  OR2_X1 U15208 ( .A1(n15087), .A2(n14837), .ZN(n12981) );
  INV_X1 U15209 ( .A(n14870), .ZN(n14527) );
  NAND2_X1 U15210 ( .A1(n14860), .A2(n14527), .ZN(n14833) );
  OR2_X1 U15211 ( .A1(n14860), .A2(n14527), .ZN(n12745) );
  INV_X1 U15212 ( .A(n12941), .ZN(n12747) );
  OR2_X1 U15213 ( .A1(n12942), .A2(n12747), .ZN(n15023) );
  NOR2_X1 U15214 ( .A1(n12749), .A2(n12748), .ZN(n12760) );
  AND4_X1 U15215 ( .A1(n12752), .A2(n12751), .A3(n15386), .A4(n12750), .ZN(
        n12755) );
  NAND4_X1 U15216 ( .A1(n12755), .A2(n12754), .A3(n15367), .A4(n12753), .ZN(
        n12757) );
  NOR2_X1 U15217 ( .A1(n12757), .A2(n12756), .ZN(n12759) );
  AND4_X1 U15218 ( .A1(n12761), .A2(n12760), .A3(n12759), .A4(n12758), .ZN(
        n12764) );
  NAND4_X1 U15219 ( .A1(n15023), .A2(n12764), .A3(n12763), .A4(n12762), .ZN(
        n12766) );
  INV_X1 U15220 ( .A(n15016), .ZN(n14554) );
  XNOR2_X1 U15221 ( .A(n15166), .B(n14554), .ZN(n15039) );
  OR4_X1 U15222 ( .A1(n15055), .A2(n12766), .A3(n15039), .A4(n12765), .ZN(
        n12768) );
  INV_X1 U15223 ( .A(n14995), .ZN(n14996) );
  NAND2_X1 U15224 ( .A1(n12767), .A2(n12914), .ZN(n14981) );
  NAND2_X1 U15225 ( .A1(n14955), .A2(n14964), .ZN(n12947) );
  NAND2_X1 U15226 ( .A1(n12949), .A2(n12947), .ZN(n14947) );
  XNOR2_X1 U15227 ( .A(n15143), .B(n14942), .ZN(n14973) );
  INV_X1 U15228 ( .A(n14973), .ZN(n14961) );
  AND4_X1 U15229 ( .A1(n14926), .A2(n6668), .A3(n14947), .A4(n14961), .ZN(
        n12769) );
  XNOR2_X1 U15230 ( .A(n15121), .B(n14930), .ZN(n14910) );
  XNOR2_X1 U15231 ( .A(n15111), .B(n14907), .ZN(n14885) );
  AND4_X1 U15232 ( .A1(n14853), .A2(n12769), .A3(n14910), .A4(n14885), .ZN(
        n12770) );
  XNOR2_X1 U15233 ( .A(n14879), .B(n14887), .ZN(n14880) );
  NAND4_X1 U15234 ( .A1(n12956), .A2(n12770), .A3(n7260), .A4(n14880), .ZN(
        n12771) );
  XNOR2_X1 U15235 ( .A(n12773), .B(n14809), .ZN(n12787) );
  INV_X1 U15236 ( .A(n12774), .ZN(n12778) );
  AOI22_X1 U15237 ( .A1(n12778), .A2(n12777), .B1(n12776), .B2(n12775), .ZN(
        n12785) );
  NAND2_X1 U15238 ( .A1(n12780), .A2(n12779), .ZN(n12782) );
  MUX2_X1 U15239 ( .A(n12783), .B(n12782), .S(n12781), .Z(n12784) );
  OAI211_X1 U15240 ( .C1(n12787), .C2(n12786), .A(n12785), .B(n12784), .ZN(
        n12788) );
  NAND3_X1 U15241 ( .A1(n12790), .A2(n12969), .A3(n15029), .ZN(n12791) );
  OAI211_X1 U15242 ( .C1(n15237), .C2(n12793), .A(n12791), .B(P1_B_REG_SCAN_IN), .ZN(n12792) );
  OAI21_X1 U15243 ( .B1(n12796), .B2(n12795), .A(n12794), .ZN(n12798) );
  XNOR2_X1 U15244 ( .A(n12798), .B(n12797), .ZN(n12804) );
  INV_X1 U15245 ( .A(n12799), .ZN(n12802) );
  NOR4_X1 U15246 ( .A1(P3_U3151), .A2(n9370), .A3(P3_IR_REG_30__SCAN_IN), .A4(
        P3_IR_REG_29__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U15247 ( .A1(n12802), .A2(n12801), .B1(n12800), .B2(SI_31_), .ZN(
        n12803) );
  OAI21_X1 U15248 ( .B1(n12804), .B2(n12962), .A(n12803), .ZN(P3_U3264) );
  INV_X1 U15249 ( .A(n12805), .ZN(n15225) );
  OAI222_X1 U15250 ( .A1(n10996), .A2(n15225), .B1(n12807), .B2(P2_U3088), 
        .C1(n12806), .C2(n14478), .ZN(P2_U3297) );
  OAI21_X1 U15251 ( .B1(n12810), .B2(n12809), .A(n12808), .ZN(n12811) );
  NAND2_X1 U15252 ( .A1(n12811), .A2(n14621), .ZN(n12816) );
  OAI22_X1 U15253 ( .A1(n12813), .A2(n14941), .B1(n12812), .B2(n14943), .ZN(
        n15388) );
  AOI22_X1 U15254 ( .A1(n14571), .A2(n15388), .B1(n12814), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n12815) );
  OAI211_X1 U15255 ( .C1(n15418), .C2(n14633), .A(n12816), .B(n12815), .ZN(
        P1_U3237) );
  NAND2_X1 U15256 ( .A1(n14082), .A2(n14064), .ZN(n12819) );
  NAND2_X1 U15257 ( .A1(n14322), .A2(n14065), .ZN(n12821) );
  INV_X1 U15258 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n12844) );
  AOI211_X1 U15259 ( .C1(n13875), .C2(n14038), .A(n8582), .B(n14027), .ZN(
        n12853) );
  AND2_X1 U15260 ( .A1(n12823), .A2(n12824), .ZN(n14055) );
  AND2_X1 U15261 ( .A1(n14057), .A2(n14055), .ZN(n12829) );
  NAND2_X1 U15262 ( .A1(n12825), .A2(n12824), .ZN(n12827) );
  NAND2_X1 U15263 ( .A1(n12827), .A2(n12826), .ZN(n14056) );
  NAND2_X1 U15264 ( .A1(n14056), .A2(n14057), .ZN(n12828) );
  NOR2_X1 U15265 ( .A1(n14413), .A2(n14046), .ZN(n14042) );
  INV_X1 U15266 ( .A(n14045), .ZN(n12831) );
  NAND3_X1 U15267 ( .A1(n12831), .A2(n13931), .A3(n14307), .ZN(n12843) );
  INV_X1 U15268 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n15873) );
  NAND2_X1 U15269 ( .A1(n12832), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n12835) );
  NAND2_X1 U15270 ( .A1(n12833), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n12834) );
  OAI211_X1 U15271 ( .C1(n12836), .C2(n15873), .A(n12835), .B(n12834), .ZN(
        n13960) );
  INV_X1 U15272 ( .A(n13960), .ZN(n13869) );
  OAI22_X1 U15273 ( .A1(n14065), .A2(n14116), .B1(n13869), .B2(n12837), .ZN(
        n12838) );
  INV_X1 U15274 ( .A(n12838), .ZN(n12842) );
  INV_X1 U15275 ( .A(n13931), .ZN(n12840) );
  NAND4_X1 U15276 ( .A1(n13931), .A2(n14040), .A3(n13962), .A4(n14307), .ZN(
        n12841) );
  MUX2_X1 U15277 ( .A(n12844), .B(n12846), .S(n15659), .Z(n12845) );
  OAI21_X1 U15278 ( .B1(n12857), .B2(n14461), .A(n12845), .ZN(P2_U3496) );
  INV_X1 U15279 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n12847) );
  MUX2_X1 U15280 ( .A(n12847), .B(n12846), .S(n15670), .Z(n12848) );
  OAI21_X1 U15281 ( .B1(n12857), .B2(n14401), .A(n12848), .ZN(P2_U3528) );
  NOR2_X1 U15282 ( .A1(n13874), .A2(n14275), .ZN(n12852) );
  OAI22_X1 U15283 ( .A1(n12850), .A2(n14290), .B1(n12849), .B2(n14293), .ZN(
        n12851) );
  AOI211_X1 U15284 ( .C1(n12853), .C2(n14282), .A(n12852), .B(n12851), .ZN(
        n12856) );
  NAND2_X1 U15285 ( .A1(n12854), .A2(n14293), .ZN(n12855) );
  OAI211_X1 U15286 ( .C1(n12857), .C2(n14279), .A(n12856), .B(n12855), .ZN(
        P2_U3236) );
  AOI21_X1 U15287 ( .B1(n12865), .B2(n13369), .A(n12858), .ZN(n12864) );
  INV_X1 U15288 ( .A(n12864), .ZN(n12860) );
  NAND3_X1 U15289 ( .A1(n12864), .A2(n13022), .A3(n12863), .ZN(n12872) );
  INV_X1 U15290 ( .A(n12865), .ZN(n12870) );
  NAND2_X1 U15291 ( .A1(n12866), .A2(n13369), .ZN(n12869) );
  AOI22_X1 U15292 ( .A1(n12870), .A2(n12869), .B1(n12868), .B2(n12867), .ZN(
        n12871) );
  XNOR2_X1 U15293 ( .A(n12874), .B(n9715), .ZN(n12875) );
  XNOR2_X1 U15294 ( .A(n12875), .B(n13094), .ZN(n13028) );
  NAND2_X1 U15295 ( .A1(n13027), .A2(n13028), .ZN(n12878) );
  INV_X1 U15296 ( .A(n12875), .ZN(n12876) );
  NAND2_X1 U15297 ( .A1(n12876), .A2(n13094), .ZN(n12877) );
  XNOR2_X1 U15298 ( .A(n13327), .B(n9722), .ZN(n12879) );
  XNOR2_X1 U15299 ( .A(n12879), .B(n13342), .ZN(n13088) );
  INV_X1 U15300 ( .A(n12879), .ZN(n12880) );
  NOR2_X1 U15301 ( .A1(n12880), .A2(n13342), .ZN(n12881) );
  XNOR2_X1 U15302 ( .A(n12991), .B(n9722), .ZN(n12882) );
  XNOR2_X1 U15303 ( .A(n12882), .B(n12888), .ZN(n12992) );
  INV_X1 U15304 ( .A(n12882), .ZN(n12883) );
  XNOR2_X1 U15305 ( .A(n12884), .B(n9722), .ZN(n12885) );
  NOR2_X1 U15306 ( .A1(n12886), .A2(n13072), .ZN(n12890) );
  AOI22_X1 U15307 ( .A1(n13303), .A2(n13090), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12887) );
  OAI21_X1 U15308 ( .B1(n12888), .B2(n13093), .A(n12887), .ZN(n12889) );
  AOI211_X1 U15309 ( .C1(n10178), .C2(n13096), .A(n12890), .B(n12889), .ZN(
        n12891) );
  OAI21_X1 U15310 ( .B1(n12892), .B2(n13098), .A(n12891), .ZN(P3_U3160) );
  AOI21_X1 U15311 ( .B1(n12893), .B2(n12894), .A(n13695), .ZN(n12897) );
  NOR3_X1 U15312 ( .A1(n12895), .A2(n14119), .A3(n13697), .ZN(n12896) );
  NOR2_X1 U15313 ( .A1(n12897), .A2(n12896), .ZN(n12903) );
  AOI22_X1 U15314 ( .A1(n14090), .A2(n13701), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12899) );
  OAI21_X1 U15315 ( .B1(n12900), .B2(n13703), .A(n12899), .ZN(n12901) );
  AOI21_X1 U15316 ( .B1(n13859), .B2(n13693), .A(n12901), .ZN(n12902) );
  OAI21_X1 U15317 ( .B1(n12903), .B2(n12898), .A(n12902), .ZN(P2_U3197) );
  INV_X1 U15318 ( .A(n12904), .ZN(n15228) );
  OAI222_X1 U15319 ( .A1(n10996), .A2(n15228), .B1(n12906), .B2(P2_U3088), 
        .C1(n12905), .C2(n14478), .ZN(P2_U3298) );
  NAND2_X1 U15320 ( .A1(n12908), .A2(n12907), .ZN(n15046) );
  NAND2_X1 U15321 ( .A1(n15046), .A2(n15045), .ZN(n15044) );
  NAND2_X1 U15322 ( .A1(n15044), .A2(n12909), .ZN(n15028) );
  NAND2_X1 U15323 ( .A1(n15166), .A2(n14554), .ZN(n12910) );
  INV_X1 U15324 ( .A(n15032), .ZN(n14540) );
  AND2_X1 U15325 ( .A1(n15161), .A2(n14540), .ZN(n12911) );
  OR2_X1 U15326 ( .A1(n15161), .A2(n14540), .ZN(n12912) );
  INV_X1 U15327 ( .A(n15015), .ZN(n12913) );
  OR2_X1 U15328 ( .A1(n15143), .A2(n14942), .ZN(n12915) );
  INV_X1 U15329 ( .A(n14964), .ZN(n14580) );
  INV_X1 U15330 ( .A(n14930), .ZN(n14889) );
  INV_X1 U15331 ( .A(n14887), .ZN(n14610) );
  OR2_X1 U15332 ( .A1(n14879), .A2(n14610), .ZN(n12916) );
  INV_X1 U15333 ( .A(n14907), .ZN(n14526) );
  OR2_X1 U15334 ( .A1(n15111), .A2(n14526), .ZN(n14867) );
  OAI211_X1 U15335 ( .C1(n14889), .C2(n15121), .A(n12916), .B(n14867), .ZN(
        n12918) );
  OR2_X1 U15336 ( .A1(n12918), .A2(n12917), .ZN(n12927) );
  OR2_X1 U15337 ( .A1(n12918), .A2(n14902), .ZN(n12925) );
  AND2_X1 U15338 ( .A1(n15121), .A2(n14889), .ZN(n14865) );
  NAND2_X1 U15339 ( .A1(n14865), .A2(n14867), .ZN(n12920) );
  AOI21_X1 U15340 ( .B1(n15111), .B2(n14526), .A(n14610), .ZN(n12919) );
  NAND2_X1 U15341 ( .A1(n12920), .A2(n12919), .ZN(n12921) );
  NAND2_X1 U15342 ( .A1(n12921), .A2(n14879), .ZN(n12924) );
  NAND3_X1 U15343 ( .A1(n15111), .A2(n14526), .A3(n14610), .ZN(n12923) );
  NAND4_X1 U15344 ( .A1(n14867), .A2(n14889), .A3(n14610), .A4(n15121), .ZN(
        n12922) );
  AOI21_X2 U15345 ( .B1(n12932), .B2(n15389), .A(n12931), .ZN(n15091) );
  INV_X1 U15346 ( .A(n15156), .ZN(n15007) );
  INV_X1 U15347 ( .A(n14955), .ZN(n15135) );
  INV_X1 U15348 ( .A(n14879), .ZN(n15108) );
  INV_X1 U15349 ( .A(n14860), .ZN(n15100) );
  NAND2_X1 U15350 ( .A1(n14875), .A2(n15100), .ZN(n14855) );
  AOI21_X1 U15351 ( .B1(n14841), .B2(n15087), .A(n15397), .ZN(n12933) );
  NAND2_X1 U15352 ( .A1(n12933), .A2(n14817), .ZN(n15089) );
  AOI22_X1 U15353 ( .A1(n12934), .A2(n15392), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15405), .ZN(n12936) );
  NAND2_X1 U15354 ( .A1(n15087), .A2(n14954), .ZN(n12935) );
  OAI211_X1 U15355 ( .C1(n15089), .C2(n14935), .A(n12936), .B(n12935), .ZN(
        n12937) );
  INV_X1 U15356 ( .A(n12937), .ZN(n12959) );
  NAND2_X1 U15357 ( .A1(n15175), .A2(n14638), .ZN(n15056) );
  AND2_X1 U15358 ( .A1(n15055), .A2(n15056), .ZN(n12938) );
  OR2_X1 U15359 ( .A1(n15171), .A2(n15030), .ZN(n12940) );
  OR2_X1 U15360 ( .A1(n15150), .A2(n14993), .ZN(n12944) );
  AND2_X1 U15361 ( .A1(n14978), .A2(n12944), .ZN(n12945) );
  NAND2_X1 U15362 ( .A1(n15143), .A2(n14637), .ZN(n12946) );
  INV_X1 U15363 ( .A(n12947), .ZN(n12948) );
  INV_X1 U15364 ( .A(n12949), .ZN(n14925) );
  AOI22_X1 U15365 ( .A1(n14922), .A2(n14925), .B1(n14944), .B2(n15129), .ZN(
        n12950) );
  NAND2_X1 U15366 ( .A1(n15121), .A2(n14930), .ZN(n12951) );
  OR2_X1 U15367 ( .A1(n15111), .A2(n14907), .ZN(n12952) );
  NAND2_X1 U15368 ( .A1(n14879), .A2(n14887), .ZN(n12953) );
  NAND2_X1 U15369 ( .A1(n14860), .A2(n14870), .ZN(n12954) );
  NOR2_X1 U15370 ( .A1(n15093), .A2(n14856), .ZN(n12979) );
  NAND2_X1 U15371 ( .A1(n12955), .A2(n12928), .ZN(n15086) );
  INV_X1 U15372 ( .A(n12955), .ZN(n12957) );
  NAND2_X1 U15373 ( .A1(n12957), .A2(n12956), .ZN(n15085) );
  NAND3_X1 U15374 ( .A1(n15086), .A2(n15381), .A3(n15085), .ZN(n12958) );
  OAI211_X1 U15375 ( .C1(n15091), .C2(n15405), .A(n12959), .B(n12958), .ZN(
        P1_U3265) );
  OAI222_X1 U15376 ( .A1(n12962), .A2(n12961), .B1(n13550), .B2(n12960), .C1(
        P3_U3151), .C2(n10042), .ZN(P3_U3274) );
  INV_X1 U15377 ( .A(n12963), .ZN(n12965) );
  OAI222_X1 U15378 ( .A1(n13550), .A2(n15965), .B1(n12962), .B2(n12965), .C1(
        n12964), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U15379 ( .A(n14837), .ZN(n12966) );
  NOR2_X1 U15380 ( .A1(n15087), .A2(n12966), .ZN(n15081) );
  INV_X1 U15381 ( .A(n15087), .ZN(n12967) );
  NOR2_X1 U15382 ( .A1(n12967), .A2(n14837), .ZN(n15076) );
  INV_X1 U15383 ( .A(n15076), .ZN(n15079) );
  OAI21_X1 U15384 ( .B1(n15083), .B2(n15081), .A(n15079), .ZN(n12968) );
  XNOR2_X1 U15385 ( .A(n12968), .B(n15077), .ZN(n12990) );
  NAND2_X1 U15386 ( .A1(n15392), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n12972) );
  NAND2_X1 U15387 ( .A1(n12969), .A2(P1_B_REG_SCAN_IN), .ZN(n12970) );
  AND2_X1 U15388 ( .A1(n15031), .A2(n12970), .ZN(n14821) );
  NAND2_X1 U15389 ( .A1(n14634), .A2(n14821), .ZN(n15069) );
  OAI22_X1 U15390 ( .A1(n12973), .A2(n12972), .B1(n15069), .B2(n12971), .ZN(
        n12975) );
  NAND2_X1 U15391 ( .A1(n14837), .A2(n15029), .ZN(n15070) );
  NOR2_X1 U15392 ( .A1(n15070), .A2(n15405), .ZN(n12974) );
  AOI211_X1 U15393 ( .C1(n15405), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12975), 
        .B(n12974), .ZN(n12976) );
  OAI21_X1 U15394 ( .B1(n15071), .B2(n15394), .A(n12976), .ZN(n12988) );
  INV_X1 U15395 ( .A(n12983), .ZN(n12977) );
  NOR2_X1 U15396 ( .A1(n15080), .A2(n12977), .ZN(n12978) );
  INV_X1 U15397 ( .A(n12979), .ZN(n12980) );
  NAND2_X1 U15398 ( .A1(n12981), .A2(n12980), .ZN(n12987) );
  AOI21_X1 U15399 ( .B1(n12983), .B2(n12987), .A(n15080), .ZN(n12982) );
  AOI21_X1 U15400 ( .B1(n12983), .B2(n15080), .A(n12982), .ZN(n12984) );
  XNOR2_X1 U15401 ( .A(n12993), .B(n12992), .ZN(n12994) );
  NAND2_X1 U15402 ( .A1(n12994), .A2(n13058), .ZN(n12999) );
  AOI22_X1 U15403 ( .A1(n13315), .A2(n13090), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12995) );
  OAI21_X1 U15404 ( .B1(n12996), .B2(n13093), .A(n12995), .ZN(n12997) );
  AOI21_X1 U15405 ( .B1(n13310), .B2(n13089), .A(n12997), .ZN(n12998) );
  OAI211_X1 U15406 ( .C1(n13501), .C2(n13081), .A(n12999), .B(n12998), .ZN(
        P3_U3154) );
  XNOR2_X1 U15407 ( .A(n13000), .B(n13073), .ZN(n13001) );
  XNOR2_X1 U15408 ( .A(n13002), .B(n13001), .ZN(n13007) );
  AOI22_X1 U15409 ( .A1(n13397), .A2(n13069), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13004) );
  NAND2_X1 U15410 ( .A1(n13374), .A2(n13090), .ZN(n13003) );
  OAI211_X1 U15411 ( .C1(n13031), .C2(n13072), .A(n13004), .B(n13003), .ZN(
        n13005) );
  AOI21_X1 U15412 ( .B1(n13373), .B2(n13096), .A(n13005), .ZN(n13006) );
  OAI21_X1 U15413 ( .B1(n13007), .B2(n13098), .A(n13006), .ZN(P3_U3156) );
  OAI211_X1 U15414 ( .C1(n13010), .C2(n13009), .A(n13008), .B(n13058), .ZN(
        n13015) );
  NAND2_X1 U15415 ( .A1(n13395), .A2(n13089), .ZN(n13012) );
  OAI211_X1 U15416 ( .C1(n13413), .C2(n13093), .A(n13012), .B(n13011), .ZN(
        n13013) );
  AOI21_X1 U15417 ( .B1(n13409), .B2(n13090), .A(n13013), .ZN(n13014) );
  OAI211_X1 U15418 ( .C1(n13081), .C2(n13535), .A(n13015), .B(n13014), .ZN(
        P3_U3159) );
  INV_X1 U15419 ( .A(n13016), .ZN(n13017) );
  AOI21_X1 U15420 ( .B1(n13019), .B2(n13018), .A(n13017), .ZN(n13026) );
  AOI22_X1 U15421 ( .A1(n13395), .A2(n13069), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13021) );
  NAND2_X1 U15422 ( .A1(n13401), .A2(n13090), .ZN(n13020) );
  OAI211_X1 U15423 ( .C1(n13022), .C2(n13072), .A(n13021), .B(n13020), .ZN(
        n13023) );
  AOI21_X1 U15424 ( .B1(n13024), .B2(n13096), .A(n13023), .ZN(n13025) );
  OAI21_X1 U15425 ( .B1(n13026), .B2(n13098), .A(n13025), .ZN(P3_U3163) );
  XOR2_X1 U15426 ( .A(n13028), .B(n13027), .Z(n13034) );
  NAND2_X1 U15427 ( .A1(n13342), .A2(n13089), .ZN(n13030) );
  AOI22_X1 U15428 ( .A1(n13346), .A2(n13090), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13029) );
  OAI211_X1 U15429 ( .C1(n13031), .C2(n13093), .A(n13030), .B(n13029), .ZN(
        n13032) );
  AOI21_X1 U15430 ( .B1(n13507), .B2(n13096), .A(n13032), .ZN(n13033) );
  OAI21_X1 U15431 ( .B1(n13034), .B2(n13098), .A(n13033), .ZN(P3_U3165) );
  XNOR2_X1 U15432 ( .A(n13035), .B(n13049), .ZN(n13036) );
  XNOR2_X1 U15433 ( .A(n13037), .B(n13036), .ZN(n13045) );
  NAND2_X1 U15434 ( .A1(n13089), .A2(n13102), .ZN(n13038) );
  NAND2_X1 U15435 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13236)
         );
  OAI211_X1 U15436 ( .C1(n13039), .C2(n13093), .A(n13038), .B(n13236), .ZN(
        n13040) );
  AOI21_X1 U15437 ( .B1(n13041), .B2(n13090), .A(n13040), .ZN(n13044) );
  NAND2_X1 U15438 ( .A1(n13042), .A2(n13096), .ZN(n13043) );
  OAI211_X1 U15439 ( .C1(n13045), .C2(n13098), .A(n13044), .B(n13043), .ZN(
        P3_U3166) );
  XNOR2_X1 U15440 ( .A(n13046), .B(n13102), .ZN(n13047) );
  XNOR2_X1 U15441 ( .A(n13048), .B(n13047), .ZN(n13056) );
  NAND2_X1 U15442 ( .A1(n13069), .A2(n13049), .ZN(n13050) );
  NAND2_X1 U15443 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13259)
         );
  OAI211_X1 U15444 ( .C1(n13413), .C2(n13072), .A(n13050), .B(n13259), .ZN(
        n13053) );
  NOR2_X1 U15445 ( .A1(n13051), .A2(n13081), .ZN(n13052) );
  AOI211_X1 U15446 ( .C1(n13054), .C2(n13090), .A(n13053), .B(n13052), .ZN(
        n13055) );
  OAI21_X1 U15447 ( .B1(n13056), .B2(n13098), .A(n13055), .ZN(P3_U3168) );
  INV_X1 U15448 ( .A(n13057), .ZN(n13067) );
  OAI211_X1 U15449 ( .C1(n13061), .C2(n13060), .A(n13059), .B(n13058), .ZN(
        n13066) );
  AOI22_X1 U15450 ( .A1(n13101), .A2(n13069), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13062) );
  OAI21_X1 U15451 ( .B1(n9989), .B2(n13072), .A(n13062), .ZN(n13063) );
  AOI21_X1 U15452 ( .B1(n13064), .B2(n13090), .A(n13063), .ZN(n13065) );
  OAI211_X1 U15453 ( .C1(n13067), .C2(n13081), .A(n13066), .B(n13065), .ZN(
        P3_U3173) );
  XNOR2_X1 U15454 ( .A(n13068), .B(n13397), .ZN(n13076) );
  AOI22_X1 U15455 ( .A1(n13384), .A2(n13069), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13071) );
  NAND2_X1 U15456 ( .A1(n13388), .A2(n13090), .ZN(n13070) );
  OAI211_X1 U15457 ( .C1(n13073), .C2(n13072), .A(n13071), .B(n13070), .ZN(
        n13074) );
  AOI21_X1 U15458 ( .B1(n13521), .B2(n13096), .A(n13074), .ZN(n13075) );
  OAI21_X1 U15459 ( .B1(n13076), .B2(n13098), .A(n13075), .ZN(P3_U3175) );
  XOR2_X1 U15460 ( .A(n13413), .B(n13077), .Z(n13078) );
  XNOR2_X1 U15461 ( .A(n13079), .B(n13078), .ZN(n13086) );
  NAND2_X1 U15462 ( .A1(n13101), .A2(n13089), .ZN(n13080) );
  NAND2_X1 U15463 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13272)
         );
  OAI211_X1 U15464 ( .C1(n13430), .C2(n13093), .A(n13080), .B(n13272), .ZN(
        n13084) );
  NOR2_X1 U15465 ( .A1(n13082), .A2(n13081), .ZN(n13083) );
  AOI211_X1 U15466 ( .C1(n13434), .C2(n13090), .A(n13084), .B(n13083), .ZN(
        n13085) );
  OAI21_X1 U15467 ( .B1(n13086), .B2(n13098), .A(n13085), .ZN(P3_U3178) );
  XOR2_X1 U15468 ( .A(n13088), .B(n13087), .Z(n13099) );
  NAND2_X1 U15469 ( .A1(n13324), .A2(n13089), .ZN(n13092) );
  AOI22_X1 U15470 ( .A1(n13328), .A2(n13090), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13091) );
  OAI211_X1 U15471 ( .C1(n13094), .C2(n13093), .A(n13092), .B(n13091), .ZN(
        n13095) );
  AOI21_X1 U15472 ( .B1(n13327), .B2(n13096), .A(n13095), .ZN(n13097) );
  OAI21_X1 U15473 ( .B1(n13099), .B2(n13098), .A(n13097), .ZN(P3_U3180) );
  MUX2_X1 U15474 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13290), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15475 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n13100), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U15476 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n13300), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15477 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13310), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15478 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13324), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15479 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13342), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15480 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13369), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15481 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13385), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U15482 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13397), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15483 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13384), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15484 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13395), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15485 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13101), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15486 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13102), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15487 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13103), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15488 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13104), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15489 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13105), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15490 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13106), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15491 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13107), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15492 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13108), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15493 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13109), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15494 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13110), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15495 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13111), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15496 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13112), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15497 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13113), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15498 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13114), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15499 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13115), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15500 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n7138), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15501 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n13118), .S(P3_U3897), .Z(
        P3_U3491) );
  OAI21_X1 U15502 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n13120), .A(n13119), .ZN(
        n13121) );
  AOI22_X1 U15503 ( .A1(n13279), .A2(n13122), .B1(n13209), .B2(n13121), .ZN(
        n13137) );
  AOI22_X1 U15504 ( .A1(n15694), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n13136) );
  INV_X1 U15505 ( .A(n13123), .ZN(n13127) );
  INV_X1 U15506 ( .A(n13124), .ZN(n13126) );
  NOR3_X1 U15507 ( .A1(n13127), .A2(n13126), .A3(n13125), .ZN(n13130) );
  INV_X1 U15508 ( .A(n13128), .ZN(n13129) );
  OAI21_X1 U15509 ( .B1(n13130), .B2(n13129), .A(n13248), .ZN(n13135) );
  OAI21_X1 U15510 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n13132), .A(n13131), .ZN(
        n13133) );
  NAND2_X1 U15511 ( .A1(n13284), .A2(n13133), .ZN(n13134) );
  NAND4_X1 U15512 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n13134), .ZN(
        P3_U3185) );
  AND3_X1 U15513 ( .A1(n13140), .A2(n13139), .A3(n13138), .ZN(n13141) );
  OAI21_X1 U15514 ( .B1(n13142), .B2(n13141), .A(n13209), .ZN(n13159) );
  NOR2_X1 U15515 ( .A1(n13261), .A2(n13143), .ZN(n13144) );
  AOI211_X1 U15516 ( .C1(n15694), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n13145), .B(
        n13144), .ZN(n13158) );
  NOR3_X1 U15517 ( .A1(n13148), .A2(n6827), .A3(n13147), .ZN(n13150) );
  OAI21_X1 U15518 ( .B1(n13150), .B2(n13149), .A(n13248), .ZN(n13157) );
  AND3_X1 U15519 ( .A1(n13153), .A2(n13152), .A3(n13151), .ZN(n13154) );
  OAI21_X1 U15520 ( .B1(n13155), .B2(n13154), .A(n13284), .ZN(n13156) );
  NAND4_X1 U15521 ( .A1(n13159), .A2(n13158), .A3(n13157), .A4(n13156), .ZN(
        P3_U3188) );
  AOI21_X1 U15522 ( .B1(n13161), .B2(n13160), .A(n6711), .ZN(n13173) );
  OAI21_X1 U15523 ( .B1(n13163), .B2(n13162), .A(n13182), .ZN(n13168) );
  NAND2_X1 U15524 ( .A1(n15694), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n13164) );
  OAI211_X1 U15525 ( .C1(n13261), .C2(n13166), .A(n13165), .B(n13164), .ZN(
        n13167) );
  AOI21_X1 U15526 ( .B1(n13168), .B2(n13248), .A(n13167), .ZN(n13172) );
  NAND2_X1 U15527 ( .A1(n13170), .A2(n13284), .ZN(n13171) );
  OAI211_X1 U15528 ( .C1(n13173), .C2(n13288), .A(n13172), .B(n13171), .ZN(
        P3_U3193) );
  NOR2_X1 U15529 ( .A1(n13175), .A2(n13174), .ZN(n13178) );
  INV_X1 U15530 ( .A(n13176), .ZN(n13177) );
  AOI21_X1 U15531 ( .B1(n13178), .B2(n13169), .A(n13177), .ZN(n13194) );
  INV_X1 U15532 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15253) );
  OAI21_X1 U15533 ( .B1(n13273), .B2(n15253), .A(n13179), .ZN(n13186) );
  INV_X1 U15534 ( .A(n13201), .ZN(n13184) );
  AOI21_X1 U15535 ( .B1(n13182), .B2(n13181), .A(n13180), .ZN(n13183) );
  NOR3_X1 U15536 ( .A1(n13184), .A2(n13183), .A3(n13277), .ZN(n13185) );
  AOI211_X1 U15537 ( .C1(n13187), .C2(n13279), .A(n13186), .B(n13185), .ZN(
        n13193) );
  OAI21_X1 U15538 ( .B1(n13190), .B2(n13189), .A(n13188), .ZN(n13191) );
  NAND2_X1 U15539 ( .A1(n13191), .A2(n13209), .ZN(n13192) );
  OAI211_X1 U15540 ( .C1(n13194), .C2(n13242), .A(n13193), .B(n13192), .ZN(
        P3_U3194) );
  INV_X1 U15541 ( .A(n13195), .ZN(n13196) );
  AOI21_X1 U15542 ( .B1(n15738), .B2(n13197), .A(n13196), .ZN(n13213) );
  INV_X1 U15543 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15264) );
  OAI21_X1 U15544 ( .B1(n13273), .B2(n15264), .A(n13198), .ZN(n13206) );
  AOI21_X1 U15545 ( .B1(n13201), .B2(n13200), .A(n13199), .ZN(n13202) );
  INV_X1 U15546 ( .A(n13202), .ZN(n13204) );
  AOI21_X1 U15547 ( .B1(n13204), .B2(n13203), .A(n13277), .ZN(n13205) );
  AOI211_X1 U15548 ( .C1(n13207), .C2(n13279), .A(n13206), .B(n13205), .ZN(
        n13212) );
  OAI21_X1 U15549 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n6717), .A(n13208), .ZN(
        n13210) );
  NAND2_X1 U15550 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  OAI211_X1 U15551 ( .C1(n13213), .C2(n13242), .A(n13212), .B(n13211), .ZN(
        P3_U3195) );
  XOR2_X1 U15552 ( .A(P3_REG2_REG_15__SCAN_IN), .B(n13214), .Z(n13225) );
  OAI21_X1 U15553 ( .B1(n6619), .B2(P3_REG1_REG_15__SCAN_IN), .A(n13241), .ZN(
        n13223) );
  OAI211_X1 U15554 ( .C1(n13217), .C2(n13216), .A(n13215), .B(n13248), .ZN(
        n13220) );
  AOI21_X1 U15555 ( .B1(n15694), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13218), 
        .ZN(n13219) );
  OAI211_X1 U15556 ( .C1(n13261), .C2(n13221), .A(n13220), .B(n13219), .ZN(
        n13222) );
  AOI21_X1 U15557 ( .B1(n13223), .B2(n13284), .A(n13222), .ZN(n13224) );
  OAI21_X1 U15558 ( .B1(n13225), .B2(n13288), .A(n13224), .ZN(P3_U3197) );
  OAI21_X1 U15559 ( .B1(n13228), .B2(n13227), .A(n13226), .ZN(n13229) );
  INV_X1 U15560 ( .A(n13229), .ZN(n13250) );
  INV_X1 U15561 ( .A(n13230), .ZN(n13232) );
  NAND2_X1 U15562 ( .A1(n13232), .A2(n13231), .ZN(n13233) );
  XNOR2_X1 U15563 ( .A(n13234), .B(n13233), .ZN(n13247) );
  NAND2_X1 U15564 ( .A1(n15694), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n13235) );
  OAI211_X1 U15565 ( .C1(n13261), .C2(n13237), .A(n13236), .B(n13235), .ZN(
        n13246) );
  INV_X1 U15566 ( .A(n13238), .ZN(n13240) );
  NAND3_X1 U15567 ( .A1(n13241), .A2(n13240), .A3(n13239), .ZN(n13243) );
  AOI21_X1 U15568 ( .B1(n13244), .B2(n13243), .A(n13242), .ZN(n13245) );
  AOI211_X1 U15569 ( .C1(n13248), .C2(n13247), .A(n13246), .B(n13245), .ZN(
        n13249) );
  OAI21_X1 U15570 ( .B1(n13250), .B2(n13288), .A(n13249), .ZN(P3_U3198) );
  INV_X1 U15571 ( .A(n13269), .ZN(n13251) );
  AOI21_X1 U15572 ( .B1(n13253), .B2(n13252), .A(n13251), .ZN(n13266) );
  OAI21_X1 U15573 ( .B1(n6969), .B2(P3_REG1_REG_17__SCAN_IN), .A(n13283), .ZN(
        n13264) );
  AOI211_X1 U15574 ( .C1(n13257), .C2(n13256), .A(n13277), .B(n13255), .ZN(
        n13263) );
  NAND2_X1 U15575 ( .A1(n15694), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n13258) );
  OAI211_X1 U15576 ( .C1(n13261), .C2(n13260), .A(n13259), .B(n13258), .ZN(
        n13262) );
  AOI211_X1 U15577 ( .C1(n13264), .C2(n13284), .A(n13263), .B(n13262), .ZN(
        n13265) );
  OAI21_X1 U15578 ( .B1(n13266), .B2(n13288), .A(n13265), .ZN(P3_U3199) );
  INV_X1 U15579 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15319) );
  OAI21_X1 U15580 ( .B1(n13273), .B2(n15319), .A(n13272), .ZN(n13278) );
  AND3_X1 U15581 ( .A1(n13283), .A2(n13282), .A3(n13281), .ZN(n13285) );
  OAI21_X1 U15582 ( .B1(n13286), .B2(n13285), .A(n13284), .ZN(n13287) );
  INV_X1 U15583 ( .A(n12478), .ZN(n13491) );
  AOI21_X1 U15584 ( .B1(n13489), .B2(n13405), .A(n13291), .ZN(n13294) );
  NAND2_X1 U15585 ( .A1(n15688), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13292) );
  OAI211_X1 U15586 ( .C1(n13491), .C2(n13403), .A(n13294), .B(n13292), .ZN(
        P3_U3202) );
  NAND2_X1 U15587 ( .A1(n15688), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13293) );
  OAI211_X1 U15588 ( .C1(n13494), .C2(n13403), .A(n13294), .B(n13293), .ZN(
        P3_U3203) );
  XNOR2_X1 U15589 ( .A(n13295), .B(n13296), .ZN(n13445) );
  INV_X1 U15590 ( .A(n13445), .ZN(n13307) );
  AOI21_X1 U15591 ( .B1(n13297), .B2(n13296), .A(n13428), .ZN(n13299) );
  NAND2_X1 U15592 ( .A1(n13299), .A2(n13298), .ZN(n13302) );
  AOI22_X1 U15593 ( .A1(n13300), .A2(n13396), .B1(n13352), .B2(n13324), .ZN(
        n13301) );
  NAND2_X1 U15594 ( .A1(n13302), .A2(n13301), .ZN(n13447) );
  AOI22_X1 U15595 ( .A1(n13303), .A2(n15675), .B1(n15688), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13304) );
  OAI21_X1 U15596 ( .B1(n13497), .B2(n13403), .A(n13304), .ZN(n13305) );
  AOI21_X1 U15597 ( .B1(n13447), .B2(n13405), .A(n13305), .ZN(n13306) );
  OAI21_X1 U15598 ( .B1(n13441), .B2(n13307), .A(n13306), .ZN(P3_U3205) );
  AOI22_X1 U15599 ( .A1(n13310), .A2(n13396), .B1(n13352), .B2(n13342), .ZN(
        n13314) );
  INV_X1 U15600 ( .A(n13313), .ZN(n13368) );
  INV_X1 U15601 ( .A(n13449), .ZN(n13319) );
  AOI22_X1 U15602 ( .A1(n13315), .A2(n15675), .B1(n15688), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13316) );
  OAI21_X1 U15603 ( .B1(n13501), .B2(n13403), .A(n13316), .ZN(n13317) );
  AOI21_X1 U15604 ( .B1(n13450), .B2(n13377), .A(n13317), .ZN(n13318) );
  OAI21_X1 U15605 ( .B1(n13319), .B2(n15688), .A(n13318), .ZN(P3_U3206) );
  XNOR2_X1 U15606 ( .A(n13320), .B(n13321), .ZN(n13326) );
  AOI22_X1 U15607 ( .A1(n13324), .A2(n13396), .B1(n13352), .B2(n13353), .ZN(
        n13325) );
  INV_X1 U15608 ( .A(n13452), .ZN(n13332) );
  INV_X1 U15609 ( .A(n13327), .ZN(n13504) );
  AOI22_X1 U15610 ( .A1(n13328), .A2(n15675), .B1(n15688), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13329) );
  OAI21_X1 U15611 ( .B1(n13504), .B2(n13403), .A(n13329), .ZN(n13330) );
  AOI21_X1 U15612 ( .B1(n13453), .B2(n13377), .A(n13330), .ZN(n13331) );
  OAI21_X1 U15613 ( .B1(n13332), .B2(n15688), .A(n13331), .ZN(P3_U3207) );
  OAI21_X1 U15614 ( .B1(n13334), .B2(n13338), .A(n13333), .ZN(n13335) );
  INV_X1 U15615 ( .A(n13335), .ZN(n13510) );
  NAND2_X1 U15616 ( .A1(n13337), .A2(n13336), .ZN(n13339) );
  NAND2_X1 U15617 ( .A1(n13339), .A2(n13338), .ZN(n13340) );
  NAND3_X1 U15618 ( .A1(n13341), .A2(n13398), .A3(n13340), .ZN(n13344) );
  AOI22_X1 U15619 ( .A1(n13342), .A2(n13396), .B1(n13352), .B2(n13369), .ZN(
        n13343) );
  MUX2_X1 U15620 ( .A(n13506), .B(n13345), .S(n15688), .Z(n13348) );
  AOI22_X1 U15621 ( .A1(n13507), .A2(n13438), .B1(n15675), .B2(n13346), .ZN(
        n13347) );
  OAI211_X1 U15622 ( .C1(n13510), .C2(n13441), .A(n13348), .B(n13347), .ZN(
        P3_U3208) );
  XNOR2_X1 U15623 ( .A(n13349), .B(n13351), .ZN(n13460) );
  INV_X1 U15624 ( .A(n13460), .ZN(n13364) );
  XNOR2_X1 U15625 ( .A(n13350), .B(n13351), .ZN(n13356) );
  NAND2_X1 U15626 ( .A1(n13460), .A2(n13368), .ZN(n13355) );
  AOI22_X1 U15627 ( .A1(n13353), .A2(n13396), .B1(n13352), .B2(n13385), .ZN(
        n13354) );
  OAI211_X1 U15628 ( .C1(n13356), .C2(n13428), .A(n13355), .B(n13354), .ZN(
        n13459) );
  NAND2_X1 U15629 ( .A1(n13459), .A2(n13405), .ZN(n13362) );
  OAI22_X1 U15630 ( .A1(n13358), .A2(n15681), .B1(n13405), .B2(n13357), .ZN(
        n13359) );
  AOI21_X1 U15631 ( .B1(n13360), .B2(n13438), .A(n13359), .ZN(n13361) );
  OAI211_X1 U15632 ( .C1(n13364), .C2(n13363), .A(n13362), .B(n13361), .ZN(
        P3_U3209) );
  XNOR2_X1 U15633 ( .A(n13365), .B(n13367), .ZN(n13372) );
  XNOR2_X1 U15634 ( .A(n13366), .B(n13367), .ZN(n13464) );
  NAND2_X1 U15635 ( .A1(n13464), .A2(n13368), .ZN(n13371) );
  AOI22_X1 U15636 ( .A1(n13369), .A2(n13396), .B1(n13352), .B2(n13397), .ZN(
        n13370) );
  OAI211_X1 U15637 ( .C1(n13372), .C2(n13428), .A(n13371), .B(n13370), .ZN(
        n13463) );
  INV_X1 U15638 ( .A(n13463), .ZN(n13379) );
  INV_X1 U15639 ( .A(n13373), .ZN(n13517) );
  AOI22_X1 U15640 ( .A1(n13374), .A2(n15675), .B1(n15688), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13375) );
  OAI21_X1 U15641 ( .B1(n13517), .B2(n13403), .A(n13375), .ZN(n13376) );
  AOI21_X1 U15642 ( .B1(n13464), .B2(n13377), .A(n13376), .ZN(n13378) );
  OAI21_X1 U15643 ( .B1(n13379), .B2(n15688), .A(n13378), .ZN(P3_U3210) );
  XNOR2_X1 U15644 ( .A(n13380), .B(n13381), .ZN(n13524) );
  XNOR2_X1 U15645 ( .A(n13383), .B(n13382), .ZN(n13386) );
  AOI222_X1 U15646 ( .A1(n13386), .A2(n13398), .B1(n13385), .B2(n13396), .C1(
        n13384), .C2(n13352), .ZN(n13518) );
  MUX2_X1 U15647 ( .A(n13387), .B(n13518), .S(n13405), .Z(n13390) );
  AOI22_X1 U15648 ( .A1(n13521), .A2(n13438), .B1(n15675), .B2(n13388), .ZN(
        n13389) );
  OAI211_X1 U15649 ( .C1(n13524), .C2(n13441), .A(n13390), .B(n13389), .ZN(
        P3_U3211) );
  XNOR2_X1 U15650 ( .A(n13393), .B(n13391), .ZN(n13473) );
  INV_X1 U15651 ( .A(n13473), .ZN(n13407) );
  OAI21_X1 U15652 ( .B1(n13394), .B2(n13393), .A(n13392), .ZN(n13399) );
  AOI222_X1 U15653 ( .A1(n13399), .A2(n13398), .B1(n13397), .B2(n13396), .C1(
        n13395), .C2(n13352), .ZN(n13400) );
  INV_X1 U15654 ( .A(n13400), .ZN(n13472) );
  AOI22_X1 U15655 ( .A1(n13401), .A2(n15675), .B1(n15688), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n13402) );
  OAI21_X1 U15656 ( .B1(n13528), .B2(n13403), .A(n13402), .ZN(n13404) );
  AOI21_X1 U15657 ( .B1(n13472), .B2(n13405), .A(n13404), .ZN(n13406) );
  OAI21_X1 U15658 ( .B1(n13407), .B2(n13441), .A(n13406), .ZN(P3_U3212) );
  XOR2_X1 U15659 ( .A(n13411), .B(n13408), .Z(n13530) );
  INV_X1 U15660 ( .A(n13530), .ZN(n13421) );
  INV_X1 U15661 ( .A(n13535), .ZN(n13410) );
  AOI22_X1 U15662 ( .A1(n13410), .A2(n13438), .B1(n15675), .B2(n13409), .ZN(
        n13420) );
  AOI21_X1 U15663 ( .B1(n13412), .B2(n13411), .A(n13428), .ZN(n13417) );
  OAI22_X1 U15664 ( .A1(n13414), .A2(n13433), .B1(n13413), .B2(n13431), .ZN(
        n13415) );
  AOI21_X1 U15665 ( .B1(n13417), .B2(n13416), .A(n13415), .ZN(n13532) );
  MUX2_X1 U15666 ( .A(n13532), .B(n13418), .S(n15688), .Z(n13419) );
  OAI211_X1 U15667 ( .C1(n13421), .C2(n13441), .A(n13420), .B(n13419), .ZN(
        P3_U3214) );
  OAI21_X1 U15668 ( .B1(n13423), .B2(n13427), .A(n13422), .ZN(n13541) );
  INV_X1 U15669 ( .A(n13424), .ZN(n13425) );
  AOI21_X1 U15670 ( .B1(n13427), .B2(n13426), .A(n13425), .ZN(n13429) );
  OAI222_X1 U15671 ( .A1(n13433), .A2(n13432), .B1(n13431), .B2(n13430), .C1(
        n13429), .C2(n13428), .ZN(n13483) );
  NAND2_X1 U15672 ( .A1(n13483), .A2(n13405), .ZN(n13440) );
  INV_X1 U15673 ( .A(n13434), .ZN(n13435) );
  OAI22_X1 U15674 ( .A1(n13405), .A2(n13436), .B1(n13435), .B2(n15681), .ZN(
        n13437) );
  AOI21_X1 U15675 ( .B1(n13484), .B2(n13438), .A(n13437), .ZN(n13439) );
  OAI211_X1 U15676 ( .C1(n13541), .C2(n13441), .A(n13440), .B(n13439), .ZN(
        P3_U3215) );
  NAND2_X1 U15677 ( .A1(n13489), .A2(n13486), .ZN(n13444) );
  NAND2_X1 U15678 ( .A1(n13478), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13442) );
  OAI211_X1 U15679 ( .C1(n13491), .C2(n13482), .A(n13444), .B(n13442), .ZN(
        P3_U3490) );
  NAND2_X1 U15680 ( .A1(n13478), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13443) );
  OAI211_X1 U15681 ( .C1(n13494), .C2(n13482), .A(n13444), .B(n13443), .ZN(
        P3_U3489) );
  INV_X1 U15682 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13448) );
  AND2_X1 U15683 ( .A1(n13445), .A2(n13474), .ZN(n13446) );
  NOR2_X1 U15684 ( .A1(n13447), .A2(n13446), .ZN(n13495) );
  MUX2_X1 U15685 ( .A(n15829), .B(n13498), .S(n13486), .Z(n13451) );
  INV_X1 U15686 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13454) );
  AOI21_X1 U15687 ( .B1(n13465), .B2(n13453), .A(n13452), .ZN(n13502) );
  MUX2_X1 U15688 ( .A(n13454), .B(n13502), .S(n13486), .Z(n13455) );
  OAI21_X1 U15689 ( .B1(n13504), .B2(n13482), .A(n13455), .ZN(P3_U3485) );
  INV_X1 U15690 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13456) );
  MUX2_X1 U15691 ( .A(n13456), .B(n13506), .S(n13486), .Z(n13458) );
  NAND2_X1 U15692 ( .A1(n13507), .A2(n13469), .ZN(n13457) );
  OAI211_X1 U15693 ( .C1(n13510), .C2(n13488), .A(n13458), .B(n13457), .ZN(
        P3_U3484) );
  INV_X1 U15694 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13461) );
  AOI21_X1 U15695 ( .B1(n13465), .B2(n13460), .A(n13459), .ZN(n13511) );
  MUX2_X1 U15696 ( .A(n13461), .B(n13511), .S(n13486), .Z(n13462) );
  OAI21_X1 U15697 ( .B1(n7237), .B2(n13482), .A(n13462), .ZN(P3_U3483) );
  INV_X1 U15698 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13466) );
  AOI21_X1 U15699 ( .B1(n13465), .B2(n13464), .A(n13463), .ZN(n13514) );
  MUX2_X1 U15700 ( .A(n13466), .B(n13514), .S(n13486), .Z(n13467) );
  OAI21_X1 U15701 ( .B1(n13517), .B2(n13482), .A(n13467), .ZN(P3_U3482) );
  INV_X1 U15702 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13468) );
  MUX2_X1 U15703 ( .A(n13468), .B(n13518), .S(n13486), .Z(n13471) );
  NAND2_X1 U15704 ( .A1(n13521), .A2(n13469), .ZN(n13470) );
  OAI211_X1 U15705 ( .C1(n13524), .C2(n13488), .A(n13471), .B(n13470), .ZN(
        P3_U3481) );
  INV_X1 U15706 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13475) );
  AOI21_X1 U15707 ( .B1(n13474), .B2(n13473), .A(n13472), .ZN(n13525) );
  MUX2_X1 U15708 ( .A(n13475), .B(n13525), .S(n13486), .Z(n13476) );
  OAI21_X1 U15709 ( .B1(n13528), .B2(n13482), .A(n13476), .ZN(P3_U3480) );
  NAND2_X1 U15710 ( .A1(n13530), .A2(n13477), .ZN(n13481) );
  INV_X1 U15711 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13479) );
  MUX2_X1 U15712 ( .A(n13532), .B(n13479), .S(n13478), .Z(n13480) );
  OAI211_X1 U15713 ( .C1(n13482), .C2(n13535), .A(n13481), .B(n13480), .ZN(
        P3_U3478) );
  AOI21_X1 U15714 ( .B1(n13485), .B2(n13484), .A(n13483), .ZN(n13537) );
  MUX2_X1 U15715 ( .A(n15759), .B(n13537), .S(n13486), .Z(n13487) );
  OAI21_X1 U15716 ( .B1(n13488), .B2(n13541), .A(n13487), .ZN(P3_U3477) );
  NAND2_X1 U15717 ( .A1(n13489), .A2(n15691), .ZN(n13493) );
  NAND2_X1 U15718 ( .A1(n15693), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13490) );
  OAI211_X1 U15719 ( .C1(n13491), .C2(n13536), .A(n13493), .B(n13490), .ZN(
        P3_U3458) );
  NAND2_X1 U15720 ( .A1(n15693), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13492) );
  OAI211_X1 U15721 ( .C1(n13494), .C2(n13536), .A(n13493), .B(n13492), .ZN(
        P3_U3457) );
  INV_X1 U15722 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13496) );
  INV_X1 U15723 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13499) );
  MUX2_X1 U15724 ( .A(n13499), .B(n13498), .S(n15691), .Z(n13500) );
  INV_X1 U15725 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n15731) );
  MUX2_X1 U15726 ( .A(n15731), .B(n13502), .S(n15691), .Z(n13503) );
  OAI21_X1 U15727 ( .B1(n13504), .B2(n13536), .A(n13503), .ZN(P3_U3453) );
  INV_X1 U15728 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13505) );
  MUX2_X1 U15729 ( .A(n13506), .B(n13505), .S(n15693), .Z(n13509) );
  NAND2_X1 U15730 ( .A1(n13507), .A2(n13520), .ZN(n13508) );
  OAI211_X1 U15731 ( .C1(n13510), .C2(n13540), .A(n13509), .B(n13508), .ZN(
        P3_U3452) );
  INV_X1 U15732 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13512) );
  MUX2_X1 U15733 ( .A(n13512), .B(n13511), .S(n15691), .Z(n13513) );
  OAI21_X1 U15734 ( .B1(n7237), .B2(n13536), .A(n13513), .ZN(P3_U3451) );
  INV_X1 U15735 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13515) );
  MUX2_X1 U15736 ( .A(n13515), .B(n13514), .S(n15691), .Z(n13516) );
  OAI21_X1 U15737 ( .B1(n13517), .B2(n13536), .A(n13516), .ZN(P3_U3450) );
  INV_X1 U15738 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13519) );
  MUX2_X1 U15739 ( .A(n13519), .B(n13518), .S(n15691), .Z(n13523) );
  NAND2_X1 U15740 ( .A1(n13521), .A2(n13520), .ZN(n13522) );
  OAI211_X1 U15741 ( .C1(n13524), .C2(n13540), .A(n13523), .B(n13522), .ZN(
        P3_U3449) );
  INV_X1 U15742 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13526) );
  MUX2_X1 U15743 ( .A(n13526), .B(n13525), .S(n15691), .Z(n13527) );
  OAI21_X1 U15744 ( .B1(n13528), .B2(n13536), .A(n13527), .ZN(P3_U3448) );
  NAND2_X1 U15745 ( .A1(n13530), .A2(n13529), .ZN(n13534) );
  INV_X1 U15746 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13531) );
  MUX2_X1 U15747 ( .A(n13532), .B(n13531), .S(n15693), .Z(n13533) );
  OAI211_X1 U15748 ( .C1(n13536), .C2(n13535), .A(n13534), .B(n13533), .ZN(
        P3_U3446) );
  INV_X1 U15749 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13538) );
  MUX2_X1 U15750 ( .A(n13538), .B(n13537), .S(n15691), .Z(n13539) );
  OAI21_X1 U15751 ( .B1(n13541), .B2(n13540), .A(n13539), .ZN(P3_U3444) );
  INV_X1 U15752 ( .A(SI_30_), .ZN(n13544) );
  INV_X1 U15753 ( .A(n13542), .ZN(n13543) );
  OAI222_X1 U15754 ( .A1(n13545), .A2(P3_U3151), .B1(n13550), .B2(n13544), 
        .C1(n12962), .C2(n13543), .ZN(P3_U3265) );
  INV_X1 U15755 ( .A(n13546), .ZN(n13547) );
  OAI222_X1 U15756 ( .A1(P3_U3151), .A2(n13548), .B1(n13550), .B2(n15944), 
        .C1(n12962), .C2(n13547), .ZN(P3_U3267) );
  INV_X1 U15757 ( .A(n13549), .ZN(n13552) );
  OAI222_X1 U15758 ( .A1(n7916), .A2(P3_U3151), .B1(n12962), .B2(n13552), .C1(
        n13551), .C2(n13550), .ZN(P3_U3268) );
  INV_X1 U15759 ( .A(n13553), .ZN(n13554) );
  OAI222_X1 U15760 ( .A1(P3_U3151), .A2(n13555), .B1(n13550), .B2(n15772), 
        .C1(n12962), .C2(n13554), .ZN(P3_U3269) );
  INV_X1 U15761 ( .A(n13556), .ZN(n13557) );
  OAI222_X1 U15762 ( .A1(P3_U3151), .A2(n13559), .B1(n13550), .B2(n13558), 
        .C1(n12962), .C2(n13557), .ZN(P3_U3270) );
  OAI211_X1 U15763 ( .C1(n13562), .C2(n13561), .A(n13560), .B(n13711), .ZN(
        n13567) );
  NOR2_X1 U15764 ( .A1(n14072), .A2(n13717), .ZN(n13565) );
  OAI22_X1 U15765 ( .A1(n14064), .A2(n13587), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13563), .ZN(n13564) );
  AOI211_X1 U15766 ( .C1(n13962), .C2(n13675), .A(n13565), .B(n13564), .ZN(
        n13566) );
  OAI211_X1 U15767 ( .C1(n14413), .C2(n13725), .A(n13567), .B(n13566), .ZN(
        P2_U3186) );
  OAI21_X1 U15768 ( .B1(n13570), .B2(n13569), .A(n13568), .ZN(n13571) );
  NAND2_X1 U15769 ( .A1(n13571), .A2(n13711), .ZN(n13578) );
  INV_X1 U15770 ( .A(n13572), .ZN(n13576) );
  INV_X1 U15771 ( .A(n14273), .ZN(n13573) );
  OAI22_X1 U15772 ( .A1(n13574), .A2(n13587), .B1(n13717), .B2(n13573), .ZN(
        n13575) );
  AOI211_X1 U15773 ( .C1(n13675), .C2(n14268), .A(n13576), .B(n13575), .ZN(
        n13577) );
  OAI211_X1 U15774 ( .C1(n14276), .C2(n13725), .A(n13578), .B(n13577), .ZN(
        P2_U3187) );
  NAND2_X1 U15775 ( .A1(n13661), .A2(n13579), .ZN(n13662) );
  INV_X1 U15776 ( .A(n13580), .ZN(n13581) );
  NAND2_X1 U15777 ( .A1(n13662), .A2(n13581), .ZN(n13583) );
  XNOR2_X1 U15778 ( .A(n13583), .B(n13582), .ZN(n13586) );
  OAI22_X1 U15779 ( .A1(n13586), .A2(n13695), .B1(n13665), .B2(n13697), .ZN(
        n13584) );
  OAI21_X1 U15780 ( .B1(n13586), .B2(n13585), .A(n13584), .ZN(n13591) );
  OAI22_X1 U15781 ( .A1(n14117), .A2(n13587), .B1(n13717), .B2(n14123), .ZN(
        n13589) );
  NOR2_X1 U15782 ( .A1(n14119), .A2(n13718), .ZN(n13588) );
  AOI211_X1 U15783 ( .C1(P2_REG3_REG_23__SCAN_IN), .C2(P2_U3088), .A(n13589), 
        .B(n13588), .ZN(n13590) );
  OAI211_X1 U15784 ( .C1(n14423), .C2(n13725), .A(n13591), .B(n13590), .ZN(
        P2_U3188) );
  INV_X1 U15785 ( .A(n13592), .ZN(n13611) );
  NOR2_X1 U15786 ( .A1(n13611), .A2(n13593), .ZN(n13594) );
  XNOR2_X1 U15787 ( .A(n13613), .B(n13594), .ZN(n13599) );
  AOI22_X1 U15788 ( .A1(n13969), .A2(n14304), .B1(n14302), .B2(n13971), .ZN(
        n14357) );
  INV_X1 U15789 ( .A(n14357), .ZN(n14190) );
  NOR2_X1 U15790 ( .A1(n13595), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14020) );
  AOI21_X1 U15791 ( .B1(n14190), .B2(n13666), .A(n14020), .ZN(n13596) );
  OAI21_X1 U15792 ( .B1(n14191), .B2(n13717), .A(n13596), .ZN(n13597) );
  AOI21_X1 U15793 ( .B1(n14196), .B2(n13693), .A(n13597), .ZN(n13598) );
  OAI21_X1 U15794 ( .B1(n13599), .B2(n13695), .A(n13598), .ZN(P2_U3191) );
  AOI22_X1 U15795 ( .A1(n13745), .A2(n13693), .B1(n13675), .B2(n13980), .ZN(
        n13610) );
  AOI22_X1 U15796 ( .A1(n13722), .A2(n10541), .B1(n13676), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n13609) );
  XNOR2_X1 U15797 ( .A(n13679), .B(n13678), .ZN(n13604) );
  INV_X1 U15798 ( .A(n13600), .ZN(n13601) );
  NAND2_X1 U15799 ( .A1(n13601), .A2(n13604), .ZN(n13677) );
  OAI21_X1 U15800 ( .B1(n13604), .B2(n13602), .A(n13677), .ZN(n13603) );
  NAND2_X1 U15801 ( .A1(n13603), .A2(n13711), .ZN(n13608) );
  INV_X1 U15802 ( .A(n13604), .ZN(n13605) );
  NAND3_X1 U15803 ( .A1(n13712), .A2(n13606), .A3(n13605), .ZN(n13607) );
  NAND4_X1 U15804 ( .A1(n13610), .A2(n13609), .A3(n13608), .A4(n13607), .ZN(
        P2_U3194) );
  INV_X1 U15805 ( .A(n13613), .ZN(n13651) );
  AOI21_X1 U15806 ( .B1(n13613), .B2(n13612), .A(n13611), .ZN(n13650) );
  XNOR2_X1 U15807 ( .A(n13615), .B(n13614), .ZN(n13659) );
  OAI211_X1 U15808 ( .C1(n13651), .C2(n13616), .A(n13650), .B(n13659), .ZN(
        n13655) );
  AOI21_X1 U15809 ( .B1(n13655), .B2(n13618), .A(n13617), .ZN(n13625) );
  NAND2_X1 U15810 ( .A1(n13619), .A2(n13711), .ZN(n13624) );
  OAI22_X1 U15811 ( .A1(n14117), .A2(n14118), .B1(n13620), .B2(n14116), .ZN(
        n14156) );
  AOI22_X1 U15812 ( .A1(n14156), .A2(n13666), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13621) );
  OAI21_X1 U15813 ( .B1(n14158), .B2(n13717), .A(n13621), .ZN(n13622) );
  AOI21_X1 U15814 ( .B1(n14345), .B2(n13693), .A(n13622), .ZN(n13623) );
  OAI21_X1 U15815 ( .B1(n13625), .B2(n13624), .A(n13623), .ZN(P2_U3195) );
  XNOR2_X1 U15816 ( .A(n13626), .B(n13627), .ZN(n13713) );
  OAI22_X1 U15817 ( .A1(n13713), .A2(n13710), .B1(n13627), .B2(n13626), .ZN(
        n13631) );
  NOR2_X1 U15818 ( .A1(n13629), .A2(n13628), .ZN(n13630) );
  XNOR2_X1 U15819 ( .A(n13631), .B(n13630), .ZN(n13636) );
  AOI22_X1 U15820 ( .A1(n13722), .A2(n14268), .B1(n13701), .B2(n14235), .ZN(
        n13632) );
  NAND2_X1 U15821 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n15590)
         );
  OAI211_X1 U15822 ( .C1(n13633), .C2(n13718), .A(n13632), .B(n15590), .ZN(
        n13634) );
  AOI21_X1 U15823 ( .B1(n14372), .B2(n13693), .A(n13634), .ZN(n13635) );
  OAI21_X1 U15824 ( .B1(n13636), .B2(n13695), .A(n13635), .ZN(P2_U3198) );
  OAI21_X1 U15825 ( .B1(n13639), .B2(n13637), .A(n13638), .ZN(n13640) );
  NAND2_X1 U15826 ( .A1(n13640), .A2(n13711), .ZN(n13643) );
  AOI22_X1 U15827 ( .A1(n13971), .A2(n14304), .B1(n14302), .B2(n14253), .ZN(
        n14216) );
  NAND2_X1 U15828 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15607)
         );
  OAI21_X1 U15829 ( .B1(n13703), .B2(n14216), .A(n15607), .ZN(n13641) );
  AOI21_X1 U15830 ( .B1(n13701), .B2(n14220), .A(n13641), .ZN(n13642) );
  OAI211_X1 U15831 ( .C1(n14222), .C2(n13725), .A(n13643), .B(n13642), .ZN(
        P2_U3200) );
  OAI211_X1 U15832 ( .C1(n13645), .C2(n13644), .A(n12893), .B(n13711), .ZN(
        n13649) );
  OAI22_X1 U15833 ( .A1(n13698), .A2(n14118), .B1(n13665), .B2(n14116), .ZN(
        n14101) );
  OAI22_X1 U15834 ( .A1(n14107), .A2(n13717), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13646), .ZN(n13647) );
  AOI21_X1 U15835 ( .B1(n14101), .B2(n13666), .A(n13647), .ZN(n13648) );
  OAI211_X1 U15836 ( .C1(n14418), .C2(n13725), .A(n13649), .B(n13648), .ZN(
        P2_U3201) );
  INV_X1 U15837 ( .A(n13650), .ZN(n13653) );
  NOR3_X1 U15838 ( .A1(n13651), .A2(n14153), .A3(n13697), .ZN(n13652) );
  AOI21_X1 U15839 ( .B1(n13711), .B2(n13653), .A(n13652), .ZN(n13660) );
  OAI22_X1 U15840 ( .A1(n13664), .A2(n14118), .B1(n14153), .B2(n14116), .ZN(
        n14170) );
  AOI22_X1 U15841 ( .A1(n14170), .A2(n13666), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13654) );
  OAI21_X1 U15842 ( .B1(n14176), .B2(n13717), .A(n13654), .ZN(n13657) );
  NOR2_X1 U15843 ( .A1(n13655), .A2(n13695), .ZN(n13656) );
  AOI211_X1 U15844 ( .C1(n14353), .C2(n13693), .A(n13657), .B(n13656), .ZN(
        n13658) );
  OAI21_X1 U15845 ( .B1(n13660), .B2(n13659), .A(n13658), .ZN(P2_U3205) );
  AOI22_X1 U15846 ( .A1(n13661), .A2(n13711), .B1(n13712), .B2(n13967), .ZN(
        n13671) );
  INV_X1 U15847 ( .A(n13662), .ZN(n13670) );
  INV_X1 U15848 ( .A(n13663), .ZN(n14143) );
  OAI22_X1 U15849 ( .A1(n13665), .A2(n14118), .B1(n13664), .B2(n14116), .ZN(
        n14136) );
  AOI22_X1 U15850 ( .A1(n14136), .A2(n13666), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13667) );
  OAI21_X1 U15851 ( .B1(n14143), .B2(n13717), .A(n13667), .ZN(n13668) );
  AOI21_X1 U15852 ( .B1(n14145), .B2(n13693), .A(n13668), .ZN(n13669) );
  OAI21_X1 U15853 ( .B1(n13671), .B2(n13670), .A(n13669), .ZN(P2_U3207) );
  OAI22_X1 U15854 ( .A1(n13697), .A2(n13744), .B1(n13678), .B2(n13695), .ZN(
        n13674) );
  XNOR2_X1 U15855 ( .A(n13672), .B(n13673), .ZN(n13681) );
  NAND3_X1 U15856 ( .A1(n13674), .A2(n13681), .A3(n13677), .ZN(n13688) );
  AOI22_X1 U15857 ( .A1(n13741), .A2(n13693), .B1(n13675), .B2(n13979), .ZN(
        n13687) );
  AOI22_X1 U15858 ( .A1(n13722), .A2(n13981), .B1(n13676), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n13686) );
  INV_X1 U15859 ( .A(n13677), .ZN(n13684) );
  INV_X1 U15860 ( .A(n13678), .ZN(n13680) );
  NOR2_X1 U15861 ( .A1(n13680), .A2(n13679), .ZN(n13683) );
  INV_X1 U15862 ( .A(n13681), .ZN(n13682) );
  OAI211_X1 U15863 ( .C1(n13684), .C2(n13683), .A(n13711), .B(n13682), .ZN(
        n13685) );
  NAND4_X1 U15864 ( .A1(n13688), .A2(n13687), .A3(n13686), .A4(n13685), .ZN(
        P2_U3209) );
  XNOR2_X1 U15865 ( .A(n13690), .B(n13689), .ZN(n13696) );
  NOR2_X1 U15866 ( .A1(n13717), .A2(n14206), .ZN(n13692) );
  AOI22_X1 U15867 ( .A1(n13970), .A2(n14304), .B1(n14302), .B2(n14231), .ZN(
        n14202) );
  NAND2_X1 U15868 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14003)
         );
  OAI21_X1 U15869 ( .B1(n14202), .B2(n13703), .A(n14003), .ZN(n13691) );
  AOI211_X1 U15870 ( .C1(n14365), .C2(n13693), .A(n13692), .B(n13691), .ZN(
        n13694) );
  OAI21_X1 U15871 ( .B1(n13696), .B2(n13695), .A(n13694), .ZN(P2_U3210) );
  NOR3_X1 U15872 ( .A1(n13699), .A2(n13698), .A3(n13697), .ZN(n13700) );
  AOI21_X1 U15873 ( .B1(n12898), .B2(n13711), .A(n13700), .ZN(n13709) );
  NOR2_X1 U15874 ( .A1(n14082), .A2(n13725), .ZN(n13706) );
  AOI22_X1 U15875 ( .A1(n14080), .A2(n13701), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13702) );
  OAI21_X1 U15876 ( .B1(n13704), .B2(n13703), .A(n13702), .ZN(n13705) );
  OAI21_X1 U15877 ( .B1(n13709), .B2(n6705), .A(n13708), .ZN(P2_U3212) );
  NAND2_X1 U15878 ( .A1(n13711), .A2(n13710), .ZN(n13715) );
  NAND2_X1 U15879 ( .A1(n13712), .A2(n14268), .ZN(n13714) );
  MUX2_X1 U15880 ( .A(n13715), .B(n13714), .S(n13713), .Z(n13724) );
  INV_X1 U15881 ( .A(n14260), .ZN(n13716) );
  OAI22_X1 U15882 ( .A1(n13719), .A2(n13718), .B1(n13717), .B2(n13716), .ZN(
        n13720) );
  AOI211_X1 U15883 ( .C1(n13722), .C2(n14254), .A(n13721), .B(n13720), .ZN(
        n13723) );
  OAI211_X1 U15884 ( .C1(n7850), .C2(n13725), .A(n13724), .B(n13723), .ZN(
        P2_U3213) );
  MUX2_X1 U15885 ( .A(n14082), .B(n14064), .S(n13867), .Z(n13864) );
  INV_X1 U15886 ( .A(n13864), .ZN(n13880) );
  OAI21_X1 U15887 ( .B1(n13977), .B2(n13768), .A(n13726), .ZN(n13730) );
  NAND2_X1 U15888 ( .A1(n13977), .A2(n13768), .ZN(n13728) );
  NAND2_X1 U15889 ( .A1(n13728), .A2(n13727), .ZN(n13729) );
  NAND2_X1 U15890 ( .A1(n13730), .A2(n13729), .ZN(n13731) );
  OAI21_X1 U15891 ( .B1(n13978), .B2(n13743), .A(n15632), .ZN(n13736) );
  NAND2_X1 U15892 ( .A1(n13978), .A2(n13855), .ZN(n13734) );
  NAND2_X1 U15893 ( .A1(n13734), .A2(n13733), .ZN(n13735) );
  NAND2_X1 U15894 ( .A1(n13736), .A2(n13735), .ZN(n13737) );
  NAND2_X1 U15895 ( .A1(n13907), .A2(n13737), .ZN(n13739) );
  AOI21_X1 U15896 ( .B1(n13774), .B2(n13739), .A(n13738), .ZN(n13782) );
  OAI21_X1 U15897 ( .B1(n13980), .B2(n13743), .A(n13741), .ZN(n13740) );
  INV_X1 U15898 ( .A(n13740), .ZN(n13766) );
  AOI21_X1 U15899 ( .B1(n13980), .B2(n13855), .A(n13741), .ZN(n13765) );
  AOI21_X1 U15900 ( .B1(n13744), .B2(n13743), .A(n13742), .ZN(n13763) );
  AOI21_X1 U15901 ( .B1(n13981), .B2(n13768), .A(n13745), .ZN(n13762) );
  NAND2_X1 U15902 ( .A1(n13944), .A2(n14017), .ZN(n13746) );
  AND2_X1 U15903 ( .A1(n13747), .A2(n13746), .ZN(n13751) );
  NAND3_X1 U15904 ( .A1(n13749), .A2(n13748), .A3(n13751), .ZN(n13754) );
  INV_X1 U15905 ( .A(n13750), .ZN(n13753) );
  INV_X1 U15906 ( .A(n13751), .ZN(n13752) );
  OAI22_X1 U15907 ( .A1(n13754), .A2(n13753), .B1(n13752), .B2(n13757), .ZN(
        n13755) );
  INV_X1 U15908 ( .A(n13755), .ZN(n13760) );
  NAND3_X1 U15909 ( .A1(n11232), .A2(n13756), .A3(n13768), .ZN(n13759) );
  NAND3_X1 U15910 ( .A1(n10541), .A2(n13743), .A3(n13757), .ZN(n13758) );
  NAND4_X1 U15911 ( .A1(n13904), .A2(n13760), .A3(n13759), .A4(n13758), .ZN(
        n13761) );
  OAI211_X1 U15912 ( .C1(n13763), .C2(n13762), .A(n13761), .B(n13903), .ZN(
        n13764) );
  OAI211_X1 U15913 ( .C1(n13766), .C2(n13765), .A(n13764), .B(n13910), .ZN(
        n13775) );
  OAI21_X1 U15914 ( .B1(n13979), .B2(n13768), .A(n13767), .ZN(n13772) );
  NAND2_X1 U15915 ( .A1(n13979), .A2(n13768), .ZN(n13770) );
  NAND2_X1 U15916 ( .A1(n13770), .A2(n13769), .ZN(n13771) );
  NAND2_X1 U15917 ( .A1(n13772), .A2(n13771), .ZN(n13773) );
  NAND4_X1 U15918 ( .A1(n13775), .A2(n13774), .A3(n13908), .A4(n13773), .ZN(
        n13781) );
  AOI21_X1 U15919 ( .B1(n13776), .B2(n13867), .A(n15641), .ZN(n13779) );
  AOI21_X1 U15920 ( .B1(n13976), .B2(n13855), .A(n13777), .ZN(n13778) );
  OR2_X1 U15921 ( .A1(n13779), .A2(n13778), .ZN(n13780) );
  NAND3_X1 U15922 ( .A1(n13782), .A2(n13781), .A3(n13780), .ZN(n13787) );
  AND2_X1 U15923 ( .A1(n13975), .A2(n13867), .ZN(n13784) );
  OAI21_X1 U15924 ( .B1(n13975), .B2(n13867), .A(n15650), .ZN(n13783) );
  OAI21_X1 U15925 ( .B1(n13784), .B2(n15650), .A(n13783), .ZN(n13785) );
  NAND2_X1 U15926 ( .A1(n13787), .A2(n13786), .ZN(n13792) );
  AND2_X1 U15927 ( .A1(n13974), .A2(n13855), .ZN(n13790) );
  OAI21_X1 U15928 ( .B1(n13855), .B2(n13974), .A(n13789), .ZN(n13788) );
  OAI21_X1 U15929 ( .B1(n13790), .B2(n13789), .A(n13788), .ZN(n13791) );
  NAND3_X1 U15930 ( .A1(n13792), .A2(n13791), .A3(n13902), .ZN(n13797) );
  AND2_X1 U15931 ( .A1(n13973), .A2(n13867), .ZN(n13795) );
  OAI21_X1 U15932 ( .B1(n13867), .B2(n13973), .A(n13794), .ZN(n13793) );
  OAI21_X1 U15933 ( .B1(n13795), .B2(n13794), .A(n13793), .ZN(n13796) );
  NAND3_X1 U15934 ( .A1(n13797), .A2(n13796), .A3(n13901), .ZN(n13801) );
  AND2_X1 U15935 ( .A1(n14303), .A2(n13855), .ZN(n13799) );
  OAI21_X1 U15936 ( .B1(n13855), .B2(n14303), .A(n14405), .ZN(n13798) );
  OAI21_X1 U15937 ( .B1(n13799), .B2(n14405), .A(n13798), .ZN(n13800) );
  NAND3_X1 U15938 ( .A1(n13801), .A2(n13800), .A3(n13913), .ZN(n13805) );
  AND2_X1 U15939 ( .A1(n13972), .A2(n13867), .ZN(n13803) );
  OAI21_X1 U15940 ( .B1(n13867), .B2(n13972), .A(n14399), .ZN(n13802) );
  OAI21_X1 U15941 ( .B1(n13803), .B2(n14399), .A(n13802), .ZN(n13804) );
  NAND2_X1 U15942 ( .A1(n13805), .A2(n13804), .ZN(n13807) );
  MUX2_X1 U15943 ( .A(n14305), .B(n14393), .S(n13855), .Z(n13808) );
  MUX2_X1 U15944 ( .A(n14305), .B(n14393), .S(n13867), .Z(n13806) );
  MUX2_X1 U15945 ( .A(n14269), .B(n14389), .S(n13867), .Z(n13810) );
  MUX2_X1 U15946 ( .A(n14269), .B(n14389), .S(n13855), .Z(n13809) );
  MUX2_X1 U15947 ( .A(n14254), .B(n14383), .S(n13855), .Z(n13814) );
  NAND2_X1 U15948 ( .A1(n13813), .A2(n13814), .ZN(n13812) );
  MUX2_X1 U15949 ( .A(n14254), .B(n14383), .S(n13867), .Z(n13811) );
  NAND2_X1 U15950 ( .A1(n13812), .A2(n13811), .ZN(n13818) );
  INV_X1 U15951 ( .A(n13813), .ZN(n13816) );
  INV_X1 U15952 ( .A(n13814), .ZN(n13815) );
  NAND2_X1 U15953 ( .A1(n13816), .A2(n13815), .ZN(n13817) );
  MUX2_X1 U15954 ( .A(n14268), .B(n14259), .S(n13867), .Z(n13820) );
  MUX2_X1 U15955 ( .A(n14268), .B(n14259), .S(n13855), .Z(n13819) );
  INV_X1 U15956 ( .A(n13820), .ZN(n13821) );
  MUX2_X1 U15957 ( .A(n14253), .B(n14372), .S(n13855), .Z(n13823) );
  MUX2_X1 U15958 ( .A(n14253), .B(n14372), .S(n13867), .Z(n13822) );
  MUX2_X1 U15959 ( .A(n14231), .B(n14368), .S(n13867), .Z(n13824) );
  NAND2_X1 U15960 ( .A1(n13827), .A2(n13824), .ZN(n13826) );
  MUX2_X1 U15961 ( .A(n14231), .B(n14368), .S(n13855), .Z(n13825) );
  NAND2_X1 U15962 ( .A1(n13826), .A2(n13825), .ZN(n13830) );
  INV_X1 U15963 ( .A(n13827), .ZN(n13828) );
  NAND2_X1 U15964 ( .A1(n13828), .A2(n6633), .ZN(n13829) );
  MUX2_X1 U15965 ( .A(n13971), .B(n14365), .S(n13855), .Z(n13832) );
  MUX2_X1 U15966 ( .A(n13971), .B(n14365), .S(n13867), .Z(n13831) );
  MUX2_X1 U15967 ( .A(n13970), .B(n14196), .S(n13867), .Z(n13836) );
  NAND2_X1 U15968 ( .A1(n13835), .A2(n13836), .ZN(n13834) );
  MUX2_X1 U15969 ( .A(n13970), .B(n14196), .S(n13855), .Z(n13833) );
  NAND2_X1 U15970 ( .A1(n13834), .A2(n13833), .ZN(n13840) );
  INV_X1 U15971 ( .A(n13835), .ZN(n13838) );
  INV_X1 U15972 ( .A(n13836), .ZN(n13837) );
  NAND2_X1 U15973 ( .A1(n13838), .A2(n13837), .ZN(n13839) );
  MUX2_X1 U15974 ( .A(n13969), .B(n14353), .S(n13855), .Z(n13842) );
  MUX2_X1 U15975 ( .A(n13969), .B(n14353), .S(n13867), .Z(n13841) );
  MUX2_X1 U15976 ( .A(n13968), .B(n14345), .S(n13867), .Z(n13844) );
  MUX2_X1 U15977 ( .A(n13968), .B(n14345), .S(n13855), .Z(n13843) );
  MUX2_X1 U15978 ( .A(n13967), .B(n14145), .S(n13855), .Z(n13848) );
  NAND2_X1 U15979 ( .A1(n13847), .A2(n13848), .ZN(n13846) );
  MUX2_X1 U15980 ( .A(n13967), .B(n14145), .S(n13867), .Z(n13845) );
  NAND2_X1 U15981 ( .A1(n13846), .A2(n13845), .ZN(n13852) );
  INV_X1 U15982 ( .A(n13847), .ZN(n13850) );
  INV_X1 U15983 ( .A(n13848), .ZN(n13849) );
  NAND2_X1 U15984 ( .A1(n13850), .A2(n13849), .ZN(n13851) );
  MUX2_X1 U15985 ( .A(n13966), .B(n14129), .S(n13867), .Z(n13854) );
  MUX2_X1 U15986 ( .A(n13966), .B(n14129), .S(n13855), .Z(n13853) );
  MUX2_X1 U15987 ( .A(n13965), .B(n14109), .S(n13855), .Z(n13857) );
  MUX2_X1 U15988 ( .A(n13965), .B(n14109), .S(n13867), .Z(n13856) );
  INV_X1 U15989 ( .A(n13857), .ZN(n13858) );
  MUX2_X1 U15990 ( .A(n13964), .B(n13859), .S(n13867), .Z(n13860) );
  MUX2_X1 U15991 ( .A(n13859), .B(n13964), .S(n13867), .Z(n13861) );
  INV_X1 U15992 ( .A(n13865), .ZN(n13879) );
  MUX2_X1 U15993 ( .A(n13963), .B(n13862), .S(n13867), .Z(n13863) );
  MUX2_X1 U15994 ( .A(n13866), .B(n14413), .S(n13855), .Z(n13882) );
  MUX2_X1 U15995 ( .A(n14046), .B(n14077), .S(n13867), .Z(n13881) );
  MUX2_X1 U15996 ( .A(n13960), .B(n14031), .S(n13867), .Z(n13889) );
  INV_X1 U15997 ( .A(n8541), .ZN(n13942) );
  OAI211_X1 U15998 ( .C1(n13942), .C2(n13944), .A(n13952), .B(n13941), .ZN(
        n13868) );
  INV_X1 U15999 ( .A(n13868), .ZN(n13870) );
  NAND2_X1 U16000 ( .A1(n13959), .A2(n13867), .ZN(n13892) );
  AOI21_X1 U16001 ( .B1(n13870), .B2(n13892), .A(n13869), .ZN(n13871) );
  AOI21_X1 U16002 ( .B1(n14031), .B2(n13855), .A(n13871), .ZN(n13888) );
  NAND2_X1 U16003 ( .A1(n13889), .A2(n13888), .ZN(n13890) );
  INV_X1 U16004 ( .A(n13890), .ZN(n13877) );
  NAND2_X1 U16005 ( .A1(n13872), .A2(n13959), .ZN(n13873) );
  NAND2_X1 U16006 ( .A1(n13893), .A2(n13873), .ZN(n13898) );
  MUX2_X1 U16007 ( .A(n13874), .B(n14047), .S(n13867), .Z(n13887) );
  INV_X1 U16008 ( .A(n14047), .ZN(n13961) );
  MUX2_X1 U16009 ( .A(n14065), .B(n14040), .S(n13855), .Z(n13884) );
  AOI22_X1 U16010 ( .A1(n13887), .A2(n13886), .B1(n13884), .B2(n13883), .ZN(
        n13876) );
  OAI22_X1 U16011 ( .A1(n13884), .A2(n13883), .B1(n13882), .B2(n13881), .ZN(
        n13885) );
  OAI22_X1 U16012 ( .A1(n13889), .A2(n13888), .B1(n13887), .B2(n13886), .ZN(
        n13891) );
  NAND3_X1 U16013 ( .A1(n13891), .A2(n13890), .A3(n13898), .ZN(n13895) );
  OAI211_X1 U16014 ( .C1(n14317), .C2(n13867), .A(n13893), .B(n13892), .ZN(
        n13894) );
  INV_X1 U16015 ( .A(n13949), .ZN(n13936) );
  INV_X1 U16016 ( .A(n13898), .ZN(n13933) );
  XOR2_X1 U16017 ( .A(n13960), .B(n14031), .Z(n13932) );
  XNOR2_X1 U16018 ( .A(n14196), .B(n14153), .ZN(n14186) );
  NAND2_X1 U16019 ( .A1(n13899), .A2(n14154), .ZN(n14172) );
  NOR2_X1 U16020 ( .A1(n6633), .A2(n13900), .ZN(n14214) );
  NAND2_X1 U16021 ( .A1(n13902), .A2(n13901), .ZN(n13918) );
  NAND4_X1 U16022 ( .A1(n13904), .A2(n13942), .A3(n13903), .A4(n15621), .ZN(
        n13906) );
  NOR2_X1 U16023 ( .A1(n13906), .A2(n13905), .ZN(n13912) );
  AND2_X1 U16024 ( .A1(n13908), .A2(n13907), .ZN(n13911) );
  AND4_X1 U16025 ( .A1(n13912), .A2(n13911), .A3(n13910), .A4(n13909), .ZN(
        n13916) );
  NAND4_X1 U16026 ( .A1(n13916), .A2(n13915), .A3(n13914), .A4(n13913), .ZN(
        n13917) );
  NOR4_X1 U16027 ( .A1(n14214), .A2(n13919), .A3(n13918), .A4(n13917), .ZN(
        n13922) );
  NAND2_X1 U16028 ( .A1(n13921), .A2(n13920), .ZN(n14277) );
  NAND4_X1 U16029 ( .A1(n13922), .A2(n14250), .A3(n14227), .A4(n14277), .ZN(
        n13923) );
  NOR4_X1 U16030 ( .A1(n14186), .A2(n14172), .A3(n13923), .A4(n14200), .ZN(
        n13925) );
  NAND4_X1 U16031 ( .A1(n13925), .A2(n14103), .A3(n14161), .A4(n13924), .ZN(
        n13926) );
  NOR3_X1 U16032 ( .A1(n13927), .A2(n14124), .A3(n13926), .ZN(n13929) );
  NAND4_X1 U16033 ( .A1(n14043), .A2(n13929), .A3(n13928), .A4(n14068), .ZN(
        n13930) );
  XNOR2_X1 U16034 ( .A(n13934), .B(n14017), .ZN(n13935) );
  NOR2_X1 U16035 ( .A1(n8541), .A2(n13941), .ZN(n13938) );
  OAI22_X1 U16036 ( .A1(n13938), .A2(n14017), .B1(n13937), .B2(n13954), .ZN(
        n13939) );
  INV_X1 U16037 ( .A(n13939), .ZN(n13948) );
  INV_X1 U16038 ( .A(n13940), .ZN(n13945) );
  NAND3_X1 U16039 ( .A1(n13942), .A2(n13941), .A3(n14017), .ZN(n13943) );
  OAI21_X1 U16040 ( .B1(n13945), .B2(n13944), .A(n13943), .ZN(n13946) );
  NAND2_X1 U16041 ( .A1(n13949), .A2(n13946), .ZN(n13947) );
  OAI21_X1 U16042 ( .B1(n13949), .B2(n13948), .A(n13947), .ZN(n13950) );
  NOR2_X1 U16043 ( .A1(n13951), .A2(n13950), .ZN(n13958) );
  INV_X1 U16044 ( .A(n15615), .ZN(n15617) );
  NOR4_X1 U16045 ( .A1(n15617), .A2(n14116), .A3(n13953), .A4(n13952), .ZN(
        n13956) );
  OAI21_X1 U16046 ( .B1(n13957), .B2(n13954), .A(P2_B_REG_SCAN_IN), .ZN(n13955) );
  OAI22_X1 U16047 ( .A1(n13958), .A2(n13957), .B1(n13956), .B2(n13955), .ZN(
        P2_U3328) );
  MUX2_X1 U16048 ( .A(n13959), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13982), .Z(
        P2_U3562) );
  MUX2_X1 U16049 ( .A(n13960), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13982), .Z(
        P2_U3561) );
  MUX2_X1 U16050 ( .A(n13961), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13982), .Z(
        P2_U3560) );
  MUX2_X1 U16051 ( .A(n13962), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13982), .Z(
        P2_U3559) );
  MUX2_X1 U16052 ( .A(n14046), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13982), .Z(
        P2_U3558) );
  MUX2_X1 U16053 ( .A(n13963), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13982), .Z(
        P2_U3557) );
  MUX2_X1 U16054 ( .A(n13964), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13982), .Z(
        P2_U3556) );
  MUX2_X1 U16055 ( .A(n13965), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13982), .Z(
        P2_U3555) );
  MUX2_X1 U16056 ( .A(n13966), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13982), .Z(
        P2_U3554) );
  MUX2_X1 U16057 ( .A(n13967), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13982), .Z(
        P2_U3553) );
  MUX2_X1 U16058 ( .A(n13968), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13982), .Z(
        P2_U3552) );
  MUX2_X1 U16059 ( .A(n13969), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13982), .Z(
        P2_U3551) );
  MUX2_X1 U16060 ( .A(n13970), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13982), .Z(
        P2_U3550) );
  MUX2_X1 U16061 ( .A(n13971), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13982), .Z(
        P2_U3549) );
  MUX2_X1 U16062 ( .A(n14231), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13982), .Z(
        P2_U3548) );
  INV_X2 U16063 ( .A(P2_U3947), .ZN(n13982) );
  MUX2_X1 U16064 ( .A(n14253), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13982), .Z(
        P2_U3547) );
  MUX2_X1 U16065 ( .A(n14268), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13982), .Z(
        P2_U3546) );
  MUX2_X1 U16066 ( .A(n14254), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13982), .Z(
        P2_U3545) );
  MUX2_X1 U16067 ( .A(n14269), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13982), .Z(
        P2_U3544) );
  MUX2_X1 U16068 ( .A(n14305), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13982), .Z(
        P2_U3543) );
  MUX2_X1 U16069 ( .A(n13972), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13982), .Z(
        P2_U3542) );
  MUX2_X1 U16070 ( .A(n14303), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13982), .Z(
        P2_U3541) );
  MUX2_X1 U16071 ( .A(n13973), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13982), .Z(
        P2_U3540) );
  MUX2_X1 U16072 ( .A(n13974), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13982), .Z(
        P2_U3539) );
  MUX2_X1 U16073 ( .A(n13975), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13982), .Z(
        P2_U3538) );
  MUX2_X1 U16074 ( .A(n13976), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13982), .Z(
        P2_U3537) );
  MUX2_X1 U16075 ( .A(n13977), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13982), .Z(
        P2_U3536) );
  MUX2_X1 U16076 ( .A(n13978), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13982), .Z(
        P2_U3535) );
  MUX2_X1 U16077 ( .A(n13979), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13982), .Z(
        P2_U3534) );
  MUX2_X1 U16078 ( .A(n13980), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13982), .Z(
        P2_U3533) );
  MUX2_X1 U16079 ( .A(n13981), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13982), .Z(
        P2_U3532) );
  MUX2_X1 U16080 ( .A(n10541), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13982), .Z(
        P2_U3531) );
  NAND2_X1 U16081 ( .A1(n13983), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n13986) );
  NAND2_X1 U16082 ( .A1(n13984), .A2(n13998), .ZN(n13985) );
  NAND2_X1 U16083 ( .A1(n13986), .A2(n13985), .ZN(n15578) );
  INV_X1 U16084 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n14237) );
  MUX2_X1 U16085 ( .A(n14237), .B(P2_REG2_REG_16__SCAN_IN), .S(n15585), .Z(
        n13987) );
  NAND2_X1 U16086 ( .A1(n15578), .A2(n13987), .ZN(n15601) );
  NAND2_X1 U16087 ( .A1(n13988), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n15600) );
  NAND2_X1 U16088 ( .A1(n15601), .A2(n15600), .ZN(n13991) );
  INV_X1 U16089 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13989) );
  MUX2_X1 U16090 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n13989), .S(n15598), .Z(
        n13990) );
  NAND2_X1 U16091 ( .A1(n13991), .A2(n13990), .ZN(n15604) );
  NAND2_X1 U16092 ( .A1(n15598), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13992) );
  NAND2_X1 U16093 ( .A1(n15604), .A2(n13992), .ZN(n13993) );
  OR2_X1 U16094 ( .A1(n13993), .A2(n14001), .ZN(n14010) );
  NAND2_X1 U16095 ( .A1(n13993), .A2(n14001), .ZN(n13994) );
  INV_X1 U16096 ( .A(n14011), .ZN(n13995) );
  AOI21_X1 U16097 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13996), .A(n13995), 
        .ZN(n14007) );
  AOI22_X1 U16098 ( .A1(n13999), .A2(n13998), .B1(P2_REG1_REG_15__SCAN_IN), 
        .B2(n13997), .ZN(n15583) );
  INV_X1 U16099 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14000) );
  XNOR2_X1 U16100 ( .A(n15585), .B(n14000), .ZN(n15582) );
  OAI22_X1 U16101 ( .A1(n15583), .A2(n15582), .B1(n14000), .B2(n15585), .ZN(
        n15593) );
  INV_X1 U16102 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14369) );
  XNOR2_X1 U16103 ( .A(n15598), .B(n14369), .ZN(n15594) );
  XNOR2_X1 U16104 ( .A(n14009), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n14005) );
  NAND2_X1 U16105 ( .A1(n15527), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n14002) );
  OAI211_X1 U16106 ( .C1(n15584), .C2(n14008), .A(n14003), .B(n14002), .ZN(
        n14004) );
  AOI21_X1 U16107 ( .B1(n14005), .B2(n15596), .A(n14004), .ZN(n14006) );
  OAI21_X1 U16108 ( .B1(n14007), .B2(n15579), .A(n14006), .ZN(P2_U3232) );
  INV_X1 U16109 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15922) );
  INV_X1 U16110 ( .A(n14016), .ZN(n14013) );
  NAND2_X1 U16111 ( .A1(n14011), .A2(n14010), .ZN(n14012) );
  XNOR2_X1 U16112 ( .A(n14012), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n14014) );
  AOI22_X1 U16113 ( .A1(n14013), .A2(n15596), .B1(n14014), .B2(n15603), .ZN(
        n14019) );
  NOR2_X1 U16114 ( .A1(n14014), .A2(n15579), .ZN(n14015) );
  AOI211_X1 U16115 ( .C1(n14016), .C2(n15596), .A(n14015), .B(n15595), .ZN(
        n14018) );
  MUX2_X1 U16116 ( .A(n14019), .B(n14018), .S(n14017), .Z(n14022) );
  INV_X1 U16117 ( .A(n14020), .ZN(n14021) );
  OAI211_X1 U16118 ( .C1(n7298), .C2(n15609), .A(n14022), .B(n14021), .ZN(
        P2_U3233) );
  NAND2_X1 U16119 ( .A1(n14023), .A2(n14282), .ZN(n14026) );
  INV_X1 U16120 ( .A(n14318), .ZN(n14024) );
  NOR2_X1 U16121 ( .A1(n14308), .A2(n14024), .ZN(n14032) );
  AOI21_X1 U16122 ( .B1(n14308), .B2(P2_REG2_REG_31__SCAN_IN), .A(n14032), 
        .ZN(n14025) );
  OAI211_X1 U16123 ( .C1(n14317), .C2(n14275), .A(n14026), .B(n14025), .ZN(
        P2_U3234) );
  INV_X1 U16124 ( .A(n14027), .ZN(n14030) );
  INV_X1 U16125 ( .A(n14028), .ZN(n14029) );
  NAND2_X1 U16126 ( .A1(n14319), .A2(n14282), .ZN(n14034) );
  AOI21_X1 U16127 ( .B1(n14308), .B2(P2_REG2_REG_30__SCAN_IN), .A(n14032), 
        .ZN(n14033) );
  OAI211_X1 U16128 ( .C1(n14411), .C2(n14275), .A(n14034), .B(n14033), .ZN(
        P2_U3235) );
  XOR2_X1 U16129 ( .A(n14043), .B(n14035), .Z(n14327) );
  INV_X1 U16130 ( .A(n14036), .ZN(n14073) );
  AOI21_X1 U16131 ( .B1(n14073), .B2(n14322), .A(n8582), .ZN(n14037) );
  AND2_X1 U16132 ( .A1(n14038), .A2(n14037), .ZN(n14323) );
  INV_X1 U16133 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n14039) );
  OAI22_X1 U16134 ( .A1(n14040), .A2(n14275), .B1(n14293), .B2(n14039), .ZN(
        n14041) );
  AOI21_X1 U16135 ( .B1(n14323), .B2(n14282), .A(n14041), .ZN(n14054) );
  NAND3_X1 U16136 ( .A1(n14045), .A2(n14307), .A3(n14044), .ZN(n14050) );
  NAND2_X1 U16137 ( .A1(n14046), .A2(n14302), .ZN(n14048) );
  AND2_X1 U16138 ( .A1(n14048), .A2(n7921), .ZN(n14049) );
  NOR2_X1 U16139 ( .A1(n14051), .A2(n14290), .ZN(n14052) );
  OAI21_X1 U16140 ( .B1(n14325), .B2(n14052), .A(n14293), .ZN(n14053) );
  OAI211_X1 U16141 ( .C1(n14327), .C2(n14279), .A(n14054), .B(n14053), .ZN(
        P2_U3237) );
  NAND2_X1 U16142 ( .A1(n14114), .A2(n14055), .ZN(n14061) );
  INV_X1 U16143 ( .A(n14056), .ZN(n14060) );
  INV_X1 U16144 ( .A(n14057), .ZN(n14058) );
  OR2_X1 U16145 ( .A1(n14068), .A2(n14058), .ZN(n14059) );
  AOI21_X1 U16146 ( .B1(n14061), .B2(n14060), .A(n14059), .ZN(n14062) );
  OAI22_X1 U16147 ( .A1(n14065), .A2(n14118), .B1(n14064), .B2(n14116), .ZN(
        n14066) );
  XNOR2_X1 U16148 ( .A(n14069), .B(n14068), .ZN(n14414) );
  INV_X1 U16149 ( .A(n14414), .ZN(n14070) );
  INV_X1 U16150 ( .A(n14279), .ZN(n14311) );
  NAND2_X1 U16151 ( .A1(n14070), .A2(n14311), .ZN(n14079) );
  INV_X1 U16152 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n14071) );
  OAI22_X1 U16153 ( .A1(n14072), .A2(n14290), .B1(n14071), .B2(n14293), .ZN(
        n14076) );
  OAI211_X1 U16154 ( .C1(n14413), .C2(n14074), .A(n14073), .B(n14239), .ZN(
        n14328) );
  NOR2_X1 U16155 ( .A1(n14328), .A2(n14297), .ZN(n14075) );
  AOI211_X1 U16156 ( .C1(n14295), .C2(n14077), .A(n14076), .B(n14075), .ZN(
        n14078) );
  OAI211_X1 U16157 ( .C1(n14308), .C2(n14329), .A(n14079), .B(n14078), .ZN(
        P2_U3238) );
  AOI22_X1 U16158 ( .A1(n14080), .A2(n14272), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14308), .ZN(n14081) );
  OAI21_X1 U16159 ( .B1(n14082), .B2(n14275), .A(n14081), .ZN(n14083) );
  AOI21_X1 U16160 ( .B1(n14084), .B2(n14282), .A(n14083), .ZN(n14087) );
  NAND2_X1 U16161 ( .A1(n14085), .A2(n14293), .ZN(n14086) );
  OAI211_X1 U16162 ( .C1(n14088), .C2(n14279), .A(n14087), .B(n14086), .ZN(
        P2_U3239) );
  NAND2_X1 U16163 ( .A1(n14089), .A2(n14293), .ZN(n14096) );
  AOI22_X1 U16164 ( .A1(n14090), .A2(n14272), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14308), .ZN(n14091) );
  OAI21_X1 U16165 ( .B1(n14092), .B2(n14275), .A(n14091), .ZN(n14093) );
  AOI21_X1 U16166 ( .B1(n14094), .B2(n14282), .A(n14093), .ZN(n14095) );
  OAI211_X1 U16167 ( .C1(n14097), .C2(n14279), .A(n14096), .B(n14095), .ZN(
        P2_U3240) );
  AND2_X1 U16168 ( .A1(n14121), .A2(n14098), .ZN(n14100) );
  OAI21_X1 U16169 ( .B1(n14100), .B2(n14103), .A(n14099), .ZN(n14102) );
  AOI21_X1 U16170 ( .B1(n14102), .B2(n14307), .A(n14101), .ZN(n14333) );
  XNOR2_X1 U16171 ( .A(n14104), .B(n14103), .ZN(n14419) );
  INV_X1 U16172 ( .A(n14419), .ZN(n14112) );
  OAI211_X1 U16173 ( .C1(n14128), .C2(n14418), .A(n14239), .B(n14105), .ZN(
        n14332) );
  OAI22_X1 U16174 ( .A1(n14107), .A2(n14290), .B1(n14106), .B2(n14293), .ZN(
        n14108) );
  AOI21_X1 U16175 ( .B1(n14109), .B2(n14295), .A(n14108), .ZN(n14110) );
  OAI21_X1 U16176 ( .B1(n14332), .B2(n14297), .A(n14110), .ZN(n14111) );
  AOI21_X1 U16177 ( .B1(n14112), .B2(n14311), .A(n14111), .ZN(n14113) );
  OAI21_X1 U16178 ( .B1(n14333), .B2(n14308), .A(n14113), .ZN(P2_U3241) );
  INV_X1 U16179 ( .A(n14114), .ZN(n14115) );
  AOI21_X1 U16180 ( .B1(n14115), .B2(n14124), .A(n14217), .ZN(n14122) );
  OAI22_X1 U16181 ( .A1(n14119), .A2(n14118), .B1(n14117), .B2(n14116), .ZN(
        n14120) );
  AOI21_X1 U16182 ( .B1(n14122), .B2(n14121), .A(n14120), .ZN(n14337) );
  OAI21_X1 U16183 ( .B1(n14123), .B2(n14290), .A(n14337), .ZN(n14133) );
  XNOR2_X1 U16184 ( .A(n7128), .B(n14124), .ZN(n14424) );
  NOR2_X1 U16185 ( .A1(n14424), .A2(n14279), .ZN(n14132) );
  OAI21_X1 U16186 ( .B1(n14126), .B2(n14423), .A(n14239), .ZN(n14127) );
  AOI22_X1 U16187 ( .A1(n14129), .A2(n14295), .B1(n14308), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n14130) );
  OAI21_X1 U16188 ( .B1(n14336), .B2(n14297), .A(n14130), .ZN(n14131) );
  AOI211_X1 U16189 ( .C1(n14133), .C2(n14293), .A(n14132), .B(n14131), .ZN(
        n14134) );
  INV_X1 U16190 ( .A(n14134), .ZN(P2_U3242) );
  XNOR2_X1 U16191 ( .A(n14135), .B(n14139), .ZN(n14137) );
  AOI21_X1 U16192 ( .B1(n14137), .B2(n14307), .A(n14136), .ZN(n14341) );
  OAI21_X1 U16193 ( .B1(n14140), .B2(n14139), .A(n14138), .ZN(n14429) );
  INV_X1 U16194 ( .A(n14429), .ZN(n14148) );
  INV_X1 U16195 ( .A(n14126), .ZN(n14141) );
  OAI211_X1 U16196 ( .C1(n14428), .C2(n14164), .A(n14141), .B(n14239), .ZN(
        n14340) );
  OAI22_X1 U16197 ( .A1(n14143), .A2(n14290), .B1(n14293), .B2(n14142), .ZN(
        n14144) );
  AOI21_X1 U16198 ( .B1(n14145), .B2(n14295), .A(n14144), .ZN(n14146) );
  OAI21_X1 U16199 ( .B1(n14340), .B2(n14297), .A(n14146), .ZN(n14147) );
  AOI21_X1 U16200 ( .B1(n14148), .B2(n14311), .A(n14147), .ZN(n14149) );
  OAI21_X1 U16201 ( .B1(n14341), .B2(n14308), .A(n14149), .ZN(P2_U3243) );
  NOR2_X1 U16202 ( .A1(n14185), .A2(n14152), .ZN(n14188) );
  AND2_X1 U16203 ( .A1(n14196), .A2(n14153), .ZN(n14184) );
  NOR2_X1 U16204 ( .A1(n14188), .A2(n14184), .ZN(n14169) );
  OAI21_X1 U16205 ( .B1(n14169), .B2(n14172), .A(n14154), .ZN(n14155) );
  XNOR2_X1 U16206 ( .A(n14155), .B(n14161), .ZN(n14157) );
  AOI21_X1 U16207 ( .B1(n14157), .B2(n14307), .A(n14156), .ZN(n14350) );
  OR2_X1 U16208 ( .A1(n14350), .A2(n14308), .ZN(n14168) );
  OAI22_X1 U16209 ( .A1(n14293), .A2(n14159), .B1(n14158), .B2(n14290), .ZN(
        n14160) );
  AOI21_X1 U16210 ( .B1(n14345), .B2(n14295), .A(n14160), .ZN(n14167) );
  NAND2_X1 U16211 ( .A1(n6684), .A2(n14161), .ZN(n14346) );
  NAND3_X1 U16212 ( .A1(n6626), .A2(n14311), .A3(n14346), .ZN(n14166) );
  NAND2_X1 U16213 ( .A1(n14174), .A2(n14345), .ZN(n14162) );
  NAND2_X1 U16214 ( .A1(n14162), .A2(n14239), .ZN(n14163) );
  NOR2_X1 U16215 ( .A1(n14164), .A2(n14163), .ZN(n14344) );
  NAND2_X1 U16216 ( .A1(n14344), .A2(n14282), .ZN(n14165) );
  NAND4_X1 U16217 ( .A1(n14168), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        P2_U3244) );
  XNOR2_X1 U16218 ( .A(n14169), .B(n14172), .ZN(n14171) );
  AOI21_X1 U16219 ( .B1(n14171), .B2(n14307), .A(n14170), .ZN(n14352) );
  XNOR2_X1 U16220 ( .A(n14173), .B(n14172), .ZN(n14434) );
  INV_X1 U16221 ( .A(n14434), .ZN(n14181) );
  AOI21_X1 U16222 ( .B1(n14193), .B2(n14353), .A(n8582), .ZN(n14175) );
  NAND2_X1 U16223 ( .A1(n14175), .A2(n14174), .ZN(n14351) );
  INV_X1 U16224 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n14177) );
  OAI22_X1 U16225 ( .A1(n14293), .A2(n14177), .B1(n14176), .B2(n14290), .ZN(
        n14178) );
  AOI21_X1 U16226 ( .B1(n14353), .B2(n14295), .A(n14178), .ZN(n14179) );
  OAI21_X1 U16227 ( .B1(n14351), .B2(n14297), .A(n14179), .ZN(n14180) );
  AOI21_X1 U16228 ( .B1(n14181), .B2(n14311), .A(n14180), .ZN(n14182) );
  OAI21_X1 U16229 ( .B1(n14352), .B2(n14308), .A(n14182), .ZN(P2_U3245) );
  XOR2_X1 U16230 ( .A(n14183), .B(n14186), .Z(n14358) );
  INV_X1 U16231 ( .A(n14184), .ZN(n14187) );
  AOI22_X1 U16232 ( .A1(n14188), .A2(n14187), .B1(n14186), .B2(n14185), .ZN(
        n14189) );
  NOR2_X1 U16233 ( .A1(n14189), .A2(n14217), .ZN(n14360) );
  OAI21_X1 U16234 ( .B1(n14360), .B2(n14190), .A(n14293), .ZN(n14198) );
  INV_X1 U16235 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14192) );
  OAI22_X1 U16236 ( .A1(n14293), .A2(n14192), .B1(n14191), .B2(n14290), .ZN(
        n14195) );
  OAI211_X1 U16237 ( .C1(n6702), .C2(n14440), .A(n14239), .B(n14193), .ZN(
        n14356) );
  NOR2_X1 U16238 ( .A1(n14356), .A2(n14297), .ZN(n14194) );
  AOI211_X1 U16239 ( .C1(n14295), .C2(n14196), .A(n14195), .B(n14194), .ZN(
        n14197) );
  OAI211_X1 U16240 ( .C1(n14358), .C2(n14279), .A(n14198), .B(n14197), .ZN(
        P2_U3246) );
  XOR2_X1 U16241 ( .A(n14199), .B(n14200), .Z(n14444) );
  XOR2_X1 U16242 ( .A(n14201), .B(n14200), .Z(n14203) );
  OAI21_X1 U16243 ( .B1(n14203), .B2(n14217), .A(n14202), .ZN(n14363) );
  NAND2_X1 U16244 ( .A1(n14363), .A2(n14293), .ZN(n14212) );
  INV_X1 U16245 ( .A(n14204), .ZN(n14205) );
  AOI211_X1 U16246 ( .C1(n14365), .C2(n14205), .A(n8582), .B(n6702), .ZN(
        n14364) );
  INV_X1 U16247 ( .A(n14206), .ZN(n14207) );
  AOI22_X1 U16248 ( .A1(n14308), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14207), 
        .B2(n14272), .ZN(n14208) );
  OAI21_X1 U16249 ( .B1(n14209), .B2(n14275), .A(n14208), .ZN(n14210) );
  AOI21_X1 U16250 ( .B1(n14364), .B2(n14282), .A(n14210), .ZN(n14211) );
  OAI211_X1 U16251 ( .C1(n14444), .C2(n14279), .A(n14212), .B(n14211), .ZN(
        P2_U3247) );
  XNOR2_X1 U16252 ( .A(n14213), .B(n14214), .ZN(n14447) );
  XNOR2_X1 U16253 ( .A(n14215), .B(n14214), .ZN(n14218) );
  OAI21_X1 U16254 ( .B1(n14218), .B2(n14217), .A(n14216), .ZN(n14367) );
  NAND2_X1 U16255 ( .A1(n14367), .A2(n14293), .ZN(n14225) );
  NOR2_X1 U16256 ( .A1(n14242), .A2(n14222), .ZN(n14219) );
  AOI22_X1 U16257 ( .A1(n14308), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14220), 
        .B2(n14272), .ZN(n14221) );
  OAI21_X1 U16258 ( .B1(n14222), .B2(n14275), .A(n14221), .ZN(n14223) );
  AOI21_X1 U16259 ( .B1(n6604), .B2(n14282), .A(n14223), .ZN(n14224) );
  OAI211_X1 U16260 ( .C1(n14447), .C2(n14279), .A(n14225), .B(n14224), .ZN(
        P2_U3248) );
  XNOR2_X1 U16261 ( .A(n14226), .B(n14227), .ZN(n14234) );
  NAND2_X1 U16262 ( .A1(n14228), .A2(n14227), .ZN(n14229) );
  NAND2_X1 U16263 ( .A1(n14230), .A2(n14229), .ZN(n14375) );
  AOI22_X1 U16264 ( .A1(n14302), .A2(n14268), .B1(n14231), .B2(n14304), .ZN(
        n14232) );
  OAI21_X1 U16265 ( .B1(n14375), .B2(n15642), .A(n14232), .ZN(n14233) );
  AOI21_X1 U16266 ( .B1(n14234), .B2(n14307), .A(n14233), .ZN(n14374) );
  INV_X1 U16267 ( .A(n14235), .ZN(n14236) );
  OAI22_X1 U16268 ( .A1(n14293), .A2(n14237), .B1(n14236), .B2(n14290), .ZN(
        n14238) );
  AOI21_X1 U16269 ( .B1(n14372), .B2(n14295), .A(n14238), .ZN(n14244) );
  NAND2_X1 U16270 ( .A1(n14257), .A2(n14372), .ZN(n14240) );
  NAND2_X1 U16271 ( .A1(n14240), .A2(n14239), .ZN(n14241) );
  NOR2_X1 U16272 ( .A1(n14242), .A2(n14241), .ZN(n14371) );
  NAND2_X1 U16273 ( .A1(n14371), .A2(n14282), .ZN(n14243) );
  OAI211_X1 U16274 ( .C1(n14375), .C2(n14265), .A(n14244), .B(n14243), .ZN(
        n14245) );
  INV_X1 U16275 ( .A(n14245), .ZN(n14246) );
  OAI21_X1 U16276 ( .B1(n14374), .B2(n14308), .A(n14246), .ZN(P2_U3249) );
  INV_X1 U16277 ( .A(n14247), .ZN(n14248) );
  AOI21_X1 U16278 ( .B1(n14250), .B2(n14249), .A(n14248), .ZN(n14376) );
  XNOR2_X1 U16279 ( .A(n14251), .B(n14250), .ZN(n14252) );
  NAND2_X1 U16280 ( .A1(n14252), .A2(n14307), .ZN(n14256) );
  AOI22_X1 U16281 ( .A1(n14302), .A2(n14254), .B1(n14253), .B2(n14304), .ZN(
        n14255) );
  OAI211_X1 U16282 ( .C1(n14376), .C2(n15642), .A(n14256), .B(n14255), .ZN(
        n14377) );
  NAND2_X1 U16283 ( .A1(n14377), .A2(n14293), .ZN(n14264) );
  INV_X1 U16284 ( .A(n14257), .ZN(n14258) );
  AOI211_X1 U16285 ( .C1(n14259), .C2(n14270), .A(n8582), .B(n14258), .ZN(
        n14378) );
  AOI22_X1 U16286 ( .A1(n14308), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14260), 
        .B2(n14272), .ZN(n14261) );
  OAI21_X1 U16287 ( .B1(n7850), .B2(n14275), .A(n14261), .ZN(n14262) );
  AOI21_X1 U16288 ( .B1(n14378), .B2(n14282), .A(n14262), .ZN(n14263) );
  OAI211_X1 U16289 ( .C1(n14376), .C2(n14265), .A(n14264), .B(n14263), .ZN(
        P2_U3250) );
  XOR2_X1 U16290 ( .A(n14277), .B(n14266), .Z(n14267) );
  AOI222_X1 U16291 ( .A1(n14269), .A2(n14302), .B1(n14268), .B2(n14304), .C1(
        n14307), .C2(n14267), .ZN(n14385) );
  INV_X1 U16292 ( .A(n12188), .ZN(n14271) );
  AOI211_X1 U16293 ( .C1(n14383), .C2(n14271), .A(n8582), .B(n7851), .ZN(
        n14382) );
  AOI22_X1 U16294 ( .A1(n14308), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n14273), 
        .B2(n14272), .ZN(n14274) );
  OAI21_X1 U16295 ( .B1(n14276), .B2(n14275), .A(n14274), .ZN(n14281) );
  XNOR2_X1 U16296 ( .A(n14278), .B(n14277), .ZN(n14386) );
  NOR2_X1 U16297 ( .A1(n14386), .A2(n14279), .ZN(n14280) );
  AOI211_X1 U16298 ( .C1(n14382), .C2(n14282), .A(n14281), .B(n14280), .ZN(
        n14283) );
  OAI21_X1 U16299 ( .B1(n14385), .B2(n14308), .A(n14283), .ZN(P2_U3251) );
  OR2_X1 U16300 ( .A1(n14284), .A2(n14299), .ZN(n14285) );
  NAND2_X1 U16301 ( .A1(n14286), .A2(n14285), .ZN(n14462) );
  INV_X1 U16302 ( .A(n14462), .ZN(n14312) );
  AOI21_X1 U16303 ( .B1(n14287), .B2(n14399), .A(n8582), .ZN(n14289) );
  NAND2_X1 U16304 ( .A1(n14289), .A2(n14288), .ZN(n14397) );
  OAI22_X1 U16305 ( .A1(n14293), .A2(n14292), .B1(n14291), .B2(n14290), .ZN(
        n14294) );
  AOI21_X1 U16306 ( .B1(n14295), .B2(n14399), .A(n14294), .ZN(n14296) );
  OAI21_X1 U16307 ( .B1(n14397), .B2(n14297), .A(n14296), .ZN(n14310) );
  NAND3_X1 U16308 ( .A1(n11954), .A2(n14299), .A3(n14298), .ZN(n14300) );
  NAND2_X1 U16309 ( .A1(n14301), .A2(n14300), .ZN(n14306) );
  AOI222_X1 U16310 ( .A1(n14307), .A2(n14306), .B1(n14305), .B2(n14304), .C1(
        n14303), .C2(n14302), .ZN(n14398) );
  NOR2_X1 U16311 ( .A1(n14398), .A2(n14308), .ZN(n14309) );
  AOI211_X1 U16312 ( .C1(n14312), .C2(n14311), .A(n14310), .B(n14309), .ZN(
        n14313) );
  INV_X1 U16313 ( .A(n14313), .ZN(P2_U3254) );
  INV_X1 U16314 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14315) );
  OAI21_X1 U16315 ( .B1(n14317), .B2(n14400), .A(n14316), .ZN(P2_U3530) );
  INV_X1 U16316 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14320) );
  NOR2_X1 U16317 ( .A1(n14319), .A2(n14318), .ZN(n14409) );
  OAI21_X1 U16318 ( .B1(n14411), .B2(n14400), .A(n14321), .ZN(P2_U3529) );
  OAI21_X1 U16319 ( .B1(n14327), .B2(n15655), .A(n14326), .ZN(n14412) );
  MUX2_X1 U16320 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14412), .S(n15670), .Z(
        P2_U3527) );
  OAI22_X1 U16321 ( .A1(n14414), .A2(n14401), .B1(n14413), .B2(n14400), .ZN(
        n14331) );
  MUX2_X1 U16322 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14415), .S(n15670), .Z(
        n14330) );
  OR2_X1 U16323 ( .A1(n14331), .A2(n14330), .ZN(P2_U3526) );
  NAND2_X1 U16324 ( .A1(n14333), .A2(n14332), .ZN(n14417) );
  MUX2_X1 U16325 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14417), .S(n15670), .Z(
        n14335) );
  OAI22_X1 U16326 ( .A1(n14419), .A2(n14401), .B1(n14418), .B2(n14400), .ZN(
        n14334) );
  OR2_X1 U16327 ( .A1(n14335), .A2(n14334), .ZN(P2_U3523) );
  NAND2_X1 U16328 ( .A1(n14337), .A2(n14336), .ZN(n14422) );
  MUX2_X1 U16329 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14422), .S(n15670), .Z(
        n14339) );
  OAI22_X1 U16330 ( .A1(n14424), .A2(n14401), .B1(n14423), .B2(n14400), .ZN(
        n14338) );
  OR2_X1 U16331 ( .A1(n14339), .A2(n14338), .ZN(P2_U3522) );
  NAND2_X1 U16332 ( .A1(n14341), .A2(n14340), .ZN(n14427) );
  MUX2_X1 U16333 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14427), .S(n15670), .Z(
        n14343) );
  OAI22_X1 U16334 ( .A1(n14429), .A2(n14401), .B1(n14428), .B2(n14400), .ZN(
        n14342) );
  OR2_X1 U16335 ( .A1(n14343), .A2(n14342), .ZN(P2_U3521) );
  AOI21_X1 U16336 ( .B1(n15651), .B2(n14345), .A(n14344), .ZN(n14349) );
  NAND3_X1 U16337 ( .A1(n6626), .A2(n14347), .A3(n14346), .ZN(n14348) );
  NAND3_X1 U16338 ( .A1(n14350), .A2(n14349), .A3(n14348), .ZN(n14432) );
  MUX2_X1 U16339 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14432), .S(n15670), .Z(
        P2_U3520) );
  NAND2_X1 U16340 ( .A1(n14352), .A2(n14351), .ZN(n14433) );
  MUX2_X1 U16341 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14433), .S(n15670), .Z(
        n14355) );
  OAI22_X1 U16342 ( .A1(n14434), .A2(n14401), .B1(n7855), .B2(n14400), .ZN(
        n14354) );
  OR2_X1 U16343 ( .A1(n14355), .A2(n14354), .ZN(P2_U3519) );
  INV_X1 U16344 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14361) );
  OAI211_X1 U16345 ( .C1(n14358), .C2(n15655), .A(n14357), .B(n14356), .ZN(
        n14359) );
  NOR2_X1 U16346 ( .A1(n14360), .A2(n14359), .ZN(n14437) );
  MUX2_X1 U16347 ( .A(n14361), .B(n14437), .S(n15670), .Z(n14362) );
  OAI21_X1 U16348 ( .B1(n14440), .B2(n14400), .A(n14362), .ZN(P2_U3518) );
  AOI211_X1 U16349 ( .C1(n15651), .C2(n14365), .A(n14364), .B(n14363), .ZN(
        n14441) );
  MUX2_X1 U16350 ( .A(n15922), .B(n14441), .S(n15670), .Z(n14366) );
  OAI21_X1 U16351 ( .B1(n14401), .B2(n14444), .A(n14366), .ZN(P2_U3517) );
  AOI211_X1 U16352 ( .C1(n15651), .C2(n14368), .A(n6604), .B(n14367), .ZN(
        n14445) );
  MUX2_X1 U16353 ( .A(n14369), .B(n14445), .S(n15670), .Z(n14370) );
  OAI21_X1 U16354 ( .B1(n14447), .B2(n14401), .A(n14370), .ZN(P2_U3516) );
  AOI21_X1 U16355 ( .B1(n15651), .B2(n14372), .A(n14371), .ZN(n14373) );
  OAI211_X1 U16356 ( .C1(n15636), .C2(n14375), .A(n14374), .B(n14373), .ZN(
        n14448) );
  MUX2_X1 U16357 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14448), .S(n15670), .Z(
        P2_U3515) );
  INV_X1 U16358 ( .A(n14376), .ZN(n14379) );
  AOI211_X1 U16359 ( .C1(n15646), .C2(n14379), .A(n14378), .B(n14377), .ZN(
        n14449) );
  MUX2_X1 U16360 ( .A(n14380), .B(n14449), .S(n15670), .Z(n14381) );
  OAI21_X1 U16361 ( .B1(n7850), .B2(n14400), .A(n14381), .ZN(P2_U3514) );
  AOI21_X1 U16362 ( .B1(n15651), .B2(n14383), .A(n14382), .ZN(n14384) );
  OAI211_X1 U16363 ( .C1(n15655), .C2(n14386), .A(n14385), .B(n14384), .ZN(
        n14452) );
  MUX2_X1 U16364 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14452), .S(n15670), .Z(
        P2_U3513) );
  INV_X1 U16365 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14390) );
  AOI211_X1 U16366 ( .C1(n15651), .C2(n14389), .A(n14388), .B(n14387), .ZN(
        n14453) );
  MUX2_X1 U16367 ( .A(n14390), .B(n14453), .S(n15670), .Z(n14391) );
  OAI21_X1 U16368 ( .B1(n14456), .B2(n14401), .A(n14391), .ZN(P2_U3512) );
  AOI21_X1 U16369 ( .B1(n15651), .B2(n14393), .A(n14392), .ZN(n14394) );
  OAI211_X1 U16370 ( .C1(n15655), .C2(n14396), .A(n14395), .B(n14394), .ZN(
        n14457) );
  MUX2_X1 U16371 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14457), .S(n15670), .Z(
        P2_U3511) );
  NAND2_X1 U16372 ( .A1(n14398), .A2(n14397), .ZN(n14458) );
  MUX2_X1 U16373 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14458), .S(n15670), .Z(
        n14403) );
  INV_X1 U16374 ( .A(n14399), .ZN(n14460) );
  OAI22_X1 U16375 ( .A1(n14462), .A2(n14401), .B1(n14460), .B2(n14400), .ZN(
        n14402) );
  OR2_X1 U16376 ( .A1(n14403), .A2(n14402), .ZN(P2_U3510) );
  AOI21_X1 U16377 ( .B1(n15651), .B2(n14405), .A(n14404), .ZN(n14406) );
  OAI211_X1 U16378 ( .C1(n15655), .C2(n14408), .A(n14407), .B(n14406), .ZN(
        n14465) );
  MUX2_X1 U16379 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14465), .S(n15670), .Z(
        P2_U3509) );
  OAI21_X1 U16380 ( .B1(n14411), .B2(n14459), .A(n14410), .ZN(P2_U3497) );
  MUX2_X1 U16381 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14412), .S(n15659), .Z(
        P2_U3495) );
  OAI22_X1 U16382 ( .A1(n14414), .A2(n14461), .B1(n14413), .B2(n14459), .ZN(
        n14416) );
  MUX2_X1 U16383 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14417), .S(n15659), .Z(
        n14421) );
  OAI22_X1 U16384 ( .A1(n14419), .A2(n14461), .B1(n14418), .B2(n14459), .ZN(
        n14420) );
  OR2_X1 U16385 ( .A1(n14421), .A2(n14420), .ZN(P2_U3491) );
  MUX2_X1 U16386 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14422), .S(n15659), .Z(
        n14426) );
  OAI22_X1 U16387 ( .A1(n14424), .A2(n14461), .B1(n14423), .B2(n14459), .ZN(
        n14425) );
  OR2_X1 U16388 ( .A1(n14426), .A2(n14425), .ZN(P2_U3490) );
  MUX2_X1 U16389 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14427), .S(n15659), .Z(
        n14431) );
  OAI22_X1 U16390 ( .A1(n14429), .A2(n14461), .B1(n14428), .B2(n14459), .ZN(
        n14430) );
  OR2_X1 U16391 ( .A1(n14431), .A2(n14430), .ZN(P2_U3489) );
  MUX2_X1 U16392 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14432), .S(n15659), .Z(
        P2_U3488) );
  MUX2_X1 U16393 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14433), .S(n15659), .Z(
        n14436) );
  OAI22_X1 U16394 ( .A1(n14434), .A2(n14461), .B1(n7855), .B2(n14459), .ZN(
        n14435) );
  OR2_X1 U16395 ( .A1(n14436), .A2(n14435), .ZN(P2_U3487) );
  INV_X1 U16396 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14438) );
  MUX2_X1 U16397 ( .A(n14438), .B(n14437), .S(n15659), .Z(n14439) );
  OAI21_X1 U16398 ( .B1(n14440), .B2(n14459), .A(n14439), .ZN(P2_U3486) );
  MUX2_X1 U16399 ( .A(n14442), .B(n14441), .S(n15659), .Z(n14443) );
  OAI21_X1 U16400 ( .B1(n14444), .B2(n14461), .A(n14443), .ZN(P2_U3484) );
  INV_X1 U16401 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n15735) );
  MUX2_X1 U16402 ( .A(n15735), .B(n14445), .S(n15659), .Z(n14446) );
  OAI21_X1 U16403 ( .B1(n14447), .B2(n14461), .A(n14446), .ZN(P2_U3481) );
  MUX2_X1 U16404 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14448), .S(n15659), .Z(
        P2_U3478) );
  INV_X1 U16405 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14450) );
  MUX2_X1 U16406 ( .A(n14450), .B(n14449), .S(n15659), .Z(n14451) );
  OAI21_X1 U16407 ( .B1(n7850), .B2(n14459), .A(n14451), .ZN(P2_U3475) );
  MUX2_X1 U16408 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14452), .S(n15659), .Z(
        P2_U3472) );
  INV_X1 U16409 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14454) );
  MUX2_X1 U16410 ( .A(n14454), .B(n14453), .S(n15659), .Z(n14455) );
  OAI21_X1 U16411 ( .B1(n14456), .B2(n14461), .A(n14455), .ZN(P2_U3469) );
  MUX2_X1 U16412 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14457), .S(n15659), .Z(
        P2_U3466) );
  MUX2_X1 U16413 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n14458), .S(n15659), .Z(
        n14464) );
  OAI22_X1 U16414 ( .A1(n14462), .A2(n14461), .B1(n14460), .B2(n14459), .ZN(
        n14463) );
  OR2_X1 U16415 ( .A1(n14464), .A2(n14463), .ZN(P2_U3463) );
  MUX2_X1 U16416 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n14465), .S(n15659), .Z(
        P2_U3460) );
  INV_X1 U16417 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14466) );
  NAND3_X1 U16418 ( .A1(n14466), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14468) );
  OAI22_X1 U16419 ( .A1(n8028), .A2(n14468), .B1(n14467), .B2(n14478), .ZN(
        n14469) );
  AOI21_X1 U16420 ( .B1(n12715), .B2(n14470), .A(n14469), .ZN(n14471) );
  INV_X1 U16421 ( .A(n14471), .ZN(P2_U3296) );
  AOI21_X1 U16422 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n14473), .A(n14472), 
        .ZN(n14474) );
  OAI21_X1 U16423 ( .B1(n14475), .B2(n10996), .A(n14474), .ZN(P2_U3299) );
  INV_X1 U16424 ( .A(n14476), .ZN(n14480) );
  INV_X1 U16425 ( .A(n14477), .ZN(n15235) );
  OAI222_X1 U16426 ( .A1(P2_U3088), .A2(n14480), .B1(n10996), .B2(n15235), 
        .C1(n14479), .C2(n14478), .ZN(P2_U3301) );
  MUX2_X1 U16427 ( .A(n14481), .B(n15497), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  XNOR2_X1 U16428 ( .A(n14483), .B(n14482), .ZN(n14488) );
  NAND2_X1 U16429 ( .A1(n14837), .A2(n14591), .ZN(n14485) );
  AOI22_X1 U16430 ( .A1(n14870), .A2(n14600), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(n6537), .ZN(n14484) );
  OAI211_X1 U16431 ( .C1(n14844), .C2(n14611), .A(n14485), .B(n14484), .ZN(
        n14486) );
  AOI21_X1 U16432 ( .B1(n15093), .B2(n14617), .A(n14486), .ZN(n14487) );
  OAI21_X1 U16433 ( .B1(n14488), .B2(n14619), .A(n14487), .ZN(P1_U3214) );
  INV_X1 U16434 ( .A(n14489), .ZN(n14490) );
  AOI21_X1 U16435 ( .B1(n14492), .B2(n14491), .A(n14490), .ZN(n14498) );
  AOI22_X1 U16436 ( .A1(n14600), .A2(n14639), .B1(n14630), .B2(n14493), .ZN(
        n14495) );
  OAI211_X1 U16437 ( .C1(n14541), .C2(n14613), .A(n14495), .B(n14494), .ZN(
        n14496) );
  AOI21_X1 U16438 ( .B1(n14617), .B2(n15175), .A(n14496), .ZN(n14497) );
  OAI21_X1 U16439 ( .B1(n14498), .B2(n14619), .A(n14497), .ZN(P1_U3215) );
  XOR2_X1 U16440 ( .A(n14500), .B(n14499), .Z(n14506) );
  OAI22_X1 U16441 ( .A1(n14609), .A2(n14944), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14501), .ZN(n14504) );
  INV_X1 U16442 ( .A(n14914), .ZN(n14502) );
  OAI22_X1 U16443 ( .A1(n14526), .A2(n14613), .B1(n14502), .B2(n14611), .ZN(
        n14503) );
  AOI211_X1 U16444 ( .C1(n15121), .C2(n14617), .A(n14504), .B(n14503), .ZN(
        n14505) );
  OAI21_X1 U16445 ( .B1(n14506), .B2(n14619), .A(n14505), .ZN(P1_U3216) );
  OAI211_X1 U16446 ( .C1(n14509), .C2(n14508), .A(n14507), .B(n14621), .ZN(
        n14514) );
  NAND2_X1 U16447 ( .A1(n14637), .A2(n15031), .ZN(n14511) );
  NAND2_X1 U16448 ( .A1(n15015), .A2(n15029), .ZN(n14510) );
  NAND2_X1 U16449 ( .A1(n14511), .A2(n14510), .ZN(n15149) );
  AND2_X1 U16450 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14812) );
  NOR2_X1 U16451 ( .A1(n14611), .A2(n14986), .ZN(n14512) );
  AOI211_X1 U16452 ( .C1(n14571), .C2(n15149), .A(n14812), .B(n14512), .ZN(
        n14513) );
  OAI211_X1 U16453 ( .C1(n7119), .C2(n14633), .A(n14514), .B(n14513), .ZN(
        P1_U3219) );
  OAI21_X1 U16454 ( .B1(n14517), .B2(n14516), .A(n14515), .ZN(n14518) );
  NAND2_X1 U16455 ( .A1(n14518), .A2(n14621), .ZN(n14522) );
  NOR2_X1 U16456 ( .A1(n14613), .A2(n14944), .ZN(n14520) );
  OAI22_X1 U16457 ( .A1(n14609), .A2(n14942), .B1(n14952), .B2(n14611), .ZN(
        n14519) );
  AOI211_X1 U16458 ( .C1(P1_REG3_REG_21__SCAN_IN), .C2(P1_U3086), .A(n14520), 
        .B(n14519), .ZN(n14521) );
  OAI211_X1 U16459 ( .C1(n15135), .C2(n14633), .A(n14522), .B(n14521), .ZN(
        P1_U3223) );
  XOR2_X1 U16460 ( .A(n14524), .B(n14523), .Z(n14531) );
  OAI22_X1 U16461 ( .A1(n14526), .A2(n14609), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14525), .ZN(n14529) );
  OAI22_X1 U16462 ( .A1(n14527), .A2(n14613), .B1(n14874), .B2(n14611), .ZN(
        n14528) );
  AOI211_X1 U16463 ( .C1(n14879), .C2(n14617), .A(n14529), .B(n14528), .ZN(
        n14530) );
  OAI21_X1 U16464 ( .B1(n14531), .B2(n14619), .A(n14530), .ZN(P1_U3225) );
  XNOR2_X1 U16465 ( .A(n14533), .B(n14532), .ZN(n14538) );
  XOR2_X1 U16466 ( .A(n14535), .B(n14536), .Z(n14624) );
  INV_X1 U16467 ( .A(n14534), .ZN(n14623) );
  NAND2_X1 U16468 ( .A1(n14624), .A2(n14623), .ZN(n14622) );
  OAI21_X1 U16469 ( .B1(n14536), .B2(n14535), .A(n14622), .ZN(n14537) );
  NOR2_X1 U16470 ( .A1(n14537), .A2(n14538), .ZN(n14549) );
  AOI21_X1 U16471 ( .B1(n14538), .B2(n14537), .A(n14549), .ZN(n14545) );
  OAI21_X1 U16472 ( .B1(n14613), .B2(n14540), .A(n14539), .ZN(n14543) );
  OAI22_X1 U16473 ( .A1(n14609), .A2(n14541), .B1(n15036), .B2(n14611), .ZN(
        n14542) );
  AOI211_X1 U16474 ( .C1(n14617), .C2(n15166), .A(n14543), .B(n14542), .ZN(
        n14544) );
  OAI21_X1 U16475 ( .B1(n14545), .B2(n14619), .A(n14544), .ZN(P1_U3226) );
  INV_X1 U16476 ( .A(n15161), .ZN(n15022) );
  INV_X1 U16477 ( .A(n14546), .ZN(n14548) );
  NOR3_X1 U16478 ( .A1(n14549), .A2(n14548), .A3(n14547), .ZN(n14552) );
  INV_X1 U16479 ( .A(n14550), .ZN(n14551) );
  OAI21_X1 U16480 ( .B1(n14552), .B2(n14551), .A(n14621), .ZN(n14558) );
  INV_X1 U16481 ( .A(n14553), .ZN(n14556) );
  OAI22_X1 U16482 ( .A1(n14609), .A2(n14554), .B1(n15019), .B2(n14611), .ZN(
        n14555) );
  AOI211_X1 U16483 ( .C1(n14591), .C2(n15015), .A(n14556), .B(n14555), .ZN(
        n14557) );
  OAI211_X1 U16484 ( .C1(n15022), .C2(n14633), .A(n14558), .B(n14557), .ZN(
        P1_U3228) );
  XOR2_X1 U16485 ( .A(n14560), .B(n14559), .Z(n14565) );
  OAI22_X1 U16486 ( .A1(n14889), .A2(n14609), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14561), .ZN(n14563) );
  OAI22_X1 U16487 ( .A1(n14610), .A2(n14613), .B1(n14894), .B2(n14611), .ZN(
        n14562) );
  AOI211_X1 U16488 ( .C1(n15111), .C2(n14617), .A(n14563), .B(n14562), .ZN(
        n14564) );
  OAI21_X1 U16489 ( .B1(n14565), .B2(n14619), .A(n14564), .ZN(P1_U3229) );
  XOR2_X1 U16490 ( .A(n14567), .B(n14566), .Z(n14568) );
  NAND2_X1 U16491 ( .A1(n14568), .A2(n14621), .ZN(n14576) );
  NAND2_X1 U16492 ( .A1(n14649), .A2(n15029), .ZN(n14570) );
  NAND2_X1 U16493 ( .A1(n14647), .A2(n15031), .ZN(n14569) );
  NAND2_X1 U16494 ( .A1(n14570), .A2(n14569), .ZN(n15369) );
  AND2_X1 U16495 ( .A1(n6537), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n15341) );
  AOI21_X1 U16496 ( .B1(n14571), .B2(n15369), .A(n15341), .ZN(n14575) );
  NAND2_X1 U16497 ( .A1(n14617), .A2(n14572), .ZN(n14574) );
  NAND2_X1 U16498 ( .A1(n14630), .A2(n15371), .ZN(n14573) );
  NAND4_X1 U16499 ( .A1(n14576), .A2(n14575), .A3(n14574), .A4(n14573), .ZN(
        P1_U3230) );
  OAI21_X1 U16500 ( .B1(n14578), .B2(n14577), .A(n14621), .ZN(n14585) );
  OAI22_X1 U16501 ( .A1(n14613), .A2(n14580), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14579), .ZN(n14582) );
  OAI22_X1 U16502 ( .A1(n14609), .A2(n14602), .B1(n14968), .B2(n14611), .ZN(
        n14581) );
  AOI211_X1 U16503 ( .C1(n15143), .C2(n14617), .A(n14582), .B(n14581), .ZN(
        n14583) );
  OAI21_X1 U16504 ( .B1(n14585), .B2(n14584), .A(n14583), .ZN(P1_U3233) );
  OAI21_X1 U16505 ( .B1(n14588), .B2(n14587), .A(n14586), .ZN(n14596) );
  NOR2_X1 U16506 ( .A1(n14589), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14590) );
  AOI21_X1 U16507 ( .B1(n14930), .B2(n14591), .A(n14590), .ZN(n14594) );
  INV_X1 U16508 ( .A(n14931), .ZN(n14592) );
  AOI22_X1 U16509 ( .A1(n14600), .A2(n14964), .B1(n14630), .B2(n14592), .ZN(
        n14593) );
  OAI211_X1 U16510 ( .C1(n15129), .C2(n14633), .A(n14594), .B(n14593), .ZN(
        n14595) );
  AOI21_X1 U16511 ( .B1(n14596), .B2(n14621), .A(n14595), .ZN(n14597) );
  INV_X1 U16512 ( .A(n14597), .ZN(P1_U3235) );
  XOR2_X1 U16513 ( .A(n14599), .B(n14598), .Z(n14605) );
  AOI22_X1 U16514 ( .A1(n14600), .A2(n15032), .B1(n14630), .B2(n15000), .ZN(
        n14601) );
  NAND2_X1 U16515 ( .A1(n6537), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14786) );
  OAI211_X1 U16516 ( .C1(n14602), .C2(n14613), .A(n14601), .B(n14786), .ZN(
        n14603) );
  AOI21_X1 U16517 ( .B1(n15156), .B2(n14617), .A(n14603), .ZN(n14604) );
  OAI21_X1 U16518 ( .B1(n14605), .B2(n14619), .A(n14604), .ZN(P1_U3238) );
  OAI22_X1 U16519 ( .A1(n14610), .A2(n14609), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14608), .ZN(n14616) );
  INV_X1 U16520 ( .A(n14857), .ZN(n14612) );
  OAI22_X1 U16521 ( .A1(n14614), .A2(n14613), .B1(n14612), .B2(n14611), .ZN(
        n14615) );
  AOI211_X1 U16522 ( .C1(n14860), .C2(n14617), .A(n14616), .B(n14615), .ZN(
        n14618) );
  OAI21_X1 U16523 ( .B1(n14620), .B2(n14619), .A(n14618), .ZN(P1_U3240) );
  INV_X1 U16524 ( .A(n15171), .ZN(n15054) );
  OAI211_X1 U16525 ( .C1(n14624), .C2(n14623), .A(n14622), .B(n14621), .ZN(
        n14632) );
  INV_X1 U16526 ( .A(n14625), .ZN(n15052) );
  AND2_X1 U16527 ( .A1(n14638), .A2(n15029), .ZN(n14626) );
  AOI21_X1 U16528 ( .B1(n15016), .B2(n15031), .A(n14626), .ZN(n15047) );
  OAI21_X1 U16529 ( .B1(n14628), .B2(n15047), .A(n14627), .ZN(n14629) );
  AOI21_X1 U16530 ( .B1(n15052), .B2(n14630), .A(n14629), .ZN(n14631) );
  OAI211_X1 U16531 ( .C1(n15054), .C2(n14633), .A(n14632), .B(n14631), .ZN(
        P1_U3241) );
  MUX2_X1 U16532 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14822), .S(n14666), .Z(
        P1_U3591) );
  MUX2_X1 U16533 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14634), .S(n14666), .Z(
        P1_U3590) );
  MUX2_X1 U16534 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14635), .S(n14666), .Z(
        P1_U3589) );
  MUX2_X1 U16535 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14837), .S(n14666), .Z(
        P1_U3588) );
  MUX2_X1 U16536 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14856), .S(n14666), .Z(
        P1_U3587) );
  MUX2_X1 U16537 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14870), .S(n14666), .Z(
        P1_U3586) );
  MUX2_X1 U16538 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14887), .S(n14666), .Z(
        P1_U3585) );
  MUX2_X1 U16539 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14907), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16540 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14930), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16541 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14636), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16542 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14964), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16543 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14637), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16544 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14993), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16545 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15015), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16546 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15032), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16547 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15016), .S(n14666), .Z(
        P1_U3576) );
  MUX2_X1 U16548 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15030), .S(n14666), .Z(
        P1_U3575) );
  MUX2_X1 U16549 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14638), .S(n14666), .Z(
        P1_U3574) );
  MUX2_X1 U16550 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14639), .S(n14666), .Z(
        P1_U3573) );
  MUX2_X1 U16551 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14640), .S(n14666), .Z(
        P1_U3572) );
  MUX2_X1 U16552 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14641), .S(n14666), .Z(
        P1_U3571) );
  MUX2_X1 U16553 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14642), .S(n14666), .Z(
        P1_U3570) );
  MUX2_X1 U16554 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14643), .S(n14666), .Z(
        P1_U3569) );
  MUX2_X1 U16555 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14644), .S(n14666), .Z(
        P1_U3568) );
  MUX2_X1 U16556 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14645), .S(n14666), .Z(
        P1_U3567) );
  MUX2_X1 U16557 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14646), .S(n14666), .Z(
        P1_U3566) );
  MUX2_X1 U16558 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14647), .S(n14666), .Z(
        P1_U3565) );
  MUX2_X1 U16559 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14648), .S(n14666), .Z(
        P1_U3564) );
  MUX2_X1 U16560 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14649), .S(n14666), .Z(
        P1_U3563) );
  MUX2_X1 U16561 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14650), .S(n14666), .Z(
        P1_U3562) );
  MUX2_X1 U16562 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n11669), .S(n14666), .Z(
        P1_U3561) );
  OAI211_X1 U16563 ( .C1(n14663), .C2(n14651), .A(n15338), .B(n14670), .ZN(
        n14661) );
  MUX2_X1 U16564 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10623), .S(n14656), .Z(
        n14652) );
  OAI21_X1 U16565 ( .B1(n14654), .B2(n14653), .A(n14652), .ZN(n14655) );
  NAND3_X1 U16566 ( .A1(n15332), .A2(n14678), .A3(n14655), .ZN(n14660) );
  INV_X1 U16567 ( .A(n14656), .ZN(n14657) );
  NAND2_X1 U16568 ( .A1(n15340), .A2(n14657), .ZN(n14659) );
  AOI22_X1 U16569 ( .A1(n15342), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n6537), .ZN(n14658) );
  NAND4_X1 U16570 ( .A1(n14661), .A2(n14660), .A3(n14659), .A4(n14658), .ZN(
        P1_U3244) );
  MUX2_X1 U16571 ( .A(n14663), .B(n14662), .S(n15230), .Z(n14665) );
  NAND2_X1 U16572 ( .A1(n14665), .A2(n14664), .ZN(n14667) );
  OAI211_X1 U16573 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14668), .A(n14667), .B(
        n14666), .ZN(n15347) );
  AOI22_X1 U16574 ( .A1(n15342), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14683) );
  MUX2_X1 U16575 ( .A(n10587), .B(P1_REG2_REG_2__SCAN_IN), .S(n14676), .Z(
        n14671) );
  NAND3_X1 U16576 ( .A1(n14671), .A2(n14670), .A3(n14669), .ZN(n14672) );
  NAND2_X1 U16577 ( .A1(n14688), .A2(n14672), .ZN(n14673) );
  OAI22_X1 U16578 ( .A1(n14674), .A2(n14804), .B1(n14805), .B2(n14673), .ZN(
        n14675) );
  INV_X1 U16579 ( .A(n14675), .ZN(n14682) );
  MUX2_X1 U16580 ( .A(n10626), .B(P1_REG1_REG_2__SCAN_IN), .S(n14676), .Z(
        n14679) );
  NAND3_X1 U16581 ( .A1(n14679), .A2(n14678), .A3(n14677), .ZN(n14680) );
  NAND3_X1 U16582 ( .A1(n15332), .A2(n14693), .A3(n14680), .ZN(n14681) );
  NAND4_X1 U16583 ( .A1(n15347), .A2(n14683), .A3(n14682), .A4(n14681), .ZN(
        P1_U3245) );
  OAI21_X1 U16584 ( .B1(n14815), .B2(n14685), .A(n14684), .ZN(n14686) );
  AOI21_X1 U16585 ( .B1(n14691), .B2(n15340), .A(n14686), .ZN(n14698) );
  MUX2_X1 U16586 ( .A(n10585), .B(P1_REG2_REG_3__SCAN_IN), .S(n14691), .Z(
        n14689) );
  NAND3_X1 U16587 ( .A1(n14689), .A2(n14688), .A3(n14687), .ZN(n14690) );
  NAND3_X1 U16588 ( .A1(n15338), .A2(n15335), .A3(n14690), .ZN(n14697) );
  MUX2_X1 U16589 ( .A(n10622), .B(P1_REG1_REG_3__SCAN_IN), .S(n14691), .Z(
        n14694) );
  NAND3_X1 U16590 ( .A1(n14694), .A2(n14693), .A3(n14692), .ZN(n14695) );
  NAND3_X1 U16591 ( .A1(n15332), .A2(n15329), .A3(n14695), .ZN(n14696) );
  NAND3_X1 U16592 ( .A1(n14698), .A2(n14697), .A3(n14696), .ZN(P1_U3246) );
  OAI21_X1 U16593 ( .B1(n14815), .B2(n14700), .A(n14699), .ZN(n14701) );
  AOI21_X1 U16594 ( .B1(n14706), .B2(n15340), .A(n14701), .ZN(n14712) );
  OAI21_X1 U16595 ( .B1(n14704), .B2(n14703), .A(n14702), .ZN(n14705) );
  NAND2_X1 U16596 ( .A1(n15332), .A2(n14705), .ZN(n14711) );
  MUX2_X1 U16597 ( .A(n10594), .B(P1_REG2_REG_5__SCAN_IN), .S(n14706), .Z(
        n14707) );
  NAND3_X1 U16598 ( .A1(n15337), .A2(n14708), .A3(n14707), .ZN(n14709) );
  NAND3_X1 U16599 ( .A1(n15338), .A2(n14719), .A3(n14709), .ZN(n14710) );
  NAND3_X1 U16600 ( .A1(n14712), .A2(n14711), .A3(n14710), .ZN(P1_U3248) );
  OAI21_X1 U16601 ( .B1(n14815), .B2(n14714), .A(n14713), .ZN(n14715) );
  AOI21_X1 U16602 ( .B1(n14716), .B2(n15340), .A(n14715), .ZN(n14726) );
  MUX2_X1 U16603 ( .A(n10597), .B(P1_REG2_REG_6__SCAN_IN), .S(n14716), .Z(
        n14717) );
  NAND3_X1 U16604 ( .A1(n14719), .A2(n14718), .A3(n14717), .ZN(n14720) );
  NAND3_X1 U16605 ( .A1(n15338), .A2(n14732), .A3(n14720), .ZN(n14725) );
  NAND2_X1 U16606 ( .A1(n14722), .A2(n14721), .ZN(n14723) );
  NAND3_X1 U16607 ( .A1(n15332), .A2(n14737), .A3(n14723), .ZN(n14724) );
  NAND3_X1 U16608 ( .A1(n14726), .A2(n14725), .A3(n14724), .ZN(P1_U3249) );
  INV_X1 U16609 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14728) );
  OAI21_X1 U16610 ( .B1(n14815), .B2(n14728), .A(n14727), .ZN(n14729) );
  AOI21_X1 U16611 ( .B1(n14734), .B2(n15340), .A(n14729), .ZN(n14742) );
  MUX2_X1 U16612 ( .A(n11692), .B(P1_REG2_REG_7__SCAN_IN), .S(n14734), .Z(
        n14730) );
  NAND3_X1 U16613 ( .A1(n14732), .A2(n14731), .A3(n14730), .ZN(n14733) );
  NAND3_X1 U16614 ( .A1(n15338), .A2(n14753), .A3(n14733), .ZN(n14741) );
  MUX2_X1 U16615 ( .A(n10636), .B(P1_REG1_REG_7__SCAN_IN), .S(n14734), .Z(
        n14735) );
  NAND3_X1 U16616 ( .A1(n14737), .A2(n14736), .A3(n14735), .ZN(n14738) );
  NAND3_X1 U16617 ( .A1(n15332), .A2(n14739), .A3(n14738), .ZN(n14740) );
  NAND3_X1 U16618 ( .A1(n14742), .A2(n14741), .A3(n14740), .ZN(P1_U3250) );
  INV_X1 U16619 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14744) );
  OAI21_X1 U16620 ( .B1(n14815), .B2(n14744), .A(n14743), .ZN(n14745) );
  AOI21_X1 U16621 ( .B1(n14750), .B2(n15340), .A(n14745), .ZN(n14758) );
  OAI21_X1 U16622 ( .B1(n14748), .B2(n14747), .A(n14746), .ZN(n14749) );
  NAND2_X1 U16623 ( .A1(n15332), .A2(n14749), .ZN(n14757) );
  MUX2_X1 U16624 ( .A(n11711), .B(P1_REG2_REG_8__SCAN_IN), .S(n14750), .Z(
        n14751) );
  NAND3_X1 U16625 ( .A1(n14753), .A2(n14752), .A3(n14751), .ZN(n14754) );
  NAND3_X1 U16626 ( .A1(n15338), .A2(n14755), .A3(n14754), .ZN(n14756) );
  NAND3_X1 U16627 ( .A1(n14758), .A2(n14757), .A3(n14756), .ZN(P1_U3251) );
  INV_X1 U16628 ( .A(n14759), .ZN(n14764) );
  AOI21_X1 U16629 ( .B1(n14762), .B2(n14761), .A(n14760), .ZN(n14763) );
  OAI21_X1 U16630 ( .B1(n14764), .B2(n14763), .A(n15332), .ZN(n14776) );
  OAI21_X1 U16631 ( .B1(n14815), .B2(n14766), .A(n14765), .ZN(n14767) );
  AOI21_X1 U16632 ( .B1(n14768), .B2(n15340), .A(n14767), .ZN(n14775) );
  MUX2_X1 U16633 ( .A(n10609), .B(P1_REG2_REG_11__SCAN_IN), .S(n14768), .Z(
        n14769) );
  NAND3_X1 U16634 ( .A1(n14771), .A2(n14770), .A3(n14769), .ZN(n14772) );
  NAND3_X1 U16635 ( .A1(n15338), .A2(n14773), .A3(n14772), .ZN(n14774) );
  NAND3_X1 U16636 ( .A1(n14776), .A2(n14775), .A3(n14774), .ZN(P1_U3254) );
  NAND2_X1 U16637 ( .A1(n14781), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14777) );
  XNOR2_X1 U16638 ( .A(n14797), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n14791) );
  NAND2_X1 U16639 ( .A1(n14780), .A2(n14779), .ZN(n14783) );
  NAND2_X1 U16640 ( .A1(n14781), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U16641 ( .A1(n14783), .A2(n14782), .ZN(n14793) );
  XNOR2_X1 U16642 ( .A(n14793), .B(n14787), .ZN(n14792) );
  XOR2_X1 U16643 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14792), .Z(n14784) );
  NAND2_X1 U16644 ( .A1(n15332), .A2(n14784), .ZN(n14785) );
  NAND2_X1 U16645 ( .A1(n14786), .A2(n14785), .ZN(n14789) );
  NOR2_X1 U16646 ( .A1(n14804), .A2(n14787), .ZN(n14788) );
  AOI211_X1 U16647 ( .C1(n15342), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n14789), 
        .B(n14788), .ZN(n14790) );
  OAI21_X1 U16648 ( .B1(n14791), .B2(n14805), .A(n14790), .ZN(P1_U3261) );
  NAND2_X1 U16649 ( .A1(n14792), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14795) );
  NAND2_X1 U16650 ( .A1(n14793), .A2(n14798), .ZN(n14794) );
  NAND2_X1 U16651 ( .A1(n14795), .A2(n14794), .ZN(n14796) );
  XNOR2_X1 U16652 ( .A(n14796), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14808) );
  INV_X1 U16653 ( .A(n14808), .ZN(n14803) );
  NAND2_X1 U16654 ( .A1(n14799), .A2(n14798), .ZN(n14800) );
  XNOR2_X1 U16655 ( .A(n14802), .B(n14801), .ZN(n14806) );
  AOI22_X1 U16656 ( .A1(n14803), .A2(n15332), .B1(n14806), .B2(n15338), .ZN(
        n14811) );
  OAI21_X1 U16657 ( .B1(n14806), .B2(n14805), .A(n14804), .ZN(n14807) );
  AOI21_X1 U16658 ( .B1(n14808), .B2(n15332), .A(n14807), .ZN(n14810) );
  MUX2_X1 U16659 ( .A(n14811), .B(n14810), .S(n14809), .Z(n14814) );
  INV_X1 U16660 ( .A(n14812), .ZN(n14813) );
  OAI211_X1 U16661 ( .C1(n7297), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        P1_U3262) );
  NOR2_X1 U16662 ( .A1(n15005), .A2(n14820), .ZN(n14823) );
  NAND2_X1 U16663 ( .A1(n14822), .A2(n14821), .ZN(n15066) );
  NOR2_X1 U16664 ( .A1(n15405), .A2(n15066), .ZN(n14828) );
  AOI211_X1 U16665 ( .C1(n15064), .C2(n14954), .A(n14823), .B(n14828), .ZN(
        n14824) );
  OAI21_X1 U16666 ( .B1(n15065), .B2(n14935), .A(n14824), .ZN(P1_U3263) );
  OAI211_X1 U16667 ( .C1(n14826), .C2(n15068), .A(n15377), .B(n14825), .ZN(
        n15067) );
  AND2_X1 U16668 ( .A1(n15405), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14827) );
  NOR2_X1 U16669 ( .A1(n14828), .A2(n14827), .ZN(n14831) );
  NAND2_X1 U16670 ( .A1(n14829), .A2(n14954), .ZN(n14830) );
  OAI211_X1 U16671 ( .C1(n15067), .C2(n14935), .A(n14831), .B(n14830), .ZN(
        P1_U3264) );
  INV_X1 U16672 ( .A(n15447), .ZN(n15461) );
  AND3_X1 U16673 ( .A1(n14852), .A2(n14834), .A3(n14833), .ZN(n14835) );
  OAI21_X1 U16674 ( .B1(n14836), .B2(n14835), .A(n15389), .ZN(n14839) );
  AOI22_X1 U16675 ( .A1(n14837), .A2(n15031), .B1(n15029), .B2(n14870), .ZN(
        n14838) );
  NOR2_X1 U16676 ( .A1(n15405), .A2(n14840), .ZN(n15401) );
  AOI21_X1 U16677 ( .B1(n14855), .B2(n15093), .A(n15397), .ZN(n14842) );
  NAND2_X1 U16678 ( .A1(n14842), .A2(n14841), .ZN(n15095) );
  OAI22_X1 U16679 ( .A1(n14844), .A2(n14985), .B1(n14843), .B2(n15005), .ZN(
        n14845) );
  AOI21_X1 U16680 ( .B1(n15093), .B2(n14954), .A(n14845), .ZN(n14846) );
  OAI21_X1 U16681 ( .B1(n15095), .B2(n14935), .A(n14846), .ZN(n14847) );
  AOI21_X1 U16682 ( .B1(n15096), .B2(n15401), .A(n14847), .ZN(n14848) );
  OAI21_X1 U16683 ( .B1(n15097), .B2(n15405), .A(n14848), .ZN(P1_U3266) );
  OAI21_X1 U16684 ( .B1(n14851), .B2(n14850), .A(n14849), .ZN(n15104) );
  OAI21_X1 U16685 ( .B1(n14854), .B2(n14853), .A(n14852), .ZN(n15102) );
  OAI211_X1 U16686 ( .C1(n14875), .C2(n15100), .A(n15377), .B(n14855), .ZN(
        n15099) );
  AOI22_X1 U16687 ( .A1(n14856), .A2(n15031), .B1(n15029), .B2(n14887), .ZN(
        n15098) );
  AOI22_X1 U16688 ( .A1(n14857), .A2(n15392), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15405), .ZN(n14858) );
  OAI21_X1 U16689 ( .B1(n15098), .B2(n15405), .A(n14858), .ZN(n14859) );
  AOI21_X1 U16690 ( .B1(n14860), .B2(n14954), .A(n14859), .ZN(n14861) );
  OAI21_X1 U16691 ( .B1(n15099), .B2(n14935), .A(n14861), .ZN(n14862) );
  AOI21_X1 U16692 ( .B1(n15102), .B2(n14983), .A(n14862), .ZN(n14863) );
  OAI21_X1 U16693 ( .B1(n15104), .B2(n15060), .A(n14863), .ZN(P1_U3267) );
  NAND2_X1 U16694 ( .A1(n14920), .A2(n14902), .ZN(n14864) );
  INV_X1 U16695 ( .A(n14865), .ZN(n14866) );
  XNOR2_X1 U16696 ( .A(n14868), .B(n7140), .ZN(n14869) );
  NAND2_X1 U16697 ( .A1(n14869), .A2(n15389), .ZN(n14872) );
  AOI22_X1 U16698 ( .A1(n14870), .A2(n15031), .B1(n15029), .B2(n14907), .ZN(
        n14871) );
  OAI22_X1 U16699 ( .A1(n14874), .A2(n14985), .B1(n15005), .B2(n14873), .ZN(
        n14878) );
  OAI21_X1 U16700 ( .B1(n6598), .B2(n15108), .A(n15377), .ZN(n14876) );
  OR2_X1 U16701 ( .A1(n14876), .A2(n14875), .ZN(n15106) );
  NOR2_X1 U16702 ( .A1(n15106), .A2(n14935), .ZN(n14877) );
  AOI211_X1 U16703 ( .C1(n14954), .C2(n14879), .A(n14878), .B(n14877), .ZN(
        n14882) );
  NAND3_X1 U16704 ( .A1(n7911), .A2(n15105), .A3(n15381), .ZN(n14881) );
  OAI211_X1 U16705 ( .C1(n6620), .C2(n15405), .A(n14882), .B(n14881), .ZN(
        P1_U3268) );
  XNOR2_X1 U16706 ( .A(n14883), .B(n14885), .ZN(n14891) );
  INV_X1 U16707 ( .A(n14891), .ZN(n15114) );
  INV_X1 U16708 ( .A(n15401), .ZN(n15009) );
  OAI211_X1 U16709 ( .C1(n14886), .C2(n14885), .A(n14884), .B(n15389), .ZN(
        n14893) );
  NAND2_X1 U16710 ( .A1(n14887), .A2(n15031), .ZN(n14888) );
  OAI21_X1 U16711 ( .B1(n14889), .B2(n14941), .A(n14888), .ZN(n14890) );
  AOI21_X1 U16712 ( .B1(n14891), .B2(n15461), .A(n14890), .ZN(n14892) );
  NAND2_X1 U16713 ( .A1(n14893), .A2(n14892), .ZN(n15116) );
  NAND2_X1 U16714 ( .A1(n15116), .A2(n15005), .ZN(n14901) );
  OAI22_X1 U16715 ( .A1(n15005), .A2(n14895), .B1(n14894), .B2(n14985), .ZN(
        n14899) );
  NAND2_X1 U16716 ( .A1(n14912), .A2(n15111), .ZN(n14896) );
  NAND2_X1 U16717 ( .A1(n14896), .A2(n15377), .ZN(n14897) );
  OR2_X1 U16718 ( .A1(n6598), .A2(n14897), .ZN(n15112) );
  NOR2_X1 U16719 ( .A1(n15112), .A2(n14935), .ZN(n14898) );
  AOI211_X1 U16720 ( .C1(n14954), .C2(n15111), .A(n14899), .B(n14898), .ZN(
        n14900) );
  OAI211_X1 U16721 ( .C1(n15114), .C2(n15009), .A(n14901), .B(n14900), .ZN(
        P1_U3269) );
  NAND3_X1 U16722 ( .A1(n14920), .A2(n7307), .A3(n14902), .ZN(n14903) );
  NAND2_X1 U16723 ( .A1(n14904), .A2(n14903), .ZN(n14905) );
  NAND2_X1 U16724 ( .A1(n14905), .A2(n15389), .ZN(n14909) );
  NOR2_X1 U16725 ( .A1(n14944), .A2(n14941), .ZN(n14906) );
  AOI21_X1 U16726 ( .B1(n14907), .B2(n15031), .A(n14906), .ZN(n14908) );
  NAND2_X1 U16727 ( .A1(n14909), .A2(n14908), .ZN(n15126) );
  NAND2_X1 U16728 ( .A1(n14911), .A2(n14910), .ZN(n15119) );
  AND3_X1 U16729 ( .A1(n15120), .A2(n15381), .A3(n15119), .ZN(n14918) );
  AOI21_X1 U16730 ( .B1(n14928), .B2(n15121), .A(n15397), .ZN(n14913) );
  NAND2_X1 U16731 ( .A1(n14913), .A2(n14912), .ZN(n15122) );
  AOI22_X1 U16732 ( .A1(n15405), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14914), 
        .B2(n15392), .ZN(n14916) );
  NAND2_X1 U16733 ( .A1(n15121), .A2(n14954), .ZN(n14915) );
  OAI211_X1 U16734 ( .C1(n15122), .C2(n14935), .A(n14916), .B(n14915), .ZN(
        n14917) );
  AOI211_X1 U16735 ( .C1(n15126), .C2(n15005), .A(n14918), .B(n14917), .ZN(
        n14919) );
  INV_X1 U16736 ( .A(n14919), .ZN(P1_U3270) );
  INV_X1 U16737 ( .A(n14920), .ZN(n14921) );
  AOI21_X1 U16738 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n15133) );
  NOR2_X1 U16739 ( .A1(n14924), .A2(n14947), .ZN(n14949) );
  NOR2_X1 U16740 ( .A1(n14949), .A2(n14925), .ZN(n14927) );
  XNOR2_X1 U16741 ( .A(n14927), .B(n14926), .ZN(n15131) );
  OAI211_X1 U16742 ( .C1(n14950), .C2(n15129), .A(n15377), .B(n14928), .ZN(
        n15128) );
  NOR2_X1 U16743 ( .A1(n15005), .A2(n14929), .ZN(n14933) );
  AOI22_X1 U16744 ( .A1(n14930), .A2(n15031), .B1(n15029), .B2(n14964), .ZN(
        n15127) );
  OAI22_X1 U16745 ( .A1(n15127), .A2(n15405), .B1(n14931), .B2(n14985), .ZN(
        n14932) );
  AOI211_X1 U16746 ( .C1(n7662), .C2(n14954), .A(n14933), .B(n14932), .ZN(
        n14934) );
  OAI21_X1 U16747 ( .B1(n15128), .B2(n14935), .A(n14934), .ZN(n14936) );
  AOI21_X1 U16748 ( .B1(n15131), .B2(n15381), .A(n14936), .ZN(n14937) );
  OAI21_X1 U16749 ( .B1(n15133), .B2(n14938), .A(n14937), .ZN(P1_U3271) );
  INV_X1 U16750 ( .A(n14947), .ZN(n14939) );
  XNOR2_X1 U16751 ( .A(n14940), .B(n14939), .ZN(n14946) );
  OAI22_X1 U16752 ( .A1(n14944), .A2(n14943), .B1(n14942), .B2(n14941), .ZN(
        n14945) );
  AOI21_X1 U16753 ( .B1(n14946), .B2(n15389), .A(n14945), .ZN(n15139) );
  AND2_X1 U16754 ( .A1(n14924), .A2(n14947), .ZN(n14948) );
  OR2_X1 U16755 ( .A1(n14949), .A2(n14948), .ZN(n15137) );
  OAI21_X1 U16756 ( .B1(n14966), .B2(n15135), .A(n15377), .ZN(n14951) );
  OR2_X1 U16757 ( .A1(n14951), .A2(n14950), .ZN(n15134) );
  INV_X1 U16758 ( .A(n14952), .ZN(n14953) );
  AOI22_X1 U16759 ( .A1(n15405), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14953), 
        .B2(n15392), .ZN(n14957) );
  NAND2_X1 U16760 ( .A1(n14955), .A2(n14954), .ZN(n14956) );
  OAI211_X1 U16761 ( .C1(n15134), .C2(n14962), .A(n14957), .B(n14956), .ZN(
        n14958) );
  AOI21_X1 U16762 ( .B1(n15137), .B2(n15381), .A(n14958), .ZN(n14959) );
  OAI21_X1 U16763 ( .B1(n15139), .B2(n15405), .A(n14959), .ZN(P1_U3272) );
  OAI211_X1 U16764 ( .C1(n6562), .C2(n14961), .A(n15389), .B(n14960), .ZN(
        n15145) );
  INV_X1 U16765 ( .A(n14962), .ZN(n14976) );
  INV_X1 U16766 ( .A(n14963), .ZN(n14984) );
  OAI21_X1 U16767 ( .B1(n14984), .B2(n14971), .A(n15377), .ZN(n14967) );
  AOI22_X1 U16768 ( .A1(n14964), .A2(n15031), .B1(n15029), .B2(n14993), .ZN(
        n14965) );
  OAI21_X1 U16769 ( .B1(n14967), .B2(n14966), .A(n14965), .ZN(n15142) );
  INV_X1 U16770 ( .A(n14968), .ZN(n14969) );
  AOI22_X1 U16771 ( .A1(n15405), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14969), 
        .B2(n15392), .ZN(n14970) );
  OAI21_X1 U16772 ( .B1(n14971), .B2(n15394), .A(n14970), .ZN(n14975) );
  OAI21_X1 U16773 ( .B1(n6618), .B2(n14973), .A(n14972), .ZN(n15146) );
  NOR2_X1 U16774 ( .A1(n15146), .A2(n15060), .ZN(n14974) );
  AOI211_X1 U16775 ( .C1(n14976), .C2(n15142), .A(n14975), .B(n14974), .ZN(
        n14977) );
  OAI21_X1 U16776 ( .B1(n15405), .B2(n15145), .A(n14977), .ZN(P1_U3273) );
  NAND2_X1 U16777 ( .A1(n14979), .A2(n14978), .ZN(n14980) );
  XOR2_X1 U16778 ( .A(n14981), .B(n14980), .Z(n15153) );
  XNOR2_X1 U16779 ( .A(n14982), .B(n14981), .ZN(n15147) );
  NAND2_X1 U16780 ( .A1(n15147), .A2(n14983), .ZN(n14992) );
  AOI211_X1 U16781 ( .C1(n15150), .C2(n15002), .A(n15397), .B(n14984), .ZN(
        n15148) );
  INV_X1 U16782 ( .A(n15149), .ZN(n14987) );
  OAI22_X1 U16783 ( .A1(n15405), .A2(n14987), .B1(n14986), .B2(n14985), .ZN(
        n14988) );
  AOI21_X1 U16784 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(n15405), .A(n14988), 
        .ZN(n14989) );
  OAI21_X1 U16785 ( .B1(n7119), .B2(n15394), .A(n14989), .ZN(n14990) );
  AOI21_X1 U16786 ( .B1(n15148), .B2(n15400), .A(n14990), .ZN(n14991) );
  OAI211_X1 U16787 ( .C1(n15153), .C2(n15060), .A(n14992), .B(n14991), .ZN(
        P1_U3274) );
  AND2_X1 U16788 ( .A1(n14993), .A2(n15031), .ZN(n15155) );
  XNOR2_X1 U16789 ( .A(n14994), .B(n14995), .ZN(n15008) );
  XNOR2_X1 U16790 ( .A(n14997), .B(n14996), .ZN(n14998) );
  AOI222_X1 U16791 ( .A1(n15008), .A2(n15461), .B1(n15032), .B2(n15029), .C1(
        n15389), .C2(n14998), .ZN(n15158) );
  INV_X1 U16792 ( .A(n15158), .ZN(n14999) );
  AOI211_X1 U16793 ( .C1(n15392), .C2(n15000), .A(n15155), .B(n14999), .ZN(
        n15013) );
  INV_X1 U16794 ( .A(n15001), .ZN(n15004) );
  INV_X1 U16795 ( .A(n15002), .ZN(n15003) );
  AOI211_X1 U16796 ( .C1(n15156), .C2(n15004), .A(n15397), .B(n15003), .ZN(
        n15154) );
  INV_X1 U16797 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15006) );
  OAI22_X1 U16798 ( .A1(n15007), .A2(n15394), .B1(n15006), .B2(n15005), .ZN(
        n15011) );
  INV_X1 U16799 ( .A(n15008), .ZN(n15159) );
  NOR2_X1 U16800 ( .A1(n15159), .A2(n15009), .ZN(n15010) );
  AOI211_X1 U16801 ( .C1(n15154), .C2(n15400), .A(n15011), .B(n15010), .ZN(
        n15012) );
  OAI21_X1 U16802 ( .B1(n15013), .B2(n15405), .A(n15012), .ZN(P1_U3275) );
  XNOR2_X1 U16803 ( .A(n15014), .B(n15023), .ZN(n15017) );
  AOI222_X1 U16804 ( .A1(n15389), .A2(n15017), .B1(n15016), .B2(n15029), .C1(
        n15015), .C2(n15031), .ZN(n15163) );
  XNOR2_X1 U16805 ( .A(n15034), .B(n15161), .ZN(n15018) );
  NOR2_X1 U16806 ( .A1(n15018), .A2(n15397), .ZN(n15160) );
  INV_X1 U16807 ( .A(n15019), .ZN(n15020) );
  AOI22_X1 U16808 ( .A1(n15405), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15020), 
        .B2(n15392), .ZN(n15021) );
  OAI21_X1 U16809 ( .B1(n15022), .B2(n15394), .A(n15021), .ZN(n15026) );
  XNOR2_X1 U16810 ( .A(n15024), .B(n15023), .ZN(n15164) );
  NOR2_X1 U16811 ( .A1(n15164), .A2(n15060), .ZN(n15025) );
  AOI211_X1 U16812 ( .C1(n15160), .C2(n15400), .A(n15026), .B(n15025), .ZN(
        n15027) );
  OAI21_X1 U16813 ( .B1(n15163), .B2(n15405), .A(n15027), .ZN(P1_U3276) );
  XNOR2_X1 U16814 ( .A(n15028), .B(n15039), .ZN(n15033) );
  AOI222_X1 U16815 ( .A1(n15389), .A2(n15033), .B1(n15032), .B2(n15031), .C1(
        n15030), .C2(n15029), .ZN(n15168) );
  INV_X1 U16816 ( .A(n15034), .ZN(n15035) );
  AOI211_X1 U16817 ( .C1(n15166), .C2(n15049), .A(n15397), .B(n15035), .ZN(
        n15165) );
  INV_X1 U16818 ( .A(n15036), .ZN(n15037) );
  AOI22_X1 U16819 ( .A1(n15405), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n15037), 
        .B2(n15392), .ZN(n15038) );
  OAI21_X1 U16820 ( .B1(n7663), .B2(n15394), .A(n15038), .ZN(n15042) );
  XOR2_X1 U16821 ( .A(n15040), .B(n15039), .Z(n15169) );
  NOR2_X1 U16822 ( .A1(n15169), .A2(n15060), .ZN(n15041) );
  AOI211_X1 U16823 ( .C1(n15165), .C2(n15400), .A(n15042), .B(n15041), .ZN(
        n15043) );
  OAI21_X1 U16824 ( .B1(n15168), .B2(n15405), .A(n15043), .ZN(P1_U3277) );
  OAI211_X1 U16825 ( .C1(n15046), .C2(n15045), .A(n15044), .B(n15389), .ZN(
        n15048) );
  AND2_X1 U16826 ( .A1(n15048), .A2(n15047), .ZN(n15173) );
  INV_X1 U16827 ( .A(n15049), .ZN(n15050) );
  AOI211_X1 U16828 ( .C1(n15171), .C2(n15051), .A(n15397), .B(n15050), .ZN(
        n15170) );
  AOI22_X1 U16829 ( .A1(n15405), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n15052), 
        .B2(n15392), .ZN(n15053) );
  OAI21_X1 U16830 ( .B1(n15054), .B2(n15394), .A(n15053), .ZN(n15062) );
  AOI21_X1 U16831 ( .B1(n12939), .B2(n15056), .A(n15055), .ZN(n15059) );
  INV_X1 U16832 ( .A(n15057), .ZN(n15058) );
  NOR2_X1 U16833 ( .A1(n15059), .A2(n15058), .ZN(n15174) );
  NOR2_X1 U16834 ( .A1(n15174), .A2(n15060), .ZN(n15061) );
  AOI211_X1 U16835 ( .C1(n15170), .C2(n15400), .A(n15062), .B(n15061), .ZN(
        n15063) );
  OAI21_X1 U16836 ( .B1(n15405), .B2(n15173), .A(n15063), .ZN(P1_U3278) );
  OAI211_X1 U16837 ( .C1(n14818), .C2(n15471), .A(n15065), .B(n15066), .ZN(
        n15192) );
  MUX2_X1 U16838 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15192), .S(n15492), .Z(
        P1_U3559) );
  OAI211_X1 U16839 ( .C1(n15068), .C2(n15471), .A(n15067), .B(n15066), .ZN(
        n15193) );
  MUX2_X1 U16840 ( .A(n15193), .B(P1_REG1_REG_30__SCAN_IN), .S(n7301), .Z(
        P1_U3558) );
  OAI211_X1 U16841 ( .C1(n15071), .C2(n15471), .A(n15070), .B(n15069), .ZN(
        n15072) );
  NOR2_X1 U16842 ( .A1(n15077), .A2(n15076), .ZN(n15084) );
  NAND2_X1 U16843 ( .A1(n15080), .A2(n15081), .ZN(n15078) );
  OAI211_X1 U16844 ( .C1(n15080), .C2(n15079), .A(n15078), .B(n15389), .ZN(
        n15082) );
  NAND2_X1 U16845 ( .A1(n15087), .A2(n15189), .ZN(n15088) );
  MUX2_X1 U16846 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15194), .S(n15492), .Z(
        P1_U3556) );
  INV_X1 U16847 ( .A(n15446), .ZN(n15468) );
  NAND2_X1 U16848 ( .A1(n15093), .A2(n15189), .ZN(n15094) );
  MUX2_X1 U16849 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15195), .S(n15492), .Z(
        P1_U3555) );
  OAI211_X1 U16850 ( .C1(n15100), .C2(n15471), .A(n15099), .B(n15098), .ZN(
        n15101) );
  AOI21_X1 U16851 ( .B1(n15102), .B2(n15389), .A(n15101), .ZN(n15103) );
  OAI21_X1 U16852 ( .B1(n15104), .B2(n15456), .A(n15103), .ZN(n15196) );
  MUX2_X1 U16853 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15196), .S(n15492), .Z(
        P1_U3554) );
  INV_X1 U16854 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15110) );
  NAND3_X1 U16855 ( .A1(n7911), .A2(n15105), .A3(n15476), .ZN(n15107) );
  OAI211_X1 U16856 ( .C1(n15108), .C2(n15471), .A(n15107), .B(n15106), .ZN(
        n15109) );
  INV_X1 U16857 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n15117) );
  NAND2_X1 U16858 ( .A1(n15111), .A2(n15189), .ZN(n15113) );
  OAI211_X1 U16859 ( .C1(n15114), .C2(n15446), .A(n15113), .B(n15112), .ZN(
        n15115) );
  NOR2_X1 U16860 ( .A1(n15116), .A2(n15115), .ZN(n15200) );
  MUX2_X1 U16861 ( .A(n15117), .B(n15200), .S(n15492), .Z(n15118) );
  INV_X1 U16862 ( .A(n15118), .ZN(P1_U3552) );
  NAND3_X1 U16863 ( .A1(n15120), .A2(n15119), .A3(n15476), .ZN(n15124) );
  NAND2_X1 U16864 ( .A1(n15121), .A2(n15189), .ZN(n15123) );
  NAND3_X1 U16865 ( .A1(n15124), .A2(n15123), .A3(n15122), .ZN(n15125) );
  MUX2_X1 U16866 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15203), .S(n15492), .Z(
        P1_U3551) );
  OAI211_X1 U16867 ( .C1(n15129), .C2(n15471), .A(n15128), .B(n15127), .ZN(
        n15130) );
  AOI21_X1 U16868 ( .B1(n15131), .B2(n15476), .A(n15130), .ZN(n15132) );
  OAI21_X1 U16869 ( .B1(n15133), .B2(n15355), .A(n15132), .ZN(n15204) );
  MUX2_X1 U16870 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15204), .S(n15492), .Z(
        P1_U3550) );
  INV_X1 U16871 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n15140) );
  OAI21_X1 U16872 ( .B1(n15135), .B2(n15471), .A(n15134), .ZN(n15136) );
  AOI21_X1 U16873 ( .B1(n15137), .B2(n15476), .A(n15136), .ZN(n15138) );
  AND2_X1 U16874 ( .A1(n15139), .A2(n15138), .ZN(n15205) );
  MUX2_X1 U16875 ( .A(n15140), .B(n15205), .S(n15492), .Z(n15141) );
  INV_X1 U16876 ( .A(n15141), .ZN(P1_U3549) );
  AOI21_X1 U16877 ( .B1(n15189), .B2(n15143), .A(n15142), .ZN(n15144) );
  OAI211_X1 U16878 ( .C1(n15456), .C2(n15146), .A(n15145), .B(n15144), .ZN(
        n15207) );
  MUX2_X1 U16879 ( .A(n15207), .B(P1_REG1_REG_20__SCAN_IN), .S(n7301), .Z(
        P1_U3548) );
  NAND2_X1 U16880 ( .A1(n15147), .A2(n15389), .ZN(n15152) );
  AOI211_X1 U16881 ( .C1(n15189), .C2(n15150), .A(n15149), .B(n15148), .ZN(
        n15151) );
  OAI211_X1 U16882 ( .C1(n15153), .C2(n15456), .A(n15152), .B(n15151), .ZN(
        n15208) );
  MUX2_X1 U16883 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15208), .S(n15492), .Z(
        P1_U3547) );
  AOI211_X1 U16884 ( .C1(n15189), .C2(n15156), .A(n15155), .B(n15154), .ZN(
        n15157) );
  OAI211_X1 U16885 ( .C1(n15159), .C2(n15446), .A(n15158), .B(n15157), .ZN(
        n15209) );
  MUX2_X1 U16886 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15209), .S(n15492), .Z(
        P1_U3546) );
  AOI21_X1 U16887 ( .B1(n15189), .B2(n15161), .A(n15160), .ZN(n15162) );
  OAI211_X1 U16888 ( .C1(n15456), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        n15210) );
  MUX2_X1 U16889 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15210), .S(n15492), .Z(
        P1_U3545) );
  AOI21_X1 U16890 ( .B1(n15189), .B2(n15166), .A(n15165), .ZN(n15167) );
  OAI211_X1 U16891 ( .C1(n15456), .C2(n15169), .A(n15168), .B(n15167), .ZN(
        n15211) );
  MUX2_X1 U16892 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15211), .S(n15492), .Z(
        P1_U3544) );
  AOI21_X1 U16893 ( .B1(n15189), .B2(n15171), .A(n15170), .ZN(n15172) );
  OAI211_X1 U16894 ( .C1(n15456), .C2(n15174), .A(n15173), .B(n15172), .ZN(
        n15212) );
  MUX2_X1 U16895 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15212), .S(n15492), .Z(
        P1_U3543) );
  NAND2_X1 U16896 ( .A1(n15175), .A2(n15189), .ZN(n15179) );
  NAND3_X1 U16897 ( .A1(n12939), .A2(n15176), .A3(n15476), .ZN(n15178) );
  NAND4_X1 U16898 ( .A1(n15180), .A2(n15179), .A3(n15178), .A4(n15177), .ZN(
        n15213) );
  MUX2_X1 U16899 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15213), .S(n15492), .Z(
        P1_U3542) );
  AOI211_X1 U16900 ( .C1(n15189), .C2(n15183), .A(n15182), .B(n15181), .ZN(
        n15184) );
  OAI21_X1 U16901 ( .B1(n15456), .B2(n15185), .A(n15184), .ZN(n15214) );
  MUX2_X1 U16902 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15214), .S(n15492), .Z(
        P1_U3541) );
  AOI211_X1 U16903 ( .C1(n15189), .C2(n15188), .A(n15187), .B(n15186), .ZN(
        n15190) );
  OAI21_X1 U16904 ( .B1(n15456), .B2(n15191), .A(n15190), .ZN(n15215) );
  MUX2_X1 U16905 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15215), .S(n15492), .Z(
        P1_U3540) );
  MUX2_X1 U16906 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15192), .S(n15478), .Z(
        P1_U3527) );
  MUX2_X1 U16907 ( .A(n15193), .B(P1_REG0_REG_30__SCAN_IN), .S(n15477), .Z(
        P1_U3526) );
  MUX2_X1 U16908 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15196), .S(n15478), .Z(
        P1_U3522) );
  INV_X1 U16909 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n15198) );
  INV_X1 U16910 ( .A(n15199), .ZN(P1_U3521) );
  INV_X1 U16911 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15201) );
  MUX2_X1 U16912 ( .A(n15201), .B(n15200), .S(n15478), .Z(n15202) );
  INV_X1 U16913 ( .A(n15202), .ZN(P1_U3520) );
  MUX2_X1 U16914 ( .A(n15203), .B(P1_REG0_REG_23__SCAN_IN), .S(n15477), .Z(
        P1_U3519) );
  MUX2_X1 U16915 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15204), .S(n15478), .Z(
        P1_U3518) );
  MUX2_X1 U16916 ( .A(n15718), .B(n15205), .S(n15478), .Z(n15206) );
  INV_X1 U16917 ( .A(n15206), .ZN(P1_U3517) );
  MUX2_X1 U16918 ( .A(n15207), .B(P1_REG0_REG_20__SCAN_IN), .S(n15477), .Z(
        P1_U3516) );
  MUX2_X1 U16919 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15208), .S(n15478), .Z(
        P1_U3515) );
  MUX2_X1 U16920 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15209), .S(n15478), .Z(
        P1_U3513) );
  MUX2_X1 U16921 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15210), .S(n15478), .Z(
        P1_U3510) );
  MUX2_X1 U16922 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15211), .S(n15478), .Z(
        P1_U3507) );
  MUX2_X1 U16923 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15212), .S(n15478), .Z(
        P1_U3504) );
  MUX2_X1 U16924 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15213), .S(n15478), .Z(
        P1_U3501) );
  MUX2_X1 U16925 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15214), .S(n15478), .Z(
        P1_U3498) );
  MUX2_X1 U16926 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15215), .S(n15478), .Z(
        P1_U3495) );
  INV_X1 U16927 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n15216) );
  NAND3_X1 U16928 ( .A1(n15216), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n15218) );
  OAI22_X1 U16929 ( .A1(n15219), .A2(n15218), .B1(n15217), .B2(n15232), .ZN(
        n15220) );
  AOI21_X1 U16930 ( .B1(n12715), .B2(n15221), .A(n15220), .ZN(n15222) );
  INV_X1 U16931 ( .A(n15222), .ZN(P1_U3324) );
  OAI222_X1 U16932 ( .A1(n15236), .A2(n15225), .B1(n15224), .B2(P1_U3086), 
        .C1(n15223), .C2(n15232), .ZN(P1_U3325) );
  OAI222_X1 U16933 ( .A1(n15236), .A2(n15228), .B1(n15227), .B2(n6537), .C1(
        n15226), .C2(n15232), .ZN(P1_U3326) );
  OAI222_X1 U16934 ( .A1(n15236), .A2(n15231), .B1(n15230), .B2(P1_U3086), 
        .C1(n15229), .C2(n15232), .ZN(P1_U3328) );
  OAI222_X1 U16935 ( .A1(n15236), .A2(n15235), .B1(n6537), .B2(n15234), .C1(
        n15233), .C2(n15232), .ZN(P1_U3329) );
  MUX2_X1 U16936 ( .A(n15238), .B(n15237), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16937 ( .A(n15239), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U16938 ( .A(n15240), .B(n15241), .Z(SUB_1596_U5) );
  XOR2_X1 U16939 ( .A(n15242), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U16940 ( .A(n15243), .B(n15244), .Z(SUB_1596_U59) );
  XOR2_X1 U16941 ( .A(n15246), .B(n15245), .Z(SUB_1596_U57) );
  XOR2_X1 U16942 ( .A(n15248), .B(n15247), .Z(SUB_1596_U56) );
  XOR2_X1 U16943 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n15249), .Z(SUB_1596_U70)
         );
  AND2_X1 U16944 ( .A1(n15253), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n15254) );
  OAI22_X1 U16945 ( .A1(n15255), .A2(n15254), .B1(P1_ADDR_REG_12__SCAN_IN), 
        .B2(n15253), .ZN(n15266) );
  INV_X1 U16946 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15256) );
  NAND2_X1 U16947 ( .A1(n15256), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n15267) );
  OAI21_X1 U16948 ( .B1(P3_ADDR_REG_13__SCAN_IN), .B2(n15256), .A(n15267), 
        .ZN(n15257) );
  XNOR2_X1 U16949 ( .A(n15266), .B(n15257), .ZN(n15258) );
  NAND2_X1 U16950 ( .A1(n15261), .A2(n15262), .ZN(n15260) );
  INV_X1 U16951 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15820) );
  XOR2_X1 U16952 ( .A(n15260), .B(n15820), .Z(SUB_1596_U67) );
  NAND2_X1 U16953 ( .A1(n15261), .A2(n15820), .ZN(n15263) );
  NAND2_X1 U16954 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15264), .ZN(n15265) );
  NAND2_X1 U16955 ( .A1(n15266), .A2(n15265), .ZN(n15268) );
  XNOR2_X1 U16956 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n15269) );
  XNOR2_X1 U16957 ( .A(n15279), .B(n15269), .ZN(n15271) );
  INV_X1 U16958 ( .A(n15271), .ZN(n15272) );
  NAND2_X1 U16959 ( .A1(n15275), .A2(n15276), .ZN(n15273) );
  XNOR2_X1 U16960 ( .A(n15273), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AND2_X1 U16961 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n15277), .ZN(n15278) );
  INV_X1 U16962 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15942) );
  NAND2_X1 U16963 ( .A1(n15942), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n15280) );
  INV_X1 U16964 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15281) );
  NAND2_X1 U16965 ( .A1(n15281), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n15290) );
  NAND2_X1 U16966 ( .A1(n11332), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n15282) );
  AND2_X1 U16967 ( .A1(n15290), .A2(n15282), .ZN(n15288) );
  INV_X1 U16968 ( .A(n15288), .ZN(n15283) );
  XNOR2_X1 U16969 ( .A(n15289), .B(n15283), .ZN(n15284) );
  NAND2_X1 U16970 ( .A1(n15286), .A2(n15287), .ZN(n15285) );
  XNOR2_X1 U16971 ( .A(n15285), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  INV_X1 U16972 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15771) );
  NOR2_X1 U16973 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15771), .ZN(n15299) );
  AOI21_X1 U16974 ( .B1(n15771), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n15299), 
        .ZN(n15292) );
  XNOR2_X1 U16975 ( .A(n15301), .B(n15292), .ZN(n15293) );
  NAND2_X1 U16976 ( .A1(n15294), .A2(n15293), .ZN(n15297) );
  NAND2_X1 U16977 ( .A1(n15296), .A2(n15297), .ZN(n15295) );
  XNOR2_X1 U16978 ( .A(n15295), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  INV_X1 U16979 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15592) );
  INV_X1 U16980 ( .A(n15299), .ZN(n15300) );
  NAND2_X1 U16981 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15771), .ZN(n15302) );
  NAND2_X1 U16982 ( .A1(n6617), .A2(n15306), .ZN(n15305) );
  XNOR2_X1 U16983 ( .A(n15305), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  NAND2_X1 U16984 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15319), .ZN(n15307) );
  OAI21_X1 U16985 ( .B1(n15319), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n15307), 
        .ZN(n15318) );
  NOR2_X1 U16986 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15309), .ZN(n15310) );
  XOR2_X1 U16987 ( .A(n15318), .B(n15321), .Z(n15312) );
  AOI21_X1 U16988 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15313), .A(n15317), 
        .ZN(n15314) );
  INV_X1 U16989 ( .A(n15314), .ZN(SUB_1596_U62) );
  INV_X1 U16990 ( .A(n15315), .ZN(n15316) );
  INV_X1 U16991 ( .A(n15318), .ZN(n15320) );
  AOI22_X1 U16992 ( .A1(n15321), .A2(n15320), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n15319), .ZN(n15324) );
  XNOR2_X1 U16993 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15322) );
  XNOR2_X1 U16994 ( .A(n15322), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n15323) );
  XNOR2_X1 U16995 ( .A(n15324), .B(n15323), .ZN(n15325) );
  XNOR2_X1 U16996 ( .A(n6672), .B(n15325), .ZN(SUB_1596_U4) );
  AOI21_X1 U16997 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15326) );
  OAI21_X1 U16998 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15326), 
        .ZN(U28) );
  INV_X1 U16999 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15856) );
  OAI221_X1 U17000 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n7295), .C2(n7935), .A(n15856), .ZN(U29) );
  MUX2_X1 U17001 ( .A(n10631), .B(P1_REG1_REG_4__SCAN_IN), .S(n15339), .Z(
        n15327) );
  NAND3_X1 U17002 ( .A1(n15329), .A2(n15328), .A3(n15327), .ZN(n15330) );
  NAND3_X1 U17003 ( .A1(n15332), .A2(n15331), .A3(n15330), .ZN(n15346) );
  MUX2_X1 U17004 ( .A(n10591), .B(P1_REG2_REG_4__SCAN_IN), .S(n15339), .Z(
        n15333) );
  NAND3_X1 U17005 ( .A1(n15335), .A2(n15334), .A3(n15333), .ZN(n15336) );
  NAND3_X1 U17006 ( .A1(n15338), .A2(n15337), .A3(n15336), .ZN(n15345) );
  NAND2_X1 U17007 ( .A1(n15340), .A2(n15339), .ZN(n15344) );
  AOI21_X1 U17008 ( .B1(n15342), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n15341), .ZN(
        n15343) );
  AND4_X1 U17009 ( .A1(n15346), .A2(n15345), .A3(n15344), .A4(n15343), .ZN(
        n15348) );
  NAND2_X1 U17010 ( .A1(n15348), .A2(n15347), .ZN(P1_U3247) );
  AND2_X1 U17011 ( .A1(n11681), .A2(n15351), .ZN(n15352) );
  XNOR2_X1 U17012 ( .A(n15352), .B(n7813), .ZN(n15444) );
  XNOR2_X1 U17013 ( .A(n15353), .B(n7813), .ZN(n15356) );
  OAI21_X1 U17014 ( .B1(n15356), .B2(n15355), .A(n15354), .ZN(n15357) );
  AOI21_X1 U17015 ( .B1(n15461), .B2(n15444), .A(n15357), .ZN(n15441) );
  AOI22_X1 U17016 ( .A1(n15405), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n15358), 
        .B2(n15392), .ZN(n15359) );
  OAI21_X1 U17017 ( .B1(n15394), .B2(n15440), .A(n15359), .ZN(n15360) );
  INV_X1 U17018 ( .A(n15360), .ZN(n15366) );
  INV_X1 U17019 ( .A(n15361), .ZN(n15363) );
  OAI211_X1 U17020 ( .C1(n15363), .C2(n15440), .A(n15377), .B(n15362), .ZN(
        n15439) );
  INV_X1 U17021 ( .A(n15439), .ZN(n15364) );
  AOI22_X1 U17022 ( .A1(n15444), .A2(n15401), .B1(n15400), .B2(n15364), .ZN(
        n15365) );
  OAI211_X1 U17023 ( .C1(n15405), .C2(n15441), .A(n15366), .B(n15365), .ZN(
        P1_U3287) );
  XNOR2_X1 U17024 ( .A(n15368), .B(n15367), .ZN(n15370) );
  AOI21_X1 U17025 ( .B1(n15370), .B2(n15389), .A(n15369), .ZN(n15428) );
  AOI22_X1 U17026 ( .A1(n15405), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n15371), 
        .B2(n15392), .ZN(n15372) );
  OAI21_X1 U17027 ( .B1(n15394), .B2(n15427), .A(n15372), .ZN(n15373) );
  INV_X1 U17028 ( .A(n15373), .ZN(n15383) );
  XNOR2_X1 U17029 ( .A(n15374), .B(n7247), .ZN(n15431) );
  INV_X1 U17030 ( .A(n15375), .ZN(n15379) );
  INV_X1 U17031 ( .A(n15376), .ZN(n15378) );
  OAI211_X1 U17032 ( .C1(n15427), .C2(n15379), .A(n15378), .B(n15377), .ZN(
        n15426) );
  INV_X1 U17033 ( .A(n15426), .ZN(n15380) );
  AOI22_X1 U17034 ( .A1(n15381), .A2(n15431), .B1(n15400), .B2(n15380), .ZN(
        n15382) );
  OAI211_X1 U17035 ( .C1(n15405), .C2(n15428), .A(n15383), .B(n15382), .ZN(
        P1_U3289) );
  XNOR2_X1 U17036 ( .A(n15384), .B(n15385), .ZN(n15420) );
  XNOR2_X1 U17037 ( .A(n15387), .B(n15386), .ZN(n15390) );
  AOI21_X1 U17038 ( .B1(n15390), .B2(n15389), .A(n15388), .ZN(n15417) );
  INV_X1 U17039 ( .A(n15417), .ZN(n15391) );
  AOI21_X1 U17040 ( .B1(n15461), .B2(n15420), .A(n15391), .ZN(n15404) );
  AOI22_X1 U17041 ( .A1(n15405), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n15392), .ZN(n15393) );
  OAI21_X1 U17042 ( .B1(n15394), .B2(n15418), .A(n15393), .ZN(n15395) );
  INV_X1 U17043 ( .A(n15395), .ZN(n15403) );
  AOI211_X1 U17044 ( .C1(n15399), .C2(n15398), .A(n15397), .B(n15396), .ZN(
        n15415) );
  AOI22_X1 U17045 ( .A1(n15401), .A2(n15420), .B1(n15400), .B2(n15415), .ZN(
        n15402) );
  OAI211_X1 U17046 ( .C1(n15405), .C2(n15404), .A(n15403), .B(n15402), .ZN(
        P1_U3291) );
  AND2_X1 U17047 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15407), .ZN(P1_U3294) );
  INV_X1 U17048 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15815) );
  NOR2_X1 U17049 ( .A1(n15406), .A2(n15815), .ZN(P1_U3295) );
  AND2_X1 U17050 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15407), .ZN(P1_U3296) );
  AND2_X1 U17051 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15407), .ZN(P1_U3297) );
  INV_X1 U17052 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15854) );
  NOR2_X1 U17053 ( .A1(n15406), .A2(n15854), .ZN(P1_U3298) );
  AND2_X1 U17054 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15407), .ZN(P1_U3299) );
  AND2_X1 U17055 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15407), .ZN(P1_U3300) );
  AND2_X1 U17056 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15407), .ZN(P1_U3301) );
  AND2_X1 U17057 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15407), .ZN(P1_U3302) );
  INV_X1 U17058 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15769) );
  NOR2_X1 U17059 ( .A1(n15406), .A2(n15769), .ZN(P1_U3303) );
  AND2_X1 U17060 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15407), .ZN(P1_U3304) );
  AND2_X1 U17061 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15407), .ZN(P1_U3305) );
  NOR2_X1 U17062 ( .A1(n15406), .A2(n15964), .ZN(P1_U3306) );
  AND2_X1 U17063 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15407), .ZN(P1_U3307) );
  AND2_X1 U17064 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15407), .ZN(P1_U3308) );
  AND2_X1 U17065 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15407), .ZN(P1_U3309) );
  AND2_X1 U17066 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15407), .ZN(P1_U3310) );
  AND2_X1 U17067 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15407), .ZN(P1_U3311) );
  NOR2_X1 U17068 ( .A1(n15406), .A2(n15760), .ZN(P1_U3312) );
  AND2_X1 U17069 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15407), .ZN(P1_U3313) );
  AND2_X1 U17070 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15407), .ZN(P1_U3314) );
  AND2_X1 U17071 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15407), .ZN(P1_U3315) );
  AND2_X1 U17072 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15407), .ZN(P1_U3316) );
  AND2_X1 U17073 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15407), .ZN(P1_U3317) );
  AND2_X1 U17074 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15407), .ZN(P1_U3318) );
  INV_X1 U17075 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15845) );
  NOR2_X1 U17076 ( .A1(n15406), .A2(n15845), .ZN(P1_U3319) );
  AND2_X1 U17077 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15407), .ZN(P1_U3320) );
  AND2_X1 U17078 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15407), .ZN(P1_U3321) );
  AND2_X1 U17079 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15407), .ZN(P1_U3322) );
  AND2_X1 U17080 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15407), .ZN(P1_U3323) );
  INV_X1 U17081 ( .A(n15408), .ZN(n15414) );
  OAI21_X1 U17082 ( .B1(n15410), .B2(n15471), .A(n15409), .ZN(n15413) );
  INV_X1 U17083 ( .A(n15411), .ZN(n15412) );
  AOI211_X1 U17084 ( .C1(n15476), .C2(n15414), .A(n15413), .B(n15412), .ZN(
        n15479) );
  AOI22_X1 U17085 ( .A1(n15478), .A2(n15479), .B1(n8863), .B2(n15477), .ZN(
        P1_U3462) );
  INV_X1 U17086 ( .A(n15415), .ZN(n15416) );
  OAI211_X1 U17087 ( .C1(n15418), .C2(n15471), .A(n15417), .B(n15416), .ZN(
        n15419) );
  AOI21_X1 U17088 ( .B1(n15420), .B2(n15476), .A(n15419), .ZN(n15480) );
  AOI22_X1 U17089 ( .A1(n15478), .A2(n15480), .B1(n15703), .B2(n15477), .ZN(
        P1_U3465) );
  AOI21_X1 U17090 ( .B1(n15447), .B2(n15446), .A(n15421), .ZN(n15425) );
  OAI21_X1 U17091 ( .B1(n11674), .B2(n15471), .A(n15422), .ZN(n15423) );
  NOR3_X1 U17092 ( .A1(n15425), .A2(n15424), .A3(n15423), .ZN(n15481) );
  AOI22_X1 U17093 ( .A1(n15478), .A2(n15481), .B1(n8895), .B2(n15477), .ZN(
        P1_U3468) );
  OAI21_X1 U17094 ( .B1(n15427), .B2(n15471), .A(n15426), .ZN(n15430) );
  INV_X1 U17095 ( .A(n15428), .ZN(n15429) );
  AOI211_X1 U17096 ( .C1(n15431), .C2(n15476), .A(n15430), .B(n15429), .ZN(
        n15482) );
  AOI22_X1 U17097 ( .A1(n15478), .A2(n15482), .B1(n8911), .B2(n15477), .ZN(
        P1_U3471) );
  OAI211_X1 U17098 ( .C1(n15434), .C2(n15471), .A(n15433), .B(n15432), .ZN(
        n15437) );
  AOI21_X1 U17099 ( .B1(n15447), .B2(n15446), .A(n15435), .ZN(n15436) );
  AOI211_X1 U17100 ( .C1(n15389), .C2(n15438), .A(n15437), .B(n15436), .ZN(
        n15484) );
  AOI22_X1 U17101 ( .A1(n15478), .A2(n15484), .B1(n8930), .B2(n15477), .ZN(
        P1_U3474) );
  OAI21_X1 U17102 ( .B1(n15440), .B2(n15471), .A(n15439), .ZN(n15443) );
  INV_X1 U17103 ( .A(n15441), .ZN(n15442) );
  AOI211_X1 U17104 ( .C1(n15468), .C2(n15444), .A(n15443), .B(n15442), .ZN(
        n15485) );
  AOI22_X1 U17105 ( .A1(n15478), .A2(n15485), .B1(n8948), .B2(n15477), .ZN(
        P1_U3477) );
  AOI21_X1 U17106 ( .B1(n15447), .B2(n15446), .A(n15445), .ZN(n15452) );
  INV_X1 U17107 ( .A(n15448), .ZN(n15450) );
  NOR4_X1 U17108 ( .A1(n15452), .A2(n15451), .A3(n15450), .A4(n15449), .ZN(
        n15486) );
  AOI22_X1 U17109 ( .A1(n15478), .A2(n15486), .B1(n8969), .B2(n15477), .ZN(
        P1_U3480) );
  INV_X1 U17110 ( .A(n15453), .ZN(n15454) );
  OAI211_X1 U17111 ( .C1(n15457), .C2(n15456), .A(n15455), .B(n15454), .ZN(
        n15460) );
  INV_X1 U17112 ( .A(n15458), .ZN(n15459) );
  NOR2_X1 U17113 ( .A1(n15460), .A2(n15459), .ZN(n15488) );
  AOI22_X1 U17114 ( .A1(n15478), .A2(n15488), .B1(n8992), .B2(n15477), .ZN(
        P1_U3483) );
  NAND2_X1 U17115 ( .A1(n15467), .A2(n15461), .ZN(n15462) );
  NAND4_X1 U17116 ( .A1(n15465), .A2(n15464), .A3(n15463), .A4(n15462), .ZN(
        n15466) );
  AOI21_X1 U17117 ( .B1(n15468), .B2(n15467), .A(n15466), .ZN(n15490) );
  AOI22_X1 U17118 ( .A1(n15478), .A2(n15490), .B1(n9012), .B2(n15477), .ZN(
        P1_U3486) );
  OAI211_X1 U17119 ( .C1(n15472), .C2(n15471), .A(n15470), .B(n15469), .ZN(
        n15474) );
  AOI211_X1 U17120 ( .C1(n15476), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        n15491) );
  AOI22_X1 U17121 ( .A1(n15478), .A2(n15491), .B1(n9026), .B2(n15477), .ZN(
        P1_U3489) );
  AOI22_X1 U17122 ( .A1(n15492), .A2(n15479), .B1(n10623), .B2(n7301), .ZN(
        P1_U3529) );
  AOI22_X1 U17123 ( .A1(n15492), .A2(n15480), .B1(n10626), .B2(n7301), .ZN(
        P1_U3530) );
  AOI22_X1 U17124 ( .A1(n15492), .A2(n15481), .B1(n10622), .B2(n7301), .ZN(
        P1_U3531) );
  AOI22_X1 U17125 ( .A1(n15492), .A2(n15482), .B1(n10631), .B2(n7301), .ZN(
        P1_U3532) );
  AOI22_X1 U17126 ( .A1(n15492), .A2(n15484), .B1(n15483), .B2(n7301), .ZN(
        P1_U3533) );
  AOI22_X1 U17127 ( .A1(n15492), .A2(n15485), .B1(n15756), .B2(n7301), .ZN(
        P1_U3534) );
  AOI22_X1 U17128 ( .A1(n15492), .A2(n15486), .B1(n10636), .B2(n7301), .ZN(
        P1_U3535) );
  AOI22_X1 U17129 ( .A1(n15492), .A2(n15488), .B1(n15487), .B2(n7301), .ZN(
        P1_U3536) );
  AOI22_X1 U17130 ( .A1(n15492), .A2(n15490), .B1(n15489), .B2(n7301), .ZN(
        P1_U3537) );
  AOI22_X1 U17131 ( .A1(n15492), .A2(n15491), .B1(n15943), .B2(n7301), .ZN(
        P1_U3538) );
  NOR2_X1 U17132 ( .A1(n15527), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U17133 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15603), .B1(n15596), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15496) );
  AOI22_X1 U17134 ( .A1(n15527), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15495) );
  OAI22_X1 U17135 ( .A1(n15586), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n15579), .ZN(n15493) );
  OAI21_X1 U17136 ( .B1(n15595), .B2(n15493), .A(n15497), .ZN(n15494) );
  OAI211_X1 U17137 ( .C1(n15497), .C2(n15496), .A(n15495), .B(n15494), .ZN(
        P2_U3214) );
  INV_X1 U17138 ( .A(n15498), .ZN(n15513) );
  OAI21_X1 U17139 ( .B1(n15513), .B2(n7840), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15499) );
  OAI21_X1 U17140 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_1__SCAN_IN), 
        .A(n15499), .ZN(n15511) );
  INV_X1 U17141 ( .A(n15500), .ZN(n15504) );
  OAI21_X1 U17142 ( .B1(n10487), .B2(n15502), .A(n15501), .ZN(n15503) );
  NAND3_X1 U17143 ( .A1(n15596), .A2(n15504), .A3(n15503), .ZN(n15510) );
  OAI211_X1 U17144 ( .C1(n15507), .C2(n15506), .A(n15603), .B(n15505), .ZN(
        n15509) );
  NAND2_X1 U17145 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15527), .ZN(n15508) );
  NAND4_X1 U17146 ( .A1(n15511), .A2(n15510), .A3(n15509), .A4(n15508), .ZN(
        P2_U3215) );
  OAI21_X1 U17147 ( .B1(n15513), .B2(n15512), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15514) );
  OAI21_X1 U17148 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_2__SCAN_IN), 
        .A(n15514), .ZN(n15524) );
  OAI211_X1 U17149 ( .C1(n15517), .C2(n15516), .A(n15603), .B(n15515), .ZN(
        n15523) );
  NAND2_X1 U17150 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n15527), .ZN(n15522) );
  AOI211_X1 U17151 ( .C1(n15519), .C2(n6606), .A(n15518), .B(n15586), .ZN(
        n15520) );
  INV_X1 U17152 ( .A(n15520), .ZN(n15521) );
  NAND4_X1 U17153 ( .A1(n15524), .A2(n15523), .A3(n15522), .A4(n15521), .ZN(
        P2_U3216) );
  OAI22_X1 U17154 ( .A1(n15584), .A2(n15525), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8069), .ZN(n15526) );
  AOI21_X1 U17155 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n15527), .A(n15526), .ZN(
        n15537) );
  AOI211_X1 U17156 ( .C1(n15530), .C2(n15529), .A(n15528), .B(n15586), .ZN(
        n15531) );
  INV_X1 U17157 ( .A(n15531), .ZN(n15536) );
  OAI211_X1 U17158 ( .C1(n15534), .C2(n15533), .A(n15603), .B(n15532), .ZN(
        n15535) );
  NAND3_X1 U17159 ( .A1(n15537), .A2(n15536), .A3(n15535), .ZN(P2_U3217) );
  INV_X1 U17160 ( .A(n15538), .ZN(n15542) );
  MUX2_X1 U17161 ( .A(n11870), .B(P2_REG2_REG_9__SCAN_IN), .S(n15539), .Z(
        n15541) );
  OAI21_X1 U17162 ( .B1(n15542), .B2(n15541), .A(n15540), .ZN(n15547) );
  XNOR2_X1 U17163 ( .A(n15544), .B(n15543), .ZN(n15545) );
  AOI222_X1 U17164 ( .A1(n15547), .A2(n15603), .B1(n15546), .B2(n15595), .C1(
        n15545), .C2(n15596), .ZN(n15549) );
  OAI211_X1 U17165 ( .C1(n15781), .C2(n15609), .A(n15549), .B(n15548), .ZN(
        P2_U3223) );
  INV_X1 U17166 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15551) );
  OAI21_X1 U17167 ( .B1(n15609), .B2(n15551), .A(n15550), .ZN(n15552) );
  AOI21_X1 U17168 ( .B1(n15553), .B2(n15595), .A(n15552), .ZN(n15563) );
  AOI211_X1 U17169 ( .C1(n15556), .C2(n15555), .A(n15586), .B(n15554), .ZN(
        n15557) );
  INV_X1 U17170 ( .A(n15557), .ZN(n15562) );
  OAI211_X1 U17171 ( .C1(n15560), .C2(n15559), .A(n15558), .B(n15603), .ZN(
        n15561) );
  NAND3_X1 U17172 ( .A1(n15563), .A2(n15562), .A3(n15561), .ZN(P2_U3224) );
  OAI21_X1 U17173 ( .B1(n15609), .B2(n15820), .A(n15564), .ZN(n15565) );
  AOI21_X1 U17174 ( .B1(n15566), .B2(n15595), .A(n15565), .ZN(n15577) );
  AOI21_X1 U17175 ( .B1(n15568), .B2(n15567), .A(n15579), .ZN(n15570) );
  NAND2_X1 U17176 ( .A1(n15570), .A2(n15569), .ZN(n15576) );
  AOI211_X1 U17177 ( .C1(n15573), .C2(n15572), .A(n15586), .B(n15571), .ZN(
        n15574) );
  INV_X1 U17178 ( .A(n15574), .ZN(n15575) );
  NAND3_X1 U17179 ( .A1(n15577), .A2(n15576), .A3(n15575), .ZN(P2_U3227) );
  INV_X1 U17180 ( .A(n15578), .ZN(n15581) );
  MUX2_X1 U17181 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n14237), .S(n15585), .Z(
        n15580) );
  AOI21_X1 U17182 ( .B1(n15581), .B2(n15580), .A(n15579), .ZN(n15589) );
  XNOR2_X1 U17183 ( .A(n15583), .B(n15582), .ZN(n15587) );
  OAI22_X1 U17184 ( .A1(n15587), .A2(n15586), .B1(n15585), .B2(n15584), .ZN(
        n15588) );
  AOI21_X1 U17185 ( .B1(n15589), .B2(n15601), .A(n15588), .ZN(n15591) );
  OAI211_X1 U17186 ( .C1(n15592), .C2(n15609), .A(n15591), .B(n15590), .ZN(
        P2_U3230) );
  XOR2_X1 U17187 ( .A(n15594), .B(n15593), .Z(n15597) );
  AOI22_X1 U17188 ( .A1(n15597), .A2(n15596), .B1(n15598), .B2(n15595), .ZN(
        n15606) );
  MUX2_X1 U17189 ( .A(n13989), .B(P2_REG2_REG_17__SCAN_IN), .S(n15598), .Z(
        n15599) );
  NAND3_X1 U17190 ( .A1(n15601), .A2(n15600), .A3(n15599), .ZN(n15602) );
  NAND3_X1 U17191 ( .A1(n15604), .A2(n15603), .A3(n15602), .ZN(n15605) );
  AND2_X1 U17192 ( .A1(n15606), .A2(n15605), .ZN(n15608) );
  OAI211_X1 U17193 ( .C1(n7504), .C2(n15609), .A(n15608), .B(n15607), .ZN(
        P2_U3231) );
  AND2_X1 U17194 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15611), .ZN(P2_U3266) );
  AND2_X1 U17195 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15611), .ZN(P2_U3267) );
  NOR2_X1 U17196 ( .A1(n15612), .A2(n15853), .ZN(P2_U3268) );
  AND2_X1 U17197 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15611), .ZN(P2_U3269) );
  AND2_X1 U17198 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15611), .ZN(P2_U3270) );
  AND2_X1 U17199 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15611), .ZN(P2_U3271) );
  AND2_X1 U17200 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15611), .ZN(P2_U3272) );
  AND2_X1 U17201 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15611), .ZN(P2_U3273) );
  AND2_X1 U17202 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15611), .ZN(P2_U3274) );
  AND2_X1 U17203 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15611), .ZN(P2_U3275) );
  AND2_X1 U17204 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15611), .ZN(P2_U3276) );
  AND2_X1 U17205 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15611), .ZN(P2_U3277) );
  AND2_X1 U17206 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15611), .ZN(P2_U3278) );
  INV_X1 U17207 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15898) );
  NOR2_X1 U17208 ( .A1(n15612), .A2(n15898), .ZN(P2_U3279) );
  INV_X1 U17209 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15872) );
  NOR2_X1 U17210 ( .A1(n15612), .A2(n15872), .ZN(P2_U3280) );
  NOR2_X1 U17211 ( .A1(n15612), .A2(n15842), .ZN(P2_U3281) );
  AND2_X1 U17212 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15611), .ZN(P2_U3282) );
  AND2_X1 U17213 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15611), .ZN(P2_U3283) );
  AND2_X1 U17214 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15611), .ZN(P2_U3284) );
  NOR2_X1 U17215 ( .A1(n15612), .A2(n15894), .ZN(P2_U3285) );
  AND2_X1 U17216 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15611), .ZN(P2_U3286) );
  AND2_X1 U17217 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15611), .ZN(P2_U3287) );
  AND2_X1 U17218 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15611), .ZN(P2_U3288) );
  NOR2_X1 U17219 ( .A1(n15612), .A2(n15923), .ZN(P2_U3289) );
  AND2_X1 U17220 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15611), .ZN(P2_U3290) );
  AND2_X1 U17221 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15611), .ZN(P2_U3291) );
  AND2_X1 U17222 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15611), .ZN(P2_U3292) );
  AND2_X1 U17223 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15611), .ZN(P2_U3293) );
  AND2_X1 U17224 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15611), .ZN(P2_U3294) );
  INV_X1 U17225 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15941) );
  NOR2_X1 U17226 ( .A1(n15612), .A2(n15941), .ZN(P2_U3295) );
  AOI22_X1 U17227 ( .A1(n15615), .A2(n15614), .B1(n15613), .B2(n15617), .ZN(
        P2_U3416) );
  AOI21_X1 U17228 ( .B1(n15618), .B2(n15617), .A(n15616), .ZN(P2_U3417) );
  OAI211_X1 U17229 ( .C1(n15621), .C2(n15636), .A(n15620), .B(n15619), .ZN(
        n15622) );
  INV_X1 U17230 ( .A(n15622), .ZN(n15660) );
  INV_X1 U17231 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15623) );
  AOI22_X1 U17232 ( .A1(n15659), .A2(n15660), .B1(n15623), .B2(n15657), .ZN(
        P2_U3430) );
  INV_X1 U17233 ( .A(n15624), .ZN(n15629) );
  OAI21_X1 U17234 ( .B1(n15626), .B2(n15640), .A(n15625), .ZN(n15628) );
  AOI211_X1 U17235 ( .C1(n15646), .C2(n15629), .A(n15628), .B(n15627), .ZN(
        n15662) );
  INV_X1 U17236 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15630) );
  AOI22_X1 U17237 ( .A1(n15659), .A2(n15662), .B1(n15630), .B2(n15657), .ZN(
        P2_U3436) );
  AOI21_X1 U17238 ( .B1(n15651), .B2(n15632), .A(n15631), .ZN(n15633) );
  OAI211_X1 U17239 ( .C1(n15636), .C2(n15635), .A(n15634), .B(n15633), .ZN(
        n15637) );
  INV_X1 U17240 ( .A(n15637), .ZN(n15664) );
  INV_X1 U17241 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15883) );
  AOI22_X1 U17242 ( .A1(n15659), .A2(n15664), .B1(n15883), .B2(n15657), .ZN(
        P2_U3442) );
  INV_X1 U17243 ( .A(n15643), .ZN(n15647) );
  OAI211_X1 U17244 ( .C1(n15641), .C2(n15640), .A(n15639), .B(n15638), .ZN(
        n15645) );
  NOR2_X1 U17245 ( .A1(n15643), .A2(n15642), .ZN(n15644) );
  AOI211_X1 U17246 ( .C1(n15647), .C2(n15646), .A(n15645), .B(n15644), .ZN(
        n15666) );
  INV_X1 U17247 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15648) );
  AOI22_X1 U17248 ( .A1(n15659), .A2(n15666), .B1(n15648), .B2(n15657), .ZN(
        P2_U3448) );
  AOI21_X1 U17249 ( .B1(n15651), .B2(n15650), .A(n15649), .ZN(n15652) );
  OAI211_X1 U17250 ( .C1(n15655), .C2(n15654), .A(n15653), .B(n15652), .ZN(
        n15656) );
  INV_X1 U17251 ( .A(n15656), .ZN(n15669) );
  INV_X1 U17252 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15658) );
  AOI22_X1 U17253 ( .A1(n15659), .A2(n15669), .B1(n15658), .B2(n15657), .ZN(
        P2_U3451) );
  AOI22_X1 U17254 ( .A1(n15670), .A2(n15660), .B1(n10487), .B2(n15667), .ZN(
        P2_U3499) );
  AOI22_X1 U17255 ( .A1(n15670), .A2(n15662), .B1(n15661), .B2(n15667), .ZN(
        P2_U3501) );
  AOI22_X1 U17256 ( .A1(n15670), .A2(n15664), .B1(n15663), .B2(n15667), .ZN(
        P2_U3503) );
  AOI22_X1 U17257 ( .A1(n15670), .A2(n15666), .B1(n15665), .B2(n15667), .ZN(
        P2_U3505) );
  AOI22_X1 U17258 ( .A1(n15670), .A2(n15669), .B1(n15668), .B2(n15667), .ZN(
        P2_U3506) );
  OAI22_X1 U17259 ( .A1(n15672), .A2(n15677), .B1(n15679), .B2(n15671), .ZN(
        n15673) );
  AOI211_X1 U17260 ( .C1(n15675), .C2(P3_REG3_REG_2__SCAN_IN), .A(n15674), .B(
        n15673), .ZN(n15676) );
  AOI22_X1 U17261 ( .A1(n15688), .A2(n6887), .B1(n15676), .B2(n13405), .ZN(
        P3_U3231) );
  NOR2_X1 U17262 ( .A1(n15678), .A2(n15677), .ZN(n15684) );
  OAI22_X1 U17263 ( .A1(n15682), .A2(n15681), .B1(n15680), .B2(n15679), .ZN(
        n15683) );
  NOR3_X1 U17264 ( .A1(n15685), .A2(n15684), .A3(n15683), .ZN(n15686) );
  AOI22_X1 U17265 ( .A1(n15688), .A2(n15687), .B1(n15686), .B2(n13405), .ZN(
        P3_U3232) );
  INV_X1 U17266 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15690) );
  AOI22_X1 U17267 ( .A1(n15693), .A2(n15690), .B1(n15689), .B2(n15691), .ZN(
        P3_U3393) );
  INV_X1 U17268 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15966) );
  AOI22_X1 U17269 ( .A1(n15693), .A2(n15966), .B1(n15692), .B2(n15691), .ZN(
        P3_U3396) );
  NOR2_X1 U17270 ( .A1(n15694), .A2(P3_U3897), .ZN(n15987) );
  NAND4_X1 U17271 ( .A1(n15696), .A2(n15695), .A3(P2_ADDR_REG_2__SCAN_IN), 
        .A4(P3_ADDR_REG_14__SCAN_IN), .ZN(n15701) );
  NAND4_X1 U17272 ( .A1(n15697), .A2(n9365), .A3(P3_IR_REG_20__SCAN_IN), .A4(
        P3_IR_REG_27__SCAN_IN), .ZN(n15700) );
  INV_X1 U17273 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n15929) );
  AND4_X1 U17274 ( .A1(P3_IR_REG_30__SCAN_IN), .A2(P3_REG2_REG_10__SCAN_IN), 
        .A3(n15927), .A4(n15922), .ZN(n15698) );
  NAND4_X1 U17275 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(n15943), .A3(n15929), .A4(
        n15698), .ZN(n15699) );
  NOR4_X1 U17276 ( .A1(n15701), .A2(n15700), .A3(n15699), .A4(n15941), .ZN(
        n15707) );
  NOR4_X1 U17277 ( .A1(n15702), .A2(n15925), .A3(n15944), .A4(
        P1_IR_REG_23__SCAN_IN), .ZN(n15706) );
  NOR4_X1 U17278 ( .A1(n15704), .A2(n15703), .A3(P3_ADDR_REG_7__SCAN_IN), .A4(
        P1_IR_REG_30__SCAN_IN), .ZN(n15705) );
  NAND3_X1 U17279 ( .A1(n15707), .A2(n15706), .A3(n15705), .ZN(n15708) );
  NOR4_X1 U17280 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(n15710), .A3(n15709), 
        .A4(n15708), .ZN(n15754) );
  NAND4_X1 U17281 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), 
        .A3(n15843), .A4(n7297), .ZN(n15715) );
  NAND4_X1 U17282 ( .A1(P3_REG1_REG_27__SCAN_IN), .A2(P3_ADDR_REG_8__SCAN_IN), 
        .A3(n15830), .A4(n15711), .ZN(n15714) );
  NAND4_X1 U17283 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(n15858), .ZN(n15713) );
  INV_X1 U17284 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n15839) );
  NAND4_X1 U17285 ( .A1(n15840), .A2(n15839), .A3(n12849), .A4(n15856), .ZN(
        n15712) );
  NOR4_X1 U17286 ( .A1(n15715), .A2(n15714), .A3(n15713), .A4(n15712), .ZN(
        n15753) );
  NAND4_X1 U17287 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P2_REG2_REG_16__SCAN_IN), 
        .A3(P3_DATAO_REG_16__SCAN_IN), .A4(n15820), .ZN(n15722) );
  NAND4_X1 U17288 ( .A1(P3_REG2_REG_28__SCAN_IN), .A2(P1_REG3_REG_9__SCAN_IN), 
        .A3(n15826), .A4(n15827), .ZN(n15716) );
  NOR3_X1 U17289 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(n15716), .A3(
        P1_REG2_REG_28__SCAN_IN), .ZN(n15719) );
  INV_X1 U17290 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n15717) );
  NAND3_X1 U17291 ( .A1(n15719), .A2(n15718), .A3(n15717), .ZN(n15721) );
  NAND4_X1 U17292 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(SI_11_), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P3_DATAO_REG_14__SCAN_IN), .ZN(n15720) );
  NOR3_X1 U17293 ( .A1(n15722), .A2(n15721), .A3(n15720), .ZN(n15752) );
  INV_X1 U17294 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15955) );
  NAND4_X1 U17295 ( .A1(P2_REG1_REG_28__SCAN_IN), .A2(n15956), .A3(n10597), 
        .A4(n15955), .ZN(n15750) );
  NAND4_X1 U17296 ( .A1(SI_29_), .A2(P3_REG3_REG_0__SCAN_IN), .A3(
        P3_ADDR_REG_10__SCAN_IN), .A4(n15966), .ZN(n15749) );
  NOR4_X1 U17297 ( .A1(P3_REG2_REG_20__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), 
        .A3(P2_REG2_REG_27__SCAN_IN), .A4(P2_REG0_REG_4__SCAN_IN), .ZN(n15730)
         );
  INV_X1 U17298 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n15953) );
  NOR4_X1 U17299 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n15953), .A3(n15952), .A4(
        n10591), .ZN(n15729) );
  NAND4_X1 U17300 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_DATAO_REG_0__SCAN_IN), 
        .A3(n15873), .A4(n8992), .ZN(n15727) );
  NAND4_X1 U17301 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(P3_REG2_REG_26__SCAN_IN), 
        .A3(n15682), .A4(n8323), .ZN(n15726) );
  OR4_X1 U17302 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .A3(P2_REG3_REG_25__SCAN_IN), .A4(P3_REG3_REG_25__SCAN_IN), .ZN(n15725) );
  NAND4_X1 U17303 ( .A1(n15723), .A2(n7372), .A3(P3_D_REG_19__SCAN_IN), .A4(
        P2_D_REG_17__SCAN_IN), .ZN(n15724) );
  NOR4_X1 U17304 ( .A1(n15727), .A2(n15726), .A3(n15725), .A4(n15724), .ZN(
        n15728) );
  NAND3_X1 U17305 ( .A1(n15730), .A2(n15729), .A3(n15728), .ZN(n15748) );
  NAND4_X1 U17306 ( .A1(n15732), .A2(n15731), .A3(P2_REG3_REG_10__SCAN_IN), 
        .A4(P2_REG0_REG_27__SCAN_IN), .ZN(n15733) );
  NOR3_X1 U17307 ( .A1(n15733), .A2(P1_IR_REG_27__SCAN_IN), .A3(n15898), .ZN(
        n15746) );
  INV_X1 U17308 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n15734) );
  NOR4_X1 U17309 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(n15735), .A3(n15734), .A4(
        n15756), .ZN(n15736) );
  NAND3_X1 U17310 ( .A1(P3_REG2_REG_15__SCAN_IN), .A2(P3_REG2_REG_16__SCAN_IN), 
        .A3(n15736), .ZN(n15744) );
  NOR4_X1 U17311 ( .A1(P2_REG0_REG_9__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), 
        .A3(n10609), .A4(n15781), .ZN(n15742) );
  NOR4_X1 U17312 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P3_ADDR_REG_16__SCAN_IN), 
        .A3(n15772), .A4(n15737), .ZN(n15741) );
  NOR4_X1 U17313 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P3_DATAO_REG_18__SCAN_IN), 
        .A3(n15797), .A4(n15790), .ZN(n15740) );
  NOR4_X1 U17314 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(SI_0_), .A3(
        P2_REG2_REG_9__SCAN_IN), .A4(n15738), .ZN(n15739) );
  NAND4_X1 U17315 ( .A1(n15742), .A2(n15741), .A3(n15740), .A4(n15739), .ZN(
        n15743) );
  NOR4_X1 U17316 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(P2_REG2_REG_21__SCAN_IN), 
        .A3(n15744), .A4(n15743), .ZN(n15745) );
  NAND4_X1 U17317 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(n15746), .A3(n15745), 
        .A4(n15909), .ZN(n15747) );
  NOR4_X1 U17318 ( .A1(n15750), .A2(n15749), .A3(n15748), .A4(n15747), .ZN(
        n15751) );
  NAND4_X1 U17319 ( .A1(n15754), .A2(n15753), .A3(n15752), .A4(n15751), .ZN(
        n15984) );
  AOI22_X1 U17320 ( .A1(n12231), .A2(keyinput50), .B1(keyinput42), .B2(n15756), 
        .ZN(n15755) );
  OAI221_X1 U17321 ( .B1(n12231), .B2(keyinput50), .C1(n15756), .C2(keyinput42), .A(n15755), .ZN(n15767) );
  AOI22_X1 U17322 ( .A1(n15759), .A2(keyinput87), .B1(keyinput69), .B2(n15758), 
        .ZN(n15757) );
  OAI221_X1 U17323 ( .B1(n15759), .B2(keyinput87), .C1(n15758), .C2(keyinput69), .A(n15757), .ZN(n15766) );
  XNOR2_X1 U17324 ( .A(n15760), .B(keyinput81), .ZN(n15765) );
  XNOR2_X1 U17325 ( .A(P3_IR_REG_20__SCAN_IN), .B(keyinput118), .ZN(n15763) );
  XNOR2_X1 U17326 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput107), .ZN(n15762) );
  XNOR2_X1 U17327 ( .A(P2_REG0_REG_28__SCAN_IN), .B(keyinput83), .ZN(n15761)
         );
  NAND3_X1 U17328 ( .A1(n15763), .A2(n15762), .A3(n15761), .ZN(n15764) );
  NOR4_X1 U17329 ( .A1(n15767), .A2(n15766), .A3(n15765), .A4(n15764), .ZN(
        n15809) );
  AOI22_X1 U17330 ( .A1(n15769), .A2(keyinput55), .B1(keyinput16), .B2(n10609), 
        .ZN(n15768) );
  OAI221_X1 U17331 ( .B1(n15769), .B2(keyinput55), .C1(n10609), .C2(keyinput16), .A(n15768), .ZN(n15779) );
  AOI22_X1 U17332 ( .A1(n15772), .A2(keyinput10), .B1(keyinput71), .B2(n15771), 
        .ZN(n15770) );
  OAI221_X1 U17333 ( .B1(n15772), .B2(keyinput10), .C1(n15771), .C2(keyinput71), .A(n15770), .ZN(n15778) );
  XNOR2_X1 U17334 ( .A(P2_REG0_REG_17__SCAN_IN), .B(keyinput82), .ZN(n15776)
         );
  XNOR2_X1 U17335 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput111), .ZN(n15775) );
  XNOR2_X1 U17336 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput56), .ZN(n15774)
         );
  XNOR2_X1 U17337 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput5), .ZN(n15773) );
  NAND4_X1 U17338 ( .A1(n15776), .A2(n15775), .A3(n15774), .A4(n15773), .ZN(
        n15777) );
  NOR3_X1 U17339 ( .A1(n15779), .A2(n15778), .A3(n15777), .ZN(n15808) );
  AOI22_X1 U17340 ( .A1(n15782), .A2(keyinput86), .B1(keyinput127), .B2(n15781), .ZN(n15780) );
  OAI221_X1 U17341 ( .B1(n15782), .B2(keyinput86), .C1(n15781), .C2(
        keyinput127), .A(n15780), .ZN(n15793) );
  XOR2_X1 U17342 ( .A(SI_0_), .B(keyinput41), .Z(n15785) );
  XNOR2_X1 U17343 ( .A(n15783), .B(keyinput113), .ZN(n15784) );
  NOR2_X1 U17344 ( .A1(n15785), .A2(n15784), .ZN(n15789) );
  XNOR2_X1 U17345 ( .A(keyinput65), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n15788) );
  XNOR2_X1 U17346 ( .A(P3_REG1_REG_13__SCAN_IN), .B(keyinput66), .ZN(n15787)
         );
  XNOR2_X1 U17347 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput68), .ZN(n15786) );
  NAND4_X1 U17348 ( .A1(n15789), .A2(n15788), .A3(n15787), .A4(n15786), .ZN(
        n15792) );
  XNOR2_X1 U17349 ( .A(n15790), .B(keyinput89), .ZN(n15791) );
  NOR3_X1 U17350 ( .A1(n15793), .A2(n15792), .A3(n15791), .ZN(n15807) );
  AOI22_X1 U17351 ( .A1(n12114), .A2(keyinput39), .B1(keyinput99), .B2(n15795), 
        .ZN(n15794) );
  OAI221_X1 U17352 ( .B1(n12114), .B2(keyinput39), .C1(n15795), .C2(keyinput99), .A(n15794), .ZN(n15805) );
  AOI22_X1 U17353 ( .A1(n15798), .A2(keyinput96), .B1(n15797), .B2(keyinput30), 
        .ZN(n15796) );
  OAI221_X1 U17354 ( .B1(n15798), .B2(keyinput96), .C1(n15797), .C2(keyinput30), .A(n15796), .ZN(n15804) );
  XNOR2_X1 U17355 ( .A(P1_REG0_REG_21__SCAN_IN), .B(keyinput74), .ZN(n15802)
         );
  XNOR2_X1 U17356 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput124), .ZN(n15801) );
  XNOR2_X1 U17357 ( .A(P3_IR_REG_26__SCAN_IN), .B(keyinput126), .ZN(n15800) );
  XNOR2_X1 U17358 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput33), .ZN(n15799) );
  NAND4_X1 U17359 ( .A1(n15802), .A2(n15801), .A3(n15800), .A4(n15799), .ZN(
        n15803) );
  NOR3_X1 U17360 ( .A1(n15805), .A2(n15804), .A3(n15803), .ZN(n15806) );
  NAND4_X1 U17361 ( .A1(n15809), .A2(n15808), .A3(n15807), .A4(n15806), .ZN(
        n15982) );
  XNOR2_X1 U17362 ( .A(n15810), .B(keyinput73), .ZN(n15814) );
  XNOR2_X1 U17363 ( .A(n15811), .B(keyinput106), .ZN(n15813) );
  XNOR2_X1 U17364 ( .A(keyinput34), .B(n9314), .ZN(n15812) );
  NOR3_X1 U17365 ( .A1(n15814), .A2(n15813), .A3(n15812), .ZN(n15818) );
  XOR2_X1 U17366 ( .A(n15815), .B(keyinput12), .Z(n15817) );
  XNOR2_X1 U17367 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput24), .ZN(n15816) );
  NAND3_X1 U17368 ( .A1(n15818), .A2(n15817), .A3(n15816), .ZN(n15824) );
  AOI22_X1 U17369 ( .A1(n15820), .A2(keyinput114), .B1(n14237), .B2(keyinput37), .ZN(n15819) );
  OAI221_X1 U17370 ( .B1(n15820), .B2(keyinput114), .C1(n14237), .C2(
        keyinput37), .A(n15819), .ZN(n15823) );
  XNOR2_X1 U17371 ( .A(n15821), .B(keyinput109), .ZN(n15822) );
  NOR3_X1 U17372 ( .A1(n15824), .A2(n15823), .A3(n15822), .ZN(n15869) );
  AOI22_X1 U17373 ( .A1(n15827), .A2(keyinput95), .B1(n15826), .B2(keyinput59), 
        .ZN(n15825) );
  OAI221_X1 U17374 ( .B1(n15827), .B2(keyinput95), .C1(n15826), .C2(keyinput59), .A(n15825), .ZN(n15837) );
  AOI22_X1 U17375 ( .A1(n15830), .A2(keyinput102), .B1(n15829), .B2(
        keyinput103), .ZN(n15828) );
  OAI221_X1 U17376 ( .B1(n15830), .B2(keyinput102), .C1(n15829), .C2(
        keyinput103), .A(n15828), .ZN(n15836) );
  XOR2_X1 U17377 ( .A(n10175), .B(keyinput119), .Z(n15834) );
  XNOR2_X1 U17378 ( .A(P3_IR_REG_15__SCAN_IN), .B(keyinput11), .ZN(n15833) );
  XNOR2_X1 U17379 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput57), .ZN(n15832) );
  XNOR2_X1 U17380 ( .A(P1_REG3_REG_9__SCAN_IN), .B(keyinput84), .ZN(n15831) );
  NAND4_X1 U17381 ( .A1(n15834), .A2(n15833), .A3(n15832), .A4(n15831), .ZN(
        n15835) );
  NOR3_X1 U17382 ( .A1(n15837), .A2(n15836), .A3(n15835), .ZN(n15868) );
  AOI22_X1 U17383 ( .A1(n15840), .A2(keyinput120), .B1(keyinput45), .B2(n15839), .ZN(n15838) );
  OAI221_X1 U17384 ( .B1(n15840), .B2(keyinput120), .C1(n15839), .C2(
        keyinput45), .A(n15838), .ZN(n15851) );
  AOI22_X1 U17385 ( .A1(n15843), .A2(keyinput53), .B1(keyinput80), .B2(n15842), 
        .ZN(n15841) );
  OAI221_X1 U17386 ( .B1(n15843), .B2(keyinput53), .C1(n15842), .C2(keyinput80), .A(n15841), .ZN(n15850) );
  AOI22_X1 U17387 ( .A1(n7297), .A2(keyinput29), .B1(keyinput72), .B2(n15845), 
        .ZN(n15844) );
  OAI221_X1 U17388 ( .B1(n7297), .B2(keyinput29), .C1(n15845), .C2(keyinput72), 
        .A(n15844), .ZN(n15849) );
  XNOR2_X1 U17389 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput27), .ZN(n15847)
         );
  XNOR2_X1 U17390 ( .A(P2_REG1_REG_23__SCAN_IN), .B(keyinput100), .ZN(n15846)
         );
  NAND2_X1 U17391 ( .A1(n15847), .A2(n15846), .ZN(n15848) );
  NOR4_X1 U17392 ( .A1(n15851), .A2(n15850), .A3(n15849), .A4(n15848), .ZN(
        n15867) );
  AOI22_X1 U17393 ( .A1(n15854), .A2(keyinput47), .B1(n15853), .B2(keyinput115), .ZN(n15852) );
  OAI221_X1 U17394 ( .B1(n15854), .B2(keyinput47), .C1(n15853), .C2(
        keyinput115), .A(n15852), .ZN(n15865) );
  AOI22_X1 U17395 ( .A1(n12849), .A2(keyinput91), .B1(keyinput98), .B2(n15856), 
        .ZN(n15855) );
  OAI221_X1 U17396 ( .B1(n12849), .B2(keyinput91), .C1(n15856), .C2(keyinput98), .A(n15855), .ZN(n15864) );
  AOI22_X1 U17397 ( .A1(n15859), .A2(keyinput61), .B1(keyinput22), .B2(n15858), 
        .ZN(n15857) );
  OAI221_X1 U17398 ( .B1(n15859), .B2(keyinput61), .C1(n15858), .C2(keyinput22), .A(n15857), .ZN(n15863) );
  XNOR2_X1 U17399 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput2), .ZN(n15861) );
  XNOR2_X1 U17400 ( .A(P1_REG0_REG_11__SCAN_IN), .B(keyinput104), .ZN(n15860)
         );
  NAND2_X1 U17401 ( .A1(n15861), .A2(n15860), .ZN(n15862) );
  NOR4_X1 U17402 ( .A1(n15865), .A2(n15864), .A3(n15863), .A4(n15862), .ZN(
        n15866) );
  NAND4_X1 U17403 ( .A1(n15869), .A2(n15868), .A3(n15867), .A4(n15866), .ZN(
        n15981) );
  AOI22_X1 U17404 ( .A1(n11408), .A2(keyinput79), .B1(keyinput123), .B2(n15682), .ZN(n15870) );
  OAI221_X1 U17405 ( .B1(n11408), .B2(keyinput79), .C1(n15682), .C2(
        keyinput123), .A(n15870), .ZN(n15881) );
  AOI22_X1 U17406 ( .A1(n15873), .A2(keyinput0), .B1(n15872), .B2(keyinput97), 
        .ZN(n15871) );
  OAI221_X1 U17407 ( .B1(n15873), .B2(keyinput0), .C1(n15872), .C2(keyinput97), 
        .A(n15871), .ZN(n15880) );
  AOI22_X1 U17408 ( .A1(n15875), .A2(keyinput15), .B1(n10146), .B2(keyinput18), 
        .ZN(n15874) );
  OAI221_X1 U17409 ( .B1(n15875), .B2(keyinput15), .C1(n10146), .C2(keyinput18), .A(n15874), .ZN(n15879) );
  XNOR2_X1 U17410 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(keyinput13), .ZN(n15877)
         );
  XNOR2_X1 U17411 ( .A(P1_REG0_REG_18__SCAN_IN), .B(keyinput70), .ZN(n15876)
         );
  NAND2_X1 U17412 ( .A1(n15877), .A2(n15876), .ZN(n15878) );
  NOR4_X1 U17413 ( .A1(n15881), .A2(n15880), .A3(n15879), .A4(n15878), .ZN(
        n15920) );
  AOI22_X1 U17414 ( .A1(n14071), .A2(keyinput51), .B1(keyinput85), .B2(n15883), 
        .ZN(n15882) );
  OAI221_X1 U17415 ( .B1(n14071), .B2(keyinput51), .C1(n15883), .C2(keyinput85), .A(n15882), .ZN(n15892) );
  INV_X1 U17416 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15885) );
  AOI22_X1 U17417 ( .A1(n15885), .A2(keyinput36), .B1(n8992), .B2(keyinput76), 
        .ZN(n15884) );
  OAI221_X1 U17418 ( .B1(n15885), .B2(keyinput36), .C1(n8992), .C2(keyinput76), 
        .A(n15884), .ZN(n15891) );
  XNOR2_X1 U17419 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput125), .ZN(n15889) );
  XNOR2_X1 U17420 ( .A(P3_REG2_REG_20__SCAN_IN), .B(keyinput93), .ZN(n15888)
         );
  XNOR2_X1 U17421 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput6), .ZN(n15887) );
  XNOR2_X1 U17422 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput4), .ZN(n15886) );
  NAND4_X1 U17423 ( .A1(n15889), .A2(n15888), .A3(n15887), .A4(n15886), .ZN(
        n15890) );
  NOR3_X1 U17424 ( .A1(n15892), .A2(n15891), .A3(n15890), .ZN(n15919) );
  AOI22_X1 U17425 ( .A1(n15895), .A2(keyinput62), .B1(n15894), .B2(keyinput121), .ZN(n15893) );
  OAI221_X1 U17426 ( .B1(n15895), .B2(keyinput62), .C1(n15894), .C2(
        keyinput121), .A(n15893), .ZN(n15905) );
  AOI22_X1 U17427 ( .A1(n14159), .A2(keyinput20), .B1(keyinput78), .B2(n15897), 
        .ZN(n15896) );
  OAI221_X1 U17428 ( .B1(n14159), .B2(keyinput20), .C1(n15897), .C2(keyinput78), .A(n15896), .ZN(n15904) );
  XOR2_X1 U17429 ( .A(n15898), .B(keyinput44), .Z(n15902) );
  XNOR2_X1 U17430 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput35), .ZN(n15901) );
  XNOR2_X1 U17431 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput117), .ZN(n15900)
         );
  XNOR2_X1 U17432 ( .A(P3_REG0_REG_26__SCAN_IN), .B(keyinput112), .ZN(n15899)
         );
  NAND4_X1 U17433 ( .A1(n15902), .A2(n15901), .A3(n15900), .A4(n15899), .ZN(
        n15903) );
  NOR3_X1 U17434 ( .A1(n15905), .A2(n15904), .A3(n15903), .ZN(n15918) );
  AOI22_X1 U17435 ( .A1(n8323), .A2(keyinput32), .B1(n15907), .B2(keyinput19), 
        .ZN(n15906) );
  OAI221_X1 U17436 ( .B1(n8323), .B2(keyinput32), .C1(n15907), .C2(keyinput19), 
        .A(n15906), .ZN(n15916) );
  AOI22_X1 U17437 ( .A1(n7372), .A2(keyinput94), .B1(n15909), .B2(keyinput9), 
        .ZN(n15908) );
  OAI221_X1 U17438 ( .B1(n7372), .B2(keyinput94), .C1(n15909), .C2(keyinput9), 
        .A(n15908), .ZN(n15915) );
  XOR2_X1 U17439 ( .A(n14177), .B(keyinput46), .Z(n15913) );
  XNOR2_X1 U17440 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput28), .ZN(n15912)
         );
  XNOR2_X1 U17441 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput92), .ZN(n15911) );
  XNOR2_X1 U17442 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput14), .ZN(n15910) );
  NAND4_X1 U17443 ( .A1(n15913), .A2(n15912), .A3(n15911), .A4(n15910), .ZN(
        n15914) );
  NOR3_X1 U17444 ( .A1(n15916), .A2(n15915), .A3(n15914), .ZN(n15917) );
  NAND4_X1 U17445 ( .A1(n15920), .A2(n15919), .A3(n15918), .A4(n15917), .ZN(
        n15980) );
  AOI22_X1 U17446 ( .A1(n15923), .A2(keyinput122), .B1(keyinput40), .B2(n15922), .ZN(n15921) );
  OAI221_X1 U17447 ( .B1(n15923), .B2(keyinput122), .C1(n15922), .C2(
        keyinput40), .A(n15921), .ZN(n15935) );
  AOI22_X1 U17448 ( .A1(n15703), .A2(keyinput63), .B1(n15925), .B2(keyinput54), 
        .ZN(n15924) );
  OAI221_X1 U17449 ( .B1(n15703), .B2(keyinput63), .C1(n15925), .C2(keyinput54), .A(n15924), .ZN(n15934) );
  AOI22_X1 U17450 ( .A1(n15928), .A2(keyinput60), .B1(n15927), .B2(keyinput21), 
        .ZN(n15926) );
  OAI221_X1 U17451 ( .B1(n15928), .B2(keyinput60), .C1(n15927), .C2(keyinput21), .A(n15926), .ZN(n15933) );
  XOR2_X1 U17452 ( .A(n15929), .B(keyinput116), .Z(n15931) );
  XNOR2_X1 U17453 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput48), .ZN(n15930) );
  NAND2_X1 U17454 ( .A1(n15931), .A2(n15930), .ZN(n15932) );
  NOR4_X1 U17455 ( .A1(n15935), .A2(n15934), .A3(n15933), .A4(n15932), .ZN(
        n15978) );
  XOR2_X1 U17456 ( .A(SI_1_), .B(keyinput8), .Z(n15936) );
  AOI21_X1 U17457 ( .B1(n15985), .B2(keyinput52), .A(n15936), .ZN(n15939) );
  XNOR2_X1 U17458 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput26), .ZN(n15938) );
  XNOR2_X1 U17459 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput1), .ZN(n15937) );
  NAND3_X1 U17460 ( .A1(n15939), .A2(n15938), .A3(n15937), .ZN(n15948) );
  AOI22_X1 U17461 ( .A1(n15942), .A2(keyinput3), .B1(n15941), .B2(keyinput58), 
        .ZN(n15940) );
  OAI221_X1 U17462 ( .B1(n15942), .B2(keyinput3), .C1(n15941), .C2(keyinput58), 
        .A(n15940), .ZN(n15947) );
  XNOR2_X1 U17463 ( .A(keyinput23), .B(n15943), .ZN(n15946) );
  INV_X1 U17464 ( .A(SI_28_), .ZN(n15944) );
  XNOR2_X1 U17465 ( .A(keyinput64), .B(n15944), .ZN(n15945) );
  NOR4_X1 U17466 ( .A1(n15948), .A2(n15947), .A3(n15946), .A4(n15945), .ZN(
        n15977) );
  AOI22_X1 U17467 ( .A1(n15950), .A2(keyinput90), .B1(keyinput88), .B2(n10585), 
        .ZN(n15949) );
  OAI221_X1 U17468 ( .B1(n15950), .B2(keyinput90), .C1(n10585), .C2(keyinput88), .A(n15949), .ZN(n15962) );
  AOI22_X1 U17469 ( .A1(n15953), .A2(keyinput17), .B1(n15952), .B2(keyinput110), .ZN(n15951) );
  OAI221_X1 U17470 ( .B1(n15953), .B2(keyinput17), .C1(n15952), .C2(
        keyinput110), .A(n15951), .ZN(n15961) );
  AOI22_X1 U17471 ( .A1(n15956), .A2(keyinput7), .B1(keyinput67), .B2(n15955), 
        .ZN(n15954) );
  OAI221_X1 U17472 ( .B1(n15956), .B2(keyinput7), .C1(n15955), .C2(keyinput67), 
        .A(n15954), .ZN(n15960) );
  XNOR2_X1 U17473 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(keyinput25), .ZN(n15958) );
  XNOR2_X1 U17474 ( .A(keyinput31), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n15957) );
  NAND2_X1 U17475 ( .A1(n15958), .A2(n15957), .ZN(n15959) );
  NOR4_X1 U17476 ( .A1(n15962), .A2(n15961), .A3(n15960), .A4(n15959), .ZN(
        n15976) );
  AOI22_X1 U17477 ( .A1(n15965), .A2(keyinput77), .B1(keyinput49), .B2(n15964), 
        .ZN(n15963) );
  OAI221_X1 U17478 ( .B1(n15965), .B2(keyinput77), .C1(n15964), .C2(keyinput49), .A(n15963), .ZN(n15974) );
  XNOR2_X1 U17479 ( .A(keyinput105), .B(n15966), .ZN(n15973) );
  XNOR2_X1 U17480 ( .A(keyinput101), .B(n10597), .ZN(n15972) );
  XNOR2_X1 U17481 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput108), .ZN(n15970)
         );
  XNOR2_X1 U17482 ( .A(P3_IR_REG_30__SCAN_IN), .B(keyinput38), .ZN(n15969) );
  XNOR2_X1 U17483 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput75), .ZN(n15968) );
  XNOR2_X1 U17484 ( .A(keyinput43), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n15967)
         );
  NAND4_X1 U17485 ( .A1(n15970), .A2(n15969), .A3(n15968), .A4(n15967), .ZN(
        n15971) );
  NOR4_X1 U17486 ( .A1(n15974), .A2(n15973), .A3(n15972), .A4(n15971), .ZN(
        n15975) );
  NAND4_X1 U17487 ( .A1(n15978), .A2(n15977), .A3(n15976), .A4(n15975), .ZN(
        n15979) );
  NOR4_X1 U17488 ( .A1(n15982), .A2(n15981), .A3(n15980), .A4(n15979), .ZN(
        n15983) );
  OAI221_X1 U17489 ( .B1(keyinput52), .B2(n15985), .C1(keyinput52), .C2(n15984), .A(n15983), .ZN(n15986) );
  XNOR2_X1 U17490 ( .A(n15987), .B(n15986), .ZN(P3_U3150) );
endmodule

