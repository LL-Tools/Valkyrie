

module b20_C_gen_AntiSAT_k_128_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4351, n4352, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217;

  INV_X2 U4857 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND2_X1 U4858 ( .A1(n5552), .A2(n5551), .ZN(n8987) );
  XNOR2_X1 U4859 ( .A(n4433), .B(n7000), .ZN(n6882) );
  CLKBUF_X2 U4860 ( .A(n5045), .Z(n6193) );
  INV_X1 U4861 ( .A(n8412), .ZN(n8432) );
  BUF_X2 U4863 ( .A(n4983), .Z(n9269) );
  NOR2_X1 U4864 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4872) );
  NAND2_X1 U4865 ( .A1(n9006), .A2(n5530), .ZN(n5552) );
  NAND3_X1 U4866 ( .A1(n5046), .A2(n6946), .A3(n4987), .ZN(n5032) );
  INV_X2 U4867 ( .A(n5628), .ZN(n5139) );
  INV_X1 U4868 ( .A(n5026), .ZN(n5461) );
  INV_X1 U4869 ( .A(n4962), .ZN(n4938) );
  INV_X1 U4870 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10141) );
  AND2_X1 U4871 ( .A1(n7090), .A2(n7089), .ZN(n7174) );
  INV_X2 U4872 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4837) );
  OR2_X1 U4873 ( .A1(n5829), .A2(n4837), .ZN(n5831) );
  OR2_X1 U4874 ( .A1(n5552), .A2(n5551), .ZN(n5553) );
  INV_X1 U4875 ( .A(n5033), .ZN(n5167) );
  AND2_X1 U4876 ( .A1(n9495), .A2(n9509), .ZN(n9490) );
  NAND2_X1 U4877 ( .A1(n5026), .A2(n6389), .ZN(n5083) );
  XNOR2_X1 U4878 ( .A(n8493), .B(n8509), .ZN(n8470) );
  XNOR2_X1 U4879 ( .A(n8547), .B(n8526), .ZN(n8527) );
  INV_X1 U4880 ( .A(n5827), .ZN(n8224) );
  NAND2_X1 U4881 ( .A1(n6144), .A2(n6146), .ZN(n6147) );
  OAI211_X1 U4882 ( .C1(n5026), .C2(n6451), .A(n5085), .B(n5084), .ZN(n9824)
         );
  INV_X1 U4883 ( .A(n5057), .ZN(n5619) );
  INV_X1 U4884 ( .A(n7877), .ZN(n6551) );
  AND4_X1 U4886 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n4351)
         );
  INV_X2 U4887 ( .A(n9468), .ZN(n9826) );
  AOI21_X2 U4888 ( .B1(n7405), .B2(n4792), .A(n4790), .ZN(n5360) );
  NAND2_X2 U4889 ( .A1(n5278), .A2(n5277), .ZN(n7405) );
  AND2_X2 U4890 ( .A1(n4866), .A2(n4590), .ZN(n4589) );
  INV_X1 U4891 ( .A(n5073), .ZN(n5471) );
  OAI21_X2 U4892 ( .B1(n5319), .B2(n4907), .A(n5340), .ZN(n6529) );
  NAND2_X4 U4894 ( .A1(n6130), .A2(n6131), .ZN(n5832) );
  XNOR2_X2 U4895 ( .A(n4579), .B(n5781), .ZN(n6131) );
  OAI21_X2 U4896 ( .B1(n7019), .B2(n8266), .A(n7018), .ZN(n7020) );
  OAI21_X1 U4897 ( .B1(n9103), .B2(n9102), .A(n9101), .ZN(n9105) );
  NAND2_X1 U4898 ( .A1(n9046), .A2(n5603), .ZN(n9016) );
  AOI211_X1 U4899 ( .C1(n4671), .C2(n8420), .A(n8419), .B(n8421), .ZN(n8424)
         );
  XNOR2_X1 U4900 ( .A(n7638), .B(n7637), .ZN(n7640) );
  NAND2_X1 U4901 ( .A1(n8497), .A2(n4749), .ZN(n4748) );
  AOI21_X1 U4902 ( .B1(n4568), .B2(n4570), .A(n4392), .ZN(n4566) );
  NOR2_X1 U4903 ( .A1(n4859), .A2(n4397), .ZN(n4858) );
  OR2_X1 U4904 ( .A1(n8470), .A2(n4747), .ZN(n4435) );
  NAND2_X1 U4905 ( .A1(n7981), .A2(n7980), .ZN(n8046) );
  NAND2_X1 U4906 ( .A1(n8469), .A2(n8468), .ZN(n8493) );
  XNOR2_X1 U4907 ( .A(n7425), .B(n7426), .ZN(n7244) );
  AND2_X1 U4908 ( .A1(n4447), .A2(n4446), .ZN(n4792) );
  NAND2_X1 U4909 ( .A1(n6053), .A2(n6052), .ZN(n8914) );
  NOR2_X1 U4910 ( .A1(n7471), .A2(n9611), .ZN(n9508) );
  OR2_X1 U4911 ( .A1(n7564), .A2(n5981), .ZN(n9701) );
  NAND2_X1 U4912 ( .A1(n6028), .A2(n6027), .ZN(n8938) );
  NOR2_X1 U4913 ( .A1(n5982), .A2(n5966), .ZN(n5981) );
  XNOR2_X1 U4914 ( .A(n7174), .B(n7175), .ZN(n7091) );
  NAND2_X1 U4915 ( .A1(n8357), .A2(n8340), .ZN(n8828) );
  OR2_X1 U4916 ( .A1(n7318), .A2(n8249), .ZN(n7320) );
  NAND2_X1 U4917 ( .A1(n4819), .A2(n4821), .ZN(n5484) );
  NOR2_X1 U4918 ( .A1(n9939), .A2(n9925), .ZN(n8944) );
  NAND2_X1 U4919 ( .A1(n4759), .A2(n4380), .ZN(n4758) );
  OAI21_X1 U4920 ( .B1(n6520), .B2(n5827), .A(n5955), .ZN(n9931) );
  NAND2_X2 U4921 ( .A1(n6614), .A2(n9390), .ZN(n9468) );
  NAND2_X1 U4922 ( .A1(n5252), .A2(n5251), .ZN(n7127) );
  INV_X1 U4923 ( .A(n6962), .ZN(n9851) );
  OR2_X1 U4924 ( .A1(n6875), .A2(n6952), .ZN(n7678) );
  NOR2_X1 U4925 ( .A1(n7063), .A2(n7064), .ZN(n7205) );
  NAND2_X1 U4926 ( .A1(n5205), .A2(n5204), .ZN(n6875) );
  INV_X1 U4927 ( .A(n5167), .ZN(n5681) );
  INV_X1 U4928 ( .A(n6293), .ZN(n6914) );
  AND2_X1 U4929 ( .A1(n4817), .A2(n4815), .ZN(n5340) );
  NAND4_X1 U4931 ( .A1(n5077), .A2(n5076), .A3(n5075), .A4(n5074), .ZN(n9142)
         );
  NAND4_X1 U4932 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(n4911), .ZN(n6540)
         );
  OR2_X1 U4933 ( .A1(n7795), .A2(n9269), .ZN(n6324) );
  INV_X1 U4934 ( .A(n9824), .ZN(n6587) );
  NAND2_X1 U4935 ( .A1(n4369), .A2(n5844), .ZN(n8465) );
  INV_X1 U4936 ( .A(n5035), .ZN(n5349) );
  INV_X1 U4937 ( .A(n7651), .ZN(n5452) );
  XNOR2_X1 U4938 ( .A(n4982), .B(P1_IR_REG_19__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U4939 ( .A1(n5693), .A2(n4967), .ZN(n5046) );
  NAND2_X1 U4940 ( .A1(n4975), .A2(n4974), .ZN(n5718) );
  AND2_X2 U4941 ( .A1(n7958), .A2(n4948), .ZN(n5073) );
  AND2_X2 U4942 ( .A1(n4948), .A2(n4942), .ZN(n7651) );
  NAND2_X1 U4943 ( .A1(n4986), .A2(n5710), .ZN(n7795) );
  CLKBUF_X1 U4944 ( .A(n4946), .Z(n7958) );
  MUX2_X1 U4945 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4972), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n4975) );
  AND2_X1 U4946 ( .A1(n5460), .A2(n4981), .ZN(n4982) );
  INV_X2 U4947 ( .A(n5832), .ZN(n6385) );
  OR2_X1 U4948 ( .A1(n4973), .A2(n5290), .ZN(n4969) );
  OR2_X1 U4949 ( .A1(n6787), .A2(n6788), .ZN(n6785) );
  NAND2_X1 U4950 ( .A1(n4979), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5460) );
  XNOR2_X1 U4951 ( .A(n4490), .B(n4939), .ZN(n9691) );
  INV_X1 U4952 ( .A(n5791), .ZN(n8962) );
  XNOR2_X1 U4953 ( .A(n5785), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5791) );
  AND2_X1 U4954 ( .A1(n4462), .A2(n4415), .ZN(n4801) );
  NAND2_X1 U4955 ( .A1(n4989), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4490) );
  NAND2_X1 U4956 ( .A1(n4401), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5785) );
  OR2_X1 U4957 ( .A1(n8955), .A2(n4837), .ZN(n5784) );
  INV_X1 U4958 ( .A(n5368), .ZN(n4931) );
  AND2_X1 U4959 ( .A1(n4372), .A2(n4869), .ZN(n4868) );
  NOR3_X1 U4960 ( .A1(n4936), .A2(P1_IR_REG_15__SCAN_IN), .A3(
        P1_IR_REG_25__SCAN_IN), .ZN(n4892) );
  NOR2_X1 U4961 ( .A1(n4676), .A2(n4675), .ZN(n4677) );
  AND2_X1 U4962 ( .A1(n4796), .A2(n4794), .ZN(n5817) );
  AND2_X1 U4963 ( .A1(n4867), .A2(n5745), .ZN(n4866) );
  AND3_X1 U4964 ( .A1(n4968), .A2(n4958), .A3(n4956), .ZN(n4935) );
  NOR2_X1 U4965 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5746) );
  NOR2_X1 U4966 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5747) );
  NOR2_X1 U4967 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5748) );
  NOR2_X1 U4968 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5749) );
  INV_X1 U4969 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5830) );
  NOR2_X1 U4970 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5829) );
  INV_X1 U4971 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5743) );
  NOR2_X1 U4972 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4867) );
  INV_X4 U4973 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OAI21_X2 U4974 ( .B1(n6147), .B2(P2_D_REG_0__SCAN_IN), .A(n6578), .ZN(n7019)
         );
  OAI21_X2 U4975 ( .B1(n8712), .B2(n8720), .A(n6061), .ZN(n8691) );
  XNOR2_X1 U4977 ( .A(n5831), .B(n5830), .ZN(n6708) );
  AND2_X4 U4978 ( .A1(n5787), .A2(n8962), .ZN(n5840) );
  OAI21_X2 U4979 ( .B1(n7075), .B2(n7073), .A(n7071), .ZN(n7300) );
  AOI21_X2 U4980 ( .B1(n6909), .B2(n5144), .A(n4402), .ZN(n7075) );
  AOI21_X2 U4981 ( .B1(n6555), .B2(n6556), .A(n4904), .ZN(n9057) );
  OAI22_X2 U4982 ( .A1(n6549), .A2(n6550), .B1(n5072), .B2(n5071), .ZN(n6555)
         );
  AND2_X1 U4983 ( .A1(n5046), .A2(n5013), .ZN(n5033) );
  NAND2_X1 U4984 ( .A1(n5389), .A2(SI_15_), .ZN(n5388) );
  AOI211_X1 U4985 ( .C1(n7800), .C2(n7799), .A(n7866), .B(n7798), .ZN(n4622)
         );
  NAND2_X1 U4986 ( .A1(n5643), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5730) );
  INV_X1 U4987 ( .A(n4602), .ZN(n4598) );
  NAND2_X1 U4988 ( .A1(n4608), .A2(n4603), .ZN(n4602) );
  INV_X1 U4989 ( .A(n7707), .ZN(n4603) );
  INV_X1 U4990 ( .A(n4607), .ZN(n4606) );
  OAI22_X1 U4991 ( .A1(n7689), .A2(n7690), .B1(n7698), .B2(n7699), .ZN(n4607)
         );
  NAND2_X1 U4992 ( .A1(n8763), .A2(n8412), .ZN(n4530) );
  NAND2_X1 U4993 ( .A1(n4617), .A2(n4616), .ZN(n4615) );
  INV_X1 U4994 ( .A(n7753), .ZN(n4616) );
  NOR2_X1 U4995 ( .A1(n4668), .A2(n8419), .ZN(n4663) );
  INV_X1 U4996 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5442) );
  INV_X1 U4997 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4954) );
  INV_X1 U4998 ( .A(n5394), .ZN(n4955) );
  NAND2_X1 U4999 ( .A1(n8061), .A2(n8001), .ZN(n4860) );
  INV_X1 U5000 ( .A(n5787), .ZN(n5792) );
  OR2_X1 U5001 ( .A1(n8671), .A2(n8090), .ZN(n8408) );
  NAND2_X1 U5002 ( .A1(n5763), .A2(n5762), .ZN(n6130) );
  OAI21_X1 U5003 ( .B1(n5760), .B2(n5759), .A(n5758), .ZN(n5763) );
  NAND2_X1 U5004 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5759), .ZN(n5758) );
  INV_X1 U5005 ( .A(n8413), .ZN(n4672) );
  NOR2_X1 U5006 ( .A1(n4665), .A2(n8240), .ZN(n4664) );
  INV_X1 U5007 ( .A(n8410), .ZN(n4665) );
  AOI21_X1 U5008 ( .B1(n8691), .B2(n4582), .A(n4581), .ZN(n6217) );
  NOR2_X1 U5009 ( .A1(n4584), .A2(n4360), .ZN(n4582) );
  OAI21_X1 U5010 ( .B1(n4583), .B2(n4360), .A(n4424), .ZN(n4581) );
  NOR2_X1 U5011 ( .A1(n8852), .A2(n8707), .ZN(n4587) );
  NOR2_X1 U5012 ( .A1(n8717), .A2(n4574), .ZN(n4573) );
  INV_X1 U5013 ( .A(n8730), .ZN(n4574) );
  AND4_X1 U5015 ( .A1(n5754), .A2(n5753), .A3(n5752), .A4(n5751), .ZN(n5755)
         );
  AND2_X1 U5016 ( .A1(n5923), .A2(n5922), .ZN(n5945) );
  INV_X1 U5017 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U5018 ( .A1(n4791), .A2(n4390), .ZN(n4790) );
  NAND2_X1 U5019 ( .A1(n4792), .A2(n5311), .ZN(n4791) );
  INV_X1 U5020 ( .A(n5482), .ZN(n4769) );
  NOR2_X1 U5021 ( .A1(n5382), .A2(n5381), .ZN(n5384) );
  OAI21_X1 U5022 ( .B1(n9347), .B2(n4713), .A(n4711), .ZN(n9312) );
  INV_X1 U5023 ( .A(n4714), .ZN(n4713) );
  AOI21_X1 U5024 ( .B1(n4714), .B2(n7844), .A(n4712), .ZN(n4711) );
  INV_X1 U5025 ( .A(n7910), .ZN(n4712) );
  OAI21_X1 U5026 ( .B1(n4614), .B2(n4877), .A(n6314), .ZN(n4876) );
  INV_X1 U5027 ( .A(n4881), .ZN(n4486) );
  XNOR2_X1 U5028 ( .A(n6328), .B(n6487), .ZN(n6330) );
  AND2_X1 U5029 ( .A1(n5636), .A2(n5611), .ZN(n5633) );
  OAI21_X1 U5030 ( .B1(n5340), .B2(n4419), .A(n4457), .ZN(n5389) );
  INV_X1 U5031 ( .A(n4458), .ZN(n4457) );
  OAI21_X1 U5032 ( .B1(n5339), .B2(n4419), .A(n5366), .ZN(n4458) );
  OAI21_X1 U5033 ( .B1(n5817), .B2(n6398), .A(n4495), .ZN(n5000) );
  AND2_X1 U5034 ( .A1(n4855), .A2(n4919), .ZN(n4854) );
  OR2_X1 U5035 ( .A1(n4856), .A2(n7544), .ZN(n4855) );
  NAND2_X1 U5036 ( .A1(n7521), .A2(n7520), .ZN(n7542) );
  AOI21_X1 U5037 ( .B1(n8237), .B2(n8236), .A(n6169), .ZN(n4626) );
  NAND2_X1 U5038 ( .A1(n5792), .A2(n5791), .ZN(n6124) );
  INV_X1 U5039 ( .A(n8681), .ZN(n8090) );
  INV_X1 U5040 ( .A(n8454), .ZN(n8693) );
  INV_X1 U5041 ( .A(n8222), .ZN(n6026) );
  OAI22_X1 U5042 ( .A1(n8786), .A2(n8785), .B1(n8208), .B2(n6013), .ZN(n8778)
         );
  NAND2_X1 U5043 ( .A1(n6168), .A2(n6517), .ZN(n6922) );
  INV_X1 U5044 ( .A(n6930), .ZN(n6168) );
  OR2_X1 U5045 ( .A1(n5782), .A2(n4837), .ZN(n4579) );
  INV_X1 U5046 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6115) );
  INV_X1 U5047 ( .A(n5656), .ZN(n5630) );
  OAI21_X1 U5048 ( .B1(n7793), .B2(n7792), .A(n7791), .ZN(n7800) );
  OR2_X1 U5049 ( .A1(n4948), .A2(n4942), .ZN(n5035) );
  OR2_X1 U5050 ( .A1(n5730), .A2(n5729), .ZN(n9282) );
  AOI21_X1 U5051 ( .B1(n9301), .B2(n4504), .A(n4503), .ZN(n4502) );
  INV_X1 U5052 ( .A(n7851), .ZN(n4504) );
  INV_X1 U5053 ( .A(n7852), .ZN(n4503) );
  NAND2_X1 U5054 ( .A1(n4473), .A2(n4471), .ZN(n6304) );
  AND2_X1 U5055 ( .A1(n4472), .A2(n9489), .ZN(n4471) );
  NAND2_X1 U5056 ( .A1(n7364), .A2(n4474), .ZN(n4473) );
  NAND2_X1 U5057 ( .A1(n4474), .A2(n4477), .ZN(n4472) );
  AND2_X1 U5058 ( .A1(n4885), .A2(n6302), .ZN(n4884) );
  NAND2_X1 U5059 ( .A1(n6301), .A2(n4886), .ZN(n4885) );
  INV_X1 U5060 ( .A(n6300), .ZN(n4886) );
  INV_X1 U5061 ( .A(n7782), .ZN(n5462) );
  INV_X1 U5062 ( .A(n5083), .ZN(n7781) );
  XNOR2_X1 U5063 ( .A(n4963), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5697) );
  AND2_X1 U5064 ( .A1(n5605), .A2(n5560), .ZN(n5581) );
  NAND2_X1 U5065 ( .A1(n4514), .A2(n5133), .ZN(n5157) );
  INV_X1 U5066 ( .A(n8453), .ZN(n8668) );
  AOI21_X1 U5067 ( .B1(n4606), .B2(n4382), .A(n4598), .ZN(n4596) );
  NAND2_X1 U5068 ( .A1(n4601), .A2(n4602), .ZN(n4600) );
  INV_X1 U5069 ( .A(n7689), .ZN(n4601) );
  NAND2_X1 U5070 ( .A1(n8373), .A2(n8432), .ZN(n4521) );
  NAND2_X1 U5071 ( .A1(n4532), .A2(n4533), .ZN(n4531) );
  NAND2_X1 U5072 ( .A1(n8374), .A2(n8432), .ZN(n4533) );
  NAND2_X1 U5073 ( .A1(n8371), .A2(n8412), .ZN(n4532) );
  NAND2_X1 U5074 ( .A1(n4527), .A2(n4525), .ZN(n4524) );
  OAI21_X1 U5075 ( .B1(n8373), .B2(n4523), .A(n4522), .ZN(n4525) );
  AND2_X1 U5076 ( .A1(n8386), .A2(n8412), .ZN(n4517) );
  AOI21_X1 U5077 ( .B1(n8379), .B2(n4519), .A(n8716), .ZN(n4518) );
  NOR2_X1 U5078 ( .A1(n4520), .A2(n8412), .ZN(n4519) );
  INV_X1 U5079 ( .A(n8378), .ZN(n4520) );
  AOI21_X1 U5080 ( .B1(n7731), .B2(n7730), .A(n4611), .ZN(n4610) );
  OAI21_X1 U5081 ( .B1(n7733), .B2(n7790), .A(n9472), .ZN(n4609) );
  NAND2_X1 U5082 ( .A1(n7732), .A2(n7790), .ZN(n4611) );
  NAND2_X1 U5083 ( .A1(n4615), .A2(n4612), .ZN(n7755) );
  NOR2_X1 U5084 ( .A1(n4614), .A2(n4613), .ZN(n4612) );
  NAND2_X1 U5085 ( .A1(n9851), .A2(n9138), .ZN(n7677) );
  AND2_X1 U5086 ( .A1(n4663), .A2(n8408), .ZN(n4659) );
  NOR2_X1 U5087 ( .A1(n9592), .A2(n9481), .ZN(n4706) );
  INV_X1 U5088 ( .A(n4824), .ZN(n4823) );
  NOR2_X1 U5089 ( .A1(n4826), .A2(n5445), .ZN(n4822) );
  NAND2_X1 U5090 ( .A1(n5829), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U5091 ( .A1(n4539), .A2(n4387), .ZN(n6811) );
  NAND2_X1 U5092 ( .A1(n6764), .A2(n4540), .ZN(n4539) );
  INV_X1 U5093 ( .A(n6763), .ZN(n4540) );
  NAND2_X1 U5094 ( .A1(n6769), .A2(n4903), .ZN(n6805) );
  OR2_X1 U5095 ( .A1(n6682), .A2(n6680), .ZN(n4903) );
  NAND2_X1 U5096 ( .A1(n7257), .A2(n7258), .ZN(n7432) );
  AOI21_X1 U5097 ( .B1(n8239), .B2(n4561), .A(n4385), .ZN(n4560) );
  INV_X1 U5098 ( .A(n6101), .ZN(n4561) );
  OR2_X1 U5099 ( .A1(n6180), .A2(n9703), .ZN(n5987) );
  INV_X1 U5100 ( .A(n4637), .ZN(n4635) );
  NAND2_X1 U5101 ( .A1(n4640), .A2(n8357), .ZN(n4634) );
  NAND2_X1 U5102 ( .A1(n5965), .A2(n5964), .ZN(n5982) );
  NOR2_X1 U5103 ( .A1(n8811), .A2(n4642), .ZN(n4641) );
  INV_X1 U5104 ( .A(n8331), .ZN(n4642) );
  NAND2_X1 U5105 ( .A1(n8825), .A2(n9709), .ZN(n8340) );
  AND2_X1 U5106 ( .A1(n8316), .A2(n7388), .ZN(n8314) );
  AND2_X1 U5107 ( .A1(n8248), .A2(n8313), .ZN(n4628) );
  NAND2_X1 U5108 ( .A1(n7211), .A2(n7068), .ZN(n8280) );
  NAND2_X1 U5109 ( .A1(n8280), .A2(n8289), .ZN(n8245) );
  INV_X1 U5110 ( .A(n8269), .ZN(n7015) );
  NAND2_X1 U5111 ( .A1(n6973), .A2(n5819), .ZN(n8273) );
  INV_X1 U5112 ( .A(n8423), .ZN(n8433) );
  NAND2_X1 U5113 ( .A1(n4650), .A2(n4648), .ZN(n4647) );
  OR2_X1 U5114 ( .A1(n8895), .A2(n8693), .ZN(n8403) );
  OR2_X1 U5115 ( .A1(n8914), .A2(n8708), .ZN(n8388) );
  OR2_X1 U5116 ( .A1(n8926), .A2(n8068), .ZN(n8383) );
  OR2_X1 U5117 ( .A1(n8878), .A2(n8208), .ZN(n8368) );
  NAND2_X1 U5118 ( .A1(n6165), .A2(n6164), .ZN(n6933) );
  NOR2_X1 U5119 ( .A1(n6145), .A2(n7631), .ZN(n6164) );
  INV_X1 U5120 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6139) );
  INV_X1 U5121 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U5122 ( .A1(n5830), .A2(n5750), .ZN(n4675) );
  INV_X1 U5123 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4590) );
  AND2_X1 U5124 ( .A1(n5920), .A2(n5919), .ZN(n5923) );
  INV_X1 U5125 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5919) );
  INV_X1 U5126 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4797) );
  INV_X1 U5127 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4708) );
  INV_X1 U5128 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4795) );
  XNOR2_X1 U5129 ( .A(n7945), .B(n9126), .ZN(n7830) );
  NAND2_X1 U5130 ( .A1(n9643), .A2(n4699), .ZN(n4698) );
  INV_X1 U5131 ( .A(n9386), .ZN(n4480) );
  NOR2_X1 U5132 ( .A1(n4891), .A2(n6311), .ZN(n4890) );
  INV_X1 U5133 ( .A(n6310), .ZN(n4891) );
  AOI21_X1 U5134 ( .B1(n4733), .B2(n4731), .A(n4730), .ZN(n4729) );
  INV_X1 U5135 ( .A(n4733), .ZN(n4732) );
  INV_X1 U5136 ( .A(n9430), .ZN(n4730) );
  NOR2_X1 U5137 ( .A1(n9520), .A2(n4719), .ZN(n4718) );
  INV_X1 U5138 ( .A(n7722), .ZN(n4719) );
  INV_X1 U5139 ( .A(n4485), .ZN(n4484) );
  OAI21_X1 U5140 ( .B1(n4879), .B2(n4486), .A(n7816), .ZN(n4485) );
  NOR2_X1 U5141 ( .A1(n7814), .A2(n4880), .ZN(n4879) );
  INV_X1 U5142 ( .A(n7041), .ZN(n4880) );
  AOI21_X1 U5143 ( .B1(n7120), .B2(n4882), .A(n4389), .ZN(n4881) );
  INV_X1 U5144 ( .A(n6298), .ZN(n4882) );
  OR2_X1 U5145 ( .A1(n4690), .A2(n7510), .ZN(n4689) );
  NAND2_X1 U5146 ( .A1(n9867), .A2(n4691), .ZN(n4690) );
  NAND2_X1 U5147 ( .A1(n6540), .A2(n6635), .ZN(n6544) );
  NAND2_X1 U5148 ( .A1(n6544), .A2(n6330), .ZN(n6543) );
  AND2_X1 U5149 ( .A1(n7795), .A2(n7798), .ZN(n6325) );
  OAI21_X1 U5150 ( .B1(n7640), .B2(n10129), .A(n7639), .ZN(n7780) );
  AND2_X1 U5151 ( .A1(n5633), .A2(n5632), .ZN(n5634) );
  AND2_X1 U5152 ( .A1(n4958), .A2(n4968), .ZN(n4780) );
  AND2_X1 U5153 ( .A1(n4970), .A2(n4958), .ZN(n4973) );
  AND2_X1 U5154 ( .A1(n4814), .A2(n4455), .ZN(n4454) );
  AND2_X1 U5155 ( .A1(n4818), .A2(n4907), .ZN(n4814) );
  AOI21_X1 U5156 ( .B1(n4355), .B2(n4813), .A(n4398), .ZN(n4808) );
  OAI211_X1 U5157 ( .C1(n5157), .C2(n4722), .A(n4355), .B(n4444), .ZN(n4807)
         );
  AOI21_X1 U5158 ( .B1(n4908), .B2(n4812), .A(n4811), .ZN(n4810) );
  INV_X1 U5159 ( .A(n5226), .ZN(n4811) );
  INV_X1 U5160 ( .A(n5159), .ZN(n4804) );
  AND2_X1 U5161 ( .A1(n8124), .A2(n7997), .ZN(n8065) );
  INV_X1 U5162 ( .A(n7594), .ZN(n4856) );
  AND2_X1 U5163 ( .A1(n8076), .A2(n8000), .ZN(n8125) );
  INV_X1 U5164 ( .A(n8820), .ZN(n8339) );
  INV_X1 U5165 ( .A(n8049), .ZN(n7980) );
  INV_X1 U5166 ( .A(n6130), .ZN(n6686) );
  XNOR2_X1 U5167 ( .A(n6805), .B(n6812), .ZN(n6683) );
  NOR2_X1 U5168 ( .A1(n6683), .A2(n6684), .ZN(n6808) );
  NAND2_X1 U5169 ( .A1(n4746), .A2(n4430), .ZN(n6881) );
  NAND2_X1 U5170 ( .A1(n6881), .A2(n6880), .ZN(n4433) );
  NAND2_X1 U5171 ( .A1(n4432), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4759) );
  INV_X1 U5172 ( .A(n6882), .ZN(n4432) );
  NAND2_X1 U5173 ( .A1(n4758), .A2(n4757), .ZN(n7090) );
  INV_X1 U5174 ( .A(n6989), .ZN(n4757) );
  NAND2_X1 U5175 ( .A1(n4751), .A2(n4750), .ZN(n7243) );
  INV_X1 U5176 ( .A(n7180), .ZN(n4750) );
  AND2_X1 U5177 ( .A1(n7243), .A2(n7242), .ZN(n7425) );
  XNOR2_X1 U5178 ( .A(n7432), .B(n7426), .ZN(n7259) );
  NAND2_X1 U5179 ( .A1(n7259), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U5180 ( .A1(n4741), .A2(n4740), .ZN(n8469) );
  INV_X1 U5181 ( .A(n7430), .ZN(n4740) );
  OR2_X1 U5182 ( .A1(n8525), .A2(n8524), .ZN(n8547) );
  OR2_X1 U5183 ( .A1(n6933), .A2(n7586), .ZN(n6671) );
  OR2_X1 U5184 ( .A1(n8579), .A2(n4754), .ZN(n4752) );
  NAND2_X1 U5185 ( .A1(n4755), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4754) );
  OR2_X1 U5186 ( .A1(n4358), .A2(n8601), .ZN(n4753) );
  AND2_X1 U5187 ( .A1(n4664), .A2(n4661), .ZN(n4660) );
  NAND2_X1 U5188 ( .A1(n4671), .A2(n4670), .ZN(n4669) );
  AOI21_X1 U5189 ( .B1(n4586), .B2(n6068), .A(n4400), .ZN(n4583) );
  AND2_X1 U5190 ( .A1(n8407), .A2(n8408), .ZN(n8669) );
  INV_X1 U5191 ( .A(n4647), .ZN(n4646) );
  NAND2_X1 U5192 ( .A1(n5779), .A2(n5778), .ZN(n6058) );
  NAND2_X1 U5193 ( .A1(n8351), .A2(n8348), .ZN(n8802) );
  INV_X1 U5194 ( .A(n4641), .ZN(n4640) );
  AOI21_X1 U5195 ( .B1(n4641), .B2(n4639), .A(n4638), .ZN(n4637) );
  INV_X1 U5196 ( .A(n8358), .ZN(n4638) );
  INV_X1 U5197 ( .A(n8256), .ZN(n4639) );
  NAND2_X1 U5198 ( .A1(n7559), .A2(n8256), .ZN(n7558) );
  AND4_X1 U5199 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n7607)
         );
  NOR2_X1 U5200 ( .A1(n4593), .A2(n4592), .ZN(n4591) );
  INV_X1 U5201 ( .A(n5908), .ZN(n4592) );
  AND2_X1 U5202 ( .A1(n4593), .A2(n8317), .ZN(n4674) );
  NAND2_X1 U5203 ( .A1(n7268), .A2(n4594), .ZN(n7390) );
  AND2_X1 U5204 ( .A1(n8251), .A2(n5898), .ZN(n4594) );
  OAI22_X1 U5205 ( .A1(n7281), .A2(n5873), .B1(n8463), .B2(n7239), .ZN(n7318)
         );
  XNOR2_X1 U5206 ( .A(n8464), .B(n8306), .ZN(n8287) );
  AND2_X1 U5207 ( .A1(n7139), .A2(n5836), .ZN(n5835) );
  OR2_X1 U5208 ( .A1(n5837), .A2(n6176), .ZN(n6844) );
  INV_X1 U5209 ( .A(n8466), .ZN(n6969) );
  AND2_X1 U5210 ( .A1(n4673), .A2(n4672), .ZN(n6236) );
  NAND2_X1 U5211 ( .A1(n4666), .A2(n4664), .ZN(n4673) );
  AND2_X1 U5212 ( .A1(n8403), .A2(n8404), .ZN(n8686) );
  INV_X1 U5213 ( .A(n4587), .ZN(n4585) );
  AOI21_X1 U5214 ( .B1(n4571), .B2(n4569), .A(n4391), .ZN(n4568) );
  INV_X1 U5215 ( .A(n4573), .ZN(n4569) );
  INV_X1 U5216 ( .A(n4571), .ZN(n4570) );
  NAND2_X1 U5217 ( .A1(n8432), .A2(n7023), .ZN(n9710) );
  AOI21_X1 U5218 ( .B1(n4652), .B2(n4655), .A(n4651), .ZN(n4650) );
  INV_X1 U5219 ( .A(n8388), .ZN(n4651) );
  NAND2_X1 U5220 ( .A1(n8727), .A2(n4652), .ZN(n4649) );
  AOI21_X1 U5221 ( .B1(n8731), .B2(n4572), .A(n4654), .ZN(n4571) );
  INV_X1 U5222 ( .A(n8717), .ZN(n4572) );
  NAND2_X1 U5223 ( .A1(n8741), .A2(n4573), .ZN(n4567) );
  INV_X1 U5224 ( .A(n8386), .ZN(n4655) );
  AOI21_X1 U5225 ( .B1(n8741), .B2(n8730), .A(n8731), .ZN(n8729) );
  INV_X1 U5226 ( .A(n4575), .ZN(n8743) );
  NAND2_X1 U5227 ( .A1(n8932), .A2(n8769), .ZN(n4576) );
  NOR2_X1 U5228 ( .A1(n8932), .A2(n8769), .ZN(n4577) );
  AND2_X1 U5229 ( .A1(n8945), .A2(n8768), .ZN(n6023) );
  OR2_X1 U5230 ( .A1(n8945), .A2(n8788), .ZN(n8761) );
  INV_X1 U5231 ( .A(n9710), .ZN(n8822) );
  NAND2_X1 U5232 ( .A1(n4534), .A2(n5992), .ZN(n9719) );
  NAND2_X1 U5233 ( .A1(n6827), .A2(n8224), .ZN(n4534) );
  AND2_X1 U5234 ( .A1(n5926), .A2(n5925), .ZN(n9919) );
  NAND2_X1 U5235 ( .A1(n6267), .A2(n9892), .ZN(n9933) );
  NAND2_X1 U5236 ( .A1(n6150), .A2(n6149), .ZN(n6259) );
  INV_X1 U5237 ( .A(n4834), .ZN(n4833) );
  INV_X1 U5238 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6134) );
  INV_X1 U5239 ( .A(n4836), .ZN(n4835) );
  OAI21_X1 U5240 ( .B1(n6167), .B2(n4837), .A(n6139), .ZN(n4836) );
  NOR2_X1 U5241 ( .A1(n6139), .A2(n4837), .ZN(n4834) );
  AND2_X1 U5242 ( .A1(n5799), .A2(n6115), .ZN(n4870) );
  NAND2_X1 U5243 ( .A1(n5798), .A2(n4372), .ZN(n6121) );
  INV_X1 U5244 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5799) );
  INV_X1 U5245 ( .A(n8975), .ZN(n4789) );
  NAND2_X1 U5246 ( .A1(n4782), .A2(n4787), .ZN(n4783) );
  AND2_X1 U5247 ( .A1(n5683), .A2(n5682), .ZN(n6204) );
  NOR2_X1 U5248 ( .A1(n4766), .A2(n4356), .ZN(n4763) );
  OAI21_X1 U5249 ( .B1(n4765), .B2(n4356), .A(n4393), .ZN(n4762) );
  NAND2_X1 U5250 ( .A1(n9113), .A2(n5385), .ZN(n9025) );
  OR2_X1 U5251 ( .A1(n5327), .A2(n5326), .ZN(n5351) );
  AND2_X1 U5252 ( .A1(n5473), .A2(n5472), .ZN(n5478) );
  INV_X1 U5253 ( .A(n5118), .ZN(n4778) );
  NAND2_X1 U5254 ( .A1(n9112), .A2(n9114), .ZN(n9113) );
  NOR2_X1 U5255 ( .A1(n5720), .A2(n7936), .ZN(n5725) );
  NAND2_X1 U5256 ( .A1(n7865), .A2(n7866), .ZN(n4621) );
  INV_X1 U5257 ( .A(n4622), .ZN(n4460) );
  NAND2_X1 U5258 ( .A1(n7927), .A2(n5718), .ZN(n7928) );
  OR2_X1 U5259 ( .A1(n5471), .A2(n4949), .ZN(n4950) );
  INV_X1 U5260 ( .A(n7651), .ZN(n5037) );
  AND4_X1 U5261 ( .A1(n4927), .A2(n4926), .A3(n4925), .A4(n4924), .ZN(n4928)
         );
  AND2_X1 U5262 ( .A1(n9331), .A2(n4694), .ZN(n9275) );
  NOR2_X1 U5263 ( .A1(n4695), .A2(n7945), .ZN(n4694) );
  INV_X1 U5264 ( .A(n4697), .ZN(n4695) );
  AND2_X1 U5265 ( .A1(n5731), .A2(n9282), .ZN(n9293) );
  NAND2_X1 U5266 ( .A1(n4487), .A2(n4386), .ZN(n4873) );
  AND2_X1 U5267 ( .A1(n5676), .A2(n5675), .ZN(n9304) );
  NAND2_X1 U5268 ( .A1(n9329), .A2(n9330), .ZN(n4487) );
  NAND2_X1 U5269 ( .A1(n9347), .A2(n7760), .ZN(n4710) );
  AND2_X1 U5270 ( .A1(n9338), .A2(n4715), .ZN(n4714) );
  NAND2_X1 U5271 ( .A1(n9346), .A2(n7760), .ZN(n4715) );
  NAND2_X1 U5272 ( .A1(n9363), .A2(n7834), .ZN(n9347) );
  NAND2_X1 U5273 ( .A1(n4717), .A2(n4716), .ZN(n9349) );
  INV_X1 U5274 ( .A(n9346), .ZN(n4716) );
  INV_X1 U5275 ( .A(n9347), .ZN(n4717) );
  OAI21_X1 U5276 ( .B1(n6345), .B2(n4508), .A(n4506), .ZN(n9404) );
  INV_X1 U5277 ( .A(n4507), .ZN(n4506) );
  OAI21_X1 U5278 ( .B1(n4368), .B2(n4508), .A(n9406), .ZN(n4507) );
  INV_X1 U5279 ( .A(n7749), .ZN(n4508) );
  AND2_X1 U5280 ( .A1(n7661), .A2(n7662), .ZN(n9406) );
  NAND2_X1 U5281 ( .A1(n6345), .A2(n4368), .ZN(n9417) );
  OAI21_X1 U5282 ( .B1(n6304), .B2(n4898), .A(n4895), .ZN(n9442) );
  NAND2_X1 U5283 ( .A1(n4357), .A2(n4901), .ZN(n4898) );
  AOI21_X1 U5284 ( .B1(n4357), .B2(n4896), .A(n4374), .ZN(n4895) );
  OAI21_X1 U5285 ( .B1(n9471), .B2(n7734), .A(n7735), .ZN(n9457) );
  NOR2_X1 U5286 ( .A1(n6305), .A2(n4900), .ZN(n4899) );
  INV_X1 U5287 ( .A(n6303), .ZN(n4900) );
  OR2_X1 U5288 ( .A1(n9481), .A2(n9501), .ZN(n4901) );
  AOI21_X1 U5289 ( .B1(n4475), .B2(n4476), .A(n4422), .ZN(n4474) );
  INV_X1 U5290 ( .A(n4883), .ZN(n4475) );
  NOR2_X1 U5291 ( .A1(n4887), .A2(n7820), .ZN(n4883) );
  INV_X1 U5292 ( .A(n6301), .ZN(n4887) );
  OR2_X1 U5293 ( .A1(n7486), .A2(n7229), .ZN(n7721) );
  NAND2_X1 U5294 ( .A1(n6343), .A2(n4371), .ZN(n7473) );
  NAND2_X1 U5295 ( .A1(n7364), .A2(n7363), .ZN(n7362) );
  OR2_X1 U5296 ( .A1(n7510), .A2(n7411), .ZN(n7709) );
  NAND2_X1 U5297 ( .A1(n7709), .A2(n7710), .ZN(n7816) );
  NAND2_X1 U5298 ( .A1(n7042), .A2(n7041), .ZN(n7040) );
  NOR2_X2 U5299 ( .A1(n7861), .A2(n6466), .ZN(n9500) );
  INV_X1 U5300 ( .A(n9142), .ZN(n6536) );
  INV_X1 U5301 ( .A(n9500), .ZN(n9516) );
  AND2_X1 U5302 ( .A1(n6325), .A2(n5718), .ZN(n9531) );
  NAND2_X1 U5303 ( .A1(n5670), .A2(n5669), .ZN(n9322) );
  NAND2_X1 U5304 ( .A1(n5562), .A2(n5561), .ZN(n9388) );
  NAND2_X1 U5305 ( .A1(n5512), .A2(n5511), .ZN(n9422) );
  NAND2_X1 U5306 ( .A1(n5397), .A2(n5396), .ZN(n9601) );
  NAND2_X1 U5307 ( .A1(n5348), .A2(n5347), .ZN(n9611) );
  AND2_X1 U5308 ( .A1(n6325), .A2(n7929), .ZN(n9623) );
  AND2_X1 U5309 ( .A1(n5695), .A2(n5697), .ZN(n6416) );
  NOR2_X1 U5310 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4624) );
  NAND2_X1 U5311 ( .A1(n4451), .A2(n6105), .ZN(n6229) );
  NOR2_X1 U5312 ( .A1(n4936), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n4893) );
  XNOR2_X1 U5313 ( .A(n5612), .B(n5633), .ZN(n7626) );
  XNOR2_X1 U5314 ( .A(n5587), .B(n5586), .ZN(n7589) );
  OAI21_X1 U5315 ( .B1(n5535), .B2(n5534), .A(n5533), .ZN(n5556) );
  INV_X1 U5316 ( .A(n5531), .ZN(n5532) );
  NAND2_X1 U5317 ( .A1(n4984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U5318 ( .A1(n4985), .A2(n4959), .ZN(n5710) );
  OAI21_X1 U5319 ( .B1(n5484), .B2(n5485), .A(n5486), .ZN(n5507) );
  INV_X1 U5320 ( .A(n4820), .ZN(n5459) );
  AOI21_X1 U5321 ( .B1(n5418), .B2(n4826), .A(n4824), .ZN(n4820) );
  OAI21_X1 U5322 ( .B1(n5418), .B2(n5417), .A(n5416), .ZN(n5441) );
  OAI21_X1 U5323 ( .B1(n5157), .B2(n4722), .A(n4720), .ZN(n5225) );
  AOI21_X1 U5324 ( .B1(n4721), .B2(n4801), .A(n4812), .ZN(n4720) );
  NOR2_X1 U5325 ( .A1(n4803), .A2(n5201), .ZN(n4721) );
  NAND2_X1 U5326 ( .A1(n4494), .A2(n5113), .ZN(n5131) );
  NAND2_X1 U5327 ( .A1(n4440), .A2(n4491), .ZN(n4439) );
  NAND2_X1 U5328 ( .A1(n4491), .A2(n5004), .ZN(n5081) );
  NAND2_X1 U5329 ( .A1(n4492), .A2(n5001), .ZN(n5062) );
  OR2_X1 U5330 ( .A1(n6405), .A2(n5827), .ZN(n5896) );
  INV_X1 U5331 ( .A(n8680), .ZN(n8707) );
  AND3_X1 U5332 ( .A1(n5790), .A2(n5789), .A3(n5788), .ZN(n8694) );
  AOI21_X1 U5333 ( .B1(n8196), .B2(n4564), .A(n4563), .ZN(n7025) );
  AND2_X1 U5334 ( .A1(n8205), .A2(n5819), .ZN(n4563) );
  AND2_X1 U5335 ( .A1(n6926), .A2(n6925), .ZN(n8199) );
  INV_X1 U5336 ( .A(n6686), .ZN(n8444) );
  OR2_X1 U5337 ( .A1(n4626), .A2(n4625), .ZN(n4536) );
  OR2_X1 U5338 ( .A1(n8424), .A2(n4799), .ZN(n4798) );
  XNOR2_X1 U5339 ( .A(n6118), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U5340 ( .A1(n6117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U5341 ( .A1(n6099), .A2(n6098), .ZN(n8453) );
  NAND2_X1 U5342 ( .A1(n6089), .A2(n6088), .ZN(n8681) );
  NAND2_X1 U5343 ( .A1(n6078), .A2(n6077), .ZN(n8454) );
  INV_X1 U5344 ( .A(n8694), .ZN(n8720) );
  NAND2_X1 U5345 ( .A1(n4548), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5346 ( .A1(n8630), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4547) );
  NAND2_X1 U5347 ( .A1(n4544), .A2(n4543), .ZN(n4542) );
  INV_X1 U5348 ( .A(n8639), .ZN(n4543) );
  NAND2_X1 U5349 ( .A1(n8640), .A2(n9883), .ZN(n4544) );
  AOI21_X1 U5350 ( .B1(n8657), .B2(n7282), .A(n6242), .ZN(n6243) );
  NAND2_X1 U5351 ( .A1(n8418), .A2(n8239), .ZN(n4559) );
  NAND2_X1 U5352 ( .A1(n5765), .A2(n5764), .ZN(n8712) );
  OR2_X1 U5353 ( .A1(n6275), .A2(n8952), .ZN(n6189) );
  NOR2_X1 U5354 ( .A1(n4681), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4680) );
  NAND2_X1 U5355 ( .A1(n4683), .A2(n4682), .ZN(n4681) );
  INV_X1 U5356 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4682) );
  AND2_X1 U5357 ( .A1(n5697), .A2(n4966), .ZN(n4967) );
  XNOR2_X1 U5358 ( .A(n5711), .B(n4960), .ZN(n6408) );
  NAND2_X1 U5359 ( .A1(n5710), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5711) );
  INV_X1 U5360 ( .A(n7867), .ZN(n7925) );
  INV_X1 U5361 ( .A(n9304), .ZN(n9340) );
  NAND2_X1 U5362 ( .A1(n5625), .A2(n5624), .ZN(n9339) );
  NAND2_X1 U5363 ( .A1(n5570), .A2(n5569), .ZN(n9408) );
  INV_X1 U5364 ( .A(n7229), .ZN(n9133) );
  NOR2_X1 U5365 ( .A1(n4909), .A2(n4910), .ZN(n5060) );
  NAND2_X1 U5366 ( .A1(n7651), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U5367 ( .A1(n5073), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5020) );
  OAI211_X1 U5368 ( .C1(n9311), .C2(n4501), .A(n4500), .B(n4498), .ZN(n6354)
         );
  NAND2_X1 U5369 ( .A1(n7778), .A2(n9301), .ZN(n4501) );
  AND2_X1 U5370 ( .A1(n4465), .A2(n7650), .ZN(n9638) );
  NAND2_X1 U5371 ( .A1(n8954), .A2(n7781), .ZN(n4465) );
  NOR2_X1 U5372 ( .A1(n6369), .A2(n9866), .ZN(n6572) );
  NAND2_X1 U5373 ( .A1(n6355), .A2(n9871), .ZN(n4739) );
  NAND2_X1 U5374 ( .A1(n4738), .A2(n4361), .ZN(n4489) );
  INV_X1 U5375 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9682) );
  AND2_X1 U5376 ( .A1(n7885), .A2(n7709), .ZN(n4608) );
  INV_X1 U5377 ( .A(n4596), .ZN(n4595) );
  INV_X1 U5378 ( .A(n4530), .ZN(n4523) );
  AOI21_X1 U5379 ( .B1(n4530), .B2(n8412), .A(n8381), .ZN(n4522) );
  AND2_X1 U5380 ( .A1(n4528), .A2(n8380), .ZN(n4527) );
  NAND2_X1 U5381 ( .A1(n4521), .A2(n4530), .ZN(n4526) );
  NAND2_X1 U5382 ( .A1(n4515), .A2(n8390), .ZN(n8397) );
  NAND2_X1 U5383 ( .A1(n4518), .A2(n4516), .ZN(n4515) );
  NAND2_X1 U5384 ( .A1(n8387), .A2(n4517), .ZN(n4516) );
  NAND2_X1 U5385 ( .A1(n7740), .A2(n4620), .ZN(n4619) );
  AND2_X1 U5386 ( .A1(n7746), .A2(n7786), .ZN(n4620) );
  INV_X1 U5387 ( .A(n7752), .ZN(n4613) );
  NAND2_X1 U5388 ( .A1(n7678), .A2(n7706), .ZN(n7697) );
  NAND2_X1 U5389 ( .A1(n8417), .A2(n4537), .ZN(n8428) );
  AND2_X1 U5390 ( .A1(n4806), .A2(n8416), .ZN(n4537) );
  AND2_X1 U5391 ( .A1(n5761), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5760) );
  INV_X1 U5392 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5745) );
  NOR2_X1 U5393 ( .A1(n7831), .A2(n4463), .ZN(n7869) );
  INV_X1 U5394 ( .A(n4735), .ZN(n4731) );
  NAND2_X1 U5395 ( .A1(n4828), .A2(n5416), .ZN(n4827) );
  INV_X1 U5396 ( .A(n5440), .ZN(n4828) );
  NAND2_X1 U5397 ( .A1(n4723), .A2(n4461), .ZN(n4444) );
  INV_X1 U5398 ( .A(SI_17_), .ZN(n10041) );
  INV_X1 U5399 ( .A(n8008), .ZN(n4859) );
  INV_X1 U5400 ( .A(n8189), .ZN(n4849) );
  NAND2_X1 U5401 ( .A1(n8428), .A2(n4805), .ZN(n8420) );
  NAND2_X1 U5402 ( .A1(n4806), .A2(n8426), .ZN(n4805) );
  INV_X1 U5403 ( .A(n8420), .ZN(n8436) );
  NAND2_X1 U5404 ( .A1(n4658), .A2(n4663), .ZN(n4657) );
  INV_X1 U5405 ( .A(n4660), .ZN(n4658) );
  NAND2_X1 U5406 ( .A1(n8530), .A2(n8531), .ZN(n8553) );
  OR2_X1 U5407 ( .A1(n6147), .A2(n6162), .ZN(n6247) );
  AND2_X1 U5408 ( .A1(n8938), .A2(n7991), .ZN(n8763) );
  NAND2_X1 U5409 ( .A1(n9719), .A2(n9711), .ZN(n8348) );
  OR2_X1 U5410 ( .A1(n6940), .A2(n6939), .ZN(n6927) );
  AND2_X1 U5411 ( .A1(n8448), .A2(n8443), .ZN(n6170) );
  NAND2_X1 U5412 ( .A1(n5759), .A2(n5781), .ZN(n4684) );
  INV_X1 U5413 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5781) );
  OR2_X1 U5414 ( .A1(n5953), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5946) );
  INV_X1 U5415 ( .A(n9080), .ZN(n4786) );
  NOR2_X1 U5416 ( .A1(n9284), .A2(n4698), .ZN(n4697) );
  NOR2_X1 U5417 ( .A1(n9560), .A2(n4703), .ZN(n4702) );
  INV_X1 U5418 ( .A(n4704), .ZN(n4703) );
  NOR2_X1 U5419 ( .A1(n9388), .A2(n9571), .ZN(n4704) );
  NAND2_X1 U5420 ( .A1(n5513), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5542) );
  NOR2_X1 U5421 ( .A1(n9443), .A2(n4736), .ZN(n4735) );
  INV_X1 U5422 ( .A(n7742), .ZN(n4736) );
  AOI21_X1 U5423 ( .B1(n4735), .B2(n7801), .A(n4734), .ZN(n4733) );
  INV_X1 U5424 ( .A(n7744), .ZN(n4734) );
  NOR2_X1 U5425 ( .A1(n4899), .A2(n4897), .ZN(n4896) );
  INV_X1 U5426 ( .A(n4901), .ZN(n4897) );
  NAND2_X1 U5427 ( .A1(n6536), .A2(n9824), .ZN(n6601) );
  NAND2_X1 U5428 ( .A1(n9490), .A2(n4705), .ZN(n9434) );
  AND2_X1 U5429 ( .A1(n9439), .A2(n4363), .ZN(n4705) );
  NAND2_X1 U5430 ( .A1(n9490), .A2(n4706), .ZN(n9460) );
  NAND2_X1 U5431 ( .A1(n9490), .A2(n9664), .ZN(n9478) );
  NOR2_X1 U5432 ( .A1(n6647), .A2(n6648), .ZN(n6746) );
  NOR2_X1 U5433 ( .A1(n6397), .A2(n6388), .ZN(n4686) );
  AND2_X1 U5434 ( .A1(n5664), .A2(n5640), .ZN(n5662) );
  NAND2_X1 U5435 ( .A1(n5607), .A2(n5606), .ZN(n5635) );
  NAND2_X1 U5436 ( .A1(n4469), .A2(n4467), .ZN(n5607) );
  AND2_X1 U5437 ( .A1(n4468), .A2(n5581), .ZN(n4467) );
  NAND2_X1 U5438 ( .A1(n5556), .A2(n5554), .ZN(n4469) );
  NAND2_X1 U5439 ( .A1(n5555), .A2(n5554), .ZN(n4468) );
  AOI21_X1 U5440 ( .B1(n4823), .B2(n4822), .A(n4426), .ZN(n4821) );
  INV_X1 U5441 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4978) );
  OAI21_X1 U5442 ( .B1(n4827), .B2(n4825), .A(n5439), .ZN(n4824) );
  INV_X1 U5443 ( .A(n5417), .ZN(n4825) );
  INV_X1 U5444 ( .A(n4827), .ZN(n4826) );
  NAND2_X1 U5445 ( .A1(n4931), .A2(n4930), .ZN(n5394) );
  INV_X1 U5446 ( .A(n5286), .ZN(n4818) );
  INV_X1 U5447 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4923) );
  OAI21_X1 U5448 ( .B1(n6389), .B2(n5006), .A(n5005), .ZN(n5008) );
  NAND2_X1 U5449 ( .A1(n6389), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U5450 ( .A1(n5817), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4496) );
  INV_X1 U5451 ( .A(SI_8_), .ZN(n10143) );
  INV_X1 U5452 ( .A(SI_28_), .ZN(n10071) );
  INV_X1 U5453 ( .A(SI_29_), .ZN(n10129) );
  INV_X1 U5454 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10062) );
  INV_X1 U5455 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10060) );
  NOR2_X1 U5456 ( .A1(n7460), .A2(n4862), .ZN(n4861) );
  INV_X1 U5457 ( .A(n4863), .ZN(n4862) );
  INV_X1 U5458 ( .A(n4847), .ZN(n4846) );
  OAI21_X1 U5459 ( .B1(n8038), .B2(n4848), .A(n8028), .ZN(n4847) );
  OR2_X1 U5460 ( .A1(n8027), .A2(n8668), .ZN(n8028) );
  NAND2_X1 U5461 ( .A1(n8190), .A2(n4849), .ZN(n4848) );
  OR2_X1 U5462 ( .A1(n8038), .A2(n4851), .ZN(n4850) );
  INV_X1 U5463 ( .A(n8190), .ZN(n4851) );
  INV_X1 U5464 ( .A(n8030), .ZN(n4844) );
  NAND2_X1 U5465 ( .A1(n7595), .A2(n7594), .ZN(n8157) );
  XNOR2_X1 U5466 ( .A(n7020), .B(n5820), .ZN(n7022) );
  AND2_X1 U5467 ( .A1(n8063), .A2(n7994), .ZN(n8176) );
  XNOR2_X1 U5468 ( .A(n8626), .B(n8445), .ZN(n7023) );
  NAND2_X1 U5469 ( .A1(n8429), .A2(n4800), .ZN(n4799) );
  INV_X1 U5470 ( .A(n8430), .ZN(n4800) );
  AND2_X1 U5471 ( .A1(n8265), .A2(n8437), .ZN(n4625) );
  AND2_X1 U5472 ( .A1(n8235), .A2(n6240), .ZN(n8228) );
  AND4_X1 U5473 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n8068)
         );
  INV_X1 U5474 ( .A(n5839), .ZN(n6029) );
  OAI21_X1 U5475 ( .B1(n6676), .B2(n6732), .A(n6677), .ZN(n6728) );
  NAND2_X1 U5476 ( .A1(n4760), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6730) );
  INV_X1 U5477 ( .A(n6728), .ZN(n4760) );
  NAND2_X1 U5478 ( .A1(n5829), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6689) );
  INV_X1 U5479 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10165) );
  OAI21_X1 U5480 ( .B1(n6784), .B2(n6694), .A(n4541), .ZN(n6764) );
  OR2_X1 U5481 ( .A1(n6693), .A2(n6792), .ZN(n4541) );
  XNOR2_X1 U5482 ( .A(n6811), .B(n6807), .ZN(n6696) );
  INV_X1 U5483 ( .A(n6805), .ZN(n6806) );
  INV_X1 U5484 ( .A(n4433), .ZN(n6984) );
  OR2_X1 U5485 ( .A1(n7176), .A2(n7177), .ZN(n4751) );
  OR2_X1 U5486 ( .A1(n7428), .A2(n7427), .ZN(n4741) );
  NAND2_X1 U5487 ( .A1(n7434), .A2(n7435), .ZN(n7437) );
  INV_X1 U5488 ( .A(n8498), .ZN(n4749) );
  NAND2_X1 U5489 ( .A1(n8510), .A2(n8511), .ZN(n8512) );
  NAND2_X1 U5490 ( .A1(n8512), .A2(n8513), .ZN(n8530) );
  XNOR2_X1 U5491 ( .A(n8553), .B(n8565), .ZN(n8532) );
  INV_X1 U5492 ( .A(n8552), .ZN(n4745) );
  INV_X1 U5493 ( .A(n8547), .ZN(n8548) );
  NAND2_X1 U5494 ( .A1(n8556), .A2(n8557), .ZN(n8581) );
  XNOR2_X1 U5495 ( .A(n8610), .B(n8605), .ZN(n8583) );
  NAND2_X1 U5496 ( .A1(n8581), .A2(n4538), .ZN(n8610) );
  OR2_X1 U5497 ( .A1(n8582), .A2(n8879), .ZN(n4538) );
  NAND2_X1 U5498 ( .A1(n8583), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8612) );
  OR2_X1 U5499 ( .A1(n8579), .A2(n8580), .ZN(n4756) );
  NOR2_X1 U5500 ( .A1(n8418), .A2(n4556), .ZN(n4555) );
  INV_X1 U5501 ( .A(n4560), .ZN(n4556) );
  OAI21_X1 U5502 ( .B1(n8418), .B2(n4376), .A(n4558), .ZN(n4557) );
  NAND2_X1 U5503 ( .A1(n8418), .A2(n4560), .ZN(n4558) );
  OR2_X1 U5504 ( .A1(n6092), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6110) );
  OR2_X1 U5505 ( .A1(n6058), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6064) );
  OR2_X1 U5506 ( .A1(n6046), .A2(n5777), .ZN(n6056) );
  NAND2_X1 U5507 ( .A1(n5776), .A2(n10060), .ZN(n6046) );
  INV_X1 U5508 ( .A(n6032), .ZN(n5776) );
  NAND2_X1 U5509 ( .A1(n5775), .A2(n10062), .ZN(n6030) );
  INV_X1 U5510 ( .A(n6017), .ZN(n5775) );
  OR2_X1 U5511 ( .A1(n6030), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6032) );
  INV_X1 U5512 ( .A(n5993), .ZN(n5774) );
  OR2_X1 U5513 ( .A1(n6007), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6017) );
  OR2_X1 U5514 ( .A1(n5975), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5993) );
  INV_X1 U5515 ( .A(n4633), .ZN(n4632) );
  OAI21_X1 U5516 ( .B1(n4635), .B2(n4634), .A(n8340), .ZN(n4633) );
  INV_X1 U5517 ( .A(n5982), .ZN(n5983) );
  OR2_X1 U5518 ( .A1(n5938), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5956) );
  INV_X1 U5519 ( .A(n8821), .ZN(n8167) );
  OR2_X1 U5520 ( .A1(n5927), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5938) );
  OR2_X1 U5521 ( .A1(n5899), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5909) );
  INV_X1 U5522 ( .A(n4630), .ZN(n4629) );
  OAI21_X1 U5523 ( .B1(n8311), .B2(n4631), .A(n8314), .ZN(n4630) );
  OR2_X1 U5524 ( .A1(n5874), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5886) );
  AND2_X1 U5525 ( .A1(n8290), .A2(n8307), .ZN(n8248) );
  NAND2_X1 U5526 ( .A1(n6969), .A2(n7021), .ZN(n8270) );
  NAND2_X1 U5527 ( .A1(n6263), .A2(n6262), .ZN(n6268) );
  AND2_X1 U5528 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  NAND2_X1 U5529 ( .A1(n4644), .A2(n4643), .ZN(n8687) );
  AOI21_X1 U5530 ( .B1(n4645), .B2(n4647), .A(n8399), .ZN(n4643) );
  AOI21_X1 U5531 ( .B1(n4646), .B2(n4653), .A(n8396), .ZN(n4645) );
  NAND2_X1 U5532 ( .A1(n8766), .A2(n4902), .ZN(n4578) );
  OR2_X1 U5533 ( .A1(n8188), .A2(n7991), .ZN(n4902) );
  OR2_X1 U5534 ( .A1(n8381), .A2(n8241), .ZN(n8753) );
  INV_X1 U5535 ( .A(n8366), .ZN(n8777) );
  AND2_X1 U5536 ( .A1(n8368), .A2(n8367), .ZN(n8785) );
  AND2_X2 U5537 ( .A1(n5833), .A2(n4359), .ZN(n9891) );
  OR2_X1 U5538 ( .A1(n8222), .A2(n5828), .ZN(n5833) );
  INV_X1 U5539 ( .A(n9907), .ZN(n9892) );
  INV_X1 U5540 ( .A(n6927), .ZN(n6924) );
  OR2_X1 U5541 ( .A1(n7017), .A2(n8412), .ZN(n6978) );
  NAND2_X1 U5542 ( .A1(n6933), .A2(n6580), .ZN(n6939) );
  XNOR2_X1 U5543 ( .A(n6166), .B(n6167), .ZN(n6932) );
  INV_X1 U5544 ( .A(n4684), .ZN(n4683) );
  XNOR2_X1 U5545 ( .A(n6143), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6146) );
  NOR2_X1 U5546 ( .A1(n5924), .A2(n5945), .ZN(n7196) );
  NOR2_X1 U5547 ( .A1(n4678), .A2(n4679), .ZN(n5869) );
  NAND2_X1 U5548 ( .A1(n5830), .A2(n5743), .ZN(n4678) );
  INV_X1 U5549 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5744) );
  XNOR2_X1 U5550 ( .A(n5660), .B(n5658), .ZN(n9017) );
  INV_X1 U5551 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5401) );
  OR2_X1 U5552 ( .A1(n5402), .A2(n5401), .ZN(n5427) );
  NAND2_X1 U5553 ( .A1(n4450), .A2(n9047), .ZN(n9046) );
  NAND2_X1 U5554 ( .A1(n4404), .A2(n4769), .ZN(n4765) );
  OR2_X1 U5555 ( .A1(n9038), .A2(n4768), .ZN(n4767) );
  NAND2_X1 U5556 ( .A1(n4769), .A2(n5438), .ZN(n4766) );
  INV_X1 U5557 ( .A(n7479), .ZN(n4446) );
  NAND2_X1 U5558 ( .A1(n5312), .A2(n4448), .ZN(n4447) );
  INV_X1 U5559 ( .A(n7406), .ZN(n4448) );
  NAND2_X1 U5560 ( .A1(n7405), .A2(n7406), .ZN(n7404) );
  NAND2_X1 U5561 ( .A1(n4785), .A2(n4786), .ZN(n8985) );
  INV_X1 U5562 ( .A(n9078), .ZN(n4785) );
  OAI22_X1 U5563 ( .A1(n6535), .A2(n5656), .B1(n6328), .B2(n5086), .ZN(n5034)
         );
  XNOR2_X1 U5564 ( .A(n5031), .B(n5628), .ZN(n5054) );
  NAND2_X1 U5565 ( .A1(n9837), .A2(n5045), .ZN(n5029) );
  XNOR2_X1 U5566 ( .A(n5070), .B(n5628), .ZN(n5072) );
  NAND2_X1 U5567 ( .A1(n5425), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5465) );
  INV_X1 U5568 ( .A(n5427), .ZN(n5425) );
  INV_X1 U5569 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9092) );
  INV_X1 U5570 ( .A(n6832), .ZN(n4775) );
  AND2_X1 U5571 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  NAND2_X1 U5572 ( .A1(n5372), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5402) );
  INV_X1 U5573 ( .A(n5374), .ZN(n5372) );
  AND2_X1 U5574 ( .A1(n9638), .A2(n9125), .ZN(n7867) );
  AND2_X1 U5575 ( .A1(n5302), .A2(n5301), .ZN(n7328) );
  AND2_X1 U5576 ( .A1(n5264), .A2(n5263), .ZN(n7380) );
  AND2_X1 U5577 ( .A1(n5215), .A2(n5214), .ZN(n6952) );
  AND2_X1 U5578 ( .A1(n5155), .A2(n5154), .ZN(n6740) );
  AND2_X1 U5579 ( .A1(n5106), .A2(n5105), .ZN(n6739) );
  INV_X1 U5580 ( .A(n4698), .ZN(n4696) );
  OAI21_X1 U5581 ( .B1(n7778), .B2(n4383), .A(n4499), .ZN(n4498) );
  NAND2_X1 U5582 ( .A1(n9300), .A2(n9301), .ZN(n9299) );
  AND2_X1 U5583 ( .A1(n5736), .A2(n5735), .ZN(n9315) );
  AND2_X1 U5584 ( .A1(n7916), .A2(n7851), .ZN(n9313) );
  NAND2_X1 U5585 ( .A1(n9398), .A2(n4700), .ZN(n9353) );
  AND2_X1 U5586 ( .A1(n4702), .A2(n4701), .ZN(n4700) );
  INV_X1 U5587 ( .A(n4876), .ZN(n4875) );
  AND2_X1 U5588 ( .A1(n5652), .A2(n5651), .ZN(n9350) );
  OR2_X1 U5589 ( .A1(n9332), .A2(n5057), .ZN(n5652) );
  NAND2_X1 U5590 ( .A1(n9398), .A2(n4702), .ZN(n9369) );
  NAND2_X1 U5591 ( .A1(n9378), .A2(n9387), .ZN(n9377) );
  NAND2_X1 U5592 ( .A1(n9377), .A2(n4513), .ZN(n9363) );
  AND2_X1 U5593 ( .A1(n9368), .A2(n9362), .ZN(n4513) );
  AND2_X1 U5594 ( .A1(n7751), .A2(n9362), .ZN(n9387) );
  AOI21_X1 U5595 ( .B1(n4890), .B2(n4418), .A(n4362), .ZN(n4889) );
  NAND2_X1 U5596 ( .A1(n9413), .A2(n4890), .ZN(n4888) );
  NAND2_X1 U5597 ( .A1(n9398), .A2(n9403), .ZN(n9399) );
  NAND2_X1 U5598 ( .A1(n6345), .A2(n7745), .ZN(n9415) );
  NAND2_X1 U5599 ( .A1(n5490), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5514) );
  INV_X1 U5600 ( .A(n5491), .ZN(n5490) );
  OR2_X1 U5601 ( .A1(n5467), .A2(n9001), .ZN(n5491) );
  NAND2_X1 U5602 ( .A1(n4728), .A2(n4733), .ZN(n9431) );
  NAND2_X1 U5603 ( .A1(n9457), .A2(n4735), .ZN(n4728) );
  OAI21_X1 U5604 ( .B1(n9442), .B2(n6307), .A(n6306), .ZN(n9429) );
  OR2_X1 U5605 ( .A1(n9587), .A2(n9132), .ZN(n6306) );
  OAI21_X1 U5606 ( .B1(n4718), .B2(n4512), .A(n4510), .ZN(n9497) );
  INV_X1 U5607 ( .A(n7726), .ZN(n4512) );
  NAND2_X1 U5608 ( .A1(n6343), .A2(n4511), .ZN(n4510) );
  AND2_X1 U5609 ( .A1(n4371), .A2(n7726), .ZN(n4511) );
  AND2_X1 U5610 ( .A1(n5332), .A2(n5331), .ZN(n7229) );
  NAND2_X1 U5611 ( .A1(n4482), .A2(n4481), .ZN(n7220) );
  AOI21_X1 U5612 ( .B1(n4484), .B2(n4486), .A(n4423), .ZN(n4481) );
  NAND2_X1 U5613 ( .A1(n7042), .A2(n4484), .ZN(n4482) );
  INV_X1 U5614 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5237) );
  OR2_X1 U5615 ( .A1(n7327), .A2(n7816), .ZN(n7330) );
  NAND2_X1 U5616 ( .A1(n4483), .A2(n4881), .ZN(n7326) );
  NAND2_X1 U5617 ( .A1(n7042), .A2(n4879), .ZN(n4483) );
  NAND2_X1 U5618 ( .A1(n4493), .A2(n7888), .ZN(n7115) );
  AND2_X1 U5619 ( .A1(n7886), .A2(n7814), .ZN(n4493) );
  OR2_X1 U5620 ( .A1(n5208), .A2(n7305), .ZN(n5210) );
  INV_X1 U5621 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5192) );
  OR2_X1 U5622 ( .A1(n5210), .A2(n5192), .ZN(n5257) );
  INV_X1 U5623 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5148) );
  OR2_X1 U5624 ( .A1(n5149), .A2(n5148), .ZN(n5208) );
  NAND2_X1 U5625 ( .A1(n6290), .A2(n9063), .ZN(n6651) );
  OR2_X1 U5626 ( .A1(n6599), .A2(n9063), .ZN(n6647) );
  NAND2_X1 U5627 ( .A1(n6651), .A2(n7881), .ZN(n7804) );
  NAND2_X1 U5628 ( .A1(n6567), .A2(n6587), .ZN(n6599) );
  NOR2_X1 U5629 ( .A1(n6545), .A2(n6551), .ZN(n6567) );
  NAND2_X1 U5630 ( .A1(n6287), .A2(n6543), .ZN(n6532) );
  NAND2_X1 U5631 ( .A1(n6328), .A2(n6546), .ZN(n6545) );
  INV_X1 U5632 ( .A(n9531), .ZN(n9510) );
  NAND2_X1 U5633 ( .A1(n7784), .A2(n7783), .ZN(n7945) );
  AND2_X1 U5634 ( .A1(n9125), .A2(n7946), .ZN(n9530) );
  NAND2_X1 U5635 ( .A1(n5642), .A2(n5641), .ZN(n9549) );
  NAND2_X1 U5636 ( .A1(n5371), .A2(n5370), .ZN(n9606) );
  NOR2_X1 U5637 ( .A1(n7044), .A2(n7384), .ZN(n7124) );
  INV_X1 U5638 ( .A(n9869), .ZN(n9625) );
  NAND2_X1 U5639 ( .A1(n7332), .A2(n9627), .ZN(n9869) );
  XNOR2_X1 U5640 ( .A(n7780), .B(n7779), .ZN(n8216) );
  XNOR2_X1 U5641 ( .A(n4941), .B(P1_IR_REG_29__SCAN_IN), .ZN(n4946) );
  NAND2_X1 U5642 ( .A1(n9679), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4988) );
  AND2_X1 U5643 ( .A1(n6105), .A2(n5668), .ZN(n6103) );
  OAI21_X1 U5644 ( .B1(n4984), .B2(n4961), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4781) );
  NAND2_X1 U5645 ( .A1(n4960), .A2(n4959), .ZN(n4961) );
  XNOR2_X1 U5646 ( .A(n4969), .B(n4968), .ZN(n5712) );
  INV_X1 U5647 ( .A(SI_20_), .ZN(n10170) );
  NAND2_X1 U5648 ( .A1(n4907), .A2(n4816), .ZN(n4815) );
  INV_X1 U5649 ( .A(n5313), .ZN(n4816) );
  NAND2_X1 U5650 ( .A1(n4453), .A2(n5280), .ZN(n5284) );
  NAND2_X1 U5651 ( .A1(n4809), .A2(n4810), .ZN(n5248) );
  OR2_X1 U5652 ( .A1(n5180), .A2(n4813), .ZN(n4809) );
  NAND2_X1 U5653 ( .A1(n4725), .A2(n4723), .ZN(n5180) );
  NAND2_X1 U5654 ( .A1(n5172), .A2(n4804), .ZN(n4462) );
  NAND2_X1 U5655 ( .A1(n5157), .A2(n4803), .ZN(n4725) );
  CLKBUF_X1 U5656 ( .A(n5161), .Z(n5162) );
  NOR2_X2 U5657 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4990) );
  NOR2_X2 U5658 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4991) );
  XNOR2_X1 U5659 ( .A(n5000), .B(n4999), .ZN(n5023) );
  NAND2_X1 U5660 ( .A1(n7456), .A2(n4863), .ZN(n7459) );
  NAND2_X1 U5661 ( .A1(n4845), .A2(n8190), .ZN(n8039) );
  OAI211_X1 U5662 ( .C1(n5832), .C2(n6691), .A(n5849), .B(n5848), .ZN(n7068)
         );
  OR2_X1 U5663 ( .A1(n5827), .A2(n6395), .ZN(n5848) );
  NAND2_X1 U5664 ( .A1(n4842), .A2(n4840), .ZN(n4839) );
  OR2_X1 U5665 ( .A1(n4846), .A2(n8030), .ZN(n4842) );
  NAND2_X1 U5666 ( .A1(n4846), .A2(n4841), .ZN(n4840) );
  NAND2_X1 U5667 ( .A1(n4850), .A2(n4844), .ZN(n4841) );
  OR2_X1 U5668 ( .A1(n4844), .A2(n4850), .ZN(n4843) );
  OR2_X1 U5669 ( .A1(n6412), .A2(n5827), .ZN(n5907) );
  AOI21_X1 U5670 ( .B1(n4854), .B2(n4856), .A(n7612), .ZN(n4853) );
  OR2_X1 U5671 ( .A1(n6399), .A2(n5827), .ZN(n5872) );
  NAND2_X1 U5672 ( .A1(n7545), .A2(n7544), .ZN(n7595) );
  AND2_X1 U5673 ( .A1(n8075), .A2(n8125), .ZN(n8128) );
  INV_X1 U5674 ( .A(n8465), .ZN(n7211) );
  INV_X1 U5675 ( .A(n8205), .ZN(n8120) );
  INV_X1 U5676 ( .A(n8199), .ZN(n8179) );
  OR2_X1 U5677 ( .A1(n6402), .A2(n5827), .ZN(n5884) );
  NAND2_X1 U5678 ( .A1(n6920), .A2(n9697), .ZN(n8196) );
  NAND2_X1 U5679 ( .A1(n6080), .A2(n6079), .ZN(n8671) );
  INV_X1 U5680 ( .A(n8799), .ZN(n8208) );
  NAND2_X1 U5681 ( .A1(n6942), .A2(n6941), .ZN(n8210) );
  NOR2_X1 U5682 ( .A1(n8200), .A2(n4865), .ZN(n4864) );
  INV_X1 U5683 ( .A(n7983), .ZN(n4865) );
  NAND2_X1 U5684 ( .A1(n8046), .A2(n7983), .ZN(n8201) );
  INV_X1 U5685 ( .A(n7607), .ZN(n8457) );
  NAND4_X1 U5686 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n8464)
         );
  NAND2_X1 U5687 ( .A1(n5822), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5805) );
  NAND4_X1 U5688 ( .A1(n5816), .A2(n5815), .A3(n5814), .A4(n5813), .ZN(n8466)
         );
  OR2_X1 U5689 ( .A1(n6124), .A2(n10044), .ZN(n5815) );
  NAND2_X1 U5690 ( .A1(n5839), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5816) );
  OR2_X2 U5691 ( .A1(n6671), .A2(P2_U3151), .ZN(n8609) );
  AND2_X1 U5692 ( .A1(n6673), .A2(n6672), .ZN(n9886) );
  INV_X1 U5693 ( .A(n4759), .ZN(n6986) );
  INV_X1 U5694 ( .A(n4758), .ZN(n6990) );
  INV_X1 U5695 ( .A(n4751), .ZN(n7181) );
  INV_X1 U5696 ( .A(n4741), .ZN(n7431) );
  NOR2_X1 U5697 ( .A1(n8470), .A2(n8471), .ZN(n8496) );
  NOR2_X1 U5698 ( .A1(n8527), .A2(n8528), .ZN(n8549) );
  NAND2_X1 U5699 ( .A1(n4744), .A2(n4742), .ZN(n8577) );
  NAND2_X1 U5700 ( .A1(n8550), .A2(n4745), .ZN(n4744) );
  OR2_X1 U5701 ( .A1(n8527), .A2(n4743), .ZN(n4742) );
  NAND2_X1 U5702 ( .A1(n4745), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U5703 ( .A1(n4753), .A2(n4752), .ZN(n8622) );
  NAND2_X1 U5704 ( .A1(n4552), .A2(n4551), .ZN(n4550) );
  INV_X1 U5705 ( .A(n8619), .ZN(n4552) );
  AOI21_X1 U5706 ( .B1(n8954), .B2(n8224), .A(n8223), .ZN(n8833) );
  NAND2_X1 U5707 ( .A1(n4662), .A2(n4667), .ZN(n8215) );
  NAND2_X1 U5708 ( .A1(n4666), .A2(n4660), .ZN(n4662) );
  OR2_X1 U5709 ( .A1(n6275), .A2(n8795), .ZN(n6272) );
  AND2_X1 U5710 ( .A1(n4666), .A2(n8407), .ZN(n6223) );
  NAND2_X1 U5711 ( .A1(n6091), .A2(n6090), .ZN(n8661) );
  NAND2_X1 U5712 ( .A1(n4580), .A2(n4583), .ZN(n8666) );
  AND2_X1 U5713 ( .A1(n4649), .A2(n4646), .ZN(n8698) );
  NAND2_X1 U5714 ( .A1(n6006), .A2(n6005), .ZN(n8878) );
  OAI21_X1 U5715 ( .B1(n7559), .B2(n4640), .A(n4637), .ZN(n8829) );
  NAND2_X1 U5716 ( .A1(n9932), .A2(n6186), .ZN(n9699) );
  NAND2_X1 U5717 ( .A1(n7558), .A2(n8331), .ZN(n7570) );
  AND2_X1 U5718 ( .A1(n7268), .A2(n5898), .ZN(n7391) );
  OR2_X1 U5719 ( .A1(n5827), .A2(n6392), .ZN(n5859) );
  INV_X1 U5720 ( .A(n8795), .ZN(n8830) );
  OR2_X1 U5721 ( .A1(n6268), .A2(n9699), .ZN(n8807) );
  OR2_X1 U5722 ( .A1(n6939), .A2(n6264), .ZN(n9697) );
  INV_X1 U5723 ( .A(n8807), .ZN(n8792) );
  NAND2_X2 U5724 ( .A1(n6268), .A2(n9697), .ZN(n9716) );
  OR2_X1 U5725 ( .A1(n6275), .A2(n8881), .ZN(n6280) );
  INV_X1 U5726 ( .A(n8671), .ZN(n8892) );
  NAND2_X1 U5727 ( .A1(n6070), .A2(n6069), .ZN(n8895) );
  NAND2_X1 U5728 ( .A1(n4588), .A2(n4586), .ZN(n8678) );
  NAND2_X1 U5729 ( .A1(n6063), .A2(n6062), .ZN(n8902) );
  OAI21_X1 U5730 ( .B1(n8741), .B2(n4570), .A(n4568), .ZN(n8705) );
  NAND2_X1 U5731 ( .A1(n4649), .A2(n4650), .ZN(n8703) );
  NAND2_X1 U5732 ( .A1(n4567), .A2(n4571), .ZN(n8719) );
  AOI21_X1 U5733 ( .B1(n8727), .B2(n8384), .A(n4655), .ZN(n8715) );
  NAND2_X1 U5734 ( .A1(n6045), .A2(n6044), .ZN(n8920) );
  NAND2_X1 U5735 ( .A1(n6039), .A2(n6038), .ZN(n8926) );
  NAND2_X1 U5736 ( .A1(n6016), .A2(n6015), .ZN(n8945) );
  AND2_X1 U5737 ( .A1(n9722), .A2(n9721), .ZN(n9732) );
  INV_X1 U5738 ( .A(n7543), .ZN(n7581) );
  INV_X1 U5739 ( .A(n6259), .ZN(n6491) );
  INV_X1 U5740 ( .A(n6939), .ZN(n6517) );
  AND2_X1 U5741 ( .A1(n6932), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6580) );
  AND2_X1 U5742 ( .A1(n6389), .A2(P2_U3151), .ZN(n8958) );
  INV_X1 U5743 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5783) );
  INV_X1 U5744 ( .A(n6146), .ZN(n7631) );
  INV_X1 U5745 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U5746 ( .A1(n4831), .A2(n4835), .ZN(n6140) );
  AOI22_X1 U5747 ( .A1(n4835), .A2(n4837), .B1(n4834), .B2(
        P2_IR_REG_23__SCAN_IN), .ZN(n4832) );
  OR2_X1 U5748 ( .A1(n6166), .A2(n4833), .ZN(n4830) );
  INV_X1 U5749 ( .A(n8448), .ZN(n7552) );
  INV_X1 U5750 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7490) );
  XNOR2_X1 U5751 ( .A(n6119), .B(n4869), .ZN(n8269) );
  NAND2_X1 U5752 ( .A1(n6122), .A2(n6121), .ZN(n8423) );
  INV_X1 U5753 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7315) );
  INV_X1 U5754 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7218) );
  INV_X1 U5755 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7131) );
  INV_X1 U5756 ( .A(n8495), .ZN(n8509) );
  INV_X1 U5757 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6423) );
  INV_X1 U5758 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6413) );
  INV_X1 U5759 ( .A(n7003), .ZN(n7102) );
  INV_X1 U5760 ( .A(n6807), .ZN(n6812) );
  XNOR2_X1 U5761 ( .A(n4761), .B(n5807), .ZN(n6732) );
  NAND2_X1 U5762 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4761) );
  NAND2_X1 U5763 ( .A1(n4784), .A2(n4783), .ZN(n8984) );
  AND2_X1 U5764 ( .A1(n5242), .A2(n5241), .ZN(n7411) );
  AND2_X1 U5765 ( .A1(n9104), .A2(n5690), .ZN(n6203) );
  INV_X1 U5766 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7305) );
  XNOR2_X1 U5767 ( .A(n5054), .B(n5056), .ZN(n7961) );
  AND2_X1 U5768 ( .A1(n5595), .A2(n5594), .ZN(n9382) );
  AND2_X1 U5769 ( .A1(n5618), .A2(n5645), .ZN(n9356) );
  AND2_X1 U5770 ( .A1(n5129), .A2(n5128), .ZN(n6953) );
  INV_X1 U5771 ( .A(n4777), .ZN(n4776) );
  AND2_X1 U5772 ( .A1(n5725), .A2(n5713), .ZN(n9060) );
  AND2_X1 U5773 ( .A1(n7404), .A2(n5312), .ZN(n7480) );
  NAND2_X1 U5774 ( .A1(n8987), .A2(n5553), .ZN(n9078) );
  INV_X1 U5775 ( .A(n9124), .ZN(n9096) );
  AND2_X1 U5776 ( .A1(n5725), .A2(n5714), .ZN(n9115) );
  NAND2_X1 U5777 ( .A1(n5724), .A2(n7931), .ZN(n9121) );
  NOR2_X1 U5778 ( .A1(n7932), .A2(n7931), .ZN(n7933) );
  NAND2_X1 U5779 ( .A1(n4459), .A2(n7928), .ZN(n7934) );
  NOR2_X1 U5780 ( .A1(n7930), .A2(n7929), .ZN(n7932) );
  INV_X1 U5781 ( .A(n9350), .ZN(n9128) );
  INV_X1 U5782 ( .A(n7328), .ZN(n9134) );
  INV_X1 U5783 ( .A(n7411), .ZN(n9135) );
  INV_X1 U5784 ( .A(n6952), .ZN(n9137) );
  INV_X1 U5785 ( .A(n6740), .ZN(n9138) );
  INV_X1 U5786 ( .A(n6953), .ZN(n9139) );
  INV_X1 U5787 ( .A(n6739), .ZN(n9140) );
  NAND2_X1 U5788 ( .A1(n4953), .A2(n4952), .ZN(n9141) );
  NAND2_X1 U5789 ( .A1(n5073), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U5790 ( .A1(n5349), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5040) );
  OR2_X1 U5791 ( .A1(n5057), .A2(n5036), .ZN(n5038) );
  NAND2_X1 U5792 ( .A1(n4873), .A2(n6319), .ZN(n9291) );
  NAND2_X1 U5793 ( .A1(n9349), .A2(n7760), .ZN(n9337) );
  NAND2_X1 U5794 ( .A1(n4710), .A2(n4714), .ZN(n9336) );
  NAND2_X1 U5795 ( .A1(n4878), .A2(n4614), .ZN(n9559) );
  INV_X1 U5796 ( .A(n9367), .ZN(n4878) );
  NAND2_X1 U5797 ( .A1(n9417), .A2(n7749), .ZN(n9405) );
  NAND2_X1 U5798 ( .A1(n4737), .A2(n7742), .ZN(n9444) );
  OR2_X1 U5799 ( .A1(n9457), .A2(n7801), .ZN(n4737) );
  NAND2_X1 U5800 ( .A1(n5464), .A2(n5463), .ZN(n9592) );
  NAND2_X1 U5801 ( .A1(n4894), .A2(n4901), .ZN(n9455) );
  NAND2_X1 U5802 ( .A1(n6304), .A2(n4899), .ZN(n4894) );
  NAND2_X1 U5803 ( .A1(n6304), .A2(n6303), .ZN(n9470) );
  OR2_X1 U5804 ( .A1(n7364), .A2(n4477), .ZN(n4470) );
  NAND2_X1 U5805 ( .A1(n7473), .A2(n7722), .ZN(n9519) );
  NAND2_X1 U5806 ( .A1(n7364), .A2(n4883), .ZN(n4478) );
  NAND2_X1 U5807 ( .A1(n7362), .A2(n6300), .ZN(n7470) );
  NAND2_X1 U5808 ( .A1(n7121), .A2(n7120), .ZN(n7119) );
  NAND2_X1 U5809 ( .A1(n7040), .A2(n6298), .ZN(n7121) );
  OR2_X1 U5810 ( .A1(n6356), .A2(n7936), .ZN(n9390) );
  OR2_X1 U5811 ( .A1(n9826), .A2(n6615), .ZN(n9529) );
  OR2_X1 U5812 ( .A1(n9826), .A2(n9269), .ZN(n9841) );
  INV_X1 U5813 ( .A(n9514), .ZN(n9838) );
  AND2_X1 U5814 ( .A1(n9876), .A2(n9623), .ZN(n6606) );
  INV_X1 U5815 ( .A(n7945), .ZN(n7956) );
  INV_X1 U5816 ( .A(n9322), .ZN(n9643) );
  INV_X1 U5817 ( .A(n9422), .ZN(n9657) );
  NAND2_X2 U5818 ( .A1(n6418), .A2(n6417), .ZN(n9847) );
  NAND2_X1 U5819 ( .A1(n4685), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4871) );
  AND2_X1 U5820 ( .A1(n4624), .A2(n4409), .ZN(n4623) );
  XNOR2_X1 U5821 ( .A(n6229), .B(n6228), .ZN(n8965) );
  XNOR2_X1 U5822 ( .A(n6104), .B(n6103), .ZN(n9690) );
  XNOR2_X1 U5823 ( .A(n4965), .B(n4964), .ZN(n7628) );
  NAND2_X1 U5824 ( .A1(n4466), .A2(n5554), .ZN(n5582) );
  OR2_X1 U5825 ( .A1(n5556), .A2(n5555), .ZN(n4466) );
  INV_X1 U5826 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7555) );
  OR2_X1 U5827 ( .A1(n4985), .A2(n4959), .ZN(n4986) );
  INV_X1 U5828 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7500) );
  CLKBUF_X1 U5829 ( .A(n5712), .Z(n7798) );
  INV_X1 U5830 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U5831 ( .A1(n4802), .A2(n5159), .ZN(n5173) );
  NAND2_X1 U5832 ( .A1(n5157), .A2(n5156), .ZN(n4802) );
  XNOR2_X1 U5833 ( .A(n4535), .B(n8638), .ZN(n8451) );
  XNOR2_X1 U5834 ( .A(n4546), .B(n8634), .ZN(n4545) );
  INV_X1 U5835 ( .A(n6255), .ZN(n6256) );
  OAI22_X1 U5836 ( .A1(n8654), .A2(n8855), .B1(n9950), .B2(n6254), .ZN(n6255)
         );
  OR2_X1 U5837 ( .A1(n6274), .A2(n9939), .ZN(n6190) );
  NAND2_X1 U5838 ( .A1(n6226), .A2(n6225), .ZN(P2_U3454) );
  MUX2_X1 U5839 ( .A(n9533), .B(n9635), .S(n9876), .Z(n9534) );
  MUX2_X1 U5840 ( .A(n9636), .B(n9635), .S(n9871), .Z(n9637) );
  NAND2_X1 U5841 ( .A1(n4488), .A2(n6371), .ZN(P1_U3519) );
  OAI21_X1 U5842 ( .B1(n4739), .B2(n4489), .A(n6370), .ZN(n4488) );
  AND2_X1 U5843 ( .A1(n4810), .A2(n4373), .ZN(n4355) );
  INV_X1 U5844 ( .A(n8381), .ZN(n4529) );
  AND2_X1 U5845 ( .A1(n7855), .A2(n7858), .ZN(n7778) );
  AND2_X1 U5846 ( .A1(n9070), .A2(n5503), .ZN(n4356) );
  OR2_X1 U5847 ( .A1(n9592), .A2(n9474), .ZN(n4357) );
  OR2_X1 U5848 ( .A1(n8605), .A2(n8599), .ZN(n4358) );
  AND2_X1 U5849 ( .A1(n5834), .A2(n4403), .ZN(n4359) );
  AOI21_X1 U5850 ( .B1(n5822), .B2(n8031), .A(n6114), .ZN(n8042) );
  INV_X1 U5851 ( .A(n8042), .ZN(n4670) );
  INV_X1 U5852 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4930) );
  AND2_X1 U5853 ( .A1(n8671), .A2(n8681), .ZN(n4360) );
  AND2_X1 U5854 ( .A1(n9286), .A2(n6353), .ZN(n4361) );
  INV_X1 U5855 ( .A(n8716), .ZN(n4654) );
  AND2_X1 U5856 ( .A1(n9571), .A2(n9130), .ZN(n4362) );
  AND2_X1 U5857 ( .A1(n4706), .A2(n9452), .ZN(n4363) );
  AND2_X1 U5858 ( .A1(n4361), .A2(n9876), .ZN(n4364) );
  AND2_X1 U5859 ( .A1(n7834), .A2(n7839), .ZN(n9368) );
  INV_X1 U5860 ( .A(n9368), .ZN(n4614) );
  INV_X1 U5861 ( .A(n4908), .ZN(n4813) );
  INV_X1 U5862 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U5863 ( .A1(n4931), .A2(n4893), .ZN(n4365) );
  INV_X1 U5864 ( .A(n9414), .ZN(n4509) );
  OR2_X1 U5865 ( .A1(n7044), .A2(n4690), .ZN(n4366) );
  AND4_X1 U5866 ( .A1(n5797), .A2(n5796), .A3(n5795), .A4(n5794), .ZN(n8182)
         );
  INV_X1 U5867 ( .A(n8182), .ZN(n8769) );
  NAND2_X1 U5868 ( .A1(n5869), .A2(n4866), .ZN(n5893) );
  OR2_X1 U5869 ( .A1(n8920), .A2(n8130), .ZN(n8386) );
  NAND2_X1 U5870 ( .A1(n5665), .A2(n5664), .ZN(n6104) );
  INV_X1 U5871 ( .A(n8239), .ZN(n4661) );
  INV_X1 U5872 ( .A(n5838), .ZN(n6127) );
  NAND2_X1 U5873 ( .A1(n9331), .A2(n4696), .ZN(n4367) );
  OR2_X1 U5874 ( .A1(n8825), .A2(n9709), .ZN(n8357) );
  NOR2_X1 U5875 ( .A1(n5761), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5782) );
  AND2_X1 U5876 ( .A1(n4509), .A2(n7745), .ZN(n4368) );
  NAND2_X1 U5877 ( .A1(n5811), .A2(n5820), .ZN(n6175) );
  INV_X1 U5878 ( .A(n7120), .ZN(n7814) );
  XNOR2_X1 U5879 ( .A(n4871), .B(n9682), .ZN(n4948) );
  AND3_X1 U5880 ( .A1(n5843), .A2(n5842), .A3(n5841), .ZN(n4369) );
  AND2_X1 U5881 ( .A1(n4860), .A2(n8008), .ZN(n4370) );
  XNOR2_X1 U5882 ( .A(n5784), .B(n5783), .ZN(n5787) );
  INV_X1 U5883 ( .A(n8392), .ZN(n4648) );
  INV_X1 U5884 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U5885 ( .A1(n9559), .A2(n6313), .ZN(n9345) );
  AND2_X1 U5886 ( .A1(n7821), .A2(n7721), .ZN(n4371) );
  NAND3_X1 U5887 ( .A1(n4830), .A2(n4829), .A3(n4832), .ZN(n6145) );
  AND2_X1 U5888 ( .A1(n4870), .A2(n6116), .ZN(n4372) );
  INV_X1 U5889 ( .A(n4477), .ZN(n4476) );
  NAND2_X1 U5890 ( .A1(n4884), .A2(n4375), .ZN(n4477) );
  NAND2_X1 U5891 ( .A1(n4487), .A2(n6317), .ZN(n9310) );
  XOR2_X1 U5892 ( .A(n5227), .B(SI_10_), .Z(n4373) );
  NAND2_X1 U5893 ( .A1(n6192), .A2(n6191), .ZN(n9536) );
  INV_X1 U5894 ( .A(n9536), .ZN(n4699) );
  AND2_X1 U5895 ( .A1(n9592), .A2(n9474), .ZN(n4374) );
  INV_X1 U5896 ( .A(n8252), .ZN(n4593) );
  XNOR2_X1 U5897 ( .A(n8267), .B(n8042), .ZN(n8239) );
  INV_X1 U5898 ( .A(n6985), .ZN(n7000) );
  INV_X1 U5899 ( .A(n5820), .ZN(n6973) );
  NAND4_X1 U5900 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n6843)
         );
  INV_X1 U5901 ( .A(n6843), .ZN(n4562) );
  OR2_X1 U5902 ( .A1(n9606), .A2(n9499), .ZN(n4375) );
  NAND2_X1 U5903 ( .A1(n9037), .A2(n9038), .ZN(n9036) );
  NAND2_X1 U5904 ( .A1(n4976), .A2(n5718), .ZN(n5014) );
  NAND2_X1 U5905 ( .A1(n7721), .A2(n7894), .ZN(n7363) );
  NAND2_X1 U5906 ( .A1(n8214), .A2(n8220), .ZN(n8418) );
  INV_X1 U5907 ( .A(n8418), .ZN(n4806) );
  INV_X1 U5908 ( .A(n5179), .ZN(n4812) );
  AND2_X1 U5909 ( .A1(n4560), .A2(n4661), .ZN(n4376) );
  OR2_X1 U5910 ( .A1(n4610), .A2(n4609), .ZN(n4377) );
  NAND2_X1 U5911 ( .A1(n5829), .A2(n5830), .ZN(n5845) );
  NAND2_X1 U5912 ( .A1(n5869), .A2(n5744), .ZN(n5880) );
  INV_X1 U5913 ( .A(n4653), .ZN(n4652) );
  OAI21_X1 U5914 ( .B1(n4655), .B2(n8384), .A(n4654), .ZN(n4653) );
  NAND2_X1 U5915 ( .A1(n5540), .A2(n5539), .ZN(n9571) );
  NOR2_X1 U5916 ( .A1(n8550), .A2(n8549), .ZN(n4378) );
  NAND2_X1 U5917 ( .A1(n5869), .A2(n4867), .ZN(n4379) );
  NAND2_X1 U5918 ( .A1(n5589), .A2(n5588), .ZN(n9560) );
  OR2_X1 U5919 ( .A1(n6985), .A2(n6984), .ZN(n4380) );
  NAND2_X1 U5920 ( .A1(n9036), .A2(n5438), .ZN(n8994) );
  INV_X1 U5921 ( .A(n9301), .ZN(n4505) );
  AND2_X1 U5922 ( .A1(n7854), .A2(n7852), .ZN(n9301) );
  AND2_X1 U5923 ( .A1(n5027), .A2(n4687), .ZN(n4381) );
  AND2_X1 U5924 ( .A1(n4608), .A2(n7706), .ZN(n4382) );
  INV_X1 U5925 ( .A(n9481), .ZN(n9664) );
  NAND2_X1 U5926 ( .A1(n5424), .A2(n5423), .ZN(n9481) );
  INV_X1 U5927 ( .A(n4461), .ZN(n4803) );
  OAI21_X1 U5928 ( .B1(n4804), .B2(n5156), .A(n5172), .ZN(n4461) );
  AND2_X1 U5929 ( .A1(n4502), .A2(n4505), .ZN(n4383) );
  AND2_X1 U5930 ( .A1(n4588), .A2(n4585), .ZN(n4384) );
  AND2_X1 U5931 ( .A1(n8267), .A2(n4670), .ZN(n4385) );
  AND2_X1 U5932 ( .A1(n6318), .A2(n6317), .ZN(n4386) );
  NAND2_X1 U5933 ( .A1(n6322), .A2(n6321), .ZN(n9284) );
  INV_X1 U5934 ( .A(n5438), .ZN(n4768) );
  INV_X1 U5935 ( .A(n4668), .ZN(n4667) );
  OAI21_X1 U5936 ( .B1(n8239), .B2(n4672), .A(n4669), .ZN(n4668) );
  OR2_X1 U5937 ( .A1(n6682), .A2(n9942), .ZN(n4387) );
  AND4_X1 U5938 ( .A1(n9301), .A2(n9313), .A3(n9338), .A4(n7829), .ZN(n4388)
         );
  NOR2_X1 U5939 ( .A1(n7127), .A2(n9136), .ZN(n4389) );
  INV_X1 U5940 ( .A(n5201), .ZN(n4724) );
  INV_X1 U5941 ( .A(n8986), .ZN(n4787) );
  NAND2_X1 U5942 ( .A1(n5338), .A2(n5337), .ZN(n4390) );
  INV_X1 U5943 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6167) );
  INV_X1 U5944 ( .A(n4464), .ZN(n7921) );
  OR2_X1 U5945 ( .A1(n9638), .A2(n9125), .ZN(n4464) );
  NOR2_X1 U5946 ( .A1(n8914), .A2(n8734), .ZN(n4391) );
  INV_X1 U5947 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4964) );
  NOR2_X1 U5948 ( .A1(n8908), .A2(n8694), .ZN(n4392) );
  NAND2_X1 U5949 ( .A1(n5504), .A2(n9069), .ZN(n4393) );
  OR2_X1 U5950 ( .A1(n4679), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U5951 ( .A1(n5798), .A2(n4870), .ZN(n4395) );
  NAND2_X1 U5952 ( .A1(n5798), .A2(n5799), .ZN(n4396) );
  NAND2_X1 U5953 ( .A1(n8149), .A2(n8147), .ZN(n4397) );
  AND2_X1 U5954 ( .A1(n5227), .A2(SI_10_), .ZN(n4398) );
  INV_X1 U5955 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U5956 ( .A1(n4370), .A2(n8079), .ZN(n4399) );
  AND2_X1 U5957 ( .A1(n8677), .A2(n8693), .ZN(n4400) );
  INV_X1 U5958 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4939) );
  OR2_X1 U5959 ( .A1(n5761), .A2(n4684), .ZN(n4401) );
  OAI21_X1 U5960 ( .B1(n7611), .B2(n8160), .A(n7610), .ZN(n7612) );
  NAND2_X1 U5961 ( .A1(n4479), .A2(n6312), .ZN(n9367) );
  AND2_X1 U5962 ( .A1(n5143), .A2(n5142), .ZN(n4402) );
  INV_X1 U5963 ( .A(n6328), .ZN(n9837) );
  OR2_X1 U5964 ( .A1(n5832), .A2(n4354), .ZN(n4403) );
  INV_X1 U5965 ( .A(n4722), .ZN(n4723) );
  NAND2_X1 U5966 ( .A1(n4801), .A2(n4724), .ZN(n4722) );
  NAND2_X1 U5967 ( .A1(n5483), .A2(n4767), .ZN(n4404) );
  INV_X1 U5968 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5759) );
  AND2_X1 U5969 ( .A1(n6205), .A2(n9115), .ZN(n4405) );
  OR2_X1 U5970 ( .A1(n8902), .A2(n8707), .ZN(n8398) );
  AND2_X1 U5971 ( .A1(n4637), .A2(n8357), .ZN(n4406) );
  INV_X1 U5972 ( .A(n8313), .ZN(n4631) );
  INV_X1 U5973 ( .A(n4586), .ZN(n4584) );
  NOR2_X1 U5974 ( .A1(n8686), .A2(n4587), .ZN(n4586) );
  AND2_X1 U5975 ( .A1(n5198), .A2(n5197), .ZN(n7306) );
  INV_X1 U5976 ( .A(n7306), .ZN(n4726) );
  NAND2_X1 U5977 ( .A1(n6388), .A2(n5808), .ZN(n4407) );
  NOR2_X1 U5978 ( .A1(n7871), .A2(n5718), .ZN(n4408) );
  NOR2_X1 U5979 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4409) );
  INV_X1 U5980 ( .A(n6313), .ZN(n4877) );
  AND2_X1 U5981 ( .A1(n4505), .A2(n6319), .ZN(n4410) );
  AND2_X1 U5982 ( .A1(n4846), .A2(n4844), .ZN(n4411) );
  AND2_X1 U5983 ( .A1(n4756), .A2(n4358), .ZN(n4412) );
  NAND3_X1 U5984 ( .A1(n6202), .A2(n9115), .A3(n6201), .ZN(n4413) );
  AND2_X1 U5985 ( .A1(n4787), .A2(n4786), .ZN(n4414) );
  NAND2_X1 U5986 ( .A1(n5174), .A2(SI_7_), .ZN(n4415) );
  INV_X1 U5987 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4958) );
  INV_X1 U5988 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4968) );
  OR2_X1 U5989 ( .A1(n7698), .A2(n4598), .ZN(n4416) );
  INV_X1 U5990 ( .A(n5167), .ZN(n6197) );
  AND2_X1 U5991 ( .A1(n5792), .A2(n5791), .ZN(n5822) );
  INV_X2 U5992 ( .A(n7207), .ZN(n8029) );
  XNOR2_X1 U5993 ( .A(n4781), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5693) );
  AND2_X1 U5994 ( .A1(n9398), .A2(n4704), .ZN(n4417) );
  NAND2_X1 U5995 ( .A1(n6107), .A2(n6106), .ZN(n8267) );
  INV_X1 U5996 ( .A(n8267), .ZN(n4671) );
  AND2_X1 U5997 ( .A1(n9422), .A2(n9407), .ZN(n4418) );
  AND2_X1 U5998 ( .A1(n5363), .A2(n10168), .ZN(n4419) );
  INV_X1 U5999 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4497) );
  AND2_X1 U6000 ( .A1(n7866), .A2(n5718), .ZN(n5713) );
  OAI21_X1 U6001 ( .B1(n9429), .B2(n6308), .A(n6309), .ZN(n9413) );
  INV_X1 U6002 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4959) );
  NAND2_X1 U6003 ( .A1(n4578), .A2(n6037), .ZN(n8752) );
  NAND2_X1 U6004 ( .A1(n4636), .A2(n4632), .ZN(n9696) );
  NAND2_X1 U6005 ( .A1(n4470), .A2(n4474), .ZN(n9488) );
  NAND2_X1 U6006 ( .A1(n4478), .A2(n4884), .ZN(n9507) );
  NAND2_X1 U6007 ( .A1(n5450), .A2(n5449), .ZN(n9587) );
  INV_X1 U6008 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4869) );
  NAND2_X1 U6009 ( .A1(n9025), .A2(n9027), .ZN(n9023) );
  AND2_X1 U6010 ( .A1(n7390), .A2(n5908), .ZN(n7491) );
  AND3_X1 U6011 ( .A1(n4351), .A2(n4866), .A3(n5869), .ZN(n6000) );
  NOR2_X1 U6012 ( .A1(n5384), .A2(n5383), .ZN(n9112) );
  NOR2_X1 U6013 ( .A1(n9434), .A2(n9422), .ZN(n9398) );
  AND2_X1 U6014 ( .A1(n4718), .A2(n7473), .ZN(n4420) );
  NOR2_X1 U6015 ( .A1(n8497), .A2(n8496), .ZN(n4421) );
  AND2_X1 U6016 ( .A1(n9606), .A2(n9499), .ZN(n4422) );
  NAND2_X1 U6017 ( .A1(n9490), .A2(n4363), .ZN(n4707) );
  NAND2_X1 U6018 ( .A1(n5802), .A2(n5801), .ZN(n8932) );
  NOR2_X1 U6019 ( .A1(n7510), .A2(n9135), .ZN(n4423) );
  OR2_X1 U6020 ( .A1(n8671), .A2(n8681), .ZN(n4424) );
  AND2_X1 U6021 ( .A1(n5361), .A2(n4788), .ZN(n4425) );
  AND2_X1 U6022 ( .A1(n5444), .A2(SI_18_), .ZN(n4426) );
  NAND2_X1 U6023 ( .A1(n5614), .A2(n5613), .ZN(n9355) );
  INV_X1 U6024 ( .A(n9355), .ZN(n4701) );
  OAI21_X1 U6025 ( .B1(n9413), .B2(n4418), .A(n6310), .ZN(n9397) );
  AND2_X1 U6026 ( .A1(n6343), .A2(n7721), .ZN(n4427) );
  INV_X1 U6027 ( .A(n7510), .ZN(n9677) );
  NAND2_X1 U6028 ( .A1(n5233), .A2(n5232), .ZN(n7510) );
  NAND2_X1 U6029 ( .A1(n5489), .A2(n5488), .ZN(n9582) );
  AND2_X1 U6030 ( .A1(n4823), .A2(n5458), .ZN(n4428) );
  INV_X1 U6031 ( .A(n5362), .ZN(n5361) );
  INV_X1 U6032 ( .A(n6136), .ZN(n6166) );
  NAND2_X1 U6033 ( .A1(n7277), .A2(n8248), .ZN(n7276) );
  NAND2_X1 U6034 ( .A1(n4629), .A2(n4627), .ZN(n7270) );
  OAI21_X1 U6035 ( .B1(n8270), .B2(n8244), .A(n6175), .ZN(n7134) );
  AND2_X1 U6036 ( .A1(n7320), .A2(n5885), .ZN(n7267) );
  NAND2_X1 U6037 ( .A1(n6178), .A2(n8317), .ZN(n7494) );
  NOR3_X1 U6038 ( .A1(n7044), .A2(n4689), .A3(n9622), .ZN(n4688) );
  INV_X1 U6039 ( .A(n4693), .ZN(n7335) );
  NOR2_X1 U6040 ( .A1(n7044), .A2(n4689), .ZN(n4693) );
  NAND2_X1 U6041 ( .A1(n9055), .A2(n4776), .ZN(n4429) );
  NAND2_X1 U6042 ( .A1(n4727), .A2(n5188), .ZN(n7384) );
  INV_X1 U6043 ( .A(n7384), .ZN(n4691) );
  INV_X1 U6044 ( .A(n9622), .ZN(n4692) );
  XNOR2_X1 U6045 ( .A(n7022), .B(n5819), .ZN(n7029) );
  INV_X1 U6046 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4960) );
  AND2_X1 U6047 ( .A1(n6348), .A2(n7796), .ZN(n9518) );
  INV_X1 U6048 ( .A(n9518), .ZN(n9503) );
  NAND2_X1 U6049 ( .A1(n6532), .A2(n7805), .ZN(n6531) );
  OR2_X1 U6050 ( .A1(n6808), .A2(n6809), .ZN(n4746) );
  OR2_X1 U6051 ( .A1(n9878), .A2(n6686), .ZN(n8635) );
  XNOR2_X1 U6052 ( .A(n5800), .B(n6115), .ZN(n8638) );
  INV_X1 U6053 ( .A(n8624), .ZN(n8630) );
  AND2_X1 U6054 ( .A1(n5757), .A2(n4680), .ZN(n8955) );
  AND2_X1 U6055 ( .A1(n6880), .A2(n6810), .ZN(n4430) );
  INV_X1 U6056 ( .A(n8601), .ZN(n4755) );
  OR2_X1 U6057 ( .A1(n8624), .A2(n8771), .ZN(n4431) );
  INV_X1 U6058 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4709) );
  XNOR2_X1 U6059 ( .A(n4434), .B(n8627), .ZN(n8643) );
  NAND3_X1 U6060 ( .A1(n4752), .A2(n4753), .A3(n4431), .ZN(n4434) );
  XNOR2_X1 U6061 ( .A(n8599), .B(n8605), .ZN(n8579) );
  NAND2_X1 U6062 ( .A1(n4748), .A2(n4435), .ZN(n8525) );
  NOR2_X1 U6063 ( .A1(n7244), .A2(n7247), .ZN(n7428) );
  NOR2_X1 U6064 ( .A1(n7091), .A2(n7496), .ZN(n7176) );
  NAND2_X1 U6065 ( .A1(n6681), .A2(n6765), .ZN(n6769) );
  NAND2_X1 U6066 ( .A1(n4436), .A2(n5023), .ZN(n4492) );
  XNOR2_X1 U6067 ( .A(n4436), .B(n5023), .ZN(n6397) );
  NAND2_X1 U6068 ( .A1(n5043), .A2(n4998), .ZN(n4436) );
  NAND2_X1 U6069 ( .A1(n9007), .A2(n9008), .ZN(n9006) );
  AOI21_X2 U6070 ( .B1(n4764), .B2(n4763), .A(n4762), .ZN(n9007) );
  NAND3_X1 U6071 ( .A1(n4439), .A2(n5110), .A3(n4437), .ZN(n4494) );
  NAND2_X1 U6072 ( .A1(n4438), .A2(n5009), .ZN(n4437) );
  INV_X1 U6073 ( .A(n5082), .ZN(n4438) );
  NOR2_X1 U6074 ( .A1(n4443), .A2(n4441), .ZN(n4440) );
  INV_X1 U6075 ( .A(n5004), .ZN(n4441) );
  NAND2_X1 U6076 ( .A1(n4442), .A2(n5009), .ZN(n5111) );
  NAND2_X1 U6077 ( .A1(n5081), .A2(n5082), .ZN(n4442) );
  INV_X1 U6078 ( .A(n5009), .ZN(n4443) );
  OAI211_X1 U6079 ( .C1(n6203), .C2(n4413), .A(n4445), .B(n6216), .ZN(P1_U3220) );
  NAND2_X1 U6080 ( .A1(n6203), .A2(n4405), .ZN(n4445) );
  NAND2_X2 U6081 ( .A1(n9023), .A2(n9026), .ZN(n9037) );
  AND2_X2 U6082 ( .A1(n4449), .A2(n4789), .ZN(n4788) );
  NAND2_X1 U6083 ( .A1(n5361), .A2(n4449), .ZN(n8974) );
  NAND2_X1 U6084 ( .A1(n5360), .A2(n5359), .ZN(n4449) );
  NAND2_X2 U6085 ( .A1(n9016), .A2(n9017), .ZN(n9100) );
  NAND3_X1 U6086 ( .A1(n4783), .A2(n4784), .A3(n5580), .ZN(n4450) );
  NAND2_X1 U6087 ( .A1(n6229), .A2(n6228), .ZN(n6233) );
  NAND2_X1 U6088 ( .A1(n6104), .A2(n6103), .ZN(n4451) );
  NAND2_X1 U6089 ( .A1(n4452), .A2(n5282), .ZN(n5283) );
  INV_X1 U6090 ( .A(n5281), .ZN(n4452) );
  NAND2_X1 U6091 ( .A1(n5281), .A2(SI_11_), .ZN(n4453) );
  OAI21_X1 U6092 ( .B1(n5281), .B2(n4456), .A(n4454), .ZN(n4817) );
  NAND2_X1 U6093 ( .A1(n5280), .A2(n5282), .ZN(n4455) );
  NOR2_X1 U6094 ( .A1(n5280), .A2(n5282), .ZN(n4456) );
  NAND2_X1 U6095 ( .A1(n4807), .A2(n4808), .ZN(n5281) );
  NAND2_X1 U6096 ( .A1(n5340), .A2(n5339), .ZN(n5364) );
  NAND3_X1 U6097 ( .A1(n4460), .A2(n4621), .A3(n4408), .ZN(n4459) );
  NAND3_X1 U6098 ( .A1(n4464), .A2(n4388), .A3(n7830), .ZN(n4463) );
  NAND2_X1 U6099 ( .A1(n5635), .A2(n5634), .ZN(n5637) );
  NAND2_X1 U6100 ( .A1(n9367), .A2(n6313), .ZN(n4874) );
  NAND2_X1 U6101 ( .A1(n4480), .A2(n4922), .ZN(n4479) );
  NAND2_X2 U6102 ( .A1(n5726), .A2(n9691), .ZN(n5026) );
  NAND2_X1 U6103 ( .A1(n5062), .A2(n5061), .ZN(n4491) );
  NAND2_X1 U6104 ( .A1(n7115), .A2(n7707), .ZN(n7327) );
  NAND2_X1 U6105 ( .A1(n6340), .A2(n6339), .ZN(n7886) );
  NAND2_X1 U6106 ( .A1(n5131), .A2(n5130), .ZN(n4514) );
  NAND3_X1 U6107 ( .A1(n4796), .A2(n4794), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n4495) );
  OAI21_X1 U6108 ( .B1(n5817), .B2(n4497), .A(n4496), .ZN(n5003) );
  NAND2_X1 U6109 ( .A1(n7778), .A2(n4502), .ZN(n4499) );
  NAND2_X1 U6110 ( .A1(n9311), .A2(n7851), .ZN(n9300) );
  NAND3_X1 U6111 ( .A1(n9311), .A2(n4502), .A3(n7831), .ZN(n4500) );
  NAND4_X1 U6112 ( .A1(n7694), .A2(n7677), .A3(n7678), .A4(n7706), .ZN(n7802)
         );
  NAND3_X1 U6113 ( .A1(n6355), .A2(n4738), .A3(n4364), .ZN(n6364) );
  AOI21_X1 U6114 ( .B1(n8375), .B2(n4531), .A(n4526), .ZN(n8382) );
  NAND2_X1 U6115 ( .A1(n4524), .A2(n8383), .ZN(n8385) );
  NAND3_X1 U6116 ( .A1(n8375), .A2(n4531), .A3(n4529), .ZN(n4528) );
  NAND3_X1 U6117 ( .A1(n4912), .A2(n4798), .A3(n4536), .ZN(n4535) );
  AOI21_X1 U6118 ( .B1(n4545), .B2(n8595), .A(n4542), .ZN(n8641) );
  NAND2_X1 U6119 ( .A1(n8632), .A2(n8631), .ZN(n4548) );
  OAI21_X1 U6120 ( .B1(n8621), .B2(n8642), .A(n4549), .ZN(P2_U3200) );
  AOI21_X1 U6121 ( .B1(n4553), .B2(n8595), .A(n4550), .ZN(n4549) );
  NAND2_X1 U6122 ( .A1(n8620), .A2(n8624), .ZN(n4551) );
  XNOR2_X1 U6123 ( .A(n8632), .B(n8631), .ZN(n4553) );
  NAND2_X1 U6124 ( .A1(n6102), .A2(n4555), .ZN(n4554) );
  OAI211_X1 U6125 ( .C1(n6102), .C2(n4559), .A(n4557), .B(n4554), .ZN(n6244)
         );
  NAND2_X1 U6126 ( .A1(n6102), .A2(n6101), .ZN(n6227) );
  NAND2_X1 U6127 ( .A1(n9891), .A2(n4562), .ZN(n5836) );
  XNOR2_X1 U6128 ( .A(n7207), .B(n9891), .ZN(n7059) );
  INV_X1 U6129 ( .A(n9891), .ZN(n4564) );
  NAND2_X1 U6130 ( .A1(n8741), .A2(n4568), .ZN(n4565) );
  NAND2_X1 U6131 ( .A1(n4565), .A2(n4566), .ZN(n6061) );
  OAI21_X2 U6132 ( .B1(n8752), .B2(n4577), .A(n4576), .ZN(n4575) );
  NAND2_X4 U6133 ( .A1(n5832), .A2(n6389), .ZN(n8222) );
  NAND2_X1 U6134 ( .A1(n8691), .A2(n4586), .ZN(n4580) );
  OR2_X2 U6135 ( .A1(n8691), .A2(n6068), .ZN(n4588) );
  INV_X1 U6136 ( .A(n6142), .ZN(n5757) );
  NAND4_X1 U6137 ( .A1(n4589), .A2(n5755), .A3(n4351), .A4(n4677), .ZN(n6142)
         );
  AND3_X2 U6138 ( .A1(n4589), .A2(n4351), .A3(n4677), .ZN(n5798) );
  NAND3_X1 U6139 ( .A1(n4677), .A2(n4351), .A3(n4866), .ZN(n6003) );
  OAI21_X2 U6140 ( .B1(n6529), .B2(n5827), .A(n5947), .ZN(n8825) );
  NAND2_X1 U6141 ( .A1(n7390), .A2(n4591), .ZN(n7492) );
  INV_X1 U6142 ( .A(n6330), .ZN(n6539) );
  NOR2_X1 U6143 ( .A1(n7805), .A2(n6330), .ZN(n7807) );
  OAI21_X1 U6144 ( .B1(n6330), .B2(n6544), .A(n6543), .ZN(n9835) );
  OR2_X1 U6145 ( .A1(n7700), .A2(n7698), .ZN(n4604) );
  OR2_X1 U6146 ( .A1(n7691), .A2(n4600), .ZN(n4599) );
  OR2_X1 U6147 ( .A1(n7700), .A2(n4416), .ZN(n4597) );
  OR2_X1 U6148 ( .A1(n7691), .A2(n7689), .ZN(n4605) );
  NAND3_X1 U6149 ( .A1(n4599), .A2(n4597), .A3(n4595), .ZN(n7714) );
  NAND3_X1 U6150 ( .A1(n4605), .A2(n4604), .A3(n4606), .ZN(n7708) );
  NAND3_X1 U6151 ( .A1(n4619), .A2(n9406), .A3(n4618), .ZN(n4617) );
  NAND3_X1 U6152 ( .A1(n7750), .A2(n7790), .A3(n7749), .ZN(n4618) );
  NAND2_X1 U6153 ( .A1(n4938), .A2(n4624), .ZN(n9679) );
  NAND2_X1 U6154 ( .A1(n4938), .A2(n4623), .ZN(n4685) );
  NAND2_X1 U6155 ( .A1(n4938), .A2(n4937), .ZN(n4989) );
  NAND2_X1 U6156 ( .A1(n7277), .A2(n4628), .ZN(n4627) );
  NAND2_X1 U6157 ( .A1(n7276), .A2(n8311), .ZN(n7271) );
  NAND2_X1 U6158 ( .A1(n7559), .A2(n4406), .ZN(n4636) );
  NAND2_X1 U6159 ( .A1(n8727), .A2(n4645), .ZN(n4644) );
  NAND2_X1 U6160 ( .A1(n4656), .A2(n4657), .ZN(n8230) );
  NAND2_X1 U6161 ( .A1(n8670), .A2(n4659), .ZN(n4656) );
  NAND2_X1 U6162 ( .A1(n8670), .A2(n8408), .ZN(n4666) );
  NAND2_X1 U6163 ( .A1(n6178), .A2(n4674), .ZN(n7529) );
  NAND2_X1 U6164 ( .A1(n7529), .A2(n8303), .ZN(n6179) );
  NAND4_X1 U6165 ( .A1(n4857), .A2(n5807), .A3(n5846), .A4(n5743), .ZN(n4676)
         );
  NAND3_X1 U6166 ( .A1(n4857), .A2(n5807), .A3(n5846), .ZN(n4679) );
  NAND2_X1 U6167 ( .A1(n5757), .A2(n5756), .ZN(n5761) );
  OAI21_X1 U6168 ( .B1(n9702), .B2(n5989), .A(n5988), .ZN(n8797) );
  NAND2_X1 U6169 ( .A1(n5934), .A2(n5933), .ZN(n9702) );
  NAND2_X2 U6170 ( .A1(n8743), .A2(n8742), .ZN(n8741) );
  AND2_X4 U6171 ( .A1(n5792), .A2(n8962), .ZN(n5839) );
  OR2_X1 U6172 ( .A1(n8222), .A2(n6387), .ZN(n5810) );
  NAND2_X1 U6173 ( .A1(n8279), .A2(n8281), .ZN(n6176) );
  NAND2_X1 U6174 ( .A1(n5026), .A2(n4686), .ZN(n4687) );
  INV_X1 U6175 ( .A(n4688), .ZN(n7366) );
  NAND2_X1 U6176 ( .A1(n9331), .A2(n4697), .ZN(n7944) );
  NAND2_X1 U6177 ( .A1(n9331), .A2(n9643), .ZN(n9319) );
  INV_X1 U6178 ( .A(n4707), .ZN(n9447) );
  NAND3_X1 U6179 ( .A1(n4797), .A2(n4709), .A3(n4708), .ZN(n4796) );
  NAND2_X1 U6180 ( .A1(n4725), .A2(n4801), .ZN(n5202) );
  NAND3_X1 U6181 ( .A1(n4727), .A2(n5188), .A3(n4726), .ZN(n7706) );
  NAND2_X1 U6182 ( .A1(n6421), .A2(n7781), .ZN(n4727) );
  OAI21_X1 U6183 ( .B1(n9457), .B2(n4732), .A(n4729), .ZN(n6345) );
  NAND2_X1 U6184 ( .A1(n6354), .A2(n9503), .ZN(n4738) );
  AND2_X1 U6185 ( .A1(n4738), .A2(n6353), .ZN(n9289) );
  NAND2_X1 U6186 ( .A1(n4749), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4747) );
  INV_X1 U6187 ( .A(n4756), .ZN(n8600) );
  NAND4_X1 U6188 ( .A1(n4991), .A2(n4990), .A3(n4872), .A4(n4923), .ZN(n5161)
         );
  OAI21_X1 U6189 ( .B1(n9037), .B2(n4766), .A(n4765), .ZN(n9068) );
  INV_X1 U6190 ( .A(n9037), .ZN(n4764) );
  NAND2_X1 U6191 ( .A1(n4770), .A2(n5118), .ZN(n6831) );
  NAND2_X1 U6192 ( .A1(n9055), .A2(n4779), .ZN(n4770) );
  OAI211_X2 U6193 ( .C1(n9055), .C2(n4774), .A(n4773), .B(n4771), .ZN(n6909)
         );
  NAND2_X1 U6194 ( .A1(n4772), .A2(n5118), .ZN(n4771) );
  INV_X1 U6195 ( .A(n4779), .ZN(n4772) );
  NAND2_X1 U6196 ( .A1(n4777), .A2(n4775), .ZN(n4773) );
  NOR2_X1 U6197 ( .A1(n5118), .A2(n4775), .ZN(n4774) );
  NAND2_X1 U6198 ( .A1(n4779), .A2(n4778), .ZN(n4777) );
  OR2_X1 U6199 ( .A1(n5095), .A2(n5096), .ZN(n4779) );
  NAND2_X1 U6200 ( .A1(n4970), .A2(n4780), .ZN(n4984) );
  INV_X1 U6201 ( .A(n8987), .ZN(n4782) );
  NAND3_X1 U6202 ( .A1(n5553), .A2(n8987), .A3(n4414), .ZN(n4784) );
  NOR2_X2 U6203 ( .A1(n4788), .A2(n5362), .ZN(n5382) );
  OAI21_X1 U6204 ( .B1(n7405), .B2(n5311), .A(n4792), .ZN(n4793) );
  INV_X1 U6205 ( .A(n4793), .ZN(n7478) );
  NAND3_X1 U6206 ( .A1(n4795), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4794) );
  NAND2_X1 U6207 ( .A1(n5314), .A2(n5313), .ZN(n5319) );
  NAND3_X1 U6208 ( .A1(n5284), .A2(n5283), .A3(n4818), .ZN(n5314) );
  NAND2_X1 U6209 ( .A1(n5284), .A2(n5283), .ZN(n5287) );
  NAND2_X1 U6210 ( .A1(n5392), .A2(n5391), .ZN(n5418) );
  NAND3_X1 U6211 ( .A1(n5392), .A2(n5391), .A3(n4428), .ZN(n4819) );
  NAND2_X1 U6212 ( .A1(n6166), .A2(n4835), .ZN(n4829) );
  OR2_X1 U6213 ( .A1(n6166), .A2(n4837), .ZN(n4831) );
  NAND2_X1 U6214 ( .A1(n8192), .A2(n4411), .ZN(n4838) );
  OAI211_X1 U6215 ( .C1(n8192), .C2(n4843), .A(n4839), .B(n4838), .ZN(n8037)
         );
  NAND2_X1 U6216 ( .A1(n8192), .A2(n8189), .ZN(n4845) );
  NAND2_X1 U6217 ( .A1(n4852), .A2(n4853), .ZN(n7614) );
  NAND2_X1 U6218 ( .A1(n7545), .A2(n4854), .ZN(n4852) );
  NAND2_X1 U6219 ( .A1(n4860), .A2(n4858), .ZN(n8013) );
  NAND2_X1 U6220 ( .A1(n7456), .A2(n4861), .ZN(n7521) );
  OR2_X1 U6221 ( .A1(n7457), .A2(n7461), .ZN(n4863) );
  NAND2_X1 U6222 ( .A1(n8046), .A2(n4864), .ZN(n8202) );
  AND2_X2 U6223 ( .A1(n5798), .A2(n4868), .ZN(n6135) );
  NAND3_X1 U6224 ( .A1(n4872), .A2(n4990), .A3(n4991), .ZN(n5134) );
  NAND2_X1 U6225 ( .A1(n4873), .A2(n4410), .ZN(n9290) );
  NAND2_X1 U6226 ( .A1(n4874), .A2(n4875), .ZN(n6316) );
  NAND2_X1 U6227 ( .A1(n4888), .A2(n4889), .ZN(n9386) );
  NAND2_X1 U6228 ( .A1(n4931), .A2(n4892), .ZN(n4962) );
  OAI21_X1 U6229 ( .B1(n6203), .B2(n5715), .A(n9115), .ZN(n5742) );
  AOI21_X1 U6230 ( .B1(n9104), .B2(n5692), .A(n5691), .ZN(n5715) );
  INV_X1 U6231 ( .A(n9398), .ZN(n9421) );
  NAND2_X1 U6232 ( .A1(n7138), .A2(n5835), .ZN(n6845) );
  NAND2_X1 U6233 ( .A1(n5811), .A2(n5821), .ZN(n7139) );
  OR2_X1 U6234 ( .A1(n5026), .A2(n6445), .ZN(n5065) );
  XNOR2_X1 U6235 ( .A(n6227), .B(n4661), .ZN(n6133) );
  AND2_X1 U6236 ( .A1(n7869), .A2(n7868), .ZN(n7871) );
  NAND2_X1 U6237 ( .A1(n5839), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5806) );
  OR2_X1 U6238 ( .A1(n9535), .A2(n9625), .ZN(n9542) );
  NOR2_X2 U6239 ( .A1(n6525), .A2(n5053), .ZN(n7962) );
  AND2_X1 U6240 ( .A1(n5052), .A2(n5139), .ZN(n5053) );
  CLKBUF_X1 U6241 ( .A(n6373), .Z(n7503) );
  NAND2_X1 U6242 ( .A1(n7934), .A2(n7933), .ZN(n7941) );
  XNOR2_X1 U6243 ( .A(n8215), .B(n8418), .ZN(n8657) );
  XNOR2_X1 U6244 ( .A(n4988), .B(n9681), .ZN(n5726) );
  NAND2_X1 U6245 ( .A1(n8055), .A2(n8694), .ZN(n8114) );
  XNOR2_X1 U6246 ( .A(n8014), .B(n8015), .ZN(n8055) );
  XNOR2_X1 U6247 ( .A(n6138), .B(n6137), .ZN(n6148) );
  NAND2_X1 U6248 ( .A1(n6140), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U6249 ( .A1(n8013), .A2(n8148), .ZN(n8014) );
  OR2_X1 U6250 ( .A1(n5037), .A2(n5047), .ZN(n4911) );
  XNOR2_X1 U6251 ( .A(n5248), .B(n4373), .ZN(n6425) );
  AOI22_X2 U6252 ( .A1(n7961), .A2(n7962), .B1(n5056), .B2(n5055), .ZN(n6549)
         );
  INV_X1 U6253 ( .A(n8314), .ZN(n5897) );
  INV_X1 U6254 ( .A(n8461), .ZN(n7519) );
  INV_X1 U6255 ( .A(n5718), .ZN(n7870) );
  INV_X1 U6256 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5290) );
  INV_X1 U6257 ( .A(n7991), .ZN(n8779) );
  AND4_X1 U6258 ( .A1(n6036), .A2(n6035), .A3(n6034), .A4(n6033), .ZN(n7991)
         );
  AND2_X1 U6259 ( .A1(n5093), .A2(n5092), .ZN(n4904) );
  AND2_X1 U6260 ( .A1(n6279), .A2(n6278), .ZN(n4905) );
  AND2_X1 U6261 ( .A1(n6188), .A2(n6187), .ZN(n4906) );
  INV_X1 U6262 ( .A(n8817), .ZN(n9708) );
  OR2_X1 U6263 ( .A1(n6170), .A2(n6123), .ZN(n8817) );
  AND2_X1 U6264 ( .A1(n5339), .A2(n5318), .ZN(n4907) );
  AND2_X1 U6265 ( .A1(n5226), .A2(n5184), .ZN(n4908) );
  AND2_X1 U6266 ( .A1(n5349), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4909) );
  INV_X1 U6267 ( .A(n6695), .ZN(n6682) );
  INV_X1 U6268 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5006) );
  AND2_X1 U6269 ( .A1(n5073), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4910) );
  AND2_X1 U6270 ( .A1(n6389), .A2(P1_U3086), .ZN(n7582) );
  AND2_X2 U6271 ( .A1(n4381), .A2(n5028), .ZN(n6328) );
  AND2_X2 U6272 ( .A1(n6263), .A2(n6253), .ZN(n9950) );
  NOR2_X1 U6273 ( .A1(n8442), .A2(n8441), .ZN(n4912) );
  OR2_X1 U6274 ( .A1(n8833), .A2(n8238), .ZN(n4913) );
  NOR2_X1 U6275 ( .A1(n5360), .A2(n5359), .ZN(n5362) );
  AND2_X1 U6276 ( .A1(n6280), .A2(n4905), .ZN(n4914) );
  AND2_X1 U6277 ( .A1(n6272), .A2(n4918), .ZN(n4915) );
  AND2_X1 U6278 ( .A1(n6189), .A2(n4906), .ZN(n4916) );
  AND3_X1 U6279 ( .A1(n6205), .A2(n6204), .A3(n9115), .ZN(n4917) );
  AND2_X1 U6280 ( .A1(n6271), .A2(n6270), .ZN(n4918) );
  AND2_X1 U6281 ( .A1(n7609), .A2(n7608), .ZN(n4919) );
  OR2_X1 U6282 ( .A1(n5275), .A2(n7507), .ZN(n4920) );
  AND2_X1 U6283 ( .A1(n6282), .A2(n8944), .ZN(n4921) );
  NAND2_X1 U6284 ( .A1(n9388), .A2(n9408), .ZN(n4922) );
  NAND2_X1 U6285 ( .A1(n8833), .A2(n8227), .ZN(n8225) );
  NAND2_X1 U6286 ( .A1(n8188), .A2(n7991), .ZN(n6037) );
  OR4_X1 U6287 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5705) );
  INV_X1 U6288 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4956) );
  OR2_X1 U6289 ( .A1(n8158), .A2(n8458), .ZN(n7608) );
  AOI21_X1 U6290 ( .B1(n8432), .B2(n8422), .A(n8421), .ZN(n8425) );
  NAND2_X1 U6291 ( .A1(n5983), .A2(n7565), .ZN(n5984) );
  INV_X1 U6292 ( .A(n5820), .ZN(n5821) );
  INV_X1 U6293 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5750) );
  INV_X1 U6294 ( .A(SI_14_), .ZN(n10168) );
  OR2_X1 U6295 ( .A1(n7593), .A2(n7592), .ZN(n7594) );
  AND2_X1 U6296 ( .A1(n8437), .A2(n8433), .ZN(n8236) );
  OR2_X1 U6297 ( .A1(n9716), .A2(n6269), .ZN(n6270) );
  INV_X1 U6298 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10059) );
  INV_X1 U6299 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7438) );
  NAND2_X1 U6300 ( .A1(n6277), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U6301 ( .A1(n9939), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U6302 ( .A1(n5985), .A2(n5984), .ZN(n9703) );
  OR2_X1 U6303 ( .A1(n6249), .A2(n6163), .ZN(n6930) );
  OR2_X1 U6304 ( .A1(n5026), .A2(n6447), .ZN(n5027) );
  NOR2_X1 U6305 ( .A1(n5270), .A2(n5269), .ZN(n5271) );
  OAI211_X1 U6306 ( .C1(n7300), .C2(n5224), .A(n5223), .B(n5222), .ZN(n6373)
         );
  INV_X1 U6307 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5541) );
  INV_X1 U6308 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5326) );
  INV_X1 U6309 ( .A(SI_26_), .ZN(n10164) );
  INV_X1 U6310 ( .A(SI_23_), .ZN(n5557) );
  INV_X1 U6311 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4980) );
  INV_X1 U6312 ( .A(SI_15_), .ZN(n10155) );
  INV_X1 U6313 ( .A(SI_9_), .ZN(n10173) );
  INV_X1 U6314 ( .A(n7020), .ZN(n7207) );
  NAND2_X1 U6315 ( .A1(n7518), .A2(n7519), .ZN(n7520) );
  INV_X1 U6316 ( .A(n5840), .ZN(n5786) );
  INV_X1 U6317 ( .A(n8493), .ZN(n8494) );
  INV_X1 U6318 ( .A(n8523), .ZN(n8524) );
  INV_X1 U6319 ( .A(n6056), .ZN(n5779) );
  AND2_X1 U6320 ( .A1(n6185), .A2(n6978), .ZN(n7282) );
  OR2_X1 U6321 ( .A1(n6147), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6150) );
  INV_X1 U6322 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5350) );
  INV_X1 U6323 ( .A(n5564), .ZN(n5563) );
  OR2_X1 U6324 ( .A1(n5542), .A2(n5541), .ZN(n5564) );
  OR2_X1 U6325 ( .A1(n5465), .A2(n9092), .ZN(n5467) );
  INV_X1 U6326 ( .A(n5057), .ZN(n5017) );
  OR2_X1 U6327 ( .A1(n5259), .A2(n5237), .ZN(n5296) );
  INV_X1 U6328 ( .A(n9141), .ZN(n6290) );
  AND2_X1 U6329 ( .A1(n6326), .A2(n6636), .ZN(n6327) );
  OAI21_X1 U6330 ( .B1(n5507), .B2(n10170), .A(n5506), .ZN(n5509) );
  OR2_X1 U6331 ( .A1(n5290), .A2(n4980), .ZN(n4981) );
  OR2_X1 U6332 ( .A1(n5249), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5289) );
  INV_X1 U6333 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U6334 ( .A1(n7975), .A2(n7974), .ZN(n8138) );
  INV_X1 U6335 ( .A(n8463), .ZN(n7294) );
  NAND2_X1 U6336 ( .A1(n5787), .A2(n5791), .ZN(n5812) );
  INV_X1 U6337 ( .A(n8565), .ZN(n8526) );
  INV_X1 U6338 ( .A(n6131), .ZN(n8445) );
  OR2_X1 U6339 ( .A1(n6064), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6072) );
  INV_X1 U6340 ( .A(n8768), .ZN(n8788) );
  INV_X1 U6341 ( .A(n8811), .ZN(n8328) );
  AND2_X1 U6342 ( .A1(n8412), .A2(n6251), .ZN(n6258) );
  INV_X1 U6343 ( .A(n8455), .ZN(n9711) );
  AND2_X1 U6344 ( .A1(n8332), .A2(n8331), .ZN(n8256) );
  AND2_X1 U6345 ( .A1(n8294), .A2(n8313), .ZN(n8249) );
  INV_X1 U6346 ( .A(n7282), .ZN(n6267) );
  OR2_X1 U6347 ( .A1(n7023), .A2(n8412), .ZN(n9712) );
  OR2_X1 U6348 ( .A1(n5351), .A2(n5350), .ZN(n5374) );
  INV_X1 U6349 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9001) );
  OR2_X1 U6350 ( .A1(n5617), .A2(n5616), .ZN(n5645) );
  NAND2_X1 U6351 ( .A1(n5563), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5617) );
  INV_X1 U6352 ( .A(n4352), .ZN(n6466) );
  INV_X1 U6353 ( .A(n7823), .ZN(n9472) );
  NAND2_X1 U6354 ( .A1(n7711), .A2(n7893), .ZN(n7225) );
  OR2_X1 U6355 ( .A1(n7795), .A2(n7798), .ZN(n7861) );
  INV_X1 U6356 ( .A(n9876), .ZN(n6362) );
  INV_X1 U6357 ( .A(n9871), .ZN(n6369) );
  INV_X1 U6358 ( .A(n9623), .ZN(n9866) );
  INV_X1 U6359 ( .A(n9524), .ZN(n9380) );
  NAND3_X1 U6360 ( .A1(n5046), .A2(n6408), .A3(P1_STATE_REG_SCAN_IN), .ZN(
        n7936) );
  INV_X1 U6361 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9681) );
  AOI21_X1 U6362 ( .B1(n7542), .B2(n7541), .A(n7540), .ZN(n7545) );
  AND2_X1 U6363 ( .A1(n7024), .A2(n7023), .ZN(n8205) );
  AOI22_X1 U6364 ( .A1(n7291), .A2(n7290), .B1(n7294), .B2(n7289), .ZN(n7293)
         );
  INV_X1 U6365 ( .A(n8638), .ZN(n8443) );
  INV_X1 U6366 ( .A(n9886), .ZN(n8559) );
  INV_X1 U6367 ( .A(n8635), .ZN(n8595) );
  INV_X1 U6368 ( .A(n9712), .ZN(n8819) );
  INV_X1 U6369 ( .A(n9697), .ZN(n8805) );
  INV_X1 U6370 ( .A(n9950), .ZN(n6277) );
  INV_X1 U6371 ( .A(n8855), .ZN(n8874) );
  AND2_X1 U6372 ( .A1(n6249), .A2(n6248), .ZN(n6263) );
  AND2_X1 U6373 ( .A1(n8386), .A2(n8378), .ZN(n8731) );
  INV_X1 U6374 ( .A(n9925), .ZN(n9932) );
  AND2_X1 U6375 ( .A1(n7552), .A2(n6266), .ZN(n9907) );
  OR2_X1 U6376 ( .A1(n6922), .A2(n6171), .ZN(n6174) );
  AND2_X1 U6377 ( .A1(n5972), .A2(n5990), .ZN(n8515) );
  OAI21_X1 U6378 ( .B1(n9643), .B2(n9124), .A(n5739), .ZN(n5740) );
  INV_X1 U6379 ( .A(n9121), .ZN(n9107) );
  OAI21_X2 U6380 ( .B1(n6520), .B2(n5083), .A(n5291), .ZN(n9622) );
  INV_X1 U6381 ( .A(n5478), .ZN(n9089) );
  OR2_X1 U6382 ( .A1(n5716), .A2(n6619), .ZN(n5717) );
  AND2_X1 U6383 ( .A1(n5408), .A2(n5407), .ZN(n9517) );
  INV_X1 U6384 ( .A(n9808), .ZN(n9786) );
  OR2_X1 U6385 ( .A1(n9749), .A2(n6466), .ZN(n9790) );
  INV_X1 U6386 ( .A(n9790), .ZN(n9811) );
  INV_X1 U6387 ( .A(n9798), .ZN(n9815) );
  AND2_X1 U6388 ( .A1(n7725), .A2(n7722), .ZN(n7821) );
  INV_X1 U6389 ( .A(n9529), .ZN(n9836) );
  INV_X1 U6390 ( .A(n9841), .ZN(n9527) );
  AOI21_X1 U6391 ( .B1(n6416), .B2(n5699), .A(n6420), .ZN(n6367) );
  NOR2_X1 U6392 ( .A1(n6361), .A2(n6610), .ZN(n6368) );
  INV_X1 U6393 ( .A(n8210), .ZN(n8183) );
  AND2_X1 U6394 ( .A1(n8235), .A2(n6129), .ZN(n8034) );
  INV_X1 U6395 ( .A(n8068), .ZN(n8754) );
  OR2_X1 U6396 ( .A1(P2_U3150), .A2(n6660), .ZN(n8618) );
  OR2_X1 U6397 ( .A1(n9878), .A2(n8444), .ZN(n8642) );
  AND2_X1 U6398 ( .A1(n8801), .A2(n8800), .ZN(n9722) );
  INV_X1 U6399 ( .A(n9716), .ZN(n9718) );
  NAND2_X1 U6400 ( .A1(n9716), .A2(n9715), .ZN(n8795) );
  NAND2_X1 U6401 ( .A1(n9950), .A2(n9933), .ZN(n8881) );
  NAND2_X1 U6402 ( .A1(n9950), .A2(n9932), .ZN(n8855) );
  NOR2_X1 U6403 ( .A1(n4921), .A2(n6284), .ZN(n6285) );
  NAND2_X1 U6404 ( .A1(n9937), .A2(n9933), .ZN(n8952) );
  INV_X1 U6405 ( .A(n8944), .ZN(n8907) );
  AND2_X1 U6406 ( .A1(n6174), .A2(n6173), .ZN(n9939) );
  INV_X2 U6407 ( .A(n9939), .ZN(n9937) );
  NAND2_X1 U6408 ( .A1(n6147), .A2(n6517), .ZN(n6577) );
  INV_X1 U6409 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8972) );
  INV_X1 U6410 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7553) );
  INV_X1 U6411 ( .A(n8515), .ZN(n8529) );
  NAND2_X1 U6412 ( .A1(n6388), .A2(P2_U3151), .ZN(n8960) );
  NOR2_X1 U6413 ( .A1(n4917), .A2(n6215), .ZN(n6216) );
  INV_X1 U6414 ( .A(n9560), .ZN(n9370) );
  INV_X1 U6415 ( .A(n9115), .ZN(n9098) );
  AND2_X1 U6416 ( .A1(n5717), .A2(n9390), .ZN(n9124) );
  INV_X1 U6417 ( .A(n9315), .ZN(n9127) );
  INV_X1 U6418 ( .A(n9517), .ZN(n9475) );
  OR2_X1 U6419 ( .A1(n9749), .A2(n9158), .ZN(n9798) );
  OR2_X1 U6420 ( .A1(n9749), .A2(n9738), .ZN(n9808) );
  OR2_X1 U6421 ( .A1(n9826), .A2(n6619), .ZN(n9514) );
  INV_X1 U6422 ( .A(n6606), .ZN(n9633) );
  AND2_X2 U6423 ( .A1(n6368), .A2(n6367), .ZN(n9876) );
  INV_X1 U6424 ( .A(n9388), .ZN(n9652) );
  INV_X1 U6425 ( .A(n6572), .ZN(n9676) );
  AND2_X2 U6426 ( .A1(n6368), .A2(n6613), .ZN(n9871) );
  AND2_X1 U6427 ( .A1(n7591), .A2(n7634), .ZN(n6420) );
  OR2_X1 U6428 ( .A1(n6408), .A2(P1_U3086), .ZN(n7931) );
  INV_X1 U6429 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U6430 ( .A1(n6388), .A2(P1_U3086), .ZN(n9694) );
  NAND2_X1 U6431 ( .A1(n6190), .A2(n4916), .ZN(P2_U3455) );
  AND2_X1 U6432 ( .A1(n6372), .A2(n6408), .ZN(P1_U3973) );
  INV_X1 U6433 ( .A(n5161), .ZN(n4929) );
  NOR2_X1 U6434 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4927) );
  NOR2_X1 U6435 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4926) );
  NOR2_X1 U6436 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4925) );
  NOR2_X1 U6437 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4924) );
  NAND2_X1 U6438 ( .A1(n4929), .A2(n4928), .ZN(n5368) );
  NOR2_X1 U6439 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4934) );
  NOR2_X1 U6440 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4933) );
  NOR2_X1 U6441 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4932) );
  NAND4_X1 U6442 ( .A1(n4935), .A2(n4934), .A3(n4933), .A4(n4932), .ZN(n4936)
         );
  NAND2_X1 U6443 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n4940) );
  NAND2_X1 U6444 ( .A1(n4988), .A2(n4940), .ZN(n4941) );
  INV_X1 U6445 ( .A(n4946), .ZN(n4942) );
  INV_X1 U6446 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6618) );
  INV_X1 U6447 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n4943) );
  OR2_X1 U6448 ( .A1(n5452), .A2(n4943), .ZN(n4944) );
  OAI21_X1 U6449 ( .B1(n7655), .B2(n6618), .A(n4944), .ZN(n4945) );
  INV_X1 U6450 ( .A(n4945), .ZN(n4953) );
  INV_X1 U6451 ( .A(n4948), .ZN(n4947) );
  NAND2_X2 U6452 ( .A1(n4942), .A2(n4947), .ZN(n5057) );
  NAND2_X1 U6453 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5100) );
  OAI21_X1 U6454 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n5100), .ZN(n9061) );
  INV_X1 U6455 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n4949) );
  OAI21_X1 U6456 ( .B1(n5057), .B2(n9061), .A(n4950), .ZN(n4951) );
  INV_X1 U6457 ( .A(n4951), .ZN(n4952) );
  NAND2_X1 U6458 ( .A1(n4955), .A2(n4954), .ZN(n4977) );
  NAND3_X1 U6459 ( .A1(n4980), .A2(n4978), .A3(n4956), .ZN(n4957) );
  NOR2_X2 U6460 ( .A1(n4977), .A2(n4957), .ZN(n4970) );
  NAND2_X1 U6461 ( .A1(n4962), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U6462 ( .A1(n4365), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4965) );
  INV_X1 U6463 ( .A(n7628), .ZN(n4966) );
  INV_X1 U6464 ( .A(n5712), .ZN(n4976) );
  INV_X1 U6465 ( .A(n4970), .ZN(n4971) );
  NAND2_X1 U6466 ( .A1(n4971), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4972) );
  INV_X1 U6467 ( .A(n4973), .ZN(n4974) );
  INV_X1 U6468 ( .A(n5014), .ZN(n5013) );
  NAND2_X1 U6469 ( .A1(n4977), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6470 ( .A1(n5422), .A2(n4978), .ZN(n4979) );
  NAND2_X1 U6471 ( .A1(n5013), .A2(n9269), .ZN(n6946) );
  INV_X2 U6472 ( .A(n4983), .ZN(n7866) );
  NAND2_X1 U6473 ( .A1(n5713), .A2(n7795), .ZN(n4987) );
  OR2_X1 U6474 ( .A1(n4990), .A2(n5290), .ZN(n5064) );
  OR2_X1 U6475 ( .A1(n4991), .A2(n5290), .ZN(n4992) );
  AND2_X1 U6476 ( .A1(n5064), .A2(n4992), .ZN(n4994) );
  INV_X1 U6477 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6478 ( .A1(n4994), .A2(n4993), .ZN(n5107) );
  INV_X1 U6479 ( .A(n4994), .ZN(n4995) );
  NAND2_X1 U6480 ( .A1(n4995), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U6481 ( .A1(n5107), .A2(n4996), .ZN(n9188) );
  INV_X4 U6482 ( .A(n5817), .ZN(n6389) );
  AND2_X1 U6483 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U6484 ( .A1(n6389), .A2(n4997), .ZN(n5043) );
  NAND3_X1 U6485 ( .A1(n5817), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4998) );
  INV_X1 U6486 ( .A(SI_1_), .ZN(n4999) );
  NAND2_X1 U6487 ( .A1(n5000), .A2(SI_1_), .ZN(n5001) );
  INV_X1 U6488 ( .A(SI_2_), .ZN(n5002) );
  XNOR2_X1 U6489 ( .A(n5003), .B(n5002), .ZN(n5061) );
  NAND2_X1 U6490 ( .A1(n5003), .A2(SI_2_), .ZN(n5004) );
  INV_X1 U6491 ( .A(SI_3_), .ZN(n5007) );
  XNOR2_X1 U6492 ( .A(n5008), .B(n5007), .ZN(n5082) );
  NAND2_X1 U6493 ( .A1(n5008), .A2(SI_3_), .ZN(n5009) );
  MUX2_X1 U6494 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6389), .Z(n5112) );
  INV_X1 U6495 ( .A(SI_4_), .ZN(n5010) );
  XNOR2_X1 U6496 ( .A(n5112), .B(n5010), .ZN(n5110) );
  XNOR2_X1 U6497 ( .A(n5111), .B(n5110), .ZN(n6392) );
  OR2_X1 U6498 ( .A1(n5083), .A2(n6392), .ZN(n5012) );
  INV_X1 U6499 ( .A(n6389), .ZN(n6388) );
  NAND2_X4 U6500 ( .A1(n5026), .A2(n6388), .ZN(n7782) );
  INV_X1 U6501 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6391) );
  OR2_X1 U6502 ( .A1(n7782), .A2(n6391), .ZN(n5011) );
  OAI211_X1 U6503 ( .C1(n5026), .C2(n9188), .A(n5012), .B(n5011), .ZN(n9063)
         );
  INV_X1 U6504 ( .A(n9063), .ZN(n6620) );
  OAI22_X1 U6505 ( .A1(n6290), .A2(n5656), .B1(n6620), .B2(n5167), .ZN(n5094)
         );
  INV_X1 U6506 ( .A(n5094), .ZN(n5096) );
  NAND3_X1 U6508 ( .A1(n6324), .A2(n5046), .A3(n5014), .ZN(n5015) );
  AOI22_X1 U6510 ( .A1(n9141), .A2(n5033), .B1(n9063), .B2(n6193), .ZN(n5016)
         );
  BUF_X4 U6511 ( .A(n5015), .Z(n5628) );
  XNOR2_X1 U6512 ( .A(n5016), .B(n5628), .ZN(n5095) );
  NAND2_X1 U6513 ( .A1(n5017), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5021) );
  INV_X1 U6514 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5018) );
  OR2_X1 U6515 ( .A1(n5035), .A2(n5018), .ZN(n5019) );
  NAND4_X2 U6516 ( .A1(n5022), .A2(n5021), .A3(n5020), .A4(n5019), .ZN(n6487)
         );
  NAND2_X1 U6517 ( .A1(n6487), .A2(n5033), .ZN(n5030) );
  INV_X1 U6518 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6519 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5024) );
  XNOR2_X1 U6520 ( .A(n5025), .B(n5024), .ZN(n6447) );
  INV_X1 U6521 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6398) );
  OR2_X1 U6522 ( .A1(n7782), .A2(n6398), .ZN(n5028) );
  NAND2_X1 U6523 ( .A1(n5030), .A2(n5029), .ZN(n5031) );
  INV_X1 U6524 ( .A(n6487), .ZN(n6535) );
  INV_X1 U6525 ( .A(n5033), .ZN(n5086) );
  INV_X1 U6526 ( .A(n5034), .ZN(n5056) );
  INV_X1 U6527 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5036) );
  INV_X1 U6528 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6529 ( .A1(n6389), .A2(SI_0_), .ZN(n5042) );
  INV_X1 U6530 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5041) );
  NAND2_X1 U6531 ( .A1(n5042), .A2(n5041), .ZN(n5044) );
  AND2_X1 U6532 ( .A1(n5044), .A2(n5043), .ZN(n9695) );
  MUX2_X1 U6533 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9695), .S(n5026), .Z(n6635) );
  AOI22_X1 U6534 ( .A1(n6540), .A2(n5033), .B1(n6635), .B2(n5045), .ZN(n5052)
         );
  OR2_X1 U6535 ( .A1(n5046), .A2(n5047), .ZN(n5048) );
  NAND2_X1 U6536 ( .A1(n5052), .A2(n5048), .ZN(n6523) );
  INV_X1 U6537 ( .A(n5656), .ZN(n5049) );
  NAND2_X1 U6538 ( .A1(n6540), .A2(n5049), .ZN(n5051) );
  INV_X1 U6539 ( .A(n5046), .ZN(n5723) );
  AOI22_X1 U6540 ( .A1(n6635), .A2(n5033), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5723), .ZN(n5050) );
  NAND2_X1 U6541 ( .A1(n5051), .A2(n5050), .ZN(n6522) );
  AND2_X1 U6542 ( .A1(n6523), .A2(n6522), .ZN(n6525) );
  INV_X1 U6543 ( .A(n5054), .ZN(n5055) );
  NAND2_X1 U6544 ( .A1(n5619), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6545 ( .A1(n7651), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5058) );
  NAND3_X1 U6546 ( .A1(n5060), .A2(n5059), .A3(n5058), .ZN(n9143) );
  NAND2_X1 U6547 ( .A1(n9143), .A2(n5033), .ZN(n5069) );
  XNOR2_X1 U6548 ( .A(n5062), .B(n5061), .ZN(n6394) );
  OR2_X1 U6549 ( .A1(n5083), .A2(n6394), .ZN(n5067) );
  OR2_X1 U6550 ( .A1(n7782), .A2(n4497), .ZN(n5066) );
  INV_X1 U6551 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U6552 ( .A1(n5064), .A2(n5063), .ZN(n5078) );
  OAI21_X1 U6553 ( .B1(n5064), .B2(n5063), .A(n5078), .ZN(n6445) );
  AND3_X4 U6554 ( .A1(n5067), .A2(n5066), .A3(n5065), .ZN(n7877) );
  NAND2_X1 U6555 ( .A1(n6551), .A2(n5045), .ZN(n5068) );
  NAND2_X1 U6556 ( .A1(n5069), .A2(n5068), .ZN(n5070) );
  INV_X1 U6557 ( .A(n9143), .ZN(n6557) );
  OAI22_X1 U6558 ( .A1(n6557), .A2(n5656), .B1(n7877), .B2(n5167), .ZN(n5071)
         );
  XNOR2_X1 U6559 ( .A(n5072), .B(n5071), .ZN(n6550) );
  INV_X1 U6560 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U6561 ( .A1(n5619), .A2(n9825), .ZN(n5077) );
  NAND2_X1 U6562 ( .A1(n5349), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U6563 ( .A1(n5073), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6564 ( .A1(n7651), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U6565 ( .A1(n5078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5080) );
  INV_X1 U6566 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5079) );
  XNOR2_X1 U6567 ( .A(n5080), .B(n5079), .ZN(n6451) );
  XNOR2_X1 U6568 ( .A(n5081), .B(n5082), .ZN(n6395) );
  OR2_X1 U6569 ( .A1(n5083), .A2(n6395), .ZN(n5085) );
  INV_X1 U6570 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6390) );
  OR2_X1 U6571 ( .A1(n7782), .A2(n6390), .ZN(n5084) );
  OAI22_X1 U6572 ( .A1(n6536), .A2(n5656), .B1(n6587), .B2(n5167), .ZN(n5091)
         );
  NAND2_X1 U6573 ( .A1(n9142), .A2(n5033), .ZN(n5088) );
  NAND2_X1 U6574 ( .A1(n9824), .A2(n5045), .ZN(n5087) );
  NAND2_X1 U6575 ( .A1(n5088), .A2(n5087), .ZN(n5089) );
  XNOR2_X1 U6576 ( .A(n5089), .B(n5628), .ZN(n5090) );
  XOR2_X1 U6577 ( .A(n5091), .B(n5090), .Z(n6556) );
  INV_X1 U6578 ( .A(n5090), .ZN(n5093) );
  INV_X1 U6579 ( .A(n5091), .ZN(n5092) );
  XNOR2_X1 U6580 ( .A(n5095), .B(n5094), .ZN(n9056) );
  NAND2_X1 U6581 ( .A1(n9057), .A2(n9056), .ZN(n9055) );
  INV_X1 U6582 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6433) );
  INV_X1 U6583 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6455) );
  OR2_X1 U6584 ( .A1(n5452), .A2(n6455), .ZN(n5097) );
  OAI21_X1 U6585 ( .B1(n7655), .B2(n6433), .A(n5097), .ZN(n5098) );
  INV_X1 U6586 ( .A(n5098), .ZN(n5106) );
  INV_X1 U6587 ( .A(n5100), .ZN(n5099) );
  NAND2_X1 U6588 ( .A1(n5099), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5124) );
  INV_X1 U6589 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6834) );
  NAND2_X1 U6590 ( .A1(n5100), .A2(n6834), .ZN(n5101) );
  NAND2_X1 U6591 ( .A1(n5124), .A2(n5101), .ZN(n6756) );
  INV_X1 U6592 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5102) );
  OR2_X1 U6593 ( .A1(n5471), .A2(n5102), .ZN(n5103) );
  OAI21_X1 U6594 ( .B1(n5057), .B2(n6756), .A(n5103), .ZN(n5104) );
  INV_X1 U6595 ( .A(n5104), .ZN(n5105) );
  NAND2_X1 U6596 ( .A1(n5107), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5109) );
  INV_X1 U6597 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5108) );
  XNOR2_X1 U6598 ( .A(n5109), .B(n5108), .ZN(n9201) );
  NAND2_X1 U6599 ( .A1(n5112), .A2(SI_4_), .ZN(n5113) );
  MUX2_X1 U6600 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6389), .Z(n5132) );
  INV_X1 U6601 ( .A(SI_5_), .ZN(n5114) );
  XNOR2_X1 U6602 ( .A(n5132), .B(n5114), .ZN(n5130) );
  XNOR2_X1 U6603 ( .A(n5131), .B(n5130), .ZN(n6399) );
  OR2_X1 U6604 ( .A1(n6399), .A2(n5083), .ZN(n5116) );
  INV_X1 U6605 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6400) );
  OR2_X1 U6606 ( .A1(n7782), .A2(n6400), .ZN(n5115) );
  OAI211_X1 U6607 ( .C1(n5026), .C2(n9201), .A(n5116), .B(n5115), .ZN(n6648)
         );
  AOI22_X1 U6608 ( .A1(n9140), .A2(n5033), .B1(n6648), .B2(n6193), .ZN(n5117)
         );
  XOR2_X1 U6609 ( .A(n5628), .B(n5117), .Z(n5118) );
  AOI22_X1 U6610 ( .A1(n9140), .A2(n5630), .B1(n5681), .B2(n6648), .ZN(n6832)
         );
  INV_X1 U6611 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6435) );
  INV_X1 U6612 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5119) );
  OR2_X1 U6613 ( .A1(n5471), .A2(n5119), .ZN(n5120) );
  OAI21_X1 U6614 ( .B1(n7655), .B2(n6435), .A(n5120), .ZN(n5121) );
  INV_X1 U6615 ( .A(n5121), .ZN(n5129) );
  INV_X1 U6616 ( .A(n5124), .ZN(n5122) );
  NAND2_X1 U6617 ( .A1(n5122), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5149) );
  INV_X1 U6618 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6619 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  NAND2_X1 U6620 ( .A1(n5149), .A2(n5125), .ZN(n6748) );
  INV_X1 U6621 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6457) );
  OR2_X1 U6622 ( .A1(n5452), .A2(n6457), .ZN(n5126) );
  OAI21_X1 U6623 ( .B1(n5057), .B2(n6748), .A(n5126), .ZN(n5127) );
  INV_X1 U6624 ( .A(n5127), .ZN(n5128) );
  NAND2_X1 U6625 ( .A1(n5132), .A2(SI_5_), .ZN(n5133) );
  MUX2_X1 U6626 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6389), .Z(n5158) );
  INV_X1 U6627 ( .A(SI_6_), .ZN(n10074) );
  XNOR2_X1 U6628 ( .A(n5158), .B(n10074), .ZN(n5156) );
  XNOR2_X1 U6629 ( .A(n5157), .B(n5156), .ZN(n6402) );
  OR2_X1 U6630 ( .A1(n6402), .A2(n5083), .ZN(n5137) );
  NAND2_X1 U6631 ( .A1(n5134), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5135) );
  XNOR2_X1 U6632 ( .A(n5135), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9218) );
  AOI22_X1 U6633 ( .A1(n5462), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5461), .B2(
        n9218), .ZN(n5136) );
  NAND2_X1 U6634 ( .A1(n5137), .A2(n5136), .ZN(n6293) );
  NAND2_X1 U6635 ( .A1(n6293), .A2(n6193), .ZN(n5138) );
  OAI21_X1 U6636 ( .B1(n6953), .B2(n5167), .A(n5138), .ZN(n5140) );
  XNOR2_X1 U6637 ( .A(n5140), .B(n5139), .ZN(n6907) );
  AND2_X1 U6638 ( .A1(n6293), .A2(n6197), .ZN(n5141) );
  AOI21_X1 U6639 ( .B1(n9139), .B2(n5630), .A(n5141), .ZN(n6906) );
  NAND2_X1 U6640 ( .A1(n6907), .A2(n6906), .ZN(n5144) );
  INV_X1 U6641 ( .A(n6907), .ZN(n5143) );
  INV_X1 U6642 ( .A(n6906), .ZN(n5142) );
  INV_X1 U6643 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6957) );
  INV_X1 U6644 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5145) );
  OR2_X1 U6645 ( .A1(n5452), .A2(n5145), .ZN(n5146) );
  OAI21_X1 U6646 ( .B1(n7655), .B2(n6957), .A(n5146), .ZN(n5147) );
  INV_X1 U6647 ( .A(n5147), .ZN(n5155) );
  NAND2_X1 U6648 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  NAND2_X1 U6649 ( .A1(n5208), .A2(n5150), .ZN(n7077) );
  INV_X1 U6650 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5151) );
  OR2_X1 U6651 ( .A1(n5471), .A2(n5151), .ZN(n5152) );
  OAI21_X1 U6652 ( .B1(n5057), .B2(n7077), .A(n5152), .ZN(n5153) );
  INV_X1 U6653 ( .A(n5153), .ZN(n5154) );
  NAND2_X1 U6654 ( .A1(n5158), .A2(SI_6_), .ZN(n5159) );
  MUX2_X1 U6655 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6389), .Z(n5174) );
  INV_X1 U6656 ( .A(SI_7_), .ZN(n5160) );
  XNOR2_X1 U6657 ( .A(n5174), .B(n5160), .ZN(n5172) );
  XNOR2_X1 U6658 ( .A(n5173), .B(n5172), .ZN(n6405) );
  OR2_X1 U6659 ( .A1(n6405), .A2(n5083), .ZN(n5165) );
  NAND2_X1 U6660 ( .A1(n5162), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5163) );
  XNOR2_X1 U6661 ( .A(n5163), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9231) );
  AOI22_X1 U6662 ( .A1(n5462), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5461), .B2(
        n9231), .ZN(n5164) );
  NAND2_X1 U6663 ( .A1(n5165), .A2(n5164), .ZN(n6962) );
  NAND2_X1 U6664 ( .A1(n6962), .A2(n6193), .ZN(n5166) );
  OAI21_X1 U6665 ( .B1(n6740), .B2(n5167), .A(n5166), .ZN(n5168) );
  XNOR2_X1 U6666 ( .A(n5168), .B(n5628), .ZN(n5171) );
  NAND2_X1 U6667 ( .A1(n6962), .A2(n5681), .ZN(n5169) );
  OAI21_X1 U6668 ( .B1(n6740), .B2(n5656), .A(n5169), .ZN(n5170) );
  NOR2_X1 U6669 ( .A1(n5171), .A2(n5170), .ZN(n7073) );
  NAND2_X1 U6670 ( .A1(n5171), .A2(n5170), .ZN(n7071) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5175) );
  MUX2_X1 U6672 ( .A(n6413), .B(n5175), .S(n6389), .Z(n5176) );
  NAND2_X1 U6673 ( .A1(n5176), .A2(n10143), .ZN(n5179) );
  INV_X1 U6674 ( .A(n5176), .ZN(n5177) );
  NAND2_X1 U6675 ( .A1(n5177), .A2(SI_8_), .ZN(n5178) );
  NAND2_X1 U6676 ( .A1(n5179), .A2(n5178), .ZN(n5201) );
  INV_X1 U6677 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5181) );
  MUX2_X1 U6678 ( .A(n6423), .B(n5181), .S(n6389), .Z(n5182) );
  NAND2_X1 U6679 ( .A1(n5182), .A2(n10173), .ZN(n5226) );
  INV_X1 U6680 ( .A(n5182), .ZN(n5183) );
  NAND2_X1 U6681 ( .A1(n5183), .A2(SI_9_), .ZN(n5184) );
  XNOR2_X1 U6682 ( .A(n5225), .B(n4908), .ZN(n6421) );
  NOR2_X1 U6683 ( .A1(n5162), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5230) );
  OR2_X1 U6684 ( .A1(n5230), .A2(n5290), .ZN(n5203) );
  INV_X1 U6685 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6686 ( .A1(n5203), .A2(n5185), .ZN(n5186) );
  NAND2_X1 U6687 ( .A1(n5186), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5187) );
  XNOR2_X1 U6688 ( .A(n5187), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6484) );
  AOI22_X1 U6689 ( .A1(n5462), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5461), .B2(
        n6484), .ZN(n5188) );
  INV_X1 U6690 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7043) );
  INV_X1 U6691 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5189) );
  OR2_X1 U6692 ( .A1(n5452), .A2(n5189), .ZN(n5190) );
  OAI21_X1 U6693 ( .B1(n7655), .B2(n7043), .A(n5190), .ZN(n5191) );
  INV_X1 U6694 ( .A(n5191), .ZN(n5198) );
  NAND2_X1 U6695 ( .A1(n5210), .A2(n5192), .ZN(n5193) );
  NAND2_X1 U6696 ( .A1(n5257), .A2(n5193), .ZN(n7381) );
  INV_X1 U6697 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5194) );
  OR2_X1 U6698 ( .A1(n5471), .A2(n5194), .ZN(n5195) );
  OAI21_X1 U6699 ( .B1(n5057), .B2(n7381), .A(n5195), .ZN(n5196) );
  INV_X1 U6700 ( .A(n5196), .ZN(n5197) );
  AOI22_X1 U6701 ( .A1(n7384), .A2(n6193), .B1(n6197), .B2(n4726), .ZN(n5199)
         );
  XNOR2_X1 U6702 ( .A(n5199), .B(n5628), .ZN(n7376) );
  NOR2_X1 U6703 ( .A1(n7306), .A2(n5656), .ZN(n5200) );
  AOI21_X1 U6704 ( .B1(n7384), .B2(n5681), .A(n5200), .ZN(n7375) );
  XNOR2_X1 U6705 ( .A(n5202), .B(n4724), .ZN(n6412) );
  OR2_X1 U6706 ( .A1(n6412), .A2(n5083), .ZN(n5205) );
  XNOR2_X1 U6707 ( .A(n5203), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9244) );
  AOI22_X1 U6708 ( .A1(n5462), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5461), .B2(
        n9244), .ZN(n5204) );
  INV_X1 U6709 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6873) );
  INV_X1 U6710 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6460) );
  OR2_X1 U6711 ( .A1(n5452), .A2(n6460), .ZN(n5206) );
  OAI21_X1 U6712 ( .B1(n7655), .B2(n6873), .A(n5206), .ZN(n5207) );
  INV_X1 U6713 ( .A(n5207), .ZN(n5215) );
  NAND2_X1 U6714 ( .A1(n5208), .A2(n7305), .ZN(n5209) );
  NAND2_X1 U6715 ( .A1(n5210), .A2(n5209), .ZN(n7307) );
  INV_X1 U6716 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5211) );
  OR2_X1 U6717 ( .A1(n5471), .A2(n5211), .ZN(n5212) );
  OAI21_X1 U6718 ( .B1(n5057), .B2(n7307), .A(n5212), .ZN(n5213) );
  INV_X1 U6719 ( .A(n5213), .ZN(n5214) );
  NOR2_X1 U6720 ( .A1(n6952), .A2(n5656), .ZN(n5216) );
  AOI21_X1 U6721 ( .B1(n6875), .B2(n5681), .A(n5216), .ZN(n7303) );
  NAND2_X1 U6722 ( .A1(n6875), .A2(n6193), .ZN(n5218) );
  NAND2_X1 U6723 ( .A1(n9137), .A2(n6197), .ZN(n5217) );
  NAND2_X1 U6724 ( .A1(n5218), .A2(n5217), .ZN(n5219) );
  XNOR2_X1 U6725 ( .A(n5219), .B(n5139), .ZN(n7301) );
  OAI22_X1 U6726 ( .A1(n7376), .A2(n7375), .B1(n7303), .B2(n7301), .ZN(n5224)
         );
  NAND3_X1 U6727 ( .A1(n7375), .A2(n7303), .A3(n7301), .ZN(n5223) );
  INV_X1 U6728 ( .A(n7301), .ZN(n7374) );
  INV_X1 U6729 ( .A(n7303), .ZN(n5220) );
  NOR2_X1 U6730 ( .A1(n7374), .A2(n5220), .ZN(n5221) );
  OAI21_X1 U6731 ( .B1(n5221), .B2(n7375), .A(n7376), .ZN(n5222) );
  MUX2_X1 U6732 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6389), .Z(n5227) );
  MUX2_X1 U6733 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6389), .Z(n5279) );
  XNOR2_X1 U6734 ( .A(n5279), .B(SI_11_), .ZN(n5228) );
  XNOR2_X1 U6735 ( .A(n5281), .B(n5228), .ZN(n6512) );
  NAND2_X1 U6736 ( .A1(n6512), .A2(n7781), .ZN(n5233) );
  NOR2_X1 U6737 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5229) );
  NAND2_X1 U6738 ( .A1(n5230), .A2(n5229), .ZN(n5249) );
  NAND2_X1 U6739 ( .A1(n5289), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5231) );
  XNOR2_X1 U6740 ( .A(n5231), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6514) );
  AOI22_X1 U6741 ( .A1(n5462), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5461), .B2(
        n6514), .ZN(n5232) );
  NAND2_X1 U6742 ( .A1(n7510), .A2(n6193), .ZN(n5244) );
  INV_X1 U6743 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7336) );
  INV_X1 U6744 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9631) );
  OR2_X1 U6745 ( .A1(n5452), .A2(n9631), .ZN(n5234) );
  OAI21_X1 U6746 ( .B1(n7655), .B2(n7336), .A(n5234), .ZN(n5235) );
  INV_X1 U6747 ( .A(n5235), .ZN(n5242) );
  INV_X1 U6748 ( .A(n5257), .ZN(n5236) );
  NAND2_X1 U6749 ( .A1(n5236), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6750 ( .A1(n5259), .A2(n5237), .ZN(n5238) );
  NAND2_X1 U6751 ( .A1(n5296), .A2(n5238), .ZN(n7514) );
  INV_X1 U6752 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9674) );
  OR2_X1 U6753 ( .A1(n5471), .A2(n9674), .ZN(n5239) );
  OAI21_X1 U6754 ( .B1(n5057), .B2(n7514), .A(n5239), .ZN(n5240) );
  INV_X1 U6755 ( .A(n5240), .ZN(n5241) );
  NAND2_X1 U6756 ( .A1(n9135), .A2(n5681), .ZN(n5243) );
  NAND2_X1 U6757 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  XNOR2_X1 U6758 ( .A(n5245), .B(n5628), .ZN(n7506) );
  NAND2_X1 U6759 ( .A1(n7510), .A2(n6197), .ZN(n5247) );
  NAND2_X1 U6760 ( .A1(n9135), .A2(n5630), .ZN(n5246) );
  NAND2_X1 U6761 ( .A1(n5247), .A2(n5246), .ZN(n7507) );
  NAND2_X1 U6762 ( .A1(n7506), .A2(n7507), .ZN(n7505) );
  INV_X1 U6763 ( .A(n7505), .ZN(n5270) );
  NAND2_X1 U6764 ( .A1(n6425), .A2(n7781), .ZN(n5252) );
  NAND2_X1 U6765 ( .A1(n5249), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5250) );
  XNOR2_X1 U6766 ( .A(n5250), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6500) );
  AOI22_X1 U6767 ( .A1(n5462), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5461), .B2(
        n6500), .ZN(n5251) );
  NAND2_X1 U6768 ( .A1(n7127), .A2(n6193), .ZN(n5266) );
  INV_X1 U6769 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7123) );
  INV_X1 U6770 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5253) );
  OR2_X1 U6771 ( .A1(n5452), .A2(n5253), .ZN(n5254) );
  OAI21_X1 U6772 ( .B1(n7655), .B2(n7123), .A(n5254), .ZN(n5255) );
  INV_X1 U6773 ( .A(n5255), .ZN(n5264) );
  INV_X1 U6774 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6775 ( .A1(n5257), .A2(n5256), .ZN(n5258) );
  NAND2_X1 U6776 ( .A1(n5259), .A2(n5258), .ZN(n7122) );
  INV_X1 U6777 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5260) );
  OR2_X1 U6778 ( .A1(n5471), .A2(n5260), .ZN(n5261) );
  OAI21_X1 U6779 ( .B1(n5057), .B2(n7122), .A(n5261), .ZN(n5262) );
  INV_X1 U6780 ( .A(n5262), .ZN(n5263) );
  INV_X1 U6781 ( .A(n7380), .ZN(n9136) );
  NAND2_X1 U6782 ( .A1(n9136), .A2(n6197), .ZN(n5265) );
  NAND2_X1 U6783 ( .A1(n5266), .A2(n5265), .ZN(n5267) );
  XNOR2_X1 U6784 ( .A(n5267), .B(n5139), .ZN(n7504) );
  NOR2_X1 U6785 ( .A1(n7380), .A2(n5656), .ZN(n5268) );
  AOI21_X1 U6786 ( .B1(n7127), .B2(n6197), .A(n5268), .ZN(n6374) );
  NOR2_X1 U6787 ( .A1(n7504), .A2(n6374), .ZN(n5269) );
  NAND2_X1 U6788 ( .A1(n6373), .A2(n5271), .ZN(n5278) );
  AND2_X1 U6789 ( .A1(n7504), .A2(n6374), .ZN(n5274) );
  INV_X1 U6790 ( .A(n7507), .ZN(n5273) );
  INV_X1 U6791 ( .A(n7506), .ZN(n5272) );
  OAI21_X1 U6792 ( .B1(n5274), .B2(n5273), .A(n5272), .ZN(n5276) );
  INV_X1 U6793 ( .A(n5274), .ZN(n5275) );
  AND2_X1 U6794 ( .A1(n5276), .A2(n4920), .ZN(n5277) );
  INV_X1 U6795 ( .A(n5279), .ZN(n5280) );
  INV_X1 U6796 ( .A(SI_11_), .ZN(n5282) );
  MUX2_X1 U6797 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6389), .Z(n5285) );
  NAND2_X1 U6798 ( .A1(n5285), .A2(SI_12_), .ZN(n5313) );
  OAI21_X1 U6799 ( .B1(n5285), .B2(SI_12_), .A(n5313), .ZN(n5286) );
  NAND2_X1 U6800 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  NAND2_X1 U6801 ( .A1(n5314), .A2(n5288), .ZN(n6520) );
  NOR2_X1 U6802 ( .A1(n5289), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5344) );
  OR2_X1 U6803 ( .A1(n5344), .A2(n5290), .ZN(n5320) );
  XNOR2_X1 U6804 ( .A(n5320), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7162) );
  AOI22_X1 U6805 ( .A1(n5462), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5461), .B2(
        n7162), .ZN(n5291) );
  NAND2_X1 U6806 ( .A1(n9622), .A2(n6193), .ZN(n5304) );
  INV_X1 U6807 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7222) );
  INV_X1 U6808 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6503) );
  OR2_X1 U6809 ( .A1(n5452), .A2(n6503), .ZN(n5292) );
  OAI21_X1 U6810 ( .B1(n7655), .B2(n7222), .A(n5292), .ZN(n5293) );
  INV_X1 U6811 ( .A(n5293), .ZN(n5302) );
  INV_X1 U6812 ( .A(n5296), .ZN(n5294) );
  NAND2_X1 U6813 ( .A1(n5294), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5327) );
  INV_X1 U6814 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6815 ( .A1(n5296), .A2(n5295), .ZN(n5297) );
  NAND2_X1 U6816 ( .A1(n5327), .A2(n5297), .ZN(n7408) );
  INV_X1 U6817 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5298) );
  OR2_X1 U6818 ( .A1(n5471), .A2(n5298), .ZN(n5299) );
  OAI21_X1 U6819 ( .B1(n5057), .B2(n7408), .A(n5299), .ZN(n5300) );
  INV_X1 U6820 ( .A(n5300), .ZN(n5301) );
  NAND2_X1 U6821 ( .A1(n9134), .A2(n6197), .ZN(n5303) );
  NAND2_X1 U6822 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  XNOR2_X1 U6823 ( .A(n5305), .B(n5139), .ZN(n5308) );
  INV_X1 U6824 ( .A(n5308), .ZN(n5310) );
  NOR2_X1 U6825 ( .A1(n7328), .A2(n5656), .ZN(n5306) );
  AOI21_X1 U6826 ( .B1(n9622), .B2(n5681), .A(n5306), .ZN(n5307) );
  INV_X1 U6827 ( .A(n5307), .ZN(n5309) );
  AND2_X1 U6828 ( .A1(n5308), .A2(n5307), .ZN(n5311) );
  AOI21_X1 U6829 ( .B1(n5310), .B2(n5309), .A(n5311), .ZN(n7406) );
  INV_X1 U6830 ( .A(n5311), .ZN(n5312) );
  MUX2_X1 U6831 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6389), .Z(n5315) );
  NAND2_X1 U6832 ( .A1(n5315), .A2(SI_13_), .ZN(n5339) );
  INV_X1 U6833 ( .A(n5315), .ZN(n5317) );
  INV_X1 U6834 ( .A(SI_13_), .ZN(n5316) );
  NAND2_X1 U6835 ( .A1(n5317), .A2(n5316), .ZN(n5318) );
  INV_X1 U6836 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6837 ( .A1(n5320), .A2(n5343), .ZN(n5321) );
  NAND2_X1 U6838 ( .A1(n5321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5322) );
  XNOR2_X1 U6839 ( .A(n5322), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9773) );
  AOI22_X1 U6840 ( .A1(n5462), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5461), .B2(
        n9773), .ZN(n5323) );
  OAI21_X2 U6841 ( .B1(n6529), .B2(n5083), .A(n5323), .ZN(n7486) );
  INV_X1 U6842 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7367) );
  INV_X1 U6843 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9618) );
  OR2_X1 U6844 ( .A1(n5452), .A2(n9618), .ZN(n5324) );
  OAI21_X1 U6845 ( .B1(n7655), .B2(n7367), .A(n5324), .ZN(n5325) );
  INV_X1 U6846 ( .A(n5325), .ZN(n5332) );
  NAND2_X1 U6847 ( .A1(n5327), .A2(n5326), .ZN(n5328) );
  NAND2_X1 U6848 ( .A1(n5351), .A2(n5328), .ZN(n7484) );
  INV_X1 U6849 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9669) );
  OR2_X1 U6850 ( .A1(n5471), .A2(n9669), .ZN(n5329) );
  OAI21_X1 U6851 ( .B1(n5057), .B2(n7484), .A(n5329), .ZN(n5330) );
  INV_X1 U6852 ( .A(n5330), .ZN(n5331) );
  AOI22_X1 U6853 ( .A1(n7486), .A2(n6197), .B1(n5630), .B2(n9133), .ZN(n5337)
         );
  NAND2_X1 U6854 ( .A1(n7486), .A2(n6193), .ZN(n5334) );
  NAND2_X1 U6855 ( .A1(n9133), .A2(n6197), .ZN(n5333) );
  NAND2_X1 U6856 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  XNOR2_X1 U6857 ( .A(n5335), .B(n5628), .ZN(n5336) );
  XOR2_X1 U6858 ( .A(n5337), .B(n5336), .Z(n7479) );
  INV_X1 U6859 ( .A(n5336), .ZN(n5338) );
  MUX2_X1 U6860 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6389), .Z(n5365) );
  XNOR2_X1 U6861 ( .A(n5365), .B(SI_14_), .ZN(n5341) );
  XNOR2_X1 U6862 ( .A(n5364), .B(n5341), .ZN(n6591) );
  NAND2_X1 U6863 ( .A1(n6591), .A2(n7781), .ZN(n5348) );
  INV_X1 U6864 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5342) );
  NAND3_X1 U6865 ( .A1(n5344), .A2(n5343), .A3(n5342), .ZN(n5345) );
  NAND2_X1 U6866 ( .A1(n5345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5346) );
  XNOR2_X1 U6867 ( .A(n5346), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9777) );
  AOI22_X1 U6868 ( .A1(n5462), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5461), .B2(
        n9777), .ZN(n5347) );
  NAND2_X1 U6869 ( .A1(n5349), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6870 ( .A1(n5351), .A2(n5350), .ZN(n5352) );
  AND2_X1 U6871 ( .A1(n5374), .A2(n5352), .ZN(n8981) );
  NAND2_X1 U6872 ( .A1(n5619), .A2(n8981), .ZN(n5356) );
  INV_X1 U6873 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5353) );
  OR2_X1 U6874 ( .A1(n5452), .A2(n5353), .ZN(n5355) );
  NAND2_X1 U6875 ( .A1(n5073), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5354) );
  NAND4_X1 U6876 ( .A1(n5357), .A2(n5356), .A3(n5355), .A4(n5354), .ZN(n9523)
         );
  AOI22_X1 U6877 ( .A1(n9611), .A2(n6193), .B1(n5681), .B2(n9523), .ZN(n5358)
         );
  XOR2_X1 U6878 ( .A(n5628), .B(n5358), .Z(n5359) );
  INV_X1 U6879 ( .A(n9611), .ZN(n8978) );
  INV_X1 U6880 ( .A(n9523), .ZN(n7481) );
  OAI22_X1 U6881 ( .A1(n8978), .A2(n5167), .B1(n7481), .B2(n5656), .ZN(n8975)
         );
  INV_X1 U6882 ( .A(n5365), .ZN(n5363) );
  NAND2_X1 U6883 ( .A1(n5365), .A2(SI_14_), .ZN(n5366) );
  MUX2_X1 U6884 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6389), .Z(n5386) );
  XNOR2_X1 U6885 ( .A(n5386), .B(SI_15_), .ZN(n5367) );
  XNOR2_X1 U6886 ( .A(n5389), .B(n5367), .ZN(n6827) );
  NAND2_X1 U6887 ( .A1(n6827), .A2(n7781), .ZN(n5371) );
  NAND2_X1 U6888 ( .A1(n5368), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5369) );
  XNOR2_X1 U6889 ( .A(n5369), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9804) );
  AOI22_X1 U6890 ( .A1(n5462), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5461), .B2(
        n9804), .ZN(n5370) );
  NAND2_X1 U6891 ( .A1(n5349), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5379) );
  INV_X1 U6892 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6893 ( .A1(n5374), .A2(n5373), .ZN(n5375) );
  AND2_X1 U6894 ( .A1(n5402), .A2(n5375), .ZN(n9512) );
  NAND2_X1 U6895 ( .A1(n5619), .A2(n9512), .ZN(n5378) );
  INV_X1 U6896 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9796) );
  OR2_X1 U6897 ( .A1(n5452), .A2(n9796), .ZN(n5377) );
  NAND2_X1 U6898 ( .A1(n5073), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5376) );
  NAND4_X1 U6899 ( .A1(n5379), .A2(n5378), .A3(n5377), .A4(n5376), .ZN(n9499)
         );
  AOI22_X1 U6900 ( .A1(n9606), .A2(n6193), .B1(n6197), .B2(n9499), .ZN(n5380)
         );
  XOR2_X1 U6901 ( .A(n5628), .B(n5380), .Z(n5381) );
  AOI22_X1 U6902 ( .A1(n9606), .A2(n5681), .B1(n5630), .B2(n9499), .ZN(n9114)
         );
  INV_X1 U6903 ( .A(n5384), .ZN(n5385) );
  INV_X1 U6904 ( .A(n5386), .ZN(n5387) );
  NAND2_X1 U6905 ( .A1(n5388), .A2(n5387), .ZN(n5392) );
  INV_X1 U6906 ( .A(n5389), .ZN(n5390) );
  NAND2_X1 U6907 ( .A1(n5390), .A2(n10155), .ZN(n5391) );
  MUX2_X1 U6908 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6389), .Z(n5415) );
  INV_X1 U6909 ( .A(SI_16_), .ZN(n10149) );
  XNOR2_X1 U6910 ( .A(n5415), .B(n10149), .ZN(n5393) );
  XNOR2_X1 U6911 ( .A(n5418), .B(n5393), .ZN(n6859) );
  NAND2_X1 U6912 ( .A1(n6859), .A2(n7781), .ZN(n5397) );
  NAND2_X1 U6913 ( .A1(n5394), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5395) );
  XNOR2_X1 U6914 ( .A(n5395), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7346) );
  AOI22_X1 U6915 ( .A1(n5462), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5461), .B2(
        n7346), .ZN(n5396) );
  NAND2_X1 U6916 ( .A1(n9601), .A2(n6193), .ZN(n5410) );
  INV_X1 U6917 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5399) );
  INV_X1 U6918 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7342) );
  OR2_X1 U6919 ( .A1(n5452), .A2(n7342), .ZN(n5398) );
  OAI21_X1 U6920 ( .B1(n7655), .B2(n5399), .A(n5398), .ZN(n5400) );
  INV_X1 U6921 ( .A(n5400), .ZN(n5408) );
  NAND2_X1 U6922 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  NAND2_X1 U6923 ( .A1(n5427), .A2(n5403), .ZN(n9492) );
  INV_X1 U6924 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5404) );
  OR2_X1 U6925 ( .A1(n5471), .A2(n5404), .ZN(n5405) );
  OAI21_X1 U6926 ( .B1(n5057), .B2(n9492), .A(n5405), .ZN(n5406) );
  INV_X1 U6927 ( .A(n5406), .ZN(n5407) );
  NAND2_X1 U6928 ( .A1(n9475), .A2(n6197), .ZN(n5409) );
  NAND2_X1 U6929 ( .A1(n5410), .A2(n5409), .ZN(n5411) );
  XNOR2_X1 U6930 ( .A(n5411), .B(n5139), .ZN(n5414) );
  NOR2_X1 U6931 ( .A1(n9517), .A2(n5656), .ZN(n5412) );
  AOI21_X1 U6932 ( .B1(n9601), .B2(n6197), .A(n5412), .ZN(n5413) );
  OR2_X1 U6933 ( .A1(n5414), .A2(n5413), .ZN(n9027) );
  NAND2_X1 U6934 ( .A1(n5414), .A2(n5413), .ZN(n9026) );
  NOR2_X1 U6935 ( .A1(n5415), .A2(SI_16_), .ZN(n5417) );
  NAND2_X1 U6936 ( .A1(n5415), .A2(SI_16_), .ZN(n5416) );
  MUX2_X1 U6937 ( .A(n7131), .B(n7133), .S(n6389), .Z(n5419) );
  NAND2_X1 U6938 ( .A1(n5419), .A2(n10041), .ZN(n5439) );
  INV_X1 U6939 ( .A(n5419), .ZN(n5420) );
  NAND2_X1 U6940 ( .A1(n5420), .A2(SI_17_), .ZN(n5421) );
  NAND2_X1 U6941 ( .A1(n5439), .A2(n5421), .ZN(n5440) );
  XNOR2_X1 U6942 ( .A(n5441), .B(n5440), .ZN(n7130) );
  NAND2_X1 U6943 ( .A1(n7130), .A2(n7781), .ZN(n5424) );
  XNOR2_X1 U6944 ( .A(n5422), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9259) );
  AOI22_X1 U6945 ( .A1(n5462), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5461), .B2(
        n9259), .ZN(n5423) );
  INV_X1 U6946 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6947 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  AND2_X1 U6948 ( .A1(n5465), .A2(n5428), .ZN(n9482) );
  NAND2_X1 U6949 ( .A1(n9482), .A2(n5619), .ZN(n5432) );
  INV_X1 U6950 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9598) );
  OR2_X1 U6951 ( .A1(n5452), .A2(n9598), .ZN(n5431) );
  NAND2_X1 U6952 ( .A1(n5349), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6953 ( .A1(n5073), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5429) );
  NAND4_X1 U6954 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), .ZN(n9501)
         );
  INV_X1 U6955 ( .A(n9501), .ZN(n9031) );
  OAI22_X1 U6956 ( .A1(n9664), .A2(n5167), .B1(n9031), .B2(n5656), .ZN(n5436)
         );
  NAND2_X1 U6957 ( .A1(n9481), .A2(n6193), .ZN(n5434) );
  NAND2_X1 U6958 ( .A1(n9501), .A2(n5681), .ZN(n5433) );
  NAND2_X1 U6959 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  XNOR2_X1 U6960 ( .A(n5435), .B(n5628), .ZN(n5437) );
  XOR2_X1 U6961 ( .A(n5436), .B(n5437), .Z(n9038) );
  OR2_X1 U6962 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  MUX2_X1 U6963 ( .A(n7218), .B(n5442), .S(n6389), .Z(n5443) );
  XNOR2_X1 U6964 ( .A(n5443), .B(SI_18_), .ZN(n5458) );
  INV_X1 U6965 ( .A(n5458), .ZN(n5445) );
  INV_X1 U6966 ( .A(n5443), .ZN(n5444) );
  MUX2_X1 U6967 ( .A(n7315), .B(n7313), .S(n6389), .Z(n5446) );
  INV_X1 U6968 ( .A(SI_19_), .ZN(n10073) );
  NAND2_X1 U6969 ( .A1(n5446), .A2(n10073), .ZN(n5486) );
  INV_X1 U6970 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U6971 ( .A1(n5447), .A2(SI_19_), .ZN(n5448) );
  NAND2_X1 U6972 ( .A1(n5486), .A2(n5448), .ZN(n5485) );
  XNOR2_X1 U6973 ( .A(n5484), .B(n5485), .ZN(n7312) );
  NAND2_X1 U6974 ( .A1(n7312), .A2(n7781), .ZN(n5450) );
  AOI22_X1 U6975 ( .A1(n5462), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9269), .B2(
        n5461), .ZN(n5449) );
  NAND2_X1 U6976 ( .A1(n9587), .A2(n6193), .ZN(n5456) );
  NAND2_X1 U6977 ( .A1(n5467), .A2(n9001), .ZN(n5451) );
  NAND2_X1 U6978 ( .A1(n5491), .A2(n5451), .ZN(n9448) );
  AOI22_X1 U6979 ( .A1(n5349), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n5073), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5454) );
  INV_X1 U6980 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9263) );
  OR2_X1 U6981 ( .A1(n5452), .A2(n9263), .ZN(n5453) );
  OAI211_X1 U6982 ( .C1(n9448), .C2(n5057), .A(n5454), .B(n5453), .ZN(n9132)
         );
  NAND2_X1 U6983 ( .A1(n9132), .A2(n5681), .ZN(n5455) );
  NAND2_X1 U6984 ( .A1(n5456), .A2(n5455), .ZN(n5457) );
  XNOR2_X1 U6985 ( .A(n5457), .B(n5628), .ZN(n8997) );
  AOI22_X1 U6986 ( .A1(n9587), .A2(n5681), .B1(n5630), .B2(n9132), .ZN(n8996)
         );
  INV_X1 U6987 ( .A(n8996), .ZN(n5477) );
  XNOR2_X1 U6988 ( .A(n5459), .B(n5458), .ZN(n7154) );
  NAND2_X1 U6989 ( .A1(n7154), .A2(n7781), .ZN(n5464) );
  XNOR2_X1 U6990 ( .A(n5460), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9812) );
  AOI22_X1 U6991 ( .A1(n5462), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5461), .B2(
        n9812), .ZN(n5463) );
  NAND2_X1 U6992 ( .A1(n9592), .A2(n5681), .ZN(n5473) );
  INV_X1 U6993 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6994 ( .A1(n5465), .A2(n9092), .ZN(n5466) );
  NAND2_X1 U6995 ( .A1(n5467), .A2(n5466), .ZN(n9462) );
  OR2_X1 U6996 ( .A1(n9462), .A2(n5057), .ZN(n5469) );
  AOI22_X1 U6997 ( .A1(n5349), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n7651), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5468) );
  OAI211_X1 U6998 ( .C1(n5471), .C2(n5470), .A(n5469), .B(n5468), .ZN(n9474)
         );
  NAND2_X1 U6999 ( .A1(n9474), .A2(n5630), .ZN(n5472) );
  NAND2_X1 U7000 ( .A1(n9592), .A2(n6193), .ZN(n5475) );
  NAND2_X1 U7001 ( .A1(n9474), .A2(n6197), .ZN(n5474) );
  NAND2_X1 U7002 ( .A1(n5475), .A2(n5474), .ZN(n5476) );
  XNOR2_X1 U7003 ( .A(n5476), .B(n5139), .ZN(n8995) );
  INV_X1 U7004 ( .A(n8995), .ZN(n5480) );
  AOI22_X1 U7005 ( .A1(n8997), .A2(n5477), .B1(n9089), .B2(n5480), .ZN(n5483)
         );
  AOI21_X1 U7006 ( .B1(n8995), .B2(n5478), .A(n8996), .ZN(n5481) );
  NAND2_X1 U7007 ( .A1(n8996), .A2(n5478), .ZN(n5479) );
  OAI22_X1 U7008 ( .A1(n5481), .A2(n8997), .B1(n5480), .B2(n5479), .ZN(n5482)
         );
  MUX2_X1 U7009 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6389), .Z(n5505) );
  XNOR2_X1 U7010 ( .A(n5505), .B(n10170), .ZN(n5487) );
  XNOR2_X1 U7011 ( .A(n5507), .B(n5487), .ZN(n7401) );
  NAND2_X1 U7012 ( .A1(n7401), .A2(n7781), .ZN(n5489) );
  INV_X1 U7013 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7400) );
  OR2_X1 U7014 ( .A1(n7782), .A2(n7400), .ZN(n5488) );
  NAND2_X1 U7015 ( .A1(n9582), .A2(n6193), .ZN(n5500) );
  INV_X1 U7016 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U7017 ( .A1(n5491), .A2(n9073), .ZN(n5492) );
  AND2_X1 U7018 ( .A1(n5514), .A2(n5492), .ZN(n9436) );
  NAND2_X1 U7019 ( .A1(n9436), .A2(n5619), .ZN(n5498) );
  INV_X1 U7020 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7021 ( .A1(n7651), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U7022 ( .A1(n5073), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5493) );
  OAI211_X1 U7023 ( .C1(n7655), .C2(n5495), .A(n5494), .B(n5493), .ZN(n5496)
         );
  INV_X1 U7024 ( .A(n5496), .ZN(n5497) );
  NAND2_X1 U7025 ( .A1(n5498), .A2(n5497), .ZN(n9131) );
  NAND2_X1 U7026 ( .A1(n9131), .A2(n6197), .ZN(n5499) );
  NAND2_X1 U7027 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  XNOR2_X1 U7028 ( .A(n5501), .B(n5139), .ZN(n9070) );
  AND2_X1 U7029 ( .A1(n9131), .A2(n5630), .ZN(n5502) );
  AOI21_X1 U7030 ( .B1(n9582), .B2(n5681), .A(n5502), .ZN(n5503) );
  INV_X1 U7031 ( .A(n9070), .ZN(n5504) );
  INV_X1 U7032 ( .A(n5503), .ZN(n9069) );
  INV_X1 U7033 ( .A(n5505), .ZN(n5506) );
  NAND2_X1 U7034 ( .A1(n5507), .A2(n10170), .ZN(n5508) );
  NAND2_X1 U7035 ( .A1(n5509), .A2(n5508), .ZN(n5535) );
  MUX2_X1 U7036 ( .A(n7490), .B(n7500), .S(n6389), .Z(n5531) );
  XNOR2_X1 U7037 ( .A(n5531), .B(SI_21_), .ZN(n5510) );
  XNOR2_X1 U7038 ( .A(n5535), .B(n5510), .ZN(n7489) );
  NAND2_X1 U7039 ( .A1(n7489), .A2(n7781), .ZN(n5512) );
  OR2_X1 U7040 ( .A1(n7782), .A2(n7500), .ZN(n5511) );
  NAND2_X1 U7041 ( .A1(n9422), .A2(n6193), .ZN(n5523) );
  INV_X1 U7042 ( .A(n5514), .ZN(n5513) );
  INV_X1 U7043 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9012) );
  NAND2_X1 U7044 ( .A1(n5514), .A2(n9012), .ZN(n5515) );
  NAND2_X1 U7045 ( .A1(n5542), .A2(n5515), .ZN(n9010) );
  OR2_X1 U7046 ( .A1(n9010), .A2(n5057), .ZN(n5521) );
  INV_X1 U7047 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7048 ( .A1(n7651), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7049 ( .A1(n5073), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5516) );
  OAI211_X1 U7050 ( .C1(n7655), .C2(n5518), .A(n5517), .B(n5516), .ZN(n5519)
         );
  INV_X1 U7051 ( .A(n5519), .ZN(n5520) );
  NAND2_X1 U7052 ( .A1(n5521), .A2(n5520), .ZN(n9407) );
  NAND2_X1 U7053 ( .A1(n9407), .A2(n6197), .ZN(n5522) );
  NAND2_X1 U7054 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  XNOR2_X1 U7055 ( .A(n5524), .B(n5628), .ZN(n5528) );
  NAND2_X1 U7056 ( .A1(n9422), .A2(n5681), .ZN(n5526) );
  NAND2_X1 U7057 ( .A1(n9407), .A2(n5630), .ZN(n5525) );
  NAND2_X1 U7058 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  NOR2_X1 U7059 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  AOI21_X1 U7060 ( .B1(n5528), .B2(n5527), .A(n5529), .ZN(n9008) );
  INV_X1 U7061 ( .A(n5529), .ZN(n5530) );
  NOR2_X1 U7062 ( .A1(n5532), .A2(SI_21_), .ZN(n5534) );
  NAND2_X1 U7063 ( .A1(n5532), .A2(SI_21_), .ZN(n5533) );
  MUX2_X1 U7064 ( .A(n7553), .B(n7555), .S(n6389), .Z(n5536) );
  INV_X1 U7065 ( .A(SI_22_), .ZN(n10035) );
  NAND2_X1 U7066 ( .A1(n5536), .A2(n10035), .ZN(n5554) );
  INV_X1 U7067 ( .A(n5536), .ZN(n5537) );
  NAND2_X1 U7068 ( .A1(n5537), .A2(SI_22_), .ZN(n5538) );
  NAND2_X1 U7069 ( .A1(n5554), .A2(n5538), .ZN(n5555) );
  XNOR2_X1 U7070 ( .A(n5556), .B(n5555), .ZN(n7551) );
  NAND2_X1 U7071 ( .A1(n7551), .A2(n7781), .ZN(n5540) );
  OR2_X1 U7072 ( .A1(n7782), .A2(n7555), .ZN(n5539) );
  NAND2_X1 U7073 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  AND2_X1 U7074 ( .A1(n5564), .A2(n5543), .ZN(n9401) );
  NAND2_X1 U7075 ( .A1(n9401), .A2(n5619), .ZN(n5549) );
  INV_X1 U7076 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7077 ( .A1(n7651), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7078 ( .A1(n5073), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5544) );
  OAI211_X1 U7079 ( .C1(n7655), .C2(n5546), .A(n5545), .B(n5544), .ZN(n5547)
         );
  INV_X1 U7080 ( .A(n5547), .ZN(n5548) );
  NAND2_X1 U7081 ( .A1(n5549), .A2(n5548), .ZN(n9130) );
  AOI22_X1 U7082 ( .A1(n9571), .A2(n6193), .B1(n6197), .B2(n9130), .ZN(n5550)
         );
  XNOR2_X1 U7083 ( .A(n5550), .B(n5628), .ZN(n5551) );
  INV_X1 U7084 ( .A(n9571), .ZN(n9403) );
  INV_X1 U7085 ( .A(n9130), .ZN(n9381) );
  OAI22_X1 U7086 ( .A1(n9403), .A2(n5167), .B1(n9381), .B2(n5656), .ZN(n9080)
         );
  INV_X1 U7087 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7588) );
  INV_X1 U7088 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7584) );
  MUX2_X1 U7089 ( .A(n7588), .B(n7584), .S(n6389), .Z(n5558) );
  NAND2_X1 U7090 ( .A1(n5558), .A2(n5557), .ZN(n5605) );
  INV_X1 U7091 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U7092 ( .A1(n5559), .A2(SI_23_), .ZN(n5560) );
  XNOR2_X1 U7093 ( .A(n5582), .B(n5581), .ZN(n7585) );
  NAND2_X1 U7094 ( .A1(n7585), .A2(n7781), .ZN(n5562) );
  OR2_X1 U7095 ( .A1(n7782), .A2(n7584), .ZN(n5561) );
  NAND2_X1 U7096 ( .A1(n9388), .A2(n6193), .ZN(n5572) );
  INV_X1 U7097 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U7098 ( .A1(n5564), .A2(n8989), .ZN(n5565) );
  NAND2_X1 U7099 ( .A1(n5617), .A2(n5565), .ZN(n9391) );
  OR2_X1 U7100 ( .A1(n9391), .A2(n5057), .ZN(n5570) );
  INV_X1 U7101 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U7102 ( .A1(n5073), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7103 ( .A1(n7651), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5566) );
  OAI211_X1 U7104 ( .C1(n7655), .C2(n9389), .A(n5567), .B(n5566), .ZN(n5568)
         );
  INV_X1 U7105 ( .A(n5568), .ZN(n5569) );
  NAND2_X1 U7106 ( .A1(n9408), .A2(n5681), .ZN(n5571) );
  NAND2_X1 U7107 ( .A1(n5572), .A2(n5571), .ZN(n5573) );
  XNOR2_X1 U7108 ( .A(n5573), .B(n5139), .ZN(n5575) );
  AND2_X1 U7109 ( .A1(n9408), .A2(n5630), .ZN(n5574) );
  AOI21_X1 U7110 ( .B1(n9388), .B2(n5681), .A(n5574), .ZN(n5576) );
  NAND2_X1 U7111 ( .A1(n5575), .A2(n5576), .ZN(n5580) );
  INV_X1 U7112 ( .A(n5575), .ZN(n5578) );
  INV_X1 U7113 ( .A(n5576), .ZN(n5577) );
  NAND2_X1 U7114 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  NAND2_X1 U7115 ( .A1(n5580), .A2(n5579), .ZN(n8986) );
  INV_X1 U7116 ( .A(n5580), .ZN(n9048) );
  NAND2_X1 U7117 ( .A1(n5607), .A2(n5605), .ZN(n5587) );
  INV_X1 U7118 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7624) );
  INV_X1 U7119 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7590) );
  MUX2_X1 U7120 ( .A(n7624), .B(n7590), .S(n6389), .Z(n5584) );
  INV_X1 U7121 ( .A(SI_24_), .ZN(n5583) );
  NAND2_X1 U7122 ( .A1(n5584), .A2(n5583), .ZN(n5604) );
  INV_X1 U7123 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7124 ( .A1(n5585), .A2(SI_24_), .ZN(n5632) );
  AND2_X1 U7125 ( .A1(n5604), .A2(n5632), .ZN(n5586) );
  NAND2_X1 U7126 ( .A1(n7589), .A2(n7781), .ZN(n5589) );
  OR2_X1 U7127 ( .A1(n7782), .A2(n7590), .ZN(n5588) );
  NAND2_X1 U7128 ( .A1(n9560), .A2(n6193), .ZN(n5597) );
  XNOR2_X1 U7129 ( .A(n5617), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U7130 ( .A1(n9371), .A2(n5017), .ZN(n5595) );
  INV_X1 U7131 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7132 ( .A1(n5073), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7133 ( .A1(n7651), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5590) );
  OAI211_X1 U7134 ( .C1(n7655), .C2(n5592), .A(n5591), .B(n5590), .ZN(n5593)
         );
  INV_X1 U7135 ( .A(n5593), .ZN(n5594) );
  OR2_X1 U7136 ( .A1(n9382), .A2(n5167), .ZN(n5596) );
  NAND2_X1 U7137 ( .A1(n5597), .A2(n5596), .ZN(n5598) );
  XNOR2_X1 U7138 ( .A(n5598), .B(n5139), .ZN(n5601) );
  NOR2_X1 U7139 ( .A1(n9382), .A2(n5656), .ZN(n5599) );
  AOI21_X1 U7140 ( .B1(n9560), .B2(n5681), .A(n5599), .ZN(n5600) );
  NAND2_X1 U7141 ( .A1(n5601), .A2(n5600), .ZN(n5603) );
  OR2_X1 U7142 ( .A1(n5601), .A2(n5600), .ZN(n5602) );
  AND2_X1 U7143 ( .A1(n5603), .A2(n5602), .ZN(n9047) );
  AND2_X1 U7144 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  AND2_X1 U7145 ( .A1(n5635), .A2(n5632), .ZN(n5612) );
  INV_X1 U7146 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7635) );
  INV_X1 U7147 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7627) );
  MUX2_X1 U7148 ( .A(n7635), .B(n7627), .S(n6389), .Z(n5609) );
  INV_X1 U7149 ( .A(SI_25_), .ZN(n5608) );
  NAND2_X1 U7150 ( .A1(n5609), .A2(n5608), .ZN(n5636) );
  INV_X1 U7151 ( .A(n5609), .ZN(n5610) );
  NAND2_X1 U7152 ( .A1(n5610), .A2(SI_25_), .ZN(n5611) );
  NAND2_X1 U7153 ( .A1(n7626), .A2(n7781), .ZN(n5614) );
  OR2_X1 U7154 ( .A1(n7782), .A2(n7627), .ZN(n5613) );
  NAND2_X1 U7155 ( .A1(n9355), .A2(n6193), .ZN(n5627) );
  INV_X1 U7156 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9051) );
  INV_X1 U7157 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5615) );
  OAI21_X1 U7158 ( .B1(n5617), .B2(n9051), .A(n5615), .ZN(n5618) );
  NAND2_X1 U7159 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5616) );
  NAND2_X1 U7160 ( .A1(n9356), .A2(n5619), .ZN(n5625) );
  INV_X1 U7161 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7162 ( .A1(n7651), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7163 ( .A1(n5073), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5620) );
  OAI211_X1 U7164 ( .C1(n7655), .C2(n5622), .A(n5621), .B(n5620), .ZN(n5623)
         );
  INV_X1 U7165 ( .A(n5623), .ZN(n5624) );
  NAND2_X1 U7166 ( .A1(n9339), .A2(n6197), .ZN(n5626) );
  NAND2_X1 U7167 ( .A1(n5627), .A2(n5626), .ZN(n5629) );
  XNOR2_X1 U7168 ( .A(n5629), .B(n5628), .ZN(n5660) );
  AOI22_X1 U7169 ( .A1(n9355), .A2(n5681), .B1(n5630), .B2(n9339), .ZN(n5658)
         );
  NAND2_X1 U7170 ( .A1(n5637), .A2(n5636), .ZN(n5663) );
  INV_X1 U7171 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7630) );
  INV_X1 U7172 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7632) );
  MUX2_X1 U7173 ( .A(n7630), .B(n7632), .S(n6389), .Z(n5638) );
  NAND2_X1 U7174 ( .A1(n5638), .A2(n10164), .ZN(n5664) );
  INV_X1 U7175 ( .A(n5638), .ZN(n5639) );
  NAND2_X1 U7176 ( .A1(n5639), .A2(SI_26_), .ZN(n5640) );
  XNOR2_X1 U7177 ( .A(n5663), .B(n5662), .ZN(n7629) );
  NAND2_X1 U7178 ( .A1(n7629), .A2(n7781), .ZN(n5642) );
  OR2_X1 U7179 ( .A1(n7782), .A2(n7632), .ZN(n5641) );
  NAND2_X1 U7180 ( .A1(n9549), .A2(n6193), .ZN(n5654) );
  INV_X1 U7181 ( .A(n5645), .ZN(n5643) );
  INV_X1 U7182 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7183 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  NAND2_X1 U7184 ( .A1(n5730), .A2(n5646), .ZN(n9332) );
  INV_X1 U7185 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7186 ( .A1(n5073), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7187 ( .A1(n7651), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5647) );
  OAI211_X1 U7188 ( .C1(n7655), .C2(n5649), .A(n5648), .B(n5647), .ZN(n5650)
         );
  INV_X1 U7189 ( .A(n5650), .ZN(n5651) );
  NAND2_X1 U7190 ( .A1(n9128), .A2(n5681), .ZN(n5653) );
  NAND2_X1 U7191 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  XNOR2_X1 U7192 ( .A(n5655), .B(n5139), .ZN(n5687) );
  NOR2_X1 U7193 ( .A1(n9350), .A2(n5656), .ZN(n5657) );
  AOI21_X1 U7194 ( .B1(n9549), .B2(n5681), .A(n5657), .ZN(n5686) );
  XNOR2_X1 U7195 ( .A(n5687), .B(n5686), .ZN(n9101) );
  INV_X1 U7196 ( .A(n5658), .ZN(n5659) );
  NOR2_X1 U7197 ( .A1(n5660), .A2(n5659), .ZN(n9102) );
  NOR2_X1 U7198 ( .A1(n9101), .A2(n9102), .ZN(n5661) );
  NAND2_X2 U7199 ( .A1(n9100), .A2(n5661), .ZN(n9104) );
  NAND2_X1 U7200 ( .A1(n5663), .A2(n5662), .ZN(n5665) );
  INV_X1 U7201 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9693) );
  MUX2_X1 U7202 ( .A(n8972), .B(n9693), .S(n6389), .Z(n5666) );
  INV_X1 U7203 ( .A(SI_27_), .ZN(n10167) );
  NAND2_X1 U7204 ( .A1(n5666), .A2(n10167), .ZN(n6105) );
  INV_X1 U7205 ( .A(n5666), .ZN(n5667) );
  NAND2_X1 U7206 ( .A1(n5667), .A2(SI_27_), .ZN(n5668) );
  NAND2_X1 U7207 ( .A1(n9690), .A2(n7781), .ZN(n5670) );
  OR2_X1 U7208 ( .A1(n7782), .A2(n9693), .ZN(n5669) );
  NAND2_X1 U7209 ( .A1(n9322), .A2(n6193), .ZN(n5678) );
  XNOR2_X1 U7210 ( .A(n5730), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U7211 ( .A1(n9323), .A2(n5619), .ZN(n5676) );
  INV_X1 U7212 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7213 ( .A1(n5073), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U7214 ( .A1(n7651), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5671) );
  OAI211_X1 U7215 ( .C1(n7655), .C2(n5673), .A(n5672), .B(n5671), .ZN(n5674)
         );
  INV_X1 U7216 ( .A(n5674), .ZN(n5675) );
  OR2_X1 U7217 ( .A1(n9304), .A2(n5167), .ZN(n5677) );
  NAND2_X1 U7218 ( .A1(n5678), .A2(n5677), .ZN(n5679) );
  XNOR2_X1 U7219 ( .A(n5679), .B(n5139), .ZN(n5683) );
  INV_X1 U7220 ( .A(n5683), .ZN(n5685) );
  NOR2_X1 U7221 ( .A1(n9304), .A2(n5656), .ZN(n5680) );
  AOI21_X1 U7222 ( .B1(n9322), .B2(n6197), .A(n5680), .ZN(n5682) );
  INV_X1 U7223 ( .A(n5682), .ZN(n5684) );
  AOI21_X1 U7224 ( .B1(n5685), .B2(n5684), .A(n6204), .ZN(n5691) );
  INV_X1 U7225 ( .A(n5691), .ZN(n5689) );
  OR2_X1 U7226 ( .A1(n5687), .A2(n5686), .ZN(n5692) );
  INV_X1 U7227 ( .A(n5692), .ZN(n5688) );
  NOR2_X1 U7228 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  NAND2_X1 U7229 ( .A1(n7628), .A2(P1_B_REG_SCAN_IN), .ZN(n5694) );
  MUX2_X1 U7230 ( .A(n5694), .B(P1_B_REG_SCAN_IN), .S(n5693), .Z(n5695) );
  INV_X1 U7231 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U7232 ( .A1(n6416), .A2(n5696), .ZN(n5698) );
  INV_X1 U7233 ( .A(n5697), .ZN(n7634) );
  NAND2_X1 U7234 ( .A1(n7634), .A2(n7628), .ZN(n9678) );
  NAND2_X1 U7235 ( .A1(n5698), .A2(n9678), .ZN(n6357) );
  INV_X1 U7236 ( .A(n6357), .ZN(n6611) );
  INV_X1 U7237 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5699) );
  INV_X1 U7238 ( .A(n5693), .ZN(n7591) );
  NOR4_X1 U7239 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5708) );
  NOR4_X1 U7240 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5707) );
  NOR4_X1 U7241 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5703) );
  NOR4_X1 U7242 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5702) );
  NOR4_X1 U7243 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5701) );
  NOR4_X1 U7244 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5700) );
  NAND4_X1 U7245 ( .A1(n5703), .A2(n5702), .A3(n5701), .A4(n5700), .ZN(n5704)
         );
  NOR4_X1 U7246 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5705), .A4(n5704), .ZN(n5706) );
  NAND3_X1 U7247 ( .A1(n5708), .A2(n5707), .A3(n5706), .ZN(n5709) );
  NAND2_X1 U7248 ( .A1(n6416), .A2(n5709), .ZN(n6360) );
  NAND3_X1 U7249 ( .A1(n6611), .A2(n6367), .A3(n6360), .ZN(n5720) );
  INV_X1 U7250 ( .A(n5713), .ZN(n7929) );
  INV_X1 U7251 ( .A(n7861), .ZN(n6407) );
  NOR2_X1 U7252 ( .A1(n9623), .A2(n6407), .ZN(n5714) );
  INV_X1 U7253 ( .A(n5725), .ZN(n5716) );
  NAND2_X1 U7254 ( .A1(n6325), .A2(n7870), .ZN(n6619) );
  NAND2_X1 U7255 ( .A1(n9531), .A2(n9269), .ZN(n6356) );
  OR2_X1 U7256 ( .A1(n5718), .A2(P1_U3086), .ZN(n7398) );
  NAND2_X1 U7257 ( .A1(n9623), .A2(n7398), .ZN(n5719) );
  NAND2_X1 U7258 ( .A1(n5720), .A2(n5719), .ZN(n5722) );
  NOR2_X1 U7259 ( .A1(n7861), .A2(n5713), .ZN(n6358) );
  INV_X1 U7260 ( .A(n6358), .ZN(n5721) );
  NAND2_X1 U7261 ( .A1(n5722), .A2(n5721), .ZN(n6526) );
  OAI21_X1 U7262 ( .B1(n6526), .B2(n5723), .A(P1_STATE_REG_SCAN_IN), .ZN(n5724) );
  NOR2_X2 U7263 ( .A1(n7861), .A2(n4352), .ZN(n9524) );
  NAND2_X1 U7264 ( .A1(n9060), .A2(n9524), .ZN(n9083) );
  INV_X1 U7265 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5728) );
  OAI22_X1 U7266 ( .A1(n9350), .A2(n9083), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5728), .ZN(n5738) );
  INV_X1 U7267 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5727) );
  OAI21_X1 U7268 ( .B1(n5730), .B2(n5728), .A(n5727), .ZN(n5731) );
  NAND2_X1 U7269 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5729) );
  NAND2_X1 U7270 ( .A1(n9293), .A2(n5619), .ZN(n5736) );
  INV_X1 U7271 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U7272 ( .A1(n5073), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7273 ( .A1(n7651), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5732) );
  OAI211_X1 U7274 ( .C1(n7655), .C2(n9294), .A(n5733), .B(n5732), .ZN(n5734)
         );
  INV_X1 U7275 ( .A(n5734), .ZN(n5735) );
  NAND2_X1 U7276 ( .A1(n9060), .A2(n9500), .ZN(n9119) );
  NOR2_X1 U7277 ( .A1(n9315), .A2(n9119), .ZN(n5737) );
  AOI211_X1 U7278 ( .C1(n9323), .C2(n9121), .A(n5738), .B(n5737), .ZN(n5739)
         );
  INV_X1 U7279 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7280 ( .A1(n5742), .A2(n5741), .ZN(P1_U3214) );
  NOR2_X1 U7281 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5754) );
  NOR2_X1 U7282 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5753) );
  NOR2_X1 U7283 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5752) );
  NOR2_X1 U7284 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5751) );
  INV_X1 U7285 ( .A(n5782), .ZN(n5762) );
  NAND2_X2 U7286 ( .A1(n5832), .A2(n6388), .ZN(n5827) );
  NAND2_X1 U7287 ( .A1(n7585), .A2(n8224), .ZN(n5765) );
  OR2_X1 U7288 ( .A1(n8222), .A2(n7588), .ZN(n5764) );
  NAND2_X1 U7289 ( .A1(n10165), .A2(n10141), .ZN(n5862) );
  INV_X1 U7290 ( .A(n5862), .ZN(n5767) );
  INV_X1 U7291 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7292 ( .A1(n5767), .A2(n5766), .ZN(n5874) );
  INV_X1 U7293 ( .A(n5886), .ZN(n5768) );
  NAND2_X1 U7294 ( .A1(n5768), .A2(n10130), .ZN(n5899) );
  INV_X1 U7295 ( .A(n5909), .ZN(n5770) );
  INV_X1 U7296 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7297 ( .A1(n5770), .A2(n5769), .ZN(n5927) );
  INV_X1 U7298 ( .A(n5956), .ZN(n5771) );
  NAND2_X1 U7299 ( .A1(n5771), .A2(n7438), .ZN(n5958) );
  INV_X1 U7300 ( .A(n5958), .ZN(n5772) );
  NAND2_X1 U7301 ( .A1(n5772), .A2(n10125), .ZN(n5975) );
  INV_X1 U7302 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U7303 ( .A1(n5774), .A2(n5773), .ZN(n6007) );
  INV_X1 U7304 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U7305 ( .A1(n10038), .A2(n10059), .ZN(n5777) );
  INV_X1 U7306 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7307 ( .A1(n6058), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7308 ( .A1(n6064), .A2(n5780), .ZN(n8711) );
  NAND2_X1 U7309 ( .A1(n8711), .A2(n5822), .ZN(n5790) );
  AOI22_X1 U7310 ( .A1(n5840), .A2(P2_REG0_REG_23__SCAN_IN), .B1(n5839), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n5789) );
  INV_X2 U7311 ( .A(n5812), .ZN(n5838) );
  NAND2_X1 U7312 ( .A1(n5838), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7313 ( .A1(n5840), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5797) );
  INV_X1 U7314 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8756) );
  OR2_X1 U7315 ( .A1(n6029), .A2(n8756), .ZN(n5796) );
  NAND2_X1 U7316 ( .A1(n6032), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5793) );
  AND2_X1 U7317 ( .A1(n6046), .A2(n5793), .ZN(n8757) );
  OR2_X1 U7318 ( .A1(n6124), .A2(n8757), .ZN(n5795) );
  INV_X1 U7319 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8867) );
  OR2_X1 U7320 ( .A1(n6127), .A2(n8867), .ZN(n5794) );
  NAND2_X1 U7321 ( .A1(n7312), .A2(n8224), .ZN(n5802) );
  NAND2_X1 U7322 ( .A1(n4396), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5800) );
  AOI22_X1 U7323 ( .A1(n6026), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8443), .B2(
        n6385), .ZN(n5801) );
  INV_X1 U7324 ( .A(n8932), .ZN(n8073) );
  NAND2_X1 U7325 ( .A1(n5838), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7326 ( .A1(n5840), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5803) );
  NAND4_X2 U7327 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .ZN(n5819)
         );
  INV_X1 U7328 ( .A(n5819), .ZN(n5811) );
  INV_X1 U7329 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5807) );
  INV_X1 U7330 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6387) );
  INV_X1 U7331 ( .A(n6397), .ZN(n5808) );
  OR2_X1 U7332 ( .A1(n6385), .A2(n4407), .ZN(n5809) );
  OAI211_X2 U7333 ( .C1(n5832), .C2(n6732), .A(n5810), .B(n5809), .ZN(n5820)
         );
  NAND2_X2 U7334 ( .A1(n6175), .A2(n8273), .ZN(n8244) );
  INV_X1 U7335 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10044) );
  INV_X1 U7336 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6662) );
  OR2_X1 U7337 ( .A1(n5812), .A2(n6662), .ZN(n5814) );
  NAND2_X1 U7338 ( .A1(n5840), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7339 ( .A1(n5817), .A2(SI_0_), .ZN(n5818) );
  XNOR2_X1 U7340 ( .A(n5818), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8973) );
  MUX2_X1 U7341 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8973), .S(n5832), .Z(n7021) );
  NAND2_X1 U7342 ( .A1(n8466), .A2(n7021), .ZN(n6970) );
  NAND2_X1 U7343 ( .A1(n8244), .A2(n6970), .ZN(n7138) );
  NAND2_X1 U7344 ( .A1(n5840), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7345 ( .A1(n5839), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7346 ( .A1(n5822), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7347 ( .A1(n5838), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5823) );
  OR2_X1 U7348 ( .A1(n5827), .A2(n6394), .ZN(n5834) );
  INV_X1 U7349 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5828) );
  INV_X1 U7350 ( .A(n5836), .ZN(n5837) );
  OR2_X1 U7351 ( .A1(n6843), .A2(n9891), .ZN(n8279) );
  NAND2_X1 U7352 ( .A1(n6843), .A2(n9891), .ZN(n8281) );
  NAND2_X1 U7353 ( .A1(n5838), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7354 ( .A1(n5839), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7355 ( .A1(n5840), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5841) );
  OR2_X1 U7356 ( .A1(n6124), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7357 ( .A1(n5845), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5847) );
  INV_X1 U7358 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5846) );
  XNOR2_X1 U7359 ( .A(n5847), .B(n5846), .ZN(n6691) );
  OR2_X1 U7360 ( .A1(n8222), .A2(n5006), .ZN(n5849) );
  INV_X1 U7361 ( .A(n7068), .ZN(n7150) );
  NAND2_X1 U7362 ( .A1(n8465), .A2(n7150), .ZN(n8289) );
  NAND3_X1 U7363 ( .A1(n6845), .A2(n6844), .A3(n8245), .ZN(n5851) );
  NAND2_X1 U7364 ( .A1(n7211), .A2(n7150), .ZN(n5850) );
  NAND2_X1 U7365 ( .A1(n5851), .A2(n5850), .ZN(n7054) );
  NAND2_X1 U7366 ( .A1(n5840), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7367 ( .A1(n5839), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U7368 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5852) );
  AND2_X1 U7369 ( .A1(n5862), .A2(n5852), .ZN(n7216) );
  OR2_X1 U7370 ( .A1(n6124), .A2(n7216), .ZN(n5854) );
  NAND2_X1 U7371 ( .A1(n5838), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U7372 ( .A1(n4394), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5857) );
  XNOR2_X1 U7373 ( .A(n5857), .B(n5743), .ZN(n6695) );
  INV_X1 U7374 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6393) );
  OR2_X1 U7375 ( .A1(n8222), .A2(n6393), .ZN(n5858) );
  OAI211_X1 U7376 ( .C1(n5832), .C2(n6695), .A(n5859), .B(n5858), .ZN(n8306)
         );
  NOR2_X1 U7377 ( .A1(n8464), .A2(n8306), .ZN(n5861) );
  NAND2_X1 U7378 ( .A1(n8464), .A2(n8306), .ZN(n5860) );
  OAI21_X2 U7379 ( .B1(n7054), .B2(n5861), .A(n5860), .ZN(n7281) );
  NAND2_X1 U7380 ( .A1(n5840), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7381 ( .A1(n5839), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7382 ( .A1(n5862), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5863) );
  AND2_X1 U7383 ( .A1(n5874), .A2(n5863), .ZN(n7279) );
  OR2_X1 U7384 ( .A1(n6124), .A2(n7279), .ZN(n5866) );
  INV_X1 U7385 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5864) );
  OR2_X1 U7386 ( .A1(n6127), .A2(n5864), .ZN(n5865) );
  NAND4_X1 U7387 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(n8463)
         );
  OR2_X1 U7388 ( .A1(n5869), .A2(n4837), .ZN(n5870) );
  XNOR2_X1 U7389 ( .A(n5870), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6807) );
  INV_X1 U7390 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6396) );
  OR2_X1 U7391 ( .A1(n8222), .A2(n6396), .ZN(n5871) );
  OAI211_X1 U7392 ( .C1(n5832), .C2(n6812), .A(n5872), .B(n5871), .ZN(n7239)
         );
  AND2_X1 U7393 ( .A1(n8463), .A2(n7239), .ZN(n5873) );
  NAND2_X1 U7394 ( .A1(n5839), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U7395 ( .A1(n5838), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7396 ( .A1(n5874), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5875) );
  AND2_X1 U7397 ( .A1(n5886), .A2(n5875), .ZN(n7317) );
  OR2_X1 U7398 ( .A1(n6124), .A2(n7317), .ZN(n5877) );
  NAND2_X1 U7399 ( .A1(n5840), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5876) );
  NAND4_X1 U7400 ( .A1(n5879), .A2(n5878), .A3(n5877), .A4(n5876), .ZN(n8462)
         );
  INV_X1 U7401 ( .A(n8462), .ZN(n7461) );
  NAND2_X1 U7402 ( .A1(n5880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5881) );
  MUX2_X1 U7403 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5881), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5882) );
  NAND2_X1 U7404 ( .A1(n5882), .A2(n4379), .ZN(n6894) );
  INV_X1 U7405 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6403) );
  OR2_X1 U7406 ( .A1(n8222), .A2(n6403), .ZN(n5883) );
  OAI211_X1 U7407 ( .C1(n5832), .C2(n6894), .A(n5884), .B(n5883), .ZN(n7297)
         );
  NAND2_X1 U7408 ( .A1(n7461), .A2(n7297), .ZN(n8294) );
  INV_X1 U7409 ( .A(n7297), .ZN(n9909) );
  NAND2_X1 U7410 ( .A1(n8462), .A2(n9909), .ZN(n8313) );
  NAND2_X1 U7411 ( .A1(n8462), .A2(n7297), .ZN(n5885) );
  NAND2_X1 U7412 ( .A1(n5840), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7413 ( .A1(n5839), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7414 ( .A1(n5886), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5887) );
  AND2_X1 U7415 ( .A1(n5899), .A2(n5887), .ZN(n7465) );
  OR2_X1 U7416 ( .A1(n6124), .A2(n7465), .ZN(n5889) );
  INV_X1 U7417 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6885) );
  OR2_X1 U7418 ( .A1(n6127), .A2(n6885), .ZN(n5888) );
  NAND4_X1 U7419 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n8461)
         );
  NAND2_X1 U7420 ( .A1(n4379), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5892) );
  MUX2_X1 U7421 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5892), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5894) );
  AND2_X1 U7422 ( .A1(n5894), .A2(n5893), .ZN(n6985) );
  INV_X1 U7423 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6406) );
  OR2_X1 U7424 ( .A1(n8222), .A2(n6406), .ZN(n5895) );
  OAI211_X1 U7425 ( .C1(n5832), .C2(n7000), .A(n5896), .B(n5895), .ZN(n7464)
         );
  NAND2_X1 U7426 ( .A1(n7519), .A2(n7464), .ZN(n8316) );
  INV_X1 U7427 ( .A(n7464), .ZN(n7421) );
  NAND2_X1 U7428 ( .A1(n8461), .A2(n7421), .ZN(n7388) );
  NAND2_X1 U7429 ( .A1(n7267), .A2(n5897), .ZN(n7268) );
  NAND2_X1 U7430 ( .A1(n7519), .A2(n7421), .ZN(n5898) );
  NAND2_X1 U7431 ( .A1(n5839), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7432 ( .A1(n5840), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7433 ( .A1(n5899), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5900) );
  AND2_X1 U7434 ( .A1(n5909), .A2(n5900), .ZN(n7528) );
  OR2_X1 U7435 ( .A1(n6124), .A2(n7528), .ZN(n5902) );
  NAND2_X1 U7436 ( .A1(n5838), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5901) );
  NAND4_X1 U7437 ( .A1(n5904), .A2(n5903), .A3(n5902), .A4(n5901), .ZN(n8460)
         );
  INV_X1 U7438 ( .A(n8460), .ZN(n7538) );
  NAND2_X1 U7439 ( .A1(n5893), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5905) );
  XNOR2_X1 U7440 ( .A(n5905), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7003) );
  NAND2_X1 U7441 ( .A1(n6385), .A2(n7003), .ZN(n5906) );
  OAI211_X1 U7442 ( .C1(n8222), .C2(n6413), .A(n5907), .B(n5906), .ZN(n7525)
         );
  NAND2_X1 U7443 ( .A1(n7538), .A2(n7525), .ZN(n8317) );
  INV_X1 U7444 ( .A(n7525), .ZN(n9914) );
  NAND2_X1 U7445 ( .A1(n8460), .A2(n9914), .ZN(n8298) );
  NAND2_X1 U7446 ( .A1(n8317), .A2(n8298), .ZN(n8251) );
  NAND2_X1 U7447 ( .A1(n8460), .A2(n7525), .ZN(n5908) );
  NAND2_X1 U7448 ( .A1(n5840), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5914) );
  NAND2_X1 U7449 ( .A1(n5839), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7450 ( .A1(n5909), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5910) );
  AND2_X1 U7451 ( .A1(n5927), .A2(n5910), .ZN(n7550) );
  OR2_X1 U7452 ( .A1(n6124), .A2(n7550), .ZN(n5912) );
  INV_X1 U7453 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7093) );
  OR2_X1 U7454 ( .A1(n6127), .A2(n7093), .ZN(n5911) );
  NAND4_X1 U7455 ( .A1(n5914), .A2(n5913), .A3(n5912), .A4(n5911), .ZN(n8459)
         );
  INV_X1 U7456 ( .A(n8459), .ZN(n7592) );
  NAND2_X1 U7457 ( .A1(n6421), .A2(n8224), .ZN(n5917) );
  NOR2_X1 U7458 ( .A1(n5893), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5920) );
  OR2_X1 U7459 ( .A1(n5920), .A2(n4837), .ZN(n5915) );
  XNOR2_X1 U7460 ( .A(n5915), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7175) );
  AOI22_X1 U7461 ( .A1(n6026), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6385), .B2(
        n7175), .ZN(n5916) );
  NAND2_X1 U7462 ( .A1(n5917), .A2(n5916), .ZN(n7543) );
  NAND2_X1 U7463 ( .A1(n7592), .A2(n7543), .ZN(n8319) );
  NAND2_X1 U7464 ( .A1(n7581), .A2(n8459), .ZN(n8299) );
  NAND2_X1 U7465 ( .A1(n8319), .A2(n8299), .ZN(n8252) );
  NAND2_X1 U7466 ( .A1(n7592), .A2(n7581), .ZN(n5918) );
  NAND2_X1 U7467 ( .A1(n7492), .A2(n5918), .ZN(n7532) );
  NAND2_X1 U7468 ( .A1(n6425), .A2(n8224), .ZN(n5926) );
  NOR2_X1 U7469 ( .A1(n5923), .A2(n4837), .ZN(n5921) );
  MUX2_X1 U7470 ( .A(n4837), .B(n5921), .S(P2_IR_REG_10__SCAN_IN), .Z(n5924)
         );
  AOI22_X1 U7471 ( .A1(n6026), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6385), .B2(
        n7196), .ZN(n5925) );
  NAND2_X1 U7472 ( .A1(n5840), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7473 ( .A1(n5839), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7474 ( .A1(n5927), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5928) );
  AND2_X1 U7475 ( .A1(n5938), .A2(n5928), .ZN(n7598) );
  OR2_X1 U7476 ( .A1(n6124), .A2(n7598), .ZN(n5930) );
  NAND2_X1 U7477 ( .A1(n5838), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5929) );
  NAND4_X1 U7478 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(n8458)
         );
  OR2_X1 U7479 ( .A1(n9919), .A2(n8458), .ZN(n8330) );
  NAND2_X1 U7480 ( .A1(n9919), .A2(n8458), .ZN(n8325) );
  NAND2_X1 U7481 ( .A1(n8330), .A2(n8325), .ZN(n7530) );
  NAND2_X1 U7482 ( .A1(n7532), .A2(n7530), .ZN(n5934) );
  INV_X1 U7483 ( .A(n8458), .ZN(n7557) );
  NAND2_X1 U7484 ( .A1(n9919), .A2(n7557), .ZN(n5933) );
  NAND2_X1 U7485 ( .A1(n6512), .A2(n8224), .ZN(n5937) );
  OR2_X1 U7486 ( .A1(n5945), .A2(n4837), .ZN(n5935) );
  XNOR2_X1 U7487 ( .A(n5935), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7426) );
  AOI22_X1 U7488 ( .A1(n6026), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6385), .B2(
        n7426), .ZN(n5936) );
  NAND2_X1 U7489 ( .A1(n5937), .A2(n5936), .ZN(n8164) );
  NAND2_X1 U7490 ( .A1(n5840), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5943) );
  INV_X1 U7491 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7247) );
  OR2_X1 U7492 ( .A1(n6029), .A2(n7247), .ZN(n5942) );
  NAND2_X1 U7493 ( .A1(n5938), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5939) );
  AND2_X1 U7494 ( .A1(n5956), .A2(n5939), .ZN(n8165) );
  OR2_X1 U7495 ( .A1(n6124), .A2(n8165), .ZN(n5941) );
  INV_X1 U7496 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7246) );
  OR2_X1 U7497 ( .A1(n6127), .A2(n7246), .ZN(n5940) );
  NOR2_X1 U7498 ( .A1(n8164), .A2(n8457), .ZN(n7564) );
  INV_X1 U7499 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7500 ( .A1(n5945), .A2(n5944), .ZN(n5953) );
  NAND2_X1 U7501 ( .A1(n5946), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5968) );
  XNOR2_X1 U7502 ( .A(n5968), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8495) );
  AOI22_X1 U7503 ( .A1(n6026), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6385), .B2(
        n8495), .ZN(n5947) );
  NAND2_X1 U7504 ( .A1(n5840), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U7505 ( .A1(n5839), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7506 ( .A1(n5958), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5948) );
  AND2_X1 U7507 ( .A1(n5975), .A2(n5948), .ZN(n8826) );
  OR2_X1 U7508 ( .A1(n6124), .A2(n8826), .ZN(n5950) );
  INV_X1 U7509 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8473) );
  OR2_X1 U7510 ( .A1(n6127), .A2(n8473), .ZN(n5949) );
  NAND4_X1 U7511 ( .A1(n5952), .A2(n5951), .A3(n5950), .A4(n5949), .ZN(n8456)
         );
  INV_X1 U7512 ( .A(n8456), .ZN(n9709) );
  NAND2_X1 U7513 ( .A1(n5953), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U7514 ( .A(n5954), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8483) );
  AOI22_X1 U7515 ( .A1(n6026), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6385), .B2(
        n8483), .ZN(n5955) );
  NAND2_X1 U7516 ( .A1(n5840), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7517 ( .A1(n5839), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7518 ( .A1(n5956), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5957) );
  AND2_X1 U7519 ( .A1(n5958), .A2(n5957), .ZN(n7615) );
  OR2_X1 U7520 ( .A1(n6124), .A2(n7615), .ZN(n5960) );
  NAND2_X1 U7521 ( .A1(n5838), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5959) );
  NAND4_X1 U7522 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n8821)
         );
  NAND2_X1 U7523 ( .A1(n9931), .A2(n8821), .ZN(n8813) );
  INV_X1 U7524 ( .A(n8813), .ZN(n5963) );
  NAND2_X1 U7525 ( .A1(n8828), .A2(n5963), .ZN(n5965) );
  NAND2_X1 U7526 ( .A1(n8825), .A2(n8456), .ZN(n5964) );
  OR2_X1 U7527 ( .A1(n9931), .A2(n8167), .ZN(n8358) );
  NAND2_X1 U7528 ( .A1(n9931), .A2(n8167), .ZN(n8335) );
  NAND2_X1 U7529 ( .A1(n8358), .A2(n8335), .ZN(n8811) );
  AND2_X1 U7530 ( .A1(n8811), .A2(n8828), .ZN(n5966) );
  NAND2_X1 U7531 ( .A1(n6591), .A2(n8224), .ZN(n5974) );
  INV_X1 U7532 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7533 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  NAND2_X1 U7534 ( .A1(n5969), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5971) );
  INV_X1 U7535 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5970) );
  OR2_X1 U7536 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  NAND2_X1 U7537 ( .A1(n5971), .A2(n5970), .ZN(n5990) );
  AOI22_X1 U7538 ( .A1(n6026), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6385), .B2(
        n8515), .ZN(n5973) );
  NAND2_X1 U7539 ( .A1(n5974), .A2(n5973), .ZN(n9726) );
  INV_X1 U7540 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8500) );
  OR2_X1 U7541 ( .A1(n6029), .A2(n8500), .ZN(n5980) );
  NAND2_X1 U7542 ( .A1(n5840), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7543 ( .A1(n5975), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5976) );
  AND2_X1 U7544 ( .A1(n5993), .A2(n5976), .ZN(n9698) );
  OR2_X1 U7545 ( .A1(n6124), .A2(n9698), .ZN(n5978) );
  INV_X1 U7546 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8499) );
  OR2_X1 U7547 ( .A1(n6127), .A2(n8499), .ZN(n5977) );
  NAND4_X1 U7548 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(n8820)
         );
  XNOR2_X1 U7549 ( .A(n9726), .B(n8339), .ZN(n9705) );
  INV_X1 U7550 ( .A(n9705), .ZN(n6180) );
  OR2_X1 U7551 ( .A1(n9701), .A2(n6180), .ZN(n5989) );
  INV_X1 U7552 ( .A(n5981), .ZN(n5985) );
  NAND2_X1 U7553 ( .A1(n8164), .A2(n8457), .ZN(n7565) );
  NAND2_X1 U7554 ( .A1(n9726), .A2(n8820), .ZN(n5986) );
  AND2_X1 U7555 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  NAND2_X1 U7556 ( .A1(n5990), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5991) );
  XNOR2_X1 U7557 ( .A(n5991), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8565) );
  AOI22_X1 U7558 ( .A1(n6026), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8565), .B2(
        n6385), .ZN(n5992) );
  NAND2_X1 U7559 ( .A1(n5840), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7560 ( .A1(n5839), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7561 ( .A1(n5993), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5994) );
  AND2_X1 U7562 ( .A1(n6007), .A2(n5994), .ZN(n8204) );
  OR2_X1 U7563 ( .A1(n6124), .A2(n8204), .ZN(n5997) );
  INV_X1 U7564 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5995) );
  OR2_X1 U7565 ( .A1(n6127), .A2(n5995), .ZN(n5996) );
  NAND4_X1 U7566 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(n8455)
         );
  OR2_X1 U7567 ( .A1(n9719), .A2(n9711), .ZN(n8351) );
  AOI22_X1 U7568 ( .A1(n8797), .A2(n8802), .B1(n8455), .B2(n9719), .ZN(n8786)
         );
  NAND2_X1 U7569 ( .A1(n6859), .A2(n8224), .ZN(n6006) );
  NOR2_X1 U7570 ( .A1(n6000), .A2(n4837), .ZN(n6001) );
  MUX2_X1 U7571 ( .A(n4837), .B(n6001), .S(P2_IR_REG_16__SCAN_IN), .Z(n6002)
         );
  INV_X1 U7572 ( .A(n6002), .ZN(n6004) );
  AND2_X1 U7573 ( .A1(n6004), .A2(n6003), .ZN(n8582) );
  AOI22_X1 U7574 ( .A1(n6026), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6385), .B2(
        n8582), .ZN(n6005) );
  NAND2_X1 U7575 ( .A1(n5840), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6012) );
  INV_X1 U7576 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8790) );
  OR2_X1 U7577 ( .A1(n6029), .A2(n8790), .ZN(n6011) );
  NAND2_X1 U7578 ( .A1(n6007), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6008) );
  AND2_X1 U7579 ( .A1(n6017), .A2(n6008), .ZN(n8789) );
  OR2_X1 U7580 ( .A1(n6124), .A2(n8789), .ZN(n6010) );
  INV_X1 U7581 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8879) );
  OR2_X1 U7582 ( .A1(n6127), .A2(n8879), .ZN(n6009) );
  NAND4_X1 U7583 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n8799)
         );
  NAND2_X1 U7584 ( .A1(n8878), .A2(n8208), .ZN(n8367) );
  INV_X1 U7585 ( .A(n8878), .ZN(n6013) );
  NAND2_X1 U7586 ( .A1(n7130), .A2(n8224), .ZN(n6016) );
  NAND2_X1 U7587 ( .A1(n6003), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6014) );
  XNOR2_X1 U7588 ( .A(n6014), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8605) );
  AOI22_X1 U7589 ( .A1(n6026), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6385), .B2(
        n8605), .ZN(n6015) );
  NAND2_X1 U7590 ( .A1(n5840), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7591 ( .A1(n5839), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7592 ( .A1(n6017), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6018) );
  AND2_X1 U7593 ( .A1(n6030), .A2(n6018), .ZN(n8107) );
  OR2_X1 U7594 ( .A1(n6124), .A2(n8107), .ZN(n6020) );
  INV_X1 U7595 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8873) );
  OR2_X1 U7596 ( .A1(n6127), .A2(n8873), .ZN(n6019) );
  NAND4_X1 U7597 ( .A1(n6022), .A2(n6021), .A3(n6020), .A4(n6019), .ZN(n8768)
         );
  NAND2_X1 U7598 ( .A1(n8945), .A2(n8788), .ZN(n8242) );
  NAND2_X1 U7599 ( .A1(n8761), .A2(n8242), .ZN(n8366) );
  AOI21_X1 U7600 ( .B1(n8778), .B2(n8366), .A(n6023), .ZN(n8766) );
  NAND2_X1 U7601 ( .A1(n7154), .A2(n8224), .ZN(n6028) );
  INV_X1 U7602 ( .A(n5798), .ZN(n6024) );
  NAND2_X1 U7603 ( .A1(n6024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6025) );
  XNOR2_X1 U7604 ( .A(n6025), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8624) );
  AOI22_X1 U7605 ( .A1(n6026), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6385), .B2(
        n8624), .ZN(n6027) );
  INV_X1 U7606 ( .A(n8938), .ZN(n8188) );
  NAND2_X1 U7607 ( .A1(n5840), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6036) );
  INV_X1 U7608 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8771) );
  OR2_X1 U7609 ( .A1(n6029), .A2(n8771), .ZN(n6035) );
  NAND2_X1 U7610 ( .A1(n6030), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6031) );
  AND2_X1 U7611 ( .A1(n6032), .A2(n6031), .ZN(n8772) );
  OR2_X1 U7612 ( .A1(n6124), .A2(n8772), .ZN(n6034) );
  INV_X1 U7613 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8870) );
  OR2_X1 U7614 ( .A1(n6127), .A2(n8870), .ZN(n6033) );
  NAND2_X1 U7615 ( .A1(n7401), .A2(n8224), .ZN(n6039) );
  INV_X1 U7616 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7402) );
  OR2_X1 U7617 ( .A1(n8222), .A2(n7402), .ZN(n6038) );
  NAND2_X1 U7618 ( .A1(n5839), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6043) );
  XNOR2_X1 U7619 ( .A(n6046), .B(n10038), .ZN(n8747) );
  OR2_X1 U7620 ( .A1(n6124), .A2(n8747), .ZN(n6042) );
  INV_X1 U7621 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8864) );
  OR2_X1 U7622 ( .A1(n6127), .A2(n8864), .ZN(n6041) );
  INV_X1 U7623 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8925) );
  OR2_X1 U7624 ( .A1(n5786), .A2(n8925), .ZN(n6040) );
  NAND2_X1 U7625 ( .A1(n8926), .A2(n8068), .ZN(n8726) );
  NAND2_X1 U7626 ( .A1(n8383), .A2(n8726), .ZN(n8742) );
  INV_X1 U7627 ( .A(n8926), .ZN(n8135) );
  NAND2_X1 U7628 ( .A1(n8135), .A2(n8068), .ZN(n8730) );
  NAND2_X1 U7629 ( .A1(n7489), .A2(n8224), .ZN(n6045) );
  OR2_X1 U7630 ( .A1(n8222), .A2(n7490), .ZN(n6044) );
  NAND2_X1 U7631 ( .A1(n5840), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6051) );
  OAI21_X1 U7632 ( .B1(n6046), .B2(P2_REG3_REG_20__SCAN_IN), .A(
        P2_REG3_REG_21__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7633 ( .A1(n6047), .A2(n6056), .ZN(n8737) );
  NAND2_X1 U7634 ( .A1(n5822), .A2(n8737), .ZN(n6050) );
  NAND2_X1 U7635 ( .A1(n5839), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7636 ( .A1(n5838), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6048) );
  NAND4_X1 U7637 ( .A1(n6051), .A2(n6050), .A3(n6049), .A4(n6048), .ZN(n8744)
         );
  INV_X1 U7638 ( .A(n8744), .ZN(n8130) );
  NAND2_X1 U7639 ( .A1(n8920), .A2(n8130), .ZN(n8378) );
  NOR2_X1 U7640 ( .A1(n8920), .A2(n8744), .ZN(n8717) );
  NAND2_X1 U7641 ( .A1(n7551), .A2(n8224), .ZN(n6053) );
  OR2_X1 U7642 ( .A1(n8222), .A2(n7553), .ZN(n6052) );
  INV_X1 U7643 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U7644 ( .A1(n5840), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7645 ( .A1(n5839), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6054) );
  AND2_X1 U7646 ( .A1(n6055), .A2(n6054), .ZN(n6060) );
  NAND2_X1 U7647 ( .A1(n6056), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7648 ( .A1(n6058), .A2(n6057), .ZN(n8723) );
  NAND2_X1 U7649 ( .A1(n8723), .A2(n5822), .ZN(n6059) );
  OAI211_X1 U7650 ( .C1(n6127), .C2(n8858), .A(n6060), .B(n6059), .ZN(n8734)
         );
  INV_X1 U7651 ( .A(n8734), .ZN(n8708) );
  NAND2_X1 U7652 ( .A1(n8914), .A2(n8708), .ZN(n8389) );
  NAND2_X1 U7653 ( .A1(n8388), .A2(n8389), .ZN(n8716) );
  INV_X1 U7654 ( .A(n8712), .ZN(n8908) );
  NAND2_X1 U7655 ( .A1(n7589), .A2(n8224), .ZN(n6063) );
  OR2_X1 U7656 ( .A1(n8222), .A2(n7624), .ZN(n6062) );
  INV_X1 U7657 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U7658 ( .A1(n6064), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7659 ( .A1(n6072), .A2(n6065), .ZN(n8696) );
  NAND2_X1 U7660 ( .A1(n8696), .A2(n5822), .ZN(n6067) );
  AOI22_X1 U7661 ( .A1(n5838), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n5839), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n6066) );
  OAI211_X1 U7662 ( .C1(n5786), .C2(n8901), .A(n6067), .B(n6066), .ZN(n8680)
         );
  NOR2_X1 U7663 ( .A1(n8902), .A2(n8680), .ZN(n6068) );
  INV_X1 U7664 ( .A(n8902), .ZN(n8852) );
  NAND2_X1 U7665 ( .A1(n7626), .A2(n8224), .ZN(n6070) );
  OR2_X1 U7666 ( .A1(n8222), .A2(n7635), .ZN(n6069) );
  INV_X1 U7667 ( .A(n6072), .ZN(n6071) );
  NAND2_X1 U7668 ( .A1(n6071), .A2(n10076), .ZN(n6083) );
  NAND2_X1 U7669 ( .A1(n6072), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7670 ( .A1(n6083), .A2(n6073), .ZN(n8685) );
  NAND2_X1 U7671 ( .A1(n8685), .A2(n5822), .ZN(n6078) );
  INV_X1 U7672 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U7673 ( .A1(n5839), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7674 ( .A1(n5840), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6074) );
  OAI211_X1 U7675 ( .C1(n6127), .C2(n8848), .A(n6075), .B(n6074), .ZN(n6076)
         );
  INV_X1 U7676 ( .A(n6076), .ZN(n6077) );
  NAND2_X1 U7677 ( .A1(n8895), .A2(n8693), .ZN(n8404) );
  INV_X1 U7678 ( .A(n8895), .ZN(n8677) );
  NAND2_X1 U7679 ( .A1(n7629), .A2(n8224), .ZN(n6080) );
  OR2_X1 U7680 ( .A1(n8222), .A2(n7630), .ZN(n6079) );
  INV_X1 U7681 ( .A(n6083), .ZN(n6082) );
  INV_X1 U7682 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7683 ( .A1(n6082), .A2(n6081), .ZN(n6092) );
  NAND2_X1 U7684 ( .A1(n6083), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7685 ( .A1(n6092), .A2(n6084), .ZN(n8672) );
  NAND2_X1 U7686 ( .A1(n8672), .A2(n5822), .ZN(n6089) );
  INV_X1 U7687 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8846) );
  NAND2_X1 U7688 ( .A1(n5840), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7689 ( .A1(n5839), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6085) );
  OAI211_X1 U7690 ( .C1(n8846), .C2(n6127), .A(n6086), .B(n6085), .ZN(n6087)
         );
  INV_X1 U7691 ( .A(n6087), .ZN(n6088) );
  NAND2_X1 U7692 ( .A1(n9690), .A2(n8224), .ZN(n6091) );
  OR2_X1 U7693 ( .A1(n8222), .A2(n8972), .ZN(n6090) );
  INV_X1 U7694 ( .A(n8661), .ZN(n8840) );
  NAND2_X1 U7695 ( .A1(n6092), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7696 ( .A1(n6110), .A2(n6093), .ZN(n8660) );
  NAND2_X1 U7697 ( .A1(n8660), .A2(n5822), .ZN(n6099) );
  INV_X1 U7698 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7699 ( .A1(n5840), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7700 ( .A1(n5839), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6094) );
  OAI211_X1 U7701 ( .C1(n6096), .C2(n6127), .A(n6095), .B(n6094), .ZN(n6097)
         );
  INV_X1 U7702 ( .A(n6097), .ZN(n6098) );
  NAND2_X1 U7703 ( .A1(n8840), .A2(n8668), .ZN(n6100) );
  NAND2_X1 U7704 ( .A1(n6217), .A2(n6100), .ZN(n6102) );
  NAND2_X1 U7705 ( .A1(n8661), .A2(n8453), .ZN(n6101) );
  MUX2_X1 U7706 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6389), .Z(n6230) );
  XNOR2_X1 U7707 ( .A(n6230), .B(n10071), .ZN(n6228) );
  NAND2_X1 U7708 ( .A1(n8965), .A2(n8224), .ZN(n6107) );
  INV_X1 U7709 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8968) );
  OR2_X1 U7710 ( .A1(n8222), .A2(n8968), .ZN(n6106) );
  INV_X1 U7711 ( .A(n6110), .ZN(n6109) );
  INV_X1 U7712 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7713 ( .A1(n6109), .A2(n6108), .ZN(n8644) );
  NAND2_X1 U7714 ( .A1(n6110), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7715 ( .A1(n8644), .A2(n6111), .ZN(n8031) );
  INV_X1 U7716 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7717 ( .A1(n5840), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7718 ( .A1(n5839), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6112) );
  OAI211_X1 U7719 ( .C1(n6276), .C2(n6127), .A(n6113), .B(n6112), .ZN(n6114)
         );
  INV_X1 U7720 ( .A(n6135), .ZN(n6117) );
  NAND2_X1 U7721 ( .A1(n6121), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7722 ( .A1(n4395), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6120) );
  MUX2_X1 U7723 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6120), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6122) );
  NOR2_X1 U7724 ( .A1(n8269), .A2(n8423), .ZN(n6123) );
  OR2_X1 U7725 ( .A1(n8644), .A2(n6124), .ZN(n8235) );
  INV_X1 U7726 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7727 ( .A1(n5840), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7728 ( .A1(n5839), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6125) );
  OAI211_X1 U7729 ( .C1(n6254), .C2(n6127), .A(n6126), .B(n6125), .ZN(n6128)
         );
  INV_X1 U7730 ( .A(n6128), .ZN(n6129) );
  INV_X2 U7731 ( .A(n6686), .ZN(n8626) );
  OAI22_X1 U7732 ( .A1(n8034), .A2(n9712), .B1(n8668), .B2(n9710), .ZN(n6132)
         );
  AOI21_X1 U7733 ( .B1(n6133), .B2(n8817), .A(n6132), .ZN(n6274) );
  AOI21_X1 U7734 ( .B1(n6135), .B2(n6134), .A(n4837), .ZN(n6136) );
  XNOR2_X1 U7735 ( .A(n6145), .B(P2_B_REG_SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7736 ( .A1(n6148), .A2(n6141), .ZN(n6144) );
  NAND2_X1 U7737 ( .A1(n6142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7738 ( .A1(n6145), .A2(n7631), .ZN(n6578) );
  INV_X1 U7739 ( .A(n7019), .ZN(n6151) );
  NAND2_X1 U7740 ( .A1(n6148), .A2(n7631), .ZN(n6149) );
  NAND2_X1 U7741 ( .A1(n6151), .A2(n6491), .ZN(n6249) );
  NOR2_X1 U7742 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6155) );
  NOR4_X1 U7743 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6154) );
  NOR4_X1 U7744 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6153) );
  NOR4_X1 U7745 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6152) );
  NAND4_X1 U7746 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(n6161)
         );
  NOR4_X1 U7747 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6159) );
  NOR4_X1 U7748 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6158) );
  NOR4_X1 U7749 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6157) );
  NOR4_X1 U7750 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6156) );
  NAND4_X1 U7751 ( .A1(n6159), .A2(n6158), .A3(n6157), .A4(n6156), .ZN(n6160)
         );
  NOR2_X1 U7752 ( .A1(n6161), .A2(n6160), .ZN(n6162) );
  INV_X1 U7753 ( .A(n6247), .ZN(n6163) );
  INV_X1 U7754 ( .A(n6148), .ZN(n6165) );
  NAND2_X1 U7755 ( .A1(n8423), .A2(n8638), .ZN(n7017) );
  NAND2_X1 U7756 ( .A1(n8269), .A2(n8433), .ZN(n8266) );
  INV_X1 U7757 ( .A(n8266), .ZN(n6169) );
  NAND2_X1 U7758 ( .A1(n6170), .A2(n6169), .ZN(n6923) );
  AND2_X1 U7759 ( .A1(n6978), .A2(n6923), .ZN(n6171) );
  NAND3_X1 U7760 ( .A1(n7019), .A2(n6259), .A3(n6247), .ZN(n6940) );
  NAND2_X1 U7761 ( .A1(n7552), .A2(n8269), .ZN(n9925) );
  AND2_X1 U7762 ( .A1(n8412), .A2(n9925), .ZN(n6172) );
  NAND2_X1 U7763 ( .A1(n6923), .A2(n6172), .ZN(n6921) );
  NAND2_X1 U7764 ( .A1(n8423), .A2(n8443), .ZN(n6186) );
  NAND2_X1 U7765 ( .A1(n6921), .A2(n9699), .ZN(n6929) );
  NAND2_X1 U7766 ( .A1(n6924), .A2(n6929), .ZN(n6173) );
  INV_X1 U7767 ( .A(n6176), .ZN(n7135) );
  NAND2_X1 U7768 ( .A1(n7134), .A2(n7135), .ZN(n7136) );
  NAND2_X1 U7769 ( .A1(n7136), .A2(n8279), .ZN(n6842) );
  INV_X1 U7770 ( .A(n8245), .ZN(n6846) );
  NAND2_X1 U7771 ( .A1(n6842), .A2(n6846), .ZN(n6841) );
  NAND2_X1 U7772 ( .A1(n6841), .A2(n8280), .ZN(n6177) );
  NAND2_X1 U7773 ( .A1(n6177), .A2(n8287), .ZN(n7051) );
  INV_X1 U7774 ( .A(n8464), .ZN(n7236) );
  NAND2_X1 U7775 ( .A1(n7236), .A2(n8306), .ZN(n8291) );
  NAND2_X1 U7776 ( .A1(n7051), .A2(n8291), .ZN(n7277) );
  NAND2_X1 U7777 ( .A1(n7294), .A2(n7239), .ZN(n8290) );
  INV_X1 U7778 ( .A(n7239), .ZN(n9903) );
  NAND2_X1 U7779 ( .A1(n8463), .A2(n9903), .ZN(n8307) );
  AND2_X1 U7780 ( .A1(n8294), .A2(n8290), .ZN(n8311) );
  AND2_X1 U7781 ( .A1(n8298), .A2(n7388), .ZN(n8296) );
  NAND2_X1 U7782 ( .A1(n7270), .A2(n8296), .ZN(n6178) );
  AND2_X1 U7783 ( .A1(n8325), .A2(n8299), .ZN(n8303) );
  NAND2_X1 U7784 ( .A1(n6179), .A2(n8330), .ZN(n7559) );
  OR2_X1 U7785 ( .A1(n8164), .A2(n7607), .ZN(n8332) );
  NAND2_X1 U7786 ( .A1(n8164), .A2(n7607), .ZN(n8331) );
  INV_X1 U7787 ( .A(n8357), .ZN(n8346) );
  AND2_X1 U7788 ( .A1(n9726), .A2(n8339), .ZN(n8342) );
  AOI21_X1 U7789 ( .B1(n9696), .B2(n6180), .A(n8342), .ZN(n8803) );
  INV_X1 U7790 ( .A(n8351), .ZN(n6181) );
  AOI21_X1 U7791 ( .B1(n8803), .B2(n8348), .A(n6181), .ZN(n8784) );
  INV_X1 U7792 ( .A(n8367), .ZN(n6182) );
  OAI21_X1 U7793 ( .B1(n8784), .B2(n6182), .A(n8368), .ZN(n8776) );
  NAND2_X1 U7794 ( .A1(n8776), .A2(n8242), .ZN(n8762) );
  OR2_X1 U7795 ( .A1(n8938), .A2(n7991), .ZN(n8372) );
  AND2_X1 U7796 ( .A1(n8372), .A2(n8761), .ZN(n8371) );
  AOI21_X1 U7797 ( .B1(n8762), .B2(n8371), .A(n8763), .ZN(n8751) );
  NAND2_X1 U7798 ( .A1(n8932), .A2(n8182), .ZN(n8380) );
  NOR2_X1 U7799 ( .A1(n8932), .A2(n8182), .ZN(n8381) );
  AOI21_X1 U7800 ( .B1(n8751), .B2(n8380), .A(n8381), .ZN(n8740) );
  NAND2_X1 U7801 ( .A1(n8740), .A2(n8383), .ZN(n8727) );
  AND2_X1 U7802 ( .A1(n8378), .A2(n8726), .ZN(n8384) );
  NOR2_X1 U7803 ( .A1(n8712), .A2(n8694), .ZN(n8392) );
  NAND2_X1 U7804 ( .A1(n8902), .A2(n8707), .ZN(n8394) );
  NAND2_X1 U7805 ( .A1(n8712), .A2(n8694), .ZN(n8391) );
  NAND2_X1 U7806 ( .A1(n8394), .A2(n8391), .ZN(n8396) );
  INV_X1 U7807 ( .A(n8403), .ZN(n6183) );
  AOI21_X1 U7808 ( .B1(n8687), .B2(n8404), .A(n6183), .ZN(n8670) );
  AND2_X1 U7809 ( .A1(n8671), .A2(n8090), .ZN(n8240) );
  XNOR2_X1 U7810 ( .A(n8661), .B(n8453), .ZN(n8410) );
  NOR2_X1 U7811 ( .A1(n8661), .A2(n8668), .ZN(n8413) );
  XNOR2_X1 U7812 ( .A(n6236), .B(n8239), .ZN(n6275) );
  OAI211_X1 U7813 ( .C1(n8448), .C2(n8423), .A(n9925), .B(n8638), .ZN(n6184)
         );
  INV_X1 U7814 ( .A(n6184), .ZN(n6185) );
  INV_X1 U7815 ( .A(n6186), .ZN(n6266) );
  NAND2_X1 U7816 ( .A1(n8267), .A2(n8944), .ZN(n6188) );
  NAND2_X1 U7817 ( .A1(n8965), .A2(n7781), .ZN(n6192) );
  INV_X1 U7818 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7969) );
  OR2_X1 U7819 ( .A1(n7782), .A2(n7969), .ZN(n6191) );
  NAND2_X1 U7820 ( .A1(n9536), .A2(n6193), .ZN(n6195) );
  NAND2_X1 U7821 ( .A1(n9127), .A2(n6197), .ZN(n6194) );
  NAND2_X1 U7822 ( .A1(n6195), .A2(n6194), .ZN(n6196) );
  XNOR2_X1 U7823 ( .A(n6196), .B(n5139), .ZN(n6200) );
  NAND2_X1 U7824 ( .A1(n9536), .A2(n6197), .ZN(n6198) );
  OAI21_X1 U7825 ( .B1(n9315), .B2(n5656), .A(n6198), .ZN(n6199) );
  XNOR2_X1 U7826 ( .A(n6200), .B(n6199), .ZN(n6205) );
  INV_X1 U7827 ( .A(n6205), .ZN(n6202) );
  INV_X1 U7828 ( .A(n6204), .ZN(n6201) );
  NOR2_X1 U7829 ( .A1(n9304), .A2(n9083), .ZN(n6213) );
  INV_X1 U7830 ( .A(n9282), .ZN(n6209) );
  INV_X1 U7831 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U7832 ( .A1(n5073), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7833 ( .A1(n7651), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6206) );
  OAI211_X1 U7834 ( .C1(n7655), .C2(n9281), .A(n6207), .B(n6206), .ZN(n6208)
         );
  AOI21_X1 U7835 ( .B1(n6209), .B2(n5619), .A(n6208), .ZN(n9303) );
  NAND2_X1 U7836 ( .A1(P1_U3086), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7837 ( .A1(n9293), .A2(n9121), .ZN(n6210) );
  OAI211_X1 U7838 ( .C1(n9303), .C2(n9119), .A(n6211), .B(n6210), .ZN(n6212)
         );
  AOI211_X1 U7839 ( .C1(n9536), .C2(n9096), .A(n6213), .B(n6212), .ZN(n6214)
         );
  INV_X1 U7840 ( .A(n6214), .ZN(n6215) );
  XNOR2_X1 U7841 ( .A(n6217), .B(n8410), .ZN(n6218) );
  NAND2_X1 U7842 ( .A1(n6218), .A2(n8817), .ZN(n6221) );
  OAI22_X1 U7843 ( .A1(n8042), .A2(n9712), .B1(n9710), .B2(n8090), .ZN(n6219)
         );
  INV_X1 U7844 ( .A(n6219), .ZN(n6220) );
  NAND2_X1 U7845 ( .A1(n6221), .A2(n6220), .ZN(n8839) );
  MUX2_X1 U7846 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8839), .S(n9937), .Z(n6222)
         );
  INV_X1 U7847 ( .A(n6222), .ZN(n6226) );
  XOR2_X1 U7848 ( .A(n8410), .B(n6223), .Z(n8662) );
  INV_X1 U7849 ( .A(n8662), .ZN(n8841) );
  OAI22_X1 U7850 ( .A1(n8841), .A2(n8952), .B1(n8840), .B2(n8907), .ZN(n6224)
         );
  INV_X1 U7851 ( .A(n6224), .ZN(n6225) );
  INV_X1 U7852 ( .A(n6230), .ZN(n6231) );
  NAND2_X1 U7853 ( .A1(n6231), .A2(n10071), .ZN(n6232) );
  NAND2_X1 U7854 ( .A1(n6233), .A2(n6232), .ZN(n7638) );
  INV_X1 U7855 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8961) );
  INV_X1 U7856 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7960) );
  MUX2_X1 U7857 ( .A(n8961), .B(n7960), .S(n6389), .Z(n7637) );
  XNOR2_X1 U7858 ( .A(n7640), .B(SI_29_), .ZN(n7959) );
  NAND2_X1 U7859 ( .A1(n7959), .A2(n8224), .ZN(n6235) );
  OR2_X1 U7860 ( .A1(n8222), .A2(n8961), .ZN(n6234) );
  NAND2_X1 U7861 ( .A1(n6235), .A2(n6234), .ZN(n6282) );
  OR2_X1 U7862 ( .A1(n6282), .A2(n8034), .ZN(n8214) );
  NAND2_X1 U7863 ( .A1(n6282), .A2(n8034), .ZN(n8220) );
  NAND2_X1 U7864 ( .A1(n5838), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7865 ( .A1(n5840), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7866 ( .A1(n5839), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6237) );
  AND3_X1 U7867 ( .A1(n6239), .A2(n6238), .A3(n6237), .ZN(n6240) );
  NAND2_X1 U7868 ( .A1(n5832), .A2(P2_B_REG_SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7869 ( .A1(n8819), .A2(n6241), .ZN(n8645) );
  OAI22_X1 U7870 ( .A1(n8042), .A2(n9710), .B1(n8228), .B2(n8645), .ZN(n6242)
         );
  OAI21_X1 U7871 ( .B1(n6244), .B2(n9708), .A(n6243), .ZN(n8651) );
  INV_X1 U7872 ( .A(n8657), .ZN(n6245) );
  NOR2_X1 U7873 ( .A1(n6245), .A2(n9892), .ZN(n6246) );
  NOR2_X1 U7874 ( .A1(n8651), .A2(n6246), .ZN(n6286) );
  NAND2_X1 U7875 ( .A1(n8432), .A2(n7017), .ZN(n6931) );
  AND3_X1 U7876 ( .A1(n6517), .A2(n6247), .A3(n6931), .ZN(n6248) );
  NAND2_X1 U7877 ( .A1(n9907), .A2(n8269), .ZN(n6264) );
  INV_X1 U7878 ( .A(n6264), .ZN(n6250) );
  NOR2_X1 U7879 ( .A1(n7019), .A2(n6250), .ZN(n6252) );
  NAND3_X1 U7880 ( .A1(n8448), .A2(n8433), .A3(n8638), .ZN(n6251) );
  MUX2_X1 U7881 ( .A(n6491), .B(n6252), .S(n6258), .Z(n6253) );
  INV_X1 U7882 ( .A(n6282), .ZN(n8654) );
  OAI21_X1 U7883 ( .B1(n6286), .B2(n6277), .A(n6256), .ZN(P2_U3488) );
  INV_X1 U7884 ( .A(n6258), .ZN(n6257) );
  NAND2_X1 U7885 ( .A1(n7019), .A2(n6257), .ZN(n6261) );
  NAND2_X1 U7886 ( .A1(n6259), .A2(n6258), .ZN(n6260) );
  INV_X1 U7887 ( .A(n9716), .ZN(n6265) );
  OR2_X1 U7888 ( .A1(n6274), .A2(n6265), .ZN(n6273) );
  NAND2_X1 U7889 ( .A1(n7015), .A2(n6266), .ZN(n7137) );
  NAND2_X1 U7890 ( .A1(n6267), .A2(n7137), .ZN(n9715) );
  AOI22_X1 U7891 ( .A1(n8267), .A2(n8792), .B1(n8805), .B2(n8031), .ZN(n6271)
         );
  INV_X1 U7892 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7893 ( .A1(n6273), .A2(n4915), .ZN(P2_U3205) );
  OR2_X1 U7894 ( .A1(n6274), .A2(n6277), .ZN(n6281) );
  NAND2_X1 U7895 ( .A1(n8267), .A2(n8874), .ZN(n6279) );
  NAND2_X1 U7896 ( .A1(n6281), .A2(n4914), .ZN(P2_U3487) );
  INV_X1 U7897 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6283) );
  NOR2_X1 U7898 ( .A1(n9937), .A2(n6283), .ZN(n6284) );
  OAI21_X1 U7899 ( .B1(n6286), .B2(n9939), .A(n6285), .ZN(P2_U3456) );
  NAND2_X1 U7900 ( .A1(n6535), .A2(n6328), .ZN(n6287) );
  XNOR2_X1 U7901 ( .A(n9143), .B(n7877), .ZN(n7805) );
  NAND2_X1 U7902 ( .A1(n6557), .A2(n7877), .ZN(n6288) );
  NAND2_X1 U7903 ( .A1(n6531), .A2(n6288), .ZN(n6563) );
  NAND2_X1 U7904 ( .A1(n9142), .A2(n6587), .ZN(n7882) );
  NAND2_X1 U7905 ( .A1(n6601), .A2(n7882), .ZN(n6564) );
  NAND2_X1 U7906 ( .A1(n6563), .A2(n6564), .ZN(n6562) );
  NAND2_X1 U7907 ( .A1(n6536), .A2(n6587), .ZN(n6289) );
  NAND2_X1 U7908 ( .A1(n6562), .A2(n6289), .ZN(n6597) );
  NAND2_X1 U7909 ( .A1(n9141), .A2(n6620), .ZN(n7881) );
  NAND2_X1 U7910 ( .A1(n6597), .A2(n7804), .ZN(n6596) );
  NAND2_X1 U7911 ( .A1(n6290), .A2(n6620), .ZN(n6291) );
  NAND2_X1 U7912 ( .A1(n6596), .A2(n6291), .ZN(n6646) );
  NAND2_X1 U7913 ( .A1(n6739), .A2(n6648), .ZN(n7674) );
  INV_X1 U7914 ( .A(n6648), .ZN(n6835) );
  NAND2_X1 U7915 ( .A1(n9140), .A2(n6835), .ZN(n7883) );
  NAND2_X1 U7916 ( .A1(n7674), .A2(n7883), .ZN(n7810) );
  NAND2_X1 U7917 ( .A1(n6646), .A2(n7810), .ZN(n6645) );
  NAND2_X1 U7918 ( .A1(n6739), .A2(n6835), .ZN(n6292) );
  NAND2_X1 U7919 ( .A1(n6645), .A2(n6292), .ZN(n6745) );
  NAND2_X1 U7920 ( .A1(n6953), .A2(n6293), .ZN(n7675) );
  NAND2_X1 U7921 ( .A1(n6914), .A2(n9139), .ZN(n7694) );
  NAND2_X1 U7922 ( .A1(n7675), .A2(n7694), .ZN(n6744) );
  NAND2_X1 U7923 ( .A1(n6745), .A2(n6744), .ZN(n6743) );
  NAND2_X1 U7924 ( .A1(n6953), .A2(n6914), .ZN(n6294) );
  NAND2_X1 U7925 ( .A1(n6743), .A2(n6294), .ZN(n6947) );
  XNOR2_X1 U7926 ( .A(n6962), .B(n6740), .ZN(n7696) );
  NAND2_X1 U7927 ( .A1(n6947), .A2(n7696), .ZN(n6296) );
  OR2_X1 U7928 ( .A1(n9138), .A2(n6962), .ZN(n6295) );
  NAND2_X1 U7929 ( .A1(n6296), .A2(n6295), .ZN(n6862) );
  NAND2_X1 U7930 ( .A1(n6875), .A2(n6952), .ZN(n7681) );
  NAND2_X1 U7931 ( .A1(n7678), .A2(n7681), .ZN(n6866) );
  NAND2_X1 U7932 ( .A1(n6862), .A2(n6866), .ZN(n6861) );
  OR2_X1 U7933 ( .A1(n6875), .A2(n9137), .ZN(n6297) );
  NAND2_X1 U7934 ( .A1(n6861), .A2(n6297), .ZN(n7042) );
  NAND2_X1 U7935 ( .A1(n7384), .A2(n7306), .ZN(n7701) );
  NAND2_X1 U7936 ( .A1(n7706), .A2(n7701), .ZN(n7041) );
  OR2_X1 U7937 ( .A1(n7384), .A2(n4726), .ZN(n6298) );
  OR2_X1 U7938 ( .A1(n7127), .A2(n7380), .ZN(n7885) );
  NAND2_X1 U7939 ( .A1(n7127), .A2(n7380), .ZN(n7707) );
  NAND2_X1 U7940 ( .A1(n7885), .A2(n7707), .ZN(n7120) );
  NAND2_X1 U7941 ( .A1(n7510), .A2(n7411), .ZN(n7710) );
  OR2_X1 U7942 ( .A1(n9622), .A2(n7328), .ZN(n7711) );
  NAND2_X1 U7943 ( .A1(n9622), .A2(n7328), .ZN(n7893) );
  NAND2_X1 U7944 ( .A1(n7220), .A2(n7225), .ZN(n7219) );
  OR2_X1 U7945 ( .A1(n9622), .A2(n9134), .ZN(n6299) );
  NAND2_X1 U7946 ( .A1(n7219), .A2(n6299), .ZN(n7364) );
  NAND2_X1 U7947 ( .A1(n7486), .A2(n7229), .ZN(n7894) );
  OR2_X1 U7948 ( .A1(n7486), .A2(n9133), .ZN(n6300) );
  NAND2_X1 U7949 ( .A1(n9611), .A2(n9523), .ZN(n6301) );
  OR2_X1 U7950 ( .A1(n9611), .A2(n9523), .ZN(n6302) );
  OR2_X1 U7951 ( .A1(n9601), .A2(n9517), .ZN(n7730) );
  NAND2_X1 U7952 ( .A1(n9601), .A2(n9517), .ZN(n7732) );
  NAND2_X1 U7953 ( .A1(n7730), .A2(n7732), .ZN(n9489) );
  NAND2_X1 U7954 ( .A1(n9601), .A2(n9475), .ZN(n6303) );
  AND2_X1 U7955 ( .A1(n9481), .A2(n9501), .ZN(n6305) );
  AND2_X1 U7956 ( .A1(n9587), .A2(n9132), .ZN(n6307) );
  NOR2_X1 U7957 ( .A1(n9582), .A2(n9131), .ZN(n6308) );
  NAND2_X1 U7958 ( .A1(n9582), .A2(n9131), .ZN(n6309) );
  OR2_X1 U7959 ( .A1(n9422), .A2(n9407), .ZN(n6310) );
  NOR2_X1 U7960 ( .A1(n9571), .A2(n9130), .ZN(n6311) );
  OR2_X1 U7961 ( .A1(n9388), .A2(n9408), .ZN(n6312) );
  OR2_X1 U7962 ( .A1(n9560), .A2(n9382), .ZN(n7834) );
  NAND2_X1 U7963 ( .A1(n9560), .A2(n9382), .ZN(n7839) );
  INV_X1 U7964 ( .A(n9382), .ZN(n9129) );
  NAND2_X1 U7965 ( .A1(n9560), .A2(n9129), .ZN(n6313) );
  OR2_X1 U7966 ( .A1(n9355), .A2(n9339), .ZN(n6314) );
  NAND2_X1 U7967 ( .A1(n9355), .A2(n9339), .ZN(n6315) );
  NAND2_X1 U7968 ( .A1(n6316), .A2(n6315), .ZN(n9329) );
  OR2_X1 U7969 ( .A1(n9549), .A2(n9350), .ZN(n7845) );
  NAND2_X1 U7970 ( .A1(n9549), .A2(n9350), .ZN(n7910) );
  NAND2_X1 U7971 ( .A1(n7845), .A2(n7910), .ZN(n9330) );
  NAND2_X1 U7972 ( .A1(n9549), .A2(n9128), .ZN(n6317) );
  OR2_X1 U7973 ( .A1(n9322), .A2(n9304), .ZN(n7916) );
  NAND2_X1 U7974 ( .A1(n9322), .A2(n9304), .ZN(n7851) );
  INV_X1 U7975 ( .A(n9313), .ZN(n6318) );
  OR2_X1 U7976 ( .A1(n9322), .A2(n9340), .ZN(n6319) );
  OR2_X1 U7977 ( .A1(n9536), .A2(n9315), .ZN(n7854) );
  NAND2_X1 U7978 ( .A1(n9536), .A2(n9315), .ZN(n7852) );
  NAND2_X1 U7979 ( .A1(n9536), .A2(n9127), .ZN(n6320) );
  NAND2_X1 U7980 ( .A1(n9290), .A2(n6320), .ZN(n6323) );
  NAND2_X1 U7981 ( .A1(n7959), .A2(n7781), .ZN(n6322) );
  OR2_X1 U7982 ( .A1(n7782), .A2(n7960), .ZN(n6321) );
  OR2_X1 U7983 ( .A1(n9284), .A2(n9303), .ZN(n7855) );
  NAND2_X1 U7984 ( .A1(n9284), .A2(n9303), .ZN(n7858) );
  XNOR2_X1 U7985 ( .A(n6323), .B(n7778), .ZN(n9280) );
  NAND2_X1 U7986 ( .A1(n6407), .A2(n5713), .ZN(n7935) );
  NAND2_X1 U7987 ( .A1(n6324), .A2(n7929), .ZN(n6326) );
  INV_X1 U7988 ( .A(n6325), .ZN(n6636) );
  NAND2_X1 U7989 ( .A1(n7935), .A2(n6327), .ZN(n7332) );
  NAND2_X1 U7990 ( .A1(n7795), .A2(n9269), .ZN(n7790) );
  OR2_X1 U7991 ( .A1(n7790), .A2(n7870), .ZN(n9627) );
  NAND2_X1 U7992 ( .A1(n9280), .A2(n9869), .ZN(n6355) );
  INV_X1 U7993 ( .A(n9582), .ZN(n9439) );
  INV_X1 U7994 ( .A(n9601), .ZN(n9495) );
  AND2_X1 U7995 ( .A1(n6746), .A2(n6914), .ZN(n6959) );
  NAND2_X1 U7996 ( .A1(n6959), .A2(n9851), .ZN(n6958) );
  OR2_X1 U7997 ( .A1(n6958), .A2(n6875), .ZN(n7044) );
  INV_X1 U7998 ( .A(n7127), .ZN(n9867) );
  OR2_X1 U7999 ( .A1(n7366), .A2(n7486), .ZN(n7471) );
  INV_X1 U8000 ( .A(n9606), .ZN(n9515) );
  AND2_X1 U8001 ( .A1(n9508), .A2(n9515), .ZN(n9509) );
  NOR2_X2 U8002 ( .A1(n9549), .A2(n9353), .ZN(n9331) );
  AOI21_X1 U8003 ( .B1(n9284), .B2(n4367), .A(n9510), .ZN(n6329) );
  NAND2_X1 U8004 ( .A1(n6329), .A2(n7944), .ZN(n9286) );
  INV_X1 U8005 ( .A(n7363), .ZN(n7820) );
  INV_X1 U8006 ( .A(n6635), .ZN(n6546) );
  NOR2_X1 U8007 ( .A1(n6540), .A2(n6546), .ZN(n6538) );
  NAND2_X1 U8008 ( .A1(n6539), .A2(n6538), .ZN(n6332) );
  NAND2_X1 U8009 ( .A1(n6535), .A2(n9837), .ZN(n6331) );
  NAND2_X1 U8010 ( .A1(n6332), .A2(n6331), .ZN(n6533) );
  INV_X1 U8011 ( .A(n7805), .ZN(n6333) );
  NAND2_X1 U8012 ( .A1(n6533), .A2(n6333), .ZN(n6335) );
  NAND2_X1 U8013 ( .A1(n6557), .A2(n6551), .ZN(n6334) );
  NAND2_X1 U8014 ( .A1(n6335), .A2(n6334), .ZN(n6600) );
  INV_X1 U8015 ( .A(n6601), .ZN(n6336) );
  OAI211_X1 U8016 ( .C1(n6600), .C2(n6336), .A(n7881), .B(n7882), .ZN(n7670)
         );
  INV_X1 U8017 ( .A(n6651), .ZN(n7692) );
  NOR2_X1 U8018 ( .A1(n7810), .A2(n7692), .ZN(n6337) );
  NAND2_X1 U8019 ( .A1(n7670), .A2(n6337), .ZN(n6649) );
  NAND2_X1 U8020 ( .A1(n6649), .A2(n7883), .ZN(n6864) );
  NAND2_X1 U8021 ( .A1(n6962), .A2(n6740), .ZN(n6868) );
  AND2_X1 U8022 ( .A1(n7681), .A2(n6868), .ZN(n7683) );
  OR2_X1 U8023 ( .A1(n7697), .A2(n7683), .ZN(n6339) );
  AND2_X1 U8024 ( .A1(n7701), .A2(n7675), .ZN(n6338) );
  AND2_X1 U8025 ( .A1(n6339), .A2(n6338), .ZN(n7815) );
  NAND2_X1 U8026 ( .A1(n6864), .A2(n7815), .ZN(n7888) );
  AND2_X1 U8027 ( .A1(n7802), .A2(n7701), .ZN(n6340) );
  INV_X1 U8028 ( .A(n7709), .ZN(n6341) );
  NOR2_X1 U8029 ( .A1(n7225), .A2(n6341), .ZN(n6342) );
  NAND2_X1 U8030 ( .A1(n7330), .A2(n6342), .ZN(n7357) );
  NAND3_X1 U8031 ( .A1(n7820), .A2(n7357), .A3(n7893), .ZN(n6343) );
  OR2_X1 U8032 ( .A1(n9611), .A2(n7481), .ZN(n7725) );
  NAND2_X1 U8033 ( .A1(n9611), .A2(n7481), .ZN(n7722) );
  INV_X1 U8034 ( .A(n9499), .ZN(n8977) );
  OR2_X1 U8035 ( .A1(n9606), .A2(n8977), .ZN(n7726) );
  NAND2_X1 U8036 ( .A1(n9606), .A2(n8977), .ZN(n7728) );
  NAND2_X1 U8037 ( .A1(n7726), .A2(n7728), .ZN(n9520) );
  INV_X1 U8038 ( .A(n9489), .ZN(n9498) );
  NAND2_X1 U8039 ( .A1(n9497), .A2(n9498), .ZN(n9496) );
  NAND2_X1 U8040 ( .A1(n9496), .A2(n7732), .ZN(n9471) );
  AND2_X1 U8041 ( .A1(n9481), .A2(n9031), .ZN(n7734) );
  OR2_X1 U8042 ( .A1(n9481), .A2(n9031), .ZN(n7735) );
  INV_X1 U8043 ( .A(n9474), .ZN(n9042) );
  OR2_X1 U8044 ( .A1(n9592), .A2(n9042), .ZN(n7743) );
  NAND2_X1 U8045 ( .A1(n9592), .A2(n9042), .ZN(n7742) );
  NAND2_X1 U8046 ( .A1(n7743), .A2(n7742), .ZN(n7801) );
  INV_X1 U8047 ( .A(n9132), .ZN(n6344) );
  OR2_X1 U8048 ( .A1(n9587), .A2(n6344), .ZN(n7744) );
  NAND2_X1 U8049 ( .A1(n9587), .A2(n6344), .ZN(n7904) );
  NAND2_X1 U8050 ( .A1(n7744), .A2(n7904), .ZN(n9443) );
  XNOR2_X1 U8051 ( .A(n9582), .B(n9131), .ZN(n9430) );
  INV_X1 U8052 ( .A(n9131), .ZN(n7664) );
  OR2_X1 U8053 ( .A1(n9582), .A2(n7664), .ZN(n7745) );
  INV_X1 U8054 ( .A(n9407), .ZN(n9084) );
  XNOR2_X1 U8055 ( .A(n9422), .B(n9084), .ZN(n9414) );
  NAND2_X1 U8056 ( .A1(n9422), .A2(n9084), .ZN(n7749) );
  OR2_X1 U8057 ( .A1(n9571), .A2(n9381), .ZN(n7661) );
  NAND2_X1 U8058 ( .A1(n9571), .A2(n9381), .ZN(n7662) );
  NAND2_X1 U8059 ( .A1(n9404), .A2(n7662), .ZN(n9378) );
  INV_X1 U8060 ( .A(n9408), .ZN(n6346) );
  OR2_X1 U8061 ( .A1(n9388), .A2(n6346), .ZN(n7751) );
  NAND2_X1 U8062 ( .A1(n9388), .A2(n6346), .ZN(n9362) );
  INV_X1 U8063 ( .A(n9339), .ZN(n6347) );
  OR2_X1 U8064 ( .A1(n9355), .A2(n6347), .ZN(n7761) );
  NAND2_X1 U8065 ( .A1(n9355), .A2(n6347), .ZN(n7760) );
  NAND2_X1 U8066 ( .A1(n7761), .A2(n7760), .ZN(n9346) );
  INV_X1 U8067 ( .A(n9330), .ZN(n9338) );
  NAND2_X1 U8068 ( .A1(n9312), .A2(n9313), .ZN(n9311) );
  INV_X1 U8069 ( .A(n7778), .ZN(n7831) );
  OR2_X1 U8070 ( .A1(n7795), .A2(n7866), .ZN(n6348) );
  NAND2_X1 U8071 ( .A1(n4976), .A2(n7870), .ZN(n7796) );
  INV_X1 U8072 ( .A(n9691), .ZN(n9738) );
  NAND2_X1 U8073 ( .A1(n9738), .A2(P1_B_REG_SCAN_IN), .ZN(n6349) );
  AND2_X1 U8074 ( .A1(n9500), .A2(n6349), .ZN(n7946) );
  INV_X1 U8075 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U8076 ( .A1(n7651), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U8077 ( .A1(n5073), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6350) );
  OAI211_X1 U8078 ( .C1(n7655), .C2(n6352), .A(n6351), .B(n6350), .ZN(n9126)
         );
  AOI22_X1 U8079 ( .A1(n9127), .A2(n9524), .B1(n7946), .B2(n9126), .ZN(n6353)
         );
  NAND2_X1 U8080 ( .A1(n6357), .A2(n6356), .ZN(n6361) );
  NOR2_X1 U8081 ( .A1(n7936), .A2(n6358), .ZN(n6359) );
  NAND2_X1 U8082 ( .A1(n6360), .A2(n6359), .ZN(n6610) );
  OR2_X1 U8083 ( .A1(n9876), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8084 ( .A1(n6364), .A2(n6363), .ZN(n6366) );
  NAND2_X1 U8085 ( .A1(n9284), .A2(n6606), .ZN(n6365) );
  NAND2_X1 U8086 ( .A1(n6366), .A2(n6365), .ZN(P1_U3551) );
  INV_X1 U8087 ( .A(n6367), .ZN(n6613) );
  OR2_X1 U8088 ( .A1(n9871), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U8089 ( .A1(n9284), .A2(n6572), .ZN(n6371) );
  NOR2_X1 U8090 ( .A1(n5046), .A2(P1_U3086), .ZN(n6372) );
  XNOR2_X1 U8091 ( .A(n7503), .B(n7504), .ZN(n6376) );
  INV_X1 U8092 ( .A(n6374), .ZN(n6375) );
  NOR2_X1 U8093 ( .A1(n6376), .A2(n6375), .ZN(n7502) );
  AOI21_X1 U8094 ( .B1(n6376), .B2(n6375), .A(n7502), .ZN(n6377) );
  NOR2_X1 U8095 ( .A1(n6377), .A2(n9098), .ZN(n6383) );
  AND2_X1 U8096 ( .A1(n9096), .A2(n7127), .ZN(n6382) );
  INV_X1 U8097 ( .A(n7122), .ZN(n6378) );
  AND2_X1 U8098 ( .A1(n9121), .A2(n6378), .ZN(n6381) );
  OR2_X1 U8099 ( .A1(n9083), .A2(n7306), .ZN(n6379) );
  NAND2_X1 U8100 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6467) );
  OAI211_X1 U8101 ( .C1(n9119), .C2(n7411), .A(n6379), .B(n6467), .ZN(n6380)
         );
  OR4_X1 U8102 ( .A1(n6383), .A2(n6382), .A3(n6381), .A4(n6380), .ZN(P1_U3217)
         );
  INV_X1 U8103 ( .A(n6932), .ZN(n7586) );
  NAND2_X1 U8104 ( .A1(n8432), .A2(n6932), .ZN(n6384) );
  NAND2_X1 U8105 ( .A1(n6671), .A2(n6384), .ZN(n6685) );
  OR2_X1 U8106 ( .A1(n6685), .A2(n6385), .ZN(n6386) );
  NAND2_X1 U8107 ( .A1(n6386), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X2 U8108 ( .A(n8958), .ZN(n7957) );
  OAI222_X1 U8109 ( .A1(n7957), .A2(n6387), .B1(n8960), .B2(n6397), .C1(
        P2_U3151), .C2(n6732), .ZN(P2_U3294) );
  INV_X2 U8110 ( .A(n7582), .ZN(n9688) );
  OAI222_X1 U8111 ( .A1(n9694), .A2(n4497), .B1(n9688), .B2(n6394), .C1(
        P1_U3086), .C2(n6445), .ZN(P1_U3353) );
  OAI222_X1 U8112 ( .A1(n9694), .A2(n6390), .B1(n9688), .B2(n6395), .C1(
        P1_U3086), .C2(n6451), .ZN(P1_U3352) );
  OAI222_X1 U8113 ( .A1(n9694), .A2(n6391), .B1(n9688), .B2(n6392), .C1(
        P1_U3086), .C2(n9188), .ZN(P1_U3351) );
  INV_X1 U8114 ( .A(n8960), .ZN(n8969) );
  INV_X1 U8115 ( .A(n8969), .ZN(n8964) );
  OAI222_X1 U8116 ( .A1(n7957), .A2(n6393), .B1(n8964), .B2(n6392), .C1(
        P2_U3151), .C2(n6695), .ZN(P2_U3291) );
  OAI222_X1 U8117 ( .A1(n7957), .A2(n5828), .B1(n8964), .B2(n6394), .C1(
        P2_U3151), .C2(n4354), .ZN(P2_U3293) );
  OAI222_X1 U8118 ( .A1(n7957), .A2(n5006), .B1(n8964), .B2(n6395), .C1(
        P2_U3151), .C2(n6691), .ZN(P2_U3292) );
  OAI222_X1 U8119 ( .A1(n7957), .A2(n6396), .B1(n8964), .B2(n6399), .C1(
        P2_U3151), .C2(n6812), .ZN(P2_U3290) );
  OAI222_X1 U8120 ( .A1(n9694), .A2(n6398), .B1(n9688), .B2(n6397), .C1(
        P1_U3086), .C2(n6447), .ZN(P1_U3354) );
  OAI222_X1 U8121 ( .A1(n9694), .A2(n6400), .B1(n9688), .B2(n6399), .C1(
        P1_U3086), .C2(n9201), .ZN(P1_U3350) );
  INV_X1 U8122 ( .A(n9694), .ZN(n7155) );
  AOI22_X1 U8123 ( .A1(n7155), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9218), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6401) );
  OAI21_X1 U8124 ( .B1(n6402), .B2(n9688), .A(n6401), .ZN(P1_U3349) );
  OAI222_X1 U8125 ( .A1(n7957), .A2(n6403), .B1(n8964), .B2(n6402), .C1(
        P2_U3151), .C2(n6894), .ZN(P2_U3289) );
  AOI22_X1 U8126 ( .A1(n9231), .A2(P1_STATE_REG_SCAN_IN), .B1(n7155), .B2(
        P2_DATAO_REG_7__SCAN_IN), .ZN(n6404) );
  OAI21_X1 U8127 ( .B1(n6405), .B2(n9688), .A(n6404), .ZN(P1_U3348) );
  OAI222_X1 U8128 ( .A1(n7957), .A2(n6406), .B1(n8964), .B2(n6405), .C1(
        P2_U3151), .C2(n7000), .ZN(P2_U3288) );
  NAND2_X1 U8129 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  AND2_X1 U8130 ( .A1(n6409), .A2(n5026), .ZN(n6440) );
  INV_X1 U8131 ( .A(n6440), .ZN(n6410) );
  NAND2_X1 U8132 ( .A1(n7936), .A2(n7931), .ZN(n6441) );
  AND2_X1 U8133 ( .A1(n6410), .A2(n6441), .ZN(n9746) );
  NOR2_X1 U8134 ( .A1(n9746), .A2(P1_U3973), .ZN(P1_U3085) );
  AOI22_X1 U8135 ( .A1(n9244), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7155), .ZN(n6411) );
  OAI21_X1 U8136 ( .B1(n6412), .B2(n9688), .A(n6411), .ZN(P1_U3347) );
  OAI222_X1 U8137 ( .A1(n7957), .A2(n6413), .B1(n8964), .B2(n6412), .C1(
        P2_U3151), .C2(n7102), .ZN(P2_U3287) );
  INV_X1 U8138 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8139 ( .A1(n6540), .A2(P1_U3973), .ZN(n6414) );
  OAI21_X1 U8140 ( .B1(P1_U3973), .B2(n6415), .A(n6414), .ZN(P1_U3554) );
  INV_X1 U8141 ( .A(n6416), .ZN(n6418) );
  INV_X1 U8142 ( .A(n7936), .ZN(n6417) );
  NAND2_X1 U8143 ( .A1(n9847), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6419) );
  OAI21_X1 U8144 ( .B1(n9847), .B2(n6420), .A(n6419), .ZN(P1_U3439) );
  INV_X1 U8145 ( .A(n6421), .ZN(n6424) );
  AOI22_X1 U8146 ( .A1(n6484), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n7155), .ZN(n6422) );
  OAI21_X1 U8147 ( .B1(n6424), .B2(n9688), .A(n6422), .ZN(P1_U3346) );
  INV_X1 U8148 ( .A(n7175), .ZN(n7190) );
  OAI222_X1 U8149 ( .A1(n8964), .A2(n6424), .B1(n7190), .B2(P2_U3151), .C1(
        n6423), .C2(n7957), .ZN(P2_U3286) );
  INV_X1 U8150 ( .A(n6425), .ZN(n6428) );
  AOI22_X1 U8151 ( .A1(n6500), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7155), .ZN(n6426) );
  OAI21_X1 U8152 ( .B1(n6428), .B2(n9688), .A(n6426), .ZN(P1_U3345) );
  INV_X1 U8153 ( .A(n7196), .ZN(n7256) );
  INV_X1 U8154 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6427) );
  OAI222_X1 U8155 ( .A1(n8964), .A2(n6428), .B1(n7256), .B2(P2_U3151), .C1(
        n6427), .C2(n7957), .ZN(P2_U3285) );
  XNOR2_X1 U8156 ( .A(n6500), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6444) );
  INV_X1 U8157 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6627) );
  MUX2_X1 U8158 ( .A(n6627), .B(P1_REG2_REG_2__SCAN_IN), .S(n6445), .Z(n9171)
         );
  MUX2_X1 U8159 ( .A(n5018), .B(P1_REG2_REG_1__SCAN_IN), .S(n6447), .Z(n9147)
         );
  NAND2_X1 U8160 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9159) );
  INV_X1 U8161 ( .A(n9159), .ZN(n9146) );
  NAND2_X1 U8162 ( .A1(n9147), .A2(n9146), .ZN(n9145) );
  INV_X1 U8163 ( .A(n6447), .ZN(n9151) );
  NAND2_X1 U8164 ( .A1(n9151), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U8165 ( .A1(n9145), .A2(n6429), .ZN(n9170) );
  NAND2_X1 U8166 ( .A1(n9171), .A2(n9170), .ZN(n9169) );
  INV_X1 U8167 ( .A(n6445), .ZN(n9165) );
  NAND2_X1 U8168 ( .A1(n9165), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U8169 ( .A1(n9169), .A2(n6430), .ZN(n9183) );
  XNOR2_X1 U8170 ( .A(n6451), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9184) );
  NAND2_X1 U8171 ( .A1(n9183), .A2(n9184), .ZN(n9182) );
  INV_X1 U8172 ( .A(n6451), .ZN(n9178) );
  NAND2_X1 U8173 ( .A1(n9178), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U8174 ( .A1(n9182), .A2(n6431), .ZN(n9192) );
  MUX2_X1 U8175 ( .A(n6618), .B(P1_REG2_REG_4__SCAN_IN), .S(n9188), .Z(n9193)
         );
  NAND2_X1 U8176 ( .A1(n9192), .A2(n9193), .ZN(n9191) );
  INV_X1 U8177 ( .A(n9188), .ZN(n6453) );
  NAND2_X1 U8178 ( .A1(n6453), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U8179 ( .A1(n9191), .A2(n6432), .ZN(n9210) );
  XNOR2_X1 U8180 ( .A(n9201), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U8181 ( .A1(n9210), .A2(n9211), .ZN(n9209) );
  OR2_X1 U8182 ( .A1(n9201), .A2(n6433), .ZN(n6434) );
  NAND2_X1 U8183 ( .A1(n9209), .A2(n6434), .ZN(n9223) );
  XNOR2_X1 U8184 ( .A(n9218), .B(n6435), .ZN(n9224) );
  NAND2_X1 U8185 ( .A1(n9223), .A2(n9224), .ZN(n9222) );
  NAND2_X1 U8186 ( .A1(n9218), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U8187 ( .A1(n9222), .A2(n6436), .ZN(n9233) );
  MUX2_X1 U8188 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6957), .S(n9231), .Z(n9234)
         );
  NAND2_X1 U8189 ( .A1(n9233), .A2(n9234), .ZN(n9232) );
  NAND2_X1 U8190 ( .A1(n9231), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8191 ( .A1(n9232), .A2(n6437), .ZN(n9246) );
  XNOR2_X1 U8192 ( .A(n9244), .B(n6873), .ZN(n9247) );
  NAND2_X1 U8193 ( .A1(n9246), .A2(n9247), .ZN(n9245) );
  NAND2_X1 U8194 ( .A1(n9244), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U8195 ( .A1(n9245), .A2(n6438), .ZN(n6475) );
  XNOR2_X1 U8196 ( .A(n6484), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6476) );
  OR2_X1 U8197 ( .A1(n6475), .A2(n6476), .ZN(n6473) );
  OR2_X1 U8198 ( .A1(n6484), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8199 ( .A1(n6473), .A2(n6439), .ZN(n6443) );
  NAND2_X1 U8200 ( .A1(n6441), .A2(n6440), .ZN(n9749) );
  OR2_X1 U8201 ( .A1(n4352), .A2(n9691), .ZN(n9158) );
  OR2_X1 U8202 ( .A1(n6443), .A2(n6444), .ZN(n6495) );
  INV_X1 U8203 ( .A(n6495), .ZN(n6442) );
  AOI211_X1 U8204 ( .C1(n6444), .C2(n6443), .A(n9798), .B(n6442), .ZN(n6472)
         );
  XNOR2_X1 U8205 ( .A(n6500), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n6465) );
  INV_X1 U8206 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6446) );
  MUX2_X1 U8207 ( .A(n6446), .B(P1_REG1_REG_2__SCAN_IN), .S(n6445), .Z(n9168)
         );
  INV_X1 U8208 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6448) );
  MUX2_X1 U8209 ( .A(n6448), .B(P1_REG1_REG_1__SCAN_IN), .S(n6447), .Z(n9150)
         );
  AND2_X1 U8210 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9149) );
  NAND2_X1 U8211 ( .A1(n9150), .A2(n9149), .ZN(n9148) );
  NAND2_X1 U8212 ( .A1(n9151), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U8213 ( .A1(n9148), .A2(n6449), .ZN(n9167) );
  NAND2_X1 U8214 ( .A1(n9168), .A2(n9167), .ZN(n9166) );
  NAND2_X1 U8215 ( .A1(n9165), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8216 ( .A1(n9166), .A2(n6450), .ZN(n9180) );
  XNOR2_X1 U8217 ( .A(n6451), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9181) );
  NAND2_X1 U8218 ( .A1(n9180), .A2(n9181), .ZN(n9179) );
  NAND2_X1 U8219 ( .A1(n9178), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6452) );
  NAND2_X1 U8220 ( .A1(n9179), .A2(n6452), .ZN(n9195) );
  MUX2_X1 U8221 ( .A(n4943), .B(P1_REG1_REG_4__SCAN_IN), .S(n9188), .Z(n9196)
         );
  NAND2_X1 U8222 ( .A1(n9195), .A2(n9196), .ZN(n9194) );
  NAND2_X1 U8223 ( .A1(n6453), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U8224 ( .A1(n9194), .A2(n6454), .ZN(n9207) );
  XNOR2_X1 U8225 ( .A(n9201), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9208) );
  NAND2_X1 U8226 ( .A1(n9207), .A2(n9208), .ZN(n9206) );
  OR2_X1 U8227 ( .A1(n9201), .A2(n6455), .ZN(n6456) );
  NAND2_X1 U8228 ( .A1(n9206), .A2(n6456), .ZN(n9220) );
  XNOR2_X1 U8229 ( .A(n9218), .B(n6457), .ZN(n9221) );
  NAND2_X1 U8230 ( .A1(n9220), .A2(n9221), .ZN(n9219) );
  NAND2_X1 U8231 ( .A1(n9218), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8232 ( .A1(n9219), .A2(n6458), .ZN(n9236) );
  MUX2_X1 U8233 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n5145), .S(n9231), .Z(n9237)
         );
  NAND2_X1 U8234 ( .A1(n9236), .A2(n9237), .ZN(n9235) );
  NAND2_X1 U8235 ( .A1(n9231), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U8236 ( .A1(n9235), .A2(n6459), .ZN(n9249) );
  XNOR2_X1 U8237 ( .A(n9244), .B(n6460), .ZN(n9250) );
  NAND2_X1 U8238 ( .A1(n9249), .A2(n9250), .ZN(n9248) );
  NAND2_X1 U8239 ( .A1(n9244), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U8240 ( .A1(n9248), .A2(n6461), .ZN(n6478) );
  XNOR2_X1 U8241 ( .A(n6484), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n6477) );
  OR2_X1 U8242 ( .A1(n6478), .A2(n6477), .ZN(n6480) );
  OR2_X1 U8243 ( .A1(n6484), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8244 ( .A1(n6480), .A2(n6462), .ZN(n6464) );
  OR2_X1 U8245 ( .A1(n6464), .A2(n6465), .ZN(n6502) );
  INV_X1 U8246 ( .A(n6502), .ZN(n6463) );
  AOI211_X1 U8247 ( .C1(n6465), .C2(n6464), .A(n9808), .B(n6463), .ZN(n6471)
         );
  INV_X1 U8248 ( .A(n6500), .ZN(n6469) );
  NAND2_X1 U8249 ( .A1(n9746), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n6468) );
  OAI211_X1 U8250 ( .C1(n9790), .C2(n6469), .A(n6468), .B(n6467), .ZN(n6470)
         );
  OR3_X1 U8251 ( .A1(n6472), .A2(n6471), .A3(n6470), .ZN(P1_U3253) );
  INV_X1 U8252 ( .A(n6473), .ZN(n6474) );
  AOI21_X1 U8253 ( .B1(n6476), .B2(n6475), .A(n6474), .ZN(n6486) );
  NAND2_X1 U8254 ( .A1(n6478), .A2(n6477), .ZN(n6479) );
  AOI21_X1 U8255 ( .B1(n6480), .B2(n6479), .A(n9808), .ZN(n6483) );
  INV_X1 U8256 ( .A(n9746), .ZN(n9823) );
  INV_X1 U8257 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U8258 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7379) );
  OAI21_X1 U8259 ( .B1(n9823), .B2(n6481), .A(n7379), .ZN(n6482) );
  AOI211_X1 U8260 ( .C1(n9811), .C2(n6484), .A(n6483), .B(n6482), .ZN(n6485)
         );
  OAI21_X1 U8261 ( .B1(n6486), .B2(n9798), .A(n6485), .ZN(P1_U3252) );
  INV_X1 U8262 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6490) );
  AND2_X1 U8263 ( .A1(n6540), .A2(n6546), .ZN(n7876) );
  OR2_X1 U8264 ( .A1(n7876), .A2(n6538), .ZN(n7803) );
  OAI21_X1 U8265 ( .B1(n9503), .B2(n9869), .A(n7803), .ZN(n6488) );
  NAND2_X1 U8266 ( .A1(n6487), .A2(n9500), .ZN(n6637) );
  OAI211_X1 U8267 ( .C1(n6636), .C2(n6546), .A(n6488), .B(n6637), .ZN(n9634)
         );
  NAND2_X1 U8268 ( .A1(n9634), .A2(n9871), .ZN(n6489) );
  OAI21_X1 U8269 ( .B1(n9871), .B2(n6490), .A(n6489), .ZN(P1_U3453) );
  INV_X1 U8270 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U8271 ( .A1(n6491), .A2(n6517), .ZN(n6492) );
  OAI21_X1 U8272 ( .B1(n6517), .B2(n6493), .A(n6492), .ZN(P2_U3377) );
  INV_X1 U8273 ( .A(n7162), .ZN(n6519) );
  AOI22_X1 U8274 ( .A1(n7162), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7222), .B2(
        n6519), .ZN(n6499) );
  NAND2_X1 U8275 ( .A1(n6500), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U8276 ( .A1(n6495), .A2(n6494), .ZN(n9751) );
  OR2_X1 U8277 ( .A1(n6514), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U8278 ( .A1(n6514), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6496) );
  AND2_X1 U8279 ( .A1(n6497), .A2(n6496), .ZN(n9750) );
  AND2_X1 U8280 ( .A1(n9751), .A2(n9750), .ZN(n9753) );
  AOI21_X1 U8281 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6514), .A(n9753), .ZN(
        n6498) );
  NAND2_X1 U8282 ( .A1(n6499), .A2(n6498), .ZN(n7161) );
  OAI21_X1 U8283 ( .B1(n6499), .B2(n6498), .A(n7161), .ZN(n6510) );
  NAND2_X1 U8284 ( .A1(n6500), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6501) );
  NAND2_X1 U8285 ( .A1(n6502), .A2(n6501), .ZN(n9755) );
  XNOR2_X1 U8286 ( .A(n6514), .B(n9631), .ZN(n9754) );
  AND2_X1 U8287 ( .A1(n9755), .A2(n9754), .ZN(n9757) );
  AOI21_X1 U8288 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6514), .A(n9757), .ZN(
        n6505) );
  AOI22_X1 U8289 ( .A1(n7162), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n6503), .B2(
        n6519), .ZN(n6504) );
  NAND2_X1 U8290 ( .A1(n6505), .A2(n6504), .ZN(n7157) );
  OAI21_X1 U8291 ( .B1(n6505), .B2(n6504), .A(n7157), .ZN(n6506) );
  NAND2_X1 U8292 ( .A1(n6506), .A2(n9786), .ZN(n6508) );
  AND2_X1 U8293 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7409) );
  AOI21_X1 U8294 ( .B1(n9746), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7409), .ZN(
        n6507) );
  OAI211_X1 U8295 ( .C1(n9790), .C2(n6519), .A(n6508), .B(n6507), .ZN(n6509)
         );
  AOI21_X1 U8296 ( .B1(n9815), .B2(n6510), .A(n6509), .ZN(n6511) );
  INV_X1 U8297 ( .A(n6511), .ZN(P1_U3255) );
  INV_X1 U8298 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6513) );
  INV_X1 U8299 ( .A(n6512), .ZN(n6515) );
  INV_X1 U8300 ( .A(n7426), .ZN(n7433) );
  OAI222_X1 U8301 ( .A1(n7957), .A2(n6513), .B1(n8960), .B2(n6515), .C1(
        P2_U3151), .C2(n7433), .ZN(P2_U3284) );
  INV_X1 U8302 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6516) );
  INV_X1 U8303 ( .A(n6514), .ZN(n9760) );
  OAI222_X1 U8304 ( .A1(n9694), .A2(n6516), .B1(n9688), .B2(n6515), .C1(
        P1_U3086), .C2(n9760), .ZN(P1_U3344) );
  AND2_X1 U8305 ( .A1(n6577), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8306 ( .A1(n6577), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8307 ( .A1(n6577), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8308 ( .A1(n6577), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8309 ( .A1(n6577), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8310 ( .A1(n6577), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8311 ( .A1(n6577), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8312 ( .A1(n6577), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8313 ( .A1(n6577), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8314 ( .A1(n6577), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8315 ( .A1(n6577), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  INV_X1 U8316 ( .A(n8483), .ZN(n7443) );
  INV_X1 U8317 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6518) );
  OAI222_X1 U8318 ( .A1(n8960), .A2(n6520), .B1(n7443), .B2(P2_U3151), .C1(
        n6518), .C2(n7957), .ZN(P2_U3283) );
  INV_X1 U8319 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6521) );
  OAI222_X1 U8320 ( .A1(n9694), .A2(n6521), .B1(n9688), .B2(n6520), .C1(n6519), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8321 ( .A(n9119), .ZN(n9109) );
  AOI22_X1 U8322 ( .A1(n9109), .A2(n6487), .B1(n9096), .B2(n6635), .ZN(n6528)
         );
  NOR2_X1 U8323 ( .A1(n6523), .A2(n6522), .ZN(n6524) );
  NOR2_X1 U8324 ( .A1(n6525), .A2(n6524), .ZN(n9156) );
  OR2_X1 U8325 ( .A1(n6526), .A2(n7936), .ZN(n7964) );
  AOI22_X1 U8326 ( .A1(n9156), .A2(n9115), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n7964), .ZN(n6527) );
  NAND2_X1 U8327 ( .A1(n6528), .A2(n6527), .ZN(P1_U3232) );
  AOI22_X1 U8328 ( .A1(n9773), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7155), .ZN(n6530) );
  OAI21_X1 U8329 ( .B1(n6529), .B2(n9688), .A(n6530), .ZN(P1_U3342) );
  OAI21_X1 U8330 ( .B1(n6532), .B2(n7805), .A(n6531), .ZN(n6626) );
  AOI211_X1 U8331 ( .C1(n6551), .C2(n6545), .A(n9510), .B(n6567), .ZN(n6630)
         );
  XNOR2_X1 U8332 ( .A(n6533), .B(n7805), .ZN(n6534) );
  OAI222_X1 U8333 ( .A1(n9516), .A2(n6536), .B1(n9380), .B2(n6535), .C1(n9518), 
        .C2(n6534), .ZN(n6631) );
  AOI211_X1 U8334 ( .C1(n9869), .C2(n6626), .A(n6630), .B(n6631), .ZN(n6576)
         );
  AOI22_X1 U8335 ( .A1(n6606), .A2(n6551), .B1(n6362), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6537) );
  OAI21_X1 U8336 ( .B1(n6576), .B2(n6362), .A(n6537), .ZN(P1_U3524) );
  XNOR2_X1 U8337 ( .A(n6539), .B(n6538), .ZN(n6542) );
  INV_X1 U8338 ( .A(n6540), .ZN(n6541) );
  OAI22_X1 U8339 ( .A1(n6557), .A2(n9516), .B1(n6541), .B2(n9380), .ZN(n7965)
         );
  AOI21_X1 U8340 ( .B1(n6542), .B2(n9503), .A(n7965), .ZN(n9846) );
  NAND2_X1 U8341 ( .A1(n9835), .A2(n9869), .ZN(n6547) );
  OAI211_X1 U8342 ( .C1(n6546), .C2(n6328), .A(n9531), .B(n6545), .ZN(n9842)
         );
  AND3_X1 U8343 ( .A1(n9846), .A2(n6547), .A3(n9842), .ZN(n6585) );
  AOI22_X1 U8344 ( .A1(n6606), .A2(n9837), .B1(n6362), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n6548) );
  OAI21_X1 U8345 ( .B1(n6585), .B2(n6362), .A(n6548), .ZN(P1_U3523) );
  XOR2_X1 U8346 ( .A(n6550), .B(n6549), .Z(n6554) );
  AOI22_X1 U8347 ( .A1(n9096), .A2(n6551), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n7964), .ZN(n6553) );
  INV_X1 U8348 ( .A(n9083), .ZN(n9117) );
  AOI22_X1 U8349 ( .A1(n9117), .A2(n6487), .B1(n9109), .B2(n9142), .ZN(n6552)
         );
  OAI211_X1 U8350 ( .C1(n6554), .C2(n9098), .A(n6553), .B(n6552), .ZN(P1_U3237) );
  XOR2_X1 U8351 ( .A(n6556), .B(n6555), .Z(n6560) );
  OAI22_X1 U8352 ( .A1(n6557), .A2(n9380), .B1(n6290), .B2(n9516), .ZN(n6565)
         );
  AOI22_X1 U8353 ( .A1(n9096), .A2(n9824), .B1(n9060), .B2(n6565), .ZN(n6559)
         );
  MUX2_X1 U8354 ( .A(P1_STATE_REG_SCAN_IN), .B(n9107), .S(n9825), .Z(n6558) );
  OAI211_X1 U8355 ( .C1(n6560), .C2(n9098), .A(n6559), .B(n6558), .ZN(P1_U3218) );
  INV_X1 U8356 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6561) );
  OAI222_X1 U8357 ( .A1(n8960), .A2(n6529), .B1(n8509), .B2(P2_U3151), .C1(
        n6561), .C2(n7957), .ZN(P2_U3282) );
  OAI21_X1 U8358 ( .B1(n6563), .B2(n6564), .A(n6562), .ZN(n9831) );
  INV_X1 U8359 ( .A(n9831), .ZN(n6568) );
  INV_X1 U8360 ( .A(n6564), .ZN(n7806) );
  XNOR2_X1 U8361 ( .A(n6600), .B(n7806), .ZN(n6566) );
  AOI21_X1 U8362 ( .B1(n6566), .B2(n9503), .A(n6565), .ZN(n9833) );
  OAI211_X1 U8363 ( .C1(n6567), .C2(n6587), .A(n6599), .B(n9531), .ZN(n9829)
         );
  OAI211_X1 U8364 ( .C1(n6568), .C2(n9625), .A(n9833), .B(n9829), .ZN(n6589)
         );
  INV_X1 U8365 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6569) );
  OAI22_X1 U8366 ( .A1(n9633), .A2(n6587), .B1(n9876), .B2(n6569), .ZN(n6570)
         );
  AOI21_X1 U8367 ( .B1(n6589), .B2(n9876), .A(n6570), .ZN(n6571) );
  INV_X1 U8368 ( .A(n6571), .ZN(P1_U3525) );
  INV_X1 U8369 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6573) );
  OAI22_X1 U8370 ( .A1(n9676), .A2(n7877), .B1(n9871), .B2(n6573), .ZN(n6574)
         );
  INV_X1 U8371 ( .A(n6574), .ZN(n6575) );
  OAI21_X1 U8372 ( .B1(n6576), .B2(n6369), .A(n6575), .ZN(P1_U3459) );
  INV_X1 U8373 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6581) );
  INV_X1 U8374 ( .A(n6578), .ZN(n6579) );
  AOI22_X1 U8375 ( .A1(n6577), .A2(n6581), .B1(n6580), .B2(n6579), .ZN(
        P2_U3376) );
  INV_X1 U8376 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6582) );
  OAI22_X1 U8377 ( .A1(n9676), .A2(n6328), .B1(n9871), .B2(n6582), .ZN(n6583)
         );
  INV_X1 U8378 ( .A(n6583), .ZN(n6584) );
  OAI21_X1 U8379 ( .B1(n6585), .B2(n6369), .A(n6584), .ZN(P1_U3456) );
  INV_X1 U8380 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6586) );
  OAI22_X1 U8381 ( .A1(n9676), .A2(n6587), .B1(n9871), .B2(n6586), .ZN(n6588)
         );
  AOI21_X1 U8382 ( .B1(n6589), .B2(n9871), .A(n6588), .ZN(n6590) );
  INV_X1 U8383 ( .A(n6590), .ZN(P1_U3462) );
  INV_X1 U8384 ( .A(n6591), .ZN(n6643) );
  AOI22_X1 U8385 ( .A1(n9777), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7155), .ZN(n6592) );
  OAI21_X1 U8386 ( .B1(n6643), .B2(n9688), .A(n6592), .ZN(P1_U3341) );
  INV_X1 U8387 ( .A(n7021), .ZN(n6945) );
  NAND2_X1 U8388 ( .A1(n8466), .A2(n6945), .ZN(n8274) );
  NAND2_X1 U8389 ( .A1(n8274), .A2(n8270), .ZN(n8246) );
  OR2_X1 U8390 ( .A1(n9933), .A2(n8817), .ZN(n6593) );
  NAND2_X1 U8391 ( .A1(n8246), .A2(n6593), .ZN(n6594) );
  NAND2_X1 U8392 ( .A1(n5819), .A2(n8819), .ZN(n6979) );
  OAI211_X1 U8393 ( .C1(n6945), .C2(n9925), .A(n6594), .B(n6979), .ZN(n6965)
         );
  NAND2_X1 U8394 ( .A1(n9950), .A2(n6965), .ZN(n6595) );
  OAI21_X1 U8395 ( .B1(n9950), .B2(n6662), .A(n6595), .ZN(P2_U3459) );
  OAI21_X1 U8396 ( .B1(n6597), .B2(n7804), .A(n6596), .ZN(n6609) );
  INV_X1 U8397 ( .A(n6647), .ZN(n6598) );
  AOI211_X1 U8398 ( .C1(n9063), .C2(n6599), .A(n9510), .B(n6598), .ZN(n6622)
         );
  NAND2_X1 U8399 ( .A1(n6600), .A2(n7882), .ZN(n6602) );
  NAND2_X1 U8400 ( .A1(n6602), .A2(n6601), .ZN(n7671) );
  XNOR2_X1 U8401 ( .A(n7671), .B(n7804), .ZN(n6603) );
  AOI22_X1 U8402 ( .A1(n9140), .A2(n9500), .B1(n9524), .B2(n9142), .ZN(n9058)
         );
  OAI21_X1 U8403 ( .B1(n6603), .B2(n9518), .A(n9058), .ZN(n6616) );
  AOI211_X1 U8404 ( .C1(n9869), .C2(n6609), .A(n6622), .B(n6616), .ZN(n6608)
         );
  OAI22_X1 U8405 ( .A1(n9676), .A2(n6620), .B1(n9871), .B2(n4949), .ZN(n6604)
         );
  INV_X1 U8406 ( .A(n6604), .ZN(n6605) );
  OAI21_X1 U8407 ( .B1(n6608), .B2(n6369), .A(n6605), .ZN(P1_U3465) );
  AOI22_X1 U8408 ( .A1(n6606), .A2(n9063), .B1(n6362), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6607) );
  OAI21_X1 U8409 ( .B1(n6608), .B2(n6362), .A(n6607), .ZN(P1_U3526) );
  AND2_X1 U8410 ( .A1(n6577), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8411 ( .A1(n6577), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8412 ( .A1(n6577), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8413 ( .A1(n6577), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8414 ( .A1(n6577), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8415 ( .A1(n6577), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8416 ( .A1(n6577), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8417 ( .A1(n6577), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8418 ( .A1(n6577), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8419 ( .A1(n6577), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8420 ( .A1(n6577), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8421 ( .A1(n6577), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8422 ( .A1(n6577), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8423 ( .A1(n6577), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8424 ( .A1(n6577), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8425 ( .A1(n6577), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8426 ( .A1(n6577), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8427 ( .A1(n6577), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8428 ( .A1(n6577), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8429 ( .A(n6609), .ZN(n6625) );
  INV_X1 U8430 ( .A(n6610), .ZN(n6612) );
  NAND3_X1 U8431 ( .A1(n6613), .A2(n6612), .A3(n6611), .ZN(n6614) );
  AND2_X1 U8432 ( .A1(n7332), .A2(n6946), .ZN(n6615) );
  INV_X1 U8433 ( .A(n6616), .ZN(n6617) );
  MUX2_X1 U8434 ( .A(n6618), .B(n6617), .S(n9468), .Z(n6624) );
  OAI22_X1 U8435 ( .A1(n9514), .A2(n6620), .B1(n9061), .B2(n9390), .ZN(n6621)
         );
  AOI21_X1 U8436 ( .B1(n6622), .B2(n9527), .A(n6621), .ZN(n6623) );
  OAI211_X1 U8437 ( .C1(n6625), .C2(n9529), .A(n6624), .B(n6623), .ZN(P1_U3289) );
  INV_X1 U8438 ( .A(n6626), .ZN(n6634) );
  NOR2_X1 U8439 ( .A1(n9514), .A2(n7877), .ZN(n6629) );
  INV_X1 U8440 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9162) );
  OAI22_X1 U8441 ( .A1(n9468), .A2(n6627), .B1(n9162), .B2(n9390), .ZN(n6628)
         );
  AOI211_X1 U8442 ( .C1(n6630), .C2(n9527), .A(n6629), .B(n6628), .ZN(n6633)
         );
  NAND2_X1 U8443 ( .A1(n6631), .A2(n9468), .ZN(n6632) );
  OAI211_X1 U8444 ( .C1(n6634), .C2(n9529), .A(n6633), .B(n6632), .ZN(P1_U3291) );
  INV_X1 U8445 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6642) );
  NOR2_X1 U8446 ( .A1(n9841), .A2(n9510), .ZN(n9276) );
  OAI21_X1 U8447 ( .B1(n9276), .B2(n9838), .A(n6635), .ZN(n6641) );
  NAND3_X1 U8448 ( .A1(n7803), .A2(n7935), .A3(n6636), .ZN(n6638) );
  OAI211_X1 U8449 ( .C1(n5036), .C2(n9390), .A(n6638), .B(n6637), .ZN(n6639)
         );
  NAND2_X1 U8450 ( .A1(n6639), .A2(n9468), .ZN(n6640) );
  OAI211_X1 U8451 ( .C1(n9468), .C2(n6642), .A(n6641), .B(n6640), .ZN(P1_U3293) );
  INV_X1 U8452 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6644) );
  OAI222_X1 U8453 ( .A1(n7957), .A2(n6644), .B1(n8960), .B2(n6643), .C1(
        P2_U3151), .C2(n8529), .ZN(P2_U3281) );
  OAI21_X1 U8454 ( .B1(n6646), .B2(n7810), .A(n6645), .ZN(n6754) );
  AOI211_X1 U8455 ( .C1(n6648), .C2(n6647), .A(n9510), .B(n6746), .ZN(n6755)
         );
  NAND2_X1 U8456 ( .A1(n6649), .A2(n9503), .ZN(n6654) );
  INV_X1 U8457 ( .A(n7810), .ZN(n6650) );
  AOI21_X1 U8458 ( .B1(n7670), .B2(n6651), .A(n6650), .ZN(n6653) );
  AOI22_X1 U8459 ( .A1(n9500), .A2(n9139), .B1(n9141), .B2(n9524), .ZN(n6652)
         );
  OAI21_X1 U8460 ( .B1(n6654), .B2(n6653), .A(n6652), .ZN(n6760) );
  AOI211_X1 U8461 ( .C1(n9869), .C2(n6754), .A(n6755), .B(n6760), .ZN(n6659)
         );
  OAI22_X1 U8462 ( .A1(n9676), .A2(n6835), .B1(n9871), .B2(n5102), .ZN(n6655)
         );
  INV_X1 U8463 ( .A(n6655), .ZN(n6656) );
  OAI21_X1 U8464 ( .B1(n6659), .B2(n6369), .A(n6656), .ZN(P1_U3468) );
  OAI22_X1 U8465 ( .A1(n9633), .A2(n6835), .B1(n9876), .B2(n6455), .ZN(n6657)
         );
  INV_X1 U8466 ( .A(n6657), .ZN(n6658) );
  OAI21_X1 U8467 ( .B1(n6659), .B2(n6362), .A(n6658), .ZN(P1_U3527) );
  INV_X1 U8468 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6703) );
  INV_X1 U8469 ( .A(n6671), .ZN(n6660) );
  MUX2_X1 U8470 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8444), .Z(n6796) );
  XNOR2_X1 U8471 ( .A(n6796), .B(n6812), .ZN(n6798) );
  MUX2_X1 U8472 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8444), .Z(n6669) );
  MUX2_X1 U8473 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8626), .Z(n6663) );
  INV_X1 U8474 ( .A(n6732), .ZN(n6661) );
  XNOR2_X1 U8475 ( .A(n6663), .B(n6661), .ZN(n6734) );
  INV_X1 U8476 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6675) );
  MUX2_X1 U8477 ( .A(n6675), .B(n6662), .S(n8626), .Z(n9880) );
  NAND2_X1 U8478 ( .A1(n9880), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9879) );
  AND2_X1 U8479 ( .A1(n6663), .A2(n6732), .ZN(n6664) );
  AOI21_X1 U8480 ( .B1(n6734), .B2(n9879), .A(n6664), .ZN(n6718) );
  MUX2_X1 U8481 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8626), .Z(n6665) );
  XNOR2_X1 U8482 ( .A(n6665), .B(n4354), .ZN(n6716) );
  INV_X1 U8483 ( .A(n4354), .ZN(n6667) );
  INV_X1 U8484 ( .A(n6665), .ZN(n6666) );
  OAI22_X1 U8485 ( .A1(n6718), .A2(n6716), .B1(n6667), .B2(n6666), .ZN(n6782)
         );
  MUX2_X1 U8486 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8444), .Z(n6668) );
  XNOR2_X1 U8487 ( .A(n6668), .B(n6691), .ZN(n6783) );
  NOR2_X1 U8488 ( .A1(n6782), .A2(n6783), .ZN(n6781) );
  NOR2_X1 U8489 ( .A1(n6668), .A2(n6691), .ZN(n6775) );
  XNOR2_X1 U8490 ( .A(n6669), .B(n6695), .ZN(n6774) );
  NOR3_X1 U8491 ( .A1(n6781), .A2(n6775), .A3(n6774), .ZN(n6773) );
  AOI21_X1 U8492 ( .B1(n6669), .B2(n6695), .A(n6773), .ZN(n6799) );
  XOR2_X1 U8493 ( .A(n6798), .B(n6799), .Z(n6670) );
  NOR2_X2 U8494 ( .A1(n8609), .A2(n8445), .ZN(n9883) );
  NAND2_X1 U8495 ( .A1(n6670), .A2(n9883), .ZN(n6702) );
  OR2_X1 U8496 ( .A1(n8444), .A2(P2_U3151), .ZN(n8970) );
  OR3_X1 U8497 ( .A1(n6685), .A2(n8445), .A3(n8970), .ZN(n6673) );
  OR2_X1 U8498 ( .A1(n6131), .A2(P2_U3151), .ZN(n8966) );
  OR2_X1 U8499 ( .A1(n6671), .A2(n8966), .ZN(n6672) );
  NOR2_X1 U8500 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5766), .ZN(n7238) );
  INV_X1 U8501 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6684) );
  INV_X1 U8502 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6674) );
  MUX2_X1 U8503 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6674), .S(n6708), .Z(n6706)
         );
  NOR2_X1 U8504 ( .A1(n6675), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6676) );
  INV_X1 U8505 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6972) );
  NAND2_X1 U8506 ( .A1(n6730), .A2(n6677), .ZN(n6705) );
  NAND2_X1 U8507 ( .A1(n6706), .A2(n6705), .ZN(n6704) );
  NAND2_X1 U8508 ( .A1(n4354), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6678) );
  NAND2_X1 U8509 ( .A1(n6704), .A2(n6678), .ZN(n6679) );
  NAND2_X1 U8510 ( .A1(n6679), .A2(n6691), .ZN(n6766) );
  OAI21_X1 U8511 ( .B1(n6679), .B2(n6691), .A(n6766), .ZN(n6787) );
  INV_X1 U8512 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8513 ( .A1(n6785), .A2(n6766), .ZN(n6681) );
  INV_X1 U8514 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6680) );
  MUX2_X1 U8515 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6680), .S(n6695), .Z(n6765)
         );
  AOI21_X1 U8516 ( .B1(n6684), .B2(n6683), .A(n6808), .ZN(n6699) );
  OR2_X1 U8517 ( .A1(n6685), .A2(n8966), .ZN(n9878) );
  INV_X1 U8518 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6687) );
  MUX2_X1 U8519 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6687), .S(n4354), .Z(n6711)
         );
  AND2_X1 U8520 ( .A1(n4857), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6688) );
  OAI21_X1 U8521 ( .B1(n6732), .B2(n6688), .A(n6689), .ZN(n6726) );
  INV_X1 U8522 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6727) );
  OR2_X1 U8523 ( .A1(n6726), .A2(n6727), .ZN(n6724) );
  NAND2_X1 U8524 ( .A1(n6724), .A2(n6689), .ZN(n6710) );
  NAND2_X1 U8525 ( .A1(n6711), .A2(n6710), .ZN(n6709) );
  NAND2_X1 U8526 ( .A1(n4354), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U8527 ( .A1(n6709), .A2(n6690), .ZN(n6692) );
  XNOR2_X1 U8528 ( .A(n6692), .B(n6691), .ZN(n6784) );
  INV_X1 U8529 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6694) );
  INV_X1 U8530 ( .A(n6691), .ZN(n6792) );
  INV_X1 U8531 ( .A(n6692), .ZN(n6693) );
  INV_X1 U8532 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9942) );
  MUX2_X1 U8533 ( .A(n9942), .B(P2_REG1_REG_4__SCAN_IN), .S(n6695), .Z(n6763)
         );
  NAND2_X1 U8534 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n6696), .ZN(n6813) );
  OAI21_X1 U8535 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n6696), .A(n6813), .ZN(
        n6697) );
  INV_X1 U8536 ( .A(n6697), .ZN(n6698) );
  OAI22_X1 U8537 ( .A1(n6699), .A2(n8642), .B1(n8635), .B2(n6698), .ZN(n6700)
         );
  AOI211_X1 U8538 ( .C1(n6807), .C2(n8559), .A(n7238), .B(n6700), .ZN(n6701)
         );
  OAI211_X1 U8539 ( .C1(n6703), .C2(n8618), .A(n6702), .B(n6701), .ZN(P2_U3187) );
  INV_X1 U8540 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6722) );
  INV_X1 U8541 ( .A(n8642), .ZN(n6820) );
  OAI21_X1 U8542 ( .B1(n6706), .B2(n6705), .A(n6704), .ZN(n6715) );
  INV_X1 U8543 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6707) );
  OAI22_X1 U8544 ( .A1(n9886), .A2(n4354), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6707), .ZN(n6714) );
  OAI21_X1 U8545 ( .B1(n6711), .B2(n6710), .A(n6709), .ZN(n6712) );
  AND2_X1 U8546 ( .A1(n8595), .A2(n6712), .ZN(n6713) );
  AOI211_X1 U8547 ( .C1(n6820), .C2(n6715), .A(n6714), .B(n6713), .ZN(n6721)
         );
  INV_X1 U8548 ( .A(n6716), .ZN(n6717) );
  XNOR2_X1 U8549 ( .A(n6718), .B(n6717), .ZN(n6719) );
  NAND2_X1 U8550 ( .A1(n9883), .A2(n6719), .ZN(n6720) );
  OAI211_X1 U8551 ( .C1(n6722), .C2(n8618), .A(n6721), .B(n6720), .ZN(P2_U3184) );
  INV_X2 U8552 ( .A(P1_U3973), .ZN(n9144) );
  NAND2_X1 U8553 ( .A1(n9144), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6723) );
  OAI21_X1 U8554 ( .B1(n9303), .B2(n9144), .A(n6723), .ZN(P1_U3583) );
  INV_X1 U8555 ( .A(n6724), .ZN(n6725) );
  AOI21_X1 U8556 ( .B1(n6727), .B2(n6726), .A(n6725), .ZN(n6738) );
  INV_X1 U8557 ( .A(n8618), .ZN(n9877) );
  NAND2_X1 U8558 ( .A1(n6728), .A2(n6972), .ZN(n6729) );
  AND2_X1 U8559 ( .A1(n6730), .A2(n6729), .ZN(n6731) );
  OAI22_X1 U8560 ( .A1(n9886), .A2(n6732), .B1(n8642), .B2(n6731), .ZN(n6733)
         );
  AOI21_X1 U8561 ( .B1(n9877), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n6733), .ZN(
        n6737) );
  XOR2_X1 U8562 ( .A(n9879), .B(n6734), .Z(n6735) );
  AOI22_X1 U8563 ( .A1(n9883), .A2(n6735), .B1(P2_U3151), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6736) );
  OAI211_X1 U8564 ( .C1(n6738), .C2(n8635), .A(n6737), .B(n6736), .ZN(P2_U3183) );
  XOR2_X1 U8565 ( .A(n6744), .B(n6864), .Z(n6742) );
  OAI22_X1 U8566 ( .A1(n6740), .A2(n9516), .B1(n6739), .B2(n9380), .ZN(n6910)
         );
  INV_X1 U8567 ( .A(n6910), .ZN(n6741) );
  OAI21_X1 U8568 ( .B1(n6742), .B2(n9518), .A(n6741), .ZN(n6851) );
  INV_X1 U8569 ( .A(n6851), .ZN(n6753) );
  OAI21_X1 U8570 ( .B1(n6745), .B2(n6744), .A(n6743), .ZN(n6853) );
  OAI21_X1 U8571 ( .B1(n6746), .B2(n6914), .A(n9531), .ZN(n6747) );
  NOR2_X1 U8572 ( .A1(n6747), .A2(n6959), .ZN(n6852) );
  NAND2_X1 U8573 ( .A1(n6852), .A2(n9527), .ZN(n6750) );
  INV_X1 U8574 ( .A(n6748), .ZN(n6911) );
  INV_X1 U8575 ( .A(n9390), .ZN(n9834) );
  AOI22_X1 U8576 ( .A1(n9826), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n6911), .B2(
        n9834), .ZN(n6749) );
  OAI211_X1 U8577 ( .C1(n6914), .C2(n9514), .A(n6750), .B(n6749), .ZN(n6751)
         );
  AOI21_X1 U8578 ( .B1(n6853), .B2(n9836), .A(n6751), .ZN(n6752) );
  OAI21_X1 U8579 ( .B1(n6753), .B2(n9826), .A(n6752), .ZN(P1_U3287) );
  INV_X1 U8580 ( .A(n6754), .ZN(n6762) );
  NAND2_X1 U8581 ( .A1(n6755), .A2(n9527), .ZN(n6758) );
  INV_X1 U8582 ( .A(n6756), .ZN(n6838) );
  AOI22_X1 U8583 ( .A1(n9826), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6838), .B2(
        n9834), .ZN(n6757) );
  OAI211_X1 U8584 ( .C1(n6835), .C2(n9514), .A(n6758), .B(n6757), .ZN(n6759)
         );
  AOI21_X1 U8585 ( .B1(n9468), .B2(n6760), .A(n6759), .ZN(n6761) );
  OAI21_X1 U8586 ( .B1(n6762), .B2(n9529), .A(n6761), .ZN(P1_U3288) );
  INV_X1 U8587 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6780) );
  NOR2_X1 U8588 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10141), .ZN(n7213) );
  XNOR2_X1 U8589 ( .A(n6764), .B(n6763), .ZN(n6771) );
  INV_X1 U8590 ( .A(n6765), .ZN(n6767) );
  NAND3_X1 U8591 ( .A1(n6785), .A2(n6767), .A3(n6766), .ZN(n6768) );
  AND2_X1 U8592 ( .A1(n6769), .A2(n6768), .ZN(n6770) );
  OAI22_X1 U8593 ( .A1(n6771), .A2(n8635), .B1(n8642), .B2(n6770), .ZN(n6772)
         );
  AOI211_X1 U8594 ( .C1(n6682), .C2(n8559), .A(n7213), .B(n6772), .ZN(n6779)
         );
  INV_X1 U8595 ( .A(n6773), .ZN(n6777) );
  OAI21_X1 U8596 ( .B1(n6781), .B2(n6775), .A(n6774), .ZN(n6776) );
  NAND3_X1 U8597 ( .A1(n6777), .A2(n9883), .A3(n6776), .ZN(n6778) );
  OAI211_X1 U8598 ( .C1(n6780), .C2(n8618), .A(n6779), .B(n6778), .ZN(P2_U3186) );
  AOI21_X1 U8599 ( .B1(n6783), .B2(n6782), .A(n6781), .ZN(n6795) );
  INV_X1 U8600 ( .A(n9883), .ZN(n8591) );
  NOR2_X1 U8601 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10165), .ZN(n7067) );
  XNOR2_X1 U8602 ( .A(n6784), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6790) );
  INV_X1 U8603 ( .A(n6785), .ZN(n6786) );
  AOI21_X1 U8604 ( .B1(n6788), .B2(n6787), .A(n6786), .ZN(n6789) );
  OAI22_X1 U8605 ( .A1(n6790), .A2(n8635), .B1(n8642), .B2(n6789), .ZN(n6791)
         );
  AOI211_X1 U8606 ( .C1(n6792), .C2(n8559), .A(n7067), .B(n6791), .ZN(n6794)
         );
  NAND2_X1 U8607 ( .A1(n9877), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n6793) );
  OAI211_X1 U8608 ( .C1(n6795), .C2(n8591), .A(n6794), .B(n6793), .ZN(P2_U3185) );
  INV_X1 U8609 ( .A(n6796), .ZN(n6797) );
  OAI22_X1 U8610 ( .A1(n6799), .A2(n6798), .B1(n6807), .B2(n6797), .ZN(n6804)
         );
  INV_X1 U8611 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6800) );
  INV_X1 U8612 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6815) );
  MUX2_X1 U8613 ( .A(n6800), .B(n6815), .S(n8444), .Z(n6802) );
  INV_X1 U8614 ( .A(n6894), .ZN(n6801) );
  NAND2_X1 U8615 ( .A1(n6802), .A2(n6801), .ZN(n6884) );
  OAI21_X1 U8616 ( .B1(n6802), .B2(n6801), .A(n6884), .ZN(n6803) );
  NOR2_X1 U8617 ( .A1(n6804), .A2(n6803), .ZN(n6891) );
  AOI21_X1 U8618 ( .B1(n6804), .B2(n6803), .A(n6891), .ZN(n6826) );
  NOR2_X1 U8619 ( .A1(n6807), .A2(n6806), .ZN(n6809) );
  NAND2_X1 U8620 ( .A1(n6894), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6880) );
  OR2_X1 U8621 ( .A1(n6894), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6810) );
  OAI21_X1 U8622 ( .B1(n4746), .B2(n4430), .A(n6881), .ZN(n6819) );
  NAND2_X1 U8623 ( .A1(n6812), .A2(n6811), .ZN(n6814) );
  NAND2_X1 U8624 ( .A1(n6814), .A2(n6813), .ZN(n6817) );
  MUX2_X1 U8625 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6815), .S(n6894), .Z(n6816)
         );
  NAND2_X1 U8626 ( .A1(n6816), .A2(n6817), .ZN(n6895) );
  OAI21_X1 U8627 ( .B1(n6817), .B2(n6816), .A(n6895), .ZN(n6818) );
  AOI22_X1 U8628 ( .A1(n6820), .A2(n6819), .B1(n8595), .B2(n6818), .ZN(n6823)
         );
  INV_X1 U8629 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6821) );
  NOR2_X1 U8630 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6821), .ZN(n7296) );
  INV_X1 U8631 ( .A(n7296), .ZN(n6822) );
  OAI211_X1 U8632 ( .C1(n9886), .C2(n6894), .A(n6823), .B(n6822), .ZN(n6824)
         );
  AOI21_X1 U8633 ( .B1(n9877), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6824), .ZN(
        n6825) );
  OAI21_X1 U8634 ( .B1(n6826), .B2(n8591), .A(n6825), .ZN(P2_U3188) );
  INV_X1 U8635 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6828) );
  INV_X1 U8636 ( .A(n6827), .ZN(n6829) );
  OAI222_X1 U8637 ( .A1(n7957), .A2(n6828), .B1(n8960), .B2(n6829), .C1(
        P2_U3151), .C2(n8526), .ZN(P2_U3280) );
  INV_X1 U8638 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6830) );
  INV_X1 U8639 ( .A(n9804), .ZN(n7164) );
  OAI222_X1 U8640 ( .A1(n9694), .A2(n6830), .B1(n9688), .B2(n6829), .C1(
        P1_U3086), .C2(n7164), .ZN(P1_U3340) );
  NAND2_X1 U8641 ( .A1(n4429), .A2(n6831), .ZN(n6833) );
  XNOR2_X1 U8642 ( .A(n6833), .B(n6832), .ZN(n6840) );
  OAI22_X1 U8643 ( .A1(n9124), .A2(n6835), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6834), .ZN(n6837) );
  OAI22_X1 U8644 ( .A1(n6953), .A2(n9119), .B1(n9083), .B2(n6290), .ZN(n6836)
         );
  AOI211_X1 U8645 ( .C1(n6838), .C2(n9121), .A(n6837), .B(n6836), .ZN(n6839)
         );
  OAI21_X1 U8646 ( .B1(n6840), .B2(n9098), .A(n6839), .ZN(P1_U3227) );
  OAI21_X1 U8647 ( .B1(n6842), .B2(n6846), .A(n6841), .ZN(n7087) );
  AND2_X1 U8648 ( .A1(n6845), .A2(n6844), .ZN(n6847) );
  XNOR2_X1 U8649 ( .A(n6847), .B(n6846), .ZN(n6848) );
  OAI222_X1 U8650 ( .A1(n9712), .A2(n7236), .B1(n9710), .B2(n4562), .C1(n9708), 
        .C2(n6848), .ZN(n7084) );
  AOI21_X1 U8651 ( .B1(n9933), .B2(n7087), .A(n7084), .ZN(n7153) );
  OAI22_X1 U8652 ( .A1(n8855), .A2(n7150), .B1(n9950), .B2(n6694), .ZN(n6849)
         );
  INV_X1 U8653 ( .A(n6849), .ZN(n6850) );
  OAI21_X1 U8654 ( .B1(n7153), .B2(n6277), .A(n6850), .ZN(P2_U3462) );
  AOI211_X1 U8655 ( .C1(n9869), .C2(n6853), .A(n6852), .B(n6851), .ZN(n6858)
         );
  OAI22_X1 U8656 ( .A1(n9676), .A2(n6914), .B1(n9871), .B2(n5119), .ZN(n6854)
         );
  INV_X1 U8657 ( .A(n6854), .ZN(n6855) );
  OAI21_X1 U8658 ( .B1(n6858), .B2(n6369), .A(n6855), .ZN(P1_U3471) );
  OAI22_X1 U8659 ( .A1(n9633), .A2(n6914), .B1(n9876), .B2(n6457), .ZN(n6856)
         );
  INV_X1 U8660 ( .A(n6856), .ZN(n6857) );
  OAI21_X1 U8661 ( .B1(n6858), .B2(n6362), .A(n6857), .ZN(P1_U3528) );
  INV_X1 U8662 ( .A(n6859), .ZN(n6918) );
  INV_X1 U8663 ( .A(n8582), .ZN(n8578) );
  INV_X1 U8664 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6860) );
  OAI222_X1 U8665 ( .A1(n8960), .A2(n6918), .B1(n8578), .B2(P2_U3151), .C1(
        n6860), .C2(n7957), .ZN(P2_U3279) );
  OAI21_X1 U8666 ( .B1(n6862), .B2(n6866), .A(n6861), .ZN(n9859) );
  INV_X1 U8667 ( .A(n9859), .ZN(n6879) );
  INV_X1 U8668 ( .A(n7694), .ZN(n6863) );
  OR2_X1 U8669 ( .A1(n6864), .A2(n6863), .ZN(n6865) );
  NAND2_X1 U8670 ( .A1(n6865), .A2(n7675), .ZN(n6951) );
  INV_X1 U8671 ( .A(n7696), .ZN(n6950) );
  NAND2_X1 U8672 ( .A1(n6951), .A2(n6950), .ZN(n6949) );
  INV_X1 U8673 ( .A(n6866), .ZN(n6867) );
  NAND3_X1 U8674 ( .A1(n6949), .A2(n6867), .A3(n6868), .ZN(n7037) );
  NAND2_X1 U8675 ( .A1(n7037), .A2(n9503), .ZN(n6871) );
  AOI21_X1 U8676 ( .B1(n6949), .B2(n6868), .A(n6867), .ZN(n6870) );
  AOI22_X1 U8677 ( .A1(n9500), .A2(n4726), .B1(n9138), .B2(n9524), .ZN(n6869)
         );
  OAI21_X1 U8678 ( .B1(n6871), .B2(n6870), .A(n6869), .ZN(n9857) );
  INV_X1 U8679 ( .A(n6958), .ZN(n6872) );
  INV_X1 U8680 ( .A(n6875), .ZN(n9856) );
  OAI211_X1 U8681 ( .C1(n6872), .C2(n9856), .A(n9531), .B(n7044), .ZN(n9855)
         );
  OAI22_X1 U8682 ( .A1(n9468), .A2(n6873), .B1(n7307), .B2(n9390), .ZN(n6874)
         );
  AOI21_X1 U8683 ( .B1(n9838), .B2(n6875), .A(n6874), .ZN(n6876) );
  OAI21_X1 U8684 ( .B1(n9855), .B2(n9841), .A(n6876), .ZN(n6877) );
  AOI21_X1 U8685 ( .B1(n9857), .B2(n9468), .A(n6877), .ZN(n6878) );
  OAI21_X1 U8686 ( .B1(n6879), .B2(n9529), .A(n6878), .ZN(P1_U3285) );
  INV_X1 U8687 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6883) );
  AOI21_X1 U8688 ( .B1(n6883), .B2(n6882), .A(n6986), .ZN(n6905) );
  INV_X1 U8689 ( .A(n6884), .ZN(n6890) );
  MUX2_X1 U8690 ( .A(n6883), .B(n6885), .S(n8444), .Z(n6886) );
  NAND2_X1 U8691 ( .A1(n6886), .A2(n6985), .ZN(n6996) );
  INV_X1 U8692 ( .A(n6886), .ZN(n6887) );
  NAND2_X1 U8693 ( .A1(n6887), .A2(n7000), .ZN(n6888) );
  AND2_X1 U8694 ( .A1(n6996), .A2(n6888), .ZN(n6889) );
  OAI21_X1 U8695 ( .B1(n6891), .B2(n6890), .A(n6889), .ZN(n6997) );
  INV_X1 U8696 ( .A(n6997), .ZN(n6893) );
  NOR3_X1 U8697 ( .A1(n6891), .A2(n6890), .A3(n6889), .ZN(n6892) );
  OAI21_X1 U8698 ( .B1(n6893), .B2(n6892), .A(n9883), .ZN(n6904) );
  NAND2_X1 U8699 ( .A1(n6894), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8700 ( .A1(n6896), .A2(n6895), .ZN(n6999) );
  XNOR2_X1 U8701 ( .A(n6999), .B(n6985), .ZN(n6897) );
  NAND2_X1 U8702 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(n6897), .ZN(n7001) );
  OAI21_X1 U8703 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n6897), .A(n7001), .ZN(
        n6902) );
  INV_X1 U8704 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10130) );
  NOR2_X1 U8705 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10130), .ZN(n7463) );
  INV_X1 U8706 ( .A(n7463), .ZN(n6898) );
  OAI21_X1 U8707 ( .B1(n9886), .B2(n7000), .A(n6898), .ZN(n6901) );
  INV_X1 U8708 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6899) );
  NOR2_X1 U8709 ( .A1(n8618), .A2(n6899), .ZN(n6900) );
  AOI211_X1 U8710 ( .C1(n8595), .C2(n6902), .A(n6901), .B(n6900), .ZN(n6903)
         );
  OAI211_X1 U8711 ( .C1(n6905), .C2(n8642), .A(n6904), .B(n6903), .ZN(P2_U3189) );
  XNOR2_X1 U8712 ( .A(n6907), .B(n6906), .ZN(n6908) );
  XNOR2_X1 U8713 ( .A(n6909), .B(n6908), .ZN(n6916) );
  AOI22_X1 U8714 ( .A1(n9060), .A2(n6910), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n6913) );
  NAND2_X1 U8715 ( .A1(n9121), .A2(n6911), .ZN(n6912) );
  OAI211_X1 U8716 ( .C1(n6914), .C2(n9124), .A(n6913), .B(n6912), .ZN(n6915)
         );
  AOI21_X1 U8717 ( .B1(n6916), .B2(n9115), .A(n6915), .ZN(n6917) );
  INV_X1 U8718 ( .A(n6917), .ZN(P1_U3239) );
  INV_X1 U8719 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6919) );
  INV_X1 U8720 ( .A(n7346), .ZN(n7341) );
  OAI222_X1 U8721 ( .A1(n9694), .A2(n6919), .B1(n9688), .B2(n6918), .C1(n7341), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  OR2_X1 U8722 ( .A1(n6922), .A2(n9925), .ZN(n6920) );
  INV_X1 U8723 ( .A(n8196), .ZN(n8213) );
  OR2_X1 U8724 ( .A1(n6922), .A2(n6921), .ZN(n6926) );
  INV_X1 U8725 ( .A(n6923), .ZN(n6935) );
  NAND2_X1 U8726 ( .A1(n6924), .A2(n6935), .ZN(n6925) );
  NOR2_X1 U8727 ( .A1(n6927), .A2(n6978), .ZN(n7024) );
  INV_X1 U8728 ( .A(n7023), .ZN(n6928) );
  NAND2_X2 U8729 ( .A1(n7024), .A2(n6928), .ZN(n8207) );
  INV_X1 U8730 ( .A(n8207), .ZN(n8117) );
  AOI22_X1 U8731 ( .A1(n8179), .A2(n8246), .B1(n8117), .B2(n5819), .ZN(n6944)
         );
  NAND2_X1 U8732 ( .A1(n6930), .A2(n6929), .ZN(n6937) );
  NAND3_X1 U8733 ( .A1(n6933), .A2(n6932), .A3(n6931), .ZN(n6934) );
  AOI21_X1 U8734 ( .B1(n6940), .B2(n6935), .A(n6934), .ZN(n6936) );
  NAND2_X1 U8735 ( .A1(n6937), .A2(n6936), .ZN(n6938) );
  NAND2_X1 U8736 ( .A1(n6938), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6942) );
  NOR2_X1 U8737 ( .A1(n6939), .A2(n6978), .ZN(n8446) );
  NAND2_X1 U8738 ( .A1(n6940), .A2(n8446), .ZN(n6941) );
  NAND2_X1 U8739 ( .A1(n8183), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8740 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n7033), .ZN(n6943) );
  OAI211_X1 U8741 ( .C1(n8213), .C2(n6945), .A(n6944), .B(n6943), .ZN(P2_U3172) );
  INV_X1 U8742 ( .A(n6946), .ZN(n7334) );
  XNOR2_X1 U8743 ( .A(n6947), .B(n7696), .ZN(n9849) );
  INV_X1 U8744 ( .A(n7332), .ZN(n6948) );
  NAND2_X1 U8745 ( .A1(n9849), .A2(n6948), .ZN(n6956) );
  OAI21_X1 U8746 ( .B1(n6951), .B2(n6950), .A(n6949), .ZN(n6954) );
  OAI22_X1 U8747 ( .A1(n6953), .A2(n9380), .B1(n6952), .B2(n9516), .ZN(n7076)
         );
  AOI21_X1 U8748 ( .B1(n6954), .B2(n9503), .A(n7076), .ZN(n6955) );
  NAND2_X1 U8749 ( .A1(n6956), .A2(n6955), .ZN(n9854) );
  AOI21_X1 U8750 ( .B1(n7334), .B2(n9849), .A(n9854), .ZN(n6964) );
  OAI22_X1 U8751 ( .A1(n9468), .A2(n6957), .B1(n7077), .B2(n9390), .ZN(n6961)
         );
  OAI211_X1 U8752 ( .C1(n6959), .C2(n9851), .A(n9531), .B(n6958), .ZN(n9850)
         );
  NOR2_X1 U8753 ( .A1(n9850), .A2(n9841), .ZN(n6960) );
  AOI211_X1 U8754 ( .C1(n9838), .C2(n6962), .A(n6961), .B(n6960), .ZN(n6963)
         );
  OAI21_X1 U8755 ( .B1(n6964), .B2(n9826), .A(n6963), .ZN(P1_U3286) );
  INV_X1 U8756 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U8757 ( .A1(n9937), .A2(n6965), .ZN(n6966) );
  OAI21_X1 U8758 ( .B1(n9937), .B2(n6967), .A(n6966), .ZN(P2_U3390) );
  INV_X1 U8759 ( .A(n8270), .ZN(n6968) );
  XNOR2_X1 U8760 ( .A(n6968), .B(n8244), .ZN(n9887) );
  XOR2_X1 U8761 ( .A(n8244), .B(n6970), .Z(n6971) );
  OAI222_X1 U8762 ( .A1(n9710), .A2(n6969), .B1(n9712), .B2(n4562), .C1(n9708), 
        .C2(n6971), .ZN(n9889) );
  NOR2_X1 U8763 ( .A1(n9716), .A2(n6972), .ZN(n6976) );
  INV_X1 U8764 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6974) );
  OAI22_X1 U8765 ( .A1(n8807), .A2(n6973), .B1(n6974), .B2(n9697), .ZN(n6975)
         );
  AOI211_X1 U8766 ( .C1(n9716), .C2(n9889), .A(n6976), .B(n6975), .ZN(n6977)
         );
  OAI21_X1 U8767 ( .B1(n9887), .B2(n8795), .A(n6977), .ZN(P2_U3232) );
  NAND3_X1 U8768 ( .A1(n8246), .A2(n9925), .A3(n6978), .ZN(n6980) );
  OAI211_X1 U8769 ( .C1(n9697), .C2(n10044), .A(n6980), .B(n6979), .ZN(n6981)
         );
  MUX2_X1 U8770 ( .A(P2_REG2_REG_0__SCAN_IN), .B(n6981), .S(n9716), .Z(n6982)
         );
  AOI21_X1 U8771 ( .B1(n8792), .B2(n7021), .A(n6982), .ZN(n6983) );
  INV_X1 U8772 ( .A(n6983), .ZN(P2_U3233) );
  NAND2_X1 U8773 ( .A1(n7102), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7089) );
  INV_X1 U8774 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U8775 ( .A1(n7003), .A2(n6991), .ZN(n6987) );
  NAND2_X1 U8776 ( .A1(n7089), .A2(n6987), .ZN(n6989) );
  INV_X1 U8777 ( .A(n7090), .ZN(n6988) );
  AOI21_X1 U8778 ( .B1(n6990), .B2(n6989), .A(n6988), .ZN(n7014) );
  INV_X1 U8779 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7004) );
  MUX2_X1 U8780 ( .A(n6991), .B(n7004), .S(n8444), .Z(n6992) );
  NAND2_X1 U8781 ( .A1(n6992), .A2(n7003), .ZN(n7092) );
  INV_X1 U8782 ( .A(n6992), .ZN(n6993) );
  NAND2_X1 U8783 ( .A1(n6993), .A2(n7102), .ZN(n6994) );
  NAND2_X1 U8784 ( .A1(n7092), .A2(n6994), .ZN(n6995) );
  AOI21_X1 U8785 ( .B1(n6997), .B2(n6996), .A(n6995), .ZN(n7099) );
  AND3_X1 U8786 ( .A1(n6997), .A2(n6996), .A3(n6995), .ZN(n6998) );
  OAI21_X1 U8787 ( .B1(n7099), .B2(n6998), .A(n9883), .ZN(n7013) );
  NAND2_X1 U8788 ( .A1(n7000), .A2(n6999), .ZN(n7002) );
  NAND2_X1 U8789 ( .A1(n7002), .A2(n7001), .ZN(n7006) );
  MUX2_X1 U8790 ( .A(n7004), .B(P2_REG1_REG_8__SCAN_IN), .S(n7003), .Z(n7005)
         );
  NAND2_X1 U8791 ( .A1(n7005), .A2(n7006), .ZN(n7103) );
  OAI21_X1 U8792 ( .B1(n7006), .B2(n7005), .A(n7103), .ZN(n7011) );
  INV_X1 U8793 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10157) );
  NOR2_X1 U8794 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10157), .ZN(n7524) );
  INV_X1 U8795 ( .A(n7524), .ZN(n7007) );
  OAI21_X1 U8796 ( .B1(n9886), .B2(n7102), .A(n7007), .ZN(n7010) );
  INV_X1 U8797 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7008) );
  NOR2_X1 U8798 ( .A1(n8618), .A2(n7008), .ZN(n7009) );
  AOI211_X1 U8799 ( .C1(n8595), .C2(n7011), .A(n7010), .B(n7009), .ZN(n7012)
         );
  OAI211_X1 U8800 ( .C1(n7014), .C2(n8642), .A(n7013), .B(n7012), .ZN(P2_U3190) );
  NAND2_X1 U8801 ( .A1(n7015), .A2(n8423), .ZN(n7016) );
  AND2_X1 U8802 ( .A1(n7017), .A2(n7016), .ZN(n7018) );
  XOR2_X1 U8803 ( .A(n6843), .B(n7059), .Z(n7061) );
  OAI21_X1 U8804 ( .B1(n7020), .B2(n7021), .A(n8270), .ZN(n7030) );
  AOI22_X1 U8805 ( .A1(n7029), .A2(n7030), .B1(n5811), .B2(n7022), .ZN(n7062)
         );
  XOR2_X1 U8806 ( .A(n7061), .B(n7062), .Z(n7028) );
  OAI21_X1 U8807 ( .B1(n7211), .B2(n8207), .A(n7025), .ZN(n7026) );
  AOI21_X1 U8808 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7033), .A(n7026), .ZN(
        n7027) );
  OAI21_X1 U8809 ( .B1(n7028), .B2(n8199), .A(n7027), .ZN(P2_U3177) );
  XOR2_X1 U8810 ( .A(n7029), .B(n7030), .Z(n7035) );
  AOI22_X1 U8811 ( .A1(n8205), .A2(n8466), .B1(n8196), .B2(n5820), .ZN(n7031)
         );
  OAI21_X1 U8812 ( .B1(n4562), .B2(n8207), .A(n7031), .ZN(n7032) );
  AOI21_X1 U8813 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7033), .A(n7032), .ZN(
        n7034) );
  OAI21_X1 U8814 ( .B1(n8199), .B2(n7035), .A(n7034), .ZN(P2_U3162) );
  NAND2_X1 U8815 ( .A1(n8609), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7036) );
  OAI21_X1 U8816 ( .B1(n8034), .B2(n8609), .A(n7036), .ZN(P2_U3520) );
  NAND2_X1 U8817 ( .A1(n7037), .A2(n7678), .ZN(n7038) );
  XNOR2_X1 U8818 ( .A(n7038), .B(n7041), .ZN(n7039) );
  AOI22_X1 U8819 ( .A1(n7039), .A2(n9503), .B1(n9524), .B2(n9137), .ZN(n9861)
         );
  OAI21_X1 U8820 ( .B1(n7042), .B2(n7041), .A(n7040), .ZN(n9863) );
  NAND2_X1 U8821 ( .A1(n9863), .A2(n9836), .ZN(n7050) );
  OAI22_X1 U8822 ( .A1(n9468), .A2(n7043), .B1(n7381), .B2(n9390), .ZN(n7048)
         );
  XNOR2_X1 U8823 ( .A(n7044), .B(n4691), .ZN(n7046) );
  NOR2_X1 U8824 ( .A1(n7380), .A2(n9516), .ZN(n7045) );
  AOI21_X1 U8825 ( .B1(n7046), .B2(n9531), .A(n7045), .ZN(n9860) );
  NOR2_X1 U8826 ( .A1(n9860), .A2(n9841), .ZN(n7047) );
  AOI211_X1 U8827 ( .C1(n9838), .C2(n7384), .A(n7048), .B(n7047), .ZN(n7049)
         );
  OAI211_X1 U8828 ( .C1(n9861), .C2(n9826), .A(n7050), .B(n7049), .ZN(P1_U3284) );
  INV_X1 U8829 ( .A(n8280), .ZN(n8309) );
  NOR2_X1 U8830 ( .A1(n8309), .A2(n8287), .ZN(n7053) );
  INV_X1 U8831 ( .A(n7051), .ZN(n7052) );
  AOI21_X1 U8832 ( .B1(n7053), .B2(n6841), .A(n7052), .ZN(n9899) );
  XOR2_X1 U8833 ( .A(n8287), .B(n7054), .Z(n7055) );
  AOI222_X1 U8834 ( .A1(n8817), .A2(n7055), .B1(n8465), .B2(n8822), .C1(n8463), 
        .C2(n8819), .ZN(n9897) );
  MUX2_X1 U8835 ( .A(n6680), .B(n9897), .S(n9716), .Z(n7058) );
  INV_X1 U8836 ( .A(n7216), .ZN(n7056) );
  AOI22_X1 U8837 ( .A1(n8792), .A2(n8306), .B1(n8805), .B2(n7056), .ZN(n7057)
         );
  OAI211_X1 U8838 ( .C1(n9899), .C2(n8795), .A(n7058), .B(n7057), .ZN(P2_U3229) );
  XNOR2_X1 U8839 ( .A(n7020), .B(n7068), .ZN(n7204) );
  XOR2_X1 U8840 ( .A(n8465), .B(n7204), .Z(n7064) );
  INV_X1 U8841 ( .A(n7059), .ZN(n7060) );
  OAI22_X1 U8842 ( .A1(n7062), .A2(n7061), .B1(n7060), .B2(n6843), .ZN(n7063)
         );
  AOI211_X1 U8843 ( .C1(n7064), .C2(n7063), .A(n8199), .B(n7205), .ZN(n7065)
         );
  INV_X1 U8844 ( .A(n7065), .ZN(n7070) );
  OAI22_X1 U8845 ( .A1(n8120), .A2(n4562), .B1(n7236), .B2(n8207), .ZN(n7066)
         );
  AOI211_X1 U8846 ( .C1(n7068), .C2(n8196), .A(n7067), .B(n7066), .ZN(n7069)
         );
  OAI211_X1 U8847 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8183), .A(n7070), .B(
        n7069), .ZN(P2_U3158) );
  INV_X1 U8848 ( .A(n7071), .ZN(n7072) );
  NOR2_X1 U8849 ( .A1(n7073), .A2(n7072), .ZN(n7074) );
  XNOR2_X1 U8850 ( .A(n7075), .B(n7074), .ZN(n7082) );
  AOI22_X1 U8851 ( .A1(n9060), .A2(n7076), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7080) );
  INV_X1 U8852 ( .A(n7077), .ZN(n7078) );
  NAND2_X1 U8853 ( .A1(n9121), .A2(n7078), .ZN(n7079) );
  OAI211_X1 U8854 ( .C1(n9851), .C2(n9124), .A(n7080), .B(n7079), .ZN(n7081)
         );
  AOI21_X1 U8855 ( .B1(n7082), .B2(n9115), .A(n7081), .ZN(n7083) );
  INV_X1 U8856 ( .A(n7083), .ZN(P1_U3213) );
  OAI22_X1 U8857 ( .A1(n8807), .A2(n7150), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9697), .ZN(n7086) );
  MUX2_X1 U8858 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7084), .S(n9716), .Z(n7085)
         );
  AOI211_X1 U8859 ( .C1(n8830), .C2(n7087), .A(n7086), .B(n7085), .ZN(n7088)
         );
  INV_X1 U8860 ( .A(n7088), .ZN(P2_U3230) );
  INV_X1 U8861 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7496) );
  AOI21_X1 U8862 ( .B1(n7496), .B2(n7091), .A(n7176), .ZN(n7113) );
  INV_X1 U8863 ( .A(n7092), .ZN(n7098) );
  MUX2_X1 U8864 ( .A(n7496), .B(n7093), .S(n8444), .Z(n7094) );
  NAND2_X1 U8865 ( .A1(n7094), .A2(n7175), .ZN(n7186) );
  INV_X1 U8866 ( .A(n7094), .ZN(n7095) );
  NAND2_X1 U8867 ( .A1(n7095), .A2(n7190), .ZN(n7096) );
  AND2_X1 U8868 ( .A1(n7186), .A2(n7096), .ZN(n7097) );
  OAI21_X1 U8869 ( .B1(n7099), .B2(n7098), .A(n7097), .ZN(n7187) );
  INV_X1 U8870 ( .A(n7187), .ZN(n7101) );
  NOR3_X1 U8871 ( .A1(n7099), .A2(n7098), .A3(n7097), .ZN(n7100) );
  OAI21_X1 U8872 ( .B1(n7101), .B2(n7100), .A(n9883), .ZN(n7112) );
  INV_X1 U8873 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U8874 ( .A1(n7102), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7104) );
  NAND2_X1 U8875 ( .A1(n7104), .A2(n7103), .ZN(n7189) );
  XNOR2_X1 U8876 ( .A(n7189), .B(n7175), .ZN(n7105) );
  NAND2_X1 U8877 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n7105), .ZN(n7191) );
  OAI21_X1 U8878 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n7105), .A(n7191), .ZN(
        n7106) );
  NAND2_X1 U8879 ( .A1(n7106), .A2(n8595), .ZN(n7108) );
  NOR2_X1 U8880 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5769), .ZN(n7547) );
  AOI21_X1 U8881 ( .B1(n8559), .B2(n7175), .A(n7547), .ZN(n7107) );
  OAI211_X1 U8882 ( .C1(n7109), .C2(n8618), .A(n7108), .B(n7107), .ZN(n7110)
         );
  INV_X1 U8883 ( .A(n7110), .ZN(n7111) );
  OAI211_X1 U8884 ( .C1(n7113), .C2(n8642), .A(n7112), .B(n7111), .ZN(P2_U3191) );
  NAND2_X1 U8885 ( .A1(n7888), .A2(n7886), .ZN(n7114) );
  NAND2_X1 U8886 ( .A1(n7114), .A2(n7120), .ZN(n7116) );
  NAND2_X1 U8887 ( .A1(n7116), .A2(n7115), .ZN(n7118) );
  OAI22_X1 U8888 ( .A1(n7306), .A2(n9380), .B1(n7411), .B2(n9516), .ZN(n7117)
         );
  AOI21_X1 U8889 ( .B1(n7118), .B2(n9503), .A(n7117), .ZN(n9865) );
  OAI21_X1 U8890 ( .B1(n7121), .B2(n7120), .A(n7119), .ZN(n9870) );
  NAND2_X1 U8891 ( .A1(n9870), .A2(n9836), .ZN(n7129) );
  OAI22_X1 U8892 ( .A1(n9468), .A2(n7123), .B1(n7122), .B2(n9390), .ZN(n7126)
         );
  OAI211_X1 U8893 ( .C1(n9867), .C2(n7124), .A(n4366), .B(n9531), .ZN(n9864)
         );
  NOR2_X1 U8894 ( .A1(n9864), .A2(n9841), .ZN(n7125) );
  AOI211_X1 U8895 ( .C1(n9838), .C2(n7127), .A(n7126), .B(n7125), .ZN(n7128)
         );
  OAI211_X1 U8896 ( .C1(n9826), .C2(n9865), .A(n7129), .B(n7128), .ZN(P1_U3283) );
  INV_X1 U8897 ( .A(n8609), .ZN(P2_U3893) );
  INV_X1 U8898 ( .A(n7130), .ZN(n7132) );
  INV_X1 U8899 ( .A(n8605), .ZN(n8611) );
  OAI222_X1 U8900 ( .A1(n7957), .A2(n7131), .B1(n8960), .B2(n7132), .C1(
        P2_U3151), .C2(n8611), .ZN(P2_U3278) );
  INV_X1 U8901 ( .A(n9259), .ZN(n7352) );
  OAI222_X1 U8902 ( .A1(n9694), .A2(n7133), .B1(n9688), .B2(n7132), .C1(
        P1_U3086), .C2(n7352), .ZN(P1_U3338) );
  OAI21_X1 U8903 ( .B1(n7134), .B2(n7135), .A(n7136), .ZN(n7142) );
  INV_X1 U8904 ( .A(n7142), .ZN(n9893) );
  NOR2_X1 U8905 ( .A1(n9718), .A2(n7137), .ZN(n8656) );
  INV_X1 U8906 ( .A(n8656), .ZN(n7148) );
  NOR2_X1 U8907 ( .A1(n9891), .A2(n9699), .ZN(n7145) );
  NAND2_X1 U8908 ( .A1(n7138), .A2(n7139), .ZN(n7140) );
  XNOR2_X1 U8909 ( .A(n7140), .B(n7135), .ZN(n7144) );
  OAI22_X1 U8910 ( .A1(n5811), .A2(n9710), .B1(n7211), .B2(n9712), .ZN(n7141)
         );
  AOI21_X1 U8911 ( .B1(n7142), .B2(n7282), .A(n7141), .ZN(n7143) );
  OAI21_X1 U8912 ( .B1(n9708), .B2(n7144), .A(n7143), .ZN(n9895) );
  AOI211_X1 U8913 ( .C1(n8805), .C2(P2_REG3_REG_2__SCAN_IN), .A(n7145), .B(
        n9895), .ZN(n7146) );
  MUX2_X1 U8914 ( .A(n6674), .B(n7146), .S(n9716), .Z(n7147) );
  OAI21_X1 U8915 ( .B1(n9893), .B2(n7148), .A(n7147), .ZN(P2_U3231) );
  INV_X1 U8916 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7149) );
  OAI22_X1 U8917 ( .A1(n8907), .A2(n7150), .B1(n7149), .B2(n9937), .ZN(n7151)
         );
  INV_X1 U8918 ( .A(n7151), .ZN(n7152) );
  OAI21_X1 U8919 ( .B1(n7153), .B2(n9939), .A(n7152), .ZN(P2_U3399) );
  INV_X1 U8920 ( .A(n7154), .ZN(n7217) );
  AOI22_X1 U8921 ( .A1(n9812), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7155), .ZN(n7156) );
  OAI21_X1 U8922 ( .B1(n7217), .B2(n9688), .A(n7156), .ZN(P1_U3337) );
  XNOR2_X1 U8923 ( .A(n7346), .B(n7342), .ZN(n7343) );
  XNOR2_X1 U8924 ( .A(n9773), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9766) );
  OAI21_X1 U8925 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7162), .A(n7157), .ZN(
        n9767) );
  NOR2_X1 U8926 ( .A1(n9766), .A2(n9767), .ZN(n9765) );
  AOI21_X1 U8927 ( .B1(n9773), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9765), .ZN(
        n9784) );
  XNOR2_X1 U8928 ( .A(n9777), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9783) );
  NOR2_X1 U8929 ( .A1(n9784), .A2(n9783), .ZN(n9782) );
  AOI21_X1 U8930 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9777), .A(n9782), .ZN(
        n7158) );
  NOR2_X1 U8931 ( .A1(n7158), .A2(n7164), .ZN(n7159) );
  XNOR2_X1 U8932 ( .A(n7164), .B(n7158), .ZN(n9797) );
  NOR2_X1 U8933 ( .A1(n9796), .A2(n9797), .ZN(n9795) );
  NOR2_X1 U8934 ( .A1(n7159), .A2(n9795), .ZN(n7344) );
  XOR2_X1 U8935 ( .A(n7343), .B(n7344), .Z(n7173) );
  NAND2_X1 U8936 ( .A1(n9773), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7160) );
  OAI21_X1 U8937 ( .B1(n9773), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7160), .ZN(
        n9769) );
  OAI21_X1 U8938 ( .B1(n7162), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7161), .ZN(
        n9770) );
  NOR2_X1 U8939 ( .A1(n9769), .A2(n9770), .ZN(n9768) );
  AOI21_X1 U8940 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9773), .A(n9768), .ZN(
        n9779) );
  NAND2_X1 U8941 ( .A1(n9777), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7163) );
  OAI21_X1 U8942 ( .B1(n9777), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7163), .ZN(
        n9780) );
  NOR2_X1 U8943 ( .A1(n9779), .A2(n9780), .ZN(n9778) );
  AOI21_X1 U8944 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9777), .A(n9778), .ZN(
        n7165) );
  NOR2_X1 U8945 ( .A1(n7165), .A2(n7164), .ZN(n7166) );
  INV_X1 U8946 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9800) );
  XOR2_X1 U8947 ( .A(n9804), .B(n7165), .Z(n9801) );
  NOR2_X1 U8948 ( .A1(n9800), .A2(n9801), .ZN(n9799) );
  NOR2_X1 U8949 ( .A1(n7166), .A2(n9799), .ZN(n7168) );
  XNOR2_X1 U8950 ( .A(n7346), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n7167) );
  AOI21_X1 U8951 ( .B1(n7168), .B2(n7167), .A(n9798), .ZN(n7171) );
  OR2_X1 U8952 ( .A1(n7168), .A2(n7167), .ZN(n7348) );
  NAND2_X1 U8953 ( .A1(n9746), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7169) );
  NAND2_X1 U8954 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9030) );
  OAI211_X1 U8955 ( .C1(n9790), .C2(n7341), .A(n7169), .B(n9030), .ZN(n7170)
         );
  AOI21_X1 U8956 ( .B1(n7171), .B2(n7348), .A(n7170), .ZN(n7172) );
  OAI21_X1 U8957 ( .B1(n7173), .B2(n9808), .A(n7172), .ZN(P1_U3259) );
  NOR2_X1 U8958 ( .A1(n7175), .A2(n7174), .ZN(n7177) );
  INV_X1 U8959 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7534) );
  OR2_X1 U8960 ( .A1(n7196), .A2(n7534), .ZN(n7242) );
  NAND2_X1 U8961 ( .A1(n7196), .A2(n7534), .ZN(n7178) );
  NAND2_X1 U8962 ( .A1(n7242), .A2(n7178), .ZN(n7180) );
  INV_X1 U8963 ( .A(n7243), .ZN(n7179) );
  AOI21_X1 U8964 ( .B1(n7181), .B2(n7180), .A(n7179), .ZN(n7203) );
  INV_X1 U8965 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7193) );
  MUX2_X1 U8966 ( .A(n7534), .B(n7193), .S(n8444), .Z(n7182) );
  NAND2_X1 U8967 ( .A1(n7182), .A2(n7196), .ZN(n7245) );
  INV_X1 U8968 ( .A(n7182), .ZN(n7183) );
  NAND2_X1 U8969 ( .A1(n7183), .A2(n7256), .ZN(n7184) );
  NAND2_X1 U8970 ( .A1(n7245), .A2(n7184), .ZN(n7185) );
  AOI21_X1 U8971 ( .B1(n7187), .B2(n7186), .A(n7185), .ZN(n7253) );
  AND3_X1 U8972 ( .A1(n7187), .A2(n7186), .A3(n7185), .ZN(n7188) );
  OAI21_X1 U8973 ( .B1(n7253), .B2(n7188), .A(n9883), .ZN(n7202) );
  NAND2_X1 U8974 ( .A1(n7190), .A2(n7189), .ZN(n7192) );
  NAND2_X1 U8975 ( .A1(n7192), .A2(n7191), .ZN(n7195) );
  MUX2_X1 U8976 ( .A(n7193), .B(P2_REG1_REG_10__SCAN_IN), .S(n7196), .Z(n7194)
         );
  NAND2_X1 U8977 ( .A1(n7194), .A2(n7195), .ZN(n7257) );
  OAI21_X1 U8978 ( .B1(n7195), .B2(n7194), .A(n7257), .ZN(n7200) );
  INV_X1 U8979 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7198) );
  INV_X1 U8980 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10128) );
  NOR2_X1 U8981 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10128), .ZN(n7596) );
  AOI21_X1 U8982 ( .B1(n8559), .B2(n7196), .A(n7596), .ZN(n7197) );
  OAI21_X1 U8983 ( .B1(n7198), .B2(n8618), .A(n7197), .ZN(n7199) );
  AOI21_X1 U8984 ( .B1(n7200), .B2(n8595), .A(n7199), .ZN(n7201) );
  OAI211_X1 U8985 ( .C1(n7203), .C2(n8642), .A(n7202), .B(n7201), .ZN(P2_U3192) );
  INV_X1 U8986 ( .A(n7204), .ZN(n7206) );
  AOI21_X1 U8987 ( .B1(n7206), .B2(n8465), .A(n7205), .ZN(n7209) );
  XNOR2_X1 U8988 ( .A(n8029), .B(n8306), .ZN(n7232) );
  XNOR2_X1 U8989 ( .A(n7232), .B(n8464), .ZN(n7208) );
  NAND2_X1 U8990 ( .A1(n7209), .A2(n7208), .ZN(n7233) );
  OAI21_X1 U8991 ( .B1(n7209), .B2(n7208), .A(n7233), .ZN(n7210) );
  NAND2_X1 U8992 ( .A1(n7210), .A2(n8179), .ZN(n7215) );
  OAI22_X1 U8993 ( .A1(n8120), .A2(n7211), .B1(n7294), .B2(n8207), .ZN(n7212)
         );
  AOI211_X1 U8994 ( .C1(n8306), .C2(n8196), .A(n7213), .B(n7212), .ZN(n7214)
         );
  OAI211_X1 U8995 ( .C1(n7216), .C2(n8183), .A(n7215), .B(n7214), .ZN(P2_U3170) );
  OAI222_X1 U8996 ( .A1(n7957), .A2(n7218), .B1(n8630), .B2(P2_U3151), .C1(
        n8964), .C2(n7217), .ZN(P2_U3277) );
  OAI21_X1 U8997 ( .B1(n7220), .B2(n7225), .A(n7219), .ZN(n7221) );
  INV_X1 U8998 ( .A(n7221), .ZN(n9626) );
  AOI211_X1 U8999 ( .C1(n9622), .C2(n7335), .A(n9510), .B(n4688), .ZN(n9621)
         );
  NOR2_X1 U9000 ( .A1(n4692), .A2(n9514), .ZN(n7224) );
  OAI22_X1 U9001 ( .A1(n9468), .A2(n7222), .B1(n7408), .B2(n9390), .ZN(n7223)
         );
  AOI211_X1 U9002 ( .C1(n9621), .C2(n9527), .A(n7224), .B(n7223), .ZN(n7231)
         );
  INV_X1 U9003 ( .A(n7357), .ZN(n7227) );
  INV_X1 U9004 ( .A(n7225), .ZN(n7819) );
  AOI21_X1 U9005 ( .B1(n7330), .B2(n7709), .A(n7819), .ZN(n7226) );
  NOR2_X1 U9006 ( .A1(n7227), .A2(n7226), .ZN(n7228) );
  OAI222_X1 U9007 ( .A1(n9516), .A2(n7229), .B1(n9380), .B2(n7411), .C1(n9518), 
        .C2(n7228), .ZN(n9620) );
  NAND2_X1 U9008 ( .A1(n9620), .A2(n9468), .ZN(n7230) );
  OAI211_X1 U9009 ( .C1(n9626), .C2(n9529), .A(n7231), .B(n7230), .ZN(P1_U3281) );
  INV_X1 U9010 ( .A(n7232), .ZN(n7234) );
  OAI21_X1 U9011 ( .B1(n7234), .B2(n8464), .A(n7233), .ZN(n7291) );
  XNOR2_X1 U9012 ( .A(n8029), .B(n7239), .ZN(n7289) );
  XNOR2_X1 U9013 ( .A(n7289), .B(n8463), .ZN(n7290) );
  XNOR2_X1 U9014 ( .A(n7291), .B(n7290), .ZN(n7235) );
  NAND2_X1 U9015 ( .A1(n7235), .A2(n8179), .ZN(n7241) );
  OAI22_X1 U9016 ( .A1(n8120), .A2(n7236), .B1(n7461), .B2(n8207), .ZN(n7237)
         );
  AOI211_X1 U9017 ( .C1(n7239), .C2(n8196), .A(n7238), .B(n7237), .ZN(n7240)
         );
  OAI211_X1 U9018 ( .C1(n7279), .C2(n8183), .A(n7241), .B(n7240), .ZN(P2_U3167) );
  AOI21_X1 U9019 ( .B1(n7247), .B2(n7244), .A(n7428), .ZN(n7266) );
  INV_X1 U9020 ( .A(n7245), .ZN(n7252) );
  MUX2_X1 U9021 ( .A(n7247), .B(n7246), .S(n8626), .Z(n7248) );
  NAND2_X1 U9022 ( .A1(n7248), .A2(n7426), .ZN(n7447) );
  INV_X1 U9023 ( .A(n7248), .ZN(n7249) );
  NAND2_X1 U9024 ( .A1(n7249), .A2(n7433), .ZN(n7250) );
  AND2_X1 U9025 ( .A1(n7447), .A2(n7250), .ZN(n7251) );
  OAI21_X1 U9026 ( .B1(n7253), .B2(n7252), .A(n7251), .ZN(n7448) );
  INV_X1 U9027 ( .A(n7448), .ZN(n7255) );
  NOR3_X1 U9028 ( .A1(n7253), .A2(n7252), .A3(n7251), .ZN(n7254) );
  OAI21_X1 U9029 ( .B1(n7255), .B2(n7254), .A(n9883), .ZN(n7265) );
  NAND2_X1 U9030 ( .A1(n7256), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7258) );
  OAI21_X1 U9031 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7259), .A(n7434), .ZN(
        n7263) );
  INV_X1 U9032 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7261) );
  INV_X1 U9033 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10126) );
  NOR2_X1 U9034 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10126), .ZN(n8163) );
  AOI21_X1 U9035 ( .B1(n8559), .B2(n7426), .A(n8163), .ZN(n7260) );
  OAI21_X1 U9036 ( .B1(n7261), .B2(n8618), .A(n7260), .ZN(n7262) );
  AOI21_X1 U9037 ( .B1(n7263), .B2(n8595), .A(n7262), .ZN(n7264) );
  OAI211_X1 U9038 ( .C1(n7266), .C2(n8642), .A(n7265), .B(n7264), .ZN(P2_U3193) );
  OAI21_X1 U9039 ( .B1(n7267), .B2(n5897), .A(n7268), .ZN(n7269) );
  AOI222_X1 U9040 ( .A1(n8817), .A2(n7269), .B1(n8462), .B2(n8822), .C1(n8460), 
        .C2(n8819), .ZN(n7416) );
  OAI22_X1 U9041 ( .A1(n8807), .A2(n7421), .B1(n7465), .B2(n9697), .ZN(n7274)
         );
  NAND3_X1 U9042 ( .A1(n7271), .A2(n5897), .A3(n8313), .ZN(n7272) );
  NAND2_X1 U9043 ( .A1(n7270), .A2(n7272), .ZN(n7417) );
  NOR2_X1 U9044 ( .A1(n7417), .A2(n8795), .ZN(n7273) );
  AOI211_X1 U9045 ( .C1(n9718), .C2(P2_REG2_REG_7__SCAN_IN), .A(n7274), .B(
        n7273), .ZN(n7275) );
  OAI21_X1 U9046 ( .B1(n7416), .B2(n9718), .A(n7275), .ZN(P2_U3226) );
  OR2_X1 U9047 ( .A1(n7277), .A2(n8248), .ZN(n7278) );
  NAND2_X1 U9048 ( .A1(n7276), .A2(n7278), .ZN(n9906) );
  OAI22_X1 U9049 ( .A1(n8807), .A2(n9903), .B1(n7279), .B2(n9697), .ZN(n7287)
         );
  INV_X1 U9050 ( .A(n8248), .ZN(n7280) );
  XNOR2_X1 U9051 ( .A(n7281), .B(n7280), .ZN(n7285) );
  NAND2_X1 U9052 ( .A1(n9906), .A2(n7282), .ZN(n7284) );
  AOI22_X1 U9053 ( .A1(n8822), .A2(n8464), .B1(n8462), .B2(n8819), .ZN(n7283)
         );
  OAI211_X1 U9054 ( .C1(n9708), .C2(n7285), .A(n7284), .B(n7283), .ZN(n9904)
         );
  MUX2_X1 U9055 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9904), .S(n9716), .Z(n7286)
         );
  AOI211_X1 U9056 ( .C1(n8656), .C2(n9906), .A(n7287), .B(n7286), .ZN(n7288)
         );
  INV_X1 U9057 ( .A(n7288), .ZN(P2_U3228) );
  XNOR2_X1 U9058 ( .A(n8029), .B(n7297), .ZN(n7457) );
  XNOR2_X1 U9059 ( .A(n7457), .B(n8462), .ZN(n7292) );
  NAND2_X1 U9060 ( .A1(n7293), .A2(n7292), .ZN(n7456) );
  OAI211_X1 U9061 ( .C1(n7293), .C2(n7292), .A(n7456), .B(n8179), .ZN(n7299)
         );
  OAI22_X1 U9062 ( .A1(n8120), .A2(n7294), .B1(n7519), .B2(n8207), .ZN(n7295)
         );
  AOI211_X1 U9063 ( .C1(n7297), .C2(n8196), .A(n7296), .B(n7295), .ZN(n7298)
         );
  OAI211_X1 U9064 ( .C1(n7317), .C2(n8183), .A(n7299), .B(n7298), .ZN(P2_U3179) );
  XNOR2_X1 U9065 ( .A(n7300), .B(n7301), .ZN(n7302) );
  NAND2_X1 U9066 ( .A1(n7302), .A2(n7303), .ZN(n7373) );
  OAI21_X1 U9067 ( .B1(n7303), .B2(n7302), .A(n7373), .ZN(n7304) );
  NAND2_X1 U9068 ( .A1(n7304), .A2(n9115), .ZN(n7311) );
  OAI22_X1 U9069 ( .A1(n9119), .A2(n7306), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7305), .ZN(n7309) );
  NOR2_X1 U9070 ( .A1(n9107), .A2(n7307), .ZN(n7308) );
  AOI211_X1 U9071 ( .C1(n9117), .C2(n9138), .A(n7309), .B(n7308), .ZN(n7310)
         );
  OAI211_X1 U9072 ( .C1(n9856), .C2(n9124), .A(n7311), .B(n7310), .ZN(P1_U3221) );
  INV_X1 U9073 ( .A(n7312), .ZN(n7314) );
  OAI222_X1 U9074 ( .A1(n9694), .A2(n7313), .B1(n9688), .B2(n7314), .C1(
        P1_U3086), .C2(n7866), .ZN(P1_U3336) );
  OAI222_X1 U9075 ( .A1(n7957), .A2(n7315), .B1(n8960), .B2(n7314), .C1(n8638), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  NAND2_X1 U9076 ( .A1(n7276), .A2(n8290), .ZN(n7316) );
  XNOR2_X1 U9077 ( .A(n7316), .B(n8249), .ZN(n9912) );
  OAI22_X1 U9078 ( .A1(n8807), .A2(n9909), .B1(n7317), .B2(n9697), .ZN(n7324)
         );
  NAND2_X1 U9079 ( .A1(n7318), .A2(n8249), .ZN(n7319) );
  NAND3_X1 U9080 ( .A1(n7320), .A2(n8817), .A3(n7319), .ZN(n7322) );
  AOI22_X1 U9081 ( .A1(n8822), .A2(n8463), .B1(n8461), .B2(n8819), .ZN(n7321)
         );
  NAND2_X1 U9082 ( .A1(n7322), .A2(n7321), .ZN(n9910) );
  MUX2_X1 U9083 ( .A(n9910), .B(P2_REG2_REG_6__SCAN_IN), .S(n9718), .Z(n7323)
         );
  AOI211_X1 U9084 ( .C1(n8830), .C2(n9912), .A(n7324), .B(n7323), .ZN(n7325)
         );
  INV_X1 U9085 ( .A(n7325), .ZN(P2_U3227) );
  XOR2_X1 U9086 ( .A(n7326), .B(n7816), .Z(n7333) );
  INV_X1 U9087 ( .A(n7333), .ZN(n9630) );
  AOI21_X1 U9088 ( .B1(n7327), .B2(n7816), .A(n9518), .ZN(n7329) );
  OAI22_X1 U9089 ( .A1(n7380), .A2(n9380), .B1(n7328), .B2(n9516), .ZN(n7511)
         );
  AOI21_X1 U9090 ( .B1(n7330), .B2(n7329), .A(n7511), .ZN(n7331) );
  OAI21_X1 U9091 ( .B1(n7333), .B2(n7332), .A(n7331), .ZN(n9628) );
  AOI21_X1 U9092 ( .B1(n7334), .B2(n9630), .A(n9628), .ZN(n7340) );
  AOI211_X1 U9093 ( .C1(n7510), .C2(n4366), .A(n9510), .B(n4693), .ZN(n9629)
         );
  NOR2_X1 U9094 ( .A1(n9677), .A2(n9514), .ZN(n7338) );
  OAI22_X1 U9095 ( .A1(n9468), .A2(n7336), .B1(n7514), .B2(n9390), .ZN(n7337)
         );
  AOI211_X1 U9096 ( .C1(n9629), .C2(n9527), .A(n7338), .B(n7337), .ZN(n7339)
         );
  OAI21_X1 U9097 ( .B1(n7340), .B2(n9826), .A(n7339), .ZN(P1_U3282) );
  XNOR2_X1 U9098 ( .A(n9259), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9260) );
  AOI22_X1 U9099 ( .A1(n7344), .A2(n7343), .B1(n7342), .B2(n7341), .ZN(n9261)
         );
  XOR2_X1 U9100 ( .A(n9260), .B(n9261), .Z(n7356) );
  INV_X1 U9101 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7345) );
  XNOR2_X1 U9102 ( .A(n9259), .B(n7345), .ZN(n7350) );
  NAND2_X1 U9103 ( .A1(n7346), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7347) );
  AND2_X1 U9104 ( .A1(n7348), .A2(n7347), .ZN(n7349) );
  NAND2_X1 U9105 ( .A1(n7349), .A2(n7350), .ZN(n9255) );
  OAI21_X1 U9106 ( .B1(n7350), .B2(n7349), .A(n9255), .ZN(n7354) );
  NAND2_X1 U9107 ( .A1(n9746), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n7351) );
  NAND2_X1 U9108 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9040) );
  OAI211_X1 U9109 ( .C1(n9790), .C2(n7352), .A(n7351), .B(n9040), .ZN(n7353)
         );
  AOI21_X1 U9110 ( .B1(n7354), .B2(n9815), .A(n7353), .ZN(n7355) );
  OAI21_X1 U9111 ( .B1(n9808), .B2(n7356), .A(n7355), .ZN(P1_U3260) );
  NAND2_X1 U9112 ( .A1(n7357), .A2(n7893), .ZN(n7358) );
  XNOR2_X1 U9113 ( .A(n7363), .B(n7358), .ZN(n7359) );
  OR2_X1 U9114 ( .A1(n7359), .A2(n9518), .ZN(n7361) );
  AOI22_X1 U9115 ( .A1(n9134), .A2(n9524), .B1(n9500), .B2(n9523), .ZN(n7360)
         );
  NAND2_X1 U9116 ( .A1(n7361), .A2(n7360), .ZN(n9615) );
  INV_X1 U9117 ( .A(n9615), .ZN(n7372) );
  OAI21_X1 U9118 ( .B1(n7364), .B2(n7363), .A(n7362), .ZN(n9617) );
  NAND2_X1 U9119 ( .A1(n9617), .A2(n9836), .ZN(n7371) );
  INV_X1 U9120 ( .A(n7471), .ZN(n7365) );
  AOI211_X1 U9121 ( .C1(n7486), .C2(n7366), .A(n9510), .B(n7365), .ZN(n9616)
         );
  INV_X1 U9122 ( .A(n7486), .ZN(n9671) );
  NOR2_X1 U9123 ( .A1(n9671), .A2(n9514), .ZN(n7369) );
  OAI22_X1 U9124 ( .A1(n9468), .A2(n7367), .B1(n7484), .B2(n9390), .ZN(n7368)
         );
  AOI211_X1 U9125 ( .C1(n9616), .C2(n9527), .A(n7369), .B(n7368), .ZN(n7370)
         );
  OAI211_X1 U9126 ( .C1(n9826), .C2(n7372), .A(n7371), .B(n7370), .ZN(P1_U3280) );
  OAI21_X1 U9127 ( .B1(n7374), .B2(n7300), .A(n7373), .ZN(n7378) );
  XNOR2_X1 U9128 ( .A(n7376), .B(n7375), .ZN(n7377) );
  XNOR2_X1 U9129 ( .A(n7378), .B(n7377), .ZN(n7387) );
  OAI21_X1 U9130 ( .B1(n9119), .B2(n7380), .A(n7379), .ZN(n7383) );
  NOR2_X1 U9131 ( .A1(n9107), .A2(n7381), .ZN(n7382) );
  AOI211_X1 U9132 ( .C1(n9117), .C2(n9137), .A(n7383), .B(n7382), .ZN(n7386)
         );
  NAND2_X1 U9133 ( .A1(n9096), .A2(n7384), .ZN(n7385) );
  OAI211_X1 U9134 ( .C1(n7387), .C2(n9098), .A(n7386), .B(n7385), .ZN(P1_U3231) );
  NAND2_X1 U9135 ( .A1(n7270), .A2(n7388), .ZN(n7389) );
  XNOR2_X1 U9136 ( .A(n7389), .B(n8251), .ZN(n9917) );
  INV_X1 U9137 ( .A(n9917), .ZN(n7397) );
  OAI211_X1 U9138 ( .C1(n7391), .C2(n8251), .A(n7390), .B(n8817), .ZN(n7393)
         );
  AOI22_X1 U9139 ( .A1(n8822), .A2(n8461), .B1(n8459), .B2(n8819), .ZN(n7392)
         );
  NAND2_X1 U9140 ( .A1(n7393), .A2(n7392), .ZN(n9915) );
  NOR2_X1 U9141 ( .A1(n9716), .A2(n6991), .ZN(n7395) );
  OAI22_X1 U9142 ( .A1(n8807), .A2(n9914), .B1(n7528), .B2(n9697), .ZN(n7394)
         );
  AOI211_X1 U9143 ( .C1(n9915), .C2(n9716), .A(n7395), .B(n7394), .ZN(n7396)
         );
  OAI21_X1 U9144 ( .B1(n7397), .B2(n8795), .A(n7396), .ZN(P2_U3225) );
  NAND2_X1 U9145 ( .A1(n7401), .A2(n7582), .ZN(n7399) );
  OAI211_X1 U9146 ( .C1(n7400), .C2(n9694), .A(n7399), .B(n7398), .ZN(P1_U3335) );
  INV_X1 U9147 ( .A(n7401), .ZN(n7403) );
  OAI222_X1 U9148 ( .A1(n8964), .A2(n7403), .B1(P2_U3151), .B2(n8423), .C1(
        n7402), .C2(n7957), .ZN(P2_U3275) );
  OAI21_X1 U9149 ( .B1(n7406), .B2(n7405), .A(n7404), .ZN(n7407) );
  NAND2_X1 U9150 ( .A1(n7407), .A2(n9115), .ZN(n7415) );
  INV_X1 U9151 ( .A(n7408), .ZN(n7413) );
  AOI21_X1 U9152 ( .B1(n9109), .B2(n9133), .A(n7409), .ZN(n7410) );
  OAI21_X1 U9153 ( .B1(n7411), .B2(n9083), .A(n7410), .ZN(n7412) );
  AOI21_X1 U9154 ( .B1(n7413), .B2(n9121), .A(n7412), .ZN(n7414) );
  OAI211_X1 U9155 ( .C1(n4692), .C2(n9124), .A(n7415), .B(n7414), .ZN(P1_U3224) );
  INV_X1 U9156 ( .A(n9933), .ZN(n9920) );
  OAI21_X1 U9157 ( .B1(n9920), .B2(n7417), .A(n7416), .ZN(n7423) );
  OAI22_X1 U9158 ( .A1(n8855), .A2(n7421), .B1(n9950), .B2(n6885), .ZN(n7418)
         );
  AOI21_X1 U9159 ( .B1(n7423), .B2(n9950), .A(n7418), .ZN(n7419) );
  INV_X1 U9160 ( .A(n7419), .ZN(P2_U3466) );
  INV_X1 U9161 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7420) );
  OAI22_X1 U9162 ( .A1(n8907), .A2(n7421), .B1(n7420), .B2(n9937), .ZN(n7422)
         );
  AOI21_X1 U9163 ( .B1(n7423), .B2(n9937), .A(n7422), .ZN(n7424) );
  INV_X1 U9164 ( .A(n7424), .ZN(P2_U3411) );
  NOR2_X1 U9165 ( .A1(n7426), .A2(n7425), .ZN(n7427) );
  INV_X1 U9166 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8467) );
  MUX2_X1 U9167 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8467), .S(n8483), .Z(n7430)
         );
  INV_X1 U9168 ( .A(n8469), .ZN(n7429) );
  AOI21_X1 U9169 ( .B1(n7431), .B2(n7430), .A(n7429), .ZN(n7455) );
  NAND2_X1 U9170 ( .A1(n7433), .A2(n7432), .ZN(n7435) );
  INV_X1 U9171 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7441) );
  MUX2_X1 U9172 ( .A(n7441), .B(P2_REG1_REG_12__SCAN_IN), .S(n8483), .Z(n7436)
         );
  NAND2_X1 U9173 ( .A1(n7437), .A2(n7436), .ZN(n8482) );
  OAI21_X1 U9174 ( .B1(n7437), .B2(n7436), .A(n8482), .ZN(n7453) );
  INV_X1 U9175 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7440) );
  NOR2_X1 U9176 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7438), .ZN(n7616) );
  AOI21_X1 U9177 ( .B1(n8559), .B2(n8483), .A(n7616), .ZN(n7439) );
  OAI21_X1 U9178 ( .B1(n7440), .B2(n8618), .A(n7439), .ZN(n7452) );
  MUX2_X1 U9179 ( .A(n8467), .B(n7441), .S(n8444), .Z(n7442) );
  NAND2_X1 U9180 ( .A1(n7442), .A2(n8483), .ZN(n8472) );
  INV_X1 U9181 ( .A(n7442), .ZN(n7444) );
  NAND2_X1 U9182 ( .A1(n7444), .A2(n7443), .ZN(n7445) );
  NAND2_X1 U9183 ( .A1(n8472), .A2(n7445), .ZN(n7446) );
  AOI21_X1 U9184 ( .B1(n7448), .B2(n7447), .A(n7446), .ZN(n8479) );
  INV_X1 U9185 ( .A(n8479), .ZN(n7450) );
  NAND3_X1 U9186 ( .A1(n7448), .A2(n7447), .A3(n7446), .ZN(n7449) );
  AOI21_X1 U9187 ( .B1(n7450), .B2(n7449), .A(n8591), .ZN(n7451) );
  AOI211_X1 U9188 ( .C1(n8595), .C2(n7453), .A(n7452), .B(n7451), .ZN(n7454)
         );
  OAI21_X1 U9189 ( .B1(n7455), .B2(n8642), .A(n7454), .ZN(P2_U3194) );
  XNOR2_X1 U9190 ( .A(n8029), .B(n7464), .ZN(n7518) );
  XOR2_X1 U9191 ( .A(n8461), .B(n7518), .Z(n7460) );
  INV_X1 U9192 ( .A(n7521), .ZN(n7458) );
  AOI21_X1 U9193 ( .B1(n7460), .B2(n7459), .A(n7458), .ZN(n7469) );
  OAI22_X1 U9194 ( .A1(n8120), .A2(n7461), .B1(n7538), .B2(n8207), .ZN(n7462)
         );
  AOI211_X1 U9195 ( .C1(n7464), .C2(n8196), .A(n7463), .B(n7462), .ZN(n7468)
         );
  INV_X1 U9196 ( .A(n7465), .ZN(n7466) );
  NAND2_X1 U9197 ( .A1(n8210), .A2(n7466), .ZN(n7467) );
  OAI211_X1 U9198 ( .C1(n7469), .C2(n8199), .A(n7468), .B(n7467), .ZN(P2_U3153) );
  XNOR2_X1 U9199 ( .A(n7470), .B(n7821), .ZN(n9614) );
  AOI211_X1 U9200 ( .C1(n9611), .C2(n7471), .A(n9510), .B(n9508), .ZN(n9610)
         );
  AOI22_X1 U9201 ( .A1(n9826), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8981), .B2(
        n9834), .ZN(n7472) );
  OAI21_X1 U9202 ( .B1(n8978), .B2(n9514), .A(n7472), .ZN(n7476) );
  OAI21_X1 U9203 ( .B1(n7821), .B2(n4427), .A(n7473), .ZN(n7474) );
  AOI222_X1 U9204 ( .A1(n9503), .A2(n7474), .B1(n9499), .B2(n9500), .C1(n9133), 
        .C2(n9524), .ZN(n9613) );
  NOR2_X1 U9205 ( .A1(n9613), .A2(n9826), .ZN(n7475) );
  AOI211_X1 U9206 ( .C1(n9610), .C2(n9527), .A(n7476), .B(n7475), .ZN(n7477)
         );
  OAI21_X1 U9207 ( .B1(n9614), .B2(n9529), .A(n7477), .ZN(P1_U3279) );
  AOI21_X1 U9208 ( .B1(n7480), .B2(n7479), .A(n7478), .ZN(n7488) );
  NAND2_X1 U9209 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9774) );
  OAI21_X1 U9210 ( .B1(n9119), .B2(n7481), .A(n9774), .ZN(n7482) );
  AOI21_X1 U9211 ( .B1(n9117), .B2(n9134), .A(n7482), .ZN(n7483) );
  OAI21_X1 U9212 ( .B1(n9107), .B2(n7484), .A(n7483), .ZN(n7485) );
  AOI21_X1 U9213 ( .B1(n7486), .B2(n9096), .A(n7485), .ZN(n7487) );
  OAI21_X1 U9214 ( .B1(n7488), .B2(n9098), .A(n7487), .ZN(P1_U3234) );
  INV_X1 U9215 ( .A(n7489), .ZN(n7501) );
  OAI222_X1 U9216 ( .A1(n8964), .A2(n7501), .B1(P2_U3151), .B2(n8269), .C1(
        n7490), .C2(n7957), .ZN(P2_U3274) );
  OAI21_X1 U9217 ( .B1(n7491), .B2(n8252), .A(n7492), .ZN(n7493) );
  AOI222_X1 U9218 ( .A1(n8817), .A2(n7493), .B1(n8460), .B2(n8822), .C1(n8458), 
        .C2(n8819), .ZN(n7574) );
  NAND2_X1 U9219 ( .A1(n7494), .A2(n8252), .ZN(n7495) );
  AND2_X1 U9220 ( .A1(n7529), .A2(n7495), .ZN(n7576) );
  NOR2_X1 U9221 ( .A1(n8807), .A2(n7581), .ZN(n7498) );
  OAI22_X1 U9222 ( .A1(n9716), .A2(n7496), .B1(n7550), .B2(n9697), .ZN(n7497)
         );
  AOI211_X1 U9223 ( .C1(n7576), .C2(n8830), .A(n7498), .B(n7497), .ZN(n7499)
         );
  OAI21_X1 U9224 ( .B1(n7574), .B2(n9718), .A(n7499), .ZN(P2_U3224) );
  OAI222_X1 U9225 ( .A1(P1_U3086), .A2(n7798), .B1(n9688), .B2(n7501), .C1(
        n7500), .C2(n9694), .ZN(P1_U3334) );
  AOI21_X1 U9226 ( .B1(n7504), .B2(n7503), .A(n7502), .ZN(n7509) );
  OAI21_X1 U9227 ( .B1(n7507), .B2(n7506), .A(n7505), .ZN(n7508) );
  XNOR2_X1 U9228 ( .A(n7509), .B(n7508), .ZN(n7516) );
  NAND2_X1 U9229 ( .A1(n7510), .A2(n9096), .ZN(n7513) );
  AOI22_X1 U9230 ( .A1(n9060), .A2(n7511), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n7512) );
  OAI211_X1 U9231 ( .C1(n9107), .C2(n7514), .A(n7513), .B(n7512), .ZN(n7515)
         );
  AOI21_X1 U9232 ( .B1(n7516), .B2(n9115), .A(n7515), .ZN(n7517) );
  INV_X1 U9233 ( .A(n7517), .ZN(P1_U3236) );
  XNOR2_X1 U9234 ( .A(n8029), .B(n7525), .ZN(n7539) );
  XNOR2_X1 U9235 ( .A(n7539), .B(n8460), .ZN(n7541) );
  XNOR2_X1 U9236 ( .A(n7542), .B(n7541), .ZN(n7522) );
  NAND2_X1 U9237 ( .A1(n7522), .A2(n8179), .ZN(n7527) );
  OAI22_X1 U9238 ( .A1(n8120), .A2(n7519), .B1(n7592), .B2(n8207), .ZN(n7523)
         );
  AOI211_X1 U9239 ( .C1(n7525), .C2(n8196), .A(n7524), .B(n7523), .ZN(n7526)
         );
  OAI211_X1 U9240 ( .C1(n7528), .C2(n8183), .A(n7527), .B(n7526), .ZN(P2_U3161) );
  NAND2_X1 U9241 ( .A1(n7529), .A2(n8299), .ZN(n7531) );
  INV_X1 U9242 ( .A(n7530), .ZN(n8255) );
  XNOR2_X1 U9243 ( .A(n7531), .B(n8255), .ZN(n9921) );
  XNOR2_X1 U9244 ( .A(n7532), .B(n8255), .ZN(n7533) );
  OAI222_X1 U9245 ( .A1(n9710), .A2(n7592), .B1(n9712), .B2(n7607), .C1(n9708), 
        .C2(n7533), .ZN(n9923) );
  NAND2_X1 U9246 ( .A1(n9923), .A2(n9716), .ZN(n7537) );
  INV_X1 U9247 ( .A(n9919), .ZN(n7597) );
  OAI22_X1 U9248 ( .A1(n9716), .A2(n7534), .B1(n7598), .B2(n9697), .ZN(n7535)
         );
  AOI21_X1 U9249 ( .B1(n8792), .B2(n7597), .A(n7535), .ZN(n7536) );
  OAI211_X1 U9250 ( .C1(n8795), .C2(n9921), .A(n7537), .B(n7536), .ZN(P2_U3223) );
  AND2_X1 U9251 ( .A1(n7539), .A2(n7538), .ZN(n7540) );
  XNOR2_X1 U9252 ( .A(n8029), .B(n7543), .ZN(n7593) );
  XNOR2_X1 U9253 ( .A(n7593), .B(n8459), .ZN(n7544) );
  OAI211_X1 U9254 ( .C1(n7545), .C2(n7544), .A(n7595), .B(n8179), .ZN(n7549)
         );
  OAI22_X1 U9255 ( .A1(n8213), .A2(n7581), .B1(n7557), .B2(n8207), .ZN(n7546)
         );
  AOI211_X1 U9256 ( .C1(n8205), .C2(n8460), .A(n7547), .B(n7546), .ZN(n7548)
         );
  OAI211_X1 U9257 ( .C1(n7550), .C2(n8183), .A(n7549), .B(n7548), .ZN(P2_U3171) );
  INV_X1 U9258 ( .A(n7551), .ZN(n7554) );
  OAI222_X1 U9259 ( .A1(n7957), .A2(n7553), .B1(n8960), .B2(n7554), .C1(n7552), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9260 ( .A1(n9694), .A2(n7555), .B1(n9688), .B2(n7554), .C1(
        P1_U3086), .C2(n7795), .ZN(P1_U3333) );
  XNOR2_X1 U9261 ( .A(n9702), .B(n8256), .ZN(n7556) );
  OAI222_X1 U9262 ( .A1(n9710), .A2(n7557), .B1(n9712), .B2(n8167), .C1(n9708), 
        .C2(n7556), .ZN(n9927) );
  INV_X1 U9263 ( .A(n9927), .ZN(n7563) );
  OAI21_X1 U9264 ( .B1(n7559), .B2(n8256), .A(n7558), .ZN(n9929) );
  INV_X1 U9265 ( .A(n8164), .ZN(n9926) );
  NOR2_X1 U9266 ( .A1(n8807), .A2(n9926), .ZN(n7561) );
  OAI22_X1 U9267 ( .A1(n9716), .A2(n7247), .B1(n8165), .B2(n9697), .ZN(n7560)
         );
  AOI211_X1 U9268 ( .C1(n9929), .C2(n8830), .A(n7561), .B(n7560), .ZN(n7562)
         );
  OAI21_X1 U9269 ( .B1(n7563), .B2(n9718), .A(n7562), .ZN(P2_U3222) );
  OR2_X1 U9270 ( .A1(n9702), .A2(n7564), .ZN(n7566) );
  NAND2_X1 U9271 ( .A1(n7566), .A2(n7565), .ZN(n8812) );
  XNOR2_X1 U9272 ( .A(n8812), .B(n8328), .ZN(n7569) );
  NAND2_X1 U9273 ( .A1(n8456), .A2(n8819), .ZN(n7567) );
  OAI21_X1 U9274 ( .B1(n7607), .B2(n9710), .A(n7567), .ZN(n7568) );
  AOI21_X1 U9275 ( .B1(n7569), .B2(n8817), .A(n7568), .ZN(n9936) );
  XNOR2_X1 U9276 ( .A(n7570), .B(n8328), .ZN(n9934) );
  INV_X1 U9277 ( .A(n9931), .ZN(n7623) );
  NOR2_X1 U9278 ( .A1(n8807), .A2(n7623), .ZN(n7572) );
  OAI22_X1 U9279 ( .A1(n9716), .A2(n8467), .B1(n7615), .B2(n9697), .ZN(n7571)
         );
  AOI211_X1 U9280 ( .C1(n9934), .C2(n8830), .A(n7572), .B(n7571), .ZN(n7573)
         );
  OAI21_X1 U9281 ( .B1(n9936), .B2(n9718), .A(n7573), .ZN(P2_U3221) );
  INV_X1 U9282 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7577) );
  INV_X1 U9283 ( .A(n7574), .ZN(n7575) );
  AOI21_X1 U9284 ( .B1(n7576), .B2(n9933), .A(n7575), .ZN(n7579) );
  MUX2_X1 U9285 ( .A(n7577), .B(n7579), .S(n9937), .Z(n7578) );
  OAI21_X1 U9286 ( .B1(n7581), .B2(n8907), .A(n7578), .ZN(P2_U3417) );
  MUX2_X1 U9287 ( .A(n7093), .B(n7579), .S(n9950), .Z(n7580) );
  OAI21_X1 U9288 ( .B1(n7581), .B2(n8855), .A(n7580), .ZN(P2_U3468) );
  NAND2_X1 U9289 ( .A1(n7585), .A2(n7582), .ZN(n7583) );
  OAI211_X1 U9290 ( .C1(n7584), .C2(n9694), .A(n7583), .B(n7931), .ZN(P1_U3332) );
  NAND2_X1 U9291 ( .A1(n7585), .A2(n8969), .ZN(n7587) );
  NAND2_X1 U9292 ( .A1(n7586), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8450) );
  OAI211_X1 U9293 ( .C1(n7588), .C2(n7957), .A(n7587), .B(n8450), .ZN(P2_U3272) );
  INV_X1 U9294 ( .A(n7589), .ZN(n7625) );
  OAI222_X1 U9295 ( .A1(n7591), .A2(P1_U3086), .B1(n9688), .B2(n7625), .C1(
        n7590), .C2(n9694), .ZN(P1_U3331) );
  XNOR2_X1 U9296 ( .A(n8157), .B(n8458), .ZN(n8159) );
  XNOR2_X1 U9297 ( .A(n8029), .B(n9919), .ZN(n8158) );
  XNOR2_X1 U9298 ( .A(n8159), .B(n8158), .ZN(n7605) );
  AOI21_X1 U9299 ( .B1(n8205), .B2(n8459), .A(n7596), .ZN(n7603) );
  NAND2_X1 U9300 ( .A1(n8196), .A2(n7597), .ZN(n7602) );
  INV_X1 U9301 ( .A(n7598), .ZN(n7599) );
  NAND2_X1 U9302 ( .A1(n8210), .A2(n7599), .ZN(n7601) );
  OR2_X1 U9303 ( .A1(n8207), .A2(n7607), .ZN(n7600) );
  NAND4_X1 U9304 ( .A1(n7603), .A2(n7602), .A3(n7601), .A4(n7600), .ZN(n7604)
         );
  AOI21_X1 U9305 ( .B1(n7605), .B2(n8179), .A(n7604), .ZN(n7606) );
  INV_X1 U9306 ( .A(n7606), .ZN(P2_U3157) );
  XNOR2_X1 U9307 ( .A(n8029), .B(n8164), .ZN(n8160) );
  NAND2_X1 U9308 ( .A1(n8160), .A2(n7607), .ZN(n7609) );
  AOI21_X1 U9309 ( .B1(n8158), .B2(n8458), .A(n8457), .ZN(n7611) );
  NAND3_X1 U9310 ( .A1(n8158), .A2(n8458), .A3(n8457), .ZN(n7610) );
  XNOR2_X1 U9311 ( .A(n9931), .B(n8029), .ZN(n7973) );
  XNOR2_X1 U9312 ( .A(n7973), .B(n8821), .ZN(n7613) );
  NAND2_X1 U9313 ( .A1(n7614), .A2(n7613), .ZN(n7975) );
  OAI211_X1 U9314 ( .C1(n7614), .C2(n7613), .A(n7975), .B(n8179), .ZN(n7622)
         );
  INV_X1 U9315 ( .A(n7615), .ZN(n7620) );
  NAND2_X1 U9316 ( .A1(n8205), .A2(n8457), .ZN(n7618) );
  INV_X1 U9317 ( .A(n7616), .ZN(n7617) );
  OAI211_X1 U9318 ( .C1(n9709), .C2(n8207), .A(n7618), .B(n7617), .ZN(n7619)
         );
  AOI21_X1 U9319 ( .B1(n7620), .B2(n8210), .A(n7619), .ZN(n7621) );
  OAI211_X1 U9320 ( .C1(n7623), .C2(n8213), .A(n7622), .B(n7621), .ZN(P2_U3164) );
  OAI222_X1 U9321 ( .A1(n8964), .A2(n7625), .B1(P2_U3151), .B2(n6145), .C1(
        n7624), .C2(n7957), .ZN(P2_U3271) );
  INV_X1 U9322 ( .A(n7626), .ZN(n7636) );
  OAI222_X1 U9323 ( .A1(n7628), .A2(P1_U3086), .B1(n9688), .B2(n7636), .C1(
        n7627), .C2(n9694), .ZN(P1_U3330) );
  INV_X1 U9324 ( .A(n7629), .ZN(n7633) );
  OAI222_X1 U9325 ( .A1(n8964), .A2(n7633), .B1(P2_U3151), .B2(n7631), .C1(
        n7630), .C2(n7957), .ZN(P2_U3269) );
  OAI222_X1 U9326 ( .A1(n7634), .A2(P1_U3086), .B1(n9688), .B2(n7633), .C1(
        n7632), .C2(n9694), .ZN(P1_U3329) );
  OAI222_X1 U9327 ( .A1(n8964), .A2(n7636), .B1(P2_U3151), .B2(n6148), .C1(
        n7635), .C2(n7957), .ZN(P2_U3270) );
  OR2_X1 U9328 ( .A1(n7638), .A2(n7637), .ZN(n7639) );
  INV_X1 U9329 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8217) );
  INV_X1 U9330 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7972) );
  MUX2_X1 U9331 ( .A(n8217), .B(n7972), .S(n6389), .Z(n7642) );
  INV_X1 U9332 ( .A(SI_30_), .ZN(n7641) );
  NAND2_X1 U9333 ( .A1(n7642), .A2(n7641), .ZN(n7645) );
  INV_X1 U9334 ( .A(n7642), .ZN(n7643) );
  NAND2_X1 U9335 ( .A1(n7643), .A2(SI_30_), .ZN(n7644) );
  NAND2_X1 U9336 ( .A1(n7645), .A2(n7644), .ZN(n7779) );
  OAI21_X1 U9337 ( .B1(n7780), .B2(n7779), .A(n7645), .ZN(n7649) );
  MUX2_X1 U9338 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6389), .Z(n7647) );
  INV_X1 U9339 ( .A(SI_31_), .ZN(n7646) );
  XNOR2_X1 U9340 ( .A(n7647), .B(n7646), .ZN(n7648) );
  XNOR2_X1 U9341 ( .A(n7649), .B(n7648), .ZN(n8954) );
  INV_X1 U9342 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9684) );
  OR2_X1 U9343 ( .A1(n7782), .A2(n9684), .ZN(n7650) );
  INV_X1 U9344 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n7654) );
  NAND2_X1 U9345 ( .A1(n7651), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7653) );
  NAND2_X1 U9346 ( .A1(n5073), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7652) );
  OAI211_X1 U9347 ( .C1(n7655), .C2(n7654), .A(n7653), .B(n7652), .ZN(n9125)
         );
  INV_X1 U9348 ( .A(n7790), .ZN(n7786) );
  OR2_X1 U9349 ( .A1(n9304), .A2(n7786), .ZN(n7656) );
  OAI22_X1 U9350 ( .A1(n9322), .A2(n7656), .B1(n9315), .B2(n7786), .ZN(n7660)
         );
  NAND2_X1 U9351 ( .A1(n9304), .A2(n7786), .ZN(n7766) );
  OAI21_X1 U9352 ( .B1(n9127), .B2(n7766), .A(n9322), .ZN(n7659) );
  NOR2_X1 U9353 ( .A1(n7656), .A2(n9315), .ZN(n7657) );
  OR2_X1 U9354 ( .A1(n9322), .A2(n7657), .ZN(n7658) );
  AOI22_X1 U9355 ( .A1(n4699), .A2(n7660), .B1(n7659), .B2(n7658), .ZN(n7773)
         );
  NAND2_X1 U9356 ( .A1(n7751), .A2(n7661), .ZN(n7832) );
  AND2_X1 U9357 ( .A1(n9362), .A2(n7662), .ZN(n7838) );
  INV_X1 U9358 ( .A(n7838), .ZN(n7663) );
  MUX2_X1 U9359 ( .A(n7832), .B(n7663), .S(n7790), .Z(n7753) );
  NAND2_X1 U9360 ( .A1(n9582), .A2(n7664), .ZN(n7667) );
  AND2_X1 U9361 ( .A1(n7749), .A2(n7667), .ZN(n7840) );
  INV_X1 U9362 ( .A(n9587), .ZN(n9452) );
  NAND2_X1 U9363 ( .A1(n7667), .A2(n9452), .ZN(n7665) );
  NAND2_X1 U9364 ( .A1(n7665), .A2(n7790), .ZN(n7666) );
  NAND3_X1 U9365 ( .A1(n7666), .A2(n7745), .A3(n7744), .ZN(n7669) );
  NAND3_X1 U9366 ( .A1(n7667), .A2(n9132), .A3(n7790), .ZN(n7668) );
  AND2_X1 U9367 ( .A1(n7669), .A2(n7668), .ZN(n7748) );
  INV_X1 U9368 ( .A(n7748), .ZN(n7738) );
  INV_X1 U9369 ( .A(n7670), .ZN(n7673) );
  OAI21_X1 U9370 ( .B1(n7671), .B2(n7692), .A(n7881), .ZN(n7672) );
  MUX2_X1 U9371 ( .A(n7673), .B(n7672), .S(n7786), .Z(n7693) );
  INV_X1 U9372 ( .A(n7883), .ZN(n7676) );
  AND2_X1 U9373 ( .A1(n7675), .A2(n7674), .ZN(n7699) );
  OAI21_X1 U9374 ( .B1(n7693), .B2(n7676), .A(n7699), .ZN(n7691) );
  AND2_X1 U9375 ( .A1(n7678), .A2(n7677), .ZN(n7684) );
  INV_X1 U9376 ( .A(n7684), .ZN(n7680) );
  NAND2_X1 U9377 ( .A1(n7694), .A2(n7786), .ZN(n7679) );
  NOR2_X1 U9378 ( .A1(n7680), .A2(n7679), .ZN(n7690) );
  NAND2_X1 U9379 ( .A1(n7697), .A2(n7790), .ZN(n7688) );
  NAND2_X1 U9380 ( .A1(n7701), .A2(n7681), .ZN(n7682) );
  NAND2_X1 U9381 ( .A1(n7682), .A2(n7786), .ZN(n7687) );
  NAND2_X1 U9382 ( .A1(n7683), .A2(n7790), .ZN(n7686) );
  NAND3_X1 U9383 ( .A1(n7684), .A2(n7786), .A3(n7696), .ZN(n7685) );
  NAND4_X1 U9384 ( .A1(n7688), .A2(n7687), .A3(n7686), .A4(n7685), .ZN(n7689)
         );
  OAI21_X1 U9385 ( .B1(n7693), .B2(n7692), .A(n7883), .ZN(n7700) );
  NAND2_X1 U9386 ( .A1(n7694), .A2(n7790), .ZN(n7695) );
  OR3_X1 U9387 ( .A1(n7697), .A2(n7696), .A3(n7695), .ZN(n7698) );
  INV_X1 U9388 ( .A(n7701), .ZN(n7702) );
  OAI21_X1 U9389 ( .B1(n7708), .B2(n7702), .A(n7885), .ZN(n7703) );
  AND2_X1 U9390 ( .A1(n7710), .A2(n7707), .ZN(n7891) );
  NAND2_X1 U9391 ( .A1(n7703), .A2(n7891), .ZN(n7705) );
  AND2_X1 U9392 ( .A1(n7711), .A2(n7709), .ZN(n7889) );
  INV_X1 U9393 ( .A(n7893), .ZN(n7704) );
  AOI21_X1 U9394 ( .B1(n7705), .B2(n7889), .A(n7704), .ZN(n7716) );
  AND2_X1 U9395 ( .A1(n7893), .A2(n7710), .ZN(n7713) );
  INV_X1 U9396 ( .A(n7711), .ZN(n7712) );
  AOI21_X1 U9397 ( .B1(n7714), .B2(n7713), .A(n7712), .ZN(n7715) );
  MUX2_X1 U9398 ( .A(n7716), .B(n7715), .S(n7786), .Z(n7724) );
  INV_X1 U9399 ( .A(n7724), .ZN(n7717) );
  AND2_X1 U9400 ( .A1(n7728), .A2(n7722), .ZN(n7875) );
  NAND3_X1 U9401 ( .A1(n7717), .A2(n7875), .A3(n7894), .ZN(n7720) );
  NAND2_X1 U9402 ( .A1(n7725), .A2(n7721), .ZN(n7718) );
  NAND2_X1 U9403 ( .A1(n7875), .A2(n7718), .ZN(n7719) );
  AND3_X1 U9404 ( .A1(n7730), .A2(n7726), .A3(n7719), .ZN(n7900) );
  INV_X1 U9405 ( .A(n7732), .ZN(n7898) );
  AOI21_X1 U9406 ( .B1(n7720), .B2(n7900), .A(n7898), .ZN(n7733) );
  INV_X1 U9407 ( .A(n7721), .ZN(n7723) );
  OAI211_X1 U9408 ( .C1(n7724), .C2(n7723), .A(n7722), .B(n7894), .ZN(n7727)
         );
  NAND3_X1 U9409 ( .A1(n7727), .A2(n7726), .A3(n7725), .ZN(n7729) );
  NAND2_X1 U9410 ( .A1(n7729), .A2(n7728), .ZN(n7731) );
  INV_X1 U9411 ( .A(n7734), .ZN(n7741) );
  NAND2_X1 U9412 ( .A1(n7741), .A2(n7735), .ZN(n7823) );
  AND2_X1 U9413 ( .A1(n7743), .A2(n7735), .ZN(n7874) );
  NAND2_X1 U9414 ( .A1(n4377), .A2(n7874), .ZN(n7736) );
  NAND3_X1 U9415 ( .A1(n7736), .A2(n7904), .A3(n7742), .ZN(n7737) );
  NAND2_X1 U9416 ( .A1(n7738), .A2(n7737), .ZN(n7739) );
  NAND2_X1 U9417 ( .A1(n7840), .A2(n7739), .ZN(n7740) );
  NOR2_X1 U9418 ( .A1(n9422), .A2(n9084), .ZN(n7841) );
  INV_X1 U9419 ( .A(n7841), .ZN(n7746) );
  AND2_X1 U9420 ( .A1(n7742), .A2(n7741), .ZN(n7901) );
  NAND2_X1 U9421 ( .A1(n7744), .A2(n7743), .ZN(n7873) );
  AOI21_X1 U9422 ( .B1(n4377), .B2(n7901), .A(n7873), .ZN(n7747) );
  AND2_X1 U9423 ( .A1(n7746), .A2(n7745), .ZN(n7872) );
  OAI21_X1 U9424 ( .B1(n7748), .B2(n7747), .A(n7872), .ZN(n7750) );
  MUX2_X1 U9425 ( .A(n9362), .B(n7751), .S(n7790), .Z(n7752) );
  MUX2_X1 U9426 ( .A(n7834), .B(n7839), .S(n7790), .Z(n7754) );
  NAND2_X1 U9427 ( .A1(n7755), .A2(n7754), .ZN(n7763) );
  INV_X1 U9428 ( .A(n7761), .ZN(n7756) );
  OAI21_X1 U9429 ( .B1(n7763), .B2(n7756), .A(n7760), .ZN(n7757) );
  NAND2_X1 U9430 ( .A1(n7757), .A2(n7845), .ZN(n7758) );
  NAND2_X1 U9431 ( .A1(n7758), .A2(n7910), .ZN(n7759) );
  NAND4_X1 U9432 ( .A1(n7759), .A2(n7854), .A3(n7786), .A4(n7916), .ZN(n7772)
         );
  AND2_X1 U9433 ( .A1(n7910), .A2(n7790), .ZN(n7765) );
  INV_X1 U9434 ( .A(n7760), .ZN(n7844) );
  NAND2_X1 U9435 ( .A1(n7845), .A2(n7761), .ZN(n7837) );
  INV_X1 U9436 ( .A(n7837), .ZN(n7762) );
  OAI21_X1 U9437 ( .B1(n7844), .B2(n7763), .A(n7762), .ZN(n7764) );
  NAND4_X1 U9438 ( .A1(n7852), .A2(n7765), .A3(n7851), .A4(n7764), .ZN(n7771)
         );
  INV_X1 U9439 ( .A(n7766), .ZN(n7767) );
  NAND2_X1 U9440 ( .A1(n9322), .A2(n7767), .ZN(n7768) );
  OAI21_X1 U9441 ( .B1(n7790), .B2(n9127), .A(n7768), .ZN(n7769) );
  NAND2_X1 U9442 ( .A1(n7769), .A2(n9536), .ZN(n7770) );
  NAND4_X1 U9443 ( .A1(n7773), .A2(n7772), .A3(n7771), .A4(n7770), .ZN(n7777)
         );
  INV_X1 U9444 ( .A(n7858), .ZN(n7775) );
  INV_X1 U9445 ( .A(n7855), .ZN(n7774) );
  MUX2_X1 U9446 ( .A(n7775), .B(n7774), .S(n7790), .Z(n7776) );
  AOI21_X1 U9447 ( .B1(n7778), .B2(n7777), .A(n7776), .ZN(n7793) );
  NAND2_X1 U9448 ( .A1(n8216), .A2(n7781), .ZN(n7784) );
  OR2_X1 U9449 ( .A1(n7782), .A2(n7972), .ZN(n7783) );
  INV_X1 U9450 ( .A(n9638), .ZN(n9274) );
  INV_X1 U9451 ( .A(n9125), .ZN(n7785) );
  AOI22_X1 U9452 ( .A1(n7830), .A2(n9274), .B1(n7785), .B2(n7956), .ZN(n7792)
         );
  INV_X1 U9453 ( .A(n9126), .ZN(n7857) );
  OR2_X1 U9454 ( .A1(n7945), .A2(n7857), .ZN(n7922) );
  NOR2_X1 U9455 ( .A1(n9638), .A2(n7922), .ZN(n7862) );
  NOR3_X1 U9456 ( .A1(n7956), .A2(n9125), .A3(n7790), .ZN(n7789) );
  NAND3_X1 U9457 ( .A1(n7945), .A2(n7857), .A3(n7786), .ZN(n7787) );
  AOI21_X1 U9458 ( .B1(n9125), .B2(n7787), .A(n9638), .ZN(n7788) );
  AOI211_X1 U9459 ( .C1(n7862), .C2(n7790), .A(n7789), .B(n7788), .ZN(n7791)
         );
  INV_X1 U9460 ( .A(n7800), .ZN(n7794) );
  AOI21_X1 U9461 ( .B1(n7921), .B2(n9269), .A(n7794), .ZN(n7943) );
  INV_X1 U9462 ( .A(n7795), .ZN(n7799) );
  NOR2_X1 U9463 ( .A1(n7931), .A2(n7799), .ZN(n7937) );
  INV_X1 U9464 ( .A(n7796), .ZN(n7797) );
  OAI211_X1 U9465 ( .C1(n7925), .C2(n7866), .A(n7937), .B(n7797), .ZN(n7942)
         );
  INV_X1 U9466 ( .A(n9443), .ZN(n7825) );
  INV_X1 U9467 ( .A(n7801), .ZN(n9456) );
  INV_X1 U9468 ( .A(n7802), .ZN(n7813) );
  NOR2_X1 U9469 ( .A1(n7803), .A2(n4976), .ZN(n7809) );
  INV_X1 U9470 ( .A(n7804), .ZN(n7808) );
  NAND4_X1 U9471 ( .A1(n7809), .A2(n7808), .A3(n7807), .A4(n7806), .ZN(n7811)
         );
  NOR2_X1 U9472 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  NAND4_X1 U9473 ( .A1(n7815), .A2(n7814), .A3(n7813), .A4(n7812), .ZN(n7817)
         );
  NOR2_X1 U9474 ( .A1(n7817), .A2(n7816), .ZN(n7818) );
  NAND4_X1 U9475 ( .A1(n7821), .A2(n7820), .A3(n7819), .A4(n7818), .ZN(n7822)
         );
  NOR4_X1 U9476 ( .A1(n7823), .A2(n9489), .A3(n9520), .A4(n7822), .ZN(n7824)
         );
  AND4_X1 U9477 ( .A1(n9430), .A2(n7825), .A3(n9456), .A4(n7824), .ZN(n7826)
         );
  AND4_X1 U9478 ( .A1(n9387), .A2(n9406), .A3(n7826), .A4(n4509), .ZN(n7827)
         );
  NAND2_X1 U9479 ( .A1(n9368), .A2(n7827), .ZN(n7828) );
  NOR2_X1 U9480 ( .A1(n9346), .A2(n7828), .ZN(n7829) );
  NAND2_X1 U9481 ( .A1(n7832), .A2(n9362), .ZN(n7833) );
  NAND2_X1 U9482 ( .A1(n7834), .A2(n7833), .ZN(n7835) );
  AND2_X1 U9483 ( .A1(n7835), .A2(n7839), .ZN(n7836) );
  OR2_X1 U9484 ( .A1(n7837), .A2(n7836), .ZN(n7912) );
  OAI211_X1 U9485 ( .C1(n7841), .C2(n7840), .A(n7839), .B(n7838), .ZN(n7842)
         );
  INV_X1 U9486 ( .A(n7842), .ZN(n7843) );
  OR2_X1 U9487 ( .A1(n7912), .A2(n7843), .ZN(n7847) );
  NAND2_X1 U9488 ( .A1(n7845), .A2(n7844), .ZN(n7846) );
  AND2_X1 U9489 ( .A1(n7847), .A2(n7846), .ZN(n7915) );
  INV_X1 U9490 ( .A(n7912), .ZN(n7849) );
  INV_X1 U9491 ( .A(n9431), .ZN(n7848) );
  NAND3_X1 U9492 ( .A1(n7849), .A2(n7872), .A3(n7848), .ZN(n7850) );
  NAND3_X1 U9493 ( .A1(n7915), .A2(n7910), .A3(n7850), .ZN(n7853) );
  NAND2_X1 U9494 ( .A1(n7852), .A2(n7851), .ZN(n7913) );
  AOI21_X1 U9495 ( .B1(n7853), .B2(n7916), .A(n7913), .ZN(n7856) );
  NAND2_X1 U9496 ( .A1(n7855), .A2(n7854), .ZN(n7918) );
  OAI22_X1 U9497 ( .A1(n7856), .A2(n7918), .B1(n7956), .B2(n9125), .ZN(n7860)
         );
  NAND2_X1 U9498 ( .A1(n7945), .A2(n7857), .ZN(n7859) );
  NAND2_X1 U9499 ( .A1(n7859), .A2(n7858), .ZN(n7923) );
  NOR3_X1 U9500 ( .A1(n7867), .A2(n7860), .A3(n7923), .ZN(n7863) );
  NOR4_X1 U9501 ( .A1(n7863), .A2(n7921), .A3(n7862), .A4(n7861), .ZN(n7864)
         );
  AOI21_X1 U9502 ( .B1(n7869), .B2(n7925), .A(n7864), .ZN(n7865) );
  NOR2_X1 U9503 ( .A1(n7867), .A2(n7866), .ZN(n7868) );
  INV_X1 U9504 ( .A(n7872), .ZN(n7909) );
  INV_X1 U9505 ( .A(n7873), .ZN(n7907) );
  INV_X1 U9506 ( .A(n7874), .ZN(n7903) );
  INV_X1 U9507 ( .A(n7875), .ZN(n7897) );
  INV_X1 U9508 ( .A(n7876), .ZN(n7880) );
  NAND2_X1 U9509 ( .A1(n9143), .A2(n7877), .ZN(n7879) );
  NAND2_X1 U9510 ( .A1(n6487), .A2(n6328), .ZN(n7878) );
  AND4_X1 U9511 ( .A1(n7880), .A2(n7879), .A3(n7878), .A4(n4976), .ZN(n7884)
         );
  AND4_X1 U9512 ( .A1(n7884), .A2(n7883), .A3(n7882), .A4(n7881), .ZN(n7887)
         );
  OAI211_X1 U9513 ( .C1(n7888), .C2(n7887), .A(n7886), .B(n7885), .ZN(n7892)
         );
  INV_X1 U9514 ( .A(n7889), .ZN(n7890) );
  AOI21_X1 U9515 ( .B1(n7892), .B2(n7891), .A(n7890), .ZN(n7896) );
  NAND2_X1 U9516 ( .A1(n7894), .A2(n7893), .ZN(n7895) );
  OR3_X1 U9517 ( .A1(n7897), .A2(n7896), .A3(n7895), .ZN(n7899) );
  AOI21_X1 U9518 ( .B1(n7900), .B2(n7899), .A(n7898), .ZN(n7902) );
  OAI21_X1 U9519 ( .B1(n7903), .B2(n7902), .A(n7901), .ZN(n7906) );
  INV_X1 U9520 ( .A(n7904), .ZN(n7905) );
  AOI21_X1 U9521 ( .B1(n7907), .B2(n7906), .A(n7905), .ZN(n7908) );
  OR2_X1 U9522 ( .A1(n7909), .A2(n7908), .ZN(n7911) );
  OAI21_X1 U9523 ( .B1(n7912), .B2(n7911), .A(n7910), .ZN(n7914) );
  AOI21_X1 U9524 ( .B1(n7916), .B2(n7914), .A(n7913), .ZN(n7920) );
  INV_X1 U9525 ( .A(n7915), .ZN(n7917) );
  NAND2_X1 U9526 ( .A1(n7917), .A2(n7916), .ZN(n7919) );
  AOI21_X1 U9527 ( .B1(n7920), .B2(n7919), .A(n7918), .ZN(n7924) );
  OAI211_X1 U9528 ( .C1(n7924), .C2(n7923), .A(n4464), .B(n7922), .ZN(n7926)
         );
  NAND2_X1 U9529 ( .A1(n7926), .A2(n7925), .ZN(n7930) );
  NAND2_X1 U9530 ( .A1(n7930), .A2(n9269), .ZN(n7927) );
  OR3_X1 U9531 ( .A1(n7936), .A2(n7935), .A3(n9158), .ZN(n7939) );
  INV_X1 U9532 ( .A(n7937), .ZN(n7938) );
  NAND3_X1 U9533 ( .A1(n7939), .A2(P1_B_REG_SCAN_IN), .A3(n7938), .ZN(n7940)
         );
  OAI211_X1 U9534 ( .C1(n7943), .C2(n7942), .A(n7941), .B(n7940), .ZN(P1_U3242) );
  INV_X1 U9535 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n7947) );
  AOI211_X1 U9536 ( .C1(n7945), .C2(n7944), .A(n9510), .B(n9275), .ZN(n7952)
         );
  NOR2_X1 U9537 ( .A1(n7952), .A2(n9530), .ZN(n7949) );
  MUX2_X1 U9538 ( .A(n7947), .B(n7949), .S(n9871), .Z(n7948) );
  OAI21_X1 U9539 ( .B1(n7956), .B2(n9676), .A(n7948), .ZN(P1_U3520) );
  INV_X1 U9540 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7950) );
  MUX2_X1 U9541 ( .A(n7950), .B(n7949), .S(n9876), .Z(n7951) );
  OAI21_X1 U9542 ( .B1(n7956), .B2(n9633), .A(n7951), .ZN(P1_U3552) );
  NAND2_X1 U9543 ( .A1(n7952), .A2(n9527), .ZN(n7955) );
  INV_X1 U9544 ( .A(n9530), .ZN(n7953) );
  NOR2_X1 U9545 ( .A1(n9826), .A2(n7953), .ZN(n9277) );
  AOI21_X1 U9546 ( .B1(n9826), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9277), .ZN(
        n7954) );
  OAI211_X1 U9547 ( .C1(n7956), .C2(n9514), .A(n7955), .B(n7954), .ZN(P1_U3264) );
  INV_X1 U9548 ( .A(n8216), .ZN(n7971) );
  OAI222_X1 U9549 ( .A1(n7957), .A2(n8217), .B1(n8960), .B2(n7971), .C1(
        P2_U3151), .C2(n5787), .ZN(P2_U3265) );
  INV_X1 U9550 ( .A(n7959), .ZN(n8963) );
  OAI222_X1 U9551 ( .A1(n9694), .A2(n7960), .B1(P1_U3086), .B2(n7958), .C1(
        n9688), .C2(n8963), .ZN(P1_U3326) );
  XNOR2_X1 U9552 ( .A(n7962), .B(n7961), .ZN(n7963) );
  NAND2_X1 U9553 ( .A1(n7963), .A2(n9115), .ZN(n7967) );
  AOI22_X1 U9554 ( .A1(n9060), .A2(n7965), .B1(n7964), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7966) );
  OAI211_X1 U9555 ( .C1(n6328), .C2(n9124), .A(n7967), .B(n7966), .ZN(P1_U3222) );
  INV_X1 U9556 ( .A(n8965), .ZN(n7968) );
  OAI222_X1 U9557 ( .A1(n9694), .A2(n7969), .B1(n9688), .B2(n7968), .C1(n4352), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U9558 ( .A1(n7972), .A2(n9694), .B1(n9688), .B2(n7971), .C1(
        P1_U3086), .C2(n4948), .ZN(P1_U3325) );
  OR2_X1 U9559 ( .A1(n7973), .A2(n8167), .ZN(n7974) );
  XNOR2_X1 U9560 ( .A(n8825), .B(n7207), .ZN(n8136) );
  INV_X1 U9561 ( .A(n8136), .ZN(n7976) );
  NAND2_X1 U9562 ( .A1(n7976), .A2(n9709), .ZN(n7977) );
  NAND2_X1 U9563 ( .A1(n8138), .A2(n7977), .ZN(n7979) );
  NAND2_X1 U9564 ( .A1(n8136), .A2(n8456), .ZN(n7978) );
  NAND2_X1 U9565 ( .A1(n7979), .A2(n7978), .ZN(n8048) );
  INV_X1 U9566 ( .A(n8048), .ZN(n7981) );
  XNOR2_X1 U9567 ( .A(n9726), .B(n8029), .ZN(n7982) );
  XOR2_X1 U9568 ( .A(n8820), .B(n7982), .Z(n8049) );
  NAND2_X1 U9569 ( .A1(n7982), .A2(n8339), .ZN(n7983) );
  XNOR2_X1 U9570 ( .A(n9719), .B(n8029), .ZN(n7984) );
  XOR2_X1 U9571 ( .A(n8455), .B(n7984), .Z(n8200) );
  INV_X1 U9572 ( .A(n7984), .ZN(n7985) );
  NAND2_X1 U9573 ( .A1(n7985), .A2(n8455), .ZN(n7986) );
  NAND2_X1 U9574 ( .A1(n8202), .A2(n7986), .ZN(n8097) );
  XNOR2_X1 U9575 ( .A(n8878), .B(n8029), .ZN(n7987) );
  XNOR2_X1 U9576 ( .A(n7987), .B(n8799), .ZN(n8096) );
  INV_X1 U9577 ( .A(n7987), .ZN(n7988) );
  AOI22_X1 U9578 ( .A1(n8097), .A2(n8096), .B1(n7988), .B2(n8799), .ZN(n8104)
         );
  XNOR2_X1 U9579 ( .A(n8945), .B(n7207), .ZN(n7989) );
  NOR2_X1 U9580 ( .A1(n7989), .A2(n8768), .ZN(n8177) );
  AOI21_X1 U9581 ( .B1(n7989), .B2(n8768), .A(n8177), .ZN(n8105) );
  NAND2_X1 U9582 ( .A1(n8104), .A2(n8105), .ZN(n8175) );
  INV_X1 U9583 ( .A(n8177), .ZN(n7990) );
  NAND2_X1 U9584 ( .A1(n8175), .A2(n7990), .ZN(n8061) );
  XNOR2_X1 U9585 ( .A(n8938), .B(n8029), .ZN(n7992) );
  NAND2_X1 U9586 ( .A1(n7992), .A2(n7991), .ZN(n8063) );
  INV_X1 U9587 ( .A(n7992), .ZN(n7993) );
  NAND2_X1 U9588 ( .A1(n7993), .A2(n8779), .ZN(n7994) );
  XNOR2_X1 U9589 ( .A(n8932), .B(n8029), .ZN(n7995) );
  NAND2_X1 U9590 ( .A1(n7995), .A2(n8182), .ZN(n8124) );
  INV_X1 U9591 ( .A(n7995), .ZN(n7996) );
  NAND2_X1 U9592 ( .A1(n7996), .A2(n8769), .ZN(n7997) );
  XNOR2_X1 U9593 ( .A(n8926), .B(n8029), .ZN(n7998) );
  NAND2_X1 U9594 ( .A1(n7998), .A2(n8068), .ZN(n8076) );
  INV_X1 U9595 ( .A(n7998), .ZN(n7999) );
  NAND2_X1 U9596 ( .A1(n7999), .A2(n8754), .ZN(n8000) );
  XNOR2_X1 U9597 ( .A(n8920), .B(n8029), .ZN(n8009) );
  XNOR2_X1 U9598 ( .A(n8009), .B(n8744), .ZN(n8077) );
  AND2_X1 U9599 ( .A1(n8125), .A2(n8077), .ZN(n8004) );
  AND2_X1 U9600 ( .A1(n8065), .A2(n8004), .ZN(n8002) );
  AND2_X1 U9601 ( .A1(n8176), .A2(n8002), .ZN(n8001) );
  INV_X1 U9602 ( .A(n8002), .ZN(n8003) );
  OR2_X1 U9603 ( .A1(n8003), .A2(n8063), .ZN(n8007) );
  INV_X1 U9604 ( .A(n8004), .ZN(n8005) );
  OR2_X1 U9605 ( .A1(n8005), .A2(n8124), .ZN(n8006) );
  AND2_X1 U9606 ( .A1(n8007), .A2(n8006), .ZN(n8008) );
  XNOR2_X1 U9607 ( .A(n8914), .B(n7207), .ZN(n8012) );
  OR2_X1 U9608 ( .A1(n8012), .A2(n8734), .ZN(n8149) );
  NAND2_X1 U9609 ( .A1(n8009), .A2(n8130), .ZN(n8011) );
  INV_X1 U9610 ( .A(n8077), .ZN(n8010) );
  OR2_X1 U9611 ( .A1(n8010), .A2(n8076), .ZN(n8079) );
  AND2_X1 U9612 ( .A1(n8011), .A2(n8079), .ZN(n8147) );
  NAND2_X1 U9613 ( .A1(n8012), .A2(n8734), .ZN(n8148) );
  XNOR2_X1 U9614 ( .A(n8712), .B(n8029), .ZN(n8015) );
  INV_X1 U9615 ( .A(n8014), .ZN(n8016) );
  NAND2_X1 U9616 ( .A1(n8016), .A2(n8015), .ZN(n8113) );
  XNOR2_X1 U9617 ( .A(n8902), .B(n8029), .ZN(n8019) );
  NAND2_X1 U9618 ( .A1(n8019), .A2(n8707), .ZN(n8018) );
  AND2_X1 U9619 ( .A1(n8113), .A2(n8018), .ZN(n8017) );
  NAND2_X1 U9620 ( .A1(n8114), .A2(n8017), .ZN(n8087) );
  INV_X1 U9621 ( .A(n8018), .ZN(n8020) );
  XNOR2_X1 U9622 ( .A(n8019), .B(n8680), .ZN(n8116) );
  OR2_X1 U9623 ( .A1(n8020), .A2(n8116), .ZN(n8086) );
  XNOR2_X1 U9624 ( .A(n8895), .B(n8029), .ZN(n8022) );
  XNOR2_X1 U9625 ( .A(n8022), .B(n8454), .ZN(n8089) );
  AND2_X1 U9626 ( .A1(n8086), .A2(n8089), .ZN(n8021) );
  NAND2_X1 U9627 ( .A1(n8087), .A2(n8021), .ZN(n8024) );
  NAND2_X1 U9628 ( .A1(n8022), .A2(n8693), .ZN(n8023) );
  NAND2_X2 U9629 ( .A1(n8024), .A2(n8023), .ZN(n8192) );
  XNOR2_X1 U9630 ( .A(n8671), .B(n7207), .ZN(n8025) );
  NAND2_X1 U9631 ( .A1(n8025), .A2(n8681), .ZN(n8189) );
  INV_X1 U9632 ( .A(n8025), .ZN(n8026) );
  NAND2_X1 U9633 ( .A1(n8026), .A2(n8090), .ZN(n8190) );
  XNOR2_X1 U9634 ( .A(n8661), .B(n8029), .ZN(n8027) );
  XOR2_X1 U9635 ( .A(n8453), .B(n8027), .Z(n8038) );
  XOR2_X1 U9636 ( .A(n8029), .B(n8239), .Z(n8030) );
  AOI22_X1 U9637 ( .A1(n8205), .A2(n8453), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8033) );
  NAND2_X1 U9638 ( .A1(n8210), .A2(n8031), .ZN(n8032) );
  OAI211_X1 U9639 ( .C1(n8034), .C2(n8207), .A(n8033), .B(n8032), .ZN(n8035)
         );
  AOI21_X1 U9640 ( .B1(n8267), .B2(n8196), .A(n8035), .ZN(n8036) );
  OAI21_X1 U9641 ( .B1(n8037), .B2(n8199), .A(n8036), .ZN(P2_U3160) );
  XNOR2_X1 U9642 ( .A(n8039), .B(n8038), .ZN(n8045) );
  AOI22_X1 U9643 ( .A1(n8205), .A2(n8681), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8041) );
  NAND2_X1 U9644 ( .A1(n8210), .A2(n8660), .ZN(n8040) );
  OAI211_X1 U9645 ( .C1(n8042), .C2(n8207), .A(n8041), .B(n8040), .ZN(n8043)
         );
  AOI21_X1 U9646 ( .B1(n8661), .B2(n8196), .A(n8043), .ZN(n8044) );
  OAI21_X1 U9647 ( .B1(n8045), .B2(n8199), .A(n8044), .ZN(P2_U3154) );
  INV_X1 U9648 ( .A(n8046), .ZN(n8047) );
  AOI21_X1 U9649 ( .B1(n8049), .B2(n8048), .A(n8047), .ZN(n8054) );
  INV_X1 U9650 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10016) );
  NOR2_X1 U9651 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10016), .ZN(n8514) );
  NOR2_X1 U9652 ( .A1(n8207), .A2(n9711), .ZN(n8050) );
  AOI211_X1 U9653 ( .C1(n8205), .C2(n8456), .A(n8514), .B(n8050), .ZN(n8051)
         );
  OAI21_X1 U9654 ( .B1(n9698), .B2(n8183), .A(n8051), .ZN(n8052) );
  AOI21_X1 U9655 ( .B1(n9726), .B2(n8196), .A(n8052), .ZN(n8053) );
  OAI21_X1 U9656 ( .B1(n8054), .B2(n8199), .A(n8053), .ZN(P2_U3155) );
  XNOR2_X1 U9657 ( .A(n8055), .B(n8720), .ZN(n8060) );
  AOI22_X1 U9658 ( .A1(n8205), .A2(n8734), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8057) );
  NAND2_X1 U9659 ( .A1(n8210), .A2(n8711), .ZN(n8056) );
  OAI211_X1 U9660 ( .C1(n8707), .C2(n8207), .A(n8057), .B(n8056), .ZN(n8058)
         );
  AOI21_X1 U9661 ( .B1(n8712), .B2(n8196), .A(n8058), .ZN(n8059) );
  OAI21_X1 U9662 ( .B1(n8060), .B2(n8199), .A(n8059), .ZN(P2_U3156) );
  NAND2_X1 U9663 ( .A1(n8061), .A2(n8176), .ZN(n8064) );
  INV_X1 U9664 ( .A(n8064), .ZN(n8180) );
  INV_X1 U9665 ( .A(n8063), .ZN(n8062) );
  NOR3_X1 U9666 ( .A1(n8180), .A2(n8062), .A3(n8065), .ZN(n8067) );
  NAND2_X1 U9667 ( .A1(n8064), .A2(n8063), .ZN(n8066) );
  NAND2_X1 U9668 ( .A1(n8066), .A2(n8065), .ZN(n8074) );
  INV_X1 U9669 ( .A(n8074), .ZN(n8127) );
  OAI21_X1 U9670 ( .B1(n8067), .B2(n8127), .A(n8179), .ZN(n8072) );
  NAND2_X1 U9671 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8636) );
  OAI21_X1 U9672 ( .B1(n8207), .B2(n8068), .A(n8636), .ZN(n8070) );
  NOR2_X1 U9673 ( .A1(n8183), .A2(n8757), .ZN(n8069) );
  AOI211_X1 U9674 ( .C1(n8205), .C2(n8779), .A(n8070), .B(n8069), .ZN(n8071)
         );
  OAI211_X1 U9675 ( .C1(n8073), .C2(n8213), .A(n8072), .B(n8071), .ZN(P2_U3159) );
  INV_X1 U9676 ( .A(n8920), .ZN(n8085) );
  NAND2_X1 U9677 ( .A1(n8074), .A2(n8124), .ZN(n8075) );
  INV_X1 U9678 ( .A(n8076), .ZN(n8078) );
  NOR3_X1 U9679 ( .A1(n8128), .A2(n8078), .A3(n8077), .ZN(n8080) );
  OAI21_X1 U9680 ( .B1(n8080), .B2(n4399), .A(n8179), .ZN(n8084) );
  AOI22_X1 U9681 ( .A1(n8205), .A2(n8754), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8081) );
  OAI21_X1 U9682 ( .B1(n8708), .B2(n8207), .A(n8081), .ZN(n8082) );
  AOI21_X1 U9683 ( .B1(n8737), .B2(n8210), .A(n8082), .ZN(n8083) );
  OAI211_X1 U9684 ( .C1(n8085), .C2(n8213), .A(n8084), .B(n8083), .ZN(P2_U3163) );
  AND2_X1 U9685 ( .A1(n8087), .A2(n8086), .ZN(n8088) );
  XOR2_X1 U9686 ( .A(n8089), .B(n8088), .Z(n8095) );
  OAI22_X1 U9687 ( .A1(n8207), .A2(n8090), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10076), .ZN(n8092) );
  NOR2_X1 U9688 ( .A1(n8120), .A2(n8707), .ZN(n8091) );
  AOI211_X1 U9689 ( .C1(n8685), .C2(n8210), .A(n8092), .B(n8091), .ZN(n8094)
         );
  NAND2_X1 U9690 ( .A1(n8895), .A2(n8196), .ZN(n8093) );
  OAI211_X1 U9691 ( .C1(n8095), .C2(n8199), .A(n8094), .B(n8093), .ZN(P2_U3165) );
  XNOR2_X1 U9692 ( .A(n8097), .B(n8096), .ZN(n8103) );
  INV_X1 U9693 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8098) );
  NOR2_X1 U9694 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8098), .ZN(n8558) );
  NOR2_X1 U9695 ( .A1(n8207), .A2(n8788), .ZN(n8099) );
  AOI211_X1 U9696 ( .C1(n8205), .C2(n8455), .A(n8558), .B(n8099), .ZN(n8100)
         );
  OAI21_X1 U9697 ( .B1(n8789), .B2(n8183), .A(n8100), .ZN(n8101) );
  AOI21_X1 U9698 ( .B1(n8878), .B2(n8196), .A(n8101), .ZN(n8102) );
  OAI21_X1 U9699 ( .B1(n8103), .B2(n8199), .A(n8102), .ZN(P2_U3166) );
  INV_X1 U9700 ( .A(n8945), .ZN(n8112) );
  OAI21_X1 U9701 ( .B1(n8105), .B2(n8104), .A(n8175), .ZN(n8106) );
  NAND2_X1 U9702 ( .A1(n8106), .A2(n8179), .ZN(n8111) );
  INV_X1 U9703 ( .A(n8107), .ZN(n8781) );
  NOR2_X1 U9704 ( .A1(n10062), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8589) );
  AOI21_X1 U9705 ( .B1(n8117), .B2(n8779), .A(n8589), .ZN(n8108) );
  OAI21_X1 U9706 ( .B1(n8208), .B2(n8120), .A(n8108), .ZN(n8109) );
  AOI21_X1 U9707 ( .B1(n8781), .B2(n8210), .A(n8109), .ZN(n8110) );
  OAI211_X1 U9708 ( .C1(n8112), .C2(n8213), .A(n8111), .B(n8110), .ZN(P2_U3168) );
  NAND2_X1 U9709 ( .A1(n8114), .A2(n8113), .ZN(n8115) );
  XOR2_X1 U9710 ( .A(n8116), .B(n8115), .Z(n8123) );
  AOI22_X1 U9711 ( .A1(n8117), .A2(n8454), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8119) );
  NAND2_X1 U9712 ( .A1(n8210), .A2(n8696), .ZN(n8118) );
  OAI211_X1 U9713 ( .C1(n8694), .C2(n8120), .A(n8119), .B(n8118), .ZN(n8121)
         );
  AOI21_X1 U9714 ( .B1(n8902), .B2(n8196), .A(n8121), .ZN(n8122) );
  OAI21_X1 U9715 ( .B1(n8123), .B2(n8199), .A(n8122), .ZN(P2_U3169) );
  INV_X1 U9716 ( .A(n8124), .ZN(n8126) );
  NOR3_X1 U9717 ( .A1(n8127), .A2(n8126), .A3(n8125), .ZN(n8129) );
  OAI21_X1 U9718 ( .B1(n8129), .B2(n8128), .A(n8179), .ZN(n8134) );
  OAI22_X1 U9719 ( .A1(n8207), .A2(n8130), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10038), .ZN(n8132) );
  NOR2_X1 U9720 ( .A1(n8183), .A2(n8747), .ZN(n8131) );
  AOI211_X1 U9721 ( .C1(n8205), .C2(n8769), .A(n8132), .B(n8131), .ZN(n8133)
         );
  OAI211_X1 U9722 ( .C1(n8135), .C2(n8213), .A(n8134), .B(n8133), .ZN(P2_U3173) );
  XNOR2_X1 U9723 ( .A(n8136), .B(n8456), .ZN(n8137) );
  XNOR2_X1 U9724 ( .A(n8138), .B(n8137), .ZN(n8145) );
  INV_X1 U9725 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10125) );
  NOR2_X1 U9726 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10125), .ZN(n8485) );
  AOI21_X1 U9727 ( .B1(n8205), .B2(n8821), .A(n8485), .ZN(n8143) );
  NAND2_X1 U9728 ( .A1(n8196), .A2(n8825), .ZN(n8142) );
  INV_X1 U9729 ( .A(n8826), .ZN(n8139) );
  NAND2_X1 U9730 ( .A1(n8210), .A2(n8139), .ZN(n8141) );
  OR2_X1 U9731 ( .A1(n8207), .A2(n8339), .ZN(n8140) );
  NAND4_X1 U9732 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(n8144)
         );
  AOI21_X1 U9733 ( .B1(n8145), .B2(n8179), .A(n8144), .ZN(n8146) );
  INV_X1 U9734 ( .A(n8146), .ZN(P2_U3174) );
  NAND2_X1 U9735 ( .A1(n4370), .A2(n8147), .ZN(n8151) );
  NAND2_X1 U9736 ( .A1(n8149), .A2(n8148), .ZN(n8150) );
  XNOR2_X1 U9737 ( .A(n8151), .B(n8150), .ZN(n8156) );
  AOI22_X1 U9738 ( .A1(n8205), .A2(n8744), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8153) );
  NAND2_X1 U9739 ( .A1(n8210), .A2(n8723), .ZN(n8152) );
  OAI211_X1 U9740 ( .C1(n8694), .C2(n8207), .A(n8153), .B(n8152), .ZN(n8154)
         );
  AOI21_X1 U9741 ( .B1(n8914), .B2(n8196), .A(n8154), .ZN(n8155) );
  OAI21_X1 U9742 ( .B1(n8156), .B2(n8199), .A(n8155), .ZN(P2_U3175) );
  OAI22_X1 U9743 ( .A1(n8159), .A2(n8158), .B1(n8157), .B2(n8458), .ZN(n8162)
         );
  XNOR2_X1 U9744 ( .A(n8160), .B(n8457), .ZN(n8161) );
  XNOR2_X1 U9745 ( .A(n8162), .B(n8161), .ZN(n8173) );
  AOI21_X1 U9746 ( .B1(n8205), .B2(n8458), .A(n8163), .ZN(n8171) );
  NAND2_X1 U9747 ( .A1(n8196), .A2(n8164), .ZN(n8170) );
  INV_X1 U9748 ( .A(n8165), .ZN(n8166) );
  NAND2_X1 U9749 ( .A1(n8210), .A2(n8166), .ZN(n8169) );
  OR2_X1 U9750 ( .A1(n8207), .A2(n8167), .ZN(n8168) );
  NAND4_X1 U9751 ( .A1(n8171), .A2(n8170), .A3(n8169), .A4(n8168), .ZN(n8172)
         );
  AOI21_X1 U9752 ( .B1(n8173), .B2(n8179), .A(n8172), .ZN(n8174) );
  INV_X1 U9753 ( .A(n8174), .ZN(P2_U3176) );
  INV_X1 U9754 ( .A(n8175), .ZN(n8178) );
  NOR3_X1 U9755 ( .A1(n8178), .A2(n8177), .A3(n8176), .ZN(n8181) );
  OAI21_X1 U9756 ( .B1(n8181), .B2(n8180), .A(n8179), .ZN(n8187) );
  NAND2_X1 U9757 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8615) );
  OAI21_X1 U9758 ( .B1(n8207), .B2(n8182), .A(n8615), .ZN(n8185) );
  NOR2_X1 U9759 ( .A1(n8183), .A2(n8772), .ZN(n8184) );
  AOI211_X1 U9760 ( .C1(n8205), .C2(n8768), .A(n8185), .B(n8184), .ZN(n8186)
         );
  OAI211_X1 U9761 ( .C1(n8188), .C2(n8213), .A(n8187), .B(n8186), .ZN(P2_U3178) );
  NAND2_X1 U9762 ( .A1(n8190), .A2(n8189), .ZN(n8191) );
  XNOR2_X1 U9763 ( .A(n8192), .B(n8191), .ZN(n8198) );
  AOI22_X1 U9764 ( .A1(n8205), .A2(n8454), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8194) );
  NAND2_X1 U9765 ( .A1(n8210), .A2(n8672), .ZN(n8193) );
  OAI211_X1 U9766 ( .C1(n8668), .C2(n8207), .A(n8194), .B(n8193), .ZN(n8195)
         );
  AOI21_X1 U9767 ( .B1(n8671), .B2(n8196), .A(n8195), .ZN(n8197) );
  OAI21_X1 U9768 ( .B1(n8198), .B2(n8199), .A(n8197), .ZN(P2_U3180) );
  INV_X1 U9769 ( .A(n9719), .ZN(n8808) );
  AOI21_X1 U9770 ( .B1(n8201), .B2(n8200), .A(n8199), .ZN(n8203) );
  NAND2_X1 U9771 ( .A1(n8203), .A2(n8202), .ZN(n8212) );
  INV_X1 U9772 ( .A(n8204), .ZN(n8804) );
  NOR2_X1 U9773 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5773), .ZN(n8533) );
  AOI21_X1 U9774 ( .B1(n8205), .B2(n8820), .A(n8533), .ZN(n8206) );
  OAI21_X1 U9775 ( .B1(n8208), .B2(n8207), .A(n8206), .ZN(n8209) );
  AOI21_X1 U9776 ( .B1(n8804), .B2(n8210), .A(n8209), .ZN(n8211) );
  OAI211_X1 U9777 ( .C1(n8808), .C2(n8213), .A(n8212), .B(n8211), .ZN(P2_U3181) );
  INV_X1 U9778 ( .A(n8214), .ZN(n8419) );
  NAND2_X1 U9779 ( .A1(n8216), .A2(n8224), .ZN(n8219) );
  OR2_X1 U9780 ( .A1(n8222), .A2(n8217), .ZN(n8218) );
  NAND2_X1 U9781 ( .A1(n8219), .A2(n8218), .ZN(n8227) );
  NAND2_X1 U9782 ( .A1(n8227), .A2(n8228), .ZN(n8422) );
  NAND2_X1 U9783 ( .A1(n8422), .A2(n8220), .ZN(n8434) );
  INV_X1 U9784 ( .A(n8434), .ZN(n8226) );
  INV_X1 U9785 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8221) );
  NOR2_X1 U9786 ( .A1(n8222), .A2(n8221), .ZN(n8223) );
  NAND2_X1 U9787 ( .A1(n8226), .A2(n8225), .ZN(n8229) );
  INV_X1 U9788 ( .A(n8227), .ZN(n8888) );
  INV_X1 U9789 ( .A(n8228), .ZN(n8452) );
  NAND2_X1 U9790 ( .A1(n8888), .A2(n8452), .ZN(n8238) );
  OAI21_X1 U9791 ( .B1(n8230), .B2(n8229), .A(n4913), .ZN(n8237) );
  NAND2_X1 U9792 ( .A1(n5838), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8233) );
  NAND2_X1 U9793 ( .A1(n5840), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8232) );
  NAND2_X1 U9794 ( .A1(n5839), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8231) );
  AND3_X1 U9795 ( .A1(n8233), .A2(n8232), .A3(n8231), .ZN(n8234) );
  NAND2_X1 U9796 ( .A1(n8235), .A2(n8234), .ZN(n8647) );
  NAND2_X1 U9797 ( .A1(n8833), .A2(n8647), .ZN(n8437) );
  INV_X1 U9798 ( .A(n8238), .ZN(n8421) );
  INV_X1 U9799 ( .A(n8422), .ZN(n8264) );
  INV_X1 U9800 ( .A(n8240), .ZN(n8407) );
  INV_X1 U9801 ( .A(n8686), .ZN(n8679) );
  NAND2_X1 U9802 ( .A1(n8398), .A2(n8394), .ZN(n8699) );
  INV_X1 U9803 ( .A(n8391), .ZN(n8697) );
  OR2_X1 U9804 ( .A1(n8392), .A2(n8697), .ZN(n8704) );
  INV_X1 U9805 ( .A(n8380), .ZN(n8241) );
  INV_X1 U9806 ( .A(n8242), .ZN(n8243) );
  NOR2_X1 U9807 ( .A1(n8763), .A2(n8243), .ZN(n8374) );
  NAND2_X1 U9808 ( .A1(n7135), .A2(n8269), .ZN(n8247) );
  NOR4_X1 U9809 ( .A1(n8247), .A2(n8246), .A3(n8245), .A4(n8244), .ZN(n8250)
         );
  NAND4_X1 U9810 ( .A1(n8250), .A2(n8249), .A3(n8248), .A4(n8287), .ZN(n8253)
         );
  NOR4_X1 U9811 ( .A1(n8253), .A2(n8252), .A3(n8251), .A4(n5897), .ZN(n8254)
         );
  NAND4_X1 U9812 ( .A1(n8328), .A2(n8256), .A3(n8255), .A4(n8254), .ZN(n8257)
         );
  NOR4_X1 U9813 ( .A1(n8802), .A2(n8257), .A3(n9705), .A4(n8828), .ZN(n8258)
         );
  NAND4_X1 U9814 ( .A1(n8371), .A2(n8374), .A3(n8785), .A4(n8258), .ZN(n8259)
         );
  NOR3_X1 U9815 ( .A1(n8742), .A2(n8753), .A3(n8259), .ZN(n8260) );
  NAND3_X1 U9816 ( .A1(n4654), .A2(n8731), .A3(n8260), .ZN(n8261) );
  NOR4_X1 U9817 ( .A1(n8679), .A2(n8699), .A3(n8704), .A4(n8261), .ZN(n8262)
         );
  NAND4_X1 U9818 ( .A1(n4661), .A2(n8669), .A3(n8262), .A4(n8410), .ZN(n8263)
         );
  NOR4_X1 U9819 ( .A1(n8421), .A2(n8264), .A3(n8418), .A4(n8263), .ZN(n8265)
         );
  MUX2_X1 U9820 ( .A(n4670), .B(n8267), .S(n8412), .Z(n8426) );
  INV_X1 U9821 ( .A(n8274), .ZN(n8268) );
  NAND2_X1 U9822 ( .A1(n8268), .A2(n6175), .ZN(n8272) );
  NAND3_X1 U9823 ( .A1(n8270), .A2(n8269), .A3(n6175), .ZN(n8271) );
  NAND4_X1 U9824 ( .A1(n8272), .A2(n8412), .A3(n8273), .A4(n8271), .ZN(n8277)
         );
  NAND2_X1 U9825 ( .A1(n8274), .A2(n8273), .ZN(n8275) );
  NAND2_X1 U9826 ( .A1(n8275), .A2(n8432), .ZN(n8276) );
  NAND2_X1 U9827 ( .A1(n8277), .A2(n8276), .ZN(n8278) );
  OAI211_X1 U9828 ( .C1(n6175), .C2(n8412), .A(n8278), .B(n7135), .ZN(n8286)
         );
  NAND2_X1 U9829 ( .A1(n8280), .A2(n8279), .ZN(n8283) );
  NAND2_X1 U9830 ( .A1(n8289), .A2(n8281), .ZN(n8282) );
  MUX2_X1 U9831 ( .A(n8283), .B(n8282), .S(n8432), .Z(n8284) );
  INV_X1 U9832 ( .A(n8284), .ZN(n8285) );
  NAND2_X1 U9833 ( .A1(n8286), .A2(n8285), .ZN(n8288) );
  NAND2_X1 U9834 ( .A1(n8288), .A2(n8287), .ZN(n8310) );
  INV_X1 U9835 ( .A(n8289), .ZN(n8292) );
  OAI211_X1 U9836 ( .C1(n8310), .C2(n8292), .A(n8291), .B(n8290), .ZN(n8293)
         );
  NAND3_X1 U9837 ( .A1(n8293), .A2(n8313), .A3(n8307), .ZN(n8295) );
  NAND3_X1 U9838 ( .A1(n8295), .A2(n8314), .A3(n8294), .ZN(n8297) );
  NAND2_X1 U9839 ( .A1(n8297), .A2(n8296), .ZN(n8305) );
  NAND2_X1 U9840 ( .A1(n8317), .A2(n8319), .ZN(n8301) );
  NAND2_X1 U9841 ( .A1(n8299), .A2(n8298), .ZN(n8300) );
  MUX2_X1 U9842 ( .A(n8301), .B(n8300), .S(n8432), .Z(n8302) );
  INV_X1 U9843 ( .A(n8302), .ZN(n8321) );
  INV_X1 U9844 ( .A(n8303), .ZN(n8304) );
  AOI21_X1 U9845 ( .B1(n8305), .B2(n8321), .A(n8304), .ZN(n8324) );
  INV_X1 U9846 ( .A(n8306), .ZN(n9898) );
  NAND2_X1 U9847 ( .A1(n8464), .A2(n9898), .ZN(n8308) );
  OAI211_X1 U9848 ( .C1(n8310), .C2(n8309), .A(n8308), .B(n8307), .ZN(n8312)
         );
  NAND2_X1 U9849 ( .A1(n8312), .A2(n8311), .ZN(n8315) );
  NAND3_X1 U9850 ( .A1(n8315), .A2(n8314), .A3(n8313), .ZN(n8318) );
  NAND3_X1 U9851 ( .A1(n8318), .A2(n8317), .A3(n8316), .ZN(n8322) );
  NAND2_X1 U9852 ( .A1(n8330), .A2(n8319), .ZN(n8320) );
  AOI21_X1 U9853 ( .B1(n8322), .B2(n8321), .A(n8320), .ZN(n8323) );
  MUX2_X1 U9854 ( .A(n8324), .B(n8323), .S(n8432), .Z(n8334) );
  NAND2_X1 U9855 ( .A1(n8332), .A2(n8325), .ZN(n8326) );
  OAI21_X1 U9856 ( .B1(n8334), .B2(n8326), .A(n8331), .ZN(n8327) );
  NAND2_X1 U9857 ( .A1(n8327), .A2(n8432), .ZN(n8329) );
  NAND2_X1 U9858 ( .A1(n8329), .A2(n8328), .ZN(n8362) );
  NAND2_X1 U9859 ( .A1(n8331), .A2(n8330), .ZN(n8333) );
  OAI21_X1 U9860 ( .B1(n8334), .B2(n8333), .A(n8332), .ZN(n8338) );
  NAND3_X1 U9861 ( .A1(n8340), .A2(n8412), .A3(n8335), .ZN(n8336) );
  NOR2_X1 U9862 ( .A1(n8342), .A2(n8336), .ZN(n8337) );
  OAI211_X1 U9863 ( .C1(n8362), .C2(n8338), .A(n8337), .B(n8348), .ZN(n8365)
         );
  OR2_X1 U9864 ( .A1(n9726), .A2(n8339), .ZN(n8359) );
  INV_X1 U9865 ( .A(n8340), .ZN(n8341) );
  NAND3_X1 U9866 ( .A1(n8359), .A2(n8341), .A3(n8432), .ZN(n8355) );
  NAND2_X1 U9867 ( .A1(n8359), .A2(n8432), .ZN(n8344) );
  INV_X1 U9868 ( .A(n8342), .ZN(n8347) );
  NAND3_X1 U9869 ( .A1(n8348), .A2(n8347), .A3(n8412), .ZN(n8343) );
  OAI21_X1 U9870 ( .B1(n8802), .B2(n8344), .A(n8343), .ZN(n8345) );
  NAND2_X1 U9871 ( .A1(n8345), .A2(n9705), .ZN(n8354) );
  NAND4_X1 U9872 ( .A1(n8348), .A2(n8347), .A3(n8346), .A4(n8412), .ZN(n8350)
         );
  OR2_X1 U9873 ( .A1(n8348), .A2(n8412), .ZN(n8349) );
  OAI211_X1 U9874 ( .C1(n8351), .C2(n8432), .A(n8350), .B(n8349), .ZN(n8352)
         );
  INV_X1 U9875 ( .A(n8352), .ZN(n8353) );
  OAI211_X1 U9876 ( .C1(n8802), .C2(n8355), .A(n8354), .B(n8353), .ZN(n8356)
         );
  INV_X1 U9877 ( .A(n8356), .ZN(n8364) );
  NAND4_X1 U9878 ( .A1(n8359), .A2(n8432), .A3(n8358), .A4(n8357), .ZN(n8360)
         );
  NOR2_X1 U9879 ( .A1(n8802), .A2(n8360), .ZN(n8361) );
  NAND2_X1 U9880 ( .A1(n8362), .A2(n8361), .ZN(n8363) );
  NAND4_X1 U9881 ( .A1(n8365), .A2(n8364), .A3(n8785), .A4(n8363), .ZN(n8370)
         );
  MUX2_X1 U9882 ( .A(n8368), .B(n8367), .S(n8412), .Z(n8369) );
  NAND3_X1 U9883 ( .A1(n8370), .A2(n8777), .A3(n8369), .ZN(n8375) );
  INV_X1 U9884 ( .A(n8372), .ZN(n8764) );
  OR2_X1 U9885 ( .A1(n8381), .A2(n8764), .ZN(n8373) );
  INV_X1 U9886 ( .A(n8382), .ZN(n8376) );
  NAND3_X1 U9887 ( .A1(n8376), .A2(n8726), .A3(n8380), .ZN(n8377) );
  NAND3_X1 U9888 ( .A1(n8377), .A2(n8386), .A3(n8383), .ZN(n8379) );
  NAND2_X1 U9889 ( .A1(n8385), .A2(n8384), .ZN(n8387) );
  MUX2_X1 U9890 ( .A(n8389), .B(n8388), .S(n8412), .Z(n8390) );
  NAND2_X1 U9891 ( .A1(n8397), .A2(n8391), .ZN(n8393) );
  NAND3_X1 U9892 ( .A1(n8393), .A2(n8398), .A3(n4648), .ZN(n8395) );
  NAND2_X1 U9893 ( .A1(n8395), .A2(n8394), .ZN(n8402) );
  AOI21_X1 U9894 ( .B1(n8397), .B2(n4648), .A(n8396), .ZN(n8400) );
  INV_X1 U9895 ( .A(n8398), .ZN(n8399) );
  OR2_X1 U9896 ( .A1(n8400), .A2(n8399), .ZN(n8401) );
  MUX2_X1 U9897 ( .A(n8402), .B(n8401), .S(n8432), .Z(n8406) );
  MUX2_X1 U9898 ( .A(n8404), .B(n8403), .S(n8412), .Z(n8405) );
  OAI211_X1 U9899 ( .C1(n8406), .C2(n8679), .A(n8669), .B(n8405), .ZN(n8411)
         );
  MUX2_X1 U9900 ( .A(n8408), .B(n8407), .S(n8412), .Z(n8409) );
  NAND3_X1 U9901 ( .A1(n8411), .A2(n8410), .A3(n8409), .ZN(n8417) );
  AND2_X1 U9902 ( .A1(n8661), .A2(n8668), .ZN(n8414) );
  MUX2_X1 U9903 ( .A(n8414), .B(n8413), .S(n8412), .Z(n8415) );
  INV_X1 U9904 ( .A(n8415), .ZN(n8416) );
  NAND2_X1 U9905 ( .A1(n8437), .A2(n8423), .ZN(n8430) );
  INV_X1 U9906 ( .A(n8425), .ZN(n8429) );
  INV_X1 U9907 ( .A(n8426), .ZN(n8427) );
  NOR2_X1 U9908 ( .A1(n8428), .A2(n8427), .ZN(n8438) );
  NAND2_X1 U9909 ( .A1(n8429), .A2(n8438), .ZN(n8431) );
  OAI22_X1 U9910 ( .A1(n8431), .A2(n8430), .B1(n8833), .B2(n8647), .ZN(n8442)
         );
  NOR3_X1 U9911 ( .A1(n8434), .A2(n8433), .A3(n8432), .ZN(n8435) );
  OAI21_X1 U9912 ( .B1(n8436), .B2(n4670), .A(n8435), .ZN(n8440) );
  INV_X1 U9913 ( .A(n8437), .ZN(n8439) );
  NOR3_X1 U9914 ( .A1(n8440), .A2(n8439), .A3(n8438), .ZN(n8441) );
  NAND3_X1 U9915 ( .A1(n8446), .A2(n8445), .A3(n8444), .ZN(n8447) );
  OAI211_X1 U9916 ( .C1(n8448), .C2(n8450), .A(n8447), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8449) );
  OAI21_X1 U9917 ( .B1(n8451), .B2(n8450), .A(n8449), .ZN(P2_U3296) );
  MUX2_X1 U9918 ( .A(n8647), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8609), .Z(
        P2_U3522) );
  MUX2_X1 U9919 ( .A(n8452), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8609), .Z(
        P2_U3521) );
  MUX2_X1 U9920 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n4670), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9921 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8453), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9922 ( .A(n8681), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8609), .Z(
        P2_U3517) );
  MUX2_X1 U9923 ( .A(n8454), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8609), .Z(
        P2_U3516) );
  MUX2_X1 U9924 ( .A(n8680), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8609), .Z(
        P2_U3515) );
  MUX2_X1 U9925 ( .A(n8720), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8609), .Z(
        P2_U3514) );
  MUX2_X1 U9926 ( .A(n8734), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8609), .Z(
        P2_U3513) );
  MUX2_X1 U9927 ( .A(n8744), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8609), .Z(
        P2_U3512) );
  MUX2_X1 U9928 ( .A(n8754), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8609), .Z(
        P2_U3511) );
  MUX2_X1 U9929 ( .A(n8769), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8609), .Z(
        P2_U3510) );
  MUX2_X1 U9930 ( .A(n8779), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8609), .Z(
        P2_U3509) );
  MUX2_X1 U9931 ( .A(n8768), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8609), .Z(
        P2_U3508) );
  MUX2_X1 U9932 ( .A(n8799), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8609), .Z(
        P2_U3507) );
  MUX2_X1 U9933 ( .A(n8455), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8609), .Z(
        P2_U3506) );
  MUX2_X1 U9934 ( .A(n8820), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8609), .Z(
        P2_U3505) );
  MUX2_X1 U9935 ( .A(n8456), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8609), .Z(
        P2_U3504) );
  MUX2_X1 U9936 ( .A(n8821), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8609), .Z(
        P2_U3503) );
  MUX2_X1 U9937 ( .A(n8457), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8609), .Z(
        P2_U3502) );
  MUX2_X1 U9938 ( .A(n8458), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8609), .Z(
        P2_U3501) );
  MUX2_X1 U9939 ( .A(n8459), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8609), .Z(
        P2_U3500) );
  MUX2_X1 U9940 ( .A(n8460), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8609), .Z(
        P2_U3499) );
  MUX2_X1 U9941 ( .A(n8461), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8609), .Z(
        P2_U3498) );
  MUX2_X1 U9942 ( .A(n8462), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8609), .Z(
        P2_U3497) );
  MUX2_X1 U9943 ( .A(n8463), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8609), .Z(
        P2_U3496) );
  MUX2_X1 U9944 ( .A(n8464), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8609), .Z(
        P2_U3495) );
  MUX2_X1 U9945 ( .A(n8465), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8609), .Z(
        P2_U3494) );
  MUX2_X1 U9946 ( .A(n6843), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8609), .Z(
        P2_U3493) );
  MUX2_X1 U9947 ( .A(n5819), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8609), .Z(
        P2_U3492) );
  MUX2_X1 U9948 ( .A(n8466), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8609), .Z(
        P2_U3491) );
  INV_X1 U9949 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8471) );
  OR2_X1 U9950 ( .A1(n8483), .A2(n8467), .ZN(n8468) );
  AOI21_X1 U9951 ( .B1(n8471), .B2(n8470), .A(n8496), .ZN(n8492) );
  INV_X1 U9952 ( .A(n8472), .ZN(n8478) );
  MUX2_X1 U9953 ( .A(n8471), .B(n8473), .S(n8626), .Z(n8474) );
  NAND2_X1 U9954 ( .A1(n8474), .A2(n8495), .ZN(n8505) );
  INV_X1 U9955 ( .A(n8474), .ZN(n8475) );
  NAND2_X1 U9956 ( .A1(n8475), .A2(n8509), .ZN(n8476) );
  AND2_X1 U9957 ( .A1(n8505), .A2(n8476), .ZN(n8477) );
  OAI21_X1 U9958 ( .B1(n8479), .B2(n8478), .A(n8477), .ZN(n8506) );
  INV_X1 U9959 ( .A(n8506), .ZN(n8481) );
  NOR3_X1 U9960 ( .A1(n8479), .A2(n8478), .A3(n8477), .ZN(n8480) );
  OAI21_X1 U9961 ( .B1(n8481), .B2(n8480), .A(n9883), .ZN(n8491) );
  OAI21_X1 U9962 ( .B1(n8483), .B2(n7441), .A(n8482), .ZN(n8508) );
  XNOR2_X1 U9963 ( .A(n8508), .B(n8495), .ZN(n8484) );
  NAND2_X1 U9964 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n8484), .ZN(n8510) );
  OAI21_X1 U9965 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n8484), .A(n8510), .ZN(
        n8489) );
  INV_X1 U9966 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8487) );
  AOI21_X1 U9967 ( .B1(n8559), .B2(n8495), .A(n8485), .ZN(n8486) );
  OAI21_X1 U9968 ( .B1(n8487), .B2(n8618), .A(n8486), .ZN(n8488) );
  AOI21_X1 U9969 ( .B1(n8489), .B2(n8595), .A(n8488), .ZN(n8490) );
  OAI211_X1 U9970 ( .C1(n8492), .C2(n8642), .A(n8491), .B(n8490), .ZN(P2_U3195) );
  NOR2_X1 U9971 ( .A1(n8495), .A2(n8494), .ZN(n8497) );
  NAND2_X1 U9972 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8529), .ZN(n8523) );
  OAI21_X1 U9973 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8529), .A(n8523), .ZN(
        n8498) );
  AOI21_X1 U9974 ( .B1(n4421), .B2(n8498), .A(n8525), .ZN(n8522) );
  MUX2_X1 U9975 ( .A(n8500), .B(n8499), .S(n8626), .Z(n8501) );
  NAND2_X1 U9976 ( .A1(n8501), .A2(n8515), .ZN(n8536) );
  INV_X1 U9977 ( .A(n8501), .ZN(n8502) );
  NAND2_X1 U9978 ( .A1(n8502), .A2(n8529), .ZN(n8503) );
  NAND2_X1 U9979 ( .A1(n8536), .A2(n8503), .ZN(n8504) );
  AOI21_X1 U9980 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(n8538) );
  AND3_X1 U9981 ( .A1(n8506), .A2(n8505), .A3(n8504), .ZN(n8507) );
  OAI21_X1 U9982 ( .B1(n8538), .B2(n8507), .A(n9883), .ZN(n8521) );
  AOI22_X1 U9983 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8529), .B1(n8515), .B2(
        n8499), .ZN(n8513) );
  NAND2_X1 U9984 ( .A1(n8509), .A2(n8508), .ZN(n8511) );
  OAI21_X1 U9985 ( .B1(n8513), .B2(n8512), .A(n8530), .ZN(n8519) );
  INV_X1 U9986 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8517) );
  AOI21_X1 U9987 ( .B1(n8559), .B2(n8515), .A(n8514), .ZN(n8516) );
  OAI21_X1 U9988 ( .B1(n8517), .B2(n8618), .A(n8516), .ZN(n8518) );
  AOI21_X1 U9989 ( .B1(n8519), .B2(n8595), .A(n8518), .ZN(n8520) );
  OAI211_X1 U9990 ( .C1(n8522), .C2(n8642), .A(n8521), .B(n8520), .ZN(P2_U3196) );
  INV_X1 U9991 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8528) );
  AOI21_X1 U9992 ( .B1(n8528), .B2(n8527), .A(n8549), .ZN(n8546) );
  NAND2_X1 U9993 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8529), .ZN(n8531) );
  NAND2_X1 U9994 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8532), .ZN(n8554) );
  OAI21_X1 U9995 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8532), .A(n8554), .ZN(
        n8544) );
  INV_X1 U9996 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8535) );
  AOI21_X1 U9997 ( .B1(n8559), .B2(n8565), .A(n8533), .ZN(n8534) );
  OAI21_X1 U9998 ( .B1(n8535), .B2(n8618), .A(n8534), .ZN(n8543) );
  INV_X1 U9999 ( .A(n8536), .ZN(n8537) );
  NOR2_X1 U10000 ( .A1(n8538), .A2(n8537), .ZN(n8540) );
  MUX2_X1 U10001 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8626), .Z(n8562) );
  XNOR2_X1 U10002 ( .A(n8562), .B(n8526), .ZN(n8539) );
  NOR2_X1 U10003 ( .A1(n8540), .A2(n8539), .ZN(n8563) );
  AOI21_X1 U10004 ( .B1(n8540), .B2(n8539), .A(n8563), .ZN(n8541) );
  NOR2_X1 U10005 ( .A1(n8541), .A2(n8591), .ZN(n8542) );
  AOI211_X1 U10006 ( .C1(n8595), .C2(n8544), .A(n8543), .B(n8542), .ZN(n8545)
         );
  OAI21_X1 U10007 ( .B1(n8546), .B2(n8642), .A(n8545), .ZN(P2_U3197) );
  NOR2_X1 U10008 ( .A1(n8565), .A2(n8548), .ZN(n8550) );
  NAND2_X1 U10009 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8578), .ZN(n8551) );
  OAI21_X1 U10010 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8578), .A(n8551), .ZN(
        n8552) );
  AOI21_X1 U10011 ( .B1(n4378), .B2(n8552), .A(n8577), .ZN(n8576) );
  AOI22_X1 U10012 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8578), .B1(n8582), .B2(
        n8879), .ZN(n8557) );
  NAND2_X1 U10013 ( .A1(n8526), .A2(n8553), .ZN(n8555) );
  NAND2_X1 U10014 ( .A1(n8555), .A2(n8554), .ZN(n8556) );
  OAI21_X1 U10015 ( .B1(n8557), .B2(n8556), .A(n8581), .ZN(n8574) );
  INV_X1 U10016 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8561) );
  AOI21_X1 U10017 ( .B1(n8559), .B2(n8582), .A(n8558), .ZN(n8560) );
  OAI21_X1 U10018 ( .B1(n8561), .B2(n8618), .A(n8560), .ZN(n8573) );
  INV_X1 U10019 ( .A(n8562), .ZN(n8564) );
  AOI21_X1 U10020 ( .B1(n8565), .B2(n8564), .A(n8563), .ZN(n8568) );
  MUX2_X1 U10021 ( .A(n8790), .B(n8879), .S(n8626), .Z(n8566) );
  NOR2_X1 U10022 ( .A1(n8566), .A2(n8582), .ZN(n8569) );
  NOR2_X1 U10023 ( .A1(n8568), .A2(n8569), .ZN(n8585) );
  AND2_X1 U10024 ( .A1(n8566), .A2(n8582), .ZN(n8584) );
  INV_X1 U10025 ( .A(n8584), .ZN(n8567) );
  NAND2_X1 U10026 ( .A1(n8585), .A2(n8567), .ZN(n8571) );
  OAI21_X1 U10027 ( .B1(n8584), .B2(n8569), .A(n8568), .ZN(n8570) );
  AOI21_X1 U10028 ( .B1(n8571), .B2(n8570), .A(n8591), .ZN(n8572) );
  AOI211_X1 U10029 ( .C1(n8595), .C2(n8574), .A(n8573), .B(n8572), .ZN(n8575)
         );
  OAI21_X1 U10030 ( .B1(n8576), .B2(n8642), .A(n8575), .ZN(P2_U3198) );
  INV_X1 U10031 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8580) );
  AOI21_X1 U10032 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8578), .A(n8577), .ZN(
        n8599) );
  AOI21_X1 U10033 ( .B1(n8580), .B2(n8579), .A(n8600), .ZN(n8597) );
  OAI21_X1 U10034 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8583), .A(n8612), .ZN(
        n8594) );
  NOR2_X1 U10035 ( .A1(n8585), .A2(n8584), .ZN(n8587) );
  MUX2_X1 U10036 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8626), .Z(n8602) );
  XNOR2_X1 U10037 ( .A(n8602), .B(n8611), .ZN(n8586) );
  NOR2_X1 U10038 ( .A1(n8587), .A2(n8586), .ZN(n8603) );
  AOI21_X1 U10039 ( .B1(n8587), .B2(n8586), .A(n8603), .ZN(n8592) );
  NOR2_X1 U10040 ( .A1(n9886), .A2(n8611), .ZN(n8588) );
  AOI211_X1 U10041 ( .C1(n9877), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8589), .B(
        n8588), .ZN(n8590) );
  OAI21_X1 U10042 ( .B1(n8592), .B2(n8591), .A(n8590), .ZN(n8593) );
  AOI21_X1 U10043 ( .B1(n8595), .B2(n8594), .A(n8593), .ZN(n8596) );
  OAI21_X1 U10044 ( .B1(n8597), .B2(n8642), .A(n8596), .ZN(P2_U3199) );
  NOR2_X1 U10045 ( .A1(n8630), .A2(n8771), .ZN(n8598) );
  AOI21_X1 U10046 ( .B1(n8771), .B2(n8630), .A(n8598), .ZN(n8601) );
  AOI21_X1 U10047 ( .B1(n8601), .B2(n4412), .A(n8622), .ZN(n8621) );
  INV_X1 U10048 ( .A(n8602), .ZN(n8604) );
  AOI21_X1 U10049 ( .B1(n8605), .B2(n8604), .A(n8603), .ZN(n8607) );
  MUX2_X1 U10050 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8626), .Z(n8606) );
  NOR2_X1 U10051 ( .A1(n8607), .A2(n8606), .ZN(n8625) );
  INV_X1 U10052 ( .A(n8625), .ZN(n8608) );
  NAND2_X1 U10053 ( .A1(n8607), .A2(n8606), .ZN(n8623) );
  NAND2_X1 U10054 ( .A1(n8608), .A2(n8623), .ZN(n8614) );
  OAI21_X1 U10055 ( .B1(n8614), .B2(n8609), .A(n9886), .ZN(n8620) );
  XNOR2_X1 U10056 ( .A(n8624), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8631) );
  NAND2_X1 U10057 ( .A1(n8611), .A2(n8610), .ZN(n8613) );
  NAND2_X1 U10058 ( .A1(n8613), .A2(n8612), .ZN(n8632) );
  INV_X1 U10059 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8617) );
  NAND3_X1 U10060 ( .A1(n8614), .A2(n9883), .A3(n8630), .ZN(n8616) );
  OAI211_X1 U10061 ( .C1(n8618), .C2(n8617), .A(n8616), .B(n8615), .ZN(n8619)
         );
  XNOR2_X1 U10062 ( .A(n8638), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8627) );
  OAI21_X1 U10063 ( .B1(n8625), .B2(n8624), .A(n8623), .ZN(n8629) );
  XNOR2_X1 U10064 ( .A(n8638), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8633) );
  MUX2_X1 U10065 ( .A(n8627), .B(n8633), .S(n8626), .Z(n8628) );
  XNOR2_X1 U10066 ( .A(n8629), .B(n8628), .ZN(n8640) );
  INV_X1 U10067 ( .A(n8633), .ZN(n8634) );
  NAND2_X1 U10068 ( .A1(n9877), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8637) );
  OAI211_X1 U10069 ( .C1(n9886), .C2(n8638), .A(n8637), .B(n8636), .ZN(n8639)
         );
  OAI21_X1 U10070 ( .B1(n8643), .B2(n8642), .A(n8641), .ZN(P2_U3201) );
  OR2_X1 U10071 ( .A1(n8644), .A2(n9697), .ZN(n8653) );
  INV_X1 U10072 ( .A(n8645), .ZN(n8646) );
  NAND2_X1 U10073 ( .A1(n8647), .A2(n8646), .ZN(n8834) );
  AOI21_X1 U10074 ( .B1(n8653), .B2(n8834), .A(n9718), .ZN(n8649) );
  AOI21_X1 U10075 ( .B1(n9718), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8649), .ZN(
        n8648) );
  OAI21_X1 U10076 ( .B1(n8833), .B2(n8807), .A(n8648), .ZN(P2_U3202) );
  AOI21_X1 U10077 ( .B1(n9718), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8649), .ZN(
        n8650) );
  OAI21_X1 U10078 ( .B1(n8888), .B2(n8807), .A(n8650), .ZN(P2_U3203) );
  INV_X1 U10079 ( .A(n8651), .ZN(n8659) );
  NAND2_X1 U10080 ( .A1(n9718), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8652) );
  OAI211_X1 U10081 ( .C1(n8654), .C2(n8807), .A(n8653), .B(n8652), .ZN(n8655)
         );
  AOI21_X1 U10082 ( .B1(n8657), .B2(n8656), .A(n8655), .ZN(n8658) );
  OAI21_X1 U10083 ( .B1(n8659), .B2(n9718), .A(n8658), .ZN(P2_U3204) );
  AOI21_X1 U10084 ( .B1(n8805), .B2(n8660), .A(n8839), .ZN(n8665) );
  AOI22_X1 U10085 ( .A1(n8661), .A2(n8792), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9718), .ZN(n8664) );
  NAND2_X1 U10086 ( .A1(n8662), .A2(n8830), .ZN(n8663) );
  OAI211_X1 U10087 ( .C1(n8665), .C2(n9718), .A(n8664), .B(n8663), .ZN(
        P2_U3206) );
  XNOR2_X1 U10088 ( .A(n8666), .B(n8669), .ZN(n8667) );
  OAI222_X1 U10089 ( .A1(n9712), .A2(n8668), .B1(n9710), .B2(n8693), .C1(n9708), .C2(n8667), .ZN(n8844) );
  INV_X1 U10090 ( .A(n8844), .ZN(n8676) );
  XNOR2_X1 U10091 ( .A(n8670), .B(n8669), .ZN(n8845) );
  AOI22_X1 U10092 ( .A1(n9718), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8805), .B2(
        n8672), .ZN(n8673) );
  OAI21_X1 U10093 ( .B1(n8892), .B2(n8807), .A(n8673), .ZN(n8674) );
  AOI21_X1 U10094 ( .B1(n8845), .B2(n8830), .A(n8674), .ZN(n8675) );
  OAI21_X1 U10095 ( .B1(n8676), .B2(n9718), .A(n8675), .ZN(P2_U3207) );
  NOR2_X1 U10096 ( .A1(n8677), .A2(n9699), .ZN(n8684) );
  OAI21_X1 U10097 ( .B1(n4384), .B2(n8679), .A(n8678), .ZN(n8682) );
  AOI222_X1 U10098 ( .A1(n8817), .A2(n8682), .B1(n8681), .B2(n8819), .C1(n8680), .C2(n8822), .ZN(n8893) );
  INV_X1 U10099 ( .A(n8893), .ZN(n8683) );
  AOI211_X1 U10100 ( .C1(n8805), .C2(n8685), .A(n8684), .B(n8683), .ZN(n8690)
         );
  XNOR2_X1 U10101 ( .A(n8687), .B(n8686), .ZN(n8898) );
  INV_X1 U10102 ( .A(n8898), .ZN(n8688) );
  AOI22_X1 U10103 ( .A1(n8688), .A2(n8830), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9718), .ZN(n8689) );
  OAI21_X1 U10104 ( .B1(n8690), .B2(n9718), .A(n8689), .ZN(P2_U3208) );
  NOR2_X1 U10105 ( .A1(n8852), .A2(n9699), .ZN(n8695) );
  XOR2_X1 U10106 ( .A(n8699), .B(n8691), .Z(n8692) );
  OAI222_X1 U10107 ( .A1(n9710), .A2(n8694), .B1(n9712), .B2(n8693), .C1(n9708), .C2(n8692), .ZN(n8899) );
  AOI211_X1 U10108 ( .C1(n8805), .C2(n8696), .A(n8695), .B(n8899), .ZN(n8702)
         );
  NOR2_X1 U10109 ( .A1(n8698), .A2(n8697), .ZN(n8700) );
  XNOR2_X1 U10110 ( .A(n8700), .B(n8699), .ZN(n8851) );
  AOI22_X1 U10111 ( .A1(n8851), .A2(n8830), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9718), .ZN(n8701) );
  OAI21_X1 U10112 ( .B1(n8702), .B2(n9718), .A(n8701), .ZN(P2_U3209) );
  XOR2_X1 U10113 ( .A(n8704), .B(n8703), .Z(n8909) );
  INV_X1 U10114 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8710) );
  XOR2_X1 U10115 ( .A(n8705), .B(n8704), .Z(n8706) );
  OAI222_X1 U10116 ( .A1(n9710), .A2(n8708), .B1(n9712), .B2(n8707), .C1(n9708), .C2(n8706), .ZN(n8906) );
  INV_X1 U10117 ( .A(n8906), .ZN(n8709) );
  MUX2_X1 U10118 ( .A(n8710), .B(n8709), .S(n9716), .Z(n8714) );
  AOI22_X1 U10119 ( .A1(n8712), .A2(n8792), .B1(n8805), .B2(n8711), .ZN(n8713)
         );
  OAI211_X1 U10120 ( .C1(n8909), .C2(n8795), .A(n8714), .B(n8713), .ZN(
        P2_U3210) );
  XNOR2_X1 U10121 ( .A(n8715), .B(n8716), .ZN(n8917) );
  INV_X1 U10122 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8722) );
  OR3_X1 U10123 ( .A1(n8729), .A2(n8717), .A3(n8716), .ZN(n8718) );
  NAND2_X1 U10124 ( .A1(n8719), .A2(n8718), .ZN(n8721) );
  AOI222_X1 U10125 ( .A1(n8817), .A2(n8721), .B1(n8720), .B2(n8819), .C1(n8744), .C2(n8822), .ZN(n8912) );
  MUX2_X1 U10126 ( .A(n8722), .B(n8912), .S(n9716), .Z(n8725) );
  AOI22_X1 U10127 ( .A1(n8914), .A2(n8792), .B1(n8805), .B2(n8723), .ZN(n8724)
         );
  OAI211_X1 U10128 ( .C1(n8917), .C2(n8795), .A(n8725), .B(n8724), .ZN(
        P2_U3211) );
  NAND2_X1 U10129 ( .A1(n8727), .A2(n8726), .ZN(n8728) );
  XOR2_X1 U10130 ( .A(n8731), .B(n8728), .Z(n8923) );
  INV_X1 U10131 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8736) );
  INV_X1 U10132 ( .A(n8729), .ZN(n8733) );
  NAND3_X1 U10133 ( .A1(n8741), .A2(n8731), .A3(n8730), .ZN(n8732) );
  NAND2_X1 U10134 ( .A1(n8733), .A2(n8732), .ZN(n8735) );
  AOI222_X1 U10135 ( .A1(n8817), .A2(n8735), .B1(n8734), .B2(n8819), .C1(n8754), .C2(n8822), .ZN(n8918) );
  MUX2_X1 U10136 ( .A(n8736), .B(n8918), .S(n9716), .Z(n8739) );
  AOI22_X1 U10137 ( .A1(n8920), .A2(n8792), .B1(n8805), .B2(n8737), .ZN(n8738)
         );
  OAI211_X1 U10138 ( .C1(n8923), .C2(n8795), .A(n8739), .B(n8738), .ZN(
        P2_U3212) );
  XNOR2_X1 U10139 ( .A(n8740), .B(n8742), .ZN(n8929) );
  INV_X1 U10140 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8746) );
  OAI21_X1 U10141 ( .B1(n8743), .B2(n8742), .A(n8741), .ZN(n8745) );
  AOI222_X1 U10142 ( .A1(n8817), .A2(n8745), .B1(n8769), .B2(n8822), .C1(n8744), .C2(n8819), .ZN(n8924) );
  MUX2_X1 U10143 ( .A(n8746), .B(n8924), .S(n9716), .Z(n8750) );
  INV_X1 U10144 ( .A(n8747), .ZN(n8748) );
  AOI22_X1 U10145 ( .A1(n8926), .A2(n8792), .B1(n8748), .B2(n8805), .ZN(n8749)
         );
  OAI211_X1 U10146 ( .C1(n8929), .C2(n8795), .A(n8750), .B(n8749), .ZN(
        P2_U3213) );
  XOR2_X1 U10147 ( .A(n8751), .B(n8753), .Z(n8935) );
  XNOR2_X1 U10148 ( .A(n8752), .B(n8753), .ZN(n8755) );
  AOI222_X1 U10149 ( .A1(n8817), .A2(n8755), .B1(n8754), .B2(n8819), .C1(n8779), .C2(n8822), .ZN(n8930) );
  MUX2_X1 U10150 ( .A(n8756), .B(n8930), .S(n9716), .Z(n8760) );
  INV_X1 U10151 ( .A(n8757), .ZN(n8758) );
  AOI22_X1 U10152 ( .A1(n8932), .A2(n8792), .B1(n8805), .B2(n8758), .ZN(n8759)
         );
  OAI211_X1 U10153 ( .C1(n8935), .C2(n8795), .A(n8760), .B(n8759), .ZN(
        P2_U3214) );
  NAND2_X1 U10154 ( .A1(n8762), .A2(n8761), .ZN(n8765) );
  NOR2_X1 U10155 ( .A1(n8764), .A2(n8763), .ZN(n8767) );
  XNOR2_X1 U10156 ( .A(n8765), .B(n8767), .ZN(n8941) );
  XOR2_X1 U10157 ( .A(n8767), .B(n8766), .Z(n8770) );
  AOI222_X1 U10158 ( .A1(n8817), .A2(n8770), .B1(n8769), .B2(n8819), .C1(n8768), .C2(n8822), .ZN(n8936) );
  MUX2_X1 U10159 ( .A(n8771), .B(n8936), .S(n9716), .Z(n8775) );
  INV_X1 U10160 ( .A(n8772), .ZN(n8773) );
  AOI22_X1 U10161 ( .A1(n8938), .A2(n8792), .B1(n8805), .B2(n8773), .ZN(n8774)
         );
  OAI211_X1 U10162 ( .C1(n8941), .C2(n8795), .A(n8775), .B(n8774), .ZN(
        P2_U3215) );
  XNOR2_X1 U10163 ( .A(n8776), .B(n8777), .ZN(n8948) );
  XNOR2_X1 U10164 ( .A(n8778), .B(n8777), .ZN(n8780) );
  AOI222_X1 U10165 ( .A1(n8817), .A2(n8780), .B1(n8779), .B2(n8819), .C1(n8799), .C2(n8822), .ZN(n8942) );
  MUX2_X1 U10166 ( .A(n8580), .B(n8942), .S(n9716), .Z(n8783) );
  AOI22_X1 U10167 ( .A1(n8945), .A2(n8792), .B1(n8805), .B2(n8781), .ZN(n8782)
         );
  OAI211_X1 U10168 ( .C1(n8948), .C2(n8795), .A(n8783), .B(n8782), .ZN(
        P2_U3216) );
  XOR2_X1 U10169 ( .A(n8785), .B(n8784), .Z(n8953) );
  XNOR2_X1 U10170 ( .A(n8786), .B(n8785), .ZN(n8787) );
  OAI222_X1 U10171 ( .A1(n9712), .A2(n8788), .B1(n9710), .B2(n9711), .C1(n8787), .C2(n9708), .ZN(n8877) );
  NAND2_X1 U10172 ( .A1(n8877), .A2(n9716), .ZN(n8794) );
  OAI22_X1 U10173 ( .A1(n9716), .A2(n8790), .B1(n8789), .B2(n9697), .ZN(n8791)
         );
  AOI21_X1 U10174 ( .B1(n8878), .B2(n8792), .A(n8791), .ZN(n8793) );
  OAI211_X1 U10175 ( .C1(n8953), .C2(n8795), .A(n8794), .B(n8793), .ZN(
        P2_U3217) );
  INV_X1 U10176 ( .A(n8802), .ZN(n8796) );
  XNOR2_X1 U10177 ( .A(n8797), .B(n8796), .ZN(n8798) );
  NAND2_X1 U10178 ( .A1(n8798), .A2(n8817), .ZN(n8801) );
  AOI22_X1 U10179 ( .A1(n8822), .A2(n8820), .B1(n8799), .B2(n8819), .ZN(n8800)
         );
  XNOR2_X1 U10180 ( .A(n8803), .B(n8802), .ZN(n9720) );
  AOI22_X1 U10181 ( .A1(n9718), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8805), .B2(
        n8804), .ZN(n8806) );
  OAI21_X1 U10182 ( .B1(n8808), .B2(n8807), .A(n8806), .ZN(n8809) );
  AOI21_X1 U10183 ( .B1(n9720), .B2(n8830), .A(n8809), .ZN(n8810) );
  OAI21_X1 U10184 ( .B1(n9722), .B2(n9718), .A(n8810), .ZN(P2_U3218) );
  NAND2_X1 U10185 ( .A1(n8812), .A2(n8811), .ZN(n8814) );
  NAND2_X1 U10186 ( .A1(n8814), .A2(n8813), .ZN(n8816) );
  INV_X1 U10187 ( .A(n8828), .ZN(n8815) );
  XNOR2_X1 U10188 ( .A(n8816), .B(n8815), .ZN(n8818) );
  NAND2_X1 U10189 ( .A1(n8818), .A2(n8817), .ZN(n8824) );
  AOI22_X1 U10190 ( .A1(n8822), .A2(n8821), .B1(n8820), .B2(n8819), .ZN(n8823)
         );
  NAND2_X1 U10191 ( .A1(n8824), .A2(n8823), .ZN(n9731) );
  INV_X1 U10192 ( .A(n8825), .ZN(n9729) );
  OAI22_X1 U10193 ( .A1(n9729), .A2(n9699), .B1(n8826), .B2(n9697), .ZN(n8827)
         );
  OAI21_X1 U10194 ( .B1(n9731), .B2(n8827), .A(n9716), .ZN(n8832) );
  XNOR2_X1 U10195 ( .A(n8829), .B(n8828), .ZN(n9727) );
  AOI22_X1 U10196 ( .A1(n9727), .A2(n8830), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n9718), .ZN(n8831) );
  NAND2_X1 U10197 ( .A1(n8832), .A2(n8831), .ZN(P2_U3220) );
  INV_X1 U10198 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8836) );
  INV_X1 U10199 ( .A(n8833), .ZN(n8882) );
  NAND2_X1 U10200 ( .A1(n8882), .A2(n8874), .ZN(n8835) );
  INV_X1 U10201 ( .A(n8834), .ZN(n8883) );
  NAND2_X1 U10202 ( .A1(n8883), .A2(n9950), .ZN(n8837) );
  OAI211_X1 U10203 ( .C1(n9950), .C2(n8836), .A(n8835), .B(n8837), .ZN(
        P2_U3490) );
  NAND2_X1 U10204 ( .A1(n6277), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8838) );
  OAI211_X1 U10205 ( .C1(n8888), .C2(n8855), .A(n8838), .B(n8837), .ZN(
        P2_U3489) );
  MUX2_X1 U10206 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8839), .S(n9950), .Z(n8843) );
  OAI22_X1 U10207 ( .A1(n8841), .A2(n8881), .B1(n8840), .B2(n8855), .ZN(n8842)
         );
  OR2_X1 U10208 ( .A1(n8843), .A2(n8842), .ZN(P2_U3486) );
  AOI21_X1 U10209 ( .B1(n9933), .B2(n8845), .A(n8844), .ZN(n8889) );
  MUX2_X1 U10210 ( .A(n8846), .B(n8889), .S(n9950), .Z(n8847) );
  OAI21_X1 U10211 ( .B1(n8892), .B2(n8855), .A(n8847), .ZN(P2_U3485) );
  MUX2_X1 U10212 ( .A(n8848), .B(n8893), .S(n9950), .Z(n8850) );
  NAND2_X1 U10213 ( .A1(n8895), .A2(n8874), .ZN(n8849) );
  OAI211_X1 U10214 ( .C1(n8898), .C2(n8881), .A(n8850), .B(n8849), .ZN(
        P2_U3484) );
  MUX2_X1 U10215 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8899), .S(n9950), .Z(n8854) );
  INV_X1 U10216 ( .A(n8851), .ZN(n8905) );
  OAI22_X1 U10217 ( .A1(n8905), .A2(n8881), .B1(n8852), .B2(n8855), .ZN(n8853)
         );
  OR2_X1 U10218 ( .A1(n8854), .A2(n8853), .ZN(P2_U3483) );
  MUX2_X1 U10219 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8906), .S(n9950), .Z(n8857) );
  OAI22_X1 U10220 ( .A1(n8909), .A2(n8881), .B1(n8908), .B2(n8855), .ZN(n8856)
         );
  OR2_X1 U10221 ( .A1(n8857), .A2(n8856), .ZN(P2_U3482) );
  MUX2_X1 U10222 ( .A(n8858), .B(n8912), .S(n9950), .Z(n8860) );
  NAND2_X1 U10223 ( .A1(n8914), .A2(n8874), .ZN(n8859) );
  OAI211_X1 U10224 ( .C1(n8917), .C2(n8881), .A(n8860), .B(n8859), .ZN(
        P2_U3481) );
  INV_X1 U10225 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8861) );
  MUX2_X1 U10226 ( .A(n8861), .B(n8918), .S(n9950), .Z(n8863) );
  NAND2_X1 U10227 ( .A1(n8920), .A2(n8874), .ZN(n8862) );
  OAI211_X1 U10228 ( .C1(n8881), .C2(n8923), .A(n8863), .B(n8862), .ZN(
        P2_U3480) );
  MUX2_X1 U10229 ( .A(n8864), .B(n8924), .S(n9950), .Z(n8866) );
  NAND2_X1 U10230 ( .A1(n8926), .A2(n8874), .ZN(n8865) );
  OAI211_X1 U10231 ( .C1(n8929), .C2(n8881), .A(n8866), .B(n8865), .ZN(
        P2_U3479) );
  MUX2_X1 U10232 ( .A(n8867), .B(n8930), .S(n9950), .Z(n8869) );
  NAND2_X1 U10233 ( .A1(n8932), .A2(n8874), .ZN(n8868) );
  OAI211_X1 U10234 ( .C1(n8881), .C2(n8935), .A(n8869), .B(n8868), .ZN(
        P2_U3478) );
  MUX2_X1 U10235 ( .A(n8870), .B(n8936), .S(n9950), .Z(n8872) );
  NAND2_X1 U10236 ( .A1(n8938), .A2(n8874), .ZN(n8871) );
  OAI211_X1 U10237 ( .C1(n8941), .C2(n8881), .A(n8872), .B(n8871), .ZN(
        P2_U3477) );
  MUX2_X1 U10238 ( .A(n8873), .B(n8942), .S(n9950), .Z(n8876) );
  NAND2_X1 U10239 ( .A1(n8945), .A2(n8874), .ZN(n8875) );
  OAI211_X1 U10240 ( .C1(n8948), .C2(n8881), .A(n8876), .B(n8875), .ZN(
        P2_U3476) );
  AOI21_X1 U10241 ( .B1(n9932), .B2(n8878), .A(n8877), .ZN(n8949) );
  MUX2_X1 U10242 ( .A(n8879), .B(n8949), .S(n9950), .Z(n8880) );
  OAI21_X1 U10243 ( .B1(n8953), .B2(n8881), .A(n8880), .ZN(P2_U3475) );
  INV_X1 U10244 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8885) );
  NAND2_X1 U10245 ( .A1(n8882), .A2(n8944), .ZN(n8884) );
  NAND2_X1 U10246 ( .A1(n9937), .A2(n8883), .ZN(n8886) );
  OAI211_X1 U10247 ( .C1(n8885), .C2(n9937), .A(n8884), .B(n8886), .ZN(
        P2_U3458) );
  NAND2_X1 U10248 ( .A1(n9939), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8887) );
  OAI211_X1 U10249 ( .C1(n8888), .C2(n8907), .A(n8887), .B(n8886), .ZN(
        P2_U3457) );
  INV_X1 U10250 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8890) );
  MUX2_X1 U10251 ( .A(n8890), .B(n8889), .S(n9937), .Z(n8891) );
  OAI21_X1 U10252 ( .B1(n8892), .B2(n8907), .A(n8891), .ZN(P2_U3453) );
  INV_X1 U10253 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8894) );
  MUX2_X1 U10254 ( .A(n8894), .B(n8893), .S(n9937), .Z(n8897) );
  NAND2_X1 U10255 ( .A1(n8895), .A2(n8944), .ZN(n8896) );
  OAI211_X1 U10256 ( .C1(n8898), .C2(n8952), .A(n8897), .B(n8896), .ZN(
        P2_U3452) );
  INV_X1 U10257 ( .A(n8899), .ZN(n8900) );
  MUX2_X1 U10258 ( .A(n8901), .B(n8900), .S(n9937), .Z(n8904) );
  NAND2_X1 U10259 ( .A1(n8902), .A2(n8944), .ZN(n8903) );
  OAI211_X1 U10260 ( .C1(n8905), .C2(n8952), .A(n8904), .B(n8903), .ZN(
        P2_U3451) );
  MUX2_X1 U10261 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8906), .S(n9937), .Z(n8911) );
  OAI22_X1 U10262 ( .A1(n8909), .A2(n8952), .B1(n8908), .B2(n8907), .ZN(n8910)
         );
  OR2_X1 U10263 ( .A1(n8911), .A2(n8910), .ZN(P2_U3450) );
  INV_X1 U10264 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8913) );
  MUX2_X1 U10265 ( .A(n8913), .B(n8912), .S(n9937), .Z(n8916) );
  NAND2_X1 U10266 ( .A1(n8914), .A2(n8944), .ZN(n8915) );
  OAI211_X1 U10267 ( .C1(n8917), .C2(n8952), .A(n8916), .B(n8915), .ZN(
        P2_U3449) );
  INV_X1 U10268 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8919) );
  MUX2_X1 U10269 ( .A(n8919), .B(n8918), .S(n9937), .Z(n8922) );
  NAND2_X1 U10270 ( .A1(n8920), .A2(n8944), .ZN(n8921) );
  OAI211_X1 U10271 ( .C1(n8923), .C2(n8952), .A(n8922), .B(n8921), .ZN(
        P2_U3448) );
  MUX2_X1 U10272 ( .A(n8925), .B(n8924), .S(n9937), .Z(n8928) );
  NAND2_X1 U10273 ( .A1(n8926), .A2(n8944), .ZN(n8927) );
  OAI211_X1 U10274 ( .C1(n8929), .C2(n8952), .A(n8928), .B(n8927), .ZN(
        P2_U3447) );
  INV_X1 U10275 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8931) );
  MUX2_X1 U10276 ( .A(n8931), .B(n8930), .S(n9937), .Z(n8934) );
  NAND2_X1 U10277 ( .A1(n8932), .A2(n8944), .ZN(n8933) );
  OAI211_X1 U10278 ( .C1(n8935), .C2(n8952), .A(n8934), .B(n8933), .ZN(
        P2_U3446) );
  INV_X1 U10279 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8937) );
  MUX2_X1 U10280 ( .A(n8937), .B(n8936), .S(n9937), .Z(n8940) );
  NAND2_X1 U10281 ( .A1(n8938), .A2(n8944), .ZN(n8939) );
  OAI211_X1 U10282 ( .C1(n8941), .C2(n8952), .A(n8940), .B(n8939), .ZN(
        P2_U3444) );
  INV_X1 U10283 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8943) );
  MUX2_X1 U10284 ( .A(n8943), .B(n8942), .S(n9937), .Z(n8947) );
  NAND2_X1 U10285 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  OAI211_X1 U10286 ( .C1(n8948), .C2(n8952), .A(n8947), .B(n8946), .ZN(
        P2_U3441) );
  INV_X1 U10287 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8950) );
  MUX2_X1 U10288 ( .A(n8950), .B(n8949), .S(n9937), .Z(n8951) );
  OAI21_X1 U10289 ( .B1(n8953), .B2(n8952), .A(n8951), .ZN(P2_U3438) );
  INV_X1 U10290 ( .A(n8954), .ZN(n9689) );
  INV_X1 U10291 ( .A(n8955), .ZN(n8956) );
  NOR4_X1 U10292 ( .A1(n8956), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n4837), .ZN(n8957) );
  AOI21_X1 U10293 ( .B1(n8958), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8957), .ZN(
        n8959) );
  OAI21_X1 U10294 ( .B1(n9689), .B2(n8960), .A(n8959), .ZN(P2_U3264) );
  OAI222_X1 U10295 ( .A1(n8964), .A2(n8963), .B1(n8962), .B2(P2_U3151), .C1(
        n8961), .C2(n7957), .ZN(P2_U3266) );
  NAND2_X1 U10296 ( .A1(n8965), .A2(n8969), .ZN(n8967) );
  OAI211_X1 U10297 ( .C1(n7957), .C2(n8968), .A(n8967), .B(n8966), .ZN(
        P2_U3267) );
  NAND2_X1 U10298 ( .A1(n9690), .A2(n8969), .ZN(n8971) );
  OAI211_X1 U10299 ( .C1(n7957), .C2(n8972), .A(n8971), .B(n8970), .ZN(
        P2_U3268) );
  MUX2_X1 U10300 ( .A(n8973), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10301 ( .B1(n8975), .B2(n8974), .A(n4425), .ZN(n8983) );
  NAND2_X1 U10302 ( .A1(n9117), .A2(n9133), .ZN(n8976) );
  NAND2_X1 U10303 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9792) );
  OAI211_X1 U10304 ( .C1(n8977), .C2(n9119), .A(n8976), .B(n9792), .ZN(n8980)
         );
  NOR2_X1 U10305 ( .A1(n8978), .A2(n9124), .ZN(n8979) );
  AOI211_X1 U10306 ( .C1(n8981), .C2(n9121), .A(n8980), .B(n8979), .ZN(n8982)
         );
  OAI21_X1 U10307 ( .B1(n8983), .B2(n9098), .A(n8982), .ZN(P1_U3215) );
  AND3_X1 U10308 ( .A1(n8987), .A2(n8985), .A3(n8986), .ZN(n8988) );
  OAI21_X1 U10309 ( .B1(n8984), .B2(n8988), .A(n9115), .ZN(n8993) );
  NOR2_X1 U10310 ( .A1(n9107), .A2(n9391), .ZN(n8991) );
  OAI22_X1 U10311 ( .A1(n9382), .A2(n9119), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8989), .ZN(n8990) );
  AOI211_X1 U10312 ( .C1(n9117), .C2(n9130), .A(n8991), .B(n8990), .ZN(n8992)
         );
  OAI211_X1 U10313 ( .C1(n9652), .C2(n9124), .A(n8993), .B(n8992), .ZN(
        P1_U3216) );
  XNOR2_X1 U10314 ( .A(n8994), .B(n8995), .ZN(n9090) );
  NOR2_X1 U10315 ( .A1(n9090), .A2(n9089), .ZN(n9088) );
  AOI21_X1 U10316 ( .B1(n8995), .B2(n8994), .A(n9088), .ZN(n8999) );
  XNOR2_X1 U10317 ( .A(n8997), .B(n8996), .ZN(n8998) );
  XNOR2_X1 U10318 ( .A(n8999), .B(n8998), .ZN(n9005) );
  NOR2_X1 U10319 ( .A1(n9107), .A2(n9448), .ZN(n9003) );
  INV_X1 U10320 ( .A(n9060), .ZN(n9093) );
  AND2_X1 U10321 ( .A1(n9474), .A2(n9524), .ZN(n9000) );
  AOI21_X1 U10322 ( .B1(n9131), .B2(n9500), .A(n9000), .ZN(n9445) );
  OAI22_X1 U10323 ( .A1(n9093), .A2(n9445), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9001), .ZN(n9002) );
  AOI211_X1 U10324 ( .C1(n9587), .C2(n9096), .A(n9003), .B(n9002), .ZN(n9004)
         );
  OAI21_X1 U10325 ( .B1(n9005), .B2(n9098), .A(n9004), .ZN(P1_U3219) );
  OAI21_X1 U10326 ( .B1(n9008), .B2(n9007), .A(n9006), .ZN(n9009) );
  NAND2_X1 U10327 ( .A1(n9009), .A2(n9115), .ZN(n9015) );
  INV_X1 U10328 ( .A(n9010), .ZN(n9423) );
  AND2_X1 U10329 ( .A1(n9131), .A2(n9524), .ZN(n9011) );
  AOI21_X1 U10330 ( .B1(n9130), .B2(n9500), .A(n9011), .ZN(n9419) );
  OAI22_X1 U10331 ( .A1(n9419), .A2(n9093), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9012), .ZN(n9013) );
  AOI21_X1 U10332 ( .B1(n9423), .B2(n9121), .A(n9013), .ZN(n9014) );
  OAI211_X1 U10333 ( .C1(n9657), .C2(n9124), .A(n9015), .B(n9014), .ZN(
        P1_U3223) );
  OAI21_X1 U10334 ( .B1(n9017), .B2(n9016), .A(n9100), .ZN(n9018) );
  NAND2_X1 U10335 ( .A1(n9018), .A2(n9115), .ZN(n9022) );
  AOI22_X1 U10336 ( .A1(n9128), .A2(n9109), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9019) );
  OAI21_X1 U10337 ( .B1(n9382), .B2(n9083), .A(n9019), .ZN(n9020) );
  AOI21_X1 U10338 ( .B1(n9356), .B2(n9121), .A(n9020), .ZN(n9021) );
  OAI211_X1 U10339 ( .C1(n4701), .C2(n9124), .A(n9022), .B(n9021), .ZN(
        P1_U3225) );
  INV_X1 U10340 ( .A(n9026), .ZN(n9024) );
  NOR2_X1 U10341 ( .A1(n9023), .A2(n9024), .ZN(n9029) );
  AOI21_X1 U10342 ( .B1(n9027), .B2(n9026), .A(n9025), .ZN(n9028) );
  OAI21_X1 U10343 ( .B1(n9029), .B2(n9028), .A(n9115), .ZN(n9035) );
  OAI21_X1 U10344 ( .B1(n9119), .B2(n9031), .A(n9030), .ZN(n9033) );
  NOR2_X1 U10345 ( .A1(n9107), .A2(n9492), .ZN(n9032) );
  AOI211_X1 U10346 ( .C1(n9117), .C2(n9499), .A(n9033), .B(n9032), .ZN(n9034)
         );
  OAI211_X1 U10347 ( .C1(n9495), .C2(n9124), .A(n9035), .B(n9034), .ZN(
        P1_U3226) );
  OAI21_X1 U10348 ( .B1(n9038), .B2(n9037), .A(n9036), .ZN(n9039) );
  NAND2_X1 U10349 ( .A1(n9039), .A2(n9115), .ZN(n9045) );
  NAND2_X1 U10350 ( .A1(n9117), .A2(n9475), .ZN(n9041) );
  OAI211_X1 U10351 ( .C1(n9042), .C2(n9119), .A(n9041), .B(n9040), .ZN(n9043)
         );
  AOI21_X1 U10352 ( .B1(n9482), .B2(n9121), .A(n9043), .ZN(n9044) );
  OAI211_X1 U10353 ( .C1(n9664), .C2(n9124), .A(n9045), .B(n9044), .ZN(
        P1_U3228) );
  INV_X1 U10354 ( .A(n9046), .ZN(n9050) );
  NOR3_X1 U10355 ( .A1(n8984), .A2(n9048), .A3(n9047), .ZN(n9049) );
  OAI21_X1 U10356 ( .B1(n9050), .B2(n9049), .A(n9115), .ZN(n9054) );
  AOI22_X1 U10357 ( .A1(n9339), .A2(n9500), .B1(n9524), .B2(n9408), .ZN(n9365)
         );
  OAI22_X1 U10358 ( .A1(n9365), .A2(n9093), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9051), .ZN(n9052) );
  AOI21_X1 U10359 ( .B1(n9371), .B2(n9121), .A(n9052), .ZN(n9053) );
  OAI211_X1 U10360 ( .C1(n9370), .C2(n9124), .A(n9054), .B(n9053), .ZN(
        P1_U3229) );
  OAI211_X1 U10361 ( .C1(n9057), .C2(n9056), .A(n9055), .B(n9115), .ZN(n9067)
         );
  INV_X1 U10362 ( .A(n9058), .ZN(n9059) );
  AOI22_X1 U10363 ( .A1(n9060), .A2(n9059), .B1(P1_REG3_REG_4__SCAN_IN), .B2(
        P1_U3086), .ZN(n9066) );
  INV_X1 U10364 ( .A(n9061), .ZN(n9062) );
  NAND2_X1 U10365 ( .A1(n9121), .A2(n9062), .ZN(n9065) );
  NAND2_X1 U10366 ( .A1(n9096), .A2(n9063), .ZN(n9064) );
  NAND4_X1 U10367 ( .A1(n9067), .A2(n9066), .A3(n9065), .A4(n9064), .ZN(
        P1_U3230) );
  XNOR2_X1 U10368 ( .A(n9070), .B(n9069), .ZN(n9071) );
  XNOR2_X1 U10369 ( .A(n9068), .B(n9071), .ZN(n9077) );
  AND2_X1 U10370 ( .A1(n9132), .A2(n9524), .ZN(n9072) );
  AOI21_X1 U10371 ( .B1(n9407), .B2(n9500), .A(n9072), .ZN(n9432) );
  OAI22_X1 U10372 ( .A1(n9432), .A2(n9093), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9073), .ZN(n9075) );
  NOR2_X1 U10373 ( .A1(n9439), .A2(n9124), .ZN(n9074) );
  AOI211_X1 U10374 ( .C1(n9436), .C2(n9121), .A(n9075), .B(n9074), .ZN(n9076)
         );
  OAI21_X1 U10375 ( .B1(n9077), .B2(n9098), .A(n9076), .ZN(P1_U3233) );
  INV_X1 U10376 ( .A(n8985), .ZN(n9079) );
  AOI21_X1 U10377 ( .B1(n9080), .B2(n9078), .A(n9079), .ZN(n9087) );
  AOI22_X1 U10378 ( .A1(n9109), .A2(n9408), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9082) );
  NAND2_X1 U10379 ( .A1(n9121), .A2(n9401), .ZN(n9081) );
  OAI211_X1 U10380 ( .C1(n9084), .C2(n9083), .A(n9082), .B(n9081), .ZN(n9085)
         );
  AOI21_X1 U10381 ( .B1(n9571), .B2(n9096), .A(n9085), .ZN(n9086) );
  OAI21_X1 U10382 ( .B1(n9087), .B2(n9098), .A(n9086), .ZN(P1_U3235) );
  AOI21_X1 U10383 ( .B1(n9090), .B2(n9089), .A(n9088), .ZN(n9099) );
  NOR2_X1 U10384 ( .A1(n9107), .A2(n9462), .ZN(n9095) );
  AND2_X1 U10385 ( .A1(n9501), .A2(n9524), .ZN(n9091) );
  AOI21_X1 U10386 ( .B1(n9132), .B2(n9500), .A(n9091), .ZN(n9458) );
  OAI22_X1 U10387 ( .A1(n9093), .A2(n9458), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9092), .ZN(n9094) );
  AOI211_X1 U10388 ( .C1(n9592), .C2(n9096), .A(n9095), .B(n9094), .ZN(n9097)
         );
  OAI21_X1 U10389 ( .B1(n9099), .B2(n9098), .A(n9097), .ZN(P1_U3238) );
  INV_X1 U10390 ( .A(n9549), .ZN(n9335) );
  INV_X1 U10391 ( .A(n9100), .ZN(n9103) );
  NAND3_X1 U10392 ( .A1(n9105), .A2(n9115), .A3(n9104), .ZN(n9111) );
  AOI22_X1 U10393 ( .A1(n9339), .A2(n9117), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9106) );
  OAI21_X1 U10394 ( .B1(n9107), .B2(n9332), .A(n9106), .ZN(n9108) );
  AOI21_X1 U10395 ( .B1(n9340), .B2(n9109), .A(n9108), .ZN(n9110) );
  OAI211_X1 U10396 ( .C1(n9335), .C2(n9124), .A(n9111), .B(n9110), .ZN(
        P1_U3240) );
  OAI21_X1 U10397 ( .B1(n9112), .B2(n9114), .A(n9113), .ZN(n9116) );
  NAND2_X1 U10398 ( .A1(n9116), .A2(n9115), .ZN(n9123) );
  NAND2_X1 U10399 ( .A1(n9117), .A2(n9523), .ZN(n9118) );
  NAND2_X1 U10400 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9805) );
  OAI211_X1 U10401 ( .C1(n9517), .C2(n9119), .A(n9118), .B(n9805), .ZN(n9120)
         );
  AOI21_X1 U10402 ( .B1(n9512), .B2(n9121), .A(n9120), .ZN(n9122) );
  OAI211_X1 U10403 ( .C1(n9515), .C2(n9124), .A(n9123), .B(n9122), .ZN(
        P1_U3241) );
  MUX2_X1 U10404 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9125), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10405 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9126), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10406 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9127), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10407 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9340), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10408 ( .A(n9128), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9144), .Z(
        P1_U3580) );
  MUX2_X1 U10409 ( .A(n9339), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9144), .Z(
        P1_U3579) );
  MUX2_X1 U10410 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9129), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10411 ( .A(n9408), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9144), .Z(
        P1_U3577) );
  MUX2_X1 U10412 ( .A(n9130), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9144), .Z(
        P1_U3576) );
  MUX2_X1 U10413 ( .A(n9407), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9144), .Z(
        P1_U3575) );
  MUX2_X1 U10414 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9131), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10415 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9132), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10416 ( .A(n9474), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9144), .Z(
        P1_U3572) );
  MUX2_X1 U10417 ( .A(n9501), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9144), .Z(
        P1_U3571) );
  MUX2_X1 U10418 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9475), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10419 ( .A(n9499), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9144), .Z(
        P1_U3569) );
  MUX2_X1 U10420 ( .A(n9523), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9144), .Z(
        P1_U3568) );
  MUX2_X1 U10421 ( .A(n9133), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9144), .Z(
        P1_U3567) );
  MUX2_X1 U10422 ( .A(n9134), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9144), .Z(
        P1_U3566) );
  MUX2_X1 U10423 ( .A(n9135), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9144), .Z(
        P1_U3565) );
  MUX2_X1 U10424 ( .A(n9136), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9144), .Z(
        P1_U3564) );
  MUX2_X1 U10425 ( .A(n4726), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9144), .Z(
        P1_U3563) );
  MUX2_X1 U10426 ( .A(n9137), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9144), .Z(
        P1_U3562) );
  MUX2_X1 U10427 ( .A(n9138), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9144), .Z(
        P1_U3561) );
  MUX2_X1 U10428 ( .A(n9139), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9144), .Z(
        P1_U3560) );
  MUX2_X1 U10429 ( .A(n9140), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9144), .Z(
        P1_U3559) );
  MUX2_X1 U10430 ( .A(n9141), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9144), .Z(
        P1_U3558) );
  MUX2_X1 U10431 ( .A(n9142), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9144), .Z(
        P1_U3557) );
  MUX2_X1 U10432 ( .A(n9143), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9144), .Z(
        P1_U3556) );
  MUX2_X1 U10433 ( .A(n6487), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9144), .Z(
        P1_U3555) );
  OAI211_X1 U10434 ( .C1(n9147), .C2(n9146), .A(n9815), .B(n9145), .ZN(n9155)
         );
  OAI211_X1 U10435 ( .C1(n9150), .C2(n9149), .A(n9786), .B(n9148), .ZN(n9154)
         );
  AOI22_X1 U10436 ( .A1(n9746), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9153) );
  NAND2_X1 U10437 ( .A1(n9811), .A2(n9151), .ZN(n9152) );
  NAND4_X1 U10438 ( .A1(n9155), .A2(n9154), .A3(n9153), .A4(n9152), .ZN(
        P1_U3244) );
  NOR3_X1 U10439 ( .A1(n9156), .A2(n9738), .A3(n4352), .ZN(n9161) );
  NOR2_X1 U10440 ( .A1(n9691), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9157) );
  OR2_X1 U10441 ( .A1(n4352), .A2(n9157), .ZN(n9739) );
  INV_X1 U10442 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9741) );
  NAND2_X1 U10443 ( .A1(n9739), .A2(n9741), .ZN(n9744) );
  OAI211_X1 U10444 ( .C1(n9159), .C2(n9158), .A(P1_U3973), .B(n9744), .ZN(
        n9160) );
  OR2_X1 U10445 ( .A1(n9161), .A2(n9160), .ZN(n9200) );
  INV_X1 U10446 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9163) );
  OAI22_X1 U10447 ( .A1(n9823), .A2(n9163), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9162), .ZN(n9164) );
  AOI21_X1 U10448 ( .B1(n9165), .B2(n9811), .A(n9164), .ZN(n9174) );
  OAI211_X1 U10449 ( .C1(n9168), .C2(n9167), .A(n9786), .B(n9166), .ZN(n9173)
         );
  OAI211_X1 U10450 ( .C1(n9171), .C2(n9170), .A(n9815), .B(n9169), .ZN(n9172)
         );
  NAND4_X1 U10451 ( .A1(n9200), .A2(n9174), .A3(n9173), .A4(n9172), .ZN(
        P1_U3245) );
  INV_X1 U10452 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9176) );
  NAND2_X1 U10453 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9175) );
  OAI21_X1 U10454 ( .B1(n9823), .B2(n9176), .A(n9175), .ZN(n9177) );
  AOI21_X1 U10455 ( .B1(n9178), .B2(n9811), .A(n9177), .ZN(n9187) );
  OAI211_X1 U10456 ( .C1(n9181), .C2(n9180), .A(n9786), .B(n9179), .ZN(n9186)
         );
  OAI211_X1 U10457 ( .C1(n9184), .C2(n9183), .A(n9815), .B(n9182), .ZN(n9185)
         );
  NAND3_X1 U10458 ( .A1(n9187), .A2(n9186), .A3(n9185), .ZN(P1_U3246) );
  AND2_X1 U10459 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9190) );
  NOR2_X1 U10460 ( .A1(n9790), .A2(n9188), .ZN(n9189) );
  AOI211_X1 U10461 ( .C1(n9746), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9190), .B(
        n9189), .ZN(n9199) );
  OAI211_X1 U10462 ( .C1(n9193), .C2(n9192), .A(n9815), .B(n9191), .ZN(n9198)
         );
  OAI211_X1 U10463 ( .C1(n9196), .C2(n9195), .A(n9786), .B(n9194), .ZN(n9197)
         );
  NAND4_X1 U10464 ( .A1(n9200), .A2(n9199), .A3(n9198), .A4(n9197), .ZN(
        P1_U3247) );
  INV_X1 U10465 ( .A(n9201), .ZN(n9205) );
  INV_X1 U10466 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U10467 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9202) );
  OAI21_X1 U10468 ( .B1(n9823), .B2(n9203), .A(n9202), .ZN(n9204) );
  AOI21_X1 U10469 ( .B1(n9205), .B2(n9811), .A(n9204), .ZN(n9214) );
  OAI211_X1 U10470 ( .C1(n9208), .C2(n9207), .A(n9786), .B(n9206), .ZN(n9213)
         );
  OAI211_X1 U10471 ( .C1(n9211), .C2(n9210), .A(n9815), .B(n9209), .ZN(n9212)
         );
  NAND3_X1 U10472 ( .A1(n9214), .A2(n9213), .A3(n9212), .ZN(P1_U3248) );
  INV_X1 U10473 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9216) );
  NAND2_X1 U10474 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9215) );
  OAI21_X1 U10475 ( .B1(n9823), .B2(n9216), .A(n9215), .ZN(n9217) );
  AOI21_X1 U10476 ( .B1(n9218), .B2(n9811), .A(n9217), .ZN(n9227) );
  OAI211_X1 U10477 ( .C1(n9221), .C2(n9220), .A(n9786), .B(n9219), .ZN(n9226)
         );
  OAI211_X1 U10478 ( .C1(n9224), .C2(n9223), .A(n9815), .B(n9222), .ZN(n9225)
         );
  NAND3_X1 U10479 ( .A1(n9227), .A2(n9226), .A3(n9225), .ZN(P1_U3249) );
  INV_X1 U10480 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U10481 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9228) );
  OAI21_X1 U10482 ( .B1(n9823), .B2(n9229), .A(n9228), .ZN(n9230) );
  AOI21_X1 U10483 ( .B1(n9231), .B2(n9811), .A(n9230), .ZN(n9240) );
  OAI211_X1 U10484 ( .C1(n9234), .C2(n9233), .A(n9815), .B(n9232), .ZN(n9239)
         );
  OAI211_X1 U10485 ( .C1(n9237), .C2(n9236), .A(n9786), .B(n9235), .ZN(n9238)
         );
  NAND3_X1 U10486 ( .A1(n9240), .A2(n9239), .A3(n9238), .ZN(P1_U3250) );
  INV_X1 U10487 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U10488 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9241) );
  OAI21_X1 U10489 ( .B1(n9823), .B2(n9242), .A(n9241), .ZN(n9243) );
  AOI21_X1 U10490 ( .B1(n9244), .B2(n9811), .A(n9243), .ZN(n9253) );
  OAI211_X1 U10491 ( .C1(n9247), .C2(n9246), .A(n9815), .B(n9245), .ZN(n9252)
         );
  OAI211_X1 U10492 ( .C1(n9250), .C2(n9249), .A(n9786), .B(n9248), .ZN(n9251)
         );
  NAND3_X1 U10493 ( .A1(n9253), .A2(n9252), .A3(n9251), .ZN(P1_U3251) );
  OR2_X1 U10494 ( .A1(n9259), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9254) );
  AND2_X1 U10495 ( .A1(n9255), .A2(n9254), .ZN(n9818) );
  NAND2_X1 U10496 ( .A1(n9812), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9257) );
  OR2_X1 U10497 ( .A1(n9812), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9256) );
  AND2_X1 U10498 ( .A1(n9257), .A2(n9256), .ZN(n9817) );
  NAND2_X1 U10499 ( .A1(n9818), .A2(n9817), .ZN(n9816) );
  NAND2_X1 U10500 ( .A1(n9816), .A2(n9257), .ZN(n9258) );
  XNOR2_X1 U10501 ( .A(n9258), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9268) );
  INV_X1 U10502 ( .A(n9268), .ZN(n9265) );
  OAI22_X1 U10503 ( .A1(n9261), .A2(n9260), .B1(P1_REG1_REG_17__SCAN_IN), .B2(
        n9259), .ZN(n9810) );
  NAND2_X1 U10504 ( .A1(n9812), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9262) );
  OAI21_X1 U10505 ( .B1(n9812), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9262), .ZN(
        n9809) );
  OR2_X1 U10506 ( .A1(n9810), .A2(n9809), .ZN(n9813) );
  NAND2_X1 U10507 ( .A1(n9813), .A2(n9262), .ZN(n9264) );
  XNOR2_X1 U10508 ( .A(n9264), .B(n9263), .ZN(n9266) );
  AOI22_X1 U10509 ( .A1(n9265), .A2(n9815), .B1(n9786), .B2(n9266), .ZN(n9271)
         );
  OAI21_X1 U10510 ( .B1(n9266), .B2(n9808), .A(n9790), .ZN(n9267) );
  AOI21_X1 U10511 ( .B1(n9815), .B2(n9268), .A(n9267), .ZN(n9270) );
  MUX2_X1 U10512 ( .A(n9271), .B(n9270), .S(n9269), .Z(n9273) );
  NAND2_X1 U10513 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9272) );
  OAI211_X1 U10514 ( .C1(n4709), .C2(n9823), .A(n9273), .B(n9272), .ZN(
        P1_U3262) );
  XNOR2_X1 U10515 ( .A(n9275), .B(n9274), .ZN(n9532) );
  NAND2_X1 U10516 ( .A1(n9532), .A2(n9276), .ZN(n9279) );
  AOI21_X1 U10517 ( .B1(n9826), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9277), .ZN(
        n9278) );
  OAI211_X1 U10518 ( .C1(n9638), .C2(n9514), .A(n9279), .B(n9278), .ZN(
        P1_U3263) );
  OAI22_X1 U10519 ( .A1(n9282), .A2(n9390), .B1(n9281), .B2(n9468), .ZN(n9283)
         );
  AOI21_X1 U10520 ( .B1(n9284), .B2(n9838), .A(n9283), .ZN(n9285) );
  OAI21_X1 U10521 ( .B1(n9286), .B2(n9841), .A(n9285), .ZN(n9287) );
  AOI21_X1 U10522 ( .B1(n9280), .B2(n9836), .A(n9287), .ZN(n9288) );
  OAI21_X1 U10523 ( .B1(n9289), .B2(n9826), .A(n9288), .ZN(P1_U3356) );
  NAND2_X1 U10524 ( .A1(n9291), .A2(n9301), .ZN(n9292) );
  NAND2_X1 U10525 ( .A1(n9290), .A2(n9292), .ZN(n9535) );
  INV_X1 U10526 ( .A(n9293), .ZN(n9295) );
  OAI22_X1 U10527 ( .A1(n9295), .A2(n9390), .B1(n9294), .B2(n9468), .ZN(n9298)
         );
  NAND2_X1 U10528 ( .A1(n9536), .A2(n9319), .ZN(n9296) );
  NAND3_X1 U10529 ( .A1(n4367), .A2(n9531), .A3(n9296), .ZN(n9538) );
  NOR2_X1 U10530 ( .A1(n9538), .A2(n9841), .ZN(n9297) );
  AOI211_X1 U10531 ( .C1(n9838), .C2(n9536), .A(n9298), .B(n9297), .ZN(n9309)
         );
  OAI21_X1 U10532 ( .B1(n9301), .B2(n9300), .A(n9299), .ZN(n9302) );
  NAND2_X1 U10533 ( .A1(n9302), .A2(n9503), .ZN(n9307) );
  OAI22_X1 U10534 ( .A1(n9304), .A2(n9380), .B1(n9303), .B2(n9516), .ZN(n9305)
         );
  INV_X1 U10535 ( .A(n9305), .ZN(n9306) );
  NAND2_X1 U10536 ( .A1(n9307), .A2(n9306), .ZN(n9540) );
  NAND2_X1 U10537 ( .A1(n9540), .A2(n9468), .ZN(n9308) );
  OAI211_X1 U10538 ( .C1(n9535), .C2(n9529), .A(n9309), .B(n9308), .ZN(
        P1_U3265) );
  XNOR2_X1 U10539 ( .A(n9310), .B(n9313), .ZN(n9545) );
  INV_X1 U10540 ( .A(n9545), .ZN(n9328) );
  OAI21_X1 U10541 ( .B1(n9313), .B2(n9312), .A(n9311), .ZN(n9314) );
  NAND2_X1 U10542 ( .A1(n9314), .A2(n9503), .ZN(n9318) );
  OAI22_X1 U10543 ( .A1(n9315), .A2(n9516), .B1(n9350), .B2(n9380), .ZN(n9316)
         );
  INV_X1 U10544 ( .A(n9316), .ZN(n9317) );
  NAND2_X1 U10545 ( .A1(n9318), .A2(n9317), .ZN(n9543) );
  INV_X1 U10546 ( .A(n9331), .ZN(n9321) );
  INV_X1 U10547 ( .A(n9319), .ZN(n9320) );
  AOI211_X1 U10548 ( .C1(n9322), .C2(n9321), .A(n9510), .B(n9320), .ZN(n9544)
         );
  NAND2_X1 U10549 ( .A1(n9544), .A2(n9527), .ZN(n9325) );
  AOI22_X1 U10550 ( .A1(n9323), .A2(n9834), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9826), .ZN(n9324) );
  OAI211_X1 U10551 ( .C1(n9643), .C2(n9514), .A(n9325), .B(n9324), .ZN(n9326)
         );
  AOI21_X1 U10552 ( .B1(n9468), .B2(n9543), .A(n9326), .ZN(n9327) );
  OAI21_X1 U10553 ( .B1(n9328), .B2(n9529), .A(n9327), .ZN(P1_U3266) );
  XNOR2_X1 U10554 ( .A(n9329), .B(n9330), .ZN(n9552) );
  AOI211_X1 U10555 ( .C1(n9549), .C2(n9353), .A(n9510), .B(n9331), .ZN(n9548)
         );
  INV_X1 U10556 ( .A(n9332), .ZN(n9333) );
  AOI22_X1 U10557 ( .A1(n9333), .A2(n9834), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9826), .ZN(n9334) );
  OAI21_X1 U10558 ( .B1(n9335), .B2(n9514), .A(n9334), .ZN(n9343) );
  OAI21_X1 U10559 ( .B1(n9338), .B2(n9337), .A(n9336), .ZN(n9341) );
  AOI222_X1 U10560 ( .A1(n9503), .A2(n9341), .B1(n9340), .B2(n9500), .C1(n9339), .C2(n9524), .ZN(n9551) );
  NOR2_X1 U10561 ( .A1(n9551), .A2(n9826), .ZN(n9342) );
  AOI211_X1 U10562 ( .C1(n9548), .C2(n9527), .A(n9343), .B(n9342), .ZN(n9344)
         );
  OAI21_X1 U10563 ( .B1(n9529), .B2(n9552), .A(n9344), .ZN(P1_U3267) );
  XOR2_X1 U10564 ( .A(n9346), .B(n9345), .Z(n9555) );
  INV_X1 U10565 ( .A(n9555), .ZN(n9361) );
  NAND2_X1 U10566 ( .A1(n9347), .A2(n9346), .ZN(n9348) );
  AOI21_X1 U10567 ( .B1(n9349), .B2(n9348), .A(n9518), .ZN(n9352) );
  OAI22_X1 U10568 ( .A1(n9350), .A2(n9516), .B1(n9382), .B2(n9380), .ZN(n9351)
         );
  OR2_X1 U10569 ( .A1(n9352), .A2(n9351), .ZN(n9553) );
  INV_X1 U10570 ( .A(n9353), .ZN(n9354) );
  AOI211_X1 U10571 ( .C1(n9355), .C2(n9369), .A(n9510), .B(n9354), .ZN(n9554)
         );
  NAND2_X1 U10572 ( .A1(n9554), .A2(n9527), .ZN(n9358) );
  AOI22_X1 U10573 ( .A1(n9356), .A2(n9834), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9826), .ZN(n9357) );
  OAI211_X1 U10574 ( .C1(n4701), .C2(n9514), .A(n9358), .B(n9357), .ZN(n9359)
         );
  AOI21_X1 U10575 ( .B1(n9468), .B2(n9553), .A(n9359), .ZN(n9360) );
  OAI21_X1 U10576 ( .B1(n9361), .B2(n9529), .A(n9360), .ZN(P1_U3268) );
  AND2_X1 U10577 ( .A1(n9377), .A2(n9362), .ZN(n9364) );
  OAI211_X1 U10578 ( .C1(n9364), .C2(n9368), .A(n9363), .B(n9503), .ZN(n9366)
         );
  AND2_X1 U10579 ( .A1(n9366), .A2(n9365), .ZN(n9563) );
  NAND2_X1 U10580 ( .A1(n9367), .A2(n9368), .ZN(n9558) );
  NAND3_X1 U10581 ( .A1(n9559), .A2(n9558), .A3(n9836), .ZN(n9376) );
  OAI211_X1 U10582 ( .C1(n9370), .C2(n4417), .A(n9531), .B(n9369), .ZN(n9562)
         );
  AOI22_X1 U10583 ( .A1(n9371), .A2(n9834), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9826), .ZN(n9373) );
  NAND2_X1 U10584 ( .A1(n9560), .A2(n9838), .ZN(n9372) );
  OAI211_X1 U10585 ( .C1(n9562), .C2(n9841), .A(n9373), .B(n9372), .ZN(n9374)
         );
  INV_X1 U10586 ( .A(n9374), .ZN(n9375) );
  OAI211_X1 U10587 ( .C1(n9826), .C2(n9563), .A(n9376), .B(n9375), .ZN(
        P1_U3269) );
  OAI21_X1 U10588 ( .B1(n9387), .B2(n9378), .A(n9377), .ZN(n9379) );
  NAND2_X1 U10589 ( .A1(n9379), .A2(n9503), .ZN(n9385) );
  OAI22_X1 U10590 ( .A1(n9382), .A2(n9516), .B1(n9381), .B2(n9380), .ZN(n9383)
         );
  INV_X1 U10591 ( .A(n9383), .ZN(n9384) );
  NAND2_X1 U10592 ( .A1(n9385), .A2(n9384), .ZN(n9565) );
  INV_X1 U10593 ( .A(n9565), .ZN(n9396) );
  XNOR2_X1 U10594 ( .A(n9386), .B(n9387), .ZN(n9567) );
  NAND2_X1 U10595 ( .A1(n9567), .A2(n9836), .ZN(n9395) );
  AOI211_X1 U10596 ( .C1(n9388), .C2(n9399), .A(n9510), .B(n4417), .ZN(n9566)
         );
  NOR2_X1 U10597 ( .A1(n9652), .A2(n9514), .ZN(n9393) );
  OAI22_X1 U10598 ( .A1(n9391), .A2(n9390), .B1(n9468), .B2(n9389), .ZN(n9392)
         );
  AOI211_X1 U10599 ( .C1(n9566), .C2(n9527), .A(n9393), .B(n9392), .ZN(n9394)
         );
  OAI211_X1 U10600 ( .C1(n9826), .C2(n9396), .A(n9395), .B(n9394), .ZN(
        P1_U3270) );
  XNOR2_X1 U10601 ( .A(n9397), .B(n9406), .ZN(n9574) );
  INV_X1 U10602 ( .A(n9399), .ZN(n9400) );
  AOI211_X1 U10603 ( .C1(n9571), .C2(n9421), .A(n9510), .B(n9400), .ZN(n9570)
         );
  AOI22_X1 U10604 ( .A1(n9401), .A2(n9834), .B1(n9826), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9402) );
  OAI21_X1 U10605 ( .B1(n9403), .B2(n9514), .A(n9402), .ZN(n9411) );
  OAI21_X1 U10606 ( .B1(n9406), .B2(n9405), .A(n9404), .ZN(n9409) );
  AOI222_X1 U10607 ( .A1(n9503), .A2(n9409), .B1(n9408), .B2(n9500), .C1(n9407), .C2(n9524), .ZN(n9573) );
  NOR2_X1 U10608 ( .A1(n9573), .A2(n9826), .ZN(n9410) );
  AOI211_X1 U10609 ( .C1(n9570), .C2(n9527), .A(n9411), .B(n9410), .ZN(n9412)
         );
  OAI21_X1 U10610 ( .B1(n9574), .B2(n9529), .A(n9412), .ZN(P1_U3271) );
  XNOR2_X1 U10611 ( .A(n9413), .B(n4509), .ZN(n9577) );
  INV_X1 U10612 ( .A(n9577), .ZN(n9428) );
  NAND2_X1 U10613 ( .A1(n9415), .A2(n9414), .ZN(n9416) );
  NAND2_X1 U10614 ( .A1(n9417), .A2(n9416), .ZN(n9418) );
  NAND2_X1 U10615 ( .A1(n9418), .A2(n9503), .ZN(n9420) );
  NAND2_X1 U10616 ( .A1(n9420), .A2(n9419), .ZN(n9575) );
  AOI211_X1 U10617 ( .C1(n9422), .C2(n9434), .A(n9510), .B(n9398), .ZN(n9576)
         );
  NAND2_X1 U10618 ( .A1(n9576), .A2(n9527), .ZN(n9425) );
  AOI22_X1 U10619 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n9826), .B1(n9423), .B2(
        n9834), .ZN(n9424) );
  OAI211_X1 U10620 ( .C1(n9657), .C2(n9514), .A(n9425), .B(n9424), .ZN(n9426)
         );
  AOI21_X1 U10621 ( .B1(n9468), .B2(n9575), .A(n9426), .ZN(n9427) );
  OAI21_X1 U10622 ( .B1(n9428), .B2(n9529), .A(n9427), .ZN(P1_U3272) );
  XNOR2_X1 U10623 ( .A(n9429), .B(n9430), .ZN(n9584) );
  XNOR2_X1 U10624 ( .A(n9431), .B(n9430), .ZN(n9433) );
  OAI21_X1 U10625 ( .B1(n9433), .B2(n9518), .A(n9432), .ZN(n9580) );
  INV_X1 U10626 ( .A(n9434), .ZN(n9435) );
  AOI211_X1 U10627 ( .C1(n9582), .C2(n4707), .A(n9510), .B(n9435), .ZN(n9581)
         );
  NAND2_X1 U10628 ( .A1(n9581), .A2(n9527), .ZN(n9438) );
  AOI22_X1 U10629 ( .A1(n9826), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9436), .B2(
        n9834), .ZN(n9437) );
  OAI211_X1 U10630 ( .C1(n9439), .C2(n9514), .A(n9438), .B(n9437), .ZN(n9440)
         );
  AOI21_X1 U10631 ( .B1(n9468), .B2(n9580), .A(n9440), .ZN(n9441) );
  OAI21_X1 U10632 ( .B1(n9584), .B2(n9529), .A(n9441), .ZN(P1_U3273) );
  XNOR2_X1 U10633 ( .A(n9442), .B(n9443), .ZN(n9589) );
  XNOR2_X1 U10634 ( .A(n9444), .B(n9443), .ZN(n9446) );
  OAI21_X1 U10635 ( .B1(n9446), .B2(n9518), .A(n9445), .ZN(n9585) );
  AOI211_X1 U10636 ( .C1(n9587), .C2(n9460), .A(n9510), .B(n9447), .ZN(n9586)
         );
  NAND2_X1 U10637 ( .A1(n9586), .A2(n9527), .ZN(n9451) );
  INV_X1 U10638 ( .A(n9448), .ZN(n9449) );
  AOI22_X1 U10639 ( .A1(n9826), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9449), .B2(
        n9834), .ZN(n9450) );
  OAI211_X1 U10640 ( .C1(n9452), .C2(n9514), .A(n9451), .B(n9450), .ZN(n9453)
         );
  AOI21_X1 U10641 ( .B1(n9468), .B2(n9585), .A(n9453), .ZN(n9454) );
  OAI21_X1 U10642 ( .B1(n9589), .B2(n9529), .A(n9454), .ZN(P1_U3274) );
  XNOR2_X1 U10643 ( .A(n9455), .B(n9456), .ZN(n9594) );
  XNOR2_X1 U10644 ( .A(n9457), .B(n9456), .ZN(n9459) );
  OAI21_X1 U10645 ( .B1(n9459), .B2(n9518), .A(n9458), .ZN(n9590) );
  INV_X1 U10646 ( .A(n9592), .ZN(n9466) );
  INV_X1 U10647 ( .A(n9460), .ZN(n9461) );
  AOI211_X1 U10648 ( .C1(n9592), .C2(n9478), .A(n9510), .B(n9461), .ZN(n9591)
         );
  NAND2_X1 U10649 ( .A1(n9591), .A2(n9527), .ZN(n9465) );
  INV_X1 U10650 ( .A(n9462), .ZN(n9463) );
  AOI22_X1 U10651 ( .A1(n9826), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9463), .B2(
        n9834), .ZN(n9464) );
  OAI211_X1 U10652 ( .C1(n9466), .C2(n9514), .A(n9465), .B(n9464), .ZN(n9467)
         );
  AOI21_X1 U10653 ( .B1(n9468), .B2(n9590), .A(n9467), .ZN(n9469) );
  OAI21_X1 U10654 ( .B1(n9594), .B2(n9529), .A(n9469), .ZN(P1_U3275) );
  XNOR2_X1 U10655 ( .A(n9470), .B(n9472), .ZN(n9597) );
  INV_X1 U10656 ( .A(n9597), .ZN(n9487) );
  XNOR2_X1 U10657 ( .A(n9472), .B(n9471), .ZN(n9473) );
  NAND2_X1 U10658 ( .A1(n9473), .A2(n9503), .ZN(n9477) );
  AOI22_X1 U10659 ( .A1(n9475), .A2(n9524), .B1(n9474), .B2(n9500), .ZN(n9476)
         );
  NAND2_X1 U10660 ( .A1(n9477), .A2(n9476), .ZN(n9595) );
  INV_X1 U10661 ( .A(n9490), .ZN(n9480) );
  INV_X1 U10662 ( .A(n9478), .ZN(n9479) );
  AOI211_X1 U10663 ( .C1(n9481), .C2(n9480), .A(n9510), .B(n9479), .ZN(n9596)
         );
  NAND2_X1 U10664 ( .A1(n9596), .A2(n9527), .ZN(n9484) );
  AOI22_X1 U10665 ( .A1(n9826), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9482), .B2(
        n9834), .ZN(n9483) );
  OAI211_X1 U10666 ( .C1(n9664), .C2(n9514), .A(n9484), .B(n9483), .ZN(n9485)
         );
  AOI21_X1 U10667 ( .B1(n9468), .B2(n9595), .A(n9485), .ZN(n9486) );
  OAI21_X1 U10668 ( .B1(n9487), .B2(n9529), .A(n9486), .ZN(P1_U3276) );
  XNOR2_X1 U10669 ( .A(n9488), .B(n9489), .ZN(n9604) );
  INV_X1 U10670 ( .A(n9509), .ZN(n9491) );
  AOI211_X1 U10671 ( .C1(n9601), .C2(n9491), .A(n9510), .B(n9490), .ZN(n9600)
         );
  INV_X1 U10672 ( .A(n9492), .ZN(n9493) );
  AOI22_X1 U10673 ( .A1(n9826), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9493), .B2(
        n9834), .ZN(n9494) );
  OAI21_X1 U10674 ( .B1(n9495), .B2(n9514), .A(n9494), .ZN(n9505) );
  OAI21_X1 U10675 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9502) );
  AOI222_X1 U10676 ( .A1(n9503), .A2(n9502), .B1(n9501), .B2(n9500), .C1(n9499), .C2(n9524), .ZN(n9603) );
  NOR2_X1 U10677 ( .A1(n9603), .A2(n9826), .ZN(n9504) );
  AOI211_X1 U10678 ( .C1(n9600), .C2(n9527), .A(n9505), .B(n9504), .ZN(n9506)
         );
  OAI21_X1 U10679 ( .B1(n9529), .B2(n9604), .A(n9506), .ZN(P1_U3277) );
  XOR2_X1 U10680 ( .A(n9507), .B(n9520), .Z(n9609) );
  INV_X1 U10681 ( .A(n9508), .ZN(n9511) );
  AOI211_X1 U10682 ( .C1(n9606), .C2(n9511), .A(n9510), .B(n9509), .ZN(n9605)
         );
  AOI22_X1 U10683 ( .A1(n9826), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9512), .B2(
        n9834), .ZN(n9513) );
  OAI21_X1 U10684 ( .B1(n9515), .B2(n9514), .A(n9513), .ZN(n9526) );
  NOR2_X1 U10685 ( .A1(n9517), .A2(n9516), .ZN(n9522) );
  AOI211_X1 U10686 ( .C1(n9520), .C2(n9519), .A(n9518), .B(n4420), .ZN(n9521)
         );
  AOI211_X1 U10687 ( .C1(n9524), .C2(n9523), .A(n9522), .B(n9521), .ZN(n9608)
         );
  NOR2_X1 U10688 ( .A1(n9608), .A2(n9826), .ZN(n9525) );
  AOI211_X1 U10689 ( .C1(n9605), .C2(n9527), .A(n9526), .B(n9525), .ZN(n9528)
         );
  OAI21_X1 U10690 ( .B1(n9609), .B2(n9529), .A(n9528), .ZN(P1_U3278) );
  INV_X1 U10691 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9533) );
  AOI21_X1 U10692 ( .B1(n9532), .B2(n9531), .A(n9530), .ZN(n9635) );
  OAI21_X1 U10693 ( .B1(n9638), .B2(n9633), .A(n9534), .ZN(P1_U3553) );
  NAND2_X1 U10694 ( .A1(n9536), .A2(n9623), .ZN(n9537) );
  NAND2_X1 U10695 ( .A1(n9538), .A2(n9537), .ZN(n9539) );
  NOR2_X1 U10696 ( .A1(n9540), .A2(n9539), .ZN(n9541) );
  NAND2_X1 U10697 ( .A1(n9542), .A2(n9541), .ZN(n9639) );
  MUX2_X1 U10698 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9639), .S(n9876), .Z(
        P1_U3550) );
  INV_X1 U10699 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9546) );
  AOI211_X1 U10700 ( .C1(n9545), .C2(n9869), .A(n9544), .B(n9543), .ZN(n9640)
         );
  MUX2_X1 U10701 ( .A(n9546), .B(n9640), .S(n9876), .Z(n9547) );
  OAI21_X1 U10702 ( .B1(n9643), .B2(n9633), .A(n9547), .ZN(P1_U3549) );
  AOI21_X1 U10703 ( .B1(n9623), .B2(n9549), .A(n9548), .ZN(n9550) );
  OAI211_X1 U10704 ( .C1(n9552), .C2(n9625), .A(n9551), .B(n9550), .ZN(n9644)
         );
  MUX2_X1 U10705 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9644), .S(n9876), .Z(
        P1_U3548) );
  INV_X1 U10706 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9556) );
  AOI211_X1 U10707 ( .C1(n9555), .C2(n9869), .A(n9554), .B(n9553), .ZN(n9645)
         );
  MUX2_X1 U10708 ( .A(n9556), .B(n9645), .S(n9876), .Z(n9557) );
  OAI21_X1 U10709 ( .B1(n4701), .B2(n9633), .A(n9557), .ZN(P1_U3547) );
  NAND3_X1 U10710 ( .A1(n9559), .A2(n9558), .A3(n9869), .ZN(n9564) );
  NAND2_X1 U10711 ( .A1(n9560), .A2(n9623), .ZN(n9561) );
  NAND4_X1 U10712 ( .A1(n9564), .A2(n9563), .A3(n9562), .A4(n9561), .ZN(n9648)
         );
  MUX2_X1 U10713 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9648), .S(n9876), .Z(
        P1_U3546) );
  INV_X1 U10714 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9568) );
  AOI211_X1 U10715 ( .C1(n9567), .C2(n9869), .A(n9566), .B(n9565), .ZN(n9649)
         );
  MUX2_X1 U10716 ( .A(n9568), .B(n9649), .S(n9876), .Z(n9569) );
  OAI21_X1 U10717 ( .B1(n9652), .B2(n9633), .A(n9569), .ZN(P1_U3545) );
  AOI21_X1 U10718 ( .B1(n9623), .B2(n9571), .A(n9570), .ZN(n9572) );
  OAI211_X1 U10719 ( .C1(n9574), .C2(n9625), .A(n9573), .B(n9572), .ZN(n9653)
         );
  MUX2_X1 U10720 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9653), .S(n9876), .Z(
        P1_U3544) );
  INV_X1 U10721 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9578) );
  AOI211_X1 U10722 ( .C1(n9577), .C2(n9869), .A(n9576), .B(n9575), .ZN(n9654)
         );
  MUX2_X1 U10723 ( .A(n9578), .B(n9654), .S(n9876), .Z(n9579) );
  OAI21_X1 U10724 ( .B1(n9657), .B2(n9633), .A(n9579), .ZN(P1_U3543) );
  AOI211_X1 U10725 ( .C1(n9623), .C2(n9582), .A(n9581), .B(n9580), .ZN(n9583)
         );
  OAI21_X1 U10726 ( .B1(n9584), .B2(n9625), .A(n9583), .ZN(n9658) );
  MUX2_X1 U10727 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9658), .S(n9876), .Z(
        P1_U3542) );
  AOI211_X1 U10728 ( .C1(n9623), .C2(n9587), .A(n9586), .B(n9585), .ZN(n9588)
         );
  OAI21_X1 U10729 ( .B1(n9589), .B2(n9625), .A(n9588), .ZN(n9659) );
  MUX2_X1 U10730 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9659), .S(n9876), .Z(
        P1_U3541) );
  AOI211_X1 U10731 ( .C1(n9623), .C2(n9592), .A(n9591), .B(n9590), .ZN(n9593)
         );
  OAI21_X1 U10732 ( .B1(n9594), .B2(n9625), .A(n9593), .ZN(n9660) );
  MUX2_X1 U10733 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9660), .S(n9876), .Z(
        P1_U3540) );
  AOI211_X1 U10734 ( .C1(n9597), .C2(n9869), .A(n9596), .B(n9595), .ZN(n9661)
         );
  MUX2_X1 U10735 ( .A(n9598), .B(n9661), .S(n9876), .Z(n9599) );
  OAI21_X1 U10736 ( .B1(n9664), .B2(n9633), .A(n9599), .ZN(P1_U3539) );
  AOI21_X1 U10737 ( .B1(n9623), .B2(n9601), .A(n9600), .ZN(n9602) );
  OAI211_X1 U10738 ( .C1(n9604), .C2(n9625), .A(n9603), .B(n9602), .ZN(n9665)
         );
  MUX2_X1 U10739 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9665), .S(n9876), .Z(
        P1_U3538) );
  AOI21_X1 U10740 ( .B1(n9623), .B2(n9606), .A(n9605), .ZN(n9607) );
  OAI211_X1 U10741 ( .C1(n9609), .C2(n9625), .A(n9608), .B(n9607), .ZN(n9666)
         );
  MUX2_X1 U10742 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9666), .S(n9876), .Z(
        P1_U3537) );
  AOI21_X1 U10743 ( .B1(n9623), .B2(n9611), .A(n9610), .ZN(n9612) );
  OAI211_X1 U10744 ( .C1(n9614), .C2(n9625), .A(n9613), .B(n9612), .ZN(n9667)
         );
  MUX2_X1 U10745 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9667), .S(n9876), .Z(
        P1_U3536) );
  AOI211_X1 U10746 ( .C1(n9617), .C2(n9869), .A(n9616), .B(n9615), .ZN(n9668)
         );
  MUX2_X1 U10747 ( .A(n9618), .B(n9668), .S(n9876), .Z(n9619) );
  OAI21_X1 U10748 ( .B1(n9671), .B2(n9633), .A(n9619), .ZN(P1_U3535) );
  AOI211_X1 U10749 ( .C1(n9623), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9624)
         );
  OAI21_X1 U10750 ( .B1(n9626), .B2(n9625), .A(n9624), .ZN(n9672) );
  MUX2_X1 U10751 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9672), .S(n9876), .Z(
        P1_U3534) );
  INV_X1 U10752 ( .A(n9627), .ZN(n9848) );
  AOI211_X1 U10753 ( .C1(n9848), .C2(n9630), .A(n9629), .B(n9628), .ZN(n9673)
         );
  MUX2_X1 U10754 ( .A(n9631), .B(n9673), .S(n9876), .Z(n9632) );
  OAI21_X1 U10755 ( .B1(n9677), .B2(n9633), .A(n9632), .ZN(P1_U3533) );
  MUX2_X1 U10756 ( .A(n9634), .B(P1_REG1_REG_0__SCAN_IN), .S(n6362), .Z(
        P1_U3522) );
  INV_X1 U10757 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9636) );
  OAI21_X1 U10758 ( .B1(n9638), .B2(n9676), .A(n9637), .ZN(P1_U3521) );
  MUX2_X1 U10759 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9639), .S(n9871), .Z(
        P1_U3518) );
  INV_X1 U10760 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9641) );
  MUX2_X1 U10761 ( .A(n9641), .B(n9640), .S(n9871), .Z(n9642) );
  OAI21_X1 U10762 ( .B1(n9643), .B2(n9676), .A(n9642), .ZN(P1_U3517) );
  MUX2_X1 U10763 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9644), .S(n9871), .Z(
        P1_U3516) );
  INV_X1 U10764 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9646) );
  MUX2_X1 U10765 ( .A(n9646), .B(n9645), .S(n9871), .Z(n9647) );
  OAI21_X1 U10766 ( .B1(n4701), .B2(n9676), .A(n9647), .ZN(P1_U3515) );
  MUX2_X1 U10767 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9648), .S(n9871), .Z(
        P1_U3514) );
  INV_X1 U10768 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9650) );
  MUX2_X1 U10769 ( .A(n9650), .B(n9649), .S(n9871), .Z(n9651) );
  OAI21_X1 U10770 ( .B1(n9652), .B2(n9676), .A(n9651), .ZN(P1_U3513) );
  MUX2_X1 U10771 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9653), .S(n9871), .Z(
        P1_U3512) );
  INV_X1 U10772 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9655) );
  MUX2_X1 U10773 ( .A(n9655), .B(n9654), .S(n9871), .Z(n9656) );
  OAI21_X1 U10774 ( .B1(n9657), .B2(n9676), .A(n9656), .ZN(P1_U3511) );
  MUX2_X1 U10775 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9658), .S(n9871), .Z(
        P1_U3510) );
  MUX2_X1 U10776 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9659), .S(n9871), .Z(
        P1_U3509) );
  MUX2_X1 U10777 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9660), .S(n9871), .Z(
        P1_U3507) );
  INV_X1 U10778 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9662) );
  MUX2_X1 U10779 ( .A(n9662), .B(n9661), .S(n9871), .Z(n9663) );
  OAI21_X1 U10780 ( .B1(n9664), .B2(n9676), .A(n9663), .ZN(P1_U3504) );
  MUX2_X1 U10781 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9665), .S(n9871), .Z(
        P1_U3501) );
  MUX2_X1 U10782 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9666), .S(n9871), .Z(
        P1_U3498) );
  MUX2_X1 U10783 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9667), .S(n9871), .Z(
        P1_U3495) );
  MUX2_X1 U10784 ( .A(n9669), .B(n9668), .S(n9871), .Z(n9670) );
  OAI21_X1 U10785 ( .B1(n9671), .B2(n9676), .A(n9670), .ZN(P1_U3492) );
  MUX2_X1 U10786 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9672), .S(n9871), .Z(
        P1_U3489) );
  MUX2_X1 U10787 ( .A(n9674), .B(n9673), .S(n9871), .Z(n9675) );
  OAI21_X1 U10788 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(P1_U3486) );
  MUX2_X1 U10789 ( .A(n9678), .B(P1_D_REG_1__SCAN_IN), .S(n9847), .Z(P1_U3440)
         );
  INV_X1 U10790 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9680) );
  AND2_X1 U10791 ( .A1(n9680), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9683) );
  NAND4_X1 U10792 ( .A1(n9683), .A2(P1_IR_REG_31__SCAN_IN), .A3(n9682), .A4(
        n9681), .ZN(n9685) );
  OAI22_X1 U10793 ( .A1(n9679), .A2(n9685), .B1(n9684), .B2(n9694), .ZN(n9686)
         );
  INV_X1 U10794 ( .A(n9686), .ZN(n9687) );
  OAI21_X1 U10795 ( .B1(n9689), .B2(n9688), .A(n9687), .ZN(P1_U3324) );
  INV_X1 U10796 ( .A(n9690), .ZN(n9692) );
  OAI222_X1 U10797 ( .A1(n9694), .A2(n9693), .B1(n9688), .B2(n9692), .C1(n9691), .C2(P1_U3086), .ZN(P1_U3328) );
  MUX2_X1 U10798 ( .A(n9695), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U10799 ( .A(n9696), .B(n9705), .ZN(n9723) );
  INV_X1 U10800 ( .A(n9723), .ZN(n9714) );
  INV_X1 U10801 ( .A(n9726), .ZN(n9700) );
  OAI22_X1 U10802 ( .A1(n9700), .A2(n9699), .B1(n9698), .B2(n9697), .ZN(n9713)
         );
  OR2_X1 U10803 ( .A1(n9702), .A2(n9701), .ZN(n9704) );
  NAND2_X1 U10804 ( .A1(n9704), .A2(n9703), .ZN(n9706) );
  XNOR2_X1 U10805 ( .A(n9706), .B(n9705), .ZN(n9707) );
  OAI222_X1 U10806 ( .A1(n9712), .A2(n9711), .B1(n9710), .B2(n9709), .C1(n9708), .C2(n9707), .ZN(n9724) );
  AOI211_X1 U10807 ( .C1(n9715), .C2(n9714), .A(n9713), .B(n9724), .ZN(n9717)
         );
  AOI22_X1 U10808 ( .A1(n9718), .A2(n8500), .B1(n9717), .B2(n9716), .ZN(
        P2_U3219) );
  AOI22_X1 U10809 ( .A1(n9720), .A2(n9933), .B1(n9932), .B2(n9719), .ZN(n9721)
         );
  AOI22_X1 U10810 ( .A1(n9950), .A2(n9732), .B1(n5995), .B2(n6277), .ZN(
        P2_U3474) );
  NOR2_X1 U10811 ( .A1(n9723), .A2(n9920), .ZN(n9725) );
  AOI211_X1 U10812 ( .C1(n9932), .C2(n9726), .A(n9725), .B(n9724), .ZN(n9734)
         );
  AOI22_X1 U10813 ( .A1(n9950), .A2(n9734), .B1(n8499), .B2(n6277), .ZN(
        P2_U3473) );
  NAND2_X1 U10814 ( .A1(n9727), .A2(n9933), .ZN(n9728) );
  OAI21_X1 U10815 ( .B1(n9729), .B2(n9925), .A(n9728), .ZN(n9730) );
  NOR2_X1 U10816 ( .A1(n9731), .A2(n9730), .ZN(n9736) );
  AOI22_X1 U10817 ( .A1(n9950), .A2(n9736), .B1(n8473), .B2(n6277), .ZN(
        P2_U3472) );
  INV_X1 U10818 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9733) );
  AOI22_X1 U10819 ( .A1(n9939), .A2(n9733), .B1(n9732), .B2(n9937), .ZN(
        P2_U3435) );
  INV_X1 U10820 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9735) );
  AOI22_X1 U10821 ( .A1(n9939), .A2(n9735), .B1(n9734), .B2(n9937), .ZN(
        P2_U3432) );
  INV_X1 U10822 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9737) );
  AOI22_X1 U10823 ( .A1(n9939), .A2(n9737), .B1(n9736), .B2(n9937), .ZN(
        P2_U3429) );
  XNOR2_X1 U10824 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10825 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U10826 ( .A1(n9738), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9740) );
  OR2_X1 U10827 ( .A1(n9739), .A2(n9740), .ZN(n9743) );
  INV_X1 U10828 ( .A(n9740), .ZN(n9742) );
  MUX2_X1 U10829 ( .A(n9743), .B(n9742), .S(n9741), .Z(n9745) );
  NAND2_X1 U10830 ( .A1(n9745), .A2(n9744), .ZN(n9748) );
  AOI22_X1 U10831 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9746), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9747) );
  OAI21_X1 U10832 ( .B1(n9749), .B2(n9748), .A(n9747), .ZN(P1_U3243) );
  INV_X1 U10833 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9764) );
  NOR2_X1 U10834 ( .A1(n9751), .A2(n9750), .ZN(n9752) );
  OR3_X1 U10835 ( .A1(n9753), .A2(n9752), .A3(n9798), .ZN(n9759) );
  NOR2_X1 U10836 ( .A1(n9755), .A2(n9754), .ZN(n9756) );
  OR3_X1 U10837 ( .A1(n9757), .A2(n9756), .A3(n9808), .ZN(n9758) );
  OAI211_X1 U10838 ( .C1(n9790), .C2(n9760), .A(n9759), .B(n9758), .ZN(n9761)
         );
  INV_X1 U10839 ( .A(n9761), .ZN(n9763) );
  NAND2_X1 U10840 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9762) );
  OAI211_X1 U10841 ( .C1(n9823), .C2(n9764), .A(n9763), .B(n9762), .ZN(
        P1_U3254) );
  INV_X1 U10842 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9776) );
  AOI211_X1 U10843 ( .C1(n9767), .C2(n9766), .A(n9765), .B(n9808), .ZN(n9772)
         );
  AOI211_X1 U10844 ( .C1(n9770), .C2(n9769), .A(n9768), .B(n9798), .ZN(n9771)
         );
  AOI211_X1 U10845 ( .C1(n9811), .C2(n9773), .A(n9772), .B(n9771), .ZN(n9775)
         );
  OAI211_X1 U10846 ( .C1(n9823), .C2(n9776), .A(n9775), .B(n9774), .ZN(
        P1_U3256) );
  INV_X1 U10847 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9794) );
  INV_X1 U10848 ( .A(n9777), .ZN(n9789) );
  AOI21_X1 U10849 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(n9781) );
  NAND2_X1 U10850 ( .A1(n9815), .A2(n9781), .ZN(n9788) );
  AOI21_X1 U10851 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(n9785) );
  NAND2_X1 U10852 ( .A1(n9786), .A2(n9785), .ZN(n9787) );
  OAI211_X1 U10853 ( .C1(n9790), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9791)
         );
  INV_X1 U10854 ( .A(n9791), .ZN(n9793) );
  OAI211_X1 U10855 ( .C1(n9823), .C2(n9794), .A(n9793), .B(n9792), .ZN(
        P1_U3257) );
  INV_X1 U10856 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9807) );
  AOI211_X1 U10857 ( .C1(n9797), .C2(n9796), .A(n9795), .B(n9808), .ZN(n9803)
         );
  AOI211_X1 U10858 ( .C1(n9801), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9802)
         );
  AOI211_X1 U10859 ( .C1(n9811), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9806)
         );
  OAI211_X1 U10860 ( .C1(n9823), .C2(n9807), .A(n9806), .B(n9805), .ZN(
        P1_U3258) );
  INV_X1 U10861 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10187) );
  AOI21_X1 U10862 ( .B1(n9810), .B2(n9809), .A(n9808), .ZN(n9814) );
  AOI22_X1 U10863 ( .A1(n9814), .A2(n9813), .B1(n9812), .B2(n9811), .ZN(n9820)
         );
  OAI211_X1 U10864 ( .C1(n9818), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9819)
         );
  AND2_X1 U10865 ( .A1(n9820), .A2(n9819), .ZN(n9822) );
  NAND2_X1 U10866 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9821) );
  OAI211_X1 U10867 ( .C1(n9823), .C2(n10187), .A(n9822), .B(n9821), .ZN(
        P1_U3261) );
  NAND2_X1 U10868 ( .A1(n9838), .A2(n9824), .ZN(n9828) );
  AOI22_X1 U10869 ( .A1(n9826), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9834), .B2(
        n9825), .ZN(n9827) );
  OAI211_X1 U10870 ( .C1(n9829), .C2(n9841), .A(n9828), .B(n9827), .ZN(n9830)
         );
  AOI21_X1 U10871 ( .B1(n9831), .B2(n9836), .A(n9830), .ZN(n9832) );
  OAI21_X1 U10872 ( .B1(n9826), .B2(n9833), .A(n9832), .ZN(P1_U3290) );
  AOI22_X1 U10873 ( .A1(n9834), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n9826), .ZN(n9845) );
  NAND2_X1 U10874 ( .A1(n9836), .A2(n9835), .ZN(n9840) );
  NAND2_X1 U10875 ( .A1(n9838), .A2(n9837), .ZN(n9839) );
  OAI211_X1 U10876 ( .C1(n9842), .C2(n9841), .A(n9840), .B(n9839), .ZN(n9843)
         );
  INV_X1 U10877 ( .A(n9843), .ZN(n9844) );
  OAI211_X1 U10878 ( .C1(n9826), .C2(n9846), .A(n9845), .B(n9844), .ZN(
        P1_U3292) );
  AND2_X1 U10879 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9847), .ZN(P1_U3294) );
  AND2_X1 U10880 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9847), .ZN(P1_U3295) );
  AND2_X1 U10881 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9847), .ZN(P1_U3296) );
  AND2_X1 U10882 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9847), .ZN(P1_U3297) );
  AND2_X1 U10883 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9847), .ZN(P1_U3298) );
  AND2_X1 U10884 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9847), .ZN(P1_U3299) );
  AND2_X1 U10885 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9847), .ZN(P1_U3300) );
  AND2_X1 U10886 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9847), .ZN(P1_U3301) );
  AND2_X1 U10887 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9847), .ZN(P1_U3302) );
  AND2_X1 U10888 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9847), .ZN(P1_U3303) );
  AND2_X1 U10889 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9847), .ZN(P1_U3304) );
  AND2_X1 U10890 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9847), .ZN(P1_U3305) );
  AND2_X1 U10891 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9847), .ZN(P1_U3306) );
  AND2_X1 U10892 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9847), .ZN(P1_U3307) );
  AND2_X1 U10893 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9847), .ZN(P1_U3308) );
  AND2_X1 U10894 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9847), .ZN(P1_U3309) );
  AND2_X1 U10895 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9847), .ZN(P1_U3310) );
  AND2_X1 U10896 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9847), .ZN(P1_U3311) );
  AND2_X1 U10897 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9847), .ZN(P1_U3312) );
  AND2_X1 U10898 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9847), .ZN(P1_U3313) );
  AND2_X1 U10899 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9847), .ZN(P1_U3314) );
  AND2_X1 U10900 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9847), .ZN(P1_U3315) );
  AND2_X1 U10901 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9847), .ZN(P1_U3316) );
  AND2_X1 U10902 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9847), .ZN(P1_U3317) );
  AND2_X1 U10903 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9847), .ZN(P1_U3318) );
  AND2_X1 U10904 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9847), .ZN(P1_U3319) );
  AND2_X1 U10905 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9847), .ZN(P1_U3320) );
  AND2_X1 U10906 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9847), .ZN(P1_U3321) );
  AND2_X1 U10907 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9847), .ZN(P1_U3322) );
  AND2_X1 U10908 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9847), .ZN(P1_U3323) );
  AND2_X1 U10909 ( .A1(n9849), .A2(n9848), .ZN(n9853) );
  OAI21_X1 U10910 ( .B1(n9851), .B2(n9866), .A(n9850), .ZN(n9852) );
  NOR3_X1 U10911 ( .A1(n9854), .A2(n9853), .A3(n9852), .ZN(n9872) );
  AOI22_X1 U10912 ( .A1(n9871), .A2(n9872), .B1(n5151), .B2(n6369), .ZN(
        P1_U3474) );
  OAI21_X1 U10913 ( .B1(n9856), .B2(n9866), .A(n9855), .ZN(n9858) );
  AOI211_X1 U10914 ( .C1(n9869), .C2(n9859), .A(n9858), .B(n9857), .ZN(n9873)
         );
  AOI22_X1 U10915 ( .A1(n9871), .A2(n9873), .B1(n5211), .B2(n6369), .ZN(
        P1_U3477) );
  OAI211_X1 U10916 ( .C1(n4691), .C2(n9866), .A(n9861), .B(n9860), .ZN(n9862)
         );
  AOI21_X1 U10917 ( .B1(n9869), .B2(n9863), .A(n9862), .ZN(n9874) );
  AOI22_X1 U10918 ( .A1(n9871), .A2(n9874), .B1(n5194), .B2(n6369), .ZN(
        P1_U3480) );
  OAI211_X1 U10919 ( .C1(n9867), .C2(n9866), .A(n9865), .B(n9864), .ZN(n9868)
         );
  AOI21_X1 U10920 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n9875) );
  AOI22_X1 U10921 ( .A1(n9871), .A2(n9875), .B1(n5260), .B2(n6369), .ZN(
        P1_U3483) );
  AOI22_X1 U10922 ( .A1(n9876), .A2(n9872), .B1(n5145), .B2(n6362), .ZN(
        P1_U3529) );
  AOI22_X1 U10923 ( .A1(n9876), .A2(n9873), .B1(n6460), .B2(n6362), .ZN(
        P1_U3530) );
  AOI22_X1 U10924 ( .A1(n9876), .A2(n9874), .B1(n5189), .B2(n6362), .ZN(
        P1_U3531) );
  AOI22_X1 U10925 ( .A1(n9876), .A2(n9875), .B1(n5253), .B2(n6362), .ZN(
        P1_U3532) );
  AOI22_X1 U10926 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n9877), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n9885) );
  INV_X1 U10927 ( .A(n9878), .ZN(n9882) );
  OAI21_X1 U10928 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9880), .A(n9879), .ZN(
        n9881) );
  OAI21_X1 U10929 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(n9884) );
  OAI211_X1 U10930 ( .C1(n9886), .C2(n4857), .A(n9885), .B(n9884), .ZN(
        P2_U3182) );
  INV_X1 U10931 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9890) );
  OAI22_X1 U10932 ( .A1(n9887), .A2(n9920), .B1(n6973), .B2(n9925), .ZN(n9888)
         );
  NOR2_X1 U10933 ( .A1(n9889), .A2(n9888), .ZN(n9940) );
  AOI22_X1 U10934 ( .A1(n9939), .A2(n9890), .B1(n9940), .B2(n9937), .ZN(
        P2_U3393) );
  INV_X1 U10935 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9896) );
  OAI22_X1 U10936 ( .A1(n9893), .A2(n9892), .B1(n9891), .B2(n9925), .ZN(n9894)
         );
  NOR2_X1 U10937 ( .A1(n9895), .A2(n9894), .ZN(n9941) );
  AOI22_X1 U10938 ( .A1(n9939), .A2(n9896), .B1(n9941), .B2(n9937), .ZN(
        P2_U3396) );
  INV_X1 U10939 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9902) );
  INV_X1 U10940 ( .A(n9897), .ZN(n9901) );
  OAI22_X1 U10941 ( .A1(n9899), .A2(n9920), .B1(n9898), .B2(n9925), .ZN(n9900)
         );
  NOR2_X1 U10942 ( .A1(n9901), .A2(n9900), .ZN(n9943) );
  AOI22_X1 U10943 ( .A1(n9939), .A2(n9902), .B1(n9943), .B2(n9937), .ZN(
        P2_U3402) );
  INV_X1 U10944 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9908) );
  NOR2_X1 U10945 ( .A1(n9903), .A2(n9925), .ZN(n9905) );
  AOI211_X1 U10946 ( .C1(n9907), .C2(n9906), .A(n9905), .B(n9904), .ZN(n9944)
         );
  AOI22_X1 U10947 ( .A1(n9939), .A2(n9908), .B1(n9944), .B2(n9937), .ZN(
        P2_U3405) );
  INV_X1 U10948 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9913) );
  NOR2_X1 U10949 ( .A1(n9909), .A2(n9925), .ZN(n9911) );
  AOI211_X1 U10950 ( .C1(n9912), .C2(n9933), .A(n9911), .B(n9910), .ZN(n9945)
         );
  AOI22_X1 U10951 ( .A1(n9939), .A2(n9913), .B1(n9945), .B2(n9937), .ZN(
        P2_U3408) );
  INV_X1 U10952 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U10953 ( .A1(n9914), .A2(n9925), .ZN(n9916) );
  AOI211_X1 U10954 ( .C1(n9933), .C2(n9917), .A(n9916), .B(n9915), .ZN(n9946)
         );
  AOI22_X1 U10955 ( .A1(n9939), .A2(n9918), .B1(n9946), .B2(n9937), .ZN(
        P2_U3414) );
  INV_X1 U10956 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9924) );
  OAI22_X1 U10957 ( .A1(n9921), .A2(n9920), .B1(n9919), .B2(n9925), .ZN(n9922)
         );
  NOR2_X1 U10958 ( .A1(n9923), .A2(n9922), .ZN(n9947) );
  AOI22_X1 U10959 ( .A1(n9939), .A2(n9924), .B1(n9947), .B2(n9937), .ZN(
        P2_U3420) );
  INV_X1 U10960 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9930) );
  NOR2_X1 U10961 ( .A1(n9926), .A2(n9925), .ZN(n9928) );
  AOI211_X1 U10962 ( .C1(n9933), .C2(n9929), .A(n9928), .B(n9927), .ZN(n9948)
         );
  AOI22_X1 U10963 ( .A1(n9939), .A2(n9930), .B1(n9948), .B2(n9937), .ZN(
        P2_U3423) );
  INV_X1 U10964 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9938) );
  AOI22_X1 U10965 ( .A1(n9934), .A2(n9933), .B1(n9932), .B2(n9931), .ZN(n9935)
         );
  AND2_X1 U10966 ( .A1(n9936), .A2(n9935), .ZN(n9949) );
  AOI22_X1 U10967 ( .A1(n9939), .A2(n9938), .B1(n9949), .B2(n9937), .ZN(
        P2_U3426) );
  AOI22_X1 U10968 ( .A1(n9950), .A2(n9940), .B1(n6727), .B2(n6277), .ZN(
        P2_U3460) );
  AOI22_X1 U10969 ( .A1(n9950), .A2(n9941), .B1(n6687), .B2(n6277), .ZN(
        P2_U3461) );
  AOI22_X1 U10970 ( .A1(n9950), .A2(n9943), .B1(n9942), .B2(n6277), .ZN(
        P2_U3463) );
  AOI22_X1 U10971 ( .A1(n9950), .A2(n9944), .B1(n5864), .B2(n6277), .ZN(
        P2_U3464) );
  AOI22_X1 U10972 ( .A1(n9950), .A2(n9945), .B1(n6815), .B2(n6277), .ZN(
        P2_U3465) );
  AOI22_X1 U10973 ( .A1(n9950), .A2(n9946), .B1(n7004), .B2(n6277), .ZN(
        P2_U3467) );
  AOI22_X1 U10974 ( .A1(n9950), .A2(n9947), .B1(n7193), .B2(n6277), .ZN(
        P2_U3469) );
  AOI22_X1 U10975 ( .A1(n9950), .A2(n9948), .B1(n7246), .B2(n6277), .ZN(
        P2_U3470) );
  AOI22_X1 U10976 ( .A1(n9950), .A2(n9949), .B1(n7441), .B2(n6277), .ZN(
        P2_U3471) );
  INV_X1 U10977 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9954) );
  NAND3_X1 U10978 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9953) );
  AND2_X1 U10979 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9951) );
  NOR2_X1 U10980 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9951), .ZN(n9952) );
  INV_X1 U10981 ( .A(n9952), .ZN(n9969) );
  NAND2_X1 U10982 ( .A1(n9954), .A2(n9953), .ZN(n9968) );
  OAI222_X1 U10983 ( .A1(n9954), .A2(n9953), .B1(n9954), .B2(n9969), .C1(n9952), .C2(n9968), .ZN(ADD_1068_U5) );
  XOR2_X1 U10984 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U10985 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9955) );
  AOI21_X1 U10986 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9955), .ZN(n9976) );
  NOR2_X1 U10987 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9956) );
  AOI21_X1 U10988 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9956), .ZN(n9979) );
  NOR2_X1 U10989 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9957) );
  AOI21_X1 U10990 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9957), .ZN(n9982) );
  NOR2_X1 U10991 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9958) );
  AOI21_X1 U10992 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9958), .ZN(n9985) );
  NOR2_X1 U10993 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9959) );
  AOI21_X1 U10994 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9959), .ZN(n9988) );
  NOR2_X1 U10995 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9960) );
  AOI21_X1 U10996 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9960), .ZN(n9991) );
  NOR2_X1 U10997 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9961) );
  AOI21_X1 U10998 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9961), .ZN(n9994) );
  NOR2_X1 U10999 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9962) );
  AOI21_X1 U11000 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9962), .ZN(n9997) );
  NOR2_X1 U11001 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9963) );
  AOI21_X1 U11002 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n9963), .ZN(n10199) );
  NOR2_X1 U11003 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9964) );
  AOI21_X1 U11004 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n9964), .ZN(n10202) );
  NOR2_X1 U11005 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9965) );
  AOI21_X1 U11006 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n9965), .ZN(n10205) );
  NOR2_X1 U11007 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9966) );
  AOI21_X1 U11008 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n9966), .ZN(n10208) );
  NOR2_X1 U11009 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n9967) );
  AOI21_X1 U11010 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n9967), .ZN(n10211) );
  NAND2_X1 U11011 ( .A1(n9969), .A2(n9968), .ZN(n10196) );
  NAND2_X1 U11012 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9970) );
  OAI21_X1 U11013 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n9970), .ZN(n10195) );
  NOR2_X1 U11014 ( .A1(n10196), .A2(n10195), .ZN(n10194) );
  AOI21_X1 U11015 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10194), .ZN(n10214) );
  NAND2_X1 U11016 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9971) );
  OAI21_X1 U11017 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n9971), .ZN(n10213) );
  NOR2_X1 U11018 ( .A1(n10214), .A2(n10213), .ZN(n10212) );
  AOI21_X1 U11019 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10212), .ZN(n10217) );
  NOR2_X1 U11020 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9972) );
  AOI21_X1 U11021 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n9972), .ZN(n10216) );
  NAND2_X1 U11022 ( .A1(n10217), .A2(n10216), .ZN(n10215) );
  OAI21_X1 U11023 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10215), .ZN(n10210) );
  NAND2_X1 U11024 ( .A1(n10211), .A2(n10210), .ZN(n10209) );
  OAI21_X1 U11025 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10209), .ZN(n10207) );
  NAND2_X1 U11026 ( .A1(n10208), .A2(n10207), .ZN(n10206) );
  OAI21_X1 U11027 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10206), .ZN(n10204) );
  NAND2_X1 U11028 ( .A1(n10205), .A2(n10204), .ZN(n10203) );
  OAI21_X1 U11029 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10203), .ZN(n10201) );
  NAND2_X1 U11030 ( .A1(n10202), .A2(n10201), .ZN(n10200) );
  OAI21_X1 U11031 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10200), .ZN(n10198) );
  NAND2_X1 U11032 ( .A1(n10199), .A2(n10198), .ZN(n10197) );
  OAI21_X1 U11033 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10197), .ZN(n9996) );
  NAND2_X1 U11034 ( .A1(n9997), .A2(n9996), .ZN(n9995) );
  OAI21_X1 U11035 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9995), .ZN(n9993) );
  NAND2_X1 U11036 ( .A1(n9994), .A2(n9993), .ZN(n9992) );
  OAI21_X1 U11037 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9992), .ZN(n9990) );
  NAND2_X1 U11038 ( .A1(n9991), .A2(n9990), .ZN(n9989) );
  OAI21_X1 U11039 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9989), .ZN(n9987) );
  NAND2_X1 U11040 ( .A1(n9988), .A2(n9987), .ZN(n9986) );
  OAI21_X1 U11041 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9986), .ZN(n9984) );
  NAND2_X1 U11042 ( .A1(n9985), .A2(n9984), .ZN(n9983) );
  OAI21_X1 U11043 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9983), .ZN(n9981) );
  NAND2_X1 U11044 ( .A1(n9982), .A2(n9981), .ZN(n9980) );
  OAI21_X1 U11045 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9980), .ZN(n9978) );
  NAND2_X1 U11046 ( .A1(n9979), .A2(n9978), .ZN(n9977) );
  OAI21_X1 U11047 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9977), .ZN(n9975) );
  NAND2_X1 U11048 ( .A1(n9976), .A2(n9975), .ZN(n9974) );
  OAI21_X1 U11049 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9974), .ZN(n10186) );
  NAND2_X1 U11050 ( .A1(n10187), .A2(n10186), .ZN(n10188) );
  OAI21_X1 U11051 ( .B1(n10186), .B2(n10187), .A(n10188), .ZN(n9973) );
  XNOR2_X1 U11052 ( .A(n9973), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11053 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(ADD_1068_U56) );
  OAI21_X1 U11054 ( .B1(n9979), .B2(n9978), .A(n9977), .ZN(ADD_1068_U57) );
  OAI21_X1 U11055 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(ADD_1068_U58) );
  OAI21_X1 U11056 ( .B1(n9985), .B2(n9984), .A(n9983), .ZN(ADD_1068_U59) );
  OAI21_X1 U11057 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(ADD_1068_U60) );
  OAI21_X1 U11058 ( .B1(n9991), .B2(n9990), .A(n9989), .ZN(ADD_1068_U61) );
  OAI21_X1 U11059 ( .B1(n9994), .B2(n9993), .A(n9992), .ZN(ADD_1068_U62) );
  OAI21_X1 U11060 ( .B1(n9997), .B2(n9996), .A(n9995), .ZN(ADD_1068_U63) );
  AOI22_X1 U11061 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n9998) );
  OAI221_X1 U11062 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n9998), .ZN(n10005) );
  AOI22_X1 U11063 ( .A1(SI_8_), .A2(keyinput_f24), .B1(SI_26_), .B2(
        keyinput_f6), .ZN(n9999) );
  OAI221_X1 U11064 ( .B1(SI_8_), .B2(keyinput_f24), .C1(SI_26_), .C2(
        keyinput_f6), .A(n9999), .ZN(n10004) );
  AOI22_X1 U11065 ( .A1(SI_13_), .A2(keyinput_f19), .B1(SI_23_), .B2(
        keyinput_f9), .ZN(n10000) );
  OAI221_X1 U11066 ( .B1(SI_13_), .B2(keyinput_f19), .C1(SI_23_), .C2(
        keyinput_f9), .A(n10000), .ZN(n10003) );
  AOI22_X1 U11067 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_f56), .B1(SI_4_), .B2(keyinput_f28), .ZN(n10001) );
  OAI221_X1 U11068 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .C1(
        SI_4_), .C2(keyinput_f28), .A(n10001), .ZN(n10002) );
  NOR4_X1 U11069 ( .A1(n10005), .A2(n10004), .A3(n10003), .A4(n10002), .ZN(
        n10033) );
  XNOR2_X1 U11070 ( .A(keyinput_f0), .B(P2_WR_REG_SCAN_IN), .ZN(n10012) );
  AOI22_X1 U11071 ( .A1(SI_15_), .A2(keyinput_f17), .B1(n10130), .B2(
        keyinput_f35), .ZN(n10006) );
  OAI221_X1 U11072 ( .B1(SI_15_), .B2(keyinput_f17), .C1(n10130), .C2(
        keyinput_f35), .A(n10006), .ZN(n10011) );
  AOI22_X1 U11073 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        SI_24_), .B2(keyinput_f8), .ZN(n10007) );
  OAI221_X1 U11074 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        SI_24_), .C2(keyinput_f8), .A(n10007), .ZN(n10010) );
  AOI22_X1 U11075 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(SI_5_), 
        .B2(keyinput_f27), .ZN(n10008) );
  OAI221_X1 U11076 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(SI_5_), .C2(keyinput_f27), .A(n10008), .ZN(n10009) );
  NOR4_X1 U11077 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10032) );
  AOI22_X1 U11078 ( .A1(SI_31_), .A2(keyinput_f1), .B1(SI_9_), .B2(
        keyinput_f23), .ZN(n10013) );
  OAI221_X1 U11079 ( .B1(SI_31_), .B2(keyinput_f1), .C1(SI_9_), .C2(
        keyinput_f23), .A(n10013), .ZN(n10021) );
  AOI22_X1 U11080 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n10014) );
  OAI221_X1 U11081 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n10014), .ZN(n10020)
         );
  AOI22_X1 U11082 ( .A1(SI_25_), .A2(keyinput_f7), .B1(n10016), .B2(
        keyinput_f37), .ZN(n10015) );
  OAI221_X1 U11083 ( .B1(SI_25_), .B2(keyinput_f7), .C1(n10016), .C2(
        keyinput_f37), .A(n10015), .ZN(n10019) );
  AOI22_X1 U11084 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(
        SI_16_), .B2(keyinput_f16), .ZN(n10017) );
  OAI221_X1 U11085 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        SI_16_), .C2(keyinput_f16), .A(n10017), .ZN(n10018) );
  NOR4_X1 U11086 ( .A1(n10021), .A2(n10020), .A3(n10019), .A4(n10018), .ZN(
        n10031) );
  AOI22_X1 U11087 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        SI_10_), .B2(keyinput_f22), .ZN(n10022) );
  OAI221_X1 U11088 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        SI_10_), .C2(keyinput_f22), .A(n10022), .ZN(n10029) );
  AOI22_X1 U11089 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        SI_14_), .B2(keyinput_f18), .ZN(n10023) );
  OAI221_X1 U11090 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        SI_14_), .C2(keyinput_f18), .A(n10023), .ZN(n10028) );
  AOI22_X1 U11091 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n10024) );
  OAI221_X1 U11092 ( .B1(SI_30_), .B2(keyinput_f2), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n10024), .ZN(n10027)
         );
  AOI22_X1 U11093 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_f33), .ZN(n10025) );
  OAI221_X1 U11094 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_f33), .A(n10025), .ZN(n10026) );
  NOR4_X1 U11095 ( .A1(n10029), .A2(n10028), .A3(n10027), .A4(n10026), .ZN(
        n10030) );
  NAND4_X1 U11096 ( .A1(n10033), .A2(n10032), .A3(n10031), .A4(n10030), .ZN(
        n10087) );
  INV_X1 U11097 ( .A(SI_12_), .ZN(n10036) );
  AOI22_X1 U11098 ( .A1(n10036), .A2(keyinput_f20), .B1(n10035), .B2(
        keyinput_f10), .ZN(n10034) );
  OAI221_X1 U11099 ( .B1(n10036), .B2(keyinput_f20), .C1(n10035), .C2(
        keyinput_f10), .A(n10034), .ZN(n10048) );
  AOI22_X1 U11100 ( .A1(n10129), .A2(keyinput_f3), .B1(n10038), .B2(
        keyinput_f55), .ZN(n10037) );
  OAI221_X1 U11101 ( .B1(n10129), .B2(keyinput_f3), .C1(n10038), .C2(
        keyinput_f55), .A(n10037), .ZN(n10047) );
  AOI22_X1 U11102 ( .A1(n10041), .A2(keyinput_f15), .B1(keyinput_f34), .B2(
        P2_U3151), .ZN(n10039) );
  OAI221_X1 U11103 ( .B1(n10041), .B2(keyinput_f15), .C1(P2_U3151), .C2(
        keyinput_f34), .A(n10039), .ZN(n10046) );
  INV_X1 U11104 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10043) );
  AOI22_X1 U11105 ( .A1(n10044), .A2(keyinput_f54), .B1(n10043), .B2(
        keyinput_f60), .ZN(n10042) );
  OAI221_X1 U11106 ( .B1(n10044), .B2(keyinput_f54), .C1(n10043), .C2(
        keyinput_f60), .A(n10042), .ZN(n10045) );
  NOR4_X1 U11107 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        n10085) );
  AOI22_X1 U11108 ( .A1(n5766), .A2(keyinput_f49), .B1(keyinput_f59), .B2(
        n6707), .ZN(n10049) );
  OAI221_X1 U11109 ( .B1(n5766), .B2(keyinput_f49), .C1(n6707), .C2(
        keyinput_f59), .A(n10049), .ZN(n10057) );
  INV_X1 U11110 ( .A(SI_18_), .ZN(n10171) );
  AOI22_X1 U11111 ( .A1(n10171), .A2(keyinput_f14), .B1(n10167), .B2(
        keyinput_f5), .ZN(n10050) );
  OAI221_X1 U11112 ( .B1(n10171), .B2(keyinput_f14), .C1(n10167), .C2(
        keyinput_f5), .A(n10050), .ZN(n10056) );
  AOI22_X1 U11113 ( .A1(n10128), .A2(keyinput_f39), .B1(n10170), .B2(
        keyinput_f12), .ZN(n10051) );
  OAI221_X1 U11114 ( .B1(n10128), .B2(keyinput_f39), .C1(n10170), .C2(
        keyinput_f12), .A(n10051), .ZN(n10055) );
  XOR2_X1 U11115 ( .A(n5769), .B(keyinput_f53), .Z(n10053) );
  XNOR2_X1 U11116 ( .A(SI_2_), .B(keyinput_f30), .ZN(n10052) );
  NAND2_X1 U11117 ( .A1(n10053), .A2(n10052), .ZN(n10054) );
  NOR4_X1 U11118 ( .A1(n10057), .A2(n10056), .A3(n10055), .A4(n10054), .ZN(
        n10084) );
  AOI22_X1 U11119 ( .A1(n10060), .A2(keyinput_f41), .B1(n10059), .B2(
        keyinput_f45), .ZN(n10058) );
  OAI221_X1 U11120 ( .B1(n10060), .B2(keyinput_f41), .C1(n10059), .C2(
        keyinput_f45), .A(n10058), .ZN(n10069) );
  AOI22_X1 U11121 ( .A1(n10141), .A2(keyinput_f52), .B1(n10062), .B2(
        keyinput_f50), .ZN(n10061) );
  OAI221_X1 U11122 ( .B1(n10141), .B2(keyinput_f52), .C1(n10062), .C2(
        keyinput_f50), .A(n10061), .ZN(n10068) );
  XNOR2_X1 U11123 ( .A(SI_7_), .B(keyinput_f25), .ZN(n10066) );
  XNOR2_X1 U11124 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10065) );
  XNOR2_X1 U11125 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_f48), .ZN(n10064)
         );
  XNOR2_X1 U11126 ( .A(SI_3_), .B(keyinput_f29), .ZN(n10063) );
  NAND4_X1 U11127 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        n10067) );
  NOR3_X1 U11128 ( .A1(n10069), .A2(n10068), .A3(n10067), .ZN(n10083) );
  AOI22_X1 U11129 ( .A1(n10071), .A2(keyinput_f4), .B1(keyinput_f43), .B2(
        n10157), .ZN(n10070) );
  OAI221_X1 U11130 ( .B1(n10071), .B2(keyinput_f4), .C1(n10157), .C2(
        keyinput_f43), .A(n10070), .ZN(n10081) );
  AOI22_X1 U11131 ( .A1(n10074), .A2(keyinput_f26), .B1(n10073), .B2(
        keyinput_f13), .ZN(n10072) );
  OAI221_X1 U11132 ( .B1(n10074), .B2(keyinput_f26), .C1(n10073), .C2(
        keyinput_f13), .A(n10072), .ZN(n10080) );
  AOI22_X1 U11133 ( .A1(n10126), .A2(keyinput_f58), .B1(n10076), .B2(
        keyinput_f47), .ZN(n10075) );
  OAI221_X1 U11134 ( .B1(n10126), .B2(keyinput_f58), .C1(n10076), .C2(
        keyinput_f47), .A(n10075), .ZN(n10079) );
  INV_X1 U11135 ( .A(SI_21_), .ZN(n10150) );
  INV_X1 U11136 ( .A(SI_0_), .ZN(n10154) );
  AOI22_X1 U11137 ( .A1(n10150), .A2(keyinput_f11), .B1(keyinput_f32), .B2(
        n10154), .ZN(n10077) );
  OAI221_X1 U11138 ( .B1(n10150), .B2(keyinput_f11), .C1(n10154), .C2(
        keyinput_f32), .A(n10077), .ZN(n10078) );
  NOR4_X1 U11139 ( .A1(n10081), .A2(n10080), .A3(n10079), .A4(n10078), .ZN(
        n10082) );
  NAND4_X1 U11140 ( .A1(n10085), .A2(n10084), .A3(n10083), .A4(n10082), .ZN(
        n10086) );
  OAI22_X1 U11141 ( .A1(n10087), .A2(n10086), .B1(keyinput_f21), .B2(SI_11_), 
        .ZN(n10088) );
  AOI21_X1 U11142 ( .B1(keyinput_f21), .B2(SI_11_), .A(n10088), .ZN(n10185) );
  AOI22_X1 U11143 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_g53), .B1(SI_28_), .B2(keyinput_g4), .ZN(n10089) );
  OAI221_X1 U11144 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .C1(
        SI_28_), .C2(keyinput_g4), .A(n10089), .ZN(n10096) );
  AOI22_X1 U11145 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        SI_19_), .B2(keyinput_g13), .ZN(n10090) );
  OAI221_X1 U11146 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        SI_19_), .C2(keyinput_g13), .A(n10090), .ZN(n10095) );
  AOI22_X1 U11147 ( .A1(SI_10_), .A2(keyinput_g22), .B1(SI_24_), .B2(
        keyinput_g8), .ZN(n10091) );
  OAI221_X1 U11148 ( .B1(SI_10_), .B2(keyinput_g22), .C1(SI_24_), .C2(
        keyinput_g8), .A(n10091), .ZN(n10094) );
  AOI22_X1 U11149 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(SI_6_), 
        .B2(keyinput_g26), .ZN(n10092) );
  OAI221_X1 U11150 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(SI_6_), .C2(keyinput_g26), .A(n10092), .ZN(n10093) );
  NOR4_X1 U11151 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(
        n10123) );
  XOR2_X1 U11152 ( .A(SI_5_), .B(keyinput_g27), .Z(n10103) );
  AOI22_X1 U11153 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_g38), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n10097) );
  OAI221_X1 U11154 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n10097), .ZN(n10102)
         );
  AOI22_X1 U11155 ( .A1(SI_30_), .A2(keyinput_g2), .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n10098) );
  OAI221_X1 U11156 ( .B1(SI_30_), .B2(keyinput_g2), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n10098), .ZN(n10101)
         );
  AOI22_X1 U11157 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_23_), .B2(keyinput_g9), .ZN(n10099) );
  OAI221_X1 U11158 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        SI_23_), .C2(keyinput_g9), .A(n10099), .ZN(n10100) );
  NOR4_X1 U11159 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10122) );
  AOI22_X1 U11160 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(SI_3_), .B2(keyinput_g29), .ZN(n10104) );
  OAI221_X1 U11161 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        SI_3_), .C2(keyinput_g29), .A(n10104), .ZN(n10111) );
  AOI22_X1 U11162 ( .A1(SI_1_), .A2(keyinput_g31), .B1(SI_17_), .B2(
        keyinput_g15), .ZN(n10105) );
  OAI221_X1 U11163 ( .B1(SI_1_), .B2(keyinput_g31), .C1(SI_17_), .C2(
        keyinput_g15), .A(n10105), .ZN(n10110) );
  AOI22_X1 U11164 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        SI_22_), .B2(keyinput_g10), .ZN(n10106) );
  OAI221_X1 U11165 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        SI_22_), .C2(keyinput_g10), .A(n10106), .ZN(n10109) );
  AOI22_X1 U11166 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        SI_13_), .B2(keyinput_g19), .ZN(n10107) );
  OAI221_X1 U11167 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        SI_13_), .C2(keyinput_g19), .A(n10107), .ZN(n10108) );
  NOR4_X1 U11168 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n10121) );
  AOI22_X1 U11169 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n10112) );
  OAI221_X1 U11170 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n10112), .ZN(n10119)
         );
  AOI22_X1 U11171 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n10113) );
  OAI221_X1 U11172 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n10113), .ZN(n10118)
         );
  AOI22_X1 U11173 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .ZN(n10114) );
  OAI221_X1 U11174 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n10114), .ZN(n10117) );
  AOI22_X1 U11175 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_g45), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n10115) );
  OAI221_X1 U11176 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n10115), .ZN(n10116) );
  NOR4_X1 U11177 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(n10116), .ZN(
        n10120) );
  NAND4_X1 U11178 ( .A1(n10123), .A2(n10122), .A3(n10121), .A4(n10120), .ZN(
        n10183) );
  AOI22_X1 U11179 ( .A1(n10126), .A2(keyinput_g58), .B1(n10125), .B2(
        keyinput_g56), .ZN(n10124) );
  OAI221_X1 U11180 ( .B1(n10126), .B2(keyinput_g58), .C1(n10125), .C2(
        keyinput_g56), .A(n10124), .ZN(n10137) );
  AOI22_X1 U11181 ( .A1(n10129), .A2(keyinput_g3), .B1(n10128), .B2(
        keyinput_g39), .ZN(n10127) );
  OAI221_X1 U11182 ( .B1(n10129), .B2(keyinput_g3), .C1(n10128), .C2(
        keyinput_g39), .A(n10127), .ZN(n10136) );
  XOR2_X1 U11183 ( .A(n10130), .B(keyinput_g35), .Z(n10134) );
  XNOR2_X1 U11184 ( .A(SI_2_), .B(keyinput_g30), .ZN(n10133) );
  XNOR2_X1 U11185 ( .A(SI_4_), .B(keyinput_g28), .ZN(n10132) );
  XNOR2_X1 U11186 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_g46), .ZN(n10131)
         );
  NAND4_X1 U11187 ( .A1(n10134), .A2(n10133), .A3(n10132), .A4(n10131), .ZN(
        n10135) );
  NOR3_X1 U11188 ( .A1(n10137), .A2(n10136), .A3(n10135), .ZN(n10181) );
  AOI22_X1 U11189 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(SI_25_), .B2(keyinput_g7), .ZN(n10138) );
  OAI221_X1 U11190 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        SI_25_), .C2(keyinput_g7), .A(n10138), .ZN(n10147) );
  AOI22_X1 U11191 ( .A1(SI_7_), .A2(keyinput_g25), .B1(SI_12_), .B2(
        keyinput_g20), .ZN(n10139) );
  OAI221_X1 U11192 ( .B1(SI_7_), .B2(keyinput_g25), .C1(SI_12_), .C2(
        keyinput_g20), .A(n10139), .ZN(n10146) );
  AOI22_X1 U11193 ( .A1(n7646), .A2(keyinput_g1), .B1(n10141), .B2(
        keyinput_g52), .ZN(n10140) );
  OAI221_X1 U11194 ( .B1(n7646), .B2(keyinput_g1), .C1(n10141), .C2(
        keyinput_g52), .A(n10140), .ZN(n10145) );
  AOI22_X1 U11195 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(
        n10143), .B2(keyinput_g24), .ZN(n10142) );
  OAI221_X1 U11196 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        n10143), .C2(keyinput_g24), .A(n10142), .ZN(n10144) );
  NOR4_X1 U11197 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n10180) );
  AOI22_X1 U11198 ( .A1(n10150), .A2(keyinput_g11), .B1(keyinput_g16), .B2(
        n10149), .ZN(n10148) );
  OAI221_X1 U11199 ( .B1(n10150), .B2(keyinput_g11), .C1(n10149), .C2(
        keyinput_g16), .A(n10148), .ZN(n10162) );
  INV_X1 U11200 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U11201 ( .A1(n5773), .A2(keyinput_g63), .B1(n10152), .B2(
        keyinput_g36), .ZN(n10151) );
  OAI221_X1 U11202 ( .B1(n5773), .B2(keyinput_g63), .C1(n10152), .C2(
        keyinput_g36), .A(n10151), .ZN(n10161) );
  AOI22_X1 U11203 ( .A1(n10155), .A2(keyinput_g17), .B1(keyinput_g32), .B2(
        n10154), .ZN(n10153) );
  OAI221_X1 U11204 ( .B1(n10155), .B2(keyinput_g17), .C1(n10154), .C2(
        keyinput_g32), .A(n10153), .ZN(n10160) );
  INV_X1 U11205 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10158) );
  AOI22_X1 U11206 ( .A1(n10158), .A2(keyinput_g0), .B1(n10157), .B2(
        keyinput_g43), .ZN(n10156) );
  OAI221_X1 U11207 ( .B1(n10158), .B2(keyinput_g0), .C1(n10157), .C2(
        keyinput_g43), .A(n10156), .ZN(n10159) );
  NOR4_X1 U11208 ( .A1(n10162), .A2(n10161), .A3(n10160), .A4(n10159), .ZN(
        n10179) );
  AOI22_X1 U11209 ( .A1(n10165), .A2(keyinput_g40), .B1(n10164), .B2(
        keyinput_g6), .ZN(n10163) );
  OAI221_X1 U11210 ( .B1(n10165), .B2(keyinput_g40), .C1(n10164), .C2(
        keyinput_g6), .A(n10163), .ZN(n10177) );
  AOI22_X1 U11211 ( .A1(n10168), .A2(keyinput_g18), .B1(n10167), .B2(
        keyinput_g5), .ZN(n10166) );
  OAI221_X1 U11212 ( .B1(n10168), .B2(keyinput_g18), .C1(n10167), .C2(
        keyinput_g5), .A(n10166), .ZN(n10176) );
  AOI22_X1 U11213 ( .A1(n10171), .A2(keyinput_g14), .B1(n10170), .B2(
        keyinput_g12), .ZN(n10169) );
  OAI221_X1 U11214 ( .B1(n10171), .B2(keyinput_g14), .C1(n10170), .C2(
        keyinput_g12), .A(n10169), .ZN(n10175) );
  AOI22_X1 U11215 ( .A1(n10173), .A2(keyinput_g23), .B1(keyinput_g44), .B2(
        n6974), .ZN(n10172) );
  OAI221_X1 U11216 ( .B1(n10173), .B2(keyinput_g23), .C1(n6974), .C2(
        keyinput_g44), .A(n10172), .ZN(n10174) );
  NOR4_X1 U11217 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n10178) );
  NAND4_X1 U11218 ( .A1(n10181), .A2(n10180), .A3(n10179), .A4(n10178), .ZN(
        n10182) );
  OAI22_X1 U11219 ( .A1(SI_11_), .A2(keyinput_g21), .B1(n10183), .B2(n10182), 
        .ZN(n10184) );
  AOI211_X1 U11220 ( .C1(SI_11_), .C2(keyinput_g21), .A(n10185), .B(n10184), 
        .ZN(n10193) );
  NOR2_X1 U11221 ( .A1(n10187), .A2(n10186), .ZN(n10189) );
  OAI21_X1 U11222 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10189), .A(n10188), 
        .ZN(n10191) );
  XNOR2_X1 U11223 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10190) );
  XNOR2_X1 U11224 ( .A(n10191), .B(n10190), .ZN(n10192) );
  XNOR2_X1 U11225 ( .A(n10193), .B(n10192), .ZN(ADD_1068_U4) );
  AOI21_X1 U11226 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(ADD_1068_U54) );
  OAI21_X1 U11227 ( .B1(n10199), .B2(n10198), .A(n10197), .ZN(ADD_1068_U47) );
  OAI21_X1 U11228 ( .B1(n10202), .B2(n10201), .A(n10200), .ZN(ADD_1068_U48) );
  OAI21_X1 U11229 ( .B1(n10205), .B2(n10204), .A(n10203), .ZN(ADD_1068_U49) );
  OAI21_X1 U11230 ( .B1(n10208), .B2(n10207), .A(n10206), .ZN(ADD_1068_U50) );
  OAI21_X1 U11231 ( .B1(n10211), .B2(n10210), .A(n10209), .ZN(ADD_1068_U51) );
  AOI21_X1 U11232 ( .B1(n10214), .B2(n10213), .A(n10212), .ZN(ADD_1068_U53) );
  OAI21_X1 U11233 ( .B1(n10217), .B2(n10216), .A(n10215), .ZN(ADD_1068_U52) );
  NAND2_X1 U5014 ( .A1(n8448), .A2(n7015), .ZN(n8412) );
  CLKBUF_X3 U4976 ( .A(n5032), .Z(n5656) );
  NAND2_X1 U4862 ( .A1(n5015), .A2(n5032), .ZN(n5045) );
  CLKBUF_X2 U4885 ( .A(n5035), .Z(n7655) );
  CLKBUF_X1 U4893 ( .A(n6708), .Z(n4354) );
  CLKBUF_X1 U4930 ( .A(n5726), .Z(n4352) );
endmodule

