

module b17_C_SARLock_k_64_4 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, U355, U356, U357, U358, 
        U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, 
        U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, 
        U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, 
        U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, 
        U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, 
        U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, 
        U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, 
        U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9588, n9589, n9590, n9591, n9592, n9593, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232;

  INV_X1 U11033 ( .A(n18427), .ZN(n18436) );
  OR2_X1 U11034 ( .A1(n14623), .A2(n14557), .ZN(n14563) );
  OR2_X2 U11035 ( .A1(n16911), .A2(n9824), .ZN(n15567) );
  INV_X1 U11036 ( .A(n10350), .ZN(n10362) );
  NOR2_X1 U11037 ( .A1(n10537), .A2(n10536), .ZN(n10597) );
  NOR2_X1 U11038 ( .A1(n10537), .A2(n16217), .ZN(n10545) );
  OR2_X1 U11039 ( .A1(n10522), .A2(n10538), .ZN(n10609) );
  OAI21_X1 U11040 ( .B1(n14445), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10145), 
        .ZN(n11254) );
  INV_X1 U11041 ( .A(n12740), .ZN(n14461) );
  NAND2_X1 U11042 ( .A1(n11207), .A2(n11208), .ZN(n13653) );
  CLKBUF_X2 U11043 ( .A(n10443), .Z(n10773) );
  AND2_X1 U11045 ( .A1(n10418), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12384) );
  AND2_X2 U11046 ( .A1(n12601), .A2(n10416), .ZN(n10277) );
  AND2_X1 U11047 ( .A1(n10421), .A2(n10416), .ZN(n12202) );
  INV_X2 U11048 ( .A(n12315), .ZN(n12423) );
  AND3_X1 U11049 ( .A1(n11205), .A2(n11130), .A3(n11129), .ZN(n9832) );
  NAND2_X1 U11050 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10226), .ZN(
        n12431) );
  NAND2_X1 U11051 ( .A1(n13173), .A2(n13071), .ZN(n11135) );
  INV_X1 U11052 ( .A(n14332), .ZN(n17821) );
  AND2_X1 U11053 ( .A1(n9669), .A2(n10098), .ZN(n11132) );
  BUF_X2 U11054 ( .A(n14190), .Z(n9595) );
  NAND2_X1 U11055 ( .A1(n14970), .A2(n11116), .ZN(n13126) );
  AND4_X1 U11056 ( .A1(n11093), .A2(n11092), .A3(n11091), .A4(n11090), .ZN(
        n11098) );
  AND2_X1 U11057 ( .A1(n11050), .A2(n13297), .ZN(n13110) );
  BUF_X1 U11058 ( .A(n10459), .Z(n13721) );
  AND2_X1 U11059 ( .A1(n9665), .A2(n11065), .ZN(n11128) );
  AND4_X1 U11060 ( .A1(n10978), .A2(n10977), .A3(n10976), .A4(n10975), .ZN(
        n10987) );
  NAND3_X1 U11061 ( .A1(n10024), .A2(n10023), .A3(n10020), .ZN(n19946) );
  BUF_X1 U11062 ( .A(n10406), .Z(n19962) );
  AND2_X1 U11063 ( .A1(n10979), .A2(n13156), .ZN(n11073) );
  AND2_X1 U11064 ( .A1(n13170), .A2(n13158), .ZN(n11074) );
  AND2_X1 U11065 ( .A1(n13139), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11153) );
  AND3_X2 U11066 ( .A1(n14499), .A2(n10201), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9589) );
  AND2_X2 U11067 ( .A1(n14486), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9600) );
  INV_X1 U11068 ( .A(n11154), .ZN(n11864) );
  CLKBUF_X2 U11069 ( .A(n11160), .Z(n9618) );
  NAND2_X1 U11070 ( .A1(n11128), .A2(n13288), .ZN(n12965) );
  NAND2_X1 U11071 ( .A1(n12880), .A2(n12514), .ZN(n14422) );
  AND2_X1 U11072 ( .A1(n10226), .A2(n17035), .ZN(n12429) );
  AND2_X2 U11073 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14486) );
  INV_X1 U11074 ( .A(n11153), .ZN(n11154) );
  OAI21_X1 U11075 ( .B1(n11135), .B2(n11206), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11209) );
  INV_X1 U11076 ( .A(n13721), .ZN(n10172) );
  INV_X2 U11077 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10201) );
  AND2_X1 U11078 ( .A1(n13066), .A2(n14501), .ZN(n12024) );
  NAND2_X1 U11079 ( .A1(n12047), .A2(n12046), .ZN(n12138) );
  OR2_X1 U11080 ( .A1(n13137), .A2(n11204), .ZN(n14976) );
  AND2_X1 U11081 ( .A1(n12606), .A2(n10416), .ZN(n12366) );
  AND2_X1 U11082 ( .A1(n9600), .A2(n10416), .ZN(n12433) );
  AND2_X1 U11083 ( .A1(n12606), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12365) );
  INV_X2 U11084 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10416) );
  CLKBUF_X2 U11085 ( .A(n12010), .Z(n9612) );
  NOR2_X1 U11086 ( .A1(n14865), .A2(n14826), .ZN(n14849) );
  OR2_X1 U11087 ( .A1(n20697), .A2(n9971), .ZN(n16831) );
  NAND2_X1 U11088 ( .A1(n12643), .A2(n12642), .ZN(n12719) );
  AND2_X1 U11089 ( .A1(n13009), .A2(n13008), .ZN(n13011) );
  INV_X1 U11090 ( .A(n17047), .ZN(n12642) );
  AOI21_X1 U11091 ( .B1(n9772), .B2(n9771), .A(n9678), .ZN(n9770) );
  NAND2_X1 U11092 ( .A1(n10822), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14017) );
  CLKBUF_X2 U11093 ( .A(n15305), .Z(n19753) );
  AND2_X1 U11094 ( .A1(n14713), .A2(n14702), .ZN(n14704) );
  NAND2_X1 U11095 ( .A1(n16179), .A2(n9659), .ZN(n16989) );
  NAND2_X1 U11096 ( .A1(n10844), .A2(n9715), .ZN(n15697) );
  NOR2_X1 U11098 ( .A1(n18141), .A2(n16290), .ZN(n17273) );
  INV_X1 U11099 ( .A(n18923), .ZN(n18102) );
  NOR2_X1 U11100 ( .A1(n18482), .A2(n18693), .ZN(n18388) );
  INV_X1 U11101 ( .A(n18587), .ZN(n18573) );
  INV_X2 U11102 ( .A(n19360), .ZN(n18753) );
  INV_X1 U11103 ( .A(n13860), .ZN(n13858) );
  INV_X1 U11104 ( .A(n20687), .ZN(n20703) );
  INV_X1 U11105 ( .A(n20676), .ZN(n16601) );
  XNOR2_X1 U11106 ( .A(n14372), .B(n12039), .ZN(n14815) );
  AOI211_X1 U11107 ( .C1(n16954), .C2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15859), .B(n15858), .ZN(n15860) );
  INV_X2 U11108 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14499) );
  INV_X1 U11109 ( .A(n18580), .ZN(n18571) );
  OR2_X1 U11111 ( .A1(n16041), .A2(n15407), .ZN(n15628) );
  AND2_X1 U11112 ( .A1(n10979), .A2(n13158), .ZN(n9607) );
  NAND2_X1 U11113 ( .A1(n12047), .A2(n12046), .ZN(n9588) );
  INV_X2 U11114 ( .A(n12138), .ZN(n15123) );
  INV_X1 U11115 ( .A(n11101), .ZN(n9619) );
  NOR2_X1 U11116 ( .A1(n14167), .A2(n17648), .ZN(n16386) );
  NAND2_X2 U11117 ( .A1(n16200), .A2(n10829), .ZN(n15914) );
  NOR4_X2 U11118 ( .A1(n18026), .A2(n18155), .A3(n18153), .A4(n17949), .ZN(
        n17991) );
  NOR2_X2 U11119 ( .A1(n15332), .A2(n15690), .ZN(n15335) );
  AND2_X4 U11120 ( .A1(n16212), .A2(n14499), .ZN(n10422) );
  NOR2_X4 U11121 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16212) );
  NOR3_X2 U11122 ( .A1(n18264), .A2(n18276), .A3(n18632), .ZN(n16412) );
  NOR3_X4 U11123 ( .A1(n18923), .A2(n16557), .A3(n17091), .ZN(n17938) );
  NOR2_X2 U11124 ( .A1(n14179), .A2(n14178), .ZN(n18923) );
  NAND2_X2 U11125 ( .A1(n10528), .A2(n10199), .ZN(n10610) );
  OAI22_X2 U11126 ( .A1(n15914), .A2(n10018), .B1(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n10017), .ZN(n15898) );
  AND2_X2 U11127 ( .A1(n14486), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9590) );
  AND2_X1 U11128 ( .A1(n14486), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10419) );
  NOR2_X1 U11129 ( .A1(n14836), .A2(n15009), .ZN(n14838) );
  NAND2_X1 U11130 ( .A1(n15767), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15725) );
  NOR2_X1 U11131 ( .A1(n20108), .A2(n20576), .ZN(n20042) );
  NOR2_X1 U11132 ( .A1(n20108), .A2(n20360), .ZN(n20102) );
  NAND2_X1 U11133 ( .A1(n11378), .A2(n11377), .ZN(n12047) );
  NAND2_X1 U11134 ( .A1(n18362), .A2(n18404), .ZN(n18324) );
  NAND2_X1 U11135 ( .A1(n13035), .A2(n11262), .ZN(n13065) );
  NAND2_X1 U11136 ( .A1(n10547), .A2(n10548), .ZN(n10594) );
  NOR2_X2 U11137 ( .A1(n19534), .A2(n18582), .ZN(n18427) );
  NAND2_X1 U11138 ( .A1(n12145), .A2(n14959), .ZN(n21068) );
  OR2_X1 U11139 ( .A1(n16406), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18459) );
  NAND2_X1 U11140 ( .A1(n9822), .A2(n10496), .ZN(n10499) );
  NOR2_X2 U11141 ( .A1(n18879), .A2(n19380), .ZN(n18888) );
  INV_X4 U11142 ( .A(n17655), .ZN(n17619) );
  NOR2_X1 U11143 ( .A1(n18213), .A2(n18209), .ZN(n17133) );
  BUF_X2 U11144 ( .A(n12776), .Z(n9591) );
  INV_X2 U11145 ( .A(n11143), .ZN(n14501) );
  NAND2_X1 U11146 ( .A1(n18087), .A2(n16274), .ZN(n16434) );
  INV_X2 U11147 ( .A(n18954), .ZN(n18087) );
  NAND3_X1 U11148 ( .A1(n14265), .A2(n14264), .A3(n14263), .ZN(n19574) );
  BUF_X1 U11149 ( .A(n11027), .Z(n9614) );
  CLKBUF_X2 U11150 ( .A(n9603), .Z(n11837) );
  INV_X1 U11151 ( .A(n17708), .ZN(n17901) );
  CLKBUF_X1 U11152 ( .A(n11037), .Z(n9592) );
  CLKBUF_X2 U11153 ( .A(n11074), .Z(n11870) );
  AND3_X2 U11155 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13139) );
  INV_X2 U11156 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13141) );
  INV_X1 U11157 ( .A(n9750), .ZN(n14818) );
  AND2_X1 U11158 ( .A1(n9777), .A2(n9776), .ZN(n14407) );
  NAND2_X1 U11159 ( .A1(n9886), .A2(n15799), .ZN(n15789) );
  NOR2_X2 U11160 ( .A1(n15697), .A2(n15970), .ZN(n15682) );
  OR2_X1 U11161 ( .A1(n15800), .A2(n15748), .ZN(n9886) );
  NAND2_X1 U11162 ( .A1(n10133), .A2(n10132), .ZN(n9750) );
  NAND2_X1 U11163 ( .A1(n10781), .A2(n9778), .ZN(n9777) );
  OR2_X1 U11164 ( .A1(n10057), .A2(n10054), .ZN(n10781) );
  OAI21_X1 U11165 ( .B1(n10053), .B2(n10057), .A(n15674), .ZN(n15676) );
  XNOR2_X1 U11166 ( .A(n12616), .B(n12615), .ZN(n12774) );
  NAND2_X1 U11167 ( .A1(n9782), .A2(n9781), .ZN(n10059) );
  OR2_X1 U11168 ( .A1(n16753), .A2(n16752), .ZN(n21059) );
  NAND2_X1 U11169 ( .A1(n10069), .A2(n10068), .ZN(n10761) );
  NAND2_X1 U11170 ( .A1(n10837), .A2(n10836), .ZN(n15896) );
  NAND2_X1 U11171 ( .A1(n9870), .A2(n9871), .ZN(n9869) );
  NAND2_X1 U11172 ( .A1(n9765), .A2(n9763), .ZN(n15873) );
  OR2_X1 U11173 ( .A1(n14151), .A2(n9684), .ZN(n9870) );
  OR2_X1 U11174 ( .A1(n10142), .A2(n10141), .ZN(n9871) );
  NOR2_X1 U11175 ( .A1(n9730), .A2(n9729), .ZN(n9728) );
  AND2_X1 U11176 ( .A1(n12131), .A2(n10143), .ZN(n10142) );
  XNOR2_X1 U11177 ( .A(n9982), .B(n14502), .ZN(n15025) );
  AOI21_X1 U11178 ( .B1(n10962), .B2(n16946), .A(n10961), .ZN(n10963) );
  OR2_X1 U11179 ( .A1(n14150), .A2(n10144), .ZN(n10143) );
  NAND2_X1 U11180 ( .A1(n9751), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18228) );
  INV_X1 U11181 ( .A(n12035), .ZN(n9982) );
  XNOR2_X1 U11182 ( .A(n10076), .B(n14427), .ZN(n16899) );
  AND3_X1 U11183 ( .A1(n9808), .A2(n9809), .A3(n9702), .ZN(n12493) );
  OR2_X1 U11184 ( .A1(n15120), .A2(n12125), .ZN(n16653) );
  OR2_X1 U11185 ( .A1(n16656), .A2(n12133), .ZN(n15121) );
  AOI21_X1 U11186 ( .B1(n16690), .B2(n10127), .A(n9676), .ZN(n10126) );
  OR2_X1 U11187 ( .A1(n15638), .A2(n9811), .ZN(n9809) );
  NOR2_X1 U11188 ( .A1(n14421), .A2(n14420), .ZN(n10076) );
  XNOR2_X1 U11189 ( .A(n12104), .B(n16808), .ZN(n16690) );
  NAND2_X1 U11190 ( .A1(n12103), .A2(n12102), .ZN(n12104) );
  XNOR2_X1 U11191 ( .A(n10810), .B(n12676), .ZN(n13993) );
  XNOR2_X1 U11192 ( .A(n12047), .B(n11380), .ZN(n12106) );
  NOR2_X1 U11193 ( .A1(n16619), .A2(n14397), .ZN(n16593) );
  NOR2_X1 U11194 ( .A1(n11373), .A2(n11349), .ZN(n11366) );
  OR2_X2 U11195 ( .A1(n15578), .A2(n15450), .ZN(n15571) );
  INV_X1 U11196 ( .A(n15628), .ZN(n10161) );
  NAND2_X1 U11197 ( .A1(n9827), .A2(n11325), .ZN(n11373) );
  INV_X1 U11198 ( .A(n11326), .ZN(n9827) );
  NOR2_X1 U11199 ( .A1(n10620), .A2(n10619), .ZN(n10623) );
  AND2_X1 U11200 ( .A1(n10672), .A2(n10671), .ZN(n10823) );
  AND2_X1 U11201 ( .A1(n13065), .A2(n11270), .ZN(n9724) );
  AND4_X1 U11202 ( .A1(n10587), .A2(n10586), .A3(n10585), .A4(n10584), .ZN(
        n10589) );
  OR3_X2 U11203 ( .A1(n16645), .A2(n13079), .A3(n13078), .ZN(n14805) );
  AOI22_X1 U11204 ( .A1(n20083), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n20138), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U11205 ( .A1(n11269), .A2(n11268), .ZN(n13064) );
  NAND2_X1 U11206 ( .A1(n10547), .A2(n10199), .ZN(n10593) );
  NAND2_X1 U11207 ( .A1(n10528), .A2(n10527), .ZN(n10596) );
  INV_X1 U11208 ( .A(n10650), .ZN(n10613) );
  INV_X1 U11209 ( .A(n15480), .ZN(n10152) );
  NAND2_X1 U11210 ( .A1(n10547), .A2(n10550), .ZN(n20023) );
  OR2_X2 U11211 ( .A1(n21061), .A2(n13097), .ZN(n16695) );
  OR2_X1 U11212 ( .A1(n13531), .A2(n11290), .ZN(n11269) );
  AND2_X2 U11213 ( .A1(n10526), .A2(n13062), .ZN(n10547) );
  NAND2_X1 U11214 ( .A1(n18587), .A2(n18489), .ZN(n18582) );
  NAND2_X1 U11215 ( .A1(n10545), .A2(n14113), .ZN(n20111) );
  NAND2_X1 U11216 ( .A1(n9759), .A2(n16473), .ZN(n18374) );
  AND2_X1 U11217 ( .A1(n11263), .A2(n12050), .ZN(n11244) );
  XNOR2_X1 U11218 ( .A(n11263), .B(n12050), .ZN(n13531) );
  NAND2_X1 U11219 ( .A1(n13199), .A2(n12992), .ZN(n21049) );
  NAND2_X1 U11220 ( .A1(n16406), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18403) );
  OR2_X1 U11221 ( .A1(n11254), .A2(n11201), .ZN(n11263) );
  AND2_X1 U11222 ( .A1(n11261), .A2(n11260), .ZN(n13034) );
  NAND2_X1 U11223 ( .A1(n18501), .A2(n16405), .ZN(n16406) );
  NAND2_X1 U11224 ( .A1(n12161), .A2(n17014), .ZN(n10537) );
  AOI21_X1 U11225 ( .B1(n12161), .B2(n12172), .A(n12164), .ZN(n12165) );
  NAND2_X1 U11226 ( .A1(n10514), .A2(n10513), .ZN(n10518) );
  NOR2_X2 U11227 ( .A1(n19937), .A2(n20395), .ZN(n19938) );
  NOR2_X2 U11228 ( .A1(n19868), .A2(n20395), .ZN(n13863) );
  NAND2_X1 U11229 ( .A1(n9814), .A2(n10499), .ZN(n17014) );
  INV_X1 U11230 ( .A(n10533), .ZN(n16217) );
  AOI21_X1 U11231 ( .B1(n10533), .B2(n12172), .A(n12155), .ZN(n13055) );
  AND2_X1 U11232 ( .A1(n9820), .A2(n9817), .ZN(n14090) );
  AND2_X1 U11233 ( .A1(n10850), .A2(n10512), .ZN(n10493) );
  NAND2_X1 U11234 ( .A1(n18537), .A2(n16401), .ZN(n18530) );
  NAND2_X1 U11235 ( .A1(n10509), .A2(n10852), .ZN(n10515) );
  NAND2_X1 U11236 ( .A1(n10470), .A2(n10469), .ZN(n10496) );
  NAND3_X1 U11237 ( .A1(n10481), .A2(n10480), .A3(n10482), .ZN(n9822) );
  NAND2_X1 U11238 ( .A1(n13282), .A2(n13281), .ZN(n20697) );
  OR2_X1 U11239 ( .A1(n10508), .A2(n10507), .ZN(n10509) );
  CLKBUF_X1 U11240 ( .A(n9605), .Z(n12778) );
  AOI21_X1 U11241 ( .B1(n9605), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10488), .ZN(n10490) );
  INV_X2 U11242 ( .A(n17942), .ZN(n17935) );
  AND2_X1 U11243 ( .A1(n10477), .A2(n10476), .ZN(n10481) );
  CLKBUF_X1 U11244 ( .A(n10500), .Z(n14426) );
  NAND2_X1 U11245 ( .A1(n10439), .A2(n10473), .ZN(n10506) );
  NAND2_X1 U11246 ( .A1(n18553), .A2(n16398), .ZN(n16400) );
  AOI21_X1 U11247 ( .B1(n17033), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10447), 
        .ZN(n10448) );
  AND2_X2 U11248 ( .A1(n10083), .A2(n10082), .ZN(n10500) );
  NAND2_X1 U11249 ( .A1(n10450), .A2(n10084), .ZN(n10083) );
  AND3_X1 U11250 ( .A1(n13136), .A2(n13578), .A3(n13128), .ZN(n11121) );
  INV_X1 U11251 ( .A(n9609), .ZN(n10882) );
  NAND2_X1 U11252 ( .A1(n18564), .A2(n16394), .ZN(n16397) );
  NAND2_X1 U11253 ( .A1(n12630), .A2(n10446), .ZN(n10450) );
  OR2_X1 U11254 ( .A1(n12771), .A2(n10950), .ZN(n10473) );
  NOR2_X2 U11255 ( .A1(n15307), .A2(n19655), .ZN(n15310) );
  NOR2_X1 U11256 ( .A1(n18076), .A2(n16380), .ZN(n16379) );
  AND2_X1 U11257 ( .A1(n10403), .A2(n12622), .ZN(n13732) );
  NAND2_X1 U11258 ( .A1(n10175), .A2(n9623), .ZN(n13731) );
  OR3_X1 U11259 ( .A1(n16434), .A2(n16271), .A3(n19369), .ZN(n16433) );
  OR2_X1 U11260 ( .A1(n12798), .A2(n15843), .ZN(n15307) );
  NAND2_X1 U11261 ( .A1(n14501), .A2(n11959), .ZN(n14503) );
  OAI21_X1 U11262 ( .B1(n12719), .B2(n12644), .A(n12647), .ZN(n13009) );
  OAI21_X1 U11263 ( .B1(n10475), .B2(n12651), .A(n12650), .ZN(n13008) );
  CLKBUF_X1 U11264 ( .A(n12651), .Z(n14464) );
  NAND2_X1 U11265 ( .A1(n11128), .A2(n11948), .ZN(n13155) );
  INV_X1 U11266 ( .A(n13738), .ZN(n10465) );
  INV_X1 U11267 ( .A(n11128), .ZN(n13309) );
  AND2_X1 U11268 ( .A1(n11124), .A2(n11204), .ZN(n11123) );
  AND2_X1 U11269 ( .A1(n11226), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11909) );
  INV_X1 U11270 ( .A(n16416), .ZN(n18930) );
  AND3_X1 U11271 ( .A1(n19962), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n17047), 
        .ZN(n12514) );
  INV_X1 U11272 ( .A(n11133), .ZN(n14978) );
  OR2_X2 U11273 ( .A1(n11080), .A2(n11079), .ZN(n13288) );
  INV_X1 U11274 ( .A(n14977), .ZN(n14970) );
  NAND2_X1 U11275 ( .A1(n10445), .A2(n10444), .ZN(n13738) );
  XNOR2_X1 U11276 ( .A(n16455), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18578) );
  INV_X2 U11277 ( .A(U212), .ZN(n17220) );
  NAND4_X2 U11278 ( .A1(n11026), .A2(n11025), .A3(n11024), .A4(n11023), .ZN(
        n14977) );
  NOR2_X1 U11279 ( .A1(n11004), .A2(n11003), .ZN(n11027) );
  NAND3_X1 U11280 ( .A1(n16343), .A2(n16342), .A3(n16341), .ZN(n16455) );
  NAND2_X1 U11281 ( .A1(n10243), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10250) );
  OR2_X2 U11282 ( .A1(n17221), .A2(n17168), .ZN(n17223) );
  AND4_X1 U11283 ( .A1(n10973), .A2(n10972), .A3(n10971), .A4(n10970), .ZN(
        n10988) );
  AND4_X1 U11284 ( .A1(n10985), .A2(n10984), .A3(n10983), .A4(n10982), .ZN(
        n10986) );
  AND4_X1 U11285 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(
        n11099) );
  AND4_X1 U11286 ( .A1(n11084), .A2(n11083), .A3(n11082), .A4(n11081), .ZN(
        n11100) );
  AND4_X1 U11287 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(
        n10999) );
  AND2_X1 U11288 ( .A1(n10022), .A2(n10021), .ZN(n10020) );
  NAND2_X2 U11289 ( .A1(n10428), .A2(n10427), .ZN(n10444) );
  AND4_X1 U11290 ( .A1(n11036), .A2(n11035), .A3(n11034), .A4(n11033), .ZN(
        n11048) );
  AND4_X1 U11291 ( .A1(n11032), .A2(n11031), .A3(n11030), .A4(n11029), .ZN(
        n11049) );
  AND4_X1 U11292 ( .A1(n11105), .A2(n11104), .A3(n11103), .A4(n11102), .ZN(
        n11115) );
  AND2_X1 U11293 ( .A1(n10214), .A2(n10213), .ZN(n10377) );
  INV_X2 U11294 ( .A(n12272), .ZN(n12421) );
  NAND2_X2 U11295 ( .A1(n19584), .A2(n19450), .ZN(n19513) );
  NAND2_X1 U11296 ( .A1(n10417), .A2(n10416), .ZN(n10428) );
  AND4_X1 U11297 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(
        n11026) );
  AND4_X1 U11298 ( .A1(n11014), .A2(n11013), .A3(n11012), .A4(n11011), .ZN(
        n11025) );
  AND3_X1 U11299 ( .A1(n10078), .A2(n10077), .A3(n10416), .ZN(n10206) );
  AND4_X1 U11300 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n10417) );
  AND2_X1 U11301 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  INV_X1 U11302 ( .A(n10198), .ZN(n17816) );
  NAND2_X2 U11303 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20627), .ZN(n20556) );
  AND2_X1 U11304 ( .A1(n10026), .A2(n10025), .ZN(n10040) );
  AND3_X1 U11305 ( .A1(n10208), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10207), .ZN(n10212) );
  AND2_X1 U11306 ( .A1(n10043), .A2(n10042), .ZN(n10041) );
  BUF_X2 U11307 ( .A(n16346), .Z(n17903) );
  AND3_X1 U11308 ( .A1(n10364), .A2(n10416), .A3(n10363), .ZN(n10367) );
  AND3_X1 U11309 ( .A1(n9761), .A2(n9760), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10426) );
  AND2_X1 U11310 ( .A1(n10028), .A2(n10027), .ZN(n10032) );
  AND3_X1 U11312 ( .A1(n10370), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10369), .ZN(n10374) );
  NAND2_X2 U11313 ( .A1(n20627), .A2(n20517), .ZN(n20559) );
  BUF_X2 U11314 ( .A(n11056), .Z(n9603) );
  INV_X1 U11315 ( .A(n9617), .ZN(n9593) );
  AND2_X2 U11317 ( .A1(n10422), .A2(n10416), .ZN(n10262) );
  INV_X2 U11318 ( .A(n19585), .ZN(n19584) );
  NOR2_X4 U11319 ( .A1(n14172), .A2(n14169), .ZN(n16346) );
  INV_X2 U11320 ( .A(n11816), .ZN(n11227) );
  BUF_X2 U11321 ( .A(n10420), .Z(n12601) );
  OR2_X1 U11322 ( .A1(n17648), .A2(n14166), .ZN(n14343) );
  NOR2_X1 U11323 ( .A1(n19534), .A2(n19432), .ZN(n18129) );
  INV_X2 U11324 ( .A(n17262), .ZN(n17264) );
  AND2_X4 U11325 ( .A1(n10979), .A2(n10980), .ZN(n11175) );
  AND2_X2 U11326 ( .A1(n10974), .A2(n10979), .ZN(n11192) );
  AND2_X2 U11327 ( .A1(n9611), .A2(n10416), .ZN(n12424) );
  INV_X1 U11328 ( .A(n9613), .ZN(n9596) );
  INV_X1 U11329 ( .A(n11787), .ZN(n9597) );
  NAND2_X1 U11330 ( .A1(n19531), .A2(n19541), .ZN(n14172) );
  NAND2_X1 U11331 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19548), .ZN(
        n14169) );
  NAND2_X1 U11332 ( .A1(n19548), .A2(n19554), .ZN(n17648) );
  AND2_X2 U11333 ( .A1(n10099), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10979) );
  AND4_X2 U11334 ( .A1(n14449), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9654) );
  INV_X2 U11335 ( .A(n21048), .ZN(n9598) );
  AND2_X1 U11336 ( .A1(n13152), .A2(n11005), .ZN(n11353) );
  AND2_X1 U11337 ( .A1(n13141), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10974) );
  INV_X2 U11338 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n21204) );
  AND2_X1 U11339 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14482) );
  AND2_X1 U11340 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13152) );
  NOR2_X1 U11341 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11005) );
  AND2_X1 U11342 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13158) );
  INV_X1 U11343 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19541) );
  INV_X1 U11344 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19548) );
  NAND2_X2 U11345 ( .A1(n11051), .A2(n13110), .ZN(n11119) );
  OR2_X2 U11346 ( .A1(n12908), .A2(n12962), .ZN(n11205) );
  INV_X2 U11347 ( .A(n15725), .ZN(n10844) );
  NOR2_X2 U11348 ( .A1(n13594), .A2(n13593), .ZN(n13944) );
  AND2_X2 U11349 ( .A1(n16212), .A2(n14499), .ZN(n9599) );
  INV_X1 U11350 ( .A(n10422), .ZN(n12558) );
  INV_X1 U11351 ( .A(n11161), .ZN(n9601) );
  INV_X2 U11352 ( .A(n11015), .ZN(n11161) );
  NAND2_X1 U11353 ( .A1(n10980), .A2(n13170), .ZN(n11015) );
  NAND2_X1 U11354 ( .A1(n10485), .A2(n10484), .ZN(n10516) );
  AND2_X4 U11355 ( .A1(n13156), .A2(n13140), .ZN(n11006) );
  NAND2_X1 U11356 ( .A1(n10461), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12776) );
  BUF_X8 U11357 ( .A(n11175), .Z(n9602) );
  INV_X1 U11358 ( .A(n14422), .ZN(n9610) );
  AND2_X4 U11359 ( .A1(n17047), .A2(n21204), .ZN(n12652) );
  INV_X1 U11360 ( .A(n10500), .ZN(n9604) );
  INV_X1 U11361 ( .A(n10500), .ZN(n9605) );
  OR3_X1 U11362 ( .A1(n12908), .A2(n20633), .A3(n14963), .ZN(n13199) );
  NAND2_X1 U11363 ( .A1(n10547), .A2(n10527), .ZN(n10645) );
  NOR2_X4 U11364 ( .A1(n19394), .A2(n14166), .ZN(n14232) );
  XNOR2_X2 U11365 ( .A(n14505), .B(n14504), .ZN(n14975) );
  NOR2_X1 U11366 ( .A1(n10830), .A2(n10831), .ZN(n10832) );
  BUF_X2 U11367 ( .A(n13183), .Z(n9606) );
  XNOR2_X1 U11368 ( .A(n11254), .B(n11253), .ZN(n13183) );
  NAND2_X2 U11369 ( .A1(n10818), .A2(n10817), .ZN(n13994) );
  AND2_X1 U11370 ( .A1(n10979), .A2(n13158), .ZN(n9608) );
  AND2_X1 U11371 ( .A1(n10979), .A2(n13158), .ZN(n11037) );
  NOR2_X1 U11372 ( .A1(n10411), .A2(n16237), .ZN(n12634) );
  NOR2_X1 U11373 ( .A1(n18141), .A2(n16436), .ZN(n19358) );
  INV_X2 U11374 ( .A(n9654), .ZN(n11859) );
  NOR2_X2 U11375 ( .A1(n14614), .A2(n10117), .ZN(n14565) );
  NAND2_X2 U11376 ( .A1(n14629), .A2(n14680), .ZN(n14614) );
  AND2_X2 U11377 ( .A1(n14486), .A2(n14499), .ZN(n9611) );
  INV_X2 U11378 ( .A(n10406), .ZN(n10150) );
  XNOR2_X1 U11379 ( .A(n10499), .B(n10498), .ZN(n10533) );
  INV_X1 U11380 ( .A(n13066), .ZN(n12010) );
  AOI211_X2 U11381 ( .C1(n16499), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16117), .B(n16116), .ZN(n16118) );
  NOR2_X2 U11382 ( .A1(n13911), .A2(n13924), .ZN(n13922) );
  OR2_X2 U11383 ( .A1(n13725), .A2(n13726), .ZN(n10818) );
  OAI21_X1 U11384 ( .B1(n13725), .B2(n10350), .A(n14109), .ZN(n13724) );
  INV_X2 U11385 ( .A(n11787), .ZN(n9613) );
  NAND2_X2 U11386 ( .A1(n13334), .A2(n11301), .ZN(n12060) );
  NOR2_X4 U11388 ( .A1(n15571), .A2(n15570), .ZN(n15569) );
  NOR2_X4 U11389 ( .A1(n14547), .A2(n14549), .ZN(n14535) );
  INV_X1 U11391 ( .A(n11015), .ZN(n9616) );
  XNOR2_X2 U11392 ( .A(n13651), .B(n11301), .ZN(n12069) );
  NAND2_X4 U11393 ( .A1(n9737), .A2(n11289), .ZN(n13651) );
  INV_X2 U11394 ( .A(n11835), .ZN(n9617) );
  AND2_X4 U11395 ( .A1(n13170), .A2(n13156), .ZN(n11089) );
  NOR2_X4 U11396 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13170) );
  INV_X2 U11397 ( .A(n9619), .ZN(n9620) );
  AND2_X1 U11398 ( .A1(n10974), .A2(n13170), .ZN(n11101) );
  NAND2_X1 U11399 ( .A1(n15544), .A2(n12494), .ZN(n12517) );
  OR2_X1 U11400 ( .A1(n12493), .A2(n12492), .ZN(n12494) );
  NOR2_X1 U11401 ( .A1(n10150), .A2(n10377), .ZN(n10452) );
  NAND2_X1 U11402 ( .A1(n12770), .A2(n9671), .ZN(n10082) );
  AND2_X1 U11403 ( .A1(n14406), .A2(n9776), .ZN(n9775) );
  OR2_X1 U11404 ( .A1(n10783), .A2(n10058), .ZN(n10057) );
  INV_X1 U11405 ( .A(n10067), .ZN(n10058) );
  AOI21_X1 U11406 ( .B1(n9784), .B2(n9786), .A(n9627), .ZN(n9781) );
  NAND2_X1 U11407 ( .A1(n10761), .A2(n9784), .ZN(n9782) );
  NAND2_X1 U11408 ( .A1(n10827), .A2(n10362), .ZN(n10675) );
  OR2_X1 U11409 ( .A1(n10140), .A2(n21068), .ZN(n10137) );
  CLKBUF_X1 U11410 ( .A(n12642), .Z(n17076) );
  AND2_X1 U11411 ( .A1(n11365), .A2(n11364), .ZN(n11374) );
  OAI22_X1 U11412 ( .A1(n10581), .A2(n20023), .B1(n10650), .B2(n10580), .ZN(
        n10582) );
  OAI22_X1 U11413 ( .A1(n10579), .A2(n10593), .B1(n10594), .B2(n12495), .ZN(
        n10583) );
  AOI21_X1 U11414 ( .B1(n10506), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10486), .ZN(n10489) );
  NAND2_X1 U11415 ( .A1(n12607), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10035) );
  NAND2_X1 U11416 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10034) );
  NAND2_X1 U11417 ( .A1(n10114), .A2(n14536), .ZN(n10113) );
  INV_X1 U11418 ( .A(n14524), .ZN(n10114) );
  NOR2_X1 U11419 ( .A1(n10121), .A2(n10120), .ZN(n10119) );
  INV_X1 U11420 ( .A(n14589), .ZN(n10120) );
  NAND2_X1 U11421 ( .A1(n14727), .A2(n9721), .ZN(n14708) );
  NOR2_X1 U11422 ( .A1(n9723), .A2(n9722), .ZN(n9721) );
  INV_X1 U11423 ( .A(n10123), .ZN(n9723) );
  NAND2_X1 U11424 ( .A1(n9740), .A2(n9738), .ZN(n12141) );
  AOI21_X1 U11425 ( .B1(n16656), .B2(n9742), .A(n9739), .ZN(n9738) );
  NAND2_X1 U11426 ( .A1(n14913), .A2(n16656), .ZN(n9740) );
  INV_X1 U11427 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9739) );
  NAND2_X1 U11428 ( .A1(n14973), .A2(n9832), .ZN(n10146) );
  INV_X1 U11429 ( .A(n11226), .ZN(n11184) );
  NAND2_X1 U11430 ( .A1(n11895), .A2(n11930), .ZN(n12904) );
  AOI21_X1 U11431 ( .B1(n9934), .B2(n9933), .A(n9934), .ZN(n9932) );
  INV_X1 U11432 ( .A(n9932), .ZN(n9930) );
  AND2_X1 U11433 ( .A1(n10773), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10684) );
  INV_X1 U11434 ( .A(n10183), .ZN(n10182) );
  AND2_X1 U11435 ( .A1(n9897), .A2(n15838), .ZN(n9896) );
  AOI21_X1 U11436 ( .B1(n15862), .B2(n15743), .A(n15745), .ZN(n9900) );
  NOR2_X1 U11437 ( .A1(n10457), .A2(n10456), .ZN(n10458) );
  NAND2_X1 U11438 ( .A1(n10455), .A2(n10454), .ZN(n10457) );
  AND2_X1 U11439 ( .A1(n18496), .A2(n18598), .ZN(n16413) );
  NAND2_X1 U11440 ( .A1(n16455), .A2(n16445), .ZN(n16396) );
  OR2_X1 U11441 ( .A1(n16645), .A2(n11204), .ZN(n14378) );
  AND2_X1 U11442 ( .A1(n11264), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12040) );
  NAND2_X1 U11443 ( .A1(n14808), .A2(n15123), .ZN(n10132) );
  OR2_X1 U11444 ( .A1(n12148), .A2(n14517), .ZN(n12149) );
  OAI21_X1 U11445 ( .B1(n13183), .B2(n12066), .A(n12049), .ZN(n13093) );
  XNOR2_X1 U11446 ( .A(n12143), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10140) );
  OR2_X1 U11447 ( .A1(n20838), .A2(n15132), .ZN(n16801) );
  AND2_X1 U11448 ( .A1(n16537), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14967) );
  NAND2_X1 U11449 ( .A1(n10763), .A2(n9904), .ZN(n16884) );
  INV_X1 U11450 ( .A(n10766), .ZN(n9904) );
  NAND2_X1 U11451 ( .A1(n10680), .A2(n10348), .ZN(n14414) );
  NOR2_X1 U11452 ( .A1(n10362), .A2(n10773), .ZN(n10348) );
  OR2_X1 U11453 ( .A1(n15552), .A2(n15637), .ZN(n9811) );
  NAND2_X1 U11454 ( .A1(n9651), .A2(n9810), .ZN(n9808) );
  NOR2_X1 U11455 ( .A1(n15552), .A2(n10191), .ZN(n9810) );
  NAND2_X1 U11456 ( .A1(n9651), .A2(n12467), .ZN(n9812) );
  INV_X1 U11457 ( .A(n9778), .ZN(n9771) );
  NAND2_X1 U11458 ( .A1(n10059), .A2(n10056), .ZN(n10053) );
  AND4_X1 U11459 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10347) );
  NAND2_X1 U11460 ( .A1(n9780), .A2(n9784), .ZN(n10065) );
  OR2_X1 U11461 ( .A1(n10761), .A2(n9786), .ZN(n9780) );
  AOI21_X1 U11462 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(n9787) );
  INV_X1 U11463 ( .A(n15731), .ZN(n9788) );
  NAND2_X1 U11464 ( .A1(n16191), .A2(n9764), .ZN(n9763) );
  NAND2_X1 U11465 ( .A1(n9766), .A2(n9634), .ZN(n9765) );
  AND2_X1 U11466 ( .A1(n16190), .A2(n9634), .ZN(n9764) );
  NAND2_X1 U11467 ( .A1(n13720), .A2(n13719), .ZN(n13750) );
  XNOR2_X1 U11468 ( .A(n14090), .B(n12158), .ZN(n13054) );
  INV_X1 U11469 ( .A(n20425), .ZN(n20395) );
  NAND2_X1 U11470 ( .A1(n16379), .A2(n18072), .ZN(n17158) );
  NAND2_X1 U11471 ( .A1(n18324), .A2(n9630), .ZN(n18260) );
  INV_X1 U11472 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9754) );
  OR2_X1 U11473 ( .A1(n16645), .A2(n13080), .ZN(n14788) );
  INV_X1 U11474 ( .A(n17156), .ZN(n18068) );
  AND2_X1 U11475 ( .A1(n9853), .A2(n9852), .ZN(n11356) );
  NAND2_X1 U11476 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n9852) );
  INV_X1 U11477 ( .A(n9839), .ZN(n11307) );
  OAI21_X1 U11478 ( .B1(n11859), .B2(n9841), .A(n9840), .ZN(n9839) );
  INV_X1 U11479 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n9841) );
  NAND2_X1 U11480 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n9840) );
  AND2_X1 U11481 ( .A1(n9849), .A2(n9848), .ZN(n11190) );
  NAND2_X1 U11482 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n9848) );
  AND2_X1 U11483 ( .A1(n14449), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10981) );
  AND2_X1 U11484 ( .A1(n9851), .A2(n9850), .ZN(n11233) );
  NAND2_X1 U11485 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n9850) );
  AND2_X1 U11486 ( .A1(n10402), .A2(n10430), .ZN(n12618) );
  NAND2_X1 U11487 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10078) );
  NAND2_X1 U11488 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10077) );
  NAND2_X1 U11489 ( .A1(n11890), .A2(n11889), .ZN(n11899) );
  OAI21_X1 U11490 ( .B1(n11859), .B2(n9837), .A(n9836), .ZN(n9835) );
  NAND2_X1 U11491 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U11492 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n9842) );
  NOR2_X1 U11493 ( .A1(n10099), .A2(n20963), .ZN(n9831) );
  NAND2_X1 U11494 ( .A1(n10478), .A2(n10451), .ZN(n10174) );
  NAND2_X1 U11495 ( .A1(n10453), .A2(n10445), .ZN(n10455) );
  AOI21_X1 U11496 ( .B1(n9605), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10504), .ZN(n10508) );
  AOI22_X1 U11497 ( .A1(n9610), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10503) );
  NAND2_X1 U11498 ( .A1(n13732), .A2(n19946), .ZN(n10173) );
  NAND2_X1 U11499 ( .A1(n12607), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10043) );
  NAND2_X1 U11500 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10042) );
  AND2_X1 U11501 ( .A1(n18515), .A2(n9624), .ZN(n9996) );
  OR2_X1 U11502 ( .A1(n11531), .A2(n20963), .ZN(n11883) );
  NOR2_X1 U11503 ( .A1(n14644), .A2(n10103), .ZN(n10102) );
  INV_X1 U11504 ( .A(n10105), .ZN(n10103) );
  AND2_X1 U11505 ( .A1(n14701), .A2(n10106), .ZN(n10105) );
  INV_X1 U11506 ( .A(n14709), .ZN(n10106) );
  NOR2_X1 U11507 ( .A1(n11551), .A2(n16595), .ZN(n11552) );
  INV_X1 U11508 ( .A(n13912), .ZN(n11388) );
  XNOR2_X1 U11509 ( .A(n11366), .B(n11374), .ZN(n12097) );
  INV_X1 U11510 ( .A(n13648), .ZN(n11372) );
  INV_X1 U11511 ( .A(n11290), .ZN(n11524) );
  INV_X1 U11512 ( .A(n14553), .ZN(n9977) );
  AND2_X1 U11513 ( .A1(n14581), .A2(n14570), .ZN(n9978) );
  AND2_X1 U11514 ( .A1(n11376), .A2(n11375), .ZN(n11377) );
  INV_X1 U11515 ( .A(n11373), .ZN(n11378) );
  NOR2_X1 U11516 ( .A1(n13937), .A2(n13936), .ZN(n9984) );
  AND2_X1 U11517 ( .A1(n9847), .A2(n9846), .ZN(n11173) );
  NAND2_X1 U11518 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n9846) );
  NAND2_X1 U11519 ( .A1(n11217), .A2(n11216), .ZN(n11224) );
  OAI211_X1 U11520 ( .C1(n16537), .C2(n16513), .A(n11222), .B(n11221), .ZN(
        n11223) );
  AND2_X1 U11521 ( .A1(n13123), .A2(n13122), .ZN(n13175) );
  INV_X1 U11522 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16513) );
  NAND2_X1 U11523 ( .A1(n10357), .A2(n10776), .ZN(n14410) );
  INV_X1 U11524 ( .A(n10778), .ZN(n10357) );
  NOR2_X1 U11525 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n16871), .ZN(n10771) );
  AND2_X1 U11526 ( .A1(n10764), .A2(n14414), .ZN(n10715) );
  NOR2_X1 U11527 ( .A1(n9911), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n9910) );
  INV_X1 U11528 ( .A(n9912), .ZN(n9911) );
  AND2_X1 U11529 ( .A1(n10688), .A2(n10351), .ZN(n10695) );
  AND4_X1 U11530 ( .A1(n9907), .A2(n10673), .A3(n10639), .A4(n9908), .ZN(
        n10680) );
  INV_X1 U11531 ( .A(n10631), .ZN(n9907) );
  NOR2_X1 U11532 ( .A1(n10630), .A2(n10626), .ZN(n9908) );
  NOR2_X1 U11533 ( .A1(n10444), .A2(n19946), .ZN(n10431) );
  NOR2_X1 U11534 ( .A1(n10081), .A2(n12848), .ZN(n10080) );
  INV_X1 U11535 ( .A(n15497), .ZN(n10081) );
  OR2_X1 U11536 ( .A1(n12558), .A2(n10416), .ZN(n12272) );
  OR2_X1 U11537 ( .A1(n10221), .A2(n10416), .ZN(n12315) );
  INV_X1 U11538 ( .A(n15627), .ZN(n10162) );
  INV_X1 U11539 ( .A(n15563), .ZN(n10190) );
  INV_X1 U11540 ( .A(n10061), .ZN(n10056) );
  OAI21_X1 U11541 ( .B1(n10775), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10062), .ZN(n10061) );
  NOR2_X1 U11542 ( .A1(n10066), .A2(n10063), .ZN(n10062) );
  NOR2_X1 U11543 ( .A1(n10350), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10063) );
  AOI21_X1 U11544 ( .B1(n9787), .B2(n15730), .A(n9785), .ZN(n9784) );
  INV_X1 U11545 ( .A(n15722), .ZN(n9785) );
  NOR2_X1 U11546 ( .A1(n10087), .A2(n15420), .ZN(n10086) );
  INV_X1 U11547 ( .A(n15435), .ZN(n10087) );
  NAND2_X1 U11548 ( .A1(n10168), .A2(n15437), .ZN(n10167) );
  INV_X1 U11549 ( .A(n15650), .ZN(n10168) );
  AND2_X1 U11550 ( .A1(n9889), .A2(n9888), .ZN(n9887) );
  NAND2_X1 U11551 ( .A1(n15748), .A2(n15799), .ZN(n9888) );
  NOR2_X1 U11552 ( .A1(n15749), .A2(n9890), .ZN(n9889) );
  OR2_X1 U11553 ( .A1(n19623), .A2(n10362), .ZN(n10749) );
  AND2_X1 U11554 ( .A1(n10892), .A2(n10891), .ZN(n15582) );
  NOR2_X1 U11555 ( .A1(n10154), .A2(n15470), .ZN(n10153) );
  NAND2_X1 U11556 ( .A1(n10155), .A2(n16964), .ZN(n10154) );
  INV_X1 U11557 ( .A(n15481), .ZN(n10155) );
  OR2_X1 U11558 ( .A1(n10328), .A2(n10327), .ZN(n12687) );
  AND2_X1 U11559 ( .A1(n10625), .A2(n10362), .ZN(n9768) );
  NOR2_X1 U11560 ( .A1(n19740), .A2(n10149), .ZN(n10148) );
  INV_X1 U11561 ( .A(n13743), .ZN(n10149) );
  OR2_X1 U11562 ( .A1(n10234), .A2(n10233), .ZN(n12676) );
  NAND2_X1 U11563 ( .A1(n10016), .A2(n10574), .ZN(n10629) );
  NAND2_X1 U11564 ( .A1(n9604), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U11565 ( .A1(n12183), .A2(n21204), .ZN(n12177) );
  NAND2_X1 U11566 ( .A1(n10492), .A2(n10491), .ZN(n10512) );
  NOR2_X1 U11567 ( .A1(n17055), .A2(n17076), .ZN(n13707) );
  NAND2_X1 U11568 ( .A1(n10545), .A2(n10549), .ZN(n10614) );
  NAND2_X1 U11569 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10030) );
  NAND2_X1 U11570 ( .A1(n12605), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10031) );
  INV_X1 U11571 ( .A(n18938), .ZN(n16273) );
  INV_X1 U11572 ( .A(n16387), .ZN(n14256) );
  INV_X1 U11573 ( .A(n16334), .ZN(n14332) );
  OR2_X1 U11574 ( .A1(n17648), .A2(n14173), .ZN(n10198) );
  NOR2_X1 U11575 ( .A1(n14172), .A2(n17648), .ZN(n16387) );
  NOR2_X1 U11576 ( .A1(n18581), .A2(n9963), .ZN(n9962) );
  INV_X1 U11577 ( .A(n17492), .ZN(n9953) );
  NOR2_X1 U11578 ( .A1(n18505), .A2(n18831), .ZN(n16466) );
  NAND2_X1 U11579 ( .A1(n16399), .A2(n18080), .ZN(n16380) );
  NOR2_X1 U11580 ( .A1(n16396), .A2(n18084), .ZN(n16399) );
  INV_X1 U11581 ( .A(n16396), .ZN(n16452) );
  XNOR2_X1 U11582 ( .A(n18088), .B(n16455), .ZN(n16381) );
  AOI22_X1 U11583 ( .A1(n18916), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n14253), .B2(n14252), .ZN(n16265) );
  OR2_X1 U11584 ( .A1(n14250), .A2(n16421), .ZN(n16267) );
  AND2_X1 U11585 ( .A1(n11886), .A2(n11532), .ZN(n14981) );
  OR2_X1 U11586 ( .A1(n14030), .A2(n11457), .ZN(n11458) );
  NOR2_X1 U11587 ( .A1(n11113), .A2(n11112), .ZN(n11114) );
  NAND2_X1 U11588 ( .A1(n11715), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11759) );
  NAND2_X1 U11589 ( .A1(n10119), .A2(n10118), .ZN(n10117) );
  INV_X1 U11590 ( .A(n14578), .ZN(n10118) );
  INV_X1 U11591 ( .A(n14614), .ZN(n10116) );
  NAND2_X1 U11592 ( .A1(n12139), .A2(n15123), .ZN(n14882) );
  NAND2_X1 U11593 ( .A1(n9869), .A2(n9648), .ZN(n12139) );
  NAND2_X1 U11594 ( .A1(n13922), .A2(n10108), .ZN(n14030) );
  AND2_X1 U11595 ( .A1(n14031), .A2(n13973), .ZN(n10108) );
  INV_X1 U11596 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11383) );
  NAND2_X1 U11597 ( .A1(n11367), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11381) );
  NAND2_X1 U11598 ( .A1(n11321), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U11599 ( .A1(n13064), .A2(n13065), .ZN(n13269) );
  AND2_X1 U11600 ( .A1(n14865), .A2(n9875), .ZN(n14827) );
  NAND2_X1 U11601 ( .A1(n16656), .A2(n15009), .ZN(n9875) );
  OR2_X1 U11602 ( .A1(n16730), .A2(n15008), .ZN(n15057) );
  NAND2_X1 U11603 ( .A1(n9743), .A2(n12137), .ZN(n14915) );
  NAND2_X1 U11604 ( .A1(n14134), .A2(n9629), .ZN(n9744) );
  NAND2_X1 U11605 ( .A1(n14159), .A2(n14158), .ZN(n14729) );
  NAND2_X1 U11606 ( .A1(n9984), .A2(n9983), .ZN(n14032) );
  INV_X1 U11607 ( .A(n13980), .ZN(n9983) );
  NAND2_X1 U11608 ( .A1(n16698), .A2(n16697), .ZN(n16696) );
  AND2_X1 U11609 ( .A1(n14992), .A2(n14986), .ZN(n15132) );
  OR2_X1 U11610 ( .A1(n11183), .A2(n11200), .ZN(n10145) );
  INV_X1 U11611 ( .A(n12069), .ZN(n9746) );
  NAND2_X1 U11612 ( .A1(n11944), .A2(n11943), .ZN(n14963) );
  NAND2_X1 U11613 ( .A1(n11909), .A2(n11896), .ZN(n11944) );
  NAND2_X1 U11614 ( .A1(n11942), .A2(n11941), .ZN(n11943) );
  NOR2_X1 U11615 ( .A1(n13496), .A2(n12069), .ZN(n13504) );
  AND2_X1 U11616 ( .A1(n12069), .A2(n12060), .ZN(n13452) );
  NOR2_X1 U11617 ( .A1(n20861), .A2(n13768), .ZN(n20904) );
  NAND2_X1 U11618 ( .A1(n13150), .A2(n20963), .ZN(n9737) );
  AOI21_X1 U11619 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20864), .A(n13768), 
        .ZN(n13536) );
  NAND2_X1 U11620 ( .A1(n10442), .A2(n19936), .ZN(n12841) );
  AOI21_X1 U11621 ( .B1(n9932), .B2(n9929), .A(n9928), .ZN(n9927) );
  INV_X1 U11622 ( .A(n9933), .ZN(n9929) );
  NOR2_X1 U11623 ( .A1(n9930), .A2(n9934), .ZN(n9926) );
  NOR2_X1 U11624 ( .A1(n9930), .A2(n9935), .ZN(n9924) );
  NAND2_X1 U11625 ( .A1(n14414), .A2(n10725), .ZN(n10716) );
  OR2_X1 U11626 ( .A1(n10724), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10725) );
  AND2_X1 U11627 ( .A1(n9921), .A2(n9920), .ZN(n9919) );
  AND2_X1 U11628 ( .A1(n10351), .A2(n19783), .ZN(n9921) );
  NOR2_X1 U11629 ( .A1(n10686), .A2(n10684), .ZN(n10688) );
  AND2_X1 U11630 ( .A1(n14414), .A2(n10703), .ZN(n10701) );
  OAI21_X1 U11631 ( .B1(n12827), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12826), 
        .ZN(n15305) );
  OR2_X1 U11632 ( .A1(n17050), .A2(n12859), .ZN(n12881) );
  INV_X1 U11633 ( .A(n19737), .ZN(n19652) );
  OR2_X1 U11634 ( .A1(n12311), .A2(n12310), .ZN(n13847) );
  NAND2_X1 U11635 ( .A1(n9691), .A2(n12216), .ZN(n10183) );
  OR2_X1 U11636 ( .A1(n12201), .A2(n12200), .ZN(n12690) );
  NAND2_X1 U11637 ( .A1(n15536), .A2(n9670), .ZN(n9793) );
  INV_X1 U11638 ( .A(n12545), .ZN(n9792) );
  NAND2_X1 U11639 ( .A1(n10186), .A2(n12467), .ZN(n10185) );
  NAND2_X1 U11640 ( .A1(n15567), .A2(n10191), .ZN(n10184) );
  OR2_X1 U11641 ( .A1(n15638), .A2(n15637), .ZN(n9813) );
  NAND2_X1 U11642 ( .A1(n12725), .A2(n10163), .ZN(n16041) );
  NOR2_X1 U11643 ( .A1(n10165), .A2(n10164), .ZN(n10163) );
  INV_X1 U11644 ( .A(n16040), .ZN(n10164) );
  NAND2_X1 U11645 ( .A1(n10186), .A2(n9825), .ZN(n9823) );
  OR2_X1 U11646 ( .A1(n15328), .A2(n15700), .ZN(n15332) );
  AND2_X1 U11647 ( .A1(n15318), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15320) );
  INV_X1 U11648 ( .A(n9591), .ZN(n14424) );
  NAND2_X1 U11649 ( .A1(n9777), .A2(n9775), .ZN(n15662) );
  NAND2_X1 U11650 ( .A1(n10090), .A2(n10089), .ZN(n10088) );
  INV_X1 U11651 ( .A(n10091), .ZN(n10090) );
  NOR2_X1 U11652 ( .A1(n15546), .A2(n15373), .ZN(n10089) );
  OR2_X1 U11653 ( .A1(n15391), .A2(n10362), .ZN(n15677) );
  NOR2_X1 U11654 ( .A1(n16854), .A2(n9701), .ZN(n10783) );
  NAND2_X1 U11655 ( .A1(n9660), .A2(n9791), .ZN(n9790) );
  NOR2_X1 U11656 ( .A1(n15752), .A2(n15750), .ZN(n9791) );
  NAND2_X1 U11657 ( .A1(n10744), .A2(n9688), .ZN(n10068) );
  AND2_X1 U11658 ( .A1(n9883), .A2(n9891), .ZN(n9882) );
  INV_X1 U11659 ( .A(n15751), .ZN(n9891) );
  NAND2_X1 U11660 ( .A1(n9887), .A2(n9884), .ZN(n9883) );
  INV_X1 U11661 ( .A(n15799), .ZN(n9884) );
  INV_X1 U11662 ( .A(n9887), .ZN(n9885) );
  NAND2_X1 U11663 ( .A1(n10152), .A2(n10151), .ZN(n15453) );
  AND2_X1 U11664 ( .A1(n10153), .A2(n14099), .ZN(n10151) );
  OAI21_X1 U11665 ( .B1(n15827), .B2(n15746), .A(n15826), .ZN(n15814) );
  AOI21_X1 U11666 ( .B1(n9900), .B2(n15744), .A(n9898), .ZN(n9897) );
  INV_X1 U11667 ( .A(n15852), .ZN(n9898) );
  INV_X1 U11668 ( .A(n9900), .ZN(n9899) );
  NAND2_X1 U11669 ( .A1(n10073), .A2(n10071), .ZN(n15742) );
  OR2_X1 U11670 ( .A1(n15863), .A2(n15862), .ZN(n9901) );
  AND2_X1 U11671 ( .A1(n19682), .A2(n10697), .ZN(n16161) );
  INV_X1 U11672 ( .A(n14056), .ZN(n10159) );
  INV_X1 U11673 ( .A(n10677), .ZN(n10052) );
  NAND2_X1 U11674 ( .A1(n13722), .A2(n10049), .ZN(n10048) );
  NAND2_X1 U11675 ( .A1(n10047), .A2(n9639), .ZN(n10046) );
  INV_X1 U11676 ( .A(n13724), .ZN(n10047) );
  NAND2_X1 U11677 ( .A1(n10046), .A2(n10045), .ZN(n13999) );
  AND2_X1 U11678 ( .A1(n10048), .A2(n10050), .ZN(n10045) );
  INV_X1 U11679 ( .A(n13996), .ZN(n10050) );
  OAI22_X1 U11680 ( .A1(n10506), .A2(n10466), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10501), .ZN(n10470) );
  NOR2_X1 U11681 ( .A1(n9818), .A2(n12156), .ZN(n9816) );
  INV_X1 U11682 ( .A(n9822), .ZN(n9821) );
  NAND2_X1 U11683 ( .A1(n9795), .A2(n12160), .ZN(n13061) );
  NAND2_X1 U11684 ( .A1(n13054), .A2(n13055), .ZN(n9795) );
  OR2_X1 U11685 ( .A1(n20054), .A2(n20599), .ZN(n20360) );
  NAND2_X1 U11686 ( .A1(n10399), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10400) );
  NAND2_X1 U11687 ( .A1(n10394), .A2(n10416), .ZN(n10401) );
  AND2_X1 U11688 ( .A1(n10956), .A2(n19598), .ZN(n20425) );
  OR2_X1 U11689 ( .A1(n20054), .A2(n16223), .ZN(n20429) );
  AND2_X1 U11690 ( .A1(n9946), .A2(n9683), .ZN(n17386) );
  OR2_X1 U11691 ( .A1(n17655), .A2(n18304), .ZN(n9947) );
  BUF_X1 U11692 ( .A(n14284), .Z(n17763) );
  OAI221_X1 U11693 ( .B1(n16560), .B2(n16559), .C1(n16560), .C2(n16558), .A(
        n19572), .ZN(n16562) );
  NOR3_X1 U11694 ( .A1(n16557), .A2(n18102), .A3(n19574), .ZN(n16560) );
  NOR4_X2 U11695 ( .A1(n18923), .A2(n16434), .A3(n16270), .A4(n16272), .ZN(
        n18141) );
  NOR2_X1 U11696 ( .A1(n9951), .A2(n9952), .ZN(n9950) );
  NOR2_X1 U11697 ( .A1(n18419), .A2(n18421), .ZN(n18408) );
  INV_X1 U11698 ( .A(n18782), .ZN(n18454) );
  NOR2_X1 U11699 ( .A1(n18220), .A2(n18219), .ZN(n18218) );
  INV_X1 U11700 ( .A(n16414), .ZN(n9752) );
  INV_X1 U11701 ( .A(n18240), .ZN(n9753) );
  NAND2_X1 U11702 ( .A1(n10005), .A2(n9686), .ZN(n10004) );
  NAND2_X1 U11703 ( .A1(n18293), .A2(n18272), .ZN(n10005) );
  INV_X1 U11704 ( .A(n18260), .ZN(n18264) );
  INV_X1 U11705 ( .A(n18496), .ZN(n18404) );
  INV_X1 U11706 ( .A(n18374), .ZN(n18293) );
  NOR2_X1 U11707 ( .A1(n18373), .A2(n16410), .ZN(n18363) );
  AOI22_X1 U11708 ( .A1(n18374), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n18711), .B2(n18496), .ZN(n16409) );
  NAND2_X1 U11709 ( .A1(n18529), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10000) );
  NOR2_X1 U11710 ( .A1(n16419), .A2(n16418), .ZN(n19364) );
  INV_X1 U11711 ( .A(n14967), .ZN(n20633) );
  INV_X1 U11712 ( .A(n14815), .ZN(n9981) );
  OAI21_X1 U11713 ( .B1(n15025), .B2(n20666), .A(n9979), .ZN(n9730) );
  NOR2_X1 U11714 ( .A1(n14518), .A2(n9980), .ZN(n9979) );
  AND2_X1 U11715 ( .A1(n20684), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n9980) );
  AND2_X1 U11716 ( .A1(n13584), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13575) );
  INV_X1 U11717 ( .A(n20700), .ZN(n20666) );
  INV_X1 U11718 ( .A(n14788), .ZN(n16647) );
  NAND2_X1 U11719 ( .A1(n13107), .A2(n13076), .ZN(n13077) );
  AND2_X1 U11720 ( .A1(n13121), .A2(n13075), .ZN(n13076) );
  NOR2_X1 U11721 ( .A1(n10137), .A2(n14998), .ZN(n10135) );
  AND2_X1 U11722 ( .A1(n14535), .A2(n10109), .ZN(n12042) );
  AND2_X1 U11723 ( .A1(n10112), .A2(n10110), .ZN(n10109) );
  AND2_X1 U11724 ( .A1(n10139), .A2(n20792), .ZN(n10136) );
  AOI21_X1 U11725 ( .B1(n14808), .B2(n10134), .A(n10130), .ZN(n10129) );
  INV_X1 U11726 ( .A(n12152), .ZN(n10130) );
  NOR2_X1 U11727 ( .A1(n10137), .A2(n16656), .ZN(n10134) );
  NAND2_X1 U11728 ( .A1(n11217), .A2(n13653), .ZN(n20896) );
  NAND2_X1 U11729 ( .A1(n13415), .A2(n9745), .ZN(n15165) );
  NAND2_X1 U11730 ( .A1(n9747), .A2(n9746), .ZN(n9745) );
  INV_X1 U11731 ( .A(n13416), .ZN(n9747) );
  NOR2_X1 U11732 ( .A1(n12881), .A2(n12630), .ZN(n19599) );
  INV_X1 U11733 ( .A(n10763), .ZN(n10767) );
  AND2_X1 U11734 ( .A1(n10709), .A2(n10711), .ZN(n15446) );
  INV_X1 U11735 ( .A(n19744), .ZN(n19683) );
  INV_X1 U11736 ( .A(n19802), .ZN(n15640) );
  OR2_X1 U11737 ( .A1(n12871), .A2(n13734), .ZN(n12635) );
  NOR2_X1 U11738 ( .A1(n14090), .A2(n12990), .ZN(n16222) );
  AND2_X1 U11739 ( .A1(n19834), .A2(n12645), .ZN(n19848) );
  INV_X1 U11740 ( .A(n15933), .ZN(n16955) );
  INV_X1 U11741 ( .A(n13859), .ZN(n16946) );
  NAND2_X1 U11742 ( .A1(n9995), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9991) );
  NAND2_X1 U11743 ( .A1(n15682), .A2(n9718), .ZN(n9992) );
  OAI21_X1 U11744 ( .B1(n10781), .B2(n9773), .A(n9770), .ZN(n14418) );
  AND2_X1 U11745 ( .A1(n13750), .A2(n20621), .ZN(n17013) );
  INV_X2 U11746 ( .A(n19920), .ZN(n17009) );
  NAND2_X1 U11747 ( .A1(n13750), .A2(n13749), .ZN(n19911) );
  INV_X1 U11748 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20615) );
  INV_X1 U11749 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20605) );
  INV_X1 U11750 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20597) );
  NOR2_X2 U11751 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20585) );
  NOR2_X1 U11752 ( .A1(n20147), .A2(n20360), .ZN(n20125) );
  INV_X1 U11753 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19598) );
  NOR2_X1 U11754 ( .A1(n9968), .A2(n9967), .ZN(n9966) );
  NOR2_X1 U11755 ( .A1(n9645), .A2(n17655), .ZN(n9967) );
  INV_X1 U11756 ( .A(n9969), .ZN(n9968) );
  AOI21_X1 U11757 ( .B1(n17323), .B2(n17314), .A(n17313), .ZN(n9969) );
  AND2_X1 U11758 ( .A1(n9949), .A2(n17655), .ZN(n17400) );
  NOR2_X1 U11759 ( .A1(n19524), .A2(n17649), .ZN(n17564) );
  INV_X1 U11760 ( .A(n17564), .ZN(n17652) );
  INV_X1 U11761 ( .A(n17663), .ZN(n17650) );
  NOR2_X1 U11762 ( .A1(n9756), .A2(n17109), .ZN(n9755) );
  INV_X1 U11763 ( .A(n17122), .ZN(n9756) );
  XNOR2_X1 U11764 ( .A(n9757), .B(n17109), .ZN(n17121) );
  NAND2_X1 U11765 ( .A1(n9758), .A2(n17094), .ZN(n9757) );
  INV_X1 U11766 ( .A(n17092), .ZN(n9758) );
  OAI21_X1 U11767 ( .B1(n18218), .B2(n17159), .A(n10012), .ZN(n10011) );
  AND2_X1 U11768 ( .A1(n10014), .A2(n10013), .ZN(n10012) );
  OAI21_X1 U11769 ( .B1(n18228), .B2(n17158), .A(n17157), .ZN(n17159) );
  OR2_X1 U11770 ( .A1(n17160), .A2(n18755), .ZN(n10014) );
  NAND2_X1 U11771 ( .A1(n10009), .A2(n10008), .ZN(n10007) );
  INV_X1 U11772 ( .A(n18214), .ZN(n10008) );
  NAND2_X1 U11773 ( .A1(n18660), .A2(n18223), .ZN(n10009) );
  OR2_X1 U11774 ( .A1(n20111), .A2(n12549), .ZN(n10616) );
  AOI21_X1 U11775 ( .B1(n9616), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A(n9867), 
        .ZN(n11840) );
  NOR2_X1 U11776 ( .A1(n11859), .A2(n9868), .ZN(n9867) );
  INV_X1 U11777 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n9868) );
  AND2_X1 U11778 ( .A1(n9866), .A2(n9864), .ZN(n11820) );
  NAND2_X1 U11779 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n9864) );
  AND2_X1 U11780 ( .A1(n9863), .A2(n9862), .ZN(n11772) );
  NAND2_X1 U11781 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n9862) );
  AND2_X1 U11782 ( .A1(n9859), .A2(n9858), .ZN(n11726) );
  NAND2_X1 U11783 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n9858) );
  AND2_X1 U11784 ( .A1(n9845), .A2(n9844), .ZN(n11501) );
  NAND2_X1 U11785 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n9844) );
  INV_X1 U11786 ( .A(n10609), .ZN(n10019) );
  AOI21_X1 U11787 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n19403), .A(
        n14244), .ZN(n14245) );
  AND2_X1 U11788 ( .A1(n9861), .A2(n9860), .ZN(n11576) );
  NAND2_X1 U11789 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n9860) );
  AND2_X1 U11790 ( .A1(n9855), .A2(n9854), .ZN(n11522) );
  NAND2_X1 U11791 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U11792 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11616) );
  AND2_X1 U11793 ( .A1(n9857), .A2(n9856), .ZN(n11485) );
  NAND2_X1 U11794 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U11795 ( .A1(n9828), .A2(n13651), .ZN(n11326) );
  INV_X1 U11796 ( .A(n11301), .ZN(n9828) );
  OR2_X1 U11797 ( .A1(n9588), .A2(n12126), .ZN(n12134) );
  OR2_X1 U11798 ( .A1(n11363), .A2(n11362), .ZN(n12107) );
  OR2_X1 U11799 ( .A1(n11339), .A2(n11338), .ZN(n12099) );
  OR2_X1 U11800 ( .A1(n11314), .A2(n11313), .ZN(n12090) );
  INV_X1 U11801 ( .A(n12066), .ZN(n12105) );
  AND2_X1 U11802 ( .A1(n11125), .A2(n16528), .ZN(n13112) );
  INV_X1 U11803 ( .A(n13155), .ZN(n13127) );
  OR2_X1 U11804 ( .A1(n11198), .A2(n11197), .ZN(n12052) );
  OR2_X1 U11805 ( .A1(n11240), .A2(n11239), .ZN(n12061) );
  AND2_X1 U11806 ( .A1(n13166), .A2(n13165), .ZN(n16514) );
  NAND2_X1 U11807 ( .A1(n10220), .A2(n10219), .ZN(n10303) );
  OR2_X1 U11808 ( .A1(n10275), .A2(n10218), .ZN(n10220) );
  XNOR2_X1 U11809 ( .A(n10416), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10302) );
  NOR2_X1 U11810 ( .A1(n10303), .A2(n10302), .ZN(n10305) );
  AOI21_X1 U11811 ( .B1(n12368), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A(n9902), .ZN(n10297) );
  OAI21_X1 U11812 ( .B1(n12431), .B2(n19950), .A(n9903), .ZN(n9902) );
  NAND2_X1 U11813 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9903) );
  INV_X1 U11814 ( .A(n12429), .ZN(n12350) );
  OR2_X1 U11815 ( .A1(n10273), .A2(n10272), .ZN(n10573) );
  AND2_X1 U11816 ( .A1(n13721), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10084) );
  INV_X1 U11817 ( .A(n15786), .ZN(n9890) );
  AOI21_X1 U11818 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20588), .A(
        n10305), .ZN(n10786) );
  NAND2_X1 U11819 ( .A1(n10420), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10025) );
  NAND2_X1 U11820 ( .A1(n10420), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10027) );
  NAND4_X1 U11821 ( .A1(n10212), .A2(n10211), .A3(n10210), .A4(n10209), .ZN(
        n10213) );
  AOI22_X1 U11822 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10365) );
  NAND2_X1 U11823 ( .A1(n19554), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14171) );
  NAND2_X1 U11824 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19531), .ZN(
        n14173) );
  NAND2_X1 U11825 ( .A1(n11683), .A2(n10122), .ZN(n10121) );
  INV_X1 U11826 ( .A(n14616), .ZN(n10122) );
  INV_X1 U11827 ( .A(n11883), .ZN(n11849) );
  AND2_X1 U11828 ( .A1(n11493), .A2(n14726), .ZN(n10123) );
  INV_X1 U11829 ( .A(n9835), .ZN(n11448) );
  NAND2_X1 U11830 ( .A1(n11420), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11440) );
  NOR2_X1 U11831 ( .A1(n11405), .A2(n14137), .ZN(n11420) );
  AND2_X1 U11832 ( .A1(n9843), .A2(n9842), .ZN(n11411) );
  INV_X1 U11833 ( .A(n13525), .ZN(n9732) );
  INV_X1 U11834 ( .A(n13301), .ZN(n11255) );
  NAND2_X1 U11835 ( .A1(n11116), .A2(n14978), .ZN(n12066) );
  NOR2_X1 U11836 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n9872) );
  NOR2_X1 U11837 ( .A1(n14692), .A2(n14691), .ZN(n9975) );
  NAND2_X1 U11838 ( .A1(n11132), .A2(n9658), .ZN(n11137) );
  INV_X1 U11839 ( .A(n12044), .ZN(n11200) );
  INV_X1 U11840 ( .A(n11940), .ZN(n11941) );
  AOI21_X1 U11841 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20963), .A(
        n11939), .ZN(n11940) );
  OR2_X1 U11842 ( .A1(n11934), .A2(n12904), .ZN(n11942) );
  NAND2_X1 U11843 ( .A1(n11135), .A2(n9831), .ZN(n9829) );
  OAI21_X1 U11844 ( .B1(n11859), .B2(n9838), .A(n9834), .ZN(n9833) );
  INV_X1 U11845 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U11846 ( .A1(n11175), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11091) );
  OAI21_X1 U11847 ( .B1(n21054), .B2(n13181), .A(n15186), .ZN(n13287) );
  OR2_X1 U11848 ( .A1(n11288), .A2(n11287), .ZN(n12080) );
  AND2_X1 U11849 ( .A1(n11184), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11935) );
  AND2_X1 U11850 ( .A1(n13179), .A2(n13178), .ZN(n16518) );
  XNOR2_X1 U11851 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10939) );
  NOR2_X1 U11852 ( .A1(n9914), .A2(n9913), .ZN(n9912) );
  INV_X1 U11853 ( .A(n10353), .ZN(n9913) );
  NOR2_X1 U11854 ( .A1(n9918), .A2(n10730), .ZN(n9917) );
  INV_X1 U11855 ( .A(n15520), .ZN(n9804) );
  AND2_X1 U11856 ( .A1(n15532), .A2(n15527), .ZN(n9807) );
  NOR2_X1 U11857 ( .A1(n10187), .A2(n16904), .ZN(n10186) );
  INV_X1 U11858 ( .A(n10189), .ZN(n10187) );
  INV_X1 U11859 ( .A(n15568), .ZN(n9826) );
  NOR2_X1 U11860 ( .A1(n15734), .A2(n9945), .ZN(n9944) );
  INV_X1 U11861 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9945) );
  AND2_X1 U11862 ( .A1(n13243), .A2(n14051), .ZN(n10097) );
  NAND2_X1 U11863 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9942) );
  INV_X1 U11864 ( .A(n10573), .ZN(n12665) );
  NAND2_X1 U11865 ( .A1(n15538), .A2(n15388), .ZN(n10091) );
  NOR2_X1 U11866 ( .A1(n10780), .A2(n9779), .ZN(n9778) );
  INV_X1 U11867 ( .A(n15674), .ZN(n9779) );
  NAND2_X1 U11868 ( .A1(n10782), .A2(n21106), .ZN(n10067) );
  INV_X1 U11869 ( .A(n9787), .ZN(n9786) );
  NOR2_X1 U11870 ( .A1(n21106), .A2(n16027), .ZN(n10003) );
  INV_X1 U11871 ( .A(n15735), .ZN(n10085) );
  INV_X1 U11872 ( .A(n10071), .ZN(n10070) );
  NAND2_X1 U11873 ( .A1(n10166), .A2(n15422), .ZN(n10165) );
  INV_X1 U11874 ( .A(n10167), .ZN(n10166) );
  AND2_X1 U11875 ( .A1(n12709), .A2(n12708), .ZN(n15494) );
  NOR2_X1 U11876 ( .A1(n10698), .A2(n10072), .ZN(n10071) );
  INV_X1 U11877 ( .A(n16142), .ZN(n10072) );
  AND2_X1 U11878 ( .A1(n10096), .A2(n10097), .ZN(n10095) );
  INV_X1 U11879 ( .A(n13365), .ZN(n10096) );
  INV_X1 U11880 ( .A(n10823), .ZN(n10831) );
  NAND2_X1 U11881 ( .A1(n10015), .A2(n10592), .ZN(n10628) );
  NAND2_X1 U11882 ( .A1(n10449), .A2(n10448), .ZN(n10483) );
  NAND2_X1 U11883 ( .A1(n19962), .A2(n10377), .ZN(n12656) );
  OR2_X1 U11884 ( .A1(n10289), .A2(n10288), .ZN(n12655) );
  AOI21_X1 U11885 ( .B1(n10501), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10474), .ZN(
        n10477) );
  OR2_X1 U11886 ( .A1(n14422), .A2(n10475), .ZN(n10476) );
  AND2_X1 U11887 ( .A1(n10174), .A2(n13731), .ZN(n10479) );
  INV_X1 U11888 ( .A(n10444), .ZN(n13728) );
  NAND2_X1 U11889 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n9761) );
  NAND2_X1 U11890 ( .A1(n9611), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n9760) );
  NOR2_X1 U11891 ( .A1(n17273), .A2(n16432), .ZN(n16436) );
  NOR2_X1 U11892 ( .A1(n19394), .A2(n14173), .ZN(n16334) );
  INV_X1 U11893 ( .A(n16386), .ZN(n17847) );
  OR2_X1 U11894 ( .A1(n14167), .A2(n14171), .ZN(n16345) );
  OR2_X1 U11895 ( .A1(n14173), .A2(n14171), .ZN(n10197) );
  OR2_X1 U11896 ( .A1(n14172), .A2(n14171), .ZN(n14354) );
  NAND2_X1 U11897 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19541), .ZN(
        n14167) );
  OR3_X1 U11898 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19531), .A3(
        n19391), .ZN(n16247) );
  NAND2_X1 U11899 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18408), .ZN(
        n18376) );
  NAND2_X1 U11900 ( .A1(n9997), .A2(n9998), .ZN(n16403) );
  AOI21_X1 U11901 ( .B1(n18515), .B2(n9999), .A(n9666), .ZN(n9998) );
  INV_X1 U11902 ( .A(n10000), .ZN(n9999) );
  NOR2_X1 U11903 ( .A1(n19368), .A2(n16288), .ZN(n16268) );
  INV_X1 U11904 ( .A(n16563), .ZN(n19381) );
  AOI22_X1 U11905 ( .A1(n19359), .A2(n18753), .B1(n17090), .B2(n19364), .ZN(
        n17101) );
  OAI21_X1 U11906 ( .B1(n16436), .B2(n19415), .A(n19573), .ZN(n18100) );
  OAI21_X1 U11907 ( .B1(n16267), .B2(n16266), .A(n16265), .ZN(n17271) );
  AND2_X1 U11908 ( .A1(n12906), .A2(n12905), .ZN(n14955) );
  NAND2_X1 U11909 ( .A1(n11511), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11551) );
  NAND2_X1 U11910 ( .A1(n13944), .A2(n13929), .ZN(n20688) );
  OR2_X1 U11911 ( .A1(n13944), .A2(n13952), .ZN(n20683) );
  OR2_X1 U11912 ( .A1(n13579), .A2(n14982), .ZN(n13594) );
  NAND2_X1 U11913 ( .A1(n13928), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13579) );
  AND2_X1 U11914 ( .A1(n12007), .A2(n12006), .ZN(n14682) );
  AND2_X1 U11915 ( .A1(n11554), .A2(n11553), .ZN(n14701) );
  NOR2_X2 U11916 ( .A1(n13272), .A2(n13271), .ZN(n13282) );
  NAND2_X1 U11917 ( .A1(n13072), .A2(n14959), .ZN(n13107) );
  INV_X1 U11918 ( .A(n13576), .ZN(n13073) );
  OR3_X1 U11919 ( .A1(n13173), .A2(n20973), .A3(n14955), .ZN(n13121) );
  INV_X1 U11920 ( .A(n12039), .ZN(n10110) );
  NOR2_X1 U11921 ( .A1(n10115), .A2(n10113), .ZN(n10112) );
  INV_X1 U11922 ( .A(n14370), .ZN(n10115) );
  NAND2_X1 U11923 ( .A1(n14535), .A2(n10112), .ZN(n14372) );
  OR2_X1 U11924 ( .A1(n11809), .A2(n14527), .ZN(n11855) );
  INV_X1 U11925 ( .A(n10113), .ZN(n10111) );
  AND2_X1 U11926 ( .A1(n11760), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11761) );
  AND2_X1 U11927 ( .A1(n11714), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11715) );
  OAI21_X1 U11928 ( .B1(n11319), .B2(n14870), .A(n11737), .ZN(n14578) );
  NAND2_X1 U11929 ( .A1(n11677), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11713) );
  NAND2_X1 U11930 ( .A1(n9716), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9742) );
  AND2_X1 U11931 ( .A1(n11637), .A2(n11636), .ZN(n14680) );
  NOR2_X1 U11932 ( .A1(n10101), .A2(n14689), .ZN(n10100) );
  INV_X1 U11933 ( .A(n10102), .ZN(n10101) );
  NOR2_X1 U11934 ( .A1(n11588), .A2(n14650), .ZN(n11589) );
  NAND2_X1 U11935 ( .A1(n11552), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11588) );
  NOR2_X1 U11936 ( .A1(n11440), .A2(n14946), .ZN(n11441) );
  AND4_X1 U11937 ( .A1(n11404), .A2(n11403), .A3(n11402), .A4(n11401), .ZN(
        n13924) );
  AOI21_X1 U11938 ( .B1(n12106), .B2(n11524), .A(n11387), .ZN(n13912) );
  AOI21_X1 U11939 ( .B1(n12097), .B2(n11524), .A(n11371), .ZN(n13648) );
  NOR2_X1 U11940 ( .A1(n11342), .A2(n11345), .ZN(n11367) );
  INV_X1 U11941 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11345) );
  AND2_X1 U11942 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11291), .ZN(
        n11321) );
  NAND2_X1 U11943 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11292) );
  NAND2_X1 U11944 ( .A1(n13267), .A2(n11270), .ZN(n13278) );
  XNOR2_X1 U11945 ( .A(n12142), .B(n21093), .ZN(n10139) );
  NAND2_X1 U11946 ( .A1(n14850), .A2(n15048), .ZN(n9874) );
  INV_X1 U11947 ( .A(n14537), .ZN(n9976) );
  NAND2_X1 U11948 ( .A1(n14592), .A2(n9699), .ZN(n14551) );
  NAND2_X1 U11949 ( .A1(n14592), .A2(n9978), .ZN(n14569) );
  AND2_X1 U11950 ( .A1(n14592), .A2(n14581), .ZN(n14579) );
  INV_X1 U11951 ( .A(n14865), .ZN(n14875) );
  NOR2_X1 U11952 ( .A1(n14683), .A2(n14682), .ZN(n14684) );
  NAND2_X1 U11953 ( .A1(n14684), .A2(n14618), .ZN(n14617) );
  NAND2_X1 U11954 ( .A1(n9741), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14891) );
  INV_X1 U11955 ( .A(n14913), .ZN(n9741) );
  NAND2_X1 U11956 ( .A1(n9869), .A2(n9872), .ZN(n14890) );
  NAND2_X1 U11957 ( .A1(n9975), .A2(n9974), .ZN(n14683) );
  INV_X1 U11958 ( .A(n14635), .ZN(n9974) );
  INV_X1 U11959 ( .A(n9975), .ZN(n14694) );
  NAND2_X1 U11960 ( .A1(n14704), .A2(n14645), .ZN(n14692) );
  AND2_X1 U11961 ( .A1(n11979), .A2(n11978), .ZN(n14033) );
  NAND2_X1 U11962 ( .A1(n14134), .A2(n12121), .ZN(n14151) );
  NAND2_X1 U11963 ( .A1(n14151), .A2(n14150), .ZN(n16675) );
  AND2_X1 U11964 ( .A1(n11974), .A2(n11973), .ZN(n13936) );
  INV_X1 U11965 ( .A(n9984), .ZN(n13981) );
  NAND2_X1 U11966 ( .A1(n10125), .A2(n10126), .ZN(n16685) );
  INV_X1 U11967 ( .A(n12096), .ZN(n10127) );
  NOR2_X1 U11968 ( .A1(n16831), .A2(n13649), .ZN(n13917) );
  NAND2_X1 U11969 ( .A1(n9973), .A2(n9972), .ZN(n9971) );
  INV_X1 U11970 ( .A(n16830), .ZN(n9972) );
  OAI21_X1 U11971 ( .B1(n20813), .B2(n15151), .A(n16799), .ZN(n16829) );
  OR2_X1 U11972 ( .A1(n20847), .A2(n20839), .ZN(n16800) );
  OR2_X1 U11973 ( .A1(n11182), .A2(n11181), .ZN(n12051) );
  INV_X2 U11974 ( .A(n11935), .ZN(n11929) );
  OR2_X1 U11975 ( .A1(n11224), .A2(n11223), .ZN(n11225) );
  NAND2_X1 U11976 ( .A1(n11274), .A2(n11273), .ZN(n13420) );
  INV_X1 U11977 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13164) );
  NOR2_X1 U11978 ( .A1(n13283), .A2(n12069), .ZN(n13286) );
  NAND2_X1 U11979 ( .A1(n9690), .A2(n9746), .ZN(n13499) );
  NOR2_X1 U11980 ( .A1(n12060), .A2(n15158), .ZN(n13662) );
  INV_X1 U11981 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13870) );
  OR2_X1 U11982 ( .A1(n13538), .A2(n13663), .ZN(n20856) );
  INV_X1 U11983 ( .A(n13452), .ZN(n13535) );
  AND3_X1 U11984 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20963), .A3(n13287), 
        .ZN(n13319) );
  INV_X1 U11985 ( .A(n16848), .ZN(n13181) );
  OR2_X1 U11986 ( .A1(n14410), .A2(n14409), .ZN(n14413) );
  AOI21_X1 U11988 ( .B1(n19753), .B2(n15693), .A(n15377), .ZN(n9933) );
  NAND2_X1 U11989 ( .A1(n10356), .A2(n10355), .ZN(n10778) );
  NAND2_X1 U11990 ( .A1(n16883), .A2(n16877), .ZN(n16871) );
  NOR2_X1 U11991 ( .A1(n15628), .A2(n15627), .ZN(n15626) );
  NOR2_X1 U11992 ( .A1(n16884), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16883) );
  AND2_X1 U11993 ( .A1(n10354), .A2(n10762), .ZN(n10763) );
  NAND2_X1 U11994 ( .A1(n10716), .A2(n9912), .ZN(n10712) );
  AOI21_X1 U11995 ( .B1(n19644), .B2(n19753), .A(n15447), .ZN(n19629) );
  OAI21_X1 U11996 ( .B1(n19643), .B2(n9934), .A(n19642), .ZN(n19644) );
  AOI21_X1 U11997 ( .B1(n19662), .B2(n19753), .A(n10193), .ZN(n19643) );
  OAI21_X1 U11998 ( .B1(n9934), .B2(n19661), .A(n19660), .ZN(n19662) );
  NOR2_X1 U11999 ( .A1(n9916), .A2(n10727), .ZN(n9915) );
  INV_X1 U12000 ( .A(n9917), .ZN(n9916) );
  NAND2_X1 U12001 ( .A1(n10352), .A2(n9917), .ZN(n10733) );
  NAND2_X1 U12002 ( .A1(n10352), .A2(n10702), .ZN(n10731) );
  NAND2_X1 U12003 ( .A1(n9936), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12822) );
  INV_X1 U12004 ( .A(n12820), .ZN(n9936) );
  NAND2_X1 U12005 ( .A1(n9937), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12820) );
  INV_X1 U12006 ( .A(n12818), .ZN(n9937) );
  AND2_X1 U12007 ( .A1(n10691), .A2(n10690), .ZN(n19682) );
  AND2_X1 U12008 ( .A1(n9905), .A2(n9908), .ZN(n10674) );
  NOR2_X1 U12009 ( .A1(n10631), .A2(n9906), .ZN(n9905) );
  INV_X1 U12010 ( .A(n10639), .ZN(n9906) );
  NAND2_X1 U12011 ( .A1(n10638), .A2(n10639), .ZN(n10627) );
  NAND3_X1 U12012 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12805) );
  AND2_X1 U12013 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12804) );
  NOR3_X1 U12014 ( .A1(n15558), .A2(n15546), .A3(n10092), .ZN(n15540) );
  NOR2_X1 U12015 ( .A1(n15558), .A2(n15546), .ZN(n15548) );
  NAND2_X1 U12016 ( .A1(n15496), .A2(n9636), .ZN(n15583) );
  AOI21_X1 U12017 ( .B1(n15526), .B2(n9801), .A(n12594), .ZN(n9799) );
  NOR2_X1 U12018 ( .A1(n9804), .A2(n12590), .ZN(n9801) );
  NAND2_X1 U12019 ( .A1(n9655), .A2(n9802), .ZN(n9800) );
  NOR2_X1 U12020 ( .A1(n9804), .A2(n9803), .ZN(n9802) );
  INV_X1 U12021 ( .A(n9807), .ZN(n9803) );
  NAND2_X1 U12022 ( .A1(n9806), .A2(n9805), .ZN(n15521) );
  INV_X1 U12023 ( .A(n15609), .ZN(n10160) );
  NAND2_X1 U12024 ( .A1(n15535), .A2(n15537), .ZN(n15536) );
  XNOR2_X1 U12025 ( .A(n12493), .B(n12489), .ZN(n15543) );
  INV_X1 U12026 ( .A(n15567), .ZN(n10188) );
  AND2_X1 U12027 ( .A1(n12727), .A2(n12726), .ZN(n15650) );
  NOR2_X1 U12028 ( .A1(n15651), .A2(n15650), .ZN(n15652) );
  NAND2_X1 U12029 ( .A1(n10181), .A2(n9798), .ZN(n9797) );
  INV_X1 U12030 ( .A(n9697), .ZN(n9798) );
  AND2_X1 U12031 ( .A1(n12313), .A2(n10182), .ZN(n10181) );
  AND2_X1 U12032 ( .A1(n12700), .A2(n12699), .ZN(n16988) );
  AND2_X1 U12033 ( .A1(n12975), .A2(n20503), .ZN(n19869) );
  INV_X1 U12034 ( .A(n12759), .ZN(n13860) );
  NAND2_X1 U12035 ( .A1(n15335), .A2(n9646), .ZN(n15337) );
  AND2_X1 U12036 ( .A1(n15320), .A2(n9943), .ZN(n15329) );
  AND2_X1 U12037 ( .A1(n9635), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9943) );
  NAND2_X1 U12038 ( .A1(n15320), .A2(n9635), .ZN(n15326) );
  NAND2_X1 U12039 ( .A1(n15320), .A2(n9944), .ZN(n15324) );
  NAND2_X1 U12040 ( .A1(n15320), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15322) );
  AND2_X1 U12041 ( .A1(n15310), .A2(n9643), .ZN(n15318) );
  NAND2_X1 U12042 ( .A1(n15310), .A2(n9621), .ZN(n15316) );
  OR2_X1 U12043 ( .A1(n15466), .A2(n15576), .ZN(n15578) );
  NAND2_X1 U12044 ( .A1(n15310), .A2(n9633), .ZN(n15314) );
  INV_X1 U12045 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19655) );
  INV_X1 U12046 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15843) );
  NOR2_X1 U12047 ( .A1(n12822), .A2(n15865), .ZN(n12823) );
  INV_X1 U12048 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15865) );
  NAND2_X1 U12049 ( .A1(n12816), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12818) );
  NAND2_X1 U12050 ( .A1(n13189), .A2(n10097), .ZN(n14050) );
  NOR2_X1 U12051 ( .A1(n12810), .A2(n9939), .ZN(n12816) );
  NAND2_X1 U12052 ( .A1(n9940), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9939) );
  INV_X1 U12053 ( .A(n9942), .ZN(n9940) );
  NOR2_X1 U12054 ( .A1(n12810), .A2(n9942), .ZN(n12814) );
  AND2_X1 U12055 ( .A1(n13189), .A2(n13243), .ZN(n14052) );
  NAND2_X1 U12056 ( .A1(n9941), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12812) );
  INV_X1 U12057 ( .A(n12810), .ZN(n9941) );
  AND2_X1 U12058 ( .A1(n10860), .A2(n10859), .ZN(n13102) );
  NOR2_X1 U12059 ( .A1(n13101), .A2(n13102), .ZN(n13191) );
  NOR2_X1 U12060 ( .A1(n12805), .A2(n14004), .ZN(n12807) );
  NAND2_X1 U12061 ( .A1(n12807), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12810) );
  INV_X1 U12062 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14004) );
  AOI21_X1 U12063 ( .B1(n10849), .B2(n10854), .A(n10853), .ZN(n14001) );
  NAND2_X1 U12064 ( .A1(n15677), .A2(n15970), .ZN(n10055) );
  INV_X1 U12065 ( .A(n15665), .ZN(n9774) );
  OR2_X1 U12066 ( .A1(n9653), .A2(n10931), .ZN(n14421) );
  NAND2_X1 U12067 ( .A1(n15679), .A2(n9626), .ZN(n9776) );
  XNOR2_X1 U12068 ( .A(n15676), .B(n15675), .ZN(n15689) );
  NAND2_X1 U12069 ( .A1(n10844), .A2(n10003), .ZN(n15713) );
  NAND2_X1 U12070 ( .A1(n10844), .A2(n10843), .ZN(n15726) );
  NAND2_X1 U12071 ( .A1(n15569), .A2(n10086), .ZN(n15736) );
  NOR2_X1 U12072 ( .A1(n15651), .A2(n10165), .ZN(n16039) );
  NOR2_X1 U12073 ( .A1(n15651), .A2(n10167), .ZN(n15439) );
  AND2_X1 U12074 ( .A1(n15787), .A2(n15775), .ZN(n15762) );
  AND2_X1 U12075 ( .A1(n16055), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10006) );
  AND2_X1 U12076 ( .A1(n12724), .A2(n12723), .ZN(n15452) );
  AND2_X1 U12077 ( .A1(n16171), .A2(n16055), .ZN(n15790) );
  INV_X1 U12078 ( .A(n15582), .ZN(n10079) );
  AND2_X1 U12079 ( .A1(n12722), .A2(n12721), .ZN(n15470) );
  OR2_X1 U12080 ( .A1(n15480), .A2(n10154), .ZN(n16962) );
  OR3_X1 U12081 ( .A1(n10754), .A2(n10362), .A3(n16968), .ZN(n15825) );
  NAND2_X1 U12082 ( .A1(n9895), .A2(n9893), .ZN(n15827) );
  AND2_X1 U12083 ( .A1(n9894), .A2(n15837), .ZN(n9893) );
  AND2_X1 U12084 ( .A1(n12716), .A2(n12715), .ZN(n15481) );
  NOR2_X1 U12085 ( .A1(n15480), .A2(n15481), .ZN(n16963) );
  NAND2_X1 U12086 ( .A1(n15496), .A2(n15497), .ZN(n15495) );
  AND2_X1 U12087 ( .A1(n10878), .A2(n10877), .ZN(n13564) );
  NOR2_X1 U12088 ( .A1(n15886), .A2(n13564), .ZN(n15496) );
  NAND2_X1 U12089 ( .A1(n13189), .A2(n10093), .ZN(n15886) );
  NOR2_X1 U12090 ( .A1(n10094), .A2(n9714), .ZN(n10093) );
  INV_X1 U12091 ( .A(n10095), .ZN(n10094) );
  AND2_X1 U12092 ( .A1(n13189), .A2(n10095), .ZN(n15884) );
  NAND2_X1 U12093 ( .A1(n10687), .A2(n10683), .ZN(n9878) );
  NAND2_X1 U12094 ( .A1(n9762), .A2(n16189), .ZN(n9767) );
  INV_X1 U12095 ( .A(n9766), .ZN(n9762) );
  NOR2_X1 U12096 ( .A1(n15912), .A2(n10835), .ZN(n10018) );
  INV_X1 U12097 ( .A(n15912), .ZN(n10017) );
  AND2_X1 U12098 ( .A1(n12694), .A2(n12693), .ZN(n14056) );
  NOR3_X1 U12099 ( .A1(n10158), .A2(n14056), .A3(n10157), .ZN(n16163) );
  INV_X1 U12100 ( .A(n16178), .ZN(n10157) );
  INV_X1 U12101 ( .A(n16179), .ZN(n10158) );
  NAND2_X1 U12102 ( .A1(n16179), .A2(n16178), .ZN(n16177) );
  AND2_X1 U12103 ( .A1(n12681), .A2(n12680), .ZN(n19740) );
  NAND2_X1 U12104 ( .A1(n13744), .A2(n13743), .ZN(n19739) );
  NAND2_X1 U12105 ( .A1(n12770), .A2(n10465), .ZN(n14484) );
  XNOR2_X1 U12106 ( .A(n12660), .B(n13011), .ZN(n13372) );
  NOR2_X1 U12107 ( .A1(n9796), .A2(n13061), .ZN(n12170) );
  INV_X1 U12108 ( .A(n13059), .ZN(n9796) );
  NAND2_X1 U12109 ( .A1(n10849), .A2(n10512), .ZN(n10520) );
  INV_X1 U12110 ( .A(n20585), .ZN(n20578) );
  OR2_X1 U12111 ( .A1(n20138), .A2(n20137), .ZN(n20146) );
  NOR2_X2 U12112 ( .A1(n13860), .A2(n13859), .ZN(n19965) );
  NOR2_X2 U12113 ( .A1(n13858), .A2(n13859), .ZN(n19966) );
  NAND2_X1 U12114 ( .A1(n10029), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10023) );
  NAND2_X1 U12115 ( .A1(n10037), .A2(n10416), .ZN(n10024) );
  NAND2_X1 U12116 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20425), .ZN(n19961) );
  INV_X1 U12117 ( .A(n19961), .ZN(n19951) );
  NAND2_X1 U12118 ( .A1(n20582), .A2(n16222), .ZN(n20361) );
  NAND2_X1 U12119 ( .A1(n20582), .A2(n20609), .ZN(n20390) );
  NOR2_X1 U12120 ( .A1(n18930), .A2(n16283), .ZN(n16290) );
  OR2_X1 U12121 ( .A1(n17407), .A2(n9948), .ZN(n9946) );
  OR2_X1 U12122 ( .A1(n18304), .A2(n18313), .ZN(n9948) );
  OR2_X1 U12123 ( .A1(n17407), .A2(n18313), .ZN(n9949) );
  NOR2_X1 U12124 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17502), .ZN(n17486) );
  NOR2_X1 U12125 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17529), .ZN(n17517) );
  INV_X1 U12126 ( .A(n19394), .ZN(n19372) );
  NAND2_X1 U12127 ( .A1(n19414), .A2(n17292), .ZN(n17656) );
  AOI211_X1 U12128 ( .C1(n17816), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n16340), .B(n16339), .ZN(n16341) );
  NOR2_X1 U12129 ( .A1(n18101), .A2(n18100), .ZN(n18119) );
  NOR2_X1 U12130 ( .A1(n17271), .A2(n19413), .ZN(n18140) );
  NAND2_X1 U12131 ( .A1(n17133), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17102) );
  OR2_X1 U12132 ( .A1(n16414), .A2(n9987), .ZN(n9985) );
  AND2_X1 U12133 ( .A1(n18496), .A2(n9988), .ZN(n9987) );
  AND2_X1 U12134 ( .A1(n18300), .A2(n9694), .ZN(n18212) );
  NOR2_X1 U12135 ( .A1(n18336), .A2(n17303), .ZN(n18300) );
  NAND2_X1 U12136 ( .A1(n18327), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18336) );
  NOR2_X1 U12137 ( .A1(n18376), .A2(n18381), .ZN(n18327) );
  NAND3_X1 U12138 ( .A1(n9954), .A2(n9625), .A3(n9672), .ZN(n18419) );
  AND2_X1 U12139 ( .A1(n9954), .A2(n9625), .ZN(n18449) );
  NOR2_X1 U12140 ( .A1(n18494), .A2(n18819), .ZN(n17113) );
  NOR2_X1 U12141 ( .A1(n18520), .A2(n9956), .ZN(n9955) );
  NOR2_X1 U12142 ( .A1(n18517), .A2(n18520), .ZN(n18488) );
  AOI22_X1 U12143 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14264) );
  AOI22_X1 U12144 ( .A1(n16346), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14265) );
  NOR2_X1 U12145 ( .A1(n18228), .A2(n17154), .ZN(n16543) );
  AOI21_X1 U12146 ( .B1(n17162), .B2(n18753), .A(n17161), .ZN(n10013) );
  INV_X1 U12147 ( .A(n18403), .ZN(n9759) );
  NOR2_X1 U12148 ( .A1(n18459), .A2(n10002), .ZN(n16407) );
  NOR2_X1 U12149 ( .A1(n18779), .A2(n18708), .ZN(n18412) );
  OAI21_X1 U12150 ( .B1(n19368), .B2(n16439), .A(n19367), .ZN(n19380) );
  INV_X1 U12151 ( .A(n17113), .ZN(n18779) );
  NAND2_X1 U12152 ( .A1(n16471), .A2(n18483), .ZN(n18782) );
  NAND2_X1 U12153 ( .A1(n18926), .A2(n18710), .ZN(n19360) );
  NAND2_X1 U12154 ( .A1(n16465), .A2(n18512), .ZN(n18506) );
  XOR2_X1 U12155 ( .A(n16404), .B(n16403), .Z(n18502) );
  NAND2_X1 U12156 ( .A1(n18502), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18501) );
  XNOR2_X1 U12157 ( .A(n16381), .B(n9990), .ZN(n18566) );
  NAND2_X1 U12158 ( .A1(n18565), .A2(n18566), .ZN(n18564) );
  NAND2_X1 U12159 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19391) );
  NAND2_X1 U12160 ( .A1(n16284), .A2(n16440), .ZN(n19357) );
  INV_X1 U12161 ( .A(n19574), .ZN(n18926) );
  NOR2_X1 U12162 ( .A1(n14189), .A2(n14188), .ZN(n18934) );
  NOR2_X1 U12163 ( .A1(n14242), .A2(n14241), .ZN(n18938) );
  NOR2_X1 U12164 ( .A1(n14211), .A2(n14210), .ZN(n18942) );
  INV_X1 U12165 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19385) );
  NAND2_X1 U12166 ( .A1(n19577), .A2(n18921), .ZN(n19002) );
  NOR2_X1 U12167 ( .A1(n19574), .A2(n16285), .ZN(n19415) );
  NAND2_X1 U12168 ( .A1(n19424), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19413) );
  INV_X1 U12169 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14650) );
  INV_X1 U12170 ( .A(n20705), .ZN(n16596) );
  INV_X1 U12171 ( .A(n20702), .ZN(n20660) );
  AND2_X1 U12172 ( .A1(n13928), .A2(n13585), .ZN(n20687) );
  AND2_X1 U12173 ( .A1(n13928), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20705) );
  INV_X1 U12174 ( .A(n20683), .ZN(n16587) );
  CLKBUF_X1 U12175 ( .A(n14731), .Z(n14699) );
  INV_X1 U12176 ( .A(n14730), .ZN(n20717) );
  INV_X1 U12177 ( .A(n20721), .ZN(n14715) );
  AND2_X2 U12178 ( .A1(n11947), .A2(n14967), .ZN(n20721) );
  NAND2_X1 U12179 ( .A1(n20721), .A2(n14403), .ZN(n14730) );
  INV_X1 U12180 ( .A(n16652), .ZN(n14791) );
  NOR2_X2 U12181 ( .A1(n16647), .A2(n13081), .ZN(n14804) );
  INV_X1 U12182 ( .A(n16645), .ZN(n14802) );
  AND2_X1 U12183 ( .A1(n13041), .A2(n14953), .ZN(n20724) );
  OAI21_X1 U12184 ( .B1(n14913), .B2(n9742), .A(n16656), .ZN(n14883) );
  INV_X1 U12185 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14946) );
  INV_X1 U12186 ( .A(n16695), .ZN(n16669) );
  NOR2_X1 U12187 ( .A1(n16520), .A2(n20633), .ZN(n12145) );
  NAND2_X1 U12188 ( .A1(n11250), .A2(n11270), .ZN(n13270) );
  NAND2_X1 U12189 ( .A1(n12043), .A2(n13770), .ZN(n21063) );
  NAND2_X1 U12190 ( .A1(n14818), .A2(n10139), .ZN(n10138) );
  INV_X1 U12191 ( .A(n10140), .ZN(n9749) );
  XNOR2_X1 U12192 ( .A(n14829), .B(n14828), .ZN(n15045) );
  OAI21_X1 U12193 ( .B1(n9673), .B2(n15123), .A(n9873), .ZN(n14829) );
  OAI21_X1 U12194 ( .B1(n14827), .B2(n9719), .A(n15123), .ZN(n9873) );
  AND2_X1 U12195 ( .A1(n15076), .A2(n15005), .ZN(n16730) );
  INV_X1 U12196 ( .A(n16829), .ZN(n16778) );
  NAND2_X1 U12197 ( .A1(n16691), .A2(n16690), .ZN(n16689) );
  NAND2_X1 U12198 ( .A1(n16696), .A2(n12096), .ZN(n16691) );
  NOR2_X1 U12199 ( .A1(n16778), .A2(n16781), .ZN(n16823) );
  OR2_X1 U12200 ( .A1(n16805), .A2(n16804), .ZN(n16833) );
  AND2_X1 U12201 ( .A1(n14992), .A2(n16508), .ZN(n20838) );
  AND2_X1 U12202 ( .A1(n14992), .A2(n14979), .ZN(n20849) );
  INV_X1 U12203 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20854) );
  NOR2_X1 U12204 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20632) );
  NOR2_X1 U12205 ( .A1(n14963), .A2(n20905), .ZN(n16539) );
  INV_X1 U12206 ( .A(n15199), .ZN(n15234) );
  INV_X1 U12207 ( .A(n13817), .ZN(n13522) );
  OAI21_X1 U12208 ( .B1(n13769), .B2(n13823), .A(n20904), .ZN(n13839) );
  INV_X1 U12209 ( .A(n13781), .ZN(n13843) );
  INV_X1 U12210 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13443) );
  INV_X1 U12211 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13429) );
  INV_X1 U12212 ( .A(n15290), .ZN(n13446) );
  NOR2_X1 U12213 ( .A1(n13418), .A2(n13656), .ZN(n13450) );
  AND2_X1 U12214 ( .A1(n13452), .A2(n13451), .ZN(n20887) );
  AOI22_X1 U12215 ( .A1(n20900), .A2(n20909), .B1(n20899), .B2(n20898), .ZN(
        n20961) );
  NOR2_X1 U12216 ( .A1(n13305), .A2(n13768), .ZN(n13660) );
  NOR2_X1 U12217 ( .A1(n14789), .A2(n13768), .ZN(n13678) );
  NOR2_X1 U12218 ( .A1(n14777), .A2(n13768), .ZN(n13686) );
  NOR2_X1 U12219 ( .A1(n13494), .A2(n13768), .ZN(n13668) );
  NOR2_X1 U12220 ( .A1(n14772), .A2(n13768), .ZN(n13691) );
  INV_X1 U12221 ( .A(n15259), .ZN(n20916) );
  INV_X1 U12222 ( .A(n15264), .ZN(n20922) );
  INV_X1 U12223 ( .A(n15274), .ZN(n20934) );
  INV_X1 U12224 ( .A(n15279), .ZN(n20940) );
  OAI211_X1 U12225 ( .C1(n13872), .C2(n13903), .A(n20865), .B(n20904), .ZN(
        n13896) );
  NOR2_X1 U12226 ( .A1(n13768), .A2(n13697), .ZN(n13905) );
  NOR2_X1 U12227 ( .A1(n13768), .A2(n13914), .ZN(n13898) );
  INV_X1 U12228 ( .A(n13895), .ZN(n13906) );
  INV_X1 U12229 ( .A(n13660), .ZN(n20915) );
  INV_X1 U12230 ( .A(n13678), .ZN(n20921) );
  INV_X1 U12231 ( .A(n13682), .ZN(n20927) );
  INV_X1 U12232 ( .A(n13686), .ZN(n20933) );
  INV_X1 U12233 ( .A(n13691), .ZN(n20945) );
  INV_X1 U12234 ( .A(n15284), .ZN(n20946) );
  INV_X1 U12235 ( .A(n13898), .ZN(n20960) );
  AND2_X1 U12236 ( .A1(n20962), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16537) );
  NOR2_X1 U12237 ( .A1(n9924), .A2(n9923), .ZN(n9922) );
  INV_X1 U12238 ( .A(n9927), .ZN(n9923) );
  OAI21_X1 U12239 ( .B1(n15389), .B2(n9934), .A(n15334), .ZN(n15376) );
  AND2_X1 U12240 ( .A1(n10720), .A2(n10719), .ZN(n19649) );
  AND2_X1 U12241 ( .A1(n19599), .A2(n12835), .ZN(n19734) );
  NAND2_X1 U12242 ( .A1(n10688), .A2(n9921), .ZN(n10699) );
  NAND2_X1 U12243 ( .A1(n19753), .A2(n19757), .ZN(n14128) );
  INV_X1 U12244 ( .A(n19654), .ZN(n19732) );
  OR2_X1 U12245 ( .A1(n14130), .A2(n10180), .ZN(n10179) );
  AND2_X1 U12246 ( .A1(n19692), .A2(n12161), .ZN(n10180) );
  NOR2_X2 U12247 ( .A1(n19753), .A2(n19730), .ZN(n15465) );
  AND2_X1 U12248 ( .A1(n15341), .A2(n17075), .ZN(n19743) );
  INV_X1 U12249 ( .A(n15465), .ZN(n19665) );
  INV_X1 U12250 ( .A(n14128), .ZN(n15517) );
  NOR2_X1 U12251 ( .A1(n13363), .A2(n10183), .ZN(n19774) );
  OR2_X1 U12252 ( .A1(n12243), .A2(n12242), .ZN(n19778) );
  INV_X1 U12253 ( .A(n20599), .ZN(n16223) );
  INV_X1 U12254 ( .A(n19793), .ZN(n19788) );
  NAND2_X1 U12255 ( .A1(n9655), .A2(n15532), .ZN(n15531) );
  NAND2_X1 U12256 ( .A1(n9808), .A2(n9809), .ZN(n15551) );
  AND2_X1 U12257 ( .A1(n19834), .A2(n12762), .ZN(n19802) );
  NOR2_X1 U12258 ( .A1(n19848), .A2(n19859), .ZN(n19844) );
  NAND2_X1 U12259 ( .A1(n15640), .A2(n13007), .ZN(n19836) );
  AND2_X1 U12260 ( .A1(n19834), .A2(n12748), .ZN(n19859) );
  INV_X1 U12261 ( .A(n19836), .ZN(n19867) );
  NOR2_X1 U12264 ( .A1(n15341), .A2(n12882), .ZN(n12913) );
  XNOR2_X1 U12265 ( .A(n12825), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14430) );
  XNOR2_X1 U12266 ( .A(n14421), .B(n14420), .ZN(n15937) );
  OAI21_X1 U12267 ( .B1(n15375), .B2(n15374), .A(n9653), .ZN(n15969) );
  INV_X1 U12268 ( .A(n16942), .ZN(n16952) );
  AND2_X1 U12269 ( .A1(n16950), .A2(n15929), .ZN(n16942) );
  AND2_X1 U12270 ( .A1(n10845), .A2(n17076), .ZN(n15933) );
  AOI21_X1 U12271 ( .B1(n10775), .B2(n10350), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10060) );
  OR2_X1 U12272 ( .A1(n14457), .A2(n16021), .ZN(n16007) );
  OR2_X1 U12273 ( .A1(n16149), .A2(n14472), .ZN(n16026) );
  INV_X1 U12274 ( .A(n10770), .ZN(n10064) );
  NAND2_X1 U12275 ( .A1(n10761), .A2(n9789), .ZN(n9783) );
  AOI21_X1 U12276 ( .B1(n9882), .B2(n9885), .A(n15750), .ZN(n9879) );
  NAND2_X1 U12277 ( .A1(n16171), .A2(n10006), .ZN(n16090) );
  NAND2_X1 U12278 ( .A1(n15789), .A2(n15786), .ZN(n15774) );
  NAND2_X1 U12279 ( .A1(n9892), .A2(n9897), .ZN(n15839) );
  OR2_X1 U12280 ( .A1(n15863), .A2(n9899), .ZN(n9892) );
  AND2_X1 U12281 ( .A1(n9901), .A2(n15743), .ZN(n15853) );
  AND2_X1 U12282 ( .A1(n10073), .A2(n10074), .ZN(n16144) );
  NAND2_X1 U12283 ( .A1(n16189), .A2(n10051), .ZN(n15892) );
  NAND2_X1 U12284 ( .A1(n16189), .A2(n10677), .ZN(n15908) );
  NAND2_X1 U12285 ( .A1(n10046), .A2(n10048), .ZN(n13997) );
  OR2_X1 U12286 ( .A1(n19930), .A2(n9704), .ZN(n10178) );
  AND2_X1 U12287 ( .A1(n13750), .A2(n17051), .ZN(n19932) );
  INV_X1 U12288 ( .A(n19928), .ZN(n19909) );
  INV_X1 U12289 ( .A(n19911), .ZN(n19931) );
  OR2_X1 U12290 ( .A1(n13754), .A2(n19932), .ZN(n16497) );
  NAND2_X1 U12291 ( .A1(n10497), .A2(n9821), .ZN(n9814) );
  INV_X1 U12292 ( .A(n16222), .ZN(n20609) );
  INV_X1 U12293 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20588) );
  OAI21_X1 U12294 ( .B1(n9822), .B2(n9818), .A(n9815), .ZN(n9817) );
  AOI21_X1 U12295 ( .B1(n10470), .B2(n9628), .A(n9816), .ZN(n9815) );
  AND2_X1 U12296 ( .A1(n10177), .A2(n10176), .ZN(n17042) );
  INV_X1 U12297 ( .A(n14495), .ZN(n10176) );
  NAND2_X1 U12298 ( .A1(n12161), .A2(n17032), .ZN(n10177) );
  INV_X1 U12299 ( .A(n17055), .ZN(n10953) );
  INV_X1 U12300 ( .A(n20582), .ZN(n20570) );
  INV_X1 U12301 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17060) );
  NOR2_X2 U12302 ( .A1(n20222), .A2(n20108), .ZN(n19995) );
  NOR2_X1 U12303 ( .A1(n20147), .A2(n20576), .ZN(n20071) );
  OAI21_X1 U12304 ( .B1(n20086), .B2(n20085), .A(n20084), .ZN(n20103) );
  OAI21_X1 U12305 ( .B1(n20112), .B2(n20128), .A(n20425), .ZN(n20130) );
  INV_X1 U12306 ( .A(n20251), .ZN(n20242) );
  OAI22_X1 U12307 ( .A1(n20231), .A2(n20230), .B1(n20229), .B2(n20491), .ZN(
        n20247) );
  OR2_X1 U12308 ( .A1(n20361), .A2(n20222), .ZN(n20272) );
  INV_X1 U12309 ( .A(n20265), .ZN(n20282) );
  INV_X1 U12310 ( .A(n20272), .ZN(n20281) );
  OAI21_X1 U12311 ( .B1(n20285), .B2(n20262), .A(n20261), .ZN(n20280) );
  NOR2_X1 U12312 ( .A1(n20390), .A2(n20576), .ZN(n20297) );
  NOR2_X1 U12313 ( .A1(n20290), .A2(n20289), .ZN(n20311) );
  NOR2_X2 U12314 ( .A1(n20361), .A2(n20360), .ZN(n20418) );
  INV_X1 U12315 ( .A(n20326), .ZN(n20436) );
  INV_X1 U12316 ( .A(n20332), .ZN(n20447) );
  INV_X1 U12317 ( .A(n20373), .ZN(n20452) );
  INV_X1 U12318 ( .A(n20335), .ZN(n20453) );
  AND2_X1 U12319 ( .A1(n19946), .A2(n19951), .ZN(n20450) );
  AND2_X1 U12320 ( .A1(n19952), .A2(n19951), .ZN(n20457) );
  INV_X1 U12321 ( .A(n20341), .ZN(n20466) );
  INV_X1 U12322 ( .A(n20379), .ZN(n20467) );
  INV_X1 U12323 ( .A(n20382), .ZN(n20473) );
  INV_X1 U12324 ( .A(n20351), .ZN(n20480) );
  INV_X1 U12325 ( .A(n20388), .ZN(n20482) );
  NOR2_X2 U12326 ( .A1(n20390), .A2(n20429), .ZN(n20483) );
  NOR2_X1 U12327 ( .A1(n17079), .A2(n17080), .ZN(n20490) );
  INV_X1 U12328 ( .A(n18140), .ZN(n18101) );
  INV_X1 U12329 ( .A(n9970), .ZN(n17326) );
  NOR2_X1 U12330 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17600), .ZN(n17587) );
  AND4_X1 U12331 ( .A1(n21087), .A2(n19577), .A3(n19587), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n17651) );
  INV_X1 U12332 ( .A(n17635), .ZN(n17662) );
  NOR4_X1 U12333 ( .A1(n14268), .A2(n17674), .A3(n17732), .A4(n14267), .ZN(
        n17670) );
  NOR3_X1 U12334 ( .A1(n17503), .A2(n17842), .A3(n17857), .ZN(n17829) );
  NAND2_X1 U12335 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17874), .ZN(n17857) );
  INV_X1 U12336 ( .A(n17961), .ZN(n17954) );
  NOR2_X1 U12337 ( .A1(n18167), .A2(n17971), .ZN(n17967) );
  NOR2_X1 U12338 ( .A1(n18163), .A2(n17980), .ZN(n17975) );
  INV_X1 U12339 ( .A(n17985), .ZN(n17981) );
  NAND2_X1 U12340 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17981), .ZN(n17980) );
  NOR2_X1 U12341 ( .A1(n18087), .A2(n17990), .ZN(n17986) );
  INV_X1 U12342 ( .A(n18004), .ZN(n18000) );
  NOR2_X1 U12343 ( .A1(n18149), .A2(n18013), .ZN(n18008) );
  INV_X1 U12344 ( .A(n18019), .ZN(n18014) );
  INV_X1 U12345 ( .A(n18029), .ZN(n18018) );
  NAND2_X1 U12346 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18030), .ZN(n18026) );
  NOR2_X1 U12347 ( .A1(n18208), .A2(n18035), .ZN(n18030) );
  NOR2_X1 U12348 ( .A1(n16563), .A2(n16562), .ZN(n18049) );
  NOR3_X1 U12349 ( .A1(n18094), .A2(n18066), .A3(n18067), .ZN(n17946) );
  NOR2_X1 U12350 ( .A1(n16332), .A2(n16331), .ZN(n18084) );
  INV_X1 U12351 ( .A(n16445), .ZN(n18088) );
  INV_X1 U12352 ( .A(n16455), .ZN(n18099) );
  INV_X1 U12353 ( .A(n18061), .ZN(n18095) );
  NOR2_X1 U12354 ( .A1(n16393), .A2(n16392), .ZN(n16564) );
  NOR2_X1 U12355 ( .A1(n16562), .A2(n18173), .ZN(n17945) );
  NOR2_X2 U12356 ( .A1(n14231), .A2(n14230), .ZN(n18954) );
  CLKBUF_X1 U12358 ( .A(n18131), .Z(n18137) );
  NOR2_X1 U12359 ( .A1(n18926), .A2(n18204), .ZN(n18196) );
  OAI211_X1 U12360 ( .C1(n18926), .C2(n19568), .A(n18141), .B(n18140), .ZN(
        n18199) );
  BUF_X1 U12361 ( .A(n18199), .Z(n18204) );
  NAND2_X1 U12363 ( .A1(n9961), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9959) );
  OR2_X1 U12364 ( .A1(n17133), .A2(n17317), .ZN(n9958) );
  NAND2_X1 U12365 ( .A1(n18212), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18209) );
  NAND2_X1 U12366 ( .A1(n18300), .A2(n9622), .ZN(n18243) );
  NAND2_X1 U12367 ( .A1(n18300), .A2(n9632), .ZN(n18283) );
  AOI22_X1 U12368 ( .A1(n18498), .A2(n17113), .B1(n18550), .B2(n18782), .ZN(
        n18482) );
  NAND2_X1 U12369 ( .A1(n9954), .A2(n9955), .ZN(n18487) );
  INV_X1 U12370 ( .A(n18429), .ZN(n18498) );
  NAND2_X1 U12371 ( .A1(n18527), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18517) );
  INV_X1 U12372 ( .A(n18950), .ZN(n18949) );
  INV_X1 U12373 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18520) );
  NOR2_X1 U12374 ( .A1(n18545), .A2(n18547), .ZN(n18527) );
  INV_X1 U12375 ( .A(n18949), .ZN(n19302) );
  INV_X1 U12376 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18581) );
  NAND2_X1 U12377 ( .A1(n18364), .A2(n18436), .ZN(n18580) );
  INV_X1 U12378 ( .A(n18550), .ZN(n18591) );
  OAI21_X2 U12379 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19571), .A(n17274), 
        .ZN(n18587) );
  NOR2_X1 U12380 ( .A1(n18902), .A2(n18217), .ZN(n10010) );
  NAND2_X1 U12381 ( .A1(n18888), .A2(n19382), .ZN(n18814) );
  NAND2_X1 U12382 ( .A1(n18324), .A2(n10004), .ZN(n18265) );
  INV_X1 U12383 ( .A(n18814), .ZN(n18710) );
  NAND2_X1 U12384 ( .A1(n18516), .A2(n18515), .ZN(n18514) );
  NAND2_X1 U12385 ( .A1(n10001), .A2(n10000), .ZN(n18516) );
  NAND2_X1 U12386 ( .A1(n18530), .A2(n9624), .ZN(n10001) );
  NAND2_X1 U12387 ( .A1(n18530), .A2(n18529), .ZN(n18528) );
  NOR2_X1 U12388 ( .A1(n19589), .A2(n16433), .ZN(n18879) );
  INV_X1 U12389 ( .A(n18815), .ZN(n18892) );
  NOR2_X1 U12390 ( .A1(n16440), .A2(n16439), .ZN(n19382) );
  INV_X1 U12391 ( .A(n18896), .ZN(n18901) );
  INV_X1 U12392 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17605) );
  INV_X1 U12393 ( .A(n19413), .ZN(n19572) );
  NOR2_X1 U12394 ( .A1(n19577), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n19424) );
  NAND2_X1 U12395 ( .A1(n19448), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19585) );
  AND2_X2 U12396 ( .A1(n12794), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14738)
         );
  CLKBUF_X1 U12397 ( .A(n17252), .Z(n17258) );
  NAND2_X1 U12398 ( .A1(n9731), .A2(n9728), .ZN(P1_U2810) );
  NAND2_X1 U12399 ( .A1(n9981), .A2(n20676), .ZN(n9731) );
  INV_X1 U12400 ( .A(n14521), .ZN(n9729) );
  NAND2_X1 U12401 ( .A1(n14838), .A2(n10135), .ZN(n10128) );
  AND2_X1 U12402 ( .A1(n12767), .A2(n12766), .ZN(n12768) );
  NOR2_X1 U12403 ( .A1(n10965), .A2(n10964), .ZN(n10966) );
  INV_X1 U12404 ( .A(n10963), .ZN(n10964) );
  AOI21_X1 U12405 ( .B1(n14475), .B2(n17013), .A(n14474), .ZN(n14476) );
  OAI21_X1 U12406 ( .B1(n16899), .B2(n19911), .A(n10075), .ZN(n14474) );
  AND2_X1 U12407 ( .A1(n14473), .A2(n10192), .ZN(n10075) );
  AND2_X1 U12408 ( .A1(n9965), .A2(n9966), .ZN(n17315) );
  AOI21_X1 U12409 ( .B1(n17121), .B2(n18497), .A(n9755), .ZN(n17123) );
  AOI21_X1 U12410 ( .B1(n10011), .B2(n10010), .A(n10007), .ZN(n17164) );
  NOR2_X1 U12411 ( .A1(n14169), .A2(n14166), .ZN(n14284) );
  AND2_X1 U12412 ( .A1(n12607), .A2(n10416), .ZN(n10560) );
  NAND2_X1 U12413 ( .A1(n14797), .A2(n10105), .ZN(n14642) );
  AND2_X1 U12414 ( .A1(n9633), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9621) );
  AND2_X1 U12415 ( .A1(n9637), .A2(n9950), .ZN(n9622) );
  NAND3_X2 U12416 ( .A1(n9958), .A2(n9957), .A3(n9959), .ZN(n17655) );
  INV_X1 U12417 ( .A(n16368), .ZN(n14192) );
  NOR2_X1 U12418 ( .A1(n14167), .A2(n14169), .ZN(n14190) );
  NAND2_X1 U12419 ( .A1(n10116), .A2(n10119), .ZN(n14577) );
  NAND2_X1 U12420 ( .A1(n9732), .A2(n11372), .ZN(n13646) );
  BUF_X1 U12421 ( .A(n11006), .Z(n11842) );
  AND2_X1 U12422 ( .A1(n10440), .A2(n10451), .ZN(n9623) );
  INV_X1 U12423 ( .A(n10515), .ZN(n10849) );
  OR2_X1 U12424 ( .A1(n18529), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9624) );
  AND2_X1 U12425 ( .A1(n9955), .A2(n9953), .ZN(n9625) );
  NAND2_X1 U12426 ( .A1(n10376), .A2(n10375), .ZN(n10406) );
  AND2_X1 U12427 ( .A1(n15674), .A2(n15954), .ZN(n9626) );
  OR2_X1 U12428 ( .A1(n10770), .A2(n9703), .ZN(n9627) );
  INV_X1 U12429 ( .A(n10614), .ZN(n10665) );
  AND2_X1 U12430 ( .A1(n10469), .A2(n9819), .ZN(n9628) );
  AND2_X1 U12431 ( .A1(n12122), .A2(n12121), .ZN(n9629) );
  AND2_X1 U12432 ( .A1(n10004), .A2(n9754), .ZN(n9630) );
  NAND2_X1 U12433 ( .A1(n9753), .A2(n9752), .ZN(n9989) );
  INV_X1 U12434 ( .A(n9989), .ZN(n9751) );
  NAND2_X1 U12435 ( .A1(n10161), .A2(n9700), .ZN(n15608) );
  AND2_X1 U12436 ( .A1(n9970), .A2(n17655), .ZN(n9631) );
  NAND4_X2 U12437 ( .A1(n10347), .A2(n9668), .A3(n10346), .A4(n10345), .ZN(
        n10350) );
  NAND2_X1 U12438 ( .A1(n10188), .A2(n10189), .ZN(n15562) );
  OR2_X1 U12439 ( .A1(n15874), .A2(n16161), .ZN(n10698) );
  AND2_X1 U12440 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9632) );
  AND2_X1 U12441 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9633) );
  AND2_X1 U12442 ( .A1(n15496), .A2(n9693), .ZN(n15467) );
  NOR2_X1 U12443 ( .A1(n9877), .A2(n16160), .ZN(n9634) );
  AND2_X1 U12444 ( .A1(n9944), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9635) );
  AND2_X1 U12445 ( .A1(n10080), .A2(n15482), .ZN(n9636) );
  AND2_X1 U12446 ( .A1(n9632), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9637) );
  NAND2_X1 U12447 ( .A1(n19786), .A2(n19785), .ZN(n9638) );
  OR2_X1 U12448 ( .A1(n13722), .A2(n10049), .ZN(n9639) );
  AND2_X1 U12449 ( .A1(n10086), .A2(n10085), .ZN(n9640) );
  AND2_X1 U12450 ( .A1(n9910), .A2(n15564), .ZN(n9641) );
  AND2_X1 U12451 ( .A1(n9960), .A2(n17317), .ZN(n9642) );
  AND2_X1 U12452 ( .A1(n9621), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9643) );
  OR2_X1 U12453 ( .A1(n10687), .A2(n10683), .ZN(n9644) );
  INV_X2 U12454 ( .A(n19784), .ZN(n19796) );
  OR3_X1 U12455 ( .A1(n17619), .A2(n17319), .A3(n19428), .ZN(n9645) );
  AND2_X1 U12456 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9646) );
  AND2_X1 U12457 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13140) );
  AND2_X1 U12458 ( .A1(n10006), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9647) );
  AND2_X1 U12459 ( .A1(n9717), .A2(n9872), .ZN(n9648) );
  AND2_X1 U12460 ( .A1(n10003), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9649) );
  AND2_X1 U12461 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U12462 ( .A1(n16675), .A2(n12122), .ZN(n14921) );
  AND2_X2 U12463 ( .A1(n11117), .A2(n13288), .ZN(n11143) );
  NOR2_X1 U12464 ( .A1(n16911), .A2(n9823), .ZN(n9651) );
  OR2_X1 U12465 ( .A1(n14617), .A2(n14605), .ZN(n9652) );
  OR2_X1 U12466 ( .A1(n15558), .A2(n10088), .ZN(n9653) );
  INV_X1 U12467 ( .A(n14708), .ZN(n10104) );
  AND2_X1 U12468 ( .A1(n10974), .A2(n10981), .ZN(n11160) );
  INV_X4 U12469 ( .A(n14354), .ZN(n17883) );
  AND2_X1 U12470 ( .A1(n10169), .A2(n9793), .ZN(n9655) );
  AND2_X1 U12471 ( .A1(n10067), .A2(n10059), .ZN(n15698) );
  AND2_X1 U12472 ( .A1(n11255), .A2(n11116), .ZN(n11125) );
  NOR2_X1 U12473 ( .A1(n14614), .A2(n14616), .ZN(n14602) );
  NOR2_X1 U12474 ( .A1(n14614), .A2(n10121), .ZN(n14588) );
  NAND2_X1 U12475 ( .A1(n15521), .A2(n15520), .ZN(n15522) );
  INV_X1 U12476 ( .A(n14232), .ZN(n17790) );
  OAI21_X1 U12477 ( .B1(n15389), .B2(n9934), .A(n9933), .ZN(n9931) );
  AND2_X1 U12478 ( .A1(n10146), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9656) );
  NAND2_X1 U12479 ( .A1(n10716), .A2(n9910), .ZN(n9657) );
  NAND2_X1 U12480 ( .A1(n13126), .A2(n13309), .ZN(n9658) );
  INV_X2 U12481 ( .A(n14957), .ZN(n14982) );
  NOR2_X1 U12482 ( .A1(n14708), .A2(n14709), .ZN(n14700) );
  NOR2_X1 U12483 ( .A1(n15453), .A2(n15452), .ZN(n12725) );
  INV_X1 U12484 ( .A(n11135), .ZN(n14973) );
  AND3_X1 U12485 ( .A1(n10159), .A2(n16178), .A3(n16164), .ZN(n9659) );
  AND3_X1 U12486 ( .A1(n15776), .A2(n10760), .A3(n15786), .ZN(n9660) );
  OR3_X1 U12487 ( .A1(n15558), .A2(n10091), .A3(n15546), .ZN(n9661) );
  INV_X1 U12488 ( .A(n9603), .ZN(n11861) );
  AND2_X1 U12489 ( .A1(n10981), .A2(n13156), .ZN(n11056) );
  NAND2_X1 U12490 ( .A1(n9783), .A2(n9787), .ZN(n15721) );
  NAND2_X1 U12491 ( .A1(n9767), .A2(n9876), .ZN(n16159) );
  AND2_X1 U12492 ( .A1(n15379), .A2(n15380), .ZN(n15362) );
  NOR2_X1 U12493 ( .A1(n10783), .A2(n10060), .ZN(n9662) );
  NOR2_X1 U12494 ( .A1(n10761), .A2(n9790), .ZN(n9663) );
  NAND2_X1 U12495 ( .A1(n10352), .A2(n9915), .ZN(n9664) );
  INV_X2 U12496 ( .A(n19936), .ZN(n10451) );
  INV_X1 U12497 ( .A(n19946), .ZN(n10445) );
  AND4_X1 U12498 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n9665) );
  INV_X1 U12499 ( .A(n20111), .ZN(n10664) );
  NAND2_X2 U12500 ( .A1(n11948), .A2(n14957), .ZN(n11959) );
  XNOR2_X1 U12501 ( .A(n12517), .B(n12518), .ZN(n15535) );
  AND2_X1 U12502 ( .A1(n16402), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9666) );
  AND3_X1 U12504 ( .A1(n10131), .A2(n10129), .A3(n10128), .ZN(n9667) );
  AND4_X1 U12505 ( .A1(n10337), .A2(n10336), .A3(n10335), .A4(n10334), .ZN(
        n9668) );
  INV_X1 U12506 ( .A(n12137), .ZN(n10141) );
  OR2_X1 U12507 ( .A1(n11127), .A2(n13309), .ZN(n9669) );
  AND2_X1 U12508 ( .A1(n12520), .A2(n9792), .ZN(n9670) );
  AND2_X1 U12509 ( .A1(n10465), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9671) );
  AND2_X1 U12510 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9672) );
  AND3_X1 U12511 ( .A1(n14827), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9673) );
  INV_X1 U12512 ( .A(n9819), .ZN(n9818) );
  NAND2_X1 U12513 ( .A1(n12156), .A2(n12157), .ZN(n9819) );
  NOR2_X1 U12514 ( .A1(n15611), .A2(n15392), .ZN(n15379) );
  AND2_X1 U12515 ( .A1(n10408), .A2(n10173), .ZN(n9674) );
  NAND2_X1 U12516 ( .A1(n14797), .A2(n10102), .ZN(n10107) );
  AND2_X1 U12517 ( .A1(n10844), .A2(n9649), .ZN(n9675) );
  INV_X1 U12518 ( .A(n9986), .ZN(n18227) );
  NAND2_X1 U12519 ( .A1(n9989), .A2(n9988), .ZN(n9986) );
  AND2_X1 U12520 ( .A1(n12104), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9676) );
  NAND2_X1 U12521 ( .A1(n9881), .A2(n9887), .ZN(n9677) );
  INV_X1 U12522 ( .A(n9773), .ZN(n9772) );
  NAND2_X1 U12523 ( .A1(n9775), .A2(n9774), .ZN(n9773) );
  INV_X1 U12524 ( .A(n10655), .ZN(n10598) );
  NAND2_X1 U12525 ( .A1(n15663), .A2(n15661), .ZN(n9678) );
  INV_X1 U12526 ( .A(n12122), .ZN(n10144) );
  OR2_X1 U12527 ( .A1(n16656), .A2(n16779), .ZN(n12122) );
  OR2_X1 U12528 ( .A1(n15383), .A2(n10362), .ZN(n15679) );
  NAND2_X1 U12529 ( .A1(n15569), .A2(n15435), .ZN(n15419) );
  INV_X1 U12530 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15909) );
  AND2_X1 U12531 ( .A1(n13133), .A2(n11149), .ZN(n9679) );
  NAND3_X1 U12532 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10797) );
  AND2_X1 U12533 ( .A1(n10065), .A2(n10064), .ZN(n9680) );
  AND2_X1 U12534 ( .A1(n10148), .A2(n14021), .ZN(n9681) );
  NOR2_X1 U12535 ( .A1(n17014), .A2(n10498), .ZN(n10548) );
  AND2_X1 U12536 ( .A1(n10138), .A2(n9748), .ZN(n9682) );
  AND2_X1 U12537 ( .A1(n9947), .A2(n17655), .ZN(n9683) );
  NAND2_X1 U12538 ( .A1(n9769), .A2(n19722), .ZN(n10642) );
  OR2_X1 U12539 ( .A1(n10141), .A2(n10144), .ZN(n9684) );
  INV_X1 U12540 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17035) );
  INV_X1 U12541 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14449) );
  INV_X1 U12542 ( .A(n11257), .ZN(n11803) );
  NAND2_X1 U12543 ( .A1(n13134), .A2(n14957), .ZN(n12908) );
  NAND2_X1 U12544 ( .A1(n14727), .A2(n10123), .ZN(n14718) );
  NAND2_X1 U12545 ( .A1(n14727), .A2(n14726), .ZN(n14717) );
  INV_X1 U12546 ( .A(n11835), .ZN(n11278) );
  NAND2_X1 U12547 ( .A1(n10974), .A2(n13140), .ZN(n11835) );
  INV_X1 U12548 ( .A(n11006), .ZN(n11028) );
  AND2_X1 U12549 ( .A1(n15496), .A2(n10080), .ZN(n9685) );
  NAND2_X1 U12550 ( .A1(n13327), .A2(n11211), .ZN(n11217) );
  AND2_X1 U12551 ( .A1(n13922), .A2(n13973), .ZN(n13972) );
  NOR2_X1 U12552 ( .A1(n15493), .A2(n15494), .ZN(n12845) );
  NAND2_X1 U12553 ( .A1(n9925), .A2(n9922), .ZN(n15348) );
  OR3_X1 U12554 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n18292), .ZN(n9686) );
  INV_X1 U12555 ( .A(n15730), .ZN(n9789) );
  AND2_X1 U12556 ( .A1(n15569), .A2(n9640), .ZN(n9687) );
  OR2_X1 U12557 ( .A1(n10070), .A2(n15862), .ZN(n9688) );
  NOR2_X1 U12558 ( .A1(n16911), .A2(n16910), .ZN(n9689) );
  NAND2_X1 U12559 ( .A1(n15543), .A2(n15545), .ZN(n15544) );
  NAND2_X1 U12560 ( .A1(n16191), .A2(n16190), .ZN(n16189) );
  NAND2_X1 U12561 ( .A1(n10152), .A2(n10153), .ZN(n10156) );
  OAI21_X1 U12562 ( .B1(n11929), .B2(n15219), .A(n11315), .ZN(n11325) );
  AND2_X1 U12563 ( .A1(n19598), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12172) );
  INV_X1 U12564 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10099) );
  INV_X1 U12565 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16941) );
  OR2_X1 U12566 ( .A1(n13100), .A2(n9697), .ZN(n13363) );
  INV_X1 U12567 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20963) );
  INV_X1 U12568 ( .A(n9909), .ZN(n10638) );
  OR2_X1 U12569 ( .A1(n10630), .A2(n10631), .ZN(n9909) );
  AND2_X1 U12570 ( .A1(n13498), .A2(n12060), .ZN(n9690) );
  AND2_X1 U12571 ( .A1(n12701), .A2(n19778), .ZN(n9691) );
  AND2_X1 U12572 ( .A1(n10746), .A2(n10745), .ZN(n15750) );
  AND2_X1 U12573 ( .A1(n9915), .A2(n10739), .ZN(n9692) );
  AND2_X1 U12574 ( .A1(n9636), .A2(n10079), .ZN(n9693) );
  AND2_X1 U12575 ( .A1(n9622), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9694) );
  INV_X1 U12576 ( .A(n9877), .ZN(n9876) );
  NAND2_X1 U12577 ( .A1(n9878), .A2(n15905), .ZN(n9877) );
  AND2_X1 U12578 ( .A1(n9813), .A2(n9812), .ZN(n9695) );
  INV_X1 U12579 ( .A(n10698), .ZN(n10074) );
  AND2_X1 U12580 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9696) );
  NAND2_X1 U12581 ( .A1(n12690), .A2(n19785), .ZN(n9697) );
  INV_X1 U12582 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n9990) );
  INV_X1 U12583 ( .A(n15305), .ZN(n9934) );
  INV_X1 U12584 ( .A(n12467), .ZN(n10191) );
  AND2_X1 U12585 ( .A1(n17133), .A2(n9962), .ZN(n9698) );
  AND2_X1 U12586 ( .A1(n13191), .A2(n13190), .ZN(n13189) );
  AND2_X2 U12587 ( .A1(n12605), .A2(n10416), .ZN(n12368) );
  AND2_X2 U12588 ( .A1(n12605), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12351) );
  NAND2_X1 U12589 ( .A1(n12823), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12798) );
  AND2_X1 U12590 ( .A1(n9978), .A2(n9977), .ZN(n9699) );
  AND2_X1 U12591 ( .A1(n10162), .A2(n15618), .ZN(n9700) );
  AND2_X1 U12592 ( .A1(n15310), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15309) );
  AND2_X1 U12593 ( .A1(n10458), .A2(n12861), .ZN(n12770) );
  OR2_X1 U12594 ( .A1(n13100), .A2(n9797), .ZN(n14095) );
  INV_X1 U12595 ( .A(n10702), .ZN(n9918) );
  OR2_X1 U12596 ( .A1(n10362), .A2(n15999), .ZN(n9701) );
  INV_X1 U12597 ( .A(n10717), .ZN(n9914) );
  INV_X1 U12598 ( .A(n15705), .ZN(n10066) );
  INV_X1 U12599 ( .A(n16473), .ZN(n18693) );
  NAND2_X1 U12600 ( .A1(n12467), .A2(n12466), .ZN(n9702) );
  AND2_X1 U12601 ( .A1(n15714), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9703) );
  INV_X1 U12602 ( .A(n9825), .ZN(n9824) );
  NOR2_X1 U12603 ( .A1(n9826), .A2(n16910), .ZN(n9825) );
  INV_X1 U12604 ( .A(n15360), .ZN(n9928) );
  INV_X1 U12605 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15779) );
  INV_X1 U12606 ( .A(n16861), .ZN(n9935) );
  INV_X1 U12607 ( .A(n15538), .ZN(n10092) );
  INV_X1 U12608 ( .A(n9961), .ZN(n9960) );
  NAND2_X1 U12609 ( .A1(n9962), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9961) );
  AND2_X1 U12610 ( .A1(n15335), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10957) );
  AND2_X1 U12611 ( .A1(n19931), .A2(n12161), .ZN(n9704) );
  OR2_X1 U12612 ( .A1(n9645), .A2(n17328), .ZN(n9705) );
  OR2_X1 U12613 ( .A1(n10186), .A2(n12467), .ZN(n9706) );
  NOR2_X1 U12614 ( .A1(n14129), .A2(n10179), .ZN(n9707) );
  NOR2_X1 U12615 ( .A1(n19929), .A2(n10178), .ZN(n9708) );
  INV_X1 U12616 ( .A(n10147), .ZN(n19741) );
  NAND2_X1 U12617 ( .A1(n13744), .A2(n10148), .ZN(n10147) );
  AND2_X1 U12618 ( .A1(n9699), .A2(n9976), .ZN(n9709) );
  INV_X1 U12619 ( .A(n21068), .ZN(n20792) );
  AND2_X1 U12620 ( .A1(n9640), .A2(n15405), .ZN(n9710) );
  AND2_X1 U12621 ( .A1(n9646), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9711) );
  AND2_X1 U12622 ( .A1(n9700), .A2(n10160), .ZN(n9712) );
  INV_X1 U12623 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n9952) );
  INV_X1 U12624 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9951) );
  INV_X1 U12625 ( .A(n18517), .ZN(n9954) );
  INV_X1 U12626 ( .A(n11510), .ZN(n9722) );
  INV_X1 U12627 ( .A(n12841), .ZN(n12880) );
  AND2_X1 U12628 ( .A1(n18300), .A2(n9637), .ZN(n9713) );
  INV_X1 U12629 ( .A(n20696), .ZN(n9973) );
  AND2_X1 U12630 ( .A1(n10875), .A2(n10874), .ZN(n9714) );
  INV_X1 U12631 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10049) );
  INV_X1 U12632 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9964) );
  INV_X1 U12633 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9963) );
  AND2_X1 U12634 ( .A1(n9649), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9715) );
  AND2_X1 U12635 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n9716) );
  AND2_X1 U12636 ( .A1(n15103), .A2(n15110), .ZN(n9717) );
  INV_X1 U12637 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9988) );
  INV_X1 U12638 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9956) );
  INV_X1 U12639 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9837) );
  AND2_X1 U12640 ( .A1(n9994), .A2(n14419), .ZN(n9718) );
  OR2_X1 U12641 ( .A1(n14826), .A2(n9874), .ZN(n9719) );
  INV_X1 U12642 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n9920) );
  INV_X1 U12643 ( .A(n9995), .ZN(n9994) );
  NAND2_X1 U12644 ( .A1(n9650), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9995) );
  NOR2_X1 U12645 ( .A1(n16907), .A2(n10190), .ZN(n10189) );
  NOR2_X1 U12646 ( .A1(n15567), .A2(n16907), .ZN(n15561) );
  CLKBUF_X1 U12647 ( .A(n20768), .Z(n9720) );
  NAND2_X1 U12648 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n9866) );
  NAND2_X1 U12649 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n9863) );
  NAND2_X1 U12650 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n9861) );
  NAND2_X1 U12651 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9859) );
  NAND2_X1 U12652 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U12653 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n9857) );
  NAND2_X1 U12654 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U12655 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U12656 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n9853) );
  NAND2_X1 U12657 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U12658 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U12659 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n9847) );
  NAND3_X1 U12660 ( .A1(n11250), .A2(n9724), .A3(n13064), .ZN(n13267) );
  NOR2_X1 U12661 ( .A1(n11119), .A2(n12965), .ZN(n9727) );
  NOR2_X2 U12662 ( .A1(n9725), .A2(n11119), .ZN(n13134) );
  NAND2_X1 U12663 ( .A1(n9726), .A2(n11123), .ZN(n9725) );
  INV_X1 U12664 ( .A(n12965), .ZN(n9726) );
  NAND2_X1 U12665 ( .A1(n12144), .A2(n9727), .ZN(n13115) );
  NAND3_X1 U12666 ( .A1(n9732), .A2(n11372), .A3(n11388), .ZN(n13911) );
  NAND2_X1 U12667 ( .A1(n10146), .A2(n9696), .ZN(n9736) );
  NAND2_X1 U12668 ( .A1(n9736), .A2(n11149), .ZN(n9735) );
  NAND2_X1 U12669 ( .A1(n11148), .A2(n13133), .ZN(n9734) );
  NAND2_X2 U12670 ( .A1(n11208), .A2(n9733), .ZN(n14445) );
  NAND3_X1 U12671 ( .A1(n9736), .A2(n11148), .A3(n9679), .ZN(n9733) );
  NAND2_X2 U12672 ( .A1(n9735), .A2(n9734), .ZN(n11208) );
  NAND2_X2 U12673 ( .A1(n13164), .A2(n13139), .ZN(n11816) );
  NAND2_X1 U12674 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11002) );
  XNOR2_X2 U12675 ( .A(n13171), .B(n13420), .ZN(n13150) );
  NAND2_X2 U12676 ( .A1(n11224), .A2(n11223), .ZN(n13171) );
  NAND2_X1 U12677 ( .A1(n10142), .A2(n9744), .ZN(n9743) );
  NAND2_X1 U12678 ( .A1(n12069), .A2(n12105), .ZN(n12075) );
  NAND2_X1 U12679 ( .A1(n9750), .A2(n9749), .ZN(n9748) );
  INV_X2 U12680 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19554) );
  INV_X2 U12681 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19531) );
  AND2_X2 U12682 ( .A1(n12623), .A2(n12841), .ZN(n12630) );
  NAND2_X1 U12683 ( .A1(n10441), .A2(n10451), .ZN(n12623) );
  AND2_X4 U12684 ( .A1(n14486), .A2(n14499), .ZN(n10418) );
  NAND2_X1 U12685 ( .A1(n10051), .A2(n9644), .ZN(n9766) );
  NAND2_X1 U12686 ( .A1(n9768), .A2(n10830), .ZN(n9769) );
  NAND2_X2 U12687 ( .A1(n10622), .A2(n10621), .ZN(n10830) );
  AND2_X2 U12688 ( .A1(n10830), .A2(n10625), .ZN(n10822) );
  NAND2_X1 U12689 ( .A1(n15536), .A2(n12520), .ZN(n9794) );
  NAND2_X1 U12690 ( .A1(n9794), .A2(n12545), .ZN(n10169) );
  INV_X1 U12691 ( .A(n13100), .ZN(n19786) );
  NAND2_X1 U12692 ( .A1(n15526), .A2(n15527), .ZN(n9805) );
  NAND2_X1 U12693 ( .A1(n9655), .A2(n9807), .ZN(n9806) );
  NAND2_X1 U12694 ( .A1(n9800), .A2(n9799), .ZN(n12616) );
  INV_X1 U12695 ( .A(n9813), .ZN(n15636) );
  NAND3_X1 U12696 ( .A1(n9821), .A2(n10497), .A3(n12156), .ZN(n9820) );
  NAND3_X1 U12697 ( .A1(n16698), .A2(n16690), .A3(n16697), .ZN(n10125) );
  OAI211_X2 U12698 ( .C1(n9832), .C2(n9830), .A(n9829), .B(n11203), .ZN(n11210) );
  INV_X1 U12699 ( .A(n9831), .ZN(n9830) );
  NAND2_X1 U12700 ( .A1(n11353), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n9834) );
  INV_X1 U12701 ( .A(n9833), .ZN(n11084) );
  INV_X2 U12702 ( .A(n11859), .ZN(n9865) );
  XNOR2_X2 U12703 ( .A(n10830), .B(n10823), .ZN(n10827) );
  NAND2_X1 U12704 ( .A1(n15800), .A2(n15799), .ZN(n9881) );
  NAND2_X1 U12705 ( .A1(n9880), .A2(n9879), .ZN(n15755) );
  NAND2_X1 U12706 ( .A1(n15800), .A2(n9882), .ZN(n9880) );
  NAND2_X1 U12707 ( .A1(n15863), .A2(n9896), .ZN(n9895) );
  NAND3_X1 U12708 ( .A1(n9897), .A2(n9899), .A3(n15838), .ZN(n9894) );
  INV_X1 U12709 ( .A(n9901), .ZN(n15861) );
  NAND2_X1 U12710 ( .A1(n10716), .A2(n9641), .ZN(n10764) );
  AND2_X1 U12711 ( .A1(n10716), .A2(n10717), .ZN(n10708) );
  NAND2_X1 U12712 ( .A1(n10352), .A2(n9692), .ZN(n10724) );
  NAND2_X1 U12713 ( .A1(n10688), .A2(n9919), .ZN(n10703) );
  AOI21_X1 U12714 ( .B1(n16860), .B2(n19753), .A(n16861), .ZN(n15389) );
  NAND2_X1 U12715 ( .A1(n16860), .A2(n9926), .ZN(n9925) );
  NAND2_X1 U12716 ( .A1(n15335), .A2(n9711), .ZN(n12825) );
  INV_X1 U12717 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U12718 ( .A1(n9946), .A2(n9947), .ZN(n17399) );
  INV_X1 U12719 ( .A(n9949), .ZN(n17406) );
  NAND2_X1 U12720 ( .A1(n17133), .A2(n9642), .ZN(n9957) );
  OR2_X1 U12721 ( .A1(n17327), .A2(n9705), .ZN(n9965) );
  OR2_X1 U12722 ( .A1(n17327), .A2(n17328), .ZN(n9970) );
  NAND2_X1 U12723 ( .A1(n13068), .A2(n11953), .ZN(n13272) );
  AND2_X2 U12724 ( .A1(n14592), .A2(n9709), .ZN(n14539) );
  NOR2_X2 U12725 ( .A1(n14032), .A2(n14033), .ZN(n14159) );
  NAND2_X1 U12726 ( .A1(n11133), .A2(n16554), .ZN(n14956) );
  NOR2_X1 U12727 ( .A1(n11133), .A2(n14668), .ZN(n13591) );
  OAI21_X1 U12728 ( .B1(n11133), .B2(n14953), .A(n21051), .ZN(n14954) );
  NAND2_X1 U12729 ( .A1(n11903), .A2(n11133), .ZN(n11913) );
  NOR2_X4 U12730 ( .A1(n14982), .A2(n11133), .ZN(n13066) );
  NAND2_X1 U12731 ( .A1(n14982), .A2(n11133), .ZN(n13576) );
  NAND2_X1 U12732 ( .A1(n13116), .A2(n11133), .ZN(n13173) );
  AND2_X2 U12733 ( .A1(n13223), .A2(n11133), .ZN(n20778) );
  NOR2_X1 U12734 ( .A1(n11133), .A2(n20783), .ZN(n20768) );
  NOR2_X2 U12735 ( .A1(n18241), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18240) );
  OAI22_X1 U12736 ( .A1(n9985), .A2(n18240), .B1(n9988), .B2(n18496), .ZN(
        n18220) );
  AND2_X1 U12737 ( .A1(n15682), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15683) );
  OR2_X1 U12738 ( .A1(n15682), .A2(n14419), .ZN(n9993) );
  NAND2_X1 U12739 ( .A1(n15682), .A2(n9650), .ZN(n15668) );
  NAND3_X1 U12740 ( .A1(n9993), .A2(n9992), .A3(n9991), .ZN(n14475) );
  NAND2_X1 U12741 ( .A1(n18530), .A2(n9996), .ZN(n9997) );
  NAND3_X1 U12742 ( .A1(n18730), .A2(n18465), .A3(n18808), .ZN(n10002) );
  AND2_X2 U12743 ( .A1(n16171), .A2(n9647), .ZN(n15767) );
  NAND2_X2 U12744 ( .A1(n15896), .A2(n10840), .ZN(n16171) );
  NOR2_X2 U12745 ( .A1(n10629), .A2(n10628), .ZN(n10809) );
  NAND4_X1 U12746 ( .A1(n10591), .A2(n10590), .A3(n10588), .A4(n10589), .ZN(
        n10015) );
  NAND4_X1 U12747 ( .A1(n10557), .A2(n10559), .A3(n10556), .A4(n10558), .ZN(
        n10016) );
  INV_X1 U12748 ( .A(n15898), .ZN(n10837) );
  NAND2_X2 U12749 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19394) );
  INV_X1 U12750 ( .A(n10522), .ZN(n10528) );
  NAND2_X1 U12751 ( .A1(n10019), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10523) );
  NAND2_X1 U12752 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10028) );
  INV_X1 U12753 ( .A(n10405), .ZN(n10036) );
  INV_X1 U12754 ( .A(n10404), .ZN(n10044) );
  NAND2_X1 U12755 ( .A1(n10044), .A2(n10416), .ZN(n10021) );
  NAND2_X1 U12756 ( .A1(n10036), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10022) );
  NAND2_X1 U12757 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10026) );
  NAND4_X1 U12758 ( .A1(n10033), .A2(n10032), .A3(n10031), .A4(n10030), .ZN(
        n10029) );
  NAND4_X1 U12759 ( .A1(n10041), .A2(n10040), .A3(n10039), .A4(n10038), .ZN(
        n10037) );
  NAND2_X1 U12760 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10038) );
  NAND2_X1 U12761 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10039) );
  NOR2_X2 U12762 ( .A1(n10052), .A2(n15906), .ZN(n10051) );
  NAND3_X1 U12763 ( .A1(n10059), .A2(n10056), .A3(n10055), .ZN(n10054) );
  NAND2_X1 U12764 ( .A1(n15873), .A2(n15875), .ZN(n10073) );
  NAND3_X1 U12765 ( .A1(n15873), .A2(n10744), .A3(n15875), .ZN(n10069) );
  NAND2_X1 U12766 ( .A1(n15569), .A2(n9710), .ZN(n15556) );
  INV_X1 U12767 ( .A(n13288), .ZN(n11948) );
  OAI21_X1 U12768 ( .B1(n11123), .B2(n13288), .A(n11531), .ZN(n10098) );
  NAND2_X1 U12769 ( .A1(n10104), .A2(n10100), .ZN(n14628) );
  INV_X1 U12770 ( .A(n10107), .ZN(n14643) );
  NAND2_X1 U12771 ( .A1(n14144), .A2(n14143), .ZN(n14146) );
  XNOR2_X2 U12772 ( .A(n14030), .B(n11456), .ZN(n14144) );
  AND2_X1 U12773 ( .A1(n14535), .A2(n10111), .ZN(n14369) );
  NAND2_X1 U12774 ( .A1(n14535), .A2(n14536), .ZN(n14523) );
  NAND2_X1 U12775 ( .A1(n10124), .A2(n11212), .ZN(n12050) );
  NAND3_X1 U12776 ( .A1(n13653), .A2(n11217), .A3(n20963), .ZN(n10124) );
  NAND2_X1 U12777 ( .A1(n14838), .A2(n15038), .ZN(n10133) );
  NAND3_X1 U12778 ( .A1(n10133), .A2(n10132), .A3(n10136), .ZN(n10131) );
  NAND2_X1 U12779 ( .A1(n13744), .A2(n9681), .ZN(n14020) );
  INV_X1 U12780 ( .A(n14020), .ZN(n12686) );
  NAND2_X1 U12781 ( .A1(n10150), .A2(n10377), .ZN(n10430) );
  INV_X1 U12782 ( .A(n10156), .ZN(n14098) );
  NOR2_X2 U12783 ( .A1(n16989), .A2(n16988), .ZN(n14037) );
  NAND2_X1 U12784 ( .A1(n10161), .A2(n9712), .ZN(n15611) );
  INV_X1 U12785 ( .A(n10169), .ZN(n15526) );
  NAND2_X1 U12786 ( .A1(n10170), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10439) );
  NAND3_X1 U12787 ( .A1(n13731), .A2(n10174), .A3(n10171), .ZN(n10170) );
  NAND3_X1 U12788 ( .A1(n10173), .A2(n10408), .A3(n10172), .ZN(n10171) );
  OR2_X1 U12789 ( .A1(n10411), .A2(n10432), .ZN(n10175) );
  INV_X1 U12790 ( .A(n14095), .ZN(n12332) );
  NAND2_X1 U12791 ( .A1(n19787), .A2(n12216), .ZN(n19779) );
  OAI211_X1 U12792 ( .C1(n15567), .C2(n10185), .A(n9706), .B(n10184), .ZN(
        n15638) );
  INV_X1 U12793 ( .A(n10701), .ZN(n10352) );
  NAND2_X1 U12794 ( .A1(n14014), .A2(n14013), .ZN(n14012) );
  OAI21_X1 U12795 ( .B1(n15937), .B2(n19796), .A(n12779), .ZN(n12780) );
  INV_X1 U12796 ( .A(n10822), .ZN(n10821) );
  NOR2_X1 U12797 ( .A1(n19394), .A2(n14172), .ZN(n14168) );
  CLKBUF_X1 U12798 ( .A(n14708), .Z(n14796) );
  AND2_X1 U12799 ( .A1(n15742), .A2(n16141), .ZN(n15863) );
  XNOR2_X1 U12800 ( .A(n10629), .B(n10628), .ZN(n13725) );
  NAND2_X1 U12801 ( .A1(n10680), .A2(n10678), .ZN(n10686) );
  INV_X2 U12802 ( .A(n14332), .ZN(n17877) );
  NAND2_X1 U12803 ( .A1(n14847), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14836) );
  INV_X1 U12804 ( .A(n15682), .ZN(n15989) );
  NAND2_X1 U12805 ( .A1(n18363), .A2(n18700), .ZN(n18362) );
  AND2_X1 U12806 ( .A1(n15365), .A2(n15364), .ZN(n15957) );
  NAND2_X1 U12807 ( .A1(n15362), .A2(n15363), .ZN(n15365) );
  XNOR2_X1 U12808 ( .A(n11210), .B(n11209), .ZN(n13327) );
  CLKBUF_X1 U12809 ( .A(n13124), .Z(n15162) );
  NAND2_X1 U12810 ( .A1(n12642), .A2(n10451), .ZN(n12632) );
  NAND4_X1 U12811 ( .A1(n10519), .A2(n10516), .A3(n10850), .A4(n10515), .ZN(
        n10517) );
  NAND2_X1 U12812 ( .A1(n10519), .A2(n10516), .ZN(n10494) );
  NAND2_X2 U12813 ( .A1(n10498), .A2(n10499), .ZN(n10519) );
  AND3_X1 U12814 ( .A1(n12161), .A2(n10548), .A3(n10549), .ZN(n20352) );
  AOI22_X1 U12815 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U12816 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10207) );
  NAND2_X1 U12817 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10363) );
  NAND2_X1 U12818 ( .A1(n15467), .A2(n15468), .ZN(n15466) );
  AND2_X1 U12819 ( .A1(n19784), .A2(n16237), .ZN(n19793) );
  AND2_X1 U12820 ( .A1(n10444), .A2(n16237), .ZN(n10436) );
  CLKBUF_X1 U12821 ( .A(n13911), .Z(n13923) );
  NAND2_X1 U12822 ( .A1(n12632), .A2(n10459), .ZN(n12861) );
  NOR2_X1 U12823 ( .A1(n10459), .A2(n13738), .ZN(n10460) );
  NOR2_X1 U12824 ( .A1(n14977), .A2(n20963), .ZN(n12044) );
  NAND4_X4 U12825 ( .A1(n10989), .A2(n10988), .A3(n10987), .A4(n10986), .ZN(
        n13301) );
  NAND2_X1 U12826 ( .A1(n11225), .A2(n13171), .ZN(n13124) );
  NAND2_X1 U12827 ( .A1(n12845), .A2(n12846), .ZN(n15480) );
  NAND2_X1 U12828 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10370) );
  NAND2_X1 U12829 ( .A1(n9611), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10364) );
  NAND2_X1 U12830 ( .A1(n9611), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10208) );
  NAND2_X1 U12831 ( .A1(n14037), .A2(n14038), .ZN(n15493) );
  OR2_X1 U12832 ( .A1(n13535), .A2(n13531), .ZN(n13538) );
  NOR2_X4 U12833 ( .A1(n14167), .A2(n19394), .ZN(n16368) );
  AND2_X1 U12834 ( .A1(n16801), .A2(n15003), .ZN(n20811) );
  INV_X1 U12835 ( .A(n20811), .ZN(n15151) );
  INV_X2 U12836 ( .A(n13223), .ZN(n20783) );
  OR4_X1 U12837 ( .A1(n15971), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15943), .A4(n15941), .ZN(n10192) );
  AND2_X2 U12838 ( .A1(n12855), .A2(n17076), .ZN(n15341) );
  NOR2_X1 U12839 ( .A1(n15309), .A2(n15311), .ZN(n10193) );
  OR2_X1 U12840 ( .A1(n20721), .A2(n12036), .ZN(n10194) );
  NOR2_X2 U12841 ( .A1(n13387), .A2(n13663), .ZN(n10195) );
  NAND2_X1 U12842 ( .A1(n12141), .A2(n16656), .ZN(n14847) );
  INV_X2 U12843 ( .A(n18049), .ZN(n18098) );
  NAND2_X1 U12844 ( .A1(n13739), .A2(n10479), .ZN(n10196) );
  INV_X1 U12845 ( .A(n15905), .ZN(n10682) );
  INV_X1 U12846 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12809) );
  INV_X1 U12847 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14419) );
  INV_X1 U12848 ( .A(n14168), .ZN(n17708) );
  NOR2_X1 U12849 ( .A1(n14173), .A2(n14169), .ZN(n14170) );
  INV_X1 U12850 ( .A(n14170), .ZN(n16367) );
  INV_X1 U12851 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10683) );
  OR2_X1 U12852 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n11319) );
  NOR2_X1 U12853 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13770) );
  AND2_X2 U12854 ( .A1(n21068), .A2(n12146), .ZN(n21061) );
  INV_X1 U12855 ( .A(n13364), .ZN(n12216) );
  INV_X1 U12856 ( .A(n10419), .ZN(n14489) );
  NOR2_X1 U12857 ( .A1(n19432), .A2(n18573), .ZN(n18299) );
  INV_X1 U12858 ( .A(n18299), .ZN(n18364) );
  AND2_X1 U12859 ( .A1(n10533), .A2(n17014), .ZN(n10199) );
  AND2_X1 U12860 ( .A1(n14017), .A2(n10827), .ZN(n10200) );
  INV_X1 U12861 ( .A(n11073), .ZN(n11741) );
  NAND2_X1 U12862 ( .A1(n10501), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10502) );
  OAI21_X1 U12863 ( .B1(n11137), .B2(n13127), .A(n14982), .ZN(n11129) );
  AND2_X1 U12864 ( .A1(n20864), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11910) );
  AND2_X1 U12865 ( .A1(n20854), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11893) );
  OR2_X1 U12866 ( .A1(n10614), .A2(n12559), .ZN(n10615) );
  OR2_X1 U12867 ( .A1(n10599), .A2(n12444), .ZN(n10542) );
  AND2_X1 U12868 ( .A1(n12624), .A2(n16237), .ZN(n10403) );
  INV_X1 U12869 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11894) );
  INV_X1 U12870 ( .A(n11909), .ZN(n11915) );
  OR2_X1 U12871 ( .A1(n11931), .A2(n11893), .ZN(n11895) );
  INV_X1 U12872 ( .A(n11192), .ZN(n11159) );
  OAI22_X1 U12873 ( .A1(n10596), .A2(n10575), .B1(n10645), .B2(n19950), .ZN(
        n10578) );
  AOI22_X1 U12874 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9611), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10413) );
  NAND2_X1 U12875 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10369) );
  INV_X1 U12876 ( .A(n11713), .ZN(n11714) );
  INV_X1 U12877 ( .A(n14720), .ZN(n11493) );
  NAND2_X1 U12878 ( .A1(n11935), .A2(n12105), .ZN(n11934) );
  NAND2_X1 U12879 ( .A1(n14977), .A2(n14957), .ZN(n11226) );
  INV_X1 U12880 ( .A(n11245), .ZN(n11242) );
  INV_X1 U12881 ( .A(n12431), .ZN(n12389) );
  AND2_X1 U12882 ( .A1(n19763), .A2(n15585), .ZN(n12312) );
  AND4_X1 U12883 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10345) );
  OR2_X1 U12884 ( .A1(n11931), .A2(n11930), .ZN(n12905) );
  INV_X1 U12885 ( .A(n14603), .ZN(n11683) );
  OR2_X1 U12886 ( .A1(n11808), .A2(n11807), .ZN(n11809) );
  NOR2_X1 U12887 ( .A1(n11676), .A2(n14620), .ZN(n11677) );
  OR2_X1 U12888 ( .A1(n11167), .A2(n11166), .ZN(n12116) );
  INV_X1 U12889 ( .A(n11531), .ZN(n11532) );
  NAND2_X2 U12890 ( .A1(n11245), .A2(n11244), .ZN(n11301) );
  INV_X1 U12891 ( .A(n12609), .ZN(n12598) );
  NAND2_X1 U12892 ( .A1(n12517), .A2(n12519), .ZN(n12520) );
  OR2_X1 U12893 ( .A1(n12439), .A2(n12438), .ZN(n12461) );
  AND2_X1 U12894 ( .A1(n12312), .A2(n13847), .ZN(n12313) );
  INV_X1 U12895 ( .A(n10377), .ZN(n10443) );
  NOR2_X1 U12896 ( .A1(n15751), .A2(n10743), .ZN(n10744) );
  INV_X1 U12897 ( .A(n15893), .ZN(n10687) );
  AND2_X1 U12898 ( .A1(n12627), .A2(n12626), .ZN(n12866) );
  INV_X1 U12899 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n21139) );
  INV_X1 U12900 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n21216) );
  NAND2_X1 U12901 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14166) );
  INV_X1 U12902 ( .A(n11630), .ZN(n11631) );
  NAND2_X1 U12903 ( .A1(n13297), .A2(n13301), .ZN(n11204) );
  NAND2_X1 U12904 ( .A1(n11761), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11808) );
  OR2_X1 U12905 ( .A1(n14886), .A2(n11319), .ZN(n11681) );
  NAND2_X1 U12906 ( .A1(n11589), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11630) );
  NOR2_X1 U12907 ( .A1(n11474), .A2(n11473), .ZN(n11494) );
  AND2_X1 U12908 ( .A1(n12002), .A2(n12001), .ZN(n14691) );
  AND2_X1 U12909 ( .A1(n11963), .A2(n11962), .ZN(n20696) );
  INV_X1 U12910 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13532) );
  AOI221_X1 U12911 ( .B1(n10786), .B2(n17060), .C1(n10786), .C2(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n10785), .ZN(n10951) );
  OR2_X1 U12912 ( .A1(n12228), .A2(n12227), .ZN(n12701) );
  INV_X1 U12913 ( .A(n14097), .ZN(n12331) );
  AND2_X1 U12914 ( .A1(n13708), .A2(n10952), .ZN(n17055) );
  NAND2_X1 U12915 ( .A1(n15329), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15328) );
  INV_X1 U12916 ( .A(n16039), .ZN(n15423) );
  AND2_X1 U12917 ( .A1(n16171), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16169) );
  NAND2_X1 U12918 ( .A1(n10832), .A2(n10350), .ZN(n10838) );
  NAND2_X1 U12919 ( .A1(n14012), .A2(n10200), .ZN(n10825) );
  AND2_X1 U12920 ( .A1(n12186), .A2(n12182), .ZN(n13087) );
  AND2_X1 U12921 ( .A1(n20223), .A2(n20585), .ZN(n20227) );
  AOI21_X1 U12922 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19387), .A(
        n14243), .ZN(n14249) );
  INV_X1 U12923 ( .A(n18942), .ZN(n16270) );
  INV_X1 U12924 ( .A(n16409), .ZN(n16410) );
  NOR2_X1 U12925 ( .A1(n18507), .A2(n18506), .ZN(n18505) );
  NOR2_X1 U12926 ( .A1(n16561), .A2(n16431), .ZN(n16294) );
  NAND2_X1 U12927 ( .A1(n16269), .A2(n19358), .ZN(n16439) );
  AND2_X1 U12928 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n11631), .ZN(
        n11632) );
  INV_X1 U12929 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16595) );
  NAND2_X1 U12930 ( .A1(n13583), .A2(n13582), .ZN(n20707) );
  AND4_X1 U12931 ( .A1(n11041), .A2(n11040), .A3(n11039), .A4(n11038), .ZN(
        n11047) );
  NAND2_X1 U12932 ( .A1(n11682), .A2(n11681), .ZN(n14603) );
  AND2_X1 U12933 ( .A1(n11494), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11511) );
  INV_X1 U12934 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11473) );
  INV_X1 U12935 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14137) );
  AND2_X1 U12936 ( .A1(n11968), .A2(n11967), .ZN(n13649) );
  NAND2_X1 U12937 ( .A1(n14992), .A2(n14981), .ZN(n16799) );
  INV_X1 U12938 ( .A(n13175), .ZN(n16503) );
  AND2_X1 U12939 ( .A1(n13775), .A2(n13774), .ZN(n13840) );
  AND3_X1 U12940 ( .A1(n13661), .A2(n15158), .A3(n13334), .ZN(n13423) );
  INV_X1 U12941 ( .A(n13531), .ZN(n15158) );
  NOR2_X1 U12942 ( .A1(n20899), .A2(n13768), .ZN(n20869) );
  AND4_X1 U12943 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n11016), .ZN(
        n11024) );
  NAND2_X1 U12944 ( .A1(n17047), .A2(n19936), .ZN(n10459) );
  OR2_X1 U12945 ( .A1(n19599), .A2(n12838), .ZN(n19737) );
  INV_X1 U12946 ( .A(n12760), .ZN(n12765) );
  OAI21_X1 U12947 ( .B1(n12758), .B2(n12757), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12759) );
  INV_X1 U12948 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15880) );
  INV_X1 U12949 ( .A(n15677), .ZN(n15675) );
  INV_X1 U12950 ( .A(n15750), .ZN(n15764) );
  OR2_X1 U12951 ( .A1(n15502), .A2(n10362), .ZN(n10738) );
  OAI211_X1 U12952 ( .C1(n14012), .C2(n10827), .A(n10826), .B(n10825), .ZN(
        n16201) );
  NAND2_X1 U12953 ( .A1(n13750), .A2(n13747), .ZN(n19928) );
  NAND2_X1 U12954 ( .A1(n20569), .A2(n10955), .ZN(n10956) );
  NAND2_X1 U12955 ( .A1(n10953), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20569) );
  OR2_X1 U12956 ( .A1(n20582), .A2(n16222), .ZN(n20108) );
  OR2_X1 U12957 ( .A1(n20582), .A2(n20609), .ZN(n20147) );
  NAND2_X1 U12958 ( .A1(n20054), .A2(n20599), .ZN(n20576) );
  NAND3_X1 U12959 ( .A1(n20585), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20425), 
        .ZN(n13859) );
  INV_X1 U12960 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20491) );
  INV_X1 U12961 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18254) );
  NOR2_X1 U12962 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17429), .ZN(n17415) );
  NOR2_X1 U12963 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17453), .ZN(n17442) );
  NOR2_X1 U12964 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17478), .ZN(n17461) );
  NOR2_X1 U12965 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17580), .ZN(n17561) );
  NOR2_X1 U12966 ( .A1(n17431), .A2(n17758), .ZN(n17744) );
  OAI21_X1 U12967 ( .B1(n18926), .B2(n16285), .A(n19357), .ZN(n16558) );
  NOR2_X1 U12968 ( .A1(n18693), .A2(n18454), .ZN(n18251) );
  OR2_X1 U12969 ( .A1(n18259), .A2(n16413), .ZN(n16414) );
  NOR2_X1 U12970 ( .A1(n18496), .A2(n18495), .ZN(n18494) );
  NOR2_X1 U12971 ( .A1(n16294), .A2(n16293), .ZN(n16430) );
  INV_X1 U12972 ( .A(n18879), .ZN(n19397) );
  INV_X1 U12973 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19387) );
  OR2_X1 U12974 ( .A1(n12959), .A2(n20633), .ZN(n12992) );
  NAND2_X1 U12975 ( .A1(n11632), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11676) );
  NAND2_X1 U12976 ( .A1(n13574), .A2(n13573), .ZN(n13928) );
  AND2_X1 U12977 ( .A1(n13928), .A2(n13575), .ZN(n20676) );
  INV_X1 U12978 ( .A(n20707), .ZN(n20684) );
  NOR2_X2 U12979 ( .A1(n14378), .A2(n14738), .ZN(n16648) );
  NAND2_X1 U12980 ( .A1(n13077), .A2(n14967), .ZN(n16645) );
  AND2_X1 U12981 ( .A1(n16751), .A2(n16750), .ZN(n16753) );
  NAND2_X1 U12982 ( .A1(n11441), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11474) );
  OR2_X1 U12983 ( .A1(n11381), .A2(n11383), .ZN(n11405) );
  INV_X1 U12984 ( .A(n14963), .ZN(n14959) );
  OR2_X1 U12985 ( .A1(n12150), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16817) );
  AND2_X1 U12986 ( .A1(n14968), .A2(n14967), .ZN(n14992) );
  OR2_X1 U12987 ( .A1(n16801), .A2(n20827), .ZN(n16807) );
  INV_X1 U12988 ( .A(n20844), .ZN(n20806) );
  INV_X1 U12989 ( .A(n16799), .ZN(n20827) );
  AND2_X1 U12990 ( .A1(n15132), .A2(n20852), .ZN(n20847) );
  NAND2_X1 U12991 ( .A1(n20963), .A2(n13287), .ZN(n13768) );
  INV_X1 U12992 ( .A(n16539), .ZN(n15186) );
  OAI21_X1 U12993 ( .B1(n13285), .B2(n15192), .A(n13536), .ZN(n13316) );
  INV_X1 U12994 ( .A(n13786), .ZN(n13819) );
  INV_X1 U12995 ( .A(n9606), .ZN(n13663) );
  INV_X1 U12996 ( .A(n13770), .ZN(n20893) );
  AND2_X1 U12997 ( .A1(n13423), .A2(n13663), .ZN(n13637) );
  INV_X1 U12998 ( .A(n20856), .ZN(n20888) );
  INV_X1 U12999 ( .A(n20911), .ZN(n20956) );
  NOR2_X1 U13000 ( .A1(n14782), .A2(n13768), .ZN(n13682) );
  INV_X1 U13001 ( .A(n15254), .ZN(n20902) );
  INV_X1 U13002 ( .A(n15269), .ZN(n20928) );
  INV_X1 U13003 ( .A(n15292), .ZN(n20952) );
  INV_X1 U13004 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20905) );
  INV_X1 U13005 ( .A(n21051), .ZN(n20973) );
  INV_X1 U13006 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20972) );
  NAND2_X1 U13007 ( .A1(n12844), .A2(n12843), .ZN(n19744) );
  INV_X1 U13008 ( .A(n19748), .ZN(n19692) );
  XNOR2_X1 U13009 ( .A(n13055), .B(n13054), .ZN(n20599) );
  INV_X1 U13010 ( .A(n19834), .ZN(n19858) );
  NOR2_X1 U13011 ( .A1(n19869), .A2(n19900), .ZN(n19899) );
  INV_X1 U13012 ( .A(n12987), .ZN(n12951) );
  AND2_X1 U13013 ( .A1(n13566), .A2(n13565), .ZN(n16938) );
  INV_X1 U13014 ( .A(n16950), .ZN(n16954) );
  NOR2_X1 U13015 ( .A1(n14471), .A2(n14470), .ZN(n16998) );
  AND2_X1 U13016 ( .A1(n13750), .A2(n20620), .ZN(n19920) );
  AND2_X1 U13017 ( .A1(n13090), .A2(n13089), .ZN(n20582) );
  OAI21_X1 U13018 ( .B1(n16227), .B2(n16230), .A(n16226), .ZN(n19967) );
  NOR2_X1 U13019 ( .A1(n20222), .A2(n20147), .ZN(n20016) );
  OAI21_X1 U13020 ( .B1(n20029), .B2(n20028), .A(n20027), .ZN(n20046) );
  OAI21_X1 U13021 ( .B1(n20074), .B2(n21204), .A(n20058), .ZN(n20076) );
  NOR2_X2 U13022 ( .A1(n20429), .A2(n20108), .ZN(n20187) );
  NAND2_X1 U13023 ( .A1(n20199), .A2(n20198), .ZN(n20217) );
  INV_X1 U13024 ( .A(n20208), .ZN(n20216) );
  NAND2_X1 U13025 ( .A1(n20054), .A2(n16223), .ZN(n20222) );
  INV_X1 U13026 ( .A(n20294), .ZN(n20312) );
  NOR2_X2 U13027 ( .A1(n20361), .A2(n20576), .ZN(n20347) );
  INV_X1 U13028 ( .A(n20359), .ZN(n20384) );
  OAI21_X1 U13029 ( .B1(n20400), .B2(n20399), .A(n20398), .ZN(n20419) );
  INV_X1 U13030 ( .A(n20367), .ZN(n20441) );
  INV_X1 U13031 ( .A(n20376), .ZN(n20460) );
  NOR2_X2 U13032 ( .A1(n20361), .A2(n20429), .ZN(n20481) );
  AND2_X1 U13033 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10807), .ZN(n17073) );
  INV_X1 U13034 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20517) );
  INV_X1 U13035 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19600) );
  INV_X1 U13036 ( .A(n17101), .ZN(n19365) );
  NOR2_X1 U13037 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17392), .ZN(n17379) );
  NOR2_X1 U13038 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17408), .ZN(n17398) );
  INV_X1 U13039 ( .A(n17656), .ZN(n17638) );
  NOR2_X1 U13040 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17550), .ZN(n17534) );
  INV_X1 U13041 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17581) );
  AOI211_X1 U13042 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n19574), .A(n19414), .B(
        n17295), .ZN(n17608) );
  NOR4_X2 U13043 ( .A1(n18902), .A2(n19590), .A3(n17651), .A4(n19418), .ZN(
        n17649) );
  NOR2_X1 U13044 ( .A1(n17479), .A2(n17812), .ZN(n17788) );
  NAND2_X1 U13045 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17911), .ZN(n17890) );
  AOI21_X1 U13046 ( .B1(n16268), .B2(n14254), .A(n16296), .ZN(n16557) );
  NAND2_X1 U13047 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17975), .ZN(n17971) );
  NAND2_X1 U13048 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18014), .ZN(n18013) );
  INV_X1 U13049 ( .A(n17945), .ZN(n18094) );
  INV_X1 U13050 ( .A(n18251), .ZN(n18717) );
  INV_X1 U13051 ( .A(n18770), .ZN(n18751) );
  NOR2_X2 U13052 ( .A1(n18590), .A2(n18068), .ZN(n18497) );
  NAND2_X1 U13053 ( .A1(n18554), .A2(n18555), .ZN(n18553) );
  NOR2_X1 U13054 ( .A1(n18639), .A2(n18887), .ZN(n18660) );
  INV_X1 U13055 ( .A(n18898), .ZN(n18887) );
  INV_X1 U13056 ( .A(n18799), .ZN(n18822) );
  INV_X1 U13057 ( .A(n19382), .ZN(n19371) );
  AOI21_X2 U13058 ( .B1(n16430), .B2(n16429), .A(n19413), .ZN(n18898) );
  NOR2_X1 U13059 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19524), .ZN(
        n19549) );
  INV_X1 U13060 ( .A(n19069), .ZN(n19089) );
  INV_X1 U13061 ( .A(n19157), .ZN(n19159) );
  NOR2_X1 U13062 ( .A1(n19002), .A2(n19164), .ZN(n18950) );
  INV_X1 U13063 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19534) );
  INV_X1 U13064 ( .A(n19568), .ZN(n19575) );
  NOR2_X1 U13065 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12797), .ZN(n17252)
         );
  INV_X1 U13066 ( .A(n21049), .ZN(n13574) );
  OR3_X1 U13067 ( .A1(n14563), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14544), .ZN(
        n14545) );
  NAND2_X1 U13068 ( .A1(n16578), .A2(n14398), .ZN(n14623) );
  NAND2_X1 U13069 ( .A1(n16630), .A2(n14396), .ZN(n16619) );
  AND2_X1 U13070 ( .A1(n16601), .A2(n13577), .ZN(n14655) );
  NAND2_X1 U13071 ( .A1(n20721), .A2(n13297), .ZN(n14731) );
  OR2_X1 U13072 ( .A1(n14378), .A2(n14377), .ZN(n16652) );
  INV_X1 U13073 ( .A(n20724), .ZN(n20748) );
  NOR2_X1 U13074 ( .A1(n13199), .A2(n13198), .ZN(n13223) );
  INV_X1 U13075 ( .A(n20778), .ZN(n13247) );
  NAND2_X1 U13076 ( .A1(n14992), .A2(n14974), .ZN(n20844) );
  INV_X1 U13077 ( .A(n20849), .ZN(n20836) );
  INV_X1 U13078 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20864) );
  AOI22_X1 U13079 ( .A1(n15195), .A2(n15193), .B1(n20861), .B2(n15198), .ZN(
        n15243) );
  NAND2_X1 U13080 ( .A1(n13286), .A2(n9606), .ZN(n15238) );
  AOI22_X1 U13081 ( .A1(n13791), .A2(n13788), .B1(n20861), .B2(n15246), .ZN(
        n13822) );
  NAND2_X1 U13082 ( .A1(n13504), .A2(n13663), .ZN(n13846) );
  AOI22_X1 U13083 ( .A1(n15250), .A2(n15247), .B1(n15246), .B2(n20899), .ZN(
        n15297) );
  INV_X1 U13084 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13435) );
  AOI21_X1 U13085 ( .B1(n13604), .B2(n13605), .A(n13603), .ZN(n13645) );
  INV_X1 U13086 ( .A(n13642), .ZN(n13485) );
  AOI22_X1 U13087 ( .A1(n20862), .A2(n20870), .B1(n20861), .B2(n20860), .ZN(
        n20892) );
  OR2_X1 U13088 ( .A1(n13538), .A2(n9606), .ZN(n20911) );
  INV_X1 U13089 ( .A(n13668), .ZN(n20939) );
  INV_X1 U13090 ( .A(n13385), .ZN(n13414) );
  OR2_X1 U13091 ( .A1(n13387), .A2(n9606), .ZN(n13895) );
  INV_X1 U13092 ( .A(n13905), .ZN(n20951) );
  INV_X1 U13093 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20962) );
  INV_X1 U13094 ( .A(n21038), .ZN(n20966) );
  AND2_X1 U13095 ( .A1(n20972), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21048) );
  INV_X1 U13096 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21109) );
  NAND2_X1 U13097 ( .A1(n19599), .A2(n12850), .ZN(n19748) );
  INV_X1 U13098 ( .A(n19734), .ZN(n19684) );
  INV_X1 U13099 ( .A(n19743), .ZN(n19726) );
  AND2_X1 U13100 ( .A1(n12773), .A2(n17073), .ZN(n19784) );
  XNOR2_X1 U13101 ( .A(n13061), .B(n13060), .ZN(n20054) );
  AND2_X1 U13102 ( .A1(n12635), .A2(n17073), .ZN(n19834) );
  INV_X1 U13103 ( .A(n19848), .ZN(n19863) );
  INV_X1 U13104 ( .A(n19869), .ZN(n19902) );
  INV_X1 U13105 ( .A(n15341), .ZN(n12986) );
  NAND2_X1 U13106 ( .A1(n12860), .A2(n10959), .ZN(n16950) );
  INV_X1 U13107 ( .A(n17013), .ZN(n19926) );
  INV_X1 U13108 ( .A(n16497), .ZN(n17022) );
  INV_X1 U13109 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17068) );
  AOI211_X2 U13110 ( .C1(n16231), .C2(n16230), .A(n16229), .B(n20395), .ZN(
        n19971) );
  INV_X1 U13111 ( .A(n20016), .ZN(n19999) );
  AOI21_X1 U13112 ( .B1(n13857), .B2(n20585), .A(n13856), .ZN(n20020) );
  INV_X1 U13113 ( .A(n20042), .ZN(n20050) );
  INV_X1 U13114 ( .A(n20071), .ZN(n20079) );
  INV_X1 U13115 ( .A(n20102), .ZN(n20099) );
  INV_X1 U13116 ( .A(n20125), .ZN(n20133) );
  INV_X1 U13117 ( .A(n20187), .ZN(n20177) );
  NAND2_X1 U13118 ( .A1(n20149), .A2(n20148), .ZN(n20208) );
  OR2_X1 U13119 ( .A1(n20390), .A2(n20222), .ZN(n20251) );
  INV_X1 U13120 ( .A(n20297), .ZN(n20315) );
  OR2_X1 U13121 ( .A1(n20390), .A2(n20360), .ZN(n20387) );
  AOI211_X2 U13122 ( .C1(n20397), .C2(n20399), .A(n20396), .B(n20395), .ZN(
        n20422) );
  AOI221_X2 U13123 ( .B1(n20429), .B2(n20430), .C1(n20428), .C2(n20430), .A(
        n20427), .ZN(n20487) );
  INV_X1 U13124 ( .A(n20566), .ZN(n20497) );
  AOI21_X1 U13125 ( .B1(n19358), .B2(n19357), .A(n18101), .ZN(n19590) );
  NAND2_X1 U13126 ( .A1(n19572), .A2(n19365), .ZN(n17274) );
  INV_X1 U13127 ( .A(n17608), .ZN(n17663) );
  INV_X1 U13128 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18547) );
  NOR2_X1 U13129 ( .A1(n17673), .A2(n17691), .ZN(n17696) );
  NOR2_X1 U13130 ( .A1(n17860), .A2(n17890), .ZN(n17874) );
  NOR2_X2 U13131 ( .A1(n17941), .A2(n18954), .ZN(n17942) );
  AND2_X1 U13132 ( .A1(n18087), .A2(n17950), .ZN(n18061) );
  NOR2_X1 U13133 ( .A1(n18191), .A2(n18056), .ZN(n18059) );
  NOR2_X1 U13134 ( .A1(n16322), .A2(n16321), .ZN(n18076) );
  NOR2_X1 U13135 ( .A1(n19569), .A2(n18119), .ZN(n18131) );
  INV_X1 U13136 ( .A(n18119), .ZN(n18139) );
  INV_X1 U13137 ( .A(n18497), .ZN(n18471) );
  INV_X1 U13138 ( .A(n17106), .ZN(n18590) );
  INV_X1 U13139 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19403) );
  INV_X1 U13140 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18918) );
  AOI211_X1 U13141 ( .C1(n19572), .C2(n19379), .A(n16298), .B(n18922), .ZN(
        n19555) );
  INV_X1 U13142 ( .A(n19233), .ZN(n19231) );
  INV_X1 U13143 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19577) );
  INV_X1 U13144 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19524) );
  INV_X1 U13145 ( .A(n19521), .ZN(n19433) );
  INV_X1 U13146 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19448) );
  OAI21_X1 U13147 ( .B1(n14815), .B2(n14731), .A(n12038), .ZN(P1_U2842) );
  OAI21_X1 U13148 ( .B1(n15964), .B2(n16957), .A(n10966), .ZN(P2_U2985) );
  AND3_X4 U13149 ( .A1(n10201), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U13150 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10205) );
  AND3_X4 U13151 ( .A1(n14499), .A2(n10201), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12605) );
  AND2_X4 U13152 ( .A1(n10202), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12607) );
  AOI22_X1 U13153 ( .A1(n12605), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10204) );
  AND2_X4 U13154 ( .A1(n16212), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10421) );
  AND2_X4 U13155 ( .A1(n14482), .A2(n17035), .ZN(n10420) );
  AOI22_X1 U13156 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10203) );
  NAND4_X1 U13157 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10214) );
  AOI22_X1 U13158 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U13159 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10210) );
  AOI22_X1 U13160 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10209) );
  NAND2_X1 U13161 ( .A1(n10773), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14408) );
  NAND2_X1 U13162 ( .A1(n20615), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10802) );
  INV_X1 U13163 ( .A(n10802), .ZN(n10215) );
  NAND2_X1 U13164 ( .A1(n10939), .A2(n10215), .ZN(n10217) );
  NAND2_X1 U13165 ( .A1(n20605), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10216) );
  NAND2_X1 U13166 ( .A1(n10217), .A2(n10216), .ZN(n10275) );
  NOR2_X1 U13167 ( .A1(n14499), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10218) );
  NAND2_X1 U13168 ( .A1(n14499), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10219) );
  NAND3_X1 U13169 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10786), .A3(
        n17060), .ZN(n10800) );
  INV_X1 U13170 ( .A(n10421), .ZN(n10221) );
  AOI22_X1 U13171 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12423), .B1(
        n12202), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U13172 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U13173 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10223) );
  INV_X1 U13174 ( .A(n10418), .ZN(n10239) );
  AOI22_X1 U13175 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10222) );
  NAND4_X1 U13176 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n10234) );
  AND2_X1 U13177 ( .A1(n12607), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10295) );
  AOI22_X1 U13178 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12368), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10232) );
  AOI22_X1 U13179 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12366), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10231) );
  INV_X1 U13180 ( .A(n10797), .ZN(n10226) );
  INV_X1 U13181 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19956) );
  NAND2_X1 U13182 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12429), .ZN(
        n10227) );
  OAI21_X1 U13183 ( .B1(n12431), .B2(n19956), .A(n10227), .ZN(n10228) );
  AOI21_X1 U13184 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n10228), .ZN(n10230) );
  NAND2_X1 U13185 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10229) );
  NAND4_X1 U13186 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .ZN(
        n10233) );
  AOI22_X1 U13187 ( .A1(n10420), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10235) );
  INV_X1 U13188 ( .A(n10235), .ZN(n10238) );
  AOI22_X1 U13189 ( .A1(n12605), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10236) );
  INV_X1 U13190 ( .A(n10236), .ZN(n10237) );
  NOR2_X1 U13191 ( .A1(n10238), .A2(n10237), .ZN(n10242) );
  AOI22_X1 U13192 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9600), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U13193 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10240) );
  NAND3_X1 U13194 ( .A1(n10242), .A2(n10241), .A3(n10240), .ZN(n10243) );
  AOI22_X1 U13195 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U13196 ( .A1(n12605), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U13197 ( .A1(n10420), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U13198 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10244) );
  NAND4_X1 U13199 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10248) );
  NAND2_X1 U13200 ( .A1(n10248), .A2(n10416), .ZN(n10249) );
  NAND2_X4 U13201 ( .A1(n10250), .A2(n10249), .ZN(n17047) );
  AOI22_X1 U13202 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9611), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U13203 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U13204 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U13205 ( .A1(n12605), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10251) );
  NAND4_X1 U13206 ( .A1(n10254), .A2(n10253), .A3(n10252), .A4(n10251), .ZN(
        n10260) );
  AOI22_X1 U13207 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U13208 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U13209 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U13210 ( .A1(n12605), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10255) );
  NAND4_X1 U13211 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10259) );
  MUX2_X2 U13212 ( .A(n10260), .B(n10259), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19936) );
  MUX2_X1 U13213 ( .A(n10800), .B(n12676), .S(n10172), .Z(n10792) );
  INV_X1 U13214 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10261) );
  MUX2_X1 U13215 ( .A(n10792), .B(n10261), .S(n10773), .Z(n10639) );
  AOI22_X1 U13216 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n12423), .B1(
        n12202), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U13217 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U13218 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U13219 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10263) );
  NAND4_X1 U13220 ( .A1(n10266), .A2(n10265), .A3(n10264), .A4(n10263), .ZN(
        n10273) );
  INV_X1 U13221 ( .A(n10295), .ZN(n10565) );
  AOI22_X1 U13222 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n12351), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U13223 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12366), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10270) );
  INV_X1 U13224 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19945) );
  INV_X1 U13225 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12479) );
  OAI22_X1 U13226 ( .A1(n19945), .A2(n12431), .B1(n12479), .B2(n12350), .ZN(
        n10267) );
  AOI21_X1 U13227 ( .B1(n12368), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n10267), .ZN(n10269) );
  NAND2_X1 U13228 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10268) );
  NAND4_X1 U13229 ( .A1(n10271), .A2(n10270), .A3(n10269), .A4(n10268), .ZN(
        n10272) );
  XNOR2_X1 U13230 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10274) );
  XNOR2_X1 U13231 ( .A(n10275), .B(n10274), .ZN(n10936) );
  INV_X1 U13232 ( .A(n10936), .ZN(n10276) );
  MUX2_X1 U13233 ( .A(n10573), .B(n10276), .S(n13721), .Z(n10787) );
  INV_X1 U13234 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14126) );
  MUX2_X1 U13235 ( .A(n10787), .B(n14126), .S(n10773), .Z(n10636) );
  AOI22_X1 U13236 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12423), .B1(
        n12202), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13237 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U13238 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U13239 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10278) );
  NAND4_X1 U13240 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10289) );
  AOI22_X1 U13241 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12368), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13242 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12366), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10286) );
  INV_X1 U13243 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16234) );
  NAND2_X1 U13244 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12429), .ZN(
        n10282) );
  OAI21_X1 U13245 ( .B1(n12431), .B2(n16234), .A(n10282), .ZN(n10283) );
  AOI21_X1 U13246 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n10283), .ZN(n10285) );
  NAND2_X1 U13247 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10284) );
  NAND4_X1 U13248 ( .A1(n10287), .A2(n10286), .A3(n10285), .A4(n10284), .ZN(
        n10288) );
  NOR2_X1 U13249 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n10290) );
  MUX2_X1 U13250 ( .A(n12655), .B(n10290), .S(n10773), .Z(n10635) );
  NAND2_X1 U13251 ( .A1(n10636), .A2(n10635), .ZN(n10631) );
  AOI22_X1 U13252 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n12423), .B1(
        n12202), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13253 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__3__SCAN_IN), .B2(n12365), .ZN(n10293) );
  AOI22_X1 U13254 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13255 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10291) );
  NAND4_X1 U13256 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n10301) );
  AOI22_X1 U13257 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12351), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10299) );
  AOI22_X1 U13258 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10295), .B1(
        n12366), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10298) );
  INV_X1 U13259 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19950) );
  NAND2_X1 U13260 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10296) );
  NAND4_X1 U13261 ( .A1(n10299), .A2(n10298), .A3(n10297), .A4(n10296), .ZN(
        n10300) );
  NOR2_X1 U13262 ( .A1(n10301), .A2(n10300), .ZN(n12671) );
  AND2_X1 U13263 ( .A1(n10303), .A2(n10302), .ZN(n10304) );
  NOR2_X1 U13264 ( .A1(n10305), .A2(n10304), .ZN(n10801) );
  INV_X1 U13265 ( .A(n10801), .ZN(n10306) );
  MUX2_X1 U13266 ( .A(n12671), .B(n10306), .S(n13721), .Z(n10791) );
  MUX2_X1 U13267 ( .A(n10791), .B(P2_EBX_REG_3__SCAN_IN), .S(n10773), .Z(
        n10630) );
  AOI22_X1 U13268 ( .A1(n12423), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12202), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13269 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13270 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13271 ( .A1(n12424), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10307) );
  NAND4_X1 U13272 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10317) );
  AOI22_X1 U13273 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U13274 ( .A1(n12366), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10314) );
  INV_X1 U13275 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19960) );
  INV_X1 U13276 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10601) );
  OAI22_X1 U13277 ( .A1(n12431), .A2(n19960), .B1(n10601), .B2(n12350), .ZN(
        n10311) );
  AOI21_X1 U13278 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n10311), .ZN(n10313) );
  NAND2_X1 U13279 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10312) );
  NAND4_X1 U13280 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n10316) );
  NOR2_X1 U13281 ( .A1(n10317), .A2(n10316), .ZN(n12682) );
  MUX2_X1 U13282 ( .A(n12682), .B(P2_EBX_REG_5__SCAN_IN), .S(n10773), .Z(
        n10626) );
  AOI22_X1 U13283 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12423), .B1(
        n12202), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13284 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13285 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13286 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10318) );
  NAND4_X1 U13287 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n10328) );
  AOI22_X1 U13288 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12368), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13289 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12366), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10325) );
  INV_X1 U13290 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19970) );
  INV_X1 U13291 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10658) );
  OAI22_X1 U13292 ( .A1(n19970), .A2(n12431), .B1(n10658), .B2(n12350), .ZN(
        n10322) );
  AOI21_X1 U13293 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n10322), .ZN(n10324) );
  NAND2_X1 U13294 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10323) );
  NAND4_X1 U13295 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10327) );
  INV_X1 U13296 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n10329) );
  MUX2_X1 U13297 ( .A(n12687), .B(n10329), .S(n10773), .Z(n10673) );
  NAND2_X1 U13298 ( .A1(n12423), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10333) );
  NAND2_X1 U13299 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10332) );
  NAND2_X1 U13300 ( .A1(n12202), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10331) );
  NAND2_X1 U13301 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10330) );
  NAND2_X1 U13302 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10337) );
  NAND2_X1 U13303 ( .A1(n10277), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10336) );
  NAND2_X1 U13304 ( .A1(n12424), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10335) );
  NAND2_X1 U13305 ( .A1(n12384), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10334) );
  NAND2_X1 U13306 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10340) );
  NAND2_X1 U13307 ( .A1(n12351), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10339) );
  AOI22_X1 U13308 ( .A1(n12389), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n12429), .ZN(n10338) );
  AND3_X1 U13309 ( .A1(n10340), .A2(n10339), .A3(n10338), .ZN(n10346) );
  NAND2_X1 U13310 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10344) );
  NAND2_X1 U13311 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10343) );
  NAND2_X1 U13312 ( .A1(n12366), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10342) );
  NAND2_X1 U13313 ( .A1(n12365), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10341) );
  INV_X1 U13314 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10349) );
  MUX2_X1 U13315 ( .A(n10350), .B(n10349), .S(n10773), .Z(n10678) );
  INV_X1 U13316 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10351) );
  INV_X1 U13317 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19783) );
  NAND2_X1 U13318 ( .A1(n10773), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10702) );
  AND2_X1 U13319 ( .A1(n10773), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10730) );
  AND2_X1 U13320 ( .A1(n10773), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10727) );
  NAND2_X1 U13321 ( .A1(n10773), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U13322 ( .A1(n10773), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10717) );
  OAI21_X1 U13323 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n10773), .ZN(n10353) );
  INV_X1 U13324 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15564) );
  INV_X1 U13325 ( .A(n10715), .ZN(n10354) );
  NAND2_X1 U13326 ( .A1(n10773), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10762) );
  AND2_X1 U13327 ( .A1(n10773), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10766) );
  INV_X1 U13328 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16877) );
  INV_X1 U13329 ( .A(n10771), .ZN(n10360) );
  NAND2_X1 U13330 ( .A1(n14414), .A2(n10360), .ZN(n10356) );
  NAND2_X1 U13331 ( .A1(n10773), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10355) );
  NAND2_X1 U13332 ( .A1(n10773), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10776) );
  XOR2_X1 U13333 ( .A(n14408), .B(n14410), .Z(n10359) );
  INV_X1 U13334 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10358) );
  OAI21_X1 U13335 ( .B1(n10359), .B2(n10362), .A(n10358), .ZN(n14406) );
  INV_X1 U13336 ( .A(n10359), .ZN(n15370) );
  NAND3_X1 U13337 ( .A1(n15370), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10350), .ZN(n15661) );
  NAND2_X1 U13338 ( .A1(n14406), .A2(n15661), .ZN(n10784) );
  INV_X1 U13339 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15970) );
  NAND3_X1 U13340 ( .A1(n10773), .A2(P2_EBX_REG_27__SCAN_IN), .A3(n10360), 
        .ZN(n10361) );
  NAND2_X1 U13341 ( .A1(n10778), .A2(n10361), .ZN(n15391) );
  AOI22_X1 U13342 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U13343 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10366) );
  NAND4_X1 U13344 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10376) );
  AOI22_X1 U13345 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U13346 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13347 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10371) );
  NAND4_X1 U13348 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10375) );
  AOI22_X1 U13349 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13350 ( .A1(n12605), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13351 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13352 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10378) );
  NAND4_X1 U13353 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10382) );
  NAND2_X1 U13354 ( .A1(n10382), .A2(n10416), .ZN(n10389) );
  AOI22_X1 U13355 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13356 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13357 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U13358 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10383) );
  NAND4_X1 U13359 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10387) );
  NAND2_X1 U13360 ( .A1(n10387), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10388) );
  NAND2_X2 U13361 ( .A1(n10389), .A2(n10388), .ZN(n19952) );
  NAND2_X1 U13362 ( .A1(n12656), .A2(n19952), .ZN(n12624) );
  AOI22_X1 U13363 ( .A1(n10420), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U13364 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U13365 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10421), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13366 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10390) );
  NAND4_X1 U13367 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n10394) );
  AOI22_X1 U13368 ( .A1(n12605), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U13369 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9611), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U13370 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10395) );
  NAND4_X1 U13371 ( .A1(n10398), .A2(n10397), .A3(n10396), .A4(n10395), .ZN(
        n10399) );
  NAND2_X4 U13372 ( .A1(n10401), .A2(n10400), .ZN(n16237) );
  INV_X1 U13373 ( .A(n10452), .ZN(n10402) );
  INV_X2 U13374 ( .A(n19952), .ZN(n10435) );
  NAND2_X1 U13375 ( .A1(n12618), .A2(n10435), .ZN(n12622) );
  AOI22_X1 U13376 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U13377 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10405) );
  MUX2_X1 U13378 ( .A(n10150), .B(n16237), .S(n19952), .Z(n10407) );
  NAND2_X1 U13379 ( .A1(n10407), .A2(n10430), .ZN(n10411) );
  NAND2_X1 U13380 ( .A1(n12634), .A2(n10445), .ZN(n10408) );
  INV_X1 U13381 ( .A(n12634), .ZN(n10410) );
  AND2_X1 U13382 ( .A1(n12656), .A2(n12642), .ZN(n10409) );
  NAND2_X1 U13383 ( .A1(n10410), .A2(n10409), .ZN(n10478) );
  NAND2_X1 U13384 ( .A1(n12656), .A2(n19946), .ZN(n10454) );
  AOI22_X1 U13385 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13386 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13387 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10412) );
  AOI22_X1 U13388 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10420), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13389 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10424) );
  AOI22_X1 U13390 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10423) );
  NAND4_X1 U13391 ( .A1(n10426), .A2(n10425), .A3(n10424), .A4(n10423), .ZN(
        n10427) );
  NAND2_X1 U13392 ( .A1(n10454), .A2(n10444), .ZN(n10432) );
  NAND2_X1 U13393 ( .A1(n10435), .A2(n16237), .ZN(n10429) );
  NOR2_X2 U13394 ( .A1(n10430), .A2(n10429), .ZN(n10434) );
  NAND2_X1 U13395 ( .A1(n10434), .A2(n10431), .ZN(n10440) );
  AND2_X1 U13396 ( .A1(n10444), .A2(n19946), .ZN(n10433) );
  NAND2_X1 U13397 ( .A1(n10434), .A2(n10433), .ZN(n17046) );
  NAND3_X1 U13398 ( .A1(n17046), .A2(n10444), .A3(n17047), .ZN(n10438) );
  AND4_X2 U13399 ( .A1(n10436), .A2(n19946), .A3(n10452), .A4(n10435), .ZN(
        n10442) );
  INV_X1 U13400 ( .A(n10442), .ZN(n10437) );
  NAND2_X1 U13401 ( .A1(n10438), .A2(n10437), .ZN(n12771) );
  NAND2_X1 U13402 ( .A1(n19936), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10950) );
  NAND2_X1 U13403 ( .A1(n10506), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10449) );
  INV_X1 U13404 ( .A(n10440), .ZN(n10441) );
  NAND2_X1 U13405 ( .A1(n10443), .A2(n16237), .ZN(n12761) );
  NOR2_X1 U13406 ( .A1(n12761), .A2(n17047), .ZN(n12636) );
  NAND4_X1 U13407 ( .A1(n12636), .A2(n10451), .A3(n10465), .A4(n10150), .ZN(
        n10446) );
  INV_X2 U13408 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n20495) );
  NAND2_X1 U13409 ( .A1(n19598), .A2(n20495), .ZN(n17077) );
  NOR2_X1 U13410 ( .A1(n17077), .A2(n20605), .ZN(n10447) );
  NAND2_X1 U13411 ( .A1(n10452), .A2(n10451), .ZN(n10453) );
  NAND2_X1 U13412 ( .A1(n16237), .A2(n19952), .ZN(n10456) );
  NAND2_X1 U13413 ( .A1(n12634), .A2(n10460), .ZN(n12772) );
  INV_X1 U13414 ( .A(n12772), .ZN(n10461) );
  INV_X1 U13415 ( .A(n12776), .ZN(n10501) );
  INV_X1 U13416 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n14081) );
  INV_X1 U13417 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14076) );
  OAI22_X1 U13418 ( .A1(n14422), .A2(n14081), .B1(n20495), .B2(n14076), .ZN(
        n10462) );
  AOI21_X1 U13419 ( .B1(n10501), .B2(P2_EBX_REG_1__SCAN_IN), .A(n10462), .ZN(
        n10463) );
  AND2_X2 U13420 ( .A1(n10464), .A2(n10463), .ZN(n10485) );
  XNOR2_X2 U13421 ( .A(n10483), .B(n10485), .ZN(n10498) );
  AND3_X1 U13422 ( .A1(n10465), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10172), 
        .ZN(n10466) );
  INV_X1 U13423 ( .A(n14484), .ZN(n10468) );
  NOR2_X1 U13424 ( .A1(n17077), .A2(n20615), .ZN(n10467) );
  AOI21_X1 U13425 ( .B1(n10468), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10467), 
        .ZN(n10469) );
  NAND2_X1 U13426 ( .A1(n9605), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10482) );
  INV_X1 U13427 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n15507) );
  NAND2_X1 U13428 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10471) );
  AND2_X1 U13429 ( .A1(n17077), .A2(n10471), .ZN(n10472) );
  NAND2_X1 U13430 ( .A1(n10473), .A2(n10472), .ZN(n10474) );
  INV_X1 U13431 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10475) );
  NAND2_X1 U13432 ( .A1(n9674), .A2(n10478), .ZN(n13739) );
  NAND2_X1 U13433 ( .A1(n10196), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10480) );
  INV_X1 U13434 ( .A(n10483), .ZN(n10484) );
  OAI21_X1 U13435 ( .B1(n20597), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n20495), 
        .ZN(n10486) );
  AOI22_X1 U13436 ( .A1(n9610), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10487) );
  OAI21_X1 U13437 ( .B1(n9591), .B2(n14126), .A(n10487), .ZN(n10488) );
  NAND2_X1 U13438 ( .A1(n10489), .A2(n10490), .ZN(n10850) );
  INV_X1 U13439 ( .A(n10489), .ZN(n10492) );
  INV_X1 U13440 ( .A(n10490), .ZN(n10491) );
  OR2_X2 U13441 ( .A1(n10494), .A2(n10493), .ZN(n10495) );
  NAND2_X2 U13442 ( .A1(n10494), .A2(n10493), .ZN(n10851) );
  NAND2_X4 U13443 ( .A1(n10495), .A2(n10851), .ZN(n12161) );
  INV_X1 U13444 ( .A(n10496), .ZN(n10497) );
  NAND2_X1 U13445 ( .A1(n10503), .A2(n10502), .ZN(n10504) );
  NOR2_X1 U13446 ( .A1(n17077), .A2(n20588), .ZN(n10505) );
  AOI21_X1 U13447 ( .B1(n10506), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10505), .ZN(n10507) );
  NAND2_X1 U13448 ( .A1(n10508), .A2(n10507), .ZN(n10852) );
  INV_X1 U13449 ( .A(n10516), .ZN(n10510) );
  NAND2_X1 U13450 ( .A1(n10510), .A2(n10512), .ZN(n10511) );
  NAND3_X1 U13451 ( .A1(n10511), .A2(n10849), .A3(n10850), .ZN(n10514) );
  NAND2_X1 U13452 ( .A1(n10515), .A2(n10512), .ZN(n10513) );
  OAI211_X4 U13453 ( .C1(n10520), .C2(n10519), .A(n10518), .B(n10517), .ZN(
        n10549) );
  INV_X1 U13454 ( .A(n10549), .ZN(n14113) );
  INV_X1 U13455 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12443) );
  INV_X1 U13456 ( .A(n12161), .ZN(n10521) );
  NAND2_X1 U13457 ( .A1(n10521), .A2(n10549), .ZN(n10522) );
  INV_X1 U13458 ( .A(n17014), .ZN(n15928) );
  NAND2_X1 U13459 ( .A1(n15928), .A2(n10498), .ZN(n10546) );
  OR2_X2 U13460 ( .A1(n10522), .A2(n10546), .ZN(n10650) );
  NAND2_X1 U13461 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10524) );
  OAI211_X1 U13462 ( .C1(n20111), .C2(n12443), .A(n10524), .B(n10523), .ZN(
        n10525) );
  INV_X1 U13463 ( .A(n10525), .ZN(n10559) );
  INV_X1 U13464 ( .A(n10549), .ZN(n10526) );
  INV_X1 U13465 ( .A(n12161), .ZN(n13062) );
  NOR2_X1 U13466 ( .A1(n10533), .A2(n15928), .ZN(n10527) );
  INV_X1 U13467 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12441) );
  OAI22_X1 U13468 ( .A1(n16234), .A2(n10645), .B1(n10594), .B2(n12441), .ZN(
        n10532) );
  INV_X1 U13469 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10530) );
  INV_X1 U13470 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10529) );
  OAI22_X1 U13471 ( .A1(n10596), .A2(n10530), .B1(n10610), .B2(n10529), .ZN(
        n10531) );
  NOR2_X1 U13472 ( .A1(n10532), .A2(n10531), .ZN(n10558) );
  INV_X1 U13473 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13866) );
  INV_X1 U13474 ( .A(n10537), .ZN(n10535) );
  NOR2_X1 U13475 ( .A1(n10549), .A2(n10533), .ZN(n10534) );
  NAND2_X1 U13476 ( .A1(n10535), .A2(n10534), .ZN(n10655) );
  INV_X1 U13477 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12442) );
  OAI22_X1 U13478 ( .A1(n10593), .A2(n13866), .B1(n10655), .B2(n12442), .ZN(
        n10544) );
  NAND2_X1 U13479 ( .A1(n10549), .A2(n16217), .ZN(n10536) );
  INV_X1 U13480 ( .A(n10597), .ZN(n10654) );
  INV_X1 U13481 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12451) );
  INV_X1 U13482 ( .A(n10548), .ZN(n10538) );
  NOR2_X1 U13483 ( .A1(n10549), .A2(n10538), .ZN(n10539) );
  NAND2_X1 U13484 ( .A1(n10539), .A2(n12161), .ZN(n10599) );
  INV_X1 U13485 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12444) );
  NOR2_X1 U13486 ( .A1(n10549), .A2(n10546), .ZN(n10540) );
  NAND2_X1 U13487 ( .A1(n10540), .A2(n12161), .ZN(n10600) );
  INV_X1 U13488 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12317) );
  OR2_X1 U13489 ( .A1(n10600), .A2(n12317), .ZN(n10541) );
  OAI211_X1 U13490 ( .C1(n10654), .C2(n12451), .A(n10542), .B(n10541), .ZN(
        n10543) );
  NOR2_X1 U13491 ( .A1(n10544), .A2(n10543), .ZN(n10557) );
  INV_X1 U13492 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12452) );
  NOR2_X1 U13493 ( .A1(n10614), .A2(n12452), .ZN(n10555) );
  INV_X1 U13494 ( .A(n10546), .ZN(n10550) );
  INV_X1 U13495 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10553) );
  AOI21_X1 U13496 ( .B1(n20352), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n17076), .ZN(n10552) );
  AND3_X1 U13497 ( .A1(n12161), .A2(n10550), .A3(n10549), .ZN(n20424) );
  NAND2_X1 U13498 ( .A1(n20424), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10551) );
  OAI211_X1 U13499 ( .C1(n20023), .C2(n10553), .A(n10552), .B(n10551), .ZN(
        n10554) );
  NOR2_X1 U13500 ( .A1(n10555), .A2(n10554), .ZN(n10556) );
  AOI22_X1 U13501 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12433), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13502 ( .A1(n12202), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13503 ( .A1(n12384), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12368), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13504 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10561) );
  NAND4_X1 U13505 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n10571) );
  AOI22_X1 U13506 ( .A1(n12366), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12389), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13507 ( .A1(n10277), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13508 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12424), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13509 ( .A1(n12423), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12351), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10566) );
  NAND4_X1 U13510 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10570) );
  NOR2_X1 U13511 ( .A1(n10571), .A2(n10570), .ZN(n12644) );
  OR2_X1 U13512 ( .A1(n12644), .A2(n17047), .ZN(n15930) );
  INV_X1 U13513 ( .A(n15930), .ZN(n10572) );
  NAND2_X1 U13514 ( .A1(n10572), .A2(n12655), .ZN(n10813) );
  NAND2_X1 U13515 ( .A1(n10813), .A2(n12665), .ZN(n10574) );
  INV_X1 U13516 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10575) );
  INV_X1 U13517 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12504) );
  INV_X1 U13518 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10576) );
  OAI22_X1 U13519 ( .A1(n10609), .A2(n12504), .B1(n10610), .B2(n10576), .ZN(
        n10577) );
  NOR2_X1 U13520 ( .A1(n10578), .A2(n10577), .ZN(n10591) );
  INV_X1 U13521 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10579) );
  INV_X1 U13522 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12495) );
  INV_X1 U13523 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10581) );
  INV_X1 U13524 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10580) );
  NOR2_X1 U13525 ( .A1(n10583), .A2(n10582), .ZN(n10590) );
  NAND2_X1 U13526 ( .A1(n10598), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10587) );
  INV_X1 U13527 ( .A(n10599), .ZN(n20083) );
  INV_X1 U13528 ( .A(n10600), .ZN(n20138) );
  NAND2_X1 U13529 ( .A1(n10597), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10585) );
  AOI22_X1 U13530 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20424), .B1(
        n20352), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13531 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10664), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U13532 ( .A1(n12671), .A2(n17076), .ZN(n10592) );
  NAND2_X1 U13533 ( .A1(n10809), .A2(n12676), .ZN(n10624) );
  INV_X1 U13534 ( .A(n10624), .ZN(n10622) );
  INV_X1 U13535 ( .A(n10593), .ZN(n13861) );
  INV_X1 U13536 ( .A(n10594), .ZN(n10595) );
  AOI22_X1 U13537 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n13861), .B1(
        n10595), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10608) );
  INV_X1 U13538 ( .A(n10596), .ZN(n20197) );
  INV_X1 U13539 ( .A(n10645), .ZN(n16228) );
  AOI22_X1 U13540 ( .A1(n20197), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16228), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13541 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n10597), .B1(
        n10598), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10606) );
  INV_X1 U13542 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12550) );
  INV_X1 U13543 ( .A(n20352), .ZN(n10656) );
  INV_X1 U13544 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12560) );
  OAI22_X1 U13545 ( .A1(n10599), .A2(n12550), .B1(n10656), .B2(n12560), .ZN(
        n10604) );
  INV_X1 U13546 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10602) );
  INV_X1 U13547 ( .A(n20424), .ZN(n10659) );
  OAI22_X1 U13548 ( .A1(n10600), .A2(n10602), .B1(n10659), .B2(n10601), .ZN(
        n10603) );
  NOR2_X1 U13549 ( .A1(n10604), .A2(n10603), .ZN(n10605) );
  NAND4_X1 U13550 ( .A1(n10608), .A2(n10607), .A3(n10606), .A4(n10605), .ZN(
        n10620) );
  INV_X1 U13551 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12556) );
  INV_X1 U13552 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10611) );
  OAI22_X1 U13553 ( .A1(n10609), .A2(n12556), .B1(n10610), .B2(n10611), .ZN(
        n10612) );
  INV_X1 U13554 ( .A(n10612), .ZN(n10618) );
  INV_X1 U13555 ( .A(n20023), .ZN(n20026) );
  AOI22_X1 U13556 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n20026), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10617) );
  INV_X1 U13557 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12549) );
  INV_X1 U13558 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12559) );
  NAND4_X1 U13559 ( .A1(n10618), .A2(n10617), .A3(n10616), .A4(n10615), .ZN(
        n10619) );
  INV_X1 U13560 ( .A(n10623), .ZN(n10621) );
  NAND2_X1 U13561 ( .A1(n10624), .A2(n10623), .ZN(n10625) );
  XNOR2_X1 U13562 ( .A(n10627), .B(n10626), .ZN(n19722) );
  INV_X1 U13563 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14023) );
  XNOR2_X1 U13564 ( .A(n10642), .B(n14023), .ZN(n14011) );
  NAND2_X1 U13565 ( .A1(n10631), .A2(n10630), .ZN(n10632) );
  NAND2_X1 U13566 ( .A1(n9909), .A2(n10632), .ZN(n14109) );
  INV_X1 U13567 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14480) );
  OAI21_X1 U13568 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20615), .A(
        n10802), .ZN(n10799) );
  MUX2_X1 U13569 ( .A(n10799), .B(n12644), .S(n10172), .Z(n10790) );
  MUX2_X1 U13570 ( .A(n10790), .B(n15507), .S(n10773), .Z(n15926) );
  INV_X1 U13571 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12803) );
  NOR2_X1 U13572 ( .A1(n15926), .A2(n12803), .ZN(n12997) );
  AND3_X1 U13573 ( .A1(n10773), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10633) );
  NOR2_X1 U13574 ( .A1(n10635), .A2(n10633), .ZN(n14078) );
  NAND2_X1 U13575 ( .A1(n12997), .A2(n14078), .ZN(n12996) );
  NOR2_X1 U13576 ( .A1(n12997), .A2(n14078), .ZN(n10634) );
  AOI21_X1 U13577 ( .B1(n14480), .B2(n12996), .A(n10634), .ZN(n14440) );
  XNOR2_X1 U13578 ( .A(n10636), .B(n10635), .ZN(n14122) );
  XNOR2_X1 U13579 ( .A(n14122), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14441) );
  INV_X1 U13580 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19925) );
  NOR2_X1 U13581 ( .A1(n14122), .A2(n19925), .ZN(n10637) );
  AOI21_X1 U13582 ( .B1(n14440), .B2(n14441), .A(n10637), .ZN(n13722) );
  XNOR2_X1 U13583 ( .A(n10639), .B(n10638), .ZN(n10640) );
  INV_X1 U13584 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19906) );
  XNOR2_X1 U13585 ( .A(n10640), .B(n19906), .ZN(n13996) );
  INV_X1 U13586 ( .A(n10640), .ZN(n19733) );
  NAND2_X1 U13587 ( .A1(n19733), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10641) );
  NAND2_X1 U13588 ( .A1(n13999), .A2(n10641), .ZN(n14010) );
  NAND2_X1 U13589 ( .A1(n14011), .A2(n14010), .ZN(n14009) );
  NAND2_X1 U13590 ( .A1(n10642), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10643) );
  NAND2_X1 U13591 ( .A1(n14009), .A2(n10643), .ZN(n16191) );
  INV_X1 U13592 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10644) );
  INV_X1 U13593 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12569) );
  OAI22_X1 U13594 ( .A1(n10644), .A2(n20023), .B1(n10594), .B2(n12569), .ZN(
        n10648) );
  INV_X1 U13595 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10646) );
  OAI22_X1 U13596 ( .A1(n10646), .A2(n10593), .B1(n10645), .B2(n19970), .ZN(
        n10647) );
  NOR2_X1 U13597 ( .A1(n10648), .A2(n10647), .ZN(n10669) );
  INV_X1 U13598 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12393) );
  INV_X1 U13599 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12582) );
  OAI22_X1 U13600 ( .A1(n10596), .A2(n12393), .B1(n10610), .B2(n12582), .ZN(
        n10652) );
  INV_X1 U13601 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12580) );
  INV_X1 U13602 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10649) );
  OAI22_X1 U13603 ( .A1(n10609), .A2(n12580), .B1(n10650), .B2(n10649), .ZN(
        n10651) );
  NOR2_X1 U13604 ( .A1(n10652), .A2(n10651), .ZN(n10668) );
  INV_X1 U13605 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12396) );
  INV_X1 U13606 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10653) );
  OAI22_X1 U13607 ( .A1(n12396), .A2(n10655), .B1(n10654), .B2(n10653), .ZN(
        n10663) );
  INV_X1 U13608 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10657) );
  INV_X1 U13609 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12578) );
  OAI22_X1 U13610 ( .A1(n10600), .A2(n10657), .B1(n10656), .B2(n12578), .ZN(
        n10661) );
  INV_X1 U13611 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12570) );
  OAI22_X1 U13612 ( .A1(n10599), .A2(n12570), .B1(n10659), .B2(n10658), .ZN(
        n10660) );
  OR2_X1 U13613 ( .A1(n10661), .A2(n10660), .ZN(n10662) );
  NOR2_X1 U13614 ( .A1(n10663), .A2(n10662), .ZN(n10667) );
  AOI22_X1 U13615 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10664), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10666) );
  NAND4_X1 U13616 ( .A1(n10669), .A2(n10668), .A3(n10667), .A4(n10666), .ZN(
        n10672) );
  INV_X1 U13617 ( .A(n12687), .ZN(n10670) );
  NAND2_X1 U13618 ( .A1(n10670), .A2(n17076), .ZN(n10671) );
  XNOR2_X1 U13619 ( .A(n10674), .B(n10673), .ZN(n19712) );
  NAND2_X1 U13620 ( .A1(n10675), .A2(n19712), .ZN(n10676) );
  INV_X1 U13621 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14471) );
  XNOR2_X1 U13622 ( .A(n10676), .B(n14471), .ZN(n16190) );
  NAND2_X1 U13623 ( .A1(n10676), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10677) );
  INV_X1 U13624 ( .A(n10678), .ZN(n10679) );
  XNOR2_X1 U13625 ( .A(n10680), .B(n10679), .ZN(n19700) );
  AND2_X1 U13626 ( .A1(n19700), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15906) );
  INV_X1 U13627 ( .A(n19700), .ZN(n10681) );
  INV_X1 U13628 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10835) );
  NAND2_X1 U13629 ( .A1(n10681), .A2(n10835), .ZN(n15905) );
  INV_X1 U13630 ( .A(n10684), .ZN(n10685) );
  XNOR2_X1 U13631 ( .A(n10686), .B(n10685), .ZN(n14053) );
  AND2_X1 U13632 ( .A1(n14053), .A2(n10350), .ZN(n15893) );
  INV_X1 U13633 ( .A(n10695), .ZN(n10691) );
  NAND2_X1 U13634 ( .A1(n10773), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10689) );
  MUX2_X1 U13635 ( .A(n10689), .B(n10773), .S(n10688), .Z(n10690) );
  AOI21_X1 U13636 ( .B1(n19682), .B2(n10350), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16160) );
  NOR2_X1 U13637 ( .A1(n10695), .A2(n19783), .ZN(n10692) );
  NAND2_X1 U13638 ( .A1(n10773), .A2(n10692), .ZN(n10693) );
  NAND2_X1 U13639 ( .A1(n14414), .A2(n10693), .ZN(n10694) );
  AOI21_X1 U13640 ( .B1(n10695), .B2(n19783), .A(n10694), .ZN(n19675) );
  INV_X1 U13641 ( .A(n19675), .ZN(n10696) );
  INV_X1 U13642 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16151) );
  OAI21_X1 U13643 ( .B1(n10696), .B2(n10362), .A(n16151), .ZN(n15875) );
  AND3_X1 U13644 ( .A1(n19675), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n10350), .ZN(n15874) );
  AND2_X1 U13645 ( .A1(n10350), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10697) );
  NAND3_X1 U13646 ( .A1(n10773), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10699), 
        .ZN(n10700) );
  NAND2_X1 U13647 ( .A1(n10701), .A2(n10700), .ZN(n14045) );
  NOR2_X1 U13648 ( .A1(n14045), .A2(n10362), .ZN(n10735) );
  NAND2_X1 U13649 ( .A1(n10735), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16142) );
  NAND2_X1 U13650 ( .A1(n9918), .A2(n10703), .ZN(n10704) );
  NAND2_X1 U13651 ( .A1(n10731), .A2(n10704), .ZN(n15502) );
  INV_X1 U13652 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16133) );
  XNOR2_X1 U13653 ( .A(n10738), .B(n16133), .ZN(n15862) );
  NAND2_X1 U13654 ( .A1(n10773), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10705) );
  MUX2_X1 U13655 ( .A(n10773), .B(n10705), .S(n10712), .Z(n10706) );
  NAND2_X1 U13656 ( .A1(n10706), .A2(n9657), .ZN(n15445) );
  INV_X1 U13657 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16075) );
  OAI21_X1 U13658 ( .B1(n15445), .B2(n10362), .A(n16075), .ZN(n15763) );
  NAND2_X1 U13659 ( .A1(n10773), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10707) );
  INV_X1 U13660 ( .A(n10708), .ZN(n10719) );
  MUX2_X1 U13661 ( .A(n10773), .B(n10707), .S(n10719), .Z(n10709) );
  INV_X1 U13662 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n16913) );
  NAND2_X1 U13663 ( .A1(n10708), .A2(n16913), .ZN(n10711) );
  NAND2_X1 U13664 ( .A1(n15446), .A2(n10350), .ZN(n10710) );
  INV_X1 U13665 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15791) );
  NAND2_X1 U13666 ( .A1(n10710), .A2(n15791), .ZN(n15787) );
  NAND3_X1 U13667 ( .A1(n10711), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n10773), 
        .ZN(n10713) );
  NAND2_X1 U13668 ( .A1(n10713), .A2(n10712), .ZN(n19623) );
  INV_X1 U13669 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16088) );
  NAND2_X1 U13670 ( .A1(n10749), .A2(n16088), .ZN(n15775) );
  NAND2_X1 U13671 ( .A1(n15763), .A2(n15762), .ZN(n15751) );
  NAND3_X1 U13672 ( .A1(n9657), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n10773), .ZN(
        n10714) );
  AND2_X1 U13673 ( .A1(n10715), .A2(n10714), .ZN(n10747) );
  AOI21_X1 U13674 ( .B1(n10747), .B2(n10350), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15753) );
  INV_X1 U13675 ( .A(n10716), .ZN(n10718) );
  NAND2_X1 U13676 ( .A1(n10718), .A2(n9914), .ZN(n10720) );
  NAND2_X1 U13677 ( .A1(n19649), .A2(n10350), .ZN(n10721) );
  INV_X1 U13678 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15809) );
  NAND2_X1 U13679 ( .A1(n10721), .A2(n15809), .ZN(n15799) );
  AND2_X1 U13680 ( .A1(n10773), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10723) );
  INV_X1 U13681 ( .A(n14414), .ZN(n10722) );
  AOI21_X1 U13682 ( .B1(n10724), .B2(n10723), .A(n10722), .ZN(n10726) );
  AND2_X1 U13683 ( .A1(n10726), .A2(n10725), .ZN(n15462) );
  NAND2_X1 U13684 ( .A1(n15462), .A2(n10350), .ZN(n10752) );
  XNOR2_X1 U13685 ( .A(n10752), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15817) );
  INV_X1 U13686 ( .A(n10727), .ZN(n10728) );
  XNOR2_X1 U13687 ( .A(n10733), .B(n10728), .ZN(n15485) );
  NAND2_X1 U13688 ( .A1(n15485), .A2(n10350), .ZN(n10729) );
  INV_X1 U13689 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21218) );
  NAND2_X1 U13690 ( .A1(n10729), .A2(n21218), .ZN(n15838) );
  NAND2_X1 U13691 ( .A1(n10731), .A2(n10730), .ZN(n10732) );
  NAND2_X1 U13692 ( .A1(n10733), .A2(n10732), .ZN(n12840) );
  INV_X1 U13693 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10734) );
  OAI21_X1 U13694 ( .B1(n12840), .B2(n10362), .A(n10734), .ZN(n15852) );
  INV_X1 U13695 ( .A(n10735), .ZN(n10737) );
  INV_X1 U13696 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10736) );
  NAND2_X1 U13697 ( .A1(n10737), .A2(n10736), .ZN(n16141) );
  NAND2_X1 U13698 ( .A1(n10738), .A2(n16133), .ZN(n15743) );
  AND4_X1 U13699 ( .A1(n15838), .A2(n15852), .A3(n16141), .A4(n15743), .ZN(
        n10741) );
  XNOR2_X1 U13700 ( .A(n9664), .B(n10739), .ZN(n19668) );
  NAND2_X1 U13701 ( .A1(n19668), .A2(n10350), .ZN(n10740) );
  INV_X1 U13702 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16968) );
  NAND2_X1 U13703 ( .A1(n10740), .A2(n16968), .ZN(n15826) );
  NAND4_X1 U13704 ( .A1(n15799), .A2(n15817), .A3(n10741), .A4(n15826), .ZN(
        n10742) );
  OR2_X1 U13705 ( .A1(n15753), .A2(n10742), .ZN(n10743) );
  INV_X1 U13706 ( .A(n15445), .ZN(n10746) );
  AND2_X1 U13707 ( .A1(n10350), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10745) );
  INV_X1 U13708 ( .A(n10747), .ZN(n15430) );
  NAND2_X1 U13709 ( .A1(n10350), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10748) );
  NOR2_X1 U13710 ( .A1(n15430), .A2(n10748), .ZN(n15752) );
  INV_X1 U13711 ( .A(n10749), .ZN(n10750) );
  NAND2_X1 U13712 ( .A1(n10750), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15776) );
  AND2_X1 U13713 ( .A1(n10350), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10751) );
  NAND2_X1 U13714 ( .A1(n19649), .A2(n10751), .ZN(n15798) );
  INV_X1 U13715 ( .A(n10752), .ZN(n10753) );
  NAND2_X1 U13716 ( .A1(n10753), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15801) );
  NAND2_X1 U13717 ( .A1(n15798), .A2(n15801), .ZN(n15748) );
  INV_X1 U13718 ( .A(n19668), .ZN(n10754) );
  AND2_X1 U13719 ( .A1(n10350), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10755) );
  NAND2_X1 U13720 ( .A1(n15485), .A2(n10755), .ZN(n15837) );
  INV_X1 U13721 ( .A(n12840), .ZN(n10757) );
  AND2_X1 U13722 ( .A1(n10350), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10756) );
  NAND2_X1 U13723 ( .A1(n10757), .A2(n10756), .ZN(n15851) );
  NAND3_X1 U13724 ( .A1(n15825), .A2(n15837), .A3(n15851), .ZN(n10758) );
  NOR2_X1 U13725 ( .A1(n15748), .A2(n10758), .ZN(n10760) );
  AND2_X1 U13726 ( .A1(n10350), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10759) );
  NAND2_X1 U13727 ( .A1(n15446), .A2(n10759), .ZN(n15786) );
  INV_X1 U13728 ( .A(n10762), .ZN(n10765) );
  AOI21_X1 U13729 ( .B1(n10765), .B2(n10764), .A(n10763), .ZN(n16486) );
  AOI21_X1 U13730 ( .B1(n16486), .B2(n10350), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15730) );
  NAND3_X1 U13731 ( .A1(n16486), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n10350), .ZN(n15731) );
  NAND2_X1 U13732 ( .A1(n10767), .A2(n10766), .ZN(n10768) );
  NAND2_X1 U13733 ( .A1(n16884), .A2(n10768), .ZN(n15414) );
  NOR2_X1 U13734 ( .A1(n15414), .A2(n10362), .ZN(n10769) );
  XOR2_X1 U13735 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n10769), .Z(
        n15722) );
  INV_X1 U13736 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16028) );
  NOR3_X1 U13737 ( .A1(n15414), .A2(n10362), .A3(n16028), .ZN(n10770) );
  AND2_X1 U13738 ( .A1(n14414), .A2(n10350), .ZN(n15714) );
  INV_X1 U13739 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21106) );
  INV_X1 U13740 ( .A(n15714), .ZN(n10782) );
  INV_X1 U13741 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15998) );
  NAND2_X1 U13742 ( .A1(n10782), .A2(n15998), .ZN(n15705) );
  AND2_X1 U13743 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n16871), .ZN(n10772) );
  AOI21_X1 U13744 ( .B1(n10773), .B2(n10772), .A(n10771), .ZN(n10774) );
  NAND2_X1 U13745 ( .A1(n14414), .A2(n10774), .ZN(n16854) );
  INV_X1 U13746 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15999) );
  INV_X1 U13747 ( .A(n16854), .ZN(n10775) );
  INV_X1 U13748 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15954) );
  INV_X1 U13749 ( .A(n10776), .ZN(n10777) );
  NAND2_X1 U13750 ( .A1(n10778), .A2(n10777), .ZN(n10779) );
  NAND2_X1 U13751 ( .A1(n14410), .A2(n10779), .ZN(n15383) );
  AOI21_X1 U13752 ( .B1(n15954), .B2(n15970), .A(n15679), .ZN(n10780) );
  NOR2_X1 U13753 ( .A1(n10782), .A2(n15998), .ZN(n15706) );
  NOR2_X1 U13754 ( .A1(n10783), .A2(n15706), .ZN(n15674) );
  XOR2_X1 U13755 ( .A(n10784), .B(n14407), .Z(n15964) );
  NOR2_X1 U13756 ( .A1(n17068), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10785) );
  INV_X1 U13757 ( .A(n10951), .ZN(n10948) );
  INV_X1 U13758 ( .A(n10939), .ZN(n10789) );
  INV_X1 U13759 ( .A(n10787), .ZN(n10788) );
  OAI21_X1 U13760 ( .B1(n10790), .B2(n10789), .A(n10788), .ZN(n10794) );
  INV_X1 U13761 ( .A(n10791), .ZN(n10793) );
  NAND3_X1 U13762 ( .A1(n10794), .A2(n10793), .A3(n10792), .ZN(n10795) );
  NAND2_X1 U13763 ( .A1(n10948), .A2(n10795), .ZN(n20622) );
  AND2_X1 U13764 ( .A1(n17076), .A2(n19936), .ZN(n12617) );
  INV_X1 U13765 ( .A(n12617), .ZN(n10796) );
  OR2_X1 U13766 ( .A1(n17046), .A2(n10796), .ZN(n13727) );
  NAND2_X1 U13767 ( .A1(n17060), .A2(n10797), .ZN(n12878) );
  OR2_X1 U13768 ( .A1(n12365), .A2(n12878), .ZN(n10798) );
  INV_X1 U13769 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12874) );
  NAND2_X1 U13770 ( .A1(n10798), .A2(n12874), .ZN(n20611) );
  INV_X1 U13771 ( .A(n10799), .ZN(n10938) );
  NAND2_X1 U13772 ( .A1(n10801), .A2(n10800), .ZN(n10945) );
  NOR2_X1 U13773 ( .A1(n10936), .A2(n10945), .ZN(n10804) );
  XNOR2_X1 U13774 ( .A(n10939), .B(n10802), .ZN(n10934) );
  AND2_X1 U13775 ( .A1(n10934), .A2(n10804), .ZN(n10803) );
  OR2_X1 U13776 ( .A1(n10951), .A2(n10803), .ZN(n17050) );
  AOI21_X1 U13777 ( .B1(n10938), .B2(n10804), .A(n17050), .ZN(n10805) );
  MUX2_X1 U13778 ( .A(n20611), .B(n10805), .S(n20495), .Z(n16555) );
  NAND2_X1 U13779 ( .A1(n16555), .A2(n17047), .ZN(n10806) );
  OAI22_X1 U13780 ( .A1(n20622), .A2(n13727), .B1(n17046), .B2(n10806), .ZN(
        n13712) );
  NAND2_X1 U13781 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20495), .ZN(n20494) );
  INV_X1 U13782 ( .A(n20494), .ZN(n10807) );
  AND2_X1 U13783 ( .A1(n19936), .A2(n17073), .ZN(n10808) );
  NAND2_X1 U13784 ( .A1(n13712), .A2(n10808), .ZN(n12860) );
  OR2_X2 U13785 ( .A1(n12860), .A2(n17076), .ZN(n16957) );
  INV_X1 U13786 ( .A(n10809), .ZN(n10810) );
  AND2_X1 U13787 ( .A1(n15930), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15932) );
  XNOR2_X1 U13788 ( .A(n12644), .B(n12655), .ZN(n10811) );
  NAND2_X1 U13789 ( .A1(n15932), .A2(n10811), .ZN(n10812) );
  XOR2_X1 U13790 ( .A(n10811), .B(n15932), .Z(n13000) );
  NAND2_X1 U13791 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13000), .ZN(
        n12999) );
  NAND2_X1 U13792 ( .A1(n10812), .A2(n12999), .ZN(n10814) );
  XNOR2_X1 U13793 ( .A(n19925), .B(n10814), .ZN(n14436) );
  XNOR2_X1 U13794 ( .A(n12665), .B(n10813), .ZN(n14435) );
  NAND2_X1 U13795 ( .A1(n14436), .A2(n14435), .ZN(n14434) );
  NAND2_X1 U13796 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10814), .ZN(
        n10815) );
  NAND2_X1 U13797 ( .A1(n14434), .A2(n10815), .ZN(n10816) );
  XNOR2_X1 U13798 ( .A(n10816), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13726) );
  NAND2_X1 U13799 ( .A1(n10816), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10817) );
  OAI21_X1 U13800 ( .B1(n13993), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13994), .ZN(n10820) );
  NAND2_X1 U13801 ( .A1(n13993), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10819) );
  NAND2_X1 U13802 ( .A1(n10820), .A2(n10819), .ZN(n14014) );
  NAND2_X1 U13803 ( .A1(n10821), .A2(n14023), .ZN(n14013) );
  INV_X1 U13804 ( .A(n14017), .ZN(n10824) );
  NAND2_X1 U13805 ( .A1(n10824), .A2(n10831), .ZN(n10826) );
  NAND2_X1 U13806 ( .A1(n16201), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16200) );
  NAND2_X1 U13807 ( .A1(n14012), .A2(n14017), .ZN(n10828) );
  NAND2_X1 U13808 ( .A1(n10828), .A2(n10827), .ZN(n10829) );
  INV_X1 U13809 ( .A(n10832), .ZN(n10833) );
  NAND2_X1 U13810 ( .A1(n10833), .A2(n10362), .ZN(n10834) );
  NAND2_X1 U13811 ( .A1(n10838), .A2(n10834), .ZN(n15912) );
  XNOR2_X1 U13812 ( .A(n10838), .B(n10683), .ZN(n15899) );
  INV_X1 U13813 ( .A(n15899), .ZN(n10836) );
  INV_X1 U13814 ( .A(n10838), .ZN(n10839) );
  NAND2_X1 U13815 ( .A1(n10839), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10840) );
  NAND2_X1 U13816 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16491) );
  NOR2_X1 U13817 ( .A1(n16151), .A2(n10736), .ZN(n16150) );
  NAND2_X1 U13818 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16150), .ZN(
        n16120) );
  INV_X1 U13819 ( .A(n16120), .ZN(n10841) );
  NAND2_X1 U13820 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16978) );
  NOR2_X1 U13821 ( .A1(n21218), .A2(n16978), .ZN(n16977) );
  NAND2_X1 U13822 ( .A1(n10841), .A2(n16977), .ZN(n16108) );
  INV_X1 U13823 ( .A(n16108), .ZN(n15806) );
  NAND2_X1 U13824 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n15806), .ZN(
        n10842) );
  NOR2_X1 U13825 ( .A1(n16491), .A2(n10842), .ZN(n16096) );
  AND2_X1 U13826 ( .A1(n16096), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16055) );
  NAND2_X1 U13827 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16027) );
  INV_X1 U13828 ( .A(n16027), .ZN(n10843) );
  OAI21_X1 U13829 ( .B1(n15683), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15668), .ZN(n15951) );
  INV_X1 U13830 ( .A(n12860), .ZN(n10845) );
  NOR2_X1 U13831 ( .A1(n15951), .A2(n16955), .ZN(n10965) );
  INV_X1 U13832 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n10846) );
  INV_X1 U13833 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16949) );
  OAI22_X1 U13834 ( .A1(n9609), .A2(n10846), .B1(n20495), .B2(n16949), .ZN(
        n10848) );
  INV_X1 U13835 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16174) );
  NOR2_X1 U13836 ( .A1(n14426), .A2(n16174), .ZN(n10847) );
  AOI211_X1 U13837 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n14424), .A(n10848), .B(
        n10847), .ZN(n13365) );
  NAND2_X1 U13838 ( .A1(n10851), .A2(n10850), .ZN(n10854) );
  INV_X1 U13839 ( .A(n10852), .ZN(n10853) );
  OR2_X1 U13840 ( .A1(n10500), .A2(n19906), .ZN(n10857) );
  INV_X1 U13841 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n14003) );
  OAI22_X1 U13842 ( .A1(n14422), .A2(n14003), .B1(n20495), .B2(n14004), .ZN(
        n10855) );
  AOI21_X1 U13843 ( .B1(n14424), .B2(P2_EBX_REG_4__SCAN_IN), .A(n10855), .ZN(
        n10856) );
  NAND2_X1 U13844 ( .A1(n10857), .A2(n10856), .ZN(n14000) );
  NAND2_X1 U13845 ( .A1(n14001), .A2(n14000), .ZN(n13101) );
  OR2_X1 U13846 ( .A1(n10500), .A2(n14023), .ZN(n10860) );
  INV_X1 U13847 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n14024) );
  INV_X1 U13848 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15918) );
  OAI22_X1 U13849 ( .A1(n14422), .A2(n14024), .B1(n20495), .B2(n15918), .ZN(
        n10858) );
  AOI21_X1 U13850 ( .B1(n14424), .B2(P2_EBX_REG_5__SCAN_IN), .A(n10858), .ZN(
        n10859) );
  OR2_X1 U13851 ( .A1(n14426), .A2(n14471), .ZN(n10864) );
  INV_X1 U13852 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n10861) );
  OAI22_X1 U13853 ( .A1(n9609), .A2(n10861), .B1(n20495), .B2(n12809), .ZN(
        n10862) );
  AOI21_X1 U13854 ( .B1(n14424), .B2(P2_EBX_REG_6__SCAN_IN), .A(n10862), .ZN(
        n10863) );
  NAND2_X1 U13855 ( .A1(n10864), .A2(n10863), .ZN(n13190) );
  OR2_X1 U13856 ( .A1(n10500), .A2(n10835), .ZN(n10868) );
  INV_X1 U13857 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10865) );
  OAI22_X1 U13858 ( .A1(n9609), .A2(n10865), .B1(n20495), .B2(n15909), .ZN(
        n10866) );
  AOI21_X1 U13859 ( .B1(n14424), .B2(P2_EBX_REG_7__SCAN_IN), .A(n10866), .ZN(
        n10867) );
  NAND2_X1 U13860 ( .A1(n10868), .A2(n10867), .ZN(n13243) );
  OR2_X1 U13861 ( .A1(n10500), .A2(n10683), .ZN(n10872) );
  INV_X1 U13862 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12689) );
  INV_X1 U13863 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10869) );
  OAI22_X1 U13864 ( .A1(n9609), .A2(n12689), .B1(n20495), .B2(n10869), .ZN(
        n10870) );
  AOI21_X1 U13865 ( .B1(n14424), .B2(P2_EBX_REG_8__SCAN_IN), .A(n10870), .ZN(
        n10871) );
  NAND2_X1 U13866 ( .A1(n10872), .A2(n10871), .ZN(n14051) );
  OR2_X1 U13867 ( .A1(n14426), .A2(n16151), .ZN(n10875) );
  INV_X1 U13868 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n15879) );
  OAI22_X1 U13869 ( .A1(n9609), .A2(n15879), .B1(n20495), .B2(n15880), .ZN(
        n10873) );
  AOI21_X1 U13870 ( .B1(n14424), .B2(P2_EBX_REG_10__SCAN_IN), .A(n10873), .ZN(
        n10874) );
  OR2_X1 U13871 ( .A1(n14426), .A2(n10736), .ZN(n10878) );
  INV_X1 U13872 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12702) );
  OAI22_X1 U13873 ( .A1(n9609), .A2(n12702), .B1(n20495), .B2(n16941), .ZN(
        n10876) );
  AOI21_X1 U13874 ( .B1(n14424), .B2(P2_EBX_REG_11__SCAN_IN), .A(n10876), .ZN(
        n10877) );
  OR2_X1 U13875 ( .A1(n14426), .A2(n16133), .ZN(n10881) );
  INV_X1 U13876 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12705) );
  OAI22_X1 U13877 ( .A1(n9609), .A2(n12705), .B1(n20495), .B2(n15865), .ZN(
        n10879) );
  AOI21_X1 U13878 ( .B1(n14424), .B2(P2_EBX_REG_12__SCAN_IN), .A(n10879), .ZN(
        n10880) );
  NAND2_X1 U13879 ( .A1(n10881), .A2(n10880), .ZN(n15497) );
  INV_X1 U13880 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U13881 ( .A1(n10882), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10883) );
  OAI21_X1 U13882 ( .B1(n9591), .B2(n10884), .A(n10883), .ZN(n10885) );
  AOI21_X1 U13883 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10885), .ZN(n12848) );
  OR2_X1 U13884 ( .A1(n14426), .A2(n21218), .ZN(n10888) );
  INV_X1 U13885 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n15842) );
  OAI22_X1 U13886 ( .A1(n9609), .A2(n15842), .B1(n20495), .B2(n15843), .ZN(
        n10886) );
  AOI21_X1 U13887 ( .B1(n14424), .B2(P2_EBX_REG_14__SCAN_IN), .A(n10886), .ZN(
        n10887) );
  NAND2_X1 U13888 ( .A1(n10888), .A2(n10887), .ZN(n15482) );
  OR2_X1 U13889 ( .A1(n14426), .A2(n16968), .ZN(n10892) );
  INV_X1 U13890 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n10889) );
  OAI22_X1 U13891 ( .A1(n9609), .A2(n10889), .B1(n20495), .B2(n19655), .ZN(
        n10890) );
  AOI21_X1 U13892 ( .B1(n14424), .B2(P2_EBX_REG_15__SCAN_IN), .A(n10890), .ZN(
        n10891) );
  INV_X1 U13893 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16498) );
  OR2_X1 U13894 ( .A1(n14426), .A2(n16498), .ZN(n10895) );
  INV_X1 U13895 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n12720) );
  INV_X1 U13896 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15819) );
  OAI22_X1 U13897 ( .A1(n9609), .A2(n12720), .B1(n20495), .B2(n15819), .ZN(
        n10893) );
  AOI21_X1 U13898 ( .B1(n14424), .B2(P2_EBX_REG_16__SCAN_IN), .A(n10893), .ZN(
        n10894) );
  NAND2_X1 U13899 ( .A1(n10895), .A2(n10894), .ZN(n15468) );
  INV_X1 U13900 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13901 ( .A1(n10882), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10896) );
  OAI21_X1 U13902 ( .B1(n9591), .B2(n10897), .A(n10896), .ZN(n10898) );
  AOI21_X1 U13903 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10898), .ZN(n15576) );
  AOI22_X1 U13904 ( .A1(n10882), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10899) );
  OAI21_X1 U13905 ( .B1(n9591), .B2(n16913), .A(n10899), .ZN(n10900) );
  AOI21_X1 U13906 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10900), .ZN(n15450) );
  INV_X1 U13907 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13908 ( .A1(n10882), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10901) );
  OAI21_X1 U13909 ( .B1(n9591), .B2(n10902), .A(n10901), .ZN(n10903) );
  AOI21_X1 U13910 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10903), .ZN(n15570) );
  OR2_X1 U13911 ( .A1(n14426), .A2(n16075), .ZN(n10907) );
  INV_X1 U13912 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15768) );
  INV_X1 U13913 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10904) );
  OAI22_X1 U13914 ( .A1(n9609), .A2(n15768), .B1(n20495), .B2(n10904), .ZN(
        n10905) );
  AOI21_X1 U13915 ( .B1(n14424), .B2(P2_EBX_REG_20__SCAN_IN), .A(n10905), .ZN(
        n10906) );
  NAND2_X1 U13916 ( .A1(n10907), .A2(n10906), .ZN(n15435) );
  AOI22_X1 U13917 ( .A1(n10882), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10908) );
  OAI21_X1 U13918 ( .B1(n9591), .B2(n15564), .A(n10908), .ZN(n10909) );
  AOI21_X1 U13919 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10909), .ZN(n15420) );
  INV_X1 U13920 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16478) );
  AOI22_X1 U13921 ( .A1(n10882), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10910) );
  OAI21_X1 U13922 ( .B1(n9591), .B2(n16478), .A(n10910), .ZN(n10911) );
  AOI21_X1 U13923 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10911), .ZN(n15735) );
  OR2_X1 U13924 ( .A1(n14426), .A2(n16028), .ZN(n10914) );
  INV_X1 U13925 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20542) );
  INV_X1 U13926 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15408) );
  OAI22_X1 U13927 ( .A1(n9609), .A2(n20542), .B1(n20495), .B2(n15408), .ZN(
        n10912) );
  AOI21_X1 U13928 ( .B1(n14424), .B2(P2_EBX_REG_23__SCAN_IN), .A(n10912), .ZN(
        n10913) );
  NAND2_X1 U13929 ( .A1(n10914), .A2(n10913), .ZN(n15405) );
  INV_X1 U13930 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13931 ( .A1(n10882), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10915) );
  OAI21_X1 U13932 ( .B1(n9591), .B2(n10916), .A(n10915), .ZN(n10917) );
  AOI21_X1 U13933 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10917), .ZN(n15555) );
  OR2_X2 U13934 ( .A1(n15556), .A2(n15555), .ZN(n15558) );
  AOI22_X1 U13935 ( .A1(n10882), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10918) );
  OAI21_X1 U13936 ( .B1(n9591), .B2(n16877), .A(n10918), .ZN(n10919) );
  AOI21_X1 U13937 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10919), .ZN(n15546) );
  OR2_X1 U13938 ( .A1(n14426), .A2(n15999), .ZN(n10922) );
  INV_X1 U13939 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20548) );
  INV_X1 U13940 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15700) );
  OAI22_X1 U13941 ( .A1(n9609), .A2(n20548), .B1(n20495), .B2(n15700), .ZN(
        n10920) );
  AOI21_X1 U13942 ( .B1(n14424), .B2(P2_EBX_REG_26__SCAN_IN), .A(n10920), .ZN(
        n10921) );
  NAND2_X1 U13943 ( .A1(n10922), .A2(n10921), .ZN(n15538) );
  OR2_X1 U13944 ( .A1(n14426), .A2(n15970), .ZN(n10925) );
  INV_X1 U13945 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20551) );
  INV_X1 U13946 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15690) );
  OAI22_X1 U13947 ( .A1(n9609), .A2(n20551), .B1(n20495), .B2(n15690), .ZN(
        n10923) );
  AOI21_X1 U13948 ( .B1(n14424), .B2(P2_EBX_REG_27__SCAN_IN), .A(n10923), .ZN(
        n10924) );
  NAND2_X1 U13949 ( .A1(n10925), .A2(n10924), .ZN(n15388) );
  INV_X1 U13950 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13951 ( .A1(n10882), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10926) );
  OAI21_X1 U13952 ( .B1(n9591), .B2(n10927), .A(n10926), .ZN(n10928) );
  AOI21_X1 U13953 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10928), .ZN(n15373) );
  INV_X1 U13954 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U13955 ( .A1(n10882), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10929) );
  OAI21_X1 U13956 ( .B1(n9591), .B2(n15368), .A(n10929), .ZN(n10930) );
  AOI21_X1 U13957 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n10930), .ZN(n10931) );
  NAND2_X1 U13958 ( .A1(n9653), .A2(n10931), .ZN(n10932) );
  NAND2_X1 U13959 ( .A1(n14421), .A2(n10932), .ZN(n15960) );
  INV_X1 U13960 ( .A(n15960), .ZN(n10962) );
  NAND2_X1 U13961 ( .A1(n10950), .A2(n17047), .ZN(n10933) );
  MUX2_X1 U13962 ( .A(n13721), .B(n10933), .S(n10936), .Z(n10944) );
  OAI21_X1 U13963 ( .B1(n17047), .B2(n10938), .A(n10934), .ZN(n10935) );
  OAI21_X1 U13964 ( .B1(n17047), .B2(n10936), .A(n10935), .ZN(n10937) );
  NAND2_X1 U13965 ( .A1(n10937), .A2(n10451), .ZN(n10942) );
  NAND2_X1 U13966 ( .A1(n10939), .A2(n10938), .ZN(n10940) );
  NAND2_X1 U13967 ( .A1(n10172), .A2(n10940), .ZN(n10941) );
  NAND2_X1 U13968 ( .A1(n10942), .A2(n10941), .ZN(n10943) );
  NAND2_X1 U13969 ( .A1(n10944), .A2(n10943), .ZN(n10946) );
  MUX2_X1 U13970 ( .A(n10946), .B(n13721), .S(n10945), .Z(n10947) );
  NAND2_X1 U13971 ( .A1(n10948), .A2(n10947), .ZN(n10949) );
  MUX2_X1 U13972 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n10949), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n13708) );
  INV_X1 U13973 ( .A(n10950), .ZN(n12976) );
  NAND2_X1 U13974 ( .A1(n10951), .A2(n12976), .ZN(n10952) );
  NAND2_X1 U13975 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20606) );
  NOR2_X1 U13976 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17082) );
  INV_X1 U13977 ( .A(n17082), .ZN(n10954) );
  NAND2_X1 U13978 ( .A1(n20606), .A2(n10954), .ZN(n10955) );
  INV_X1 U13979 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15313) );
  INV_X1 U13980 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15734) );
  INV_X1 U13981 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15716) );
  OR2_X1 U13982 ( .A1(n10957), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10958) );
  NAND2_X1 U13983 ( .A1(n15337), .A2(n10958), .ZN(n15360) );
  NAND2_X1 U13984 ( .A1(n20495), .A2(n21204), .ZN(n20568) );
  INV_X1 U13985 ( .A(n20568), .ZN(n20579) );
  OR2_X1 U13986 ( .A1(n20585), .A2(n20579), .ZN(n20607) );
  NAND2_X1 U13987 ( .A1(n20607), .A2(n19598), .ZN(n10959) );
  INV_X1 U13988 ( .A(n12172), .ZN(n12157) );
  NAND2_X1 U13989 ( .A1(n21109), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12828) );
  NAND2_X1 U13990 ( .A1(n12157), .A2(n12828), .ZN(n15929) );
  NOR2_X1 U13991 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12829) );
  AND2_X2 U13992 ( .A1(n12829), .A2(n20579), .ZN(n19903) );
  INV_X2 U13993 ( .A(n19903), .ZN(n19736) );
  INV_X1 U13994 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20554) );
  NOR2_X1 U13995 ( .A1(n19736), .A2(n20554), .ZN(n15956) );
  AOI21_X1 U13996 ( .B1(n16954), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15956), .ZN(n10960) );
  OAI21_X1 U13997 ( .B1(n15360), .B2(n16952), .A(n10960), .ZN(n10961) );
  INV_X1 U13998 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13426) );
  NOR2_X2 U13999 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13141), .ZN(
        n10980) );
  NAND2_X1 U14000 ( .A1(n11175), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10968) );
  NAND2_X1 U14001 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10967) );
  OAI211_X1 U14002 ( .C1(n11816), .C2(n13426), .A(n10968), .B(n10967), .ZN(
        n10969) );
  INV_X1 U14003 ( .A(n10969), .ZN(n10989) );
  AOI22_X1 U14004 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11353), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10973) );
  NAND2_X1 U14005 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10972) );
  NAND2_X1 U14006 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10971) );
  NOR2_X4 U14007 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13156) );
  NAND2_X1 U14008 ( .A1(n11006), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10970) );
  NAND2_X1 U14009 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10978) );
  NAND2_X1 U14010 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10977) );
  NAND2_X1 U14011 ( .A1(n11074), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10976) );
  NAND2_X1 U14012 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10975) );
  NAND2_X1 U14013 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10985) );
  NAND2_X1 U14014 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10984) );
  NAND2_X1 U14015 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10983) );
  NAND2_X1 U14016 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10982) );
  AOI22_X1 U14017 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11175), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U14018 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U14019 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U14020 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11161), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10990) );
  NAND4_X1 U14021 ( .A1(n10993), .A2(n10992), .A3(n10991), .A4(n10990), .ZN(
        n11004) );
  INV_X1 U14022 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14023 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11001) );
  NAND2_X1 U14024 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11000) );
  NAND2_X1 U14025 ( .A1(n11056), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10998) );
  NAND2_X1 U14026 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10997) );
  NAND2_X1 U14027 ( .A1(n11006), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10996) );
  NAND2_X1 U14028 ( .A1(n11353), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10995) );
  NAND4_X1 U14029 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n11003) );
  INV_X1 U14030 ( .A(n11027), .ZN(n11116) );
  NAND2_X1 U14031 ( .A1(n13152), .A2(n11005), .ZN(n11787) );
  AOI22_X1 U14032 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11353), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11010) );
  NAND2_X1 U14033 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11009) );
  NAND2_X1 U14034 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11008) );
  NAND2_X1 U14035 ( .A1(n11006), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11007) );
  NAND2_X1 U14036 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11014) );
  NAND2_X1 U14037 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11013) );
  NAND2_X1 U14038 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11012) );
  NAND2_X1 U14039 ( .A1(n11074), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11011) );
  NAND2_X1 U14040 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11019) );
  NAND2_X1 U14041 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11018) );
  NAND2_X1 U14042 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11017) );
  NAND2_X1 U14043 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11016) );
  NAND2_X1 U14044 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11021) );
  NAND2_X1 U14045 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11020) );
  OAI211_X1 U14046 ( .C1(n11816), .C2(n13435), .A(n11021), .B(n11020), .ZN(
        n11022) );
  INV_X1 U14047 ( .A(n11022), .ZN(n11023) );
  NAND2_X1 U14048 ( .A1(n11125), .A2(n14970), .ZN(n11051) );
  NAND2_X1 U14049 ( .A1(n9614), .A2(n13301), .ZN(n11050) );
  AOI22_X1 U14050 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11353), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11032) );
  NAND2_X1 U14051 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11031) );
  NAND2_X1 U14052 ( .A1(n11006), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11030) );
  NAND2_X1 U14053 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11029) );
  NAND2_X1 U14054 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11036) );
  NAND2_X1 U14055 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11035) );
  NAND2_X1 U14056 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11034) );
  NAND2_X1 U14057 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11033) );
  NAND2_X1 U14058 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11041) );
  NAND2_X1 U14059 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11040) );
  NAND2_X1 U14060 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11039) );
  NAND2_X1 U14061 ( .A1(n11074), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11038) );
  INV_X1 U14062 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11044) );
  NAND2_X1 U14063 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11043) );
  NAND2_X1 U14064 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11042) );
  OAI211_X1 U14065 ( .C1(n11154), .C2(n11044), .A(n11043), .B(n11042), .ZN(
        n11045) );
  INV_X1 U14066 ( .A(n11045), .ZN(n11046) );
  NAND4_X4 U14067 ( .A1(n11049), .A2(n11048), .A3(n11047), .A4(n11046), .ZN(
        n13297) );
  AOI22_X1 U14068 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14069 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14070 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14071 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11052) );
  AOI22_X1 U14072 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9597), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11060) );
  NAND2_X1 U14073 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11059) );
  NAND2_X1 U14074 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11058) );
  NAND2_X1 U14075 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11057) );
  NAND4_X1 U14076 ( .A1(n11060), .A2(n11059), .A3(n11058), .A4(n11057), .ZN(
        n11064) );
  INV_X1 U14077 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13449) );
  NAND2_X1 U14078 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11062) );
  NAND2_X1 U14079 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11061) );
  OAI211_X1 U14080 ( .C1(n11816), .C2(n13449), .A(n11062), .B(n11061), .ZN(
        n11063) );
  NOR2_X1 U14081 ( .A1(n11064), .A2(n11063), .ZN(n11065) );
  INV_X1 U14082 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13438) );
  NAND2_X1 U14083 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11067) );
  NAND2_X1 U14084 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11066) );
  OAI211_X1 U14085 ( .C1(n11816), .C2(n13438), .A(n11067), .B(n11066), .ZN(
        n11068) );
  INV_X1 U14086 ( .A(n11068), .ZN(n11072) );
  AOI22_X1 U14087 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9597), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14088 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9603), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11070) );
  NAND2_X1 U14089 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11069) );
  NAND4_X1 U14090 ( .A1(n11072), .A2(n11071), .A3(n11070), .A4(n11069), .ZN(
        n11080) );
  AOI22_X1 U14091 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U14092 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14093 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14094 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11075) );
  NAND4_X1 U14095 ( .A1(n11078), .A2(n11077), .A3(n11076), .A4(n11075), .ZN(
        n11079) );
  NAND2_X1 U14096 ( .A1(n13297), .A2(n14977), .ZN(n11124) );
  NAND2_X1 U14097 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11083) );
  NAND2_X1 U14098 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11082) );
  NAND2_X1 U14099 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11081) );
  NAND2_X1 U14100 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11088) );
  NAND2_X1 U14101 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11087) );
  NAND2_X1 U14102 ( .A1(n11006), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11086) );
  NAND2_X1 U14103 ( .A1(n11074), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11085) );
  NAND2_X1 U14104 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11093) );
  NAND2_X1 U14105 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11092) );
  NAND2_X1 U14106 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11090) );
  NAND2_X1 U14107 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11095) );
  NAND2_X1 U14108 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11094) );
  OAI211_X1 U14109 ( .C1(n11816), .C2(n13443), .A(n11095), .B(n11094), .ZN(
        n11096) );
  INV_X1 U14110 ( .A(n11096), .ZN(n11097) );
  NAND4_X4 U14111 ( .A1(n11100), .A2(n11099), .A3(n11098), .A4(n11097), .ZN(
        n14957) );
  XNOR2_X1 U14112 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12962) );
  AOI22_X1 U14113 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14114 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14115 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11103) );
  AOI22_X1 U14116 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U14117 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11353), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11109) );
  NAND2_X1 U14118 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11108) );
  NAND2_X1 U14119 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11107) );
  NAND2_X1 U14120 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11106) );
  NAND4_X1 U14121 ( .A1(n11109), .A2(n11108), .A3(n11107), .A4(n11106), .ZN(
        n11113) );
  NAND2_X1 U14122 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11111) );
  NAND2_X1 U14123 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11110) );
  OAI211_X1 U14124 ( .C1(n11816), .C2(n13429), .A(n11111), .B(n11110), .ZN(
        n11112) );
  AND2_X4 U14125 ( .A1(n11115), .A2(n11114), .ZN(n11133) );
  NAND2_X1 U14126 ( .A1(n11133), .A2(n14957), .ZN(n16528) );
  INV_X1 U14127 ( .A(n13126), .ZN(n11118) );
  INV_X1 U14128 ( .A(n11133), .ZN(n11117) );
  NAND2_X1 U14129 ( .A1(n11118), .A2(n11143), .ZN(n13136) );
  NAND2_X1 U14130 ( .A1(n14982), .A2(n14978), .ZN(n13578) );
  NAND2_X1 U14131 ( .A1(n12965), .A2(n14957), .ZN(n13128) );
  INV_X1 U14132 ( .A(n11119), .ZN(n11120) );
  OAI211_X1 U14133 ( .C1(n14970), .C2(n13112), .A(n11121), .B(n11120), .ZN(
        n11122) );
  INV_X1 U14134 ( .A(n11122), .ZN(n11130) );
  INV_X1 U14135 ( .A(n11124), .ZN(n11126) );
  NAND2_X1 U14136 ( .A1(n11126), .A2(n11125), .ZN(n11531) );
  NAND2_X1 U14137 ( .A1(n11116), .A2(n13301), .ZN(n11127) );
  NOR2_X1 U14138 ( .A1(n13126), .A2(n14957), .ZN(n11131) );
  AND2_X2 U14139 ( .A1(n11132), .A2(n11131), .ZN(n13116) );
  INV_X1 U14140 ( .A(n12908), .ZN(n11134) );
  NAND2_X1 U14141 ( .A1(n11134), .A2(n14978), .ZN(n13071) );
  NAND2_X1 U14142 ( .A1(n20632), .A2(n20963), .ZN(n12150) );
  MUX2_X1 U14143 ( .A(n12150), .B(n16537), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11149) );
  AND2_X1 U14144 ( .A1(n11119), .A2(n14978), .ZN(n11136) );
  AOI21_X1 U14145 ( .B1(n11137), .B2(n13073), .A(n11136), .ZN(n13133) );
  INV_X1 U14146 ( .A(n13110), .ZN(n11138) );
  INV_X1 U14147 ( .A(n16528), .ZN(n12117) );
  NAND2_X1 U14148 ( .A1(n11138), .A2(n12117), .ZN(n11140) );
  OAI21_X1 U14149 ( .B1(n14982), .B2(n13309), .A(n13576), .ZN(n11139) );
  NAND4_X1 U14150 ( .A1(n11140), .A2(n20632), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n11139), .ZN(n11142) );
  NAND2_X1 U14151 ( .A1(n13127), .A2(n11255), .ZN(n11141) );
  NAND2_X1 U14152 ( .A1(n13136), .A2(n11141), .ZN(n14983) );
  NOR2_X1 U14153 ( .A1(n11142), .A2(n14983), .ZN(n11147) );
  AND2_X1 U14154 ( .A1(n13576), .A2(n14501), .ZN(n12995) );
  INV_X1 U14155 ( .A(n11125), .ZN(n13113) );
  NAND2_X1 U14156 ( .A1(n13113), .A2(n13288), .ZN(n11145) );
  INV_X1 U14157 ( .A(n13112), .ZN(n11144) );
  AOI22_X1 U14158 ( .A1(n12995), .A2(n11145), .B1(n11144), .B2(n11184), .ZN(
        n11146) );
  AND2_X1 U14159 ( .A1(n11147), .A2(n11146), .ZN(n11148) );
  INV_X1 U14160 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13624) );
  NAND2_X1 U14161 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11151) );
  NAND2_X1 U14162 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11150) );
  OAI211_X1 U14163 ( .C1(n11816), .C2(n13624), .A(n11151), .B(n11150), .ZN(
        n11152) );
  INV_X1 U14164 ( .A(n11152), .ZN(n11158) );
  AOI22_X1 U14165 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9613), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11157) );
  AOI22_X1 U14166 ( .A1(n11837), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11156) );
  NAND2_X1 U14167 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11155) );
  NAND4_X1 U14168 ( .A1(n11158), .A2(n11157), .A3(n11156), .A4(n11155), .ZN(
        n11167) );
  INV_X1 U14169 ( .A(n11159), .ZN(n11176) );
  AOI22_X1 U14170 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n11176), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U14171 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14172 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11161), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14173 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11162) );
  NAND4_X1 U14174 ( .A1(n11165), .A2(n11164), .A3(n11163), .A4(n11162), .ZN(
        n11166) );
  INV_X1 U14175 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13632) );
  INV_X2 U14176 ( .A(n11741), .ZN(n11865) );
  NAND2_X1 U14177 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11169) );
  NAND2_X1 U14178 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11168) );
  OAI211_X1 U14179 ( .C1(n11816), .C2(n13632), .A(n11169), .B(n11168), .ZN(
        n11170) );
  INV_X1 U14180 ( .A(n11170), .ZN(n11174) );
  AOI22_X1 U14181 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11172) );
  NAND2_X1 U14182 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11171) );
  NAND4_X1 U14183 ( .A1(n11174), .A2(n11173), .A3(n11172), .A4(n11171), .ZN(
        n11182) );
  AOI22_X1 U14184 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11180) );
  AOI22_X1 U14185 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11179) );
  AOI22_X1 U14186 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11178) );
  AOI22_X1 U14187 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11177) );
  NAND4_X1 U14188 ( .A1(n11180), .A2(n11179), .A3(n11178), .A4(n11177), .ZN(
        n11181) );
  XNOR2_X1 U14189 ( .A(n12116), .B(n12051), .ZN(n11183) );
  INV_X1 U14190 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15205) );
  INV_X1 U14191 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13628) );
  NAND2_X1 U14192 ( .A1(n11074), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11186) );
  NAND2_X1 U14193 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11185) );
  OAI211_X1 U14194 ( .C1(n11816), .C2(n13628), .A(n11186), .B(n11185), .ZN(
        n11187) );
  INV_X1 U14195 ( .A(n11187), .ZN(n11191) );
  AOI22_X1 U14196 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11189) );
  NAND2_X1 U14197 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11188) );
  NAND4_X1 U14198 ( .A1(n11191), .A2(n11190), .A3(n11189), .A4(n11188), .ZN(
        n11198) );
  AOI22_X1 U14199 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14200 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9592), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14201 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14202 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11193) );
  NAND4_X1 U14203 ( .A1(n11196), .A2(n11195), .A3(n11194), .A4(n11193), .ZN(
        n11197) );
  NAND3_X1 U14204 ( .A1(n14982), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n12052), 
        .ZN(n11199) );
  OAI211_X1 U14205 ( .C1(n11929), .C2(n15205), .A(n11200), .B(n11199), .ZN(
        n11201) );
  NAND2_X1 U14206 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11218) );
  OAI21_X1 U14207 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11218), .ZN(n13871) );
  OR2_X1 U14208 ( .A1(n16537), .A2(n13532), .ZN(n11213) );
  OAI21_X1 U14209 ( .B1(n12150), .B2(n13871), .A(n11213), .ZN(n11202) );
  INV_X1 U14210 ( .A(n11202), .ZN(n11203) );
  NAND3_X1 U14211 ( .A1(n13073), .A2(n13127), .A3(n9614), .ZN(n13137) );
  NAND2_X1 U14212 ( .A1(n11205), .A2(n14976), .ZN(n11206) );
  INV_X1 U14213 ( .A(n11209), .ZN(n11214) );
  XNOR2_X1 U14214 ( .A(n11210), .B(n11214), .ZN(n11207) );
  INV_X1 U14215 ( .A(n11208), .ZN(n11211) );
  NAND2_X1 U14216 ( .A1(n12044), .A2(n12052), .ZN(n11212) );
  INV_X1 U14217 ( .A(n11244), .ZN(n11243) );
  INV_X1 U14218 ( .A(n11213), .ZN(n11215) );
  OAI21_X1 U14219 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11215), .A(
        n11214), .ZN(n11216) );
  NAND2_X1 U14220 ( .A1(n9656), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11222) );
  INV_X1 U14221 ( .A(n12150), .ZN(n11220) );
  INV_X1 U14222 ( .A(n11218), .ZN(n16505) );
  NAND2_X1 U14223 ( .A1(n16505), .A2(n16513), .ZN(n13533) );
  NAND2_X1 U14224 ( .A1(n11218), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11219) );
  NAND2_X1 U14225 ( .A1(n13533), .A2(n11219), .ZN(n13606) );
  NAND2_X1 U14226 ( .A1(n11220), .A2(n13606), .ZN(n11221) );
  INV_X1 U14227 ( .A(n11227), .ZN(n13153) );
  INV_X1 U14228 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13636) );
  NAND2_X1 U14229 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11229) );
  NAND2_X1 U14230 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11228) );
  OAI211_X1 U14231 ( .C1(n13153), .C2(n13636), .A(n11229), .B(n11228), .ZN(
        n11230) );
  INV_X1 U14232 ( .A(n11230), .ZN(n11234) );
  AOI22_X1 U14233 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11232) );
  NAND2_X1 U14234 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11231) );
  NAND4_X1 U14235 ( .A1(n11234), .A2(n11233), .A3(n11232), .A4(n11231), .ZN(
        n11240) );
  INV_X1 U14236 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n21213) );
  AOI22_X1 U14237 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11238) );
  AOI22_X1 U14238 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11237) );
  AOI22_X1 U14239 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14240 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11235) );
  NAND4_X1 U14241 ( .A1(n11238), .A2(n11237), .A3(n11236), .A4(n11235), .ZN(
        n11239) );
  AOI22_X1 U14242 ( .A1(n11935), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11909), .B2(n12061), .ZN(n11241) );
  OAI21_X2 U14243 ( .B1(n13124), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11241), 
        .ZN(n11245) );
  NAND2_X1 U14244 ( .A1(n11255), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11290) );
  INV_X1 U14245 ( .A(n11204), .ZN(n13079) );
  NAND2_X1 U14246 ( .A1(n13079), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11318) );
  INV_X2 U14247 ( .A(n11319), .ZN(n13571) );
  XNOR2_X1 U14248 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14657) );
  AOI21_X1 U14249 ( .B1(n13571), .B2(n14657), .A(n12040), .ZN(n11247) );
  NOR2_X2 U14250 ( .A1(n13297), .A2(n11264), .ZN(n11257) );
  INV_X1 U14251 ( .A(n11803), .ZN(n11852) );
  NAND2_X1 U14252 ( .A1(n11852), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11246) );
  OAI211_X1 U14253 ( .C1(n11318), .C2(n13141), .A(n11247), .B(n11246), .ZN(
        n11248) );
  INV_X1 U14254 ( .A(n11248), .ZN(n11249) );
  OAI21_X2 U14255 ( .B1(n12060), .B2(n11290), .A(n11249), .ZN(n11250) );
  NAND2_X1 U14256 ( .A1(n12040), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11270) );
  INV_X1 U14257 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15200) );
  AOI21_X1 U14258 ( .B1(n14970), .B2(n12116), .A(n20963), .ZN(n11252) );
  NAND2_X1 U14259 ( .A1(n14982), .A2(n12051), .ZN(n11251) );
  OAI211_X1 U14260 ( .C1(n11929), .C2(n15200), .A(n11252), .B(n11251), .ZN(
        n11253) );
  NAND2_X1 U14261 ( .A1(n9606), .A2(n11255), .ZN(n11256) );
  NAND2_X1 U14262 ( .A1(n11256), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13033) );
  OR2_X1 U14263 ( .A1(n14445), .A2(n11290), .ZN(n11261) );
  INV_X1 U14264 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14265 ( .A1(n11257), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n11264), .ZN(n11259) );
  INV_X1 U14266 ( .A(n11318), .ZN(n11265) );
  NAND2_X1 U14267 ( .A1(n11265), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11258) );
  AND2_X1 U14268 ( .A1(n11259), .A2(n11258), .ZN(n11260) );
  OR2_X2 U14269 ( .A1(n13033), .A2(n13034), .ZN(n13035) );
  NAND2_X1 U14270 ( .A1(n13034), .A2(n13571), .ZN(n11262) );
  AOI22_X1 U14271 ( .A1(n11852), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11264), .ZN(n11267) );
  NAND2_X1 U14272 ( .A1(n11265), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11266) );
  AND2_X1 U14273 ( .A1(n11267), .A2(n11266), .ZN(n11268) );
  NAND2_X1 U14274 ( .A1(n9656), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11274) );
  NAND3_X1 U14275 ( .A1(n13870), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13421) );
  INV_X1 U14276 ( .A(n13421), .ZN(n15248) );
  NAND2_X1 U14277 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15248), .ZN(
        n13419) );
  NAND2_X1 U14278 ( .A1(n13870), .A2(n13419), .ZN(n11271) );
  NAND3_X1 U14279 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13869) );
  INV_X1 U14280 ( .A(n13869), .ZN(n13333) );
  NAND2_X1 U14281 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13333), .ZN(
        n13362) );
  NAND2_X1 U14282 ( .A1(n11271), .A2(n13362), .ZN(n13773) );
  OAI22_X1 U14283 ( .A1(n12150), .A2(n13773), .B1(n16537), .B2(n13870), .ZN(
        n11272) );
  INV_X1 U14284 ( .A(n11272), .ZN(n11273) );
  INV_X1 U14285 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13644) );
  NAND2_X1 U14286 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14287 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11275) );
  OAI211_X1 U14288 ( .C1(n11816), .C2(n13644), .A(n11276), .B(n11275), .ZN(
        n11277) );
  INV_X1 U14289 ( .A(n11277), .ZN(n11282) );
  AOI22_X1 U14290 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9613), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14291 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9616), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11280) );
  NAND2_X1 U14292 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11279) );
  NAND4_X1 U14293 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n11288) );
  AOI22_X1 U14294 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14295 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14296 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14297 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11283) );
  NAND4_X1 U14298 ( .A1(n11286), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(
        n11287) );
  AOI22_X1 U14299 ( .A1(n11935), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11909), .B2(n12080), .ZN(n11289) );
  NAND2_X1 U14300 ( .A1(n12069), .A2(n11524), .ZN(n11300) );
  INV_X1 U14301 ( .A(n11292), .ZN(n11291) );
  INV_X1 U14302 ( .A(n11321), .ZN(n11295) );
  INV_X1 U14303 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11293) );
  NAND2_X1 U14304 ( .A1(n11293), .A2(n11292), .ZN(n11294) );
  NAND2_X1 U14305 ( .A1(n11295), .A2(n11294), .ZN(n13962) );
  AOI22_X1 U14306 ( .A1(n13962), .A2(n13571), .B1(n12040), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11297) );
  NAND2_X1 U14307 ( .A1(n11852), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11296) );
  OAI211_X1 U14308 ( .C1(n11318), .C2(n13164), .A(n11297), .B(n11296), .ZN(
        n11298) );
  INV_X1 U14309 ( .A(n11298), .ZN(n11299) );
  NAND2_X1 U14310 ( .A1(n11300), .A2(n11299), .ZN(n13277) );
  NAND2_X1 U14311 ( .A1(n13278), .A2(n13277), .ZN(n13279) );
  INV_X1 U14312 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15219) );
  INV_X1 U14313 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13612) );
  NAND2_X1 U14314 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11303) );
  NAND2_X1 U14315 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11302) );
  OAI211_X1 U14316 ( .C1(n11816), .C2(n13612), .A(n11303), .B(n11302), .ZN(
        n11304) );
  INV_X1 U14317 ( .A(n11304), .ZN(n11308) );
  AOI22_X1 U14318 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U14319 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11305) );
  NAND4_X1 U14320 ( .A1(n11308), .A2(n11307), .A3(n11306), .A4(n11305), .ZN(
        n11314) );
  AOI22_X1 U14321 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14322 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14323 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14324 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11309) );
  NAND4_X1 U14325 ( .A1(n11312), .A2(n11311), .A3(n11310), .A4(n11309), .ZN(
        n11313) );
  NAND2_X1 U14326 ( .A1(n11909), .A2(n12090), .ZN(n11315) );
  XNOR2_X1 U14327 ( .A(n11326), .B(n11325), .ZN(n12079) );
  INV_X1 U14328 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n13658) );
  NAND2_X1 U14329 ( .A1(n13658), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11317) );
  NAND2_X1 U14330 ( .A1(n11852), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11316) );
  OAI211_X1 U14331 ( .C1(n11318), .C2(n11894), .A(n11317), .B(n11316), .ZN(
        n11320) );
  NAND2_X1 U14332 ( .A1(n11320), .A2(n11319), .ZN(n11323) );
  OAI21_X1 U14333 ( .B1(n11321), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11342), .ZN(n20795) );
  NAND2_X1 U14334 ( .A1(n20795), .A2(n13571), .ZN(n11322) );
  NAND2_X1 U14335 ( .A1(n11323), .A2(n11322), .ZN(n11324) );
  AOI21_X1 U14336 ( .B1(n12079), .B2(n11524), .A(n11324), .ZN(n13492) );
  NOR2_X2 U14337 ( .A1(n13279), .A2(n13492), .ZN(n13527) );
  NAND2_X1 U14338 ( .A1(n11935), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11341) );
  INV_X1 U14339 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13616) );
  NAND2_X1 U14340 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11328) );
  NAND2_X1 U14341 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11327) );
  OAI211_X1 U14342 ( .C1(n13153), .C2(n13616), .A(n11328), .B(n11327), .ZN(
        n11329) );
  INV_X1 U14343 ( .A(n11329), .ZN(n11333) );
  AOI22_X1 U14344 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9613), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14345 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U14346 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11330) );
  NAND4_X1 U14347 ( .A1(n11333), .A2(n11332), .A3(n11331), .A4(n11330), .ZN(
        n11339) );
  AOI22_X1 U14348 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9616), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14349 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14350 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14351 ( .A1(n11837), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11334) );
  NAND4_X1 U14352 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(
        n11338) );
  NAND2_X1 U14353 ( .A1(n11909), .A2(n12099), .ZN(n11340) );
  NAND2_X1 U14354 ( .A1(n11341), .A2(n11340), .ZN(n11376) );
  XNOR2_X1 U14355 ( .A(n11373), .B(n11376), .ZN(n12088) );
  NAND2_X1 U14356 ( .A1(n12088), .A2(n11524), .ZN(n11348) );
  INV_X1 U14357 ( .A(n12040), .ZN(n11436) );
  AND2_X1 U14358 ( .A1(n11342), .A2(n11345), .ZN(n11343) );
  OR2_X1 U14359 ( .A1(n11343), .A2(n11367), .ZN(n20685) );
  NAND2_X1 U14360 ( .A1(n20685), .A2(n13571), .ZN(n11344) );
  OAI21_X1 U14361 ( .B1(n11345), .B2(n11436), .A(n11344), .ZN(n11346) );
  AOI21_X1 U14362 ( .B1(n11852), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11346), .ZN(
        n11347) );
  NAND2_X1 U14363 ( .A1(n11348), .A2(n11347), .ZN(n13526) );
  NAND2_X1 U14364 ( .A1(n13527), .A2(n13526), .ZN(n13525) );
  INV_X1 U14365 ( .A(n11376), .ZN(n11349) );
  NAND2_X1 U14366 ( .A1(n11935), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11365) );
  INV_X1 U14367 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13620) );
  NAND2_X1 U14368 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11351) );
  NAND2_X1 U14369 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11350) );
  OAI211_X1 U14370 ( .C1(n13153), .C2(n13620), .A(n11351), .B(n11350), .ZN(
        n11352) );
  INV_X1 U14371 ( .A(n11352), .ZN(n11357) );
  AOI22_X1 U14372 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U14373 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11354) );
  NAND4_X1 U14374 ( .A1(n11357), .A2(n11356), .A3(n11355), .A4(n11354), .ZN(
        n11363) );
  AOI22_X1 U14375 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14376 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14377 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14378 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11358) );
  NAND4_X1 U14379 ( .A1(n11361), .A2(n11360), .A3(n11359), .A4(n11358), .ZN(
        n11362) );
  NAND2_X1 U14380 ( .A1(n11909), .A2(n12107), .ZN(n11364) );
  INV_X1 U14381 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11370) );
  OR2_X1 U14382 ( .A1(n11367), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11368) );
  NAND2_X1 U14383 ( .A1(n11381), .A2(n11368), .ZN(n20674) );
  AOI22_X1 U14384 ( .A1(n20674), .A2(n13571), .B1(n12040), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11369) );
  OAI21_X1 U14385 ( .B1(n11803), .B2(n11370), .A(n11369), .ZN(n11371) );
  INV_X1 U14386 ( .A(n11374), .ZN(n11375) );
  INV_X1 U14387 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15235) );
  INV_X1 U14388 ( .A(n12116), .ZN(n11379) );
  OAI22_X1 U14389 ( .A1(n11929), .A2(n15235), .B1(n11915), .B2(n11379), .ZN(
        n11380) );
  INV_X1 U14390 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11386) );
  NAND2_X1 U14391 ( .A1(n11381), .A2(n11383), .ZN(n11382) );
  NAND2_X1 U14392 ( .A1(n11405), .A2(n11382), .ZN(n20661) );
  NOR2_X1 U14393 ( .A1(n11436), .A2(n11383), .ZN(n11384) );
  AOI21_X1 U14394 ( .B1(n20661), .B2(n13571), .A(n11384), .ZN(n11385) );
  OAI21_X1 U14395 ( .B1(n11803), .B2(n11386), .A(n11385), .ZN(n11387) );
  NAND2_X1 U14396 ( .A1(n11852), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14397 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14398 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9592), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14399 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14400 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11389) );
  AND4_X1 U14401 ( .A1(n11392), .A2(n11391), .A3(n11390), .A4(n11389), .ZN(
        n11399) );
  AOI22_X1 U14402 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14403 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14404 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9613), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11394) );
  NAND2_X1 U14405 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11393) );
  AND3_X1 U14406 ( .A1(n11395), .A2(n11394), .A3(n11393), .ZN(n11397) );
  NAND2_X1 U14407 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11396) );
  NAND4_X1 U14408 ( .A1(n11399), .A2(n11398), .A3(n11397), .A4(n11396), .ZN(
        n11400) );
  NAND2_X1 U14409 ( .A1(n11524), .A2(n11400), .ZN(n11403) );
  XNOR2_X1 U14410 ( .A(n11405), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14139) );
  OR2_X1 U14411 ( .A1(n14139), .A2(n11319), .ZN(n11402) );
  NAND2_X1 U14412 ( .A1(n12040), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11401) );
  XOR2_X1 U14413 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11420), .Z(n13984) );
  AOI22_X1 U14414 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9617), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14415 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14416 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14417 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11406) );
  AND4_X1 U14418 ( .A1(n11409), .A2(n11408), .A3(n11407), .A4(n11406), .ZN(
        n11416) );
  AOI22_X1 U14419 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9592), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14420 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11412) );
  NAND2_X1 U14421 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11410) );
  AND3_X1 U14422 ( .A1(n11412), .A2(n11411), .A3(n11410), .ZN(n11414) );
  NAND2_X1 U14423 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11413) );
  NAND4_X1 U14424 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n11417) );
  AOI22_X1 U14425 ( .A1(n11524), .A2(n11417), .B1(n12040), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11419) );
  NAND2_X1 U14426 ( .A1(n11852), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11418) );
  OAI211_X1 U14427 ( .C1(n13984), .C2(n11319), .A(n11419), .B(n11418), .ZN(
        n13973) );
  XNOR2_X1 U14428 ( .A(n11440), .B(n14946), .ZN(n14066) );
  NAND2_X1 U14429 ( .A1(n14066), .A2(n13571), .ZN(n11439) );
  NAND2_X1 U14430 ( .A1(n11852), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14431 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14432 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14433 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14434 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11421) );
  AND4_X1 U14435 ( .A1(n11424), .A2(n11423), .A3(n11422), .A4(n11421), .ZN(
        n11432) );
  AOI22_X1 U14436 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9617), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11431) );
  NAND2_X1 U14437 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11428) );
  AOI22_X1 U14438 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9613), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11427) );
  NAND2_X1 U14439 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11426) );
  NAND2_X1 U14440 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11425) );
  AND4_X1 U14441 ( .A1(n11428), .A2(n11427), .A3(n11426), .A4(n11425), .ZN(
        n11430) );
  NAND2_X1 U14442 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11429) );
  NAND4_X1 U14443 ( .A1(n11432), .A2(n11431), .A3(n11430), .A4(n11429), .ZN(
        n11433) );
  NAND2_X1 U14444 ( .A1(n11524), .A2(n11433), .ZN(n11434) );
  OAI211_X1 U14445 ( .C1(n11436), .C2(n14946), .A(n11435), .B(n11434), .ZN(
        n11437) );
  INV_X1 U14446 ( .A(n11437), .ZN(n11438) );
  NAND2_X1 U14447 ( .A1(n11439), .A2(n11438), .ZN(n14031) );
  NAND2_X1 U14448 ( .A1(n11257), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11443) );
  OAI21_X1 U14449 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11441), .A(
        n11474), .ZN(n16682) );
  AOI22_X1 U14450 ( .A1(n13571), .A2(n16682), .B1(n12040), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11442) );
  NAND2_X1 U14451 ( .A1(n11443), .A2(n11442), .ZN(n11456) );
  AOI22_X1 U14452 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14453 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U14454 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9616), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14455 ( .A1(n11837), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11444) );
  AND4_X1 U14456 ( .A1(n11447), .A2(n11446), .A3(n11445), .A4(n11444), .ZN(
        n11454) );
  AOI22_X1 U14457 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14458 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U14459 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11449) );
  AND3_X1 U14460 ( .A1(n11450), .A2(n11449), .A3(n11448), .ZN(n11452) );
  NAND2_X1 U14461 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11451) );
  NAND4_X1 U14462 ( .A1(n11454), .A2(n11453), .A3(n11452), .A4(n11451), .ZN(
        n11455) );
  AND2_X1 U14463 ( .A1(n11524), .A2(n11455), .ZN(n14143) );
  INV_X1 U14464 ( .A(n11456), .ZN(n11457) );
  NAND2_X2 U14465 ( .A1(n14146), .A2(n11458), .ZN(n14727) );
  XOR2_X1 U14466 ( .A(n11473), .B(n11474), .Z(n16670) );
  AOI22_X1 U14467 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14468 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9592), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14469 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14470 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11459) );
  AND4_X1 U14471 ( .A1(n11462), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(
        n11469) );
  AOI22_X1 U14472 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14473 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14474 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9613), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11464) );
  NAND2_X1 U14475 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11463) );
  AND3_X1 U14476 ( .A1(n11465), .A2(n11464), .A3(n11463), .ZN(n11467) );
  NAND2_X1 U14477 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11466) );
  NAND4_X1 U14478 ( .A1(n11469), .A2(n11468), .A3(n11467), .A4(n11466), .ZN(
        n11470) );
  AOI22_X1 U14479 ( .A1(n11524), .A2(n11470), .B1(n12040), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11472) );
  NAND2_X1 U14480 ( .A1(n11257), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11471) );
  OAI211_X1 U14481 ( .C1(n16670), .C2(n11319), .A(n11472), .B(n11471), .ZN(
        n14726) );
  XNOR2_X1 U14482 ( .A(n11494), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16613) );
  AOI22_X1 U14483 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14484 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14485 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14486 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11475) );
  NAND4_X1 U14487 ( .A1(n11478), .A2(n11477), .A3(n11476), .A4(n11475), .ZN(
        n11488) );
  INV_X1 U14488 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U14489 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11480) );
  NAND2_X1 U14490 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11479) );
  OAI211_X1 U14491 ( .C1(n11816), .C2(n11481), .A(n11480), .B(n11479), .ZN(
        n11482) );
  INV_X1 U14492 ( .A(n11482), .ZN(n11486) );
  AOI22_X1 U14493 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11484) );
  NAND2_X1 U14494 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11483) );
  NAND4_X1 U14495 ( .A1(n11486), .A2(n11485), .A3(n11484), .A4(n11483), .ZN(
        n11487) );
  OAI21_X1 U14496 ( .B1(n11488), .B2(n11487), .A(n11524), .ZN(n11491) );
  NAND2_X1 U14497 ( .A1(n11257), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11490) );
  NAND2_X1 U14498 ( .A1(n12040), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11489) );
  NAND3_X1 U14499 ( .A1(n11491), .A2(n11490), .A3(n11489), .ZN(n11492) );
  AOI21_X1 U14500 ( .B1(n16613), .B2(n13571), .A(n11492), .ZN(n14720) );
  XOR2_X1 U14501 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11511), .Z(
        n16664) );
  AOI22_X1 U14502 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14503 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U14504 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11496) );
  AOI22_X1 U14505 ( .A1(n11837), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11495) );
  AND4_X1 U14506 ( .A1(n11498), .A2(n11497), .A3(n11496), .A4(n11495), .ZN(
        n11506) );
  AOI22_X1 U14507 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11505) );
  NAND2_X1 U14508 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11502) );
  NAND2_X1 U14509 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U14510 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11499) );
  AND4_X1 U14511 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(
        n11504) );
  NAND2_X1 U14512 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11503) );
  NAND4_X1 U14513 ( .A1(n11506), .A2(n11505), .A3(n11504), .A4(n11503), .ZN(
        n11507) );
  AOI22_X1 U14514 ( .A1(n11524), .A2(n11507), .B1(n12040), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11509) );
  NAND2_X1 U14515 ( .A1(n11257), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11508) );
  OAI211_X1 U14516 ( .C1(n16664), .C2(n11319), .A(n11509), .B(n11508), .ZN(
        n11510) );
  XNOR2_X1 U14517 ( .A(n11551), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16598) );
  INV_X1 U14518 ( .A(n16598), .ZN(n21062) );
  AOI22_X1 U14519 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n11176), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14520 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14521 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9616), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14522 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11512) );
  NAND4_X1 U14523 ( .A1(n11515), .A2(n11514), .A3(n11513), .A4(n11512), .ZN(
        n11526) );
  INV_X1 U14524 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11518) );
  NAND2_X1 U14525 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11517) );
  NAND2_X1 U14526 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11516) );
  OAI211_X1 U14527 ( .C1(n13153), .C2(n11518), .A(n11517), .B(n11516), .ZN(
        n11519) );
  INV_X1 U14528 ( .A(n11519), .ZN(n11523) );
  AOI22_X1 U14529 ( .A1(n11837), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11521) );
  NAND2_X1 U14530 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11520) );
  NAND4_X1 U14531 ( .A1(n11523), .A2(n11522), .A3(n11521), .A4(n11520), .ZN(
        n11525) );
  OAI21_X1 U14532 ( .B1(n11526), .B2(n11525), .A(n11524), .ZN(n11529) );
  NAND2_X1 U14533 ( .A1(n11852), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11528) );
  NAND2_X1 U14534 ( .A1(n12040), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11527) );
  NAND3_X1 U14535 ( .A1(n11529), .A2(n11528), .A3(n11527), .ZN(n11530) );
  AOI21_X1 U14536 ( .B1(n21062), .B2(n13571), .A(n11530), .ZN(n14709) );
  AOI22_X1 U14537 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14538 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9592), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14539 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14540 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11533) );
  NAND4_X1 U14541 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11546) );
  NAND2_X1 U14542 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11540) );
  NAND2_X1 U14543 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11539) );
  NAND2_X1 U14544 ( .A1(n11842), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11538) );
  NAND2_X1 U14545 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11537) );
  AND4_X1 U14546 ( .A1(n11540), .A2(n11539), .A3(n11538), .A4(n11537), .ZN(
        n11544) );
  AOI22_X1 U14547 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11543) );
  NAND2_X1 U14548 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11542) );
  NAND2_X1 U14549 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11541) );
  NAND4_X1 U14550 ( .A1(n11544), .A2(n11543), .A3(n11542), .A4(n11541), .ZN(
        n11545) );
  NOR2_X1 U14551 ( .A1(n11546), .A2(n11545), .ZN(n11550) );
  NAND2_X1 U14552 ( .A1(n13658), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14553 ( .A1(n11319), .A2(n11547), .ZN(n11548) );
  AOI21_X1 U14554 ( .B1(n11257), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11548), .ZN(
        n11549) );
  OAI21_X1 U14555 ( .B1(n11883), .B2(n11550), .A(n11549), .ZN(n11554) );
  OAI21_X1 U14556 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11552), .A(
        n11588), .ZN(n16583) );
  OR2_X1 U14557 ( .A1(n11319), .A2(n16583), .ZN(n11553) );
  AOI22_X1 U14558 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9617), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14559 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14560 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14561 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11555) );
  AND4_X1 U14562 ( .A1(n11558), .A2(n11557), .A3(n11556), .A4(n11555), .ZN(
        n11565) );
  AOI22_X1 U14563 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14564 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14565 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9613), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11560) );
  NAND2_X1 U14566 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11559) );
  AND3_X1 U14567 ( .A1(n11561), .A2(n11560), .A3(n11559), .ZN(n11563) );
  NAND2_X1 U14568 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11562) );
  NAND4_X1 U14569 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11569) );
  INV_X1 U14570 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14787) );
  INV_X1 U14571 ( .A(n11588), .ZN(n11566) );
  XNOR2_X1 U14572 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11566), .ZN(
        n14930) );
  AOI22_X1 U14573 ( .A1(n13571), .A2(n14930), .B1(n12040), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11567) );
  OAI21_X1 U14574 ( .B1(n11803), .B2(n14787), .A(n11567), .ZN(n11568) );
  AOI21_X1 U14575 ( .B1(n11849), .B2(n11569), .A(n11568), .ZN(n14644) );
  INV_X1 U14576 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U14577 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11571) );
  NAND2_X1 U14578 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11570) );
  OAI211_X1 U14579 ( .C1(n13153), .C2(n11572), .A(n11571), .B(n11570), .ZN(
        n11573) );
  INV_X1 U14580 ( .A(n11573), .ZN(n11577) );
  AOI22_X1 U14581 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11575) );
  NAND2_X1 U14582 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11574) );
  NAND4_X1 U14583 ( .A1(n11577), .A2(n11576), .A3(n11575), .A4(n11574), .ZN(
        n11583) );
  AOI22_X1 U14584 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9617), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14585 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14586 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14587 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11578) );
  NAND4_X1 U14588 ( .A1(n11581), .A2(n11580), .A3(n11579), .A4(n11578), .ZN(
        n11582) );
  NOR2_X1 U14589 ( .A1(n11583), .A2(n11582), .ZN(n11587) );
  NAND2_X1 U14590 ( .A1(n13658), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11584) );
  NAND2_X1 U14591 ( .A1(n11319), .A2(n11584), .ZN(n11585) );
  AOI21_X1 U14592 ( .B1(n11257), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11585), .ZN(
        n11586) );
  OAI21_X1 U14593 ( .B1(n11883), .B2(n11587), .A(n11586), .ZN(n11591) );
  OAI21_X1 U14594 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11589), .A(
        n11630), .ZN(n16574) );
  OR2_X1 U14595 ( .A1(n11319), .A2(n16574), .ZN(n11590) );
  NAND2_X1 U14596 ( .A1(n11591), .A2(n11590), .ZN(n14689) );
  AOI22_X1 U14597 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9602), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11599) );
  NAND2_X1 U14598 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11595) );
  NAND2_X1 U14599 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11594) );
  NAND2_X1 U14600 ( .A1(n11842), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11593) );
  NAND2_X1 U14601 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11592) );
  AND4_X1 U14602 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11598) );
  NAND2_X1 U14603 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11597) );
  NAND2_X1 U14604 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11596) );
  NAND4_X1 U14605 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(
        n11605) );
  AOI22_X1 U14606 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14607 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14608 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14609 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11600) );
  NAND4_X1 U14610 ( .A1(n11603), .A2(n11602), .A3(n11601), .A4(n11600), .ZN(
        n11604) );
  NOR2_X1 U14611 ( .A1(n11605), .A2(n11604), .ZN(n11609) );
  NAND2_X1 U14612 ( .A1(n13658), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11606) );
  NAND2_X1 U14613 ( .A1(n11319), .A2(n11606), .ZN(n11607) );
  AOI21_X1 U14614 ( .B1(n11257), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11607), .ZN(
        n11608) );
  OAI21_X1 U14615 ( .B1(n11883), .B2(n11609), .A(n11608), .ZN(n11611) );
  XNOR2_X1 U14616 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n11630), .ZN(
        n14907) );
  NAND2_X1 U14617 ( .A1(n13571), .A2(n14907), .ZN(n11610) );
  NAND2_X1 U14618 ( .A1(n11611), .A2(n11610), .ZN(n14631) );
  NOR2_X2 U14619 ( .A1(n14628), .A2(n14631), .ZN(n14629) );
  AOI22_X1 U14620 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14621 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14622 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9592), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14623 ( .A1(n11837), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11612) );
  NAND4_X1 U14624 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n11625) );
  NAND2_X1 U14625 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11619) );
  NAND2_X1 U14626 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11618) );
  NAND2_X1 U14627 ( .A1(n11842), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11617) );
  AND4_X1 U14628 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n11623) );
  AOI22_X1 U14629 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11622) );
  NAND2_X1 U14630 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11621) );
  NAND2_X1 U14631 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11620) );
  NAND4_X1 U14632 ( .A1(n11623), .A2(n11622), .A3(n11621), .A4(n11620), .ZN(
        n11624) );
  NOR2_X1 U14633 ( .A1(n11625), .A2(n11624), .ZN(n11629) );
  NAND2_X1 U14634 ( .A1(n13658), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11626) );
  NAND2_X1 U14635 ( .A1(n11319), .A2(n11626), .ZN(n11627) );
  AOI21_X1 U14636 ( .B1(n11257), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11627), .ZN(
        n11628) );
  OAI21_X1 U14637 ( .B1(n11883), .B2(n11629), .A(n11628), .ZN(n11637) );
  INV_X1 U14638 ( .A(n11632), .ZN(n11634) );
  INV_X1 U14639 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11633) );
  NAND2_X1 U14640 ( .A1(n11634), .A2(n11633), .ZN(n11635) );
  NAND2_X1 U14641 ( .A1(n11676), .A2(n11635), .ZN(n16573) );
  OR2_X1 U14642 ( .A1(n16573), .A2(n11319), .ZN(n11636) );
  INV_X1 U14643 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11640) );
  NAND2_X1 U14644 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11639) );
  NAND2_X1 U14645 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11638) );
  OAI211_X1 U14646 ( .C1(n13153), .C2(n11640), .A(n11639), .B(n11638), .ZN(
        n11641) );
  INV_X1 U14647 ( .A(n11641), .ZN(n11645) );
  AOI22_X1 U14648 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n9613), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14649 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11643) );
  NAND2_X1 U14650 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11642) );
  NAND4_X1 U14651 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11651) );
  AOI22_X1 U14652 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14653 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14654 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14655 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11646) );
  NAND4_X1 U14656 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n11650) );
  NOR2_X1 U14657 ( .A1(n11651), .A2(n11650), .ZN(n11655) );
  NAND2_X1 U14658 ( .A1(n13658), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11652) );
  NAND2_X1 U14659 ( .A1(n11319), .A2(n11652), .ZN(n11653) );
  AOI21_X1 U14660 ( .B1(n11257), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11653), .ZN(
        n11654) );
  OAI21_X1 U14661 ( .B1(n11883), .B2(n11655), .A(n11654), .ZN(n11657) );
  XNOR2_X1 U14662 ( .A(n11676), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14619) );
  NAND2_X1 U14663 ( .A1(n14619), .A2(n13571), .ZN(n11656) );
  NAND2_X1 U14664 ( .A1(n11657), .A2(n11656), .ZN(n14616) );
  INV_X1 U14665 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14666 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11659) );
  NAND2_X1 U14667 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11658) );
  OAI211_X1 U14668 ( .C1(n13153), .C2(n11660), .A(n11659), .B(n11658), .ZN(
        n11661) );
  INV_X1 U14669 ( .A(n11661), .ZN(n11665) );
  AOI22_X1 U14670 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n9613), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14671 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11663) );
  NAND2_X1 U14672 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11662) );
  NAND4_X1 U14673 ( .A1(n11665), .A2(n11664), .A3(n11663), .A4(n11662), .ZN(
        n11671) );
  AOI22_X1 U14674 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9617), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14675 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14676 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14677 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11666) );
  NAND4_X1 U14678 ( .A1(n11669), .A2(n11668), .A3(n11667), .A4(n11666), .ZN(
        n11670) );
  NOR2_X1 U14679 ( .A1(n11671), .A2(n11670), .ZN(n11675) );
  INV_X1 U14680 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20640) );
  OAI21_X1 U14681 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20640), .A(
        n13658), .ZN(n11672) );
  INV_X1 U14682 ( .A(n11672), .ZN(n11673) );
  AOI21_X1 U14683 ( .B1(n11852), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11673), .ZN(
        n11674) );
  OAI21_X1 U14684 ( .B1(n11883), .B2(n11675), .A(n11674), .ZN(n11682) );
  INV_X1 U14685 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14620) );
  INV_X1 U14686 ( .A(n11677), .ZN(n11679) );
  INV_X1 U14687 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11678) );
  NAND2_X1 U14688 ( .A1(n11679), .A2(n11678), .ZN(n11680) );
  NAND2_X1 U14689 ( .A1(n11713), .A2(n11680), .ZN(n14886) );
  INV_X1 U14690 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11691) );
  INV_X1 U14691 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11684) );
  OAI22_X1 U14692 ( .A1(n9601), .A2(n13632), .B1(n11859), .B2(n11684), .ZN(
        n11688) );
  INV_X1 U14693 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11686) );
  INV_X1 U14694 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11685) );
  OAI22_X1 U14695 ( .A1(n9593), .A2(n11686), .B1(n11861), .B2(n11685), .ZN(
        n11687) );
  AOI211_X1 U14696 ( .C1(n11864), .C2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n11688), .B(n11687), .ZN(n11690) );
  AOI22_X1 U14697 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11689) );
  OAI211_X1 U14698 ( .C1(n13153), .C2(n11691), .A(n11690), .B(n11689), .ZN(
        n11697) );
  AOI22_X1 U14699 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14700 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9592), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14701 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9613), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14702 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11692) );
  NAND4_X1 U14703 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n11696) );
  NOR2_X1 U14704 ( .A1(n11697), .A2(n11696), .ZN(n11718) );
  INV_X1 U14705 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11858) );
  INV_X1 U14706 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U14707 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14708 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9613), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11698) );
  OAI211_X1 U14709 ( .C1(n11857), .C2(n13153), .A(n11699), .B(n11698), .ZN(
        n11700) );
  INV_X1 U14710 ( .A(n11700), .ZN(n11702) );
  AOI22_X1 U14711 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11701) );
  OAI211_X1 U14712 ( .C1(n11858), .C2(n11154), .A(n11702), .B(n11701), .ZN(
        n11708) );
  AOI22_X1 U14713 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14714 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14715 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9616), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14716 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11703) );
  NAND4_X1 U14717 ( .A1(n11706), .A2(n11705), .A3(n11704), .A4(n11703), .ZN(
        n11707) );
  NOR2_X1 U14718 ( .A1(n11708), .A2(n11707), .ZN(n11719) );
  XOR2_X1 U14719 ( .A(n11718), .B(n11719), .Z(n11709) );
  NAND2_X1 U14720 ( .A1(n11709), .A2(n11849), .ZN(n11712) );
  INV_X1 U14721 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14591) );
  NOR2_X1 U14722 ( .A1(n14591), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11710) );
  AOI211_X1 U14723 ( .C1(n11852), .C2(P1_EAX_REG_23__SCAN_IN), .A(n13571), .B(
        n11710), .ZN(n11711) );
  XNOR2_X1 U14724 ( .A(n11713), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14590) );
  AOI22_X1 U14725 ( .A1(n11712), .A2(n11711), .B1(n13571), .B2(n14590), .ZN(
        n14589) );
  INV_X1 U14726 ( .A(n11715), .ZN(n11716) );
  INV_X1 U14727 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14582) );
  NAND2_X1 U14728 ( .A1(n11716), .A2(n14582), .ZN(n11717) );
  NAND2_X1 U14729 ( .A1(n11759), .A2(n11717), .ZN(n14870) );
  NOR2_X1 U14730 ( .A1(n11719), .A2(n11718), .ZN(n11739) );
  INV_X1 U14731 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11722) );
  NAND2_X1 U14732 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U14733 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11720) );
  OAI211_X1 U14734 ( .C1(n13153), .C2(n11722), .A(n11721), .B(n11720), .ZN(
        n11723) );
  INV_X1 U14735 ( .A(n11723), .ZN(n11727) );
  AOI22_X1 U14736 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11725) );
  NAND2_X1 U14737 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11724) );
  NAND4_X1 U14738 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n11733) );
  AOI22_X1 U14739 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14740 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14741 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U14742 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11728) );
  NAND4_X1 U14743 ( .A1(n11731), .A2(n11730), .A3(n11729), .A4(n11728), .ZN(
        n11732) );
  OR2_X1 U14744 ( .A1(n11733), .A2(n11732), .ZN(n11738) );
  XNOR2_X1 U14745 ( .A(n11739), .B(n11738), .ZN(n11736) );
  AOI21_X1 U14746 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n13658), .A(
        n13571), .ZN(n11735) );
  NAND2_X1 U14747 ( .A1(n11257), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n11734) );
  OAI211_X1 U14748 ( .C1(n11736), .C2(n11883), .A(n11735), .B(n11734), .ZN(
        n11737) );
  XNOR2_X1 U14749 ( .A(n11759), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14567) );
  NAND2_X1 U14750 ( .A1(n11739), .A2(n11738), .ZN(n11764) );
  INV_X1 U14751 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11747) );
  INV_X1 U14752 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13685) );
  INV_X1 U14753 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11740) );
  OAI22_X1 U14754 ( .A1(n11741), .A2(n13685), .B1(n11859), .B2(n11740), .ZN(
        n11744) );
  INV_X1 U14755 ( .A(n11870), .ZN(n11742) );
  INV_X1 U14756 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15210) );
  OAI22_X1 U14757 ( .A1(n9601), .A2(n13636), .B1(n11742), .B2(n15210), .ZN(
        n11743) );
  AOI211_X1 U14758 ( .C1(n11227), .C2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n11744), .B(n11743), .ZN(n11746) );
  AOI22_X1 U14759 ( .A1(n9602), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11745) );
  OAI211_X1 U14760 ( .C1(n11154), .C2(n11747), .A(n11746), .B(n11745), .ZN(
        n11753) );
  AOI22_X1 U14761 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14762 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14763 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14764 ( .A1(n11842), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9613), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11748) );
  NAND4_X1 U14765 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11752) );
  NOR2_X1 U14766 ( .A1(n11753), .A2(n11752), .ZN(n11765) );
  XOR2_X1 U14767 ( .A(n11764), .B(n11765), .Z(n11757) );
  INV_X1 U14768 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n11755) );
  NOR2_X1 U14769 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11754) );
  OAI22_X1 U14770 ( .A1(n11803), .A2(n11755), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11754), .ZN(n11756) );
  AOI21_X1 U14771 ( .B1(n11757), .B2(n11849), .A(n11756), .ZN(n11758) );
  AOI21_X1 U14772 ( .B1(n13571), .B2(n14567), .A(n11758), .ZN(n14566) );
  NAND2_X1 U14773 ( .A1(n14565), .A2(n14566), .ZN(n14547) );
  INV_X1 U14774 ( .A(n11759), .ZN(n11760) );
  INV_X1 U14775 ( .A(n11761), .ZN(n11762) );
  INV_X1 U14776 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14550) );
  NAND2_X1 U14777 ( .A1(n11762), .A2(n14550), .ZN(n11763) );
  NAND2_X1 U14778 ( .A1(n11808), .A2(n11763), .ZN(n14853) );
  NOR2_X1 U14779 ( .A1(n11765), .A2(n11764), .ZN(n11785) );
  INV_X1 U14780 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11768) );
  NAND2_X1 U14781 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11767) );
  NAND2_X1 U14782 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11766) );
  OAI211_X1 U14783 ( .C1(n13153), .C2(n11768), .A(n11767), .B(n11766), .ZN(
        n11769) );
  INV_X1 U14784 ( .A(n11769), .ZN(n11773) );
  AOI22_X1 U14785 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11771) );
  NAND2_X1 U14786 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11770) );
  NAND4_X1 U14787 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n11779) );
  AOI22_X1 U14788 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14789 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14790 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14791 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11774) );
  NAND4_X1 U14792 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11778) );
  OR2_X1 U14793 ( .A1(n11779), .A2(n11778), .ZN(n11784) );
  XNOR2_X1 U14794 ( .A(n11785), .B(n11784), .ZN(n11782) );
  AOI21_X1 U14795 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n13658), .A(
        n13571), .ZN(n11781) );
  NAND2_X1 U14796 ( .A1(n11257), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n11780) );
  OAI211_X1 U14797 ( .C1(n11782), .C2(n11883), .A(n11781), .B(n11780), .ZN(
        n11783) );
  OAI21_X1 U14798 ( .B1(n11319), .B2(n14853), .A(n11783), .ZN(n14549) );
  XNOR2_X1 U14799 ( .A(n11808), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14841) );
  NAND2_X1 U14800 ( .A1(n11785), .A2(n11784), .ZN(n11811) );
  INV_X1 U14801 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11794) );
  INV_X1 U14802 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11788) );
  INV_X1 U14803 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11786) );
  OAI22_X1 U14804 ( .A1(n11859), .A2(n11788), .B1(n9596), .B2(n11786), .ZN(
        n11791) );
  INV_X1 U14805 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11789) );
  OAI22_X1 U14806 ( .A1(n9601), .A2(n13612), .B1(n11861), .B2(n11789), .ZN(
        n11790) );
  AOI211_X1 U14807 ( .C1(n11864), .C2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n11791), .B(n11790), .ZN(n11793) );
  AOI22_X1 U14808 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11792) );
  OAI211_X1 U14809 ( .C1(n13153), .C2(n11794), .A(n11793), .B(n11792), .ZN(
        n11800) );
  AOI22_X1 U14810 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14811 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9592), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14812 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14813 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11795) );
  NAND4_X1 U14814 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11799) );
  NOR2_X1 U14815 ( .A1(n11800), .A2(n11799), .ZN(n11812) );
  XOR2_X1 U14816 ( .A(n11811), .B(n11812), .Z(n11805) );
  INV_X1 U14817 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n11802) );
  NOR2_X1 U14818 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11801) );
  OAI22_X1 U14819 ( .A1(n11803), .A2(n11802), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11801), .ZN(n11804) );
  AOI21_X1 U14820 ( .B1(n11805), .B2(n11849), .A(n11804), .ZN(n11806) );
  AOI21_X1 U14821 ( .B1(n13571), .B2(n14841), .A(n11806), .ZN(n14536) );
  INV_X1 U14822 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11807) );
  INV_X1 U14823 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14527) );
  NAND2_X1 U14824 ( .A1(n11809), .A2(n14527), .ZN(n11810) );
  NAND2_X1 U14825 ( .A1(n11855), .A2(n11810), .ZN(n14832) );
  NOR2_X1 U14826 ( .A1(n11812), .A2(n11811), .ZN(n11833) );
  INV_X1 U14827 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11815) );
  NAND2_X1 U14828 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11814) );
  NAND2_X1 U14829 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11813) );
  OAI211_X1 U14830 ( .C1(n11816), .C2(n11815), .A(n11814), .B(n11813), .ZN(
        n11817) );
  INV_X1 U14831 ( .A(n11817), .ZN(n11821) );
  AOI22_X1 U14832 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U14833 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11818) );
  NAND4_X1 U14834 ( .A1(n11821), .A2(n11820), .A3(n11819), .A4(n11818), .ZN(
        n11827) );
  AOI22_X1 U14835 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9602), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14836 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14837 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U14838 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11822) );
  NAND4_X1 U14839 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n11826) );
  OR2_X1 U14840 ( .A1(n11827), .A2(n11826), .ZN(n11832) );
  XNOR2_X1 U14841 ( .A(n11833), .B(n11832), .ZN(n11830) );
  AOI21_X1 U14842 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n13658), .A(
        n13571), .ZN(n11829) );
  NAND2_X1 U14843 ( .A1(n11257), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n11828) );
  OAI211_X1 U14844 ( .C1(n11830), .C2(n11883), .A(n11829), .B(n11828), .ZN(
        n11831) );
  OAI21_X1 U14845 ( .B1(n11319), .B2(n14832), .A(n11831), .ZN(n14524) );
  NAND2_X1 U14846 ( .A1(n11833), .A2(n11832), .ZN(n11877) );
  INV_X1 U14847 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13402) );
  INV_X1 U14848 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11834) );
  OAI22_X1 U14849 ( .A1(n11159), .A2(n13402), .B1(n9593), .B2(n11834), .ZN(
        n11836) );
  AOI21_X1 U14850 ( .B1(n11864), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n11836), .ZN(n11841) );
  AOI22_X1 U14851 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11839) );
  NAND2_X1 U14852 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11838) );
  NAND4_X1 U14853 ( .A1(n11841), .A2(n11840), .A3(n11839), .A4(n11838), .ZN(
        n11848) );
  AOI22_X1 U14854 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n9602), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14855 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11842), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U14856 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14857 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9597), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11843) );
  NAND4_X1 U14858 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n11847) );
  NOR2_X1 U14859 ( .A1(n11848), .A2(n11847), .ZN(n11878) );
  XOR2_X1 U14860 ( .A(n11877), .B(n11878), .Z(n11850) );
  NAND2_X1 U14861 ( .A1(n11850), .A2(n11849), .ZN(n11854) );
  INV_X1 U14862 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14392) );
  NOR2_X1 U14863 ( .A1(n14392), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11851) );
  AOI211_X1 U14864 ( .C1(n11852), .C2(P1_EAX_REG_29__SCAN_IN), .A(n13571), .B(
        n11851), .ZN(n11853) );
  XNOR2_X1 U14865 ( .A(n11855), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14391) );
  AOI22_X1 U14866 ( .A1(n11854), .A2(n11853), .B1(n13571), .B2(n14391), .ZN(
        n14370) );
  INV_X1 U14867 ( .A(n11855), .ZN(n11856) );
  NAND2_X1 U14868 ( .A1(n11856), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12148) );
  INV_X1 U14869 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14517) );
  XNOR2_X1 U14870 ( .A(n12148), .B(n14517), .ZN(n14812) );
  INV_X1 U14871 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11868) );
  OAI22_X1 U14872 ( .A1(n11859), .A2(n11858), .B1(n9596), .B2(n11857), .ZN(
        n11863) );
  INV_X1 U14873 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11860) );
  INV_X1 U14874 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13432) );
  OAI22_X1 U14875 ( .A1(n11861), .A2(n11860), .B1(n11028), .B2(n13432), .ZN(
        n11862) );
  AOI211_X1 U14876 ( .C1(n11864), .C2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n11863), .B(n11862), .ZN(n11867) );
  AOI22_X1 U14877 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n9602), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11866) );
  OAI211_X1 U14878 ( .C1(n11868), .C2(n13153), .A(n11867), .B(n11866), .ZN(
        n11876) );
  AOI22_X1 U14879 ( .A1(n11192), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9592), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14880 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9616), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14881 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14882 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11871) );
  NAND4_X1 U14883 ( .A1(n11874), .A2(n11873), .A3(n11872), .A4(n11871), .ZN(
        n11875) );
  NOR2_X1 U14884 ( .A1(n11876), .A2(n11875), .ZN(n11880) );
  NOR2_X1 U14885 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  XOR2_X1 U14886 ( .A(n11880), .B(n11879), .Z(n11884) );
  AOI21_X1 U14887 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n13658), .A(
        n13571), .ZN(n11882) );
  NAND2_X1 U14888 ( .A1(n11257), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11881) );
  OAI211_X1 U14889 ( .C1(n11884), .C2(n11883), .A(n11882), .B(n11881), .ZN(
        n11885) );
  OAI21_X1 U14890 ( .B1(n11319), .B2(n14812), .A(n11885), .ZN(n12039) );
  AND2_X1 U14891 ( .A1(n13066), .A2(n9726), .ZN(n11886) );
  XNOR2_X1 U14892 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11905) );
  NAND2_X1 U14893 ( .A1(n11910), .A2(n11905), .ZN(n11888) );
  NAND2_X1 U14894 ( .A1(n13532), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11887) );
  NAND2_X1 U14895 ( .A1(n11888), .A2(n11887), .ZN(n11902) );
  XNOR2_X1 U14896 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11900) );
  NAND2_X1 U14897 ( .A1(n11902), .A2(n11900), .ZN(n11890) );
  NAND2_X1 U14898 ( .A1(n16513), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11889) );
  XNOR2_X1 U14899 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11897) );
  NAND2_X1 U14900 ( .A1(n11899), .A2(n11897), .ZN(n11892) );
  NAND2_X1 U14901 ( .A1(n13870), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11891) );
  NAND2_X1 U14902 ( .A1(n11892), .A2(n11891), .ZN(n11931) );
  NAND2_X1 U14903 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11894), .ZN(
        n11930) );
  INV_X1 U14904 ( .A(n12904), .ZN(n11896) );
  INV_X1 U14905 ( .A(n11897), .ZN(n11898) );
  XNOR2_X1 U14906 ( .A(n11899), .B(n11898), .ZN(n12902) );
  INV_X1 U14907 ( .A(n12902), .ZN(n11928) );
  INV_X1 U14908 ( .A(n11900), .ZN(n11901) );
  XNOR2_X1 U14909 ( .A(n11902), .B(n11901), .ZN(n12901) );
  NAND2_X1 U14910 ( .A1(n9614), .A2(n14957), .ZN(n11903) );
  NOR2_X1 U14911 ( .A1(n11915), .A2(n11913), .ZN(n11926) );
  NAND2_X1 U14912 ( .A1(n11909), .A2(n12901), .ZN(n11904) );
  OAI211_X1 U14913 ( .C1(n12901), .C2(n11929), .A(n11913), .B(n11904), .ZN(
        n11925) );
  INV_X1 U14914 ( .A(n11905), .ZN(n11906) );
  XNOR2_X1 U14915 ( .A(n11906), .B(n11910), .ZN(n12900) );
  INV_X1 U14916 ( .A(n12900), .ZN(n11907) );
  OAI21_X1 U14917 ( .B1(n11909), .B2(n12066), .A(n11907), .ZN(n11919) );
  INV_X1 U14918 ( .A(n11919), .ZN(n11923) );
  NAND2_X1 U14919 ( .A1(n9614), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11932) );
  OAI21_X1 U14920 ( .B1(n12900), .B2(n11929), .A(n11932), .ZN(n11908) );
  AOI21_X1 U14921 ( .B1(n11909), .B2(n14978), .A(n11908), .ZN(n11922) );
  INV_X1 U14922 ( .A(n11922), .ZN(n11920) );
  INV_X1 U14923 ( .A(n11910), .ZN(n11912) );
  NAND2_X1 U14924 ( .A1(n14449), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11911) );
  NAND2_X1 U14925 ( .A1(n11912), .A2(n11911), .ZN(n11916) );
  INV_X1 U14926 ( .A(n11916), .ZN(n11914) );
  OAI211_X1 U14927 ( .C1(n14982), .C2(n13126), .A(n11914), .B(n11913), .ZN(
        n11918) );
  OAI21_X1 U14928 ( .B1(n11916), .B2(n11915), .A(n11934), .ZN(n11917) );
  OAI211_X1 U14929 ( .C1(n11920), .C2(n11919), .A(n11918), .B(n11917), .ZN(
        n11921) );
  OAI21_X1 U14930 ( .B1(n11923), .B2(n11922), .A(n11921), .ZN(n11924) );
  AOI22_X1 U14931 ( .A1(n12901), .A2(n11926), .B1(n11925), .B2(n11924), .ZN(
        n11927) );
  AOI21_X1 U14932 ( .B1(n11929), .B2(n11928), .A(n11927), .ZN(n11937) );
  NAND2_X1 U14933 ( .A1(n11932), .A2(n14978), .ZN(n11933) );
  OAI22_X1 U14934 ( .A1(n11934), .A2(n12902), .B1(n12905), .B2(n11933), .ZN(
        n11936) );
  OAI22_X1 U14935 ( .A1(n11937), .A2(n11936), .B1(n11935), .B2(n12905), .ZN(
        n11938) );
  INV_X1 U14936 ( .A(n11938), .ZN(n11939) );
  NAND2_X1 U14937 ( .A1(n14981), .A2(n14963), .ZN(n13120) );
  INV_X1 U14938 ( .A(n13297), .ZN(n14403) );
  NAND4_X1 U14939 ( .A1(n14970), .A2(n9614), .A3(n14403), .A4(n13301), .ZN(
        n11945) );
  NOR2_X1 U14940 ( .A1(n11945), .A2(n13155), .ZN(n13074) );
  NAND2_X1 U14941 ( .A1(n13074), .A2(n13066), .ZN(n11946) );
  NAND2_X1 U14942 ( .A1(n13120), .A2(n11946), .ZN(n11947) );
  AOI22_X1 U14943 ( .A1(n14503), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n9612), .B2(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14502) );
  NAND2_X2 U14944 ( .A1(n13066), .A2(n11143), .ZN(n12028) );
  OR2_X1 U14945 ( .A1(n12028), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n11951) );
  INV_X1 U14946 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20828) );
  NAND2_X1 U14947 ( .A1(n11959), .A2(n20828), .ZN(n11949) );
  OAI211_X1 U14948 ( .C1(n12010), .C2(P1_EBX_REG_1__SCAN_IN), .A(n14501), .B(
        n11949), .ZN(n11950) );
  NAND2_X1 U14949 ( .A1(n11951), .A2(n11950), .ZN(n11953) );
  NAND2_X1 U14950 ( .A1(n11959), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11952) );
  OAI21_X1 U14951 ( .B1(n11143), .B2(P1_EBX_REG_0__SCAN_IN), .A(n11952), .ZN(
        n13030) );
  XNOR2_X1 U14952 ( .A(n11953), .B(n13030), .ZN(n13067) );
  NAND2_X1 U14953 ( .A1(n13067), .A2(n13066), .ZN(n13068) );
  OR2_X1 U14954 ( .A1(n12028), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n11956) );
  INV_X1 U14955 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20822) );
  NAND2_X1 U14956 ( .A1(n11959), .A2(n20822), .ZN(n11954) );
  OAI211_X1 U14957 ( .C1(n9612), .C2(P1_EBX_REG_2__SCAN_IN), .A(n14501), .B(
        n11954), .ZN(n11955) );
  AND2_X1 U14958 ( .A1(n11956), .A2(n11955), .ZN(n13271) );
  MUX2_X1 U14959 ( .A(n12024), .B(n11143), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11958) );
  NOR2_X1 U14960 ( .A1(n14503), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11957) );
  NOR2_X1 U14961 ( .A1(n11958), .A2(n11957), .ZN(n13281) );
  MUX2_X1 U14962 ( .A(n12028), .B(n11959), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n11963) );
  INV_X1 U14963 ( .A(n11959), .ZN(n11960) );
  NAND2_X1 U14964 ( .A1(n9612), .A2(n11960), .ZN(n11985) );
  NAND2_X1 U14965 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n9612), .ZN(
        n11961) );
  AND2_X1 U14966 ( .A1(n11985), .A2(n11961), .ZN(n11962) );
  INV_X1 U14967 ( .A(n12024), .ZN(n12015) );
  NAND2_X1 U14968 ( .A1(n14501), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11964) );
  OAI211_X1 U14969 ( .C1(n9612), .C2(P1_EBX_REG_5__SCAN_IN), .A(n11959), .B(
        n11964), .ZN(n11965) );
  OAI21_X1 U14970 ( .B1(n12015), .B2(P1_EBX_REG_5__SCAN_IN), .A(n11965), .ZN(
        n16830) );
  MUX2_X1 U14971 ( .A(n12028), .B(n11959), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n11968) );
  NAND2_X1 U14972 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n9612), .ZN(
        n11966) );
  AND2_X1 U14973 ( .A1(n11985), .A2(n11966), .ZN(n11967) );
  INV_X1 U14974 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13919) );
  NAND2_X1 U14975 ( .A1(n12024), .A2(n13919), .ZN(n11971) );
  NAND2_X1 U14976 ( .A1(n14501), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11969) );
  OAI211_X1 U14977 ( .C1(n9612), .C2(P1_EBX_REG_7__SCAN_IN), .A(n11959), .B(
        n11969), .ZN(n11970) );
  AND2_X1 U14978 ( .A1(n11971), .A2(n11970), .ZN(n13916) );
  NAND2_X1 U14979 ( .A1(n13917), .A2(n13916), .ZN(n13937) );
  MUX2_X1 U14980 ( .A(n12028), .B(n11959), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n11974) );
  NAND2_X1 U14981 ( .A1(n9612), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11972) );
  AND2_X1 U14982 ( .A1(n11985), .A2(n11972), .ZN(n11973) );
  NAND2_X1 U14983 ( .A1(n14501), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11975) );
  OAI211_X1 U14984 ( .C1(n9612), .C2(P1_EBX_REG_9__SCAN_IN), .A(n11959), .B(
        n11975), .ZN(n11976) );
  OAI21_X1 U14985 ( .B1(n12015), .B2(P1_EBX_REG_9__SCAN_IN), .A(n11976), .ZN(
        n13980) );
  OR2_X1 U14986 ( .A1(n12028), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n11979) );
  INV_X1 U14987 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12132) );
  NAND2_X1 U14988 ( .A1(n11959), .A2(n12132), .ZN(n11977) );
  OAI211_X1 U14989 ( .C1(n9612), .C2(P1_EBX_REG_10__SCAN_IN), .A(n14501), .B(
        n11977), .ZN(n11978) );
  MUX2_X1 U14990 ( .A(n12024), .B(n11143), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11981) );
  NOR2_X1 U14991 ( .A1(n14503), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11980) );
  NOR2_X1 U14992 ( .A1(n11981), .A2(n11980), .ZN(n14158) );
  MUX2_X1 U14993 ( .A(n12024), .B(n11143), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11983) );
  NOR2_X1 U14994 ( .A1(n14503), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11982) );
  NOR2_X1 U14995 ( .A1(n11983), .A2(n11982), .ZN(n14722) );
  MUX2_X1 U14996 ( .A(n12028), .B(n11959), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11987) );
  NAND2_X1 U14997 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n9612), .ZN(
        n11984) );
  AND2_X1 U14998 ( .A1(n11985), .A2(n11984), .ZN(n11986) );
  NAND2_X1 U14999 ( .A1(n11987), .A2(n11986), .ZN(n14721) );
  NAND2_X1 U15000 ( .A1(n14722), .A2(n14721), .ZN(n11988) );
  OR2_X2 U15001 ( .A1(n14729), .A2(n11988), .ZN(n15128) );
  MUX2_X1 U15002 ( .A(n12024), .B(n11143), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11990) );
  NOR2_X1 U15003 ( .A1(n14503), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11989) );
  NOR2_X1 U15004 ( .A1(n11990), .A2(n11989), .ZN(n14711) );
  OR2_X1 U15005 ( .A1(n12028), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n11993) );
  INV_X1 U15006 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16741) );
  NAND2_X1 U15007 ( .A1(n11959), .A2(n16741), .ZN(n11991) );
  OAI211_X1 U15008 ( .C1(n9612), .C2(P1_EBX_REG_14__SCAN_IN), .A(n14501), .B(
        n11991), .ZN(n11992) );
  NAND2_X1 U15009 ( .A1(n11993), .A2(n11992), .ZN(n15127) );
  NAND2_X1 U15010 ( .A1(n14711), .A2(n15127), .ZN(n11994) );
  NOR2_X2 U15011 ( .A1(n15128), .A2(n11994), .ZN(n14713) );
  OR2_X1 U15012 ( .A1(n12028), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n11997) );
  INV_X1 U15013 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16742) );
  NAND2_X1 U15014 ( .A1(n11959), .A2(n16742), .ZN(n11995) );
  OAI211_X1 U15015 ( .C1(n9612), .C2(P1_EBX_REG_16__SCAN_IN), .A(n14501), .B(
        n11995), .ZN(n11996) );
  NAND2_X1 U15016 ( .A1(n11997), .A2(n11996), .ZN(n14702) );
  MUX2_X1 U15017 ( .A(n12024), .B(n11143), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11999) );
  NOR2_X1 U15018 ( .A1(n14503), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11998) );
  NOR2_X1 U15019 ( .A1(n11999), .A2(n11998), .ZN(n14645) );
  OR2_X1 U15020 ( .A1(n12028), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n12002) );
  INV_X1 U15021 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16729) );
  NAND2_X1 U15022 ( .A1(n11959), .A2(n16729), .ZN(n12000) );
  OAI211_X1 U15023 ( .C1(n9612), .C2(P1_EBX_REG_18__SCAN_IN), .A(n14501), .B(
        n12000), .ZN(n12001) );
  MUX2_X1 U15024 ( .A(n12024), .B(n11143), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12003) );
  INV_X1 U15025 ( .A(n12003), .ZN(n12005) );
  INV_X1 U15026 ( .A(n14503), .ZN(n13032) );
  INV_X1 U15027 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16717) );
  NAND2_X1 U15028 ( .A1(n13032), .A2(n16717), .ZN(n12004) );
  NAND2_X1 U15029 ( .A1(n12005), .A2(n12004), .ZN(n14635) );
  MUX2_X1 U15030 ( .A(n12028), .B(n11959), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12007) );
  NAND2_X1 U15031 ( .A1(n9612), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12006) );
  MUX2_X1 U15032 ( .A(n12024), .B(n11143), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12009) );
  NOR2_X1 U15033 ( .A1(n14503), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12008) );
  NOR2_X1 U15034 ( .A1(n12009), .A2(n12008), .ZN(n14618) );
  MUX2_X1 U15035 ( .A(n12028), .B(n11959), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12012) );
  NAND2_X1 U15036 ( .A1(n9612), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12011) );
  AND2_X1 U15037 ( .A1(n12012), .A2(n12011), .ZN(n14605) );
  NAND2_X1 U15038 ( .A1(n14501), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12013) );
  OAI211_X1 U15039 ( .C1(n9612), .C2(P1_EBX_REG_23__SCAN_IN), .A(n11959), .B(
        n12013), .ZN(n12014) );
  OAI21_X1 U15040 ( .B1(n12015), .B2(P1_EBX_REG_23__SCAN_IN), .A(n12014), .ZN(
        n14593) );
  NOR2_X2 U15041 ( .A1(n9652), .A2(n14593), .ZN(n14592) );
  OR2_X1 U15042 ( .A1(n12028), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n12018) );
  INV_X1 U15043 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12140) );
  NAND2_X1 U15044 ( .A1(n11959), .A2(n12140), .ZN(n12016) );
  OAI211_X1 U15045 ( .C1(n9612), .C2(P1_EBX_REG_24__SCAN_IN), .A(n14501), .B(
        n12016), .ZN(n12017) );
  NAND2_X1 U15046 ( .A1(n12018), .A2(n12017), .ZN(n14581) );
  MUX2_X1 U15047 ( .A(n12024), .B(n11143), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12020) );
  NOR2_X1 U15048 ( .A1(n14503), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12019) );
  NOR2_X1 U15049 ( .A1(n12020), .A2(n12019), .ZN(n14570) );
  OR2_X1 U15050 ( .A1(n12028), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n12023) );
  INV_X1 U15051 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14850) );
  NAND2_X1 U15052 ( .A1(n11959), .A2(n14850), .ZN(n12021) );
  OAI211_X1 U15053 ( .C1(n9612), .C2(P1_EBX_REG_26__SCAN_IN), .A(n14501), .B(
        n12021), .ZN(n12022) );
  AND2_X1 U15054 ( .A1(n12023), .A2(n12022), .ZN(n14553) );
  MUX2_X1 U15055 ( .A(n12024), .B(n11143), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12025) );
  INV_X1 U15056 ( .A(n12025), .ZN(n12027) );
  INV_X1 U15057 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15048) );
  NAND2_X1 U15058 ( .A1(n13032), .A2(n15048), .ZN(n12026) );
  NAND2_X1 U15059 ( .A1(n12027), .A2(n12026), .ZN(n14537) );
  OR2_X1 U15060 ( .A1(n12028), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n12031) );
  INV_X1 U15061 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14828) );
  NAND2_X1 U15062 ( .A1(n11959), .A2(n14828), .ZN(n12029) );
  OAI211_X1 U15063 ( .C1(n9612), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14501), .B(
        n12029), .ZN(n12030) );
  NAND2_X1 U15064 ( .A1(n12031), .A2(n12030), .ZN(n14526) );
  NAND2_X2 U15065 ( .A1(n14539), .A2(n14526), .ZN(n14525) );
  OR2_X1 U15066 ( .A1(n9612), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12032) );
  OAI21_X1 U15067 ( .B1(n14503), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12032), .ZN(n12033) );
  MUX2_X1 U15068 ( .A(n12033), .B(n12032), .S(n11143), .Z(n14381) );
  OR2_X2 U15069 ( .A1(n14525), .A2(n14381), .ZN(n14500) );
  INV_X1 U15070 ( .A(n14500), .ZN(n12034) );
  OAI22_X1 U15071 ( .A1(n12034), .A2(n14501), .B1(n12033), .B2(n14525), .ZN(
        n12035) );
  INV_X1 U15072 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n12036) );
  OAI21_X1 U15073 ( .B1(n15025), .B2(n14730), .A(n10194), .ZN(n12037) );
  INV_X1 U15074 ( .A(n12037), .ZN(n12038) );
  AOI22_X1 U15075 ( .A1(n11257), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12040), .ZN(n12041) );
  XNOR2_X1 U15076 ( .A(n12042), .B(n12041), .ZN(n14515) );
  NAND3_X1 U15077 ( .A1(n20963), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16846) );
  INV_X1 U15078 ( .A(n16846), .ZN(n12043) );
  INV_X2 U15079 ( .A(n21063), .ZN(n20791) );
  NAND2_X1 U15080 ( .A1(n14515), .A2(n20791), .ZN(n12153) );
  NAND2_X1 U15081 ( .A1(n12044), .A2(n12116), .ZN(n12045) );
  NOR2_X1 U15082 ( .A1(n12045), .A2(n12066), .ZN(n12046) );
  INV_X4 U15083 ( .A(n15123), .ZN(n16656) );
  NAND2_X1 U15084 ( .A1(n16656), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14816) );
  INV_X1 U15085 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15000) );
  NOR2_X1 U15086 ( .A1(n14816), .A2(n15000), .ZN(n12143) );
  OR2_X1 U15087 ( .A1(n16656), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14817) );
  NOR2_X1 U15088 ( .A1(n14817), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12142) );
  NAND2_X1 U15089 ( .A1(n14982), .A2(n13288), .ZN(n12062) );
  OAI21_X1 U15090 ( .B1(n16528), .B2(n12051), .A(n12062), .ZN(n12048) );
  INV_X1 U15091 ( .A(n12048), .ZN(n12049) );
  NAND2_X1 U15092 ( .A1(n13093), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12057) );
  OR2_X1 U15093 ( .A1(n12050), .A2(n12066), .ZN(n12056) );
  NAND2_X1 U15094 ( .A1(n12051), .A2(n12052), .ZN(n12071) );
  OAI21_X1 U15095 ( .B1(n12052), .B2(n12051), .A(n12071), .ZN(n12053) );
  OAI211_X1 U15096 ( .C1(n12053), .C2(n16528), .A(n9726), .B(n11116), .ZN(
        n12054) );
  INV_X1 U15097 ( .A(n12054), .ZN(n12055) );
  NAND2_X1 U15098 ( .A1(n12056), .A2(n12055), .ZN(n12058) );
  XNOR2_X1 U15099 ( .A(n12057), .B(n12058), .ZN(n13486) );
  NAND2_X1 U15100 ( .A1(n13486), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20832) );
  INV_X1 U15101 ( .A(n12057), .ZN(n13094) );
  NAND2_X1 U15102 ( .A1(n13094), .A2(n12058), .ZN(n12059) );
  NAND2_X1 U15103 ( .A1(n20832), .A2(n12059), .ZN(n12067) );
  XNOR2_X1 U15104 ( .A(n12067), .B(n20822), .ZN(n13968) );
  INV_X1 U15105 ( .A(n12061), .ZN(n12070) );
  XNOR2_X1 U15106 ( .A(n12071), .B(n12070), .ZN(n12064) );
  INV_X1 U15107 ( .A(n12062), .ZN(n12063) );
  AOI21_X1 U15108 ( .B1(n12117), .B2(n12064), .A(n12063), .ZN(n12065) );
  OAI21_X1 U15109 ( .B1(n12060), .B2(n12066), .A(n12065), .ZN(n13967) );
  NAND2_X1 U15110 ( .A1(n13968), .A2(n13967), .ZN(n13966) );
  NAND2_X1 U15111 ( .A1(n12067), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12068) );
  NAND2_X1 U15112 ( .A1(n13966), .A2(n12068), .ZN(n13959) );
  NAND2_X1 U15113 ( .A1(n12071), .A2(n12070), .ZN(n12081) );
  INV_X1 U15114 ( .A(n12080), .ZN(n12072) );
  XNOR2_X1 U15115 ( .A(n12081), .B(n12072), .ZN(n12073) );
  NAND2_X1 U15116 ( .A1(n12073), .A2(n12117), .ZN(n12074) );
  NAND2_X1 U15117 ( .A1(n12075), .A2(n12074), .ZN(n12077) );
  INV_X1 U15118 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12076) );
  XNOR2_X1 U15119 ( .A(n12077), .B(n12076), .ZN(n13958) );
  NAND2_X1 U15120 ( .A1(n13959), .A2(n13958), .ZN(n13957) );
  NAND2_X1 U15121 ( .A1(n12077), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12078) );
  NAND2_X1 U15122 ( .A1(n13957), .A2(n12078), .ZN(n20788) );
  NAND2_X1 U15123 ( .A1(n12079), .A2(n12105), .ZN(n12084) );
  NAND2_X1 U15124 ( .A1(n12081), .A2(n12080), .ZN(n12089) );
  XNOR2_X1 U15125 ( .A(n12089), .B(n12090), .ZN(n12082) );
  NAND2_X1 U15126 ( .A1(n12082), .A2(n12117), .ZN(n12083) );
  NAND2_X1 U15127 ( .A1(n12084), .A2(n12083), .ZN(n12086) );
  INV_X1 U15128 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12085) );
  XNOR2_X1 U15129 ( .A(n12086), .B(n12085), .ZN(n20787) );
  NAND2_X1 U15130 ( .A1(n20788), .A2(n20787), .ZN(n20786) );
  NAND2_X1 U15131 ( .A1(n12086), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12087) );
  NAND2_X1 U15132 ( .A1(n20786), .A2(n12087), .ZN(n16698) );
  NAND2_X1 U15133 ( .A1(n12088), .A2(n12105), .ZN(n12094) );
  INV_X1 U15134 ( .A(n12089), .ZN(n12091) );
  NAND2_X1 U15135 ( .A1(n12091), .A2(n12090), .ZN(n12098) );
  XNOR2_X1 U15136 ( .A(n12098), .B(n12099), .ZN(n12092) );
  NAND2_X1 U15137 ( .A1(n12092), .A2(n12117), .ZN(n12093) );
  NAND2_X1 U15138 ( .A1(n12094), .A2(n12093), .ZN(n12095) );
  INV_X1 U15139 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14980) );
  XNOR2_X1 U15140 ( .A(n12095), .B(n14980), .ZN(n16697) );
  NAND2_X1 U15141 ( .A1(n12095), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12096) );
  NAND2_X1 U15142 ( .A1(n12097), .A2(n12105), .ZN(n12103) );
  INV_X1 U15143 ( .A(n12098), .ZN(n12100) );
  NAND2_X1 U15144 ( .A1(n12100), .A2(n12099), .ZN(n12109) );
  XNOR2_X1 U15145 ( .A(n12109), .B(n12107), .ZN(n12101) );
  NAND2_X1 U15146 ( .A1(n12101), .A2(n12117), .ZN(n12102) );
  INV_X1 U15147 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16808) );
  NAND2_X1 U15148 ( .A1(n12106), .A2(n12105), .ZN(n12112) );
  INV_X1 U15149 ( .A(n12107), .ZN(n12108) );
  OR2_X1 U15150 ( .A1(n12109), .A2(n12108), .ZN(n12115) );
  XNOR2_X1 U15151 ( .A(n12115), .B(n12116), .ZN(n12110) );
  NAND2_X1 U15152 ( .A1(n12110), .A2(n12117), .ZN(n12111) );
  NAND2_X1 U15153 ( .A1(n12112), .A2(n12111), .ZN(n12113) );
  INV_X1 U15154 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16821) );
  XNOR2_X1 U15155 ( .A(n12113), .B(n16821), .ZN(n16684) );
  NAND2_X1 U15156 ( .A1(n16685), .A2(n16684), .ZN(n16683) );
  NAND2_X1 U15157 ( .A1(n12113), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12114) );
  NAND2_X1 U15158 ( .A1(n16683), .A2(n12114), .ZN(n14136) );
  INV_X1 U15159 ( .A(n12115), .ZN(n12118) );
  NAND3_X1 U15160 ( .A1(n12118), .A2(n12117), .A3(n12116), .ZN(n12119) );
  NAND2_X1 U15161 ( .A1(n16656), .A2(n12119), .ZN(n12120) );
  INV_X1 U15162 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16815) );
  XNOR2_X1 U15163 ( .A(n12120), .B(n16815), .ZN(n14135) );
  NAND2_X1 U15164 ( .A1(n14136), .A2(n14135), .ZN(n14134) );
  NAND2_X1 U15165 ( .A1(n12120), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12121) );
  XNOR2_X1 U15166 ( .A(n16656), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14150) );
  INV_X1 U15167 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16779) );
  XNOR2_X1 U15168 ( .A(n9588), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14939) );
  INV_X1 U15169 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15154) );
  NAND2_X1 U15170 ( .A1(n12138), .A2(n15154), .ZN(n14938) );
  NAND2_X1 U15171 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14934) );
  NAND2_X1 U15172 ( .A1(n9588), .A2(n14934), .ZN(n12123) );
  AND2_X1 U15173 ( .A1(n14938), .A2(n12123), .ZN(n12124) );
  NAND2_X1 U15174 ( .A1(n14939), .A2(n12124), .ZN(n15120) );
  AND2_X1 U15175 ( .A1(n9588), .A2(n16741), .ZN(n12125) );
  NOR2_X1 U15176 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12126) );
  INV_X1 U15177 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12128) );
  OR2_X1 U15178 ( .A1(n9588), .A2(n12128), .ZN(n12127) );
  AND2_X1 U15179 ( .A1(n12134), .A2(n12127), .ZN(n14922) );
  XNOR2_X1 U15180 ( .A(n9588), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16658) );
  NAND2_X1 U15181 ( .A1(n9588), .A2(n12128), .ZN(n12129) );
  NAND2_X1 U15182 ( .A1(n16658), .A2(n12129), .ZN(n16657) );
  AOI21_X1 U15183 ( .B1(n16653), .B2(n14922), .A(n16657), .ZN(n14923) );
  INV_X1 U15184 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14927) );
  NAND2_X1 U15185 ( .A1(n16656), .A2(n14927), .ZN(n12130) );
  AND2_X1 U15186 ( .A1(n14923), .A2(n12130), .ZN(n12131) );
  AND3_X1 U15187 ( .A1(n12132), .A2(n15154), .A3(n16776), .ZN(n12133) );
  NAND2_X1 U15188 ( .A1(n15121), .A2(n12134), .ZN(n16654) );
  NOR2_X1 U15189 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16739) );
  AND2_X1 U15190 ( .A1(n16739), .A2(n14927), .ZN(n12135) );
  NOR2_X1 U15191 ( .A1(n16656), .A2(n12135), .ZN(n12136) );
  NOR2_X1 U15192 ( .A1(n16654), .A2(n12136), .ZN(n12137) );
  XNOR2_X1 U15193 ( .A(n16656), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14914) );
  NAND2_X1 U15194 ( .A1(n14915), .A2(n14914), .ZN(n14913) );
  INV_X1 U15195 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15110) );
  INV_X1 U15196 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15103) );
  NAND2_X1 U15197 ( .A1(n12141), .A2(n14882), .ZN(n14865) );
  INV_X1 U15198 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15067) );
  INV_X1 U15199 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15089) );
  NAND3_X1 U15200 ( .A1(n15067), .A2(n12140), .A3(n15089), .ZN(n14826) );
  NOR2_X1 U15201 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15037) );
  NAND3_X1 U15202 ( .A1(n14849), .A2(n15037), .A3(n14836), .ZN(n14808) );
  AND2_X1 U15203 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14996) );
  NAND2_X1 U15204 ( .A1(n14996), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15009) );
  AND2_X1 U15205 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15038) );
  NAND2_X1 U15206 ( .A1(n11531), .A2(n14982), .ZN(n12144) );
  OR2_X1 U15207 ( .A1(n13115), .A2(n13126), .ZN(n16520) );
  NAND2_X1 U15208 ( .A1(n20893), .A2(n12150), .ZN(n21050) );
  NAND2_X1 U15209 ( .A1(n21050), .A2(n20963), .ZN(n12146) );
  NAND2_X1 U15210 ( .A1(n20963), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16527) );
  NAND2_X1 U15211 ( .A1(n20640), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12147) );
  AND2_X1 U15212 ( .A1(n16527), .A2(n12147), .ZN(n13097) );
  XNOR2_X1 U15213 ( .A(n12149), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13584) );
  INV_X1 U15214 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21030) );
  NOR2_X1 U15215 ( .A1(n16817), .A2(n21030), .ZN(n15002) );
  INV_X1 U15216 ( .A(n21061), .ZN(n14947) );
  INV_X1 U15217 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14509) );
  NOR2_X1 U15218 ( .A1(n14947), .A2(n14509), .ZN(n12151) );
  AOI211_X1 U15219 ( .C1(n16669), .C2(n13584), .A(n15002), .B(n12151), .ZN(
        n12152) );
  NAND2_X1 U15220 ( .A1(n12153), .A2(n9667), .ZN(P1_U2968) );
  NAND2_X1 U15221 ( .A1(n10150), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12183) );
  NAND2_X1 U15222 ( .A1(n12177), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12154) );
  NAND2_X1 U15223 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20615), .ZN(
        n20257) );
  NAND2_X1 U15224 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20605), .ZN(
        n20221) );
  NAND2_X1 U15225 ( .A1(n20257), .A2(n20221), .ZN(n20051) );
  NAND2_X1 U15226 ( .A1(n20585), .A2(n20051), .ZN(n20262) );
  NAND2_X1 U15227 ( .A1(n12154), .A2(n20262), .ZN(n12155) );
  AOI22_X1 U15228 ( .A1(n12177), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20585), .B2(n20615), .ZN(n12156) );
  NAND2_X1 U15229 ( .A1(n12514), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12158) );
  INV_X1 U15230 ( .A(n14090), .ZN(n12159) );
  NAND2_X1 U15231 ( .A1(n12159), .A2(n12158), .ZN(n12160) );
  NAND2_X1 U15232 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20286) );
  NAND2_X1 U15233 ( .A1(n20286), .A2(n20597), .ZN(n12162) );
  NOR2_X1 U15234 ( .A1(n20597), .A2(n20605), .ZN(n20393) );
  NAND2_X1 U15235 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20393), .ZN(
        n12173) );
  NAND2_X1 U15236 ( .A1(n12162), .A2(n12173), .ZN(n20052) );
  NAND2_X1 U15237 ( .A1(n12177), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12163) );
  OAI21_X1 U15238 ( .B1(n20052), .B2(n20578), .A(n12163), .ZN(n12164) );
  NAND2_X1 U15239 ( .A1(n12514), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12166) );
  NAND2_X1 U15240 ( .A1(n12165), .A2(n12166), .ZN(n13059) );
  INV_X1 U15241 ( .A(n12165), .ZN(n12168) );
  INV_X1 U15242 ( .A(n12166), .ZN(n12167) );
  NAND2_X1 U15243 ( .A1(n12168), .A2(n12167), .ZN(n13058) );
  INV_X1 U15244 ( .A(n13058), .ZN(n12169) );
  NOR2_X1 U15245 ( .A1(n12170), .A2(n12169), .ZN(n12171) );
  INV_X1 U15246 ( .A(n12171), .ZN(n13086) );
  NAND2_X1 U15247 ( .A1(n10549), .A2(n12172), .ZN(n12179) );
  INV_X1 U15248 ( .A(n12173), .ZN(n12174) );
  NAND2_X1 U15249 ( .A1(n12174), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20423) );
  OAI211_X1 U15250 ( .C1(n12174), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n20423), .B(n20585), .ZN(n12175) );
  INV_X1 U15251 ( .A(n12175), .ZN(n12176) );
  AOI21_X1 U15252 ( .B1(n12177), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12176), .ZN(n12178) );
  NAND2_X1 U15253 ( .A1(n12179), .A2(n12178), .ZN(n12181) );
  INV_X1 U15254 ( .A(n12514), .ZN(n12543) );
  NOR2_X1 U15255 ( .A1(n12543), .A2(n19950), .ZN(n12180) );
  NAND2_X1 U15256 ( .A1(n12181), .A2(n12180), .ZN(n12186) );
  OR2_X1 U15257 ( .A1(n12181), .A2(n12180), .ZN(n12182) );
  NAND2_X1 U15258 ( .A1(n13086), .A2(n13087), .ZN(n13090) );
  INV_X1 U15259 ( .A(n12183), .ZN(n12184) );
  NAND2_X1 U15260 ( .A1(n12184), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12185) );
  AND2_X1 U15261 ( .A1(n12186), .A2(n12185), .ZN(n12187) );
  NAND2_X1 U15262 ( .A1(n13090), .A2(n12187), .ZN(n19746) );
  NOR2_X1 U15263 ( .A1(n12543), .A2(n19956), .ZN(n19745) );
  NAND2_X1 U15264 ( .A1(n19746), .A2(n19745), .ZN(n13100) );
  INV_X1 U15265 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12188) );
  INV_X1 U15266 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n20403) );
  OAI22_X1 U15267 ( .A1(n12272), .A2(n12188), .B1(n12315), .B2(n20403), .ZN(
        n12189) );
  INV_X1 U15268 ( .A(n12189), .ZN(n12193) );
  AOI22_X1 U15269 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12424), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15270 ( .A1(n12202), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15271 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12190) );
  NAND4_X1 U15272 ( .A1(n12193), .A2(n12192), .A3(n12191), .A4(n12190), .ZN(
        n12201) );
  AOI22_X1 U15273 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15274 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12366), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12198) );
  INV_X1 U15275 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U15276 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12429), .ZN(
        n12194) );
  OAI21_X1 U15277 ( .B1(n12431), .B2(n12412), .A(n12194), .ZN(n12195) );
  AOI21_X1 U15278 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n12195), .ZN(n12197) );
  NAND2_X1 U15279 ( .A1(n12384), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12196) );
  NAND4_X1 U15280 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12196), .ZN(
        n12200) );
  INV_X1 U15281 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16240) );
  NAND2_X1 U15282 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13187) );
  NOR2_X1 U15283 ( .A1(n16240), .A2(n13187), .ZN(n19785) );
  INV_X1 U15284 ( .A(n12202), .ZN(n12316) );
  OAI22_X1 U15285 ( .A1(n12443), .A2(n12316), .B1(n12315), .B2(n12452), .ZN(
        n12203) );
  INV_X1 U15286 ( .A(n12203), .ZN(n12207) );
  AOI22_X1 U15287 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15288 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15289 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12204) );
  NAND4_X1 U15290 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12215) );
  AOI22_X1 U15291 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12368), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15292 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12366), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U15293 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12429), .ZN(
        n12208) );
  OAI21_X1 U15294 ( .B1(n12431), .B2(n12441), .A(n12208), .ZN(n12209) );
  AOI21_X1 U15295 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n12209), .ZN(n12211) );
  NAND2_X1 U15296 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12210) );
  NAND4_X1 U15297 ( .A1(n12213), .A2(n12212), .A3(n12211), .A4(n12210), .ZN(
        n12214) );
  NOR2_X1 U15298 ( .A1(n12215), .A2(n12214), .ZN(n13364) );
  AOI22_X1 U15299 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12202), .B1(
        n12423), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15300 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15301 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15302 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12217) );
  NAND4_X1 U15303 ( .A1(n12220), .A2(n12219), .A3(n12218), .A4(n12217), .ZN(
        n12228) );
  AOI22_X1 U15304 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12368), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15305 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12366), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12225) );
  NAND2_X1 U15306 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12429), .ZN(
        n12221) );
  OAI21_X1 U15307 ( .B1(n12431), .B2(n12495), .A(n12221), .ZN(n12222) );
  AOI21_X1 U15308 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n12222), .ZN(n12224) );
  NAND2_X1 U15309 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12223) );
  NAND4_X1 U15310 ( .A1(n12226), .A2(n12225), .A3(n12224), .A4(n12223), .ZN(
        n12227) );
  INV_X1 U15311 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12477) );
  INV_X1 U15312 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12229) );
  OAI22_X1 U15313 ( .A1(n12477), .A2(n12272), .B1(n12315), .B2(n12229), .ZN(
        n12230) );
  INV_X1 U15314 ( .A(n12230), .ZN(n12234) );
  AOI22_X1 U15315 ( .A1(n12202), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15316 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15317 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12368), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12231) );
  NAND4_X1 U15318 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12231), .ZN(
        n12243) );
  AOI22_X1 U15319 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n12351), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15320 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10560), .B1(
        n12366), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12240) );
  INV_X1 U15321 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12236) );
  NAND2_X1 U15322 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12429), .ZN(
        n12235) );
  OAI21_X1 U15323 ( .B1(n12431), .B2(n12236), .A(n12235), .ZN(n12237) );
  AOI21_X1 U15324 ( .B1(n12365), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n12237), .ZN(n12239) );
  NAND2_X1 U15325 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12238) );
  NAND4_X1 U15326 ( .A1(n12241), .A2(n12240), .A3(n12239), .A4(n12238), .ZN(
        n12242) );
  AOI22_X1 U15327 ( .A1(n12202), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12423), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15328 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15329 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15330 ( .A1(n12424), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12244) );
  NAND4_X1 U15331 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n12255) );
  AOI22_X1 U15332 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15333 ( .A1(n12366), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12252) );
  INV_X1 U15334 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12413) );
  NAND2_X1 U15335 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n12429), .ZN(
        n12248) );
  OAI21_X1 U15336 ( .B1(n12431), .B2(n12413), .A(n12248), .ZN(n12249) );
  AOI21_X1 U15337 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n12249), .ZN(n12251) );
  NAND2_X1 U15338 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12250) );
  NAND4_X1 U15339 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12254) );
  OR2_X1 U15340 ( .A1(n12255), .A2(n12254), .ZN(n19763) );
  INV_X1 U15341 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12257) );
  INV_X1 U15342 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12256) );
  OAI22_X1 U15343 ( .A1(n12257), .A2(n12316), .B1(n12315), .B2(n12256), .ZN(
        n12258) );
  INV_X1 U15344 ( .A(n12258), .ZN(n12262) );
  AOI22_X1 U15345 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15346 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15347 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12259) );
  NAND4_X1 U15348 ( .A1(n12262), .A2(n12261), .A3(n12260), .A4(n12259), .ZN(
        n12271) );
  AOI22_X1 U15349 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12368), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15350 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12366), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12268) );
  INV_X1 U15351 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12264) );
  NAND2_X1 U15352 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12429), .ZN(
        n12263) );
  OAI21_X1 U15353 ( .B1(n12431), .B2(n12264), .A(n12263), .ZN(n12265) );
  AOI21_X1 U15354 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n12265), .ZN(n12267) );
  NAND2_X1 U15355 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12266) );
  NAND4_X1 U15356 ( .A1(n12269), .A2(n12268), .A3(n12267), .A4(n12266), .ZN(
        n12270) );
  NOR2_X1 U15357 ( .A1(n12271), .A2(n12270), .ZN(n15588) );
  INV_X1 U15358 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12576) );
  OAI22_X1 U15359 ( .A1(n12576), .A2(n12315), .B1(n12272), .B2(n12582), .ZN(
        n12273) );
  INV_X1 U15360 ( .A(n12273), .ZN(n12277) );
  AOI22_X1 U15361 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15362 ( .A1(n12202), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15363 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12274) );
  NAND4_X1 U15364 ( .A1(n12277), .A2(n12276), .A3(n12275), .A4(n12274), .ZN(
        n12285) );
  AOI22_X1 U15365 ( .A1(n12351), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12366), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15366 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10295), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12282) );
  NAND2_X1 U15367 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12429), .ZN(
        n12278) );
  OAI21_X1 U15368 ( .B1(n12431), .B2(n12569), .A(n12278), .ZN(n12279) );
  AOI21_X1 U15369 ( .B1(n12368), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n12279), .ZN(n12281) );
  NAND2_X1 U15370 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12280) );
  NAND4_X1 U15371 ( .A1(n12283), .A2(n12282), .A3(n12281), .A4(n12280), .ZN(
        n12284) );
  NOR2_X1 U15372 ( .A1(n12285), .A2(n12284), .ZN(n19769) );
  OR2_X1 U15373 ( .A1(n15588), .A2(n19769), .ZN(n12299) );
  OAI22_X1 U15374 ( .A1(n12316), .A2(n12549), .B1(n12315), .B2(n12559), .ZN(
        n12286) );
  INV_X1 U15375 ( .A(n12286), .ZN(n12290) );
  AOI22_X1 U15376 ( .A1(n12424), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15377 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15378 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12287) );
  NAND4_X1 U15379 ( .A1(n12290), .A2(n12289), .A3(n12288), .A4(n12287), .ZN(
        n12298) );
  AOI22_X1 U15380 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15381 ( .A1(n12366), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12295) );
  INV_X1 U15382 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U15383 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12429), .ZN(
        n12291) );
  OAI21_X1 U15384 ( .B1(n12431), .B2(n12547), .A(n12291), .ZN(n12292) );
  AOI21_X1 U15385 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n12292), .ZN(n12294) );
  NAND2_X1 U15386 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12293) );
  NAND4_X1 U15387 ( .A1(n12296), .A2(n12295), .A3(n12294), .A4(n12293), .ZN(
        n12297) );
  NOR2_X1 U15388 ( .A1(n12298), .A2(n12297), .ZN(n13848) );
  NOR2_X1 U15389 ( .A1(n12299), .A2(n13848), .ZN(n15585) );
  AOI22_X1 U15390 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12421), .B1(
        n12423), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U15391 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n12365), .ZN(n12302) );
  AOI22_X1 U15392 ( .A1(n12202), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15393 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12300) );
  NAND4_X1 U15394 ( .A1(n12303), .A2(n12302), .A3(n12301), .A4(n12300), .ZN(
        n12311) );
  AOI22_X1 U15395 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12368), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15396 ( .A1(n12351), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12366), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12308) );
  INV_X1 U15397 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15398 ( .A1(n12389), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12429), .ZN(n12304) );
  OAI21_X1 U15399 ( .B1(n10565), .B2(n12531), .A(n12304), .ZN(n12305) );
  INV_X1 U15400 ( .A(n12305), .ZN(n12307) );
  NAND2_X1 U15401 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12306) );
  NAND4_X1 U15402 ( .A1(n12309), .A2(n12308), .A3(n12307), .A4(n12306), .ZN(
        n12310) );
  INV_X1 U15403 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12314) );
  OAI22_X1 U15404 ( .A1(n12317), .A2(n12316), .B1(n12315), .B2(n12314), .ZN(
        n12318) );
  INV_X1 U15405 ( .A(n12318), .ZN(n12322) );
  AOI22_X1 U15406 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15407 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15408 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12319) );
  NAND4_X1 U15409 ( .A1(n12322), .A2(n12321), .A3(n12320), .A4(n12319), .ZN(
        n12330) );
  AOI22_X1 U15410 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12368), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15411 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12365), .B1(
        n12366), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12327) );
  NAND2_X1 U15412 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12429), .ZN(
        n12323) );
  OAI21_X1 U15413 ( .B1(n12431), .B2(n13866), .A(n12323), .ZN(n12324) );
  AOI21_X1 U15414 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n12324), .ZN(n12326) );
  NAND2_X1 U15415 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12325) );
  NAND4_X1 U15416 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(
        n12329) );
  NOR2_X1 U15417 ( .A1(n12330), .A2(n12329), .ZN(n14097) );
  NAND2_X1 U15418 ( .A1(n12332), .A2(n12331), .ZN(n16911) );
  AOI22_X1 U15419 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12202), .B1(
        n12423), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15420 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15421 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15422 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12333) );
  NAND4_X1 U15423 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        n12345) );
  AOI22_X1 U15424 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12368), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15425 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12365), .B1(
        n12366), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12342) );
  INV_X1 U15426 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12338) );
  NAND2_X1 U15427 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12429), .ZN(
        n12337) );
  OAI21_X1 U15428 ( .B1(n12431), .B2(n12338), .A(n12337), .ZN(n12339) );
  AOI21_X1 U15429 ( .B1(n12351), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n12339), .ZN(n12341) );
  NAND2_X1 U15430 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12340) );
  NAND4_X1 U15431 ( .A1(n12343), .A2(n12342), .A3(n12341), .A4(n12340), .ZN(
        n12344) );
  NOR2_X1 U15432 ( .A1(n12345), .A2(n12344), .ZN(n16910) );
  AOI22_X1 U15433 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12202), .B1(
        n12423), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15434 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U15435 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12347) );
  INV_X1 U15436 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20410) );
  AOI22_X1 U15437 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12346) );
  AND4_X1 U15438 ( .A1(n12349), .A2(n12348), .A3(n12347), .A4(n12346), .ZN(
        n12357) );
  OAI22_X1 U15439 ( .A1(n10579), .A2(n12431), .B1(n12495), .B2(n12350), .ZN(
        n12353) );
  INV_X1 U15440 ( .A(n12351), .ZN(n12378) );
  INV_X1 U15441 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12505) );
  NOR2_X1 U15442 ( .A1(n12378), .A2(n12505), .ZN(n12352) );
  AOI211_X1 U15443 ( .C1(n12433), .C2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n12353), .B(n12352), .ZN(n12356) );
  AOI22_X1 U15444 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12368), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15445 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12365), .B1(
        n12366), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12354) );
  NAND4_X1 U15446 ( .A1(n12357), .A2(n12356), .A3(n12355), .A4(n12354), .ZN(
        n15568) );
  AOI22_X1 U15447 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12202), .B1(
        n12423), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15448 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15449 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15450 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12358) );
  NAND4_X1 U15451 ( .A1(n12361), .A2(n12360), .A3(n12359), .A4(n12358), .ZN(
        n12372) );
  INV_X1 U15452 ( .A(n12433), .ZN(n12392) );
  INV_X1 U15453 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12364) );
  NAND2_X1 U15454 ( .A1(n12351), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12363) );
  AOI22_X1 U15455 ( .A1(n12389), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12429), .ZN(n12362) );
  OAI211_X1 U15456 ( .C1(n12392), .C2(n12364), .A(n12363), .B(n12362), .ZN(
        n12371) );
  INV_X1 U15457 ( .A(n12365), .ZN(n12395) );
  INV_X1 U15458 ( .A(n12366), .ZN(n12394) );
  INV_X1 U15459 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12367) );
  OAI22_X1 U15460 ( .A1(n19956), .A2(n12395), .B1(n12394), .B2(n12367), .ZN(
        n12370) );
  INV_X1 U15461 ( .A(n12368), .ZN(n12397) );
  INV_X1 U15462 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12522) );
  INV_X1 U15463 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12533) );
  OAI22_X1 U15464 ( .A1(n12397), .A2(n12522), .B1(n10565), .B2(n12533), .ZN(
        n12369) );
  NOR4_X1 U15465 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n16907) );
  AOI22_X1 U15466 ( .A1(n12202), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12423), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15467 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15468 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15469 ( .A1(n12424), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12373) );
  AND4_X1 U15470 ( .A1(n12376), .A2(n12375), .A3(n12374), .A4(n12373), .ZN(
        n12383) );
  INV_X1 U15471 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15472 ( .A1(n12389), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12377) );
  OAI21_X1 U15473 ( .B1(n12378), .B2(n12557), .A(n12377), .ZN(n12379) );
  AOI21_X1 U15474 ( .B1(n12433), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n12379), .ZN(n12382) );
  AOI22_X1 U15475 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15476 ( .A1(n12366), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12380) );
  NAND4_X1 U15477 ( .A1(n12383), .A2(n12382), .A3(n12381), .A4(n12380), .ZN(
        n15563) );
  AOI22_X1 U15478 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12202), .B1(
        n12423), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U15479 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15480 ( .A1(n12421), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15481 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12385) );
  NAND4_X1 U15482 ( .A1(n12388), .A2(n12387), .A3(n12386), .A4(n12385), .ZN(
        n12401) );
  NAND2_X1 U15483 ( .A1(n12351), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12391) );
  AOI22_X1 U15484 ( .A1(n12389), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12429), .ZN(n12390) );
  OAI211_X1 U15485 ( .C1(n12392), .C2(n12582), .A(n12391), .B(n12390), .ZN(
        n12400) );
  OAI22_X1 U15486 ( .A1(n19970), .A2(n12395), .B1(n12394), .B2(n12393), .ZN(
        n12399) );
  OAI22_X1 U15487 ( .A1(n12397), .A2(n12396), .B1(n10565), .B2(n12578), .ZN(
        n12398) );
  NOR4_X1 U15488 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n12398), .ZN(
        n16904) );
  INV_X1 U15489 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12402) );
  INV_X1 U15490 ( .A(n12607), .ZN(n12577) );
  OAI22_X1 U15491 ( .A1(n12558), .A2(n12402), .B1(n12577), .B2(n20403), .ZN(
        n12406) );
  INV_X1 U15492 ( .A(n12605), .ZN(n12579) );
  INV_X1 U15493 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12404) );
  INV_X1 U15494 ( .A(n12606), .ZN(n12581) );
  INV_X1 U15495 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12403) );
  OAI22_X1 U15496 ( .A1(n12579), .A2(n12404), .B1(n12581), .B2(n12403), .ZN(
        n12405) );
  NOR2_X1 U15497 ( .A1(n12406), .A2(n12405), .ZN(n12409) );
  XNOR2_X1 U15498 ( .A(n10416), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12609) );
  INV_X1 U15499 ( .A(n10221), .ZN(n12602) );
  AOI22_X1 U15500 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15501 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9611), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12407) );
  NAND4_X1 U15502 ( .A1(n12409), .A2(n12609), .A3(n12408), .A4(n12407), .ZN(
        n12420) );
  INV_X1 U15503 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12411) );
  INV_X1 U15504 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12410) );
  OAI22_X1 U15505 ( .A1(n12579), .A2(n12411), .B1(n12577), .B2(n12410), .ZN(
        n12415) );
  INV_X1 U15506 ( .A(n12601), .ZN(n12597) );
  OAI22_X1 U15507 ( .A1(n12597), .A2(n12413), .B1(n12581), .B2(n12412), .ZN(
        n12414) );
  NOR2_X1 U15508 ( .A1(n12415), .A2(n12414), .ZN(n12418) );
  AOI22_X1 U15509 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12602), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15510 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12416) );
  NAND4_X1 U15511 ( .A1(n12418), .A2(n12417), .A3(n12416), .A4(n12598), .ZN(
        n12419) );
  AND2_X1 U15512 ( .A1(n12420), .A2(n12419), .ZN(n12464) );
  NAND2_X1 U15513 ( .A1(n17047), .A2(n12464), .ZN(n12440) );
  AOI22_X1 U15514 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12202), .B1(
        n12421), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15515 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n12365), .ZN(n12427) );
  AOI22_X1 U15516 ( .A1(n12423), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10277), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15517 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12424), .B1(
        n12384), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12425) );
  NAND4_X1 U15518 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(
        n12439) );
  AOI22_X1 U15519 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12368), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15520 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12351), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12436) );
  INV_X1 U15521 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n20019) );
  NAND2_X1 U15522 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12429), .ZN(
        n12430) );
  OAI21_X1 U15523 ( .B1(n20019), .B2(n12431), .A(n12430), .ZN(n12432) );
  AOI21_X1 U15524 ( .B1(n12366), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n12432), .ZN(n12435) );
  NAND2_X1 U15525 ( .A1(n12433), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12434) );
  NAND4_X1 U15526 ( .A1(n12437), .A2(n12436), .A3(n12435), .A4(n12434), .ZN(
        n12438) );
  XNOR2_X1 U15527 ( .A(n12440), .B(n12461), .ZN(n12467) );
  NAND2_X1 U15528 ( .A1(n17076), .A2(n12464), .ZN(n15637) );
  OAI22_X1 U15529 ( .A1(n12558), .A2(n12442), .B1(n12581), .B2(n12441), .ZN(
        n12446) );
  OAI22_X1 U15530 ( .A1(n12579), .A2(n12444), .B1(n12577), .B2(n12443), .ZN(
        n12445) );
  NOR2_X1 U15531 ( .A1(n12446), .A2(n12445), .ZN(n12449) );
  AOI22_X1 U15532 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15533 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9611), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12447) );
  NAND4_X1 U15534 ( .A1(n12449), .A2(n12448), .A3(n12447), .A4(n12598), .ZN(
        n12460) );
  INV_X1 U15535 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12450) );
  OAI22_X1 U15536 ( .A1(n12558), .A2(n12451), .B1(n12581), .B2(n12450), .ZN(
        n12455) );
  INV_X1 U15537 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12453) );
  OAI22_X1 U15538 ( .A1(n12579), .A2(n12453), .B1(n12577), .B2(n12452), .ZN(
        n12454) );
  NOR2_X1 U15539 ( .A1(n12455), .A2(n12454), .ZN(n12458) );
  AOI22_X1 U15540 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12457) );
  AOI22_X1 U15541 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9611), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12456) );
  NAND4_X1 U15542 ( .A1(n12458), .A2(n12609), .A3(n12457), .A4(n12456), .ZN(
        n12459) );
  NAND2_X1 U15543 ( .A1(n12460), .A2(n12459), .ZN(n12468) );
  NAND2_X1 U15544 ( .A1(n12461), .A2(n12464), .ZN(n12469) );
  XOR2_X1 U15545 ( .A(n12468), .B(n12469), .Z(n12462) );
  NAND2_X1 U15546 ( .A1(n12462), .A2(n12514), .ZN(n15552) );
  INV_X1 U15547 ( .A(n12468), .ZN(n12463) );
  NAND2_X1 U15548 ( .A1(n17076), .A2(n12463), .ZN(n15554) );
  INV_X1 U15549 ( .A(n12464), .ZN(n12465) );
  NOR2_X1 U15550 ( .A1(n15554), .A2(n12465), .ZN(n12466) );
  NOR2_X1 U15551 ( .A1(n12469), .A2(n12468), .ZN(n12488) );
  OAI22_X1 U15552 ( .A1(n10221), .A2(n19945), .B1(n12597), .B2(n12338), .ZN(
        n12473) );
  INV_X1 U15553 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12471) );
  INV_X1 U15554 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12470) );
  OAI22_X1 U15555 ( .A1(n14489), .A2(n12471), .B1(n10239), .B2(n12470), .ZN(
        n12472) );
  NOR2_X1 U15556 ( .A1(n12473), .A2(n12472), .ZN(n12476) );
  AOI22_X1 U15557 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15558 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12474) );
  NAND4_X1 U15559 ( .A1(n12476), .A2(n12475), .A3(n12474), .A4(n12598), .ZN(
        n12487) );
  INV_X1 U15560 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12478) );
  OAI22_X1 U15561 ( .A1(n12558), .A2(n12478), .B1(n12597), .B2(n12477), .ZN(
        n12482) );
  INV_X1 U15562 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12480) );
  OAI22_X1 U15563 ( .A1(n14489), .A2(n12480), .B1(n10239), .B2(n12479), .ZN(
        n12481) );
  NOR2_X1 U15564 ( .A1(n12482), .A2(n12481), .ZN(n12485) );
  AOI22_X1 U15565 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15566 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12483) );
  NAND4_X1 U15567 ( .A1(n12485), .A2(n12609), .A3(n12484), .A4(n12483), .ZN(
        n12486) );
  AND2_X1 U15568 ( .A1(n12487), .A2(n12486), .ZN(n12490) );
  NAND2_X1 U15569 ( .A1(n12488), .A2(n12490), .ZN(n12542) );
  OAI211_X1 U15570 ( .C1(n12488), .C2(n12490), .A(n12514), .B(n12542), .ZN(
        n12492) );
  INV_X1 U15571 ( .A(n12492), .ZN(n12489) );
  INV_X1 U15572 ( .A(n12490), .ZN(n12491) );
  NOR2_X1 U15573 ( .A1(n17047), .A2(n12491), .ZN(n15545) );
  INV_X1 U15574 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12496) );
  OAI22_X1 U15575 ( .A1(n12558), .A2(n12496), .B1(n12581), .B2(n12495), .ZN(
        n12500) );
  INV_X1 U15576 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12498) );
  INV_X1 U15577 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12497) );
  OAI22_X1 U15578 ( .A1(n12579), .A2(n12498), .B1(n12577), .B2(n12497), .ZN(
        n12499) );
  NOR2_X1 U15579 ( .A1(n12500), .A2(n12499), .ZN(n12503) );
  AOI22_X1 U15580 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15581 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12501) );
  NAND4_X1 U15582 ( .A1(n12503), .A2(n12502), .A3(n12501), .A4(n12598), .ZN(
        n12513) );
  OAI22_X1 U15583 ( .A1(n12558), .A2(n12505), .B1(n12581), .B2(n12504), .ZN(
        n12508) );
  INV_X1 U15584 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12506) );
  OAI22_X1 U15585 ( .A1(n12579), .A2(n12506), .B1(n12577), .B2(n20410), .ZN(
        n12507) );
  NOR2_X1 U15586 ( .A1(n12508), .A2(n12507), .ZN(n12511) );
  AOI22_X1 U15587 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U15588 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9611), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12509) );
  NAND4_X1 U15589 ( .A1(n12511), .A2(n12609), .A3(n12510), .A4(n12509), .ZN(
        n12512) );
  AND2_X1 U15590 ( .A1(n12513), .A2(n12512), .ZN(n12516) );
  XNOR2_X1 U15591 ( .A(n12542), .B(n12516), .ZN(n12515) );
  NAND2_X1 U15592 ( .A1(n12515), .A2(n12514), .ZN(n12518) );
  INV_X1 U15593 ( .A(n12516), .ZN(n12541) );
  NOR2_X1 U15594 ( .A1(n17047), .A2(n12541), .ZN(n15537) );
  INV_X1 U15595 ( .A(n12518), .ZN(n12519) );
  INV_X1 U15596 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12521) );
  OAI22_X1 U15597 ( .A1(n12558), .A2(n12522), .B1(n12577), .B2(n12521), .ZN(
        n12526) );
  INV_X1 U15598 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12524) );
  INV_X1 U15599 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12523) );
  OAI22_X1 U15600 ( .A1(n12579), .A2(n12524), .B1(n12581), .B2(n12523), .ZN(
        n12525) );
  NOR2_X1 U15601 ( .A1(n12526), .A2(n12525), .ZN(n12529) );
  AOI22_X1 U15602 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U15603 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12527) );
  NAND4_X1 U15604 ( .A1(n12529), .A2(n12528), .A3(n12527), .A4(n12598), .ZN(
        n12540) );
  INV_X1 U15605 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12530) );
  OAI22_X1 U15606 ( .A1(n12558), .A2(n12531), .B1(n12577), .B2(n12530), .ZN(
        n12535) );
  INV_X1 U15607 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12532) );
  OAI22_X1 U15608 ( .A1(n12579), .A2(n12533), .B1(n12581), .B2(n12532), .ZN(
        n12534) );
  NOR2_X1 U15609 ( .A1(n12535), .A2(n12534), .ZN(n12538) );
  AOI22_X1 U15610 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15611 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9611), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12536) );
  NAND4_X1 U15612 ( .A1(n12538), .A2(n12609), .A3(n12537), .A4(n12536), .ZN(
        n12539) );
  NAND2_X1 U15613 ( .A1(n12540), .A2(n12539), .ZN(n12546) );
  OR2_X1 U15614 ( .A1(n12542), .A2(n12541), .ZN(n12544) );
  NOR2_X1 U15615 ( .A1(n12544), .A2(n12546), .ZN(n15525) );
  AOI211_X1 U15616 ( .C1(n12546), .C2(n12544), .A(n12543), .B(n15525), .ZN(
        n12545) );
  NOR2_X1 U15617 ( .A1(n17047), .A2(n12546), .ZN(n15532) );
  INV_X1 U15618 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12548) );
  OAI22_X1 U15619 ( .A1(n12558), .A2(n12548), .B1(n12581), .B2(n12547), .ZN(
        n12552) );
  OAI22_X1 U15620 ( .A1(n12579), .A2(n12550), .B1(n12577), .B2(n12549), .ZN(
        n12551) );
  NOR2_X1 U15621 ( .A1(n12552), .A2(n12551), .ZN(n12555) );
  AOI22_X1 U15622 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15623 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12553) );
  NAND4_X1 U15624 ( .A1(n12555), .A2(n12554), .A3(n12553), .A4(n12598), .ZN(
        n12567) );
  OAI22_X1 U15625 ( .A1(n12558), .A2(n12557), .B1(n12581), .B2(n12556), .ZN(
        n12562) );
  OAI22_X1 U15626 ( .A1(n12579), .A2(n12560), .B1(n12577), .B2(n12559), .ZN(
        n12561) );
  NOR2_X1 U15627 ( .A1(n12562), .A2(n12561), .ZN(n12565) );
  AOI22_X1 U15628 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15629 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9611), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12563) );
  NAND4_X1 U15630 ( .A1(n12565), .A2(n12609), .A3(n12564), .A4(n12563), .ZN(
        n12566) );
  NAND2_X1 U15631 ( .A1(n12567), .A2(n12566), .ZN(n12590) );
  INV_X1 U15632 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12568) );
  OAI22_X1 U15633 ( .A1(n10221), .A2(n19970), .B1(n12577), .B2(n12568), .ZN(
        n12572) );
  OAI22_X1 U15634 ( .A1(n12579), .A2(n12570), .B1(n12581), .B2(n12569), .ZN(
        n12571) );
  NOR2_X1 U15635 ( .A1(n12572), .A2(n12571), .ZN(n12575) );
  AOI22_X1 U15636 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U15637 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12573) );
  NAND4_X1 U15638 ( .A1(n12575), .A2(n12574), .A3(n12573), .A4(n12598), .ZN(
        n12589) );
  OAI22_X1 U15639 ( .A1(n12579), .A2(n12578), .B1(n12577), .B2(n12576), .ZN(
        n12584) );
  OAI22_X1 U15640 ( .A1(n12597), .A2(n12582), .B1(n12581), .B2(n12580), .ZN(
        n12583) );
  NOR2_X1 U15641 ( .A1(n12584), .A2(n12583), .ZN(n12587) );
  AOI22_X1 U15642 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12602), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15643 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9611), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12585) );
  NAND4_X1 U15644 ( .A1(n12587), .A2(n12586), .A3(n12609), .A4(n12585), .ZN(
        n12588) );
  NAND2_X1 U15645 ( .A1(n12589), .A2(n12588), .ZN(n12593) );
  INV_X1 U15646 ( .A(n12590), .ZN(n15527) );
  AND2_X1 U15647 ( .A1(n17047), .A2(n15527), .ZN(n12591) );
  NAND2_X1 U15648 ( .A1(n15525), .A2(n12591), .ZN(n12592) );
  NOR2_X1 U15649 ( .A1(n12592), .A2(n12593), .ZN(n12594) );
  AOI21_X1 U15650 ( .B1(n12593), .B2(n12592), .A(n12594), .ZN(n15520) );
  AOI22_X1 U15651 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12596) );
  NAND2_X1 U15652 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12595) );
  OAI211_X1 U15653 ( .C1(n20019), .C2(n12597), .A(n12596), .B(n12595), .ZN(
        n12614) );
  AOI22_X1 U15654 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U15655 ( .A1(n12605), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12607), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12599) );
  NAND3_X1 U15656 ( .A1(n12600), .A2(n12599), .A3(n12598), .ZN(n12613) );
  INV_X1 U15657 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n20486) );
  AOI22_X1 U15658 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12601), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12604) );
  NAND2_X1 U15659 ( .A1(n10419), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12603) );
  OAI211_X1 U15660 ( .C1(n10239), .C2(n20486), .A(n12604), .B(n12603), .ZN(
        n12612) );
  AOI22_X1 U15661 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U15662 ( .A1(n12607), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12606), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12608) );
  NAND3_X1 U15663 ( .A1(n12610), .A2(n12609), .A3(n12608), .ZN(n12611) );
  OAI22_X1 U15664 ( .A1(n12614), .A2(n12613), .B1(n12612), .B2(n12611), .ZN(
        n12615) );
  INV_X1 U15665 ( .A(n16237), .ZN(n12748) );
  OAI21_X1 U15666 ( .B1(n12618), .B2(n12748), .A(n12617), .ZN(n13733) );
  NAND2_X1 U15667 ( .A1(n17076), .A2(n19952), .ZN(n12628) );
  NAND2_X1 U15668 ( .A1(n12628), .A2(n10451), .ZN(n12619) );
  NAND2_X1 U15669 ( .A1(n12619), .A2(n16237), .ZN(n12620) );
  NAND2_X1 U15670 ( .A1(n12620), .A2(n10444), .ZN(n12621) );
  AND4_X1 U15671 ( .A1(n13733), .A2(n13738), .A3(n12622), .A4(n12621), .ZN(
        n12627) );
  NAND2_X1 U15672 ( .A1(n12624), .A2(n10444), .ZN(n12625) );
  NAND2_X1 U15673 ( .A1(n12623), .A2(n12625), .ZN(n12626) );
  INV_X1 U15674 ( .A(n12628), .ZN(n12629) );
  NAND2_X1 U15675 ( .A1(n12866), .A2(n12629), .ZN(n14487) );
  INV_X1 U15676 ( .A(n12630), .ZN(n17049) );
  NAND2_X1 U15677 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n17069) );
  AND2_X1 U15678 ( .A1(n12861), .A2(n17069), .ZN(n12858) );
  NAND2_X1 U15679 ( .A1(n17049), .A2(n12858), .ZN(n12631) );
  OAI22_X1 U15680 ( .A1(n17055), .A2(n14487), .B1(n12631), .B2(n17050), .ZN(
        n12871) );
  NOR2_X1 U15681 ( .A1(n12632), .A2(n13738), .ZN(n12633) );
  AND2_X1 U15682 ( .A1(n12634), .A2(n12633), .ZN(n13734) );
  INV_X1 U15683 ( .A(n12656), .ZN(n12645) );
  NAND2_X1 U15684 ( .A1(n12774), .A2(n19848), .ZN(n12769) );
  NAND2_X1 U15685 ( .A1(n12636), .A2(n21204), .ZN(n12651) );
  INV_X1 U15686 ( .A(n12651), .ZN(n12742) );
  NOR2_X1 U15687 ( .A1(n16237), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12639) );
  INV_X1 U15688 ( .A(n12639), .ZN(n12740) );
  INV_X1 U15689 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12637) );
  INV_X1 U15690 ( .A(n12652), .ZN(n12739) );
  INV_X1 U15691 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15941) );
  OAI22_X1 U15692 ( .A1(n12740), .A2(n12637), .B1(n12739), .B2(n15941), .ZN(
        n12638) );
  AOI21_X1 U15693 ( .B1(n12742), .B2(P2_REIP_REG_30__SCAN_IN), .A(n12638), 
        .ZN(n12747) );
  INV_X1 U15694 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20534) );
  OR2_X1 U15695 ( .A1(n14464), .A2(n20534), .ZN(n12641) );
  AOI22_X1 U15696 ( .A1(n14461), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12640) );
  NAND2_X1 U15697 ( .A1(n12641), .A2(n12640), .ZN(n14099) );
  NOR2_X1 U15698 ( .A1(n10443), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12643) );
  INV_X1 U15699 ( .A(n12719), .ZN(n12688) );
  NAND2_X1 U15700 ( .A1(n12645), .A2(n12652), .ZN(n12663) );
  MUX2_X1 U15701 ( .A(n16237), .B(n20615), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12646) );
  AND2_X1 U15702 ( .A1(n12663), .A2(n12646), .ZN(n12647) );
  INV_X1 U15703 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12957) );
  NAND2_X1 U15704 ( .A1(n17047), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12648) );
  OAI211_X1 U15705 ( .C1(n16237), .C2(n12957), .A(n12648), .B(n21204), .ZN(
        n12649) );
  INV_X1 U15706 ( .A(n12649), .ZN(n12650) );
  OR2_X1 U15707 ( .A1(n12651), .A2(n14081), .ZN(n12654) );
  AOI22_X1 U15708 ( .A1(n12639), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12652), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12653) );
  NAND2_X1 U15709 ( .A1(n12654), .A2(n12653), .ZN(n12660) );
  INV_X1 U15710 ( .A(n12655), .ZN(n12659) );
  NAND2_X1 U15711 ( .A1(n12656), .A2(n16237), .ZN(n12657) );
  MUX2_X1 U15712 ( .A(n12657), .B(n20605), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12658) );
  OAI21_X1 U15713 ( .B1(n12659), .B2(n12719), .A(n12658), .ZN(n13371) );
  NOR2_X1 U15714 ( .A1(n13372), .A2(n13371), .ZN(n12662) );
  NOR2_X1 U15715 ( .A1(n13011), .A2(n12660), .ZN(n12661) );
  NOR2_X2 U15716 ( .A1(n12662), .A2(n12661), .ZN(n12667) );
  NAND2_X1 U15717 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12664) );
  OAI211_X1 U15718 ( .C1(n12719), .C2(n12665), .A(n12664), .B(n12663), .ZN(
        n12666) );
  XNOR2_X1 U15719 ( .A(n12667), .B(n12666), .ZN(n13370) );
  INV_X1 U15720 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19896) );
  INV_X1 U15721 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20519) );
  OAI222_X1 U15722 ( .A1(n12739), .A2(n19925), .B1(n12740), .B2(n19896), .C1(
        n12651), .C2(n20519), .ZN(n13369) );
  NOR2_X1 U15723 ( .A1(n13370), .A2(n13369), .ZN(n13368) );
  NOR2_X1 U15724 ( .A1(n12667), .A2(n12666), .ZN(n12668) );
  NOR2_X2 U15725 ( .A1(n13368), .A2(n12668), .ZN(n13744) );
  AOI22_X1 U15726 ( .A1(n12652), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12670) );
  NAND2_X1 U15727 ( .A1(n14461), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12669) );
  OAI211_X1 U15728 ( .C1(n12719), .C2(n12671), .A(n12670), .B(n12669), .ZN(
        n12672) );
  INV_X1 U15729 ( .A(n12672), .ZN(n12675) );
  INV_X1 U15730 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n12673) );
  OR2_X1 U15731 ( .A1(n12651), .A2(n12673), .ZN(n12674) );
  NAND2_X1 U15732 ( .A1(n12675), .A2(n12674), .ZN(n13743) );
  OR2_X1 U15733 ( .A1(n12651), .A2(n14003), .ZN(n12681) );
  INV_X1 U15734 ( .A(n12676), .ZN(n12677) );
  OR2_X1 U15735 ( .A1(n12719), .A2(n12677), .ZN(n12679) );
  AOI22_X1 U15736 ( .A1(n14461), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12652), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12678) );
  AND2_X1 U15737 ( .A1(n12679), .A2(n12678), .ZN(n12680) );
  AOI22_X1 U15738 ( .A1(n12742), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n14461), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12685) );
  OAI22_X1 U15739 ( .A1(n12719), .A2(n12682), .B1(n12739), .B2(n14023), .ZN(
        n12683) );
  INV_X1 U15740 ( .A(n12683), .ZN(n12684) );
  NAND2_X1 U15741 ( .A1(n12685), .A2(n12684), .ZN(n14021) );
  AOI21_X1 U15742 ( .B1(n12688), .B2(n12687), .A(n12686), .ZN(n16194) );
  AOI222_X1 U15743 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n12742), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(P2_EAX_REG_6__SCAN_IN), 
        .C2(n14461), .ZN(n16193) );
  OAI22_X2 U15744 ( .A1(n16194), .A2(n16193), .B1(n10362), .B2(n12719), .ZN(
        n16179) );
  INV_X1 U15745 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19885) );
  OAI222_X1 U15746 ( .A1(n12739), .A2(n10835), .B1(n12740), .B2(n19885), .C1(
        n14464), .C2(n10865), .ZN(n16178) );
  OR2_X1 U15747 ( .A1(n14464), .A2(n12689), .ZN(n12694) );
  INV_X1 U15748 ( .A(n12690), .ZN(n19789) );
  OR2_X1 U15749 ( .A1(n12719), .A2(n19789), .ZN(n12692) );
  AOI22_X1 U15750 ( .A1(n14461), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12652), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12691) );
  AND2_X1 U15751 ( .A1(n12692), .A2(n12691), .ZN(n12693) );
  NAND2_X1 U15752 ( .A1(n12742), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U15753 ( .A1(n14461), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12652), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12695) );
  OAI211_X1 U15754 ( .C1(n13364), .C2(n12719), .A(n12696), .B(n12695), .ZN(
        n16164) );
  OR2_X1 U15755 ( .A1(n14464), .A2(n15879), .ZN(n12700) );
  INV_X1 U15756 ( .A(n19778), .ZN(n13561) );
  OR2_X1 U15757 ( .A1(n12719), .A2(n13561), .ZN(n12698) );
  AOI22_X1 U15758 ( .A1(n14461), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12697) );
  AND2_X1 U15759 ( .A1(n12698), .A2(n12697), .ZN(n12699) );
  INV_X1 U15760 ( .A(n12701), .ZN(n13560) );
  OR2_X1 U15761 ( .A1(n14464), .A2(n12702), .ZN(n12704) );
  AOI22_X1 U15762 ( .A1(n14461), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12703) );
  OAI211_X1 U15763 ( .C1(n13560), .C2(n12719), .A(n12704), .B(n12703), .ZN(
        n14038) );
  OR2_X1 U15764 ( .A1(n12651), .A2(n12705), .ZN(n12709) );
  INV_X1 U15765 ( .A(n13847), .ZN(n19773) );
  OR2_X1 U15766 ( .A1(n12719), .A2(n19773), .ZN(n12707) );
  AOI22_X1 U15767 ( .A1(n14461), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12706) );
  AND2_X1 U15768 ( .A1(n12707), .A2(n12706), .ZN(n12708) );
  INV_X1 U15769 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n12710) );
  OR2_X1 U15770 ( .A1(n14464), .A2(n12710), .ZN(n12712) );
  AOI22_X1 U15771 ( .A1(n14461), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12711) );
  OAI211_X1 U15772 ( .C1(n13848), .C2(n12719), .A(n12712), .B(n12711), .ZN(
        n12846) );
  OR2_X1 U15773 ( .A1(n14464), .A2(n15842), .ZN(n12716) );
  OR2_X1 U15774 ( .A1(n12719), .A2(n19769), .ZN(n12714) );
  AOI22_X1 U15775 ( .A1(n14461), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12713) );
  AND2_X1 U15776 ( .A1(n12714), .A2(n12713), .ZN(n12715) );
  NAND2_X1 U15777 ( .A1(n12742), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15778 ( .A1(n14461), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12717) );
  OAI211_X1 U15779 ( .C1(n15588), .C2(n12719), .A(n12718), .B(n12717), .ZN(
        n16964) );
  OR2_X1 U15780 ( .A1(n14464), .A2(n12720), .ZN(n12722) );
  AOI22_X1 U15781 ( .A1(n14461), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12721) );
  INV_X1 U15782 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15792) );
  OR2_X1 U15783 ( .A1(n12651), .A2(n15792), .ZN(n12724) );
  AOI22_X1 U15784 ( .A1(n14461), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12723) );
  INV_X1 U15785 ( .A(n12725), .ZN(n15651) );
  INV_X1 U15786 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20537) );
  OR2_X1 U15787 ( .A1(n14464), .A2(n20537), .ZN(n12727) );
  AOI22_X1 U15788 ( .A1(n14461), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12726) );
  OR2_X1 U15789 ( .A1(n14464), .A2(n15768), .ZN(n12729) );
  AOI22_X1 U15790 ( .A1(n14461), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12728) );
  NAND2_X1 U15791 ( .A1(n12729), .A2(n12728), .ZN(n15437) );
  INV_X1 U15792 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20540) );
  OR2_X1 U15793 ( .A1(n14464), .A2(n20540), .ZN(n12731) );
  AOI22_X1 U15794 ( .A1(n14461), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12730) );
  NAND2_X1 U15795 ( .A1(n12731), .A2(n12730), .ZN(n15422) );
  INV_X1 U15796 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n15733) );
  OR2_X1 U15797 ( .A1(n14464), .A2(n15733), .ZN(n12733) );
  AOI22_X1 U15798 ( .A1(n14461), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12732) );
  NAND2_X1 U15799 ( .A1(n12733), .A2(n12732), .ZN(n16040) );
  INV_X1 U15800 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15639) );
  OAI22_X1 U15801 ( .A1(n12740), .A2(n15639), .B1(n12739), .B2(n16028), .ZN(
        n12734) );
  AOI21_X1 U15802 ( .B1(n12742), .B2(P2_REIP_REG_23__SCAN_IN), .A(n12734), 
        .ZN(n15407) );
  INV_X1 U15803 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15631) );
  OAI22_X1 U15804 ( .A1(n12740), .A2(n15631), .B1(n12739), .B2(n21106), .ZN(
        n12735) );
  AOI21_X1 U15805 ( .B1(n12742), .B2(P2_REIP_REG_24__SCAN_IN), .A(n12735), 
        .ZN(n15627) );
  INV_X1 U15806 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20546) );
  OR2_X1 U15807 ( .A1(n14464), .A2(n20546), .ZN(n12737) );
  AOI22_X1 U15808 ( .A1(n12639), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12736) );
  NAND2_X1 U15809 ( .A1(n12737), .A2(n12736), .ZN(n15618) );
  INV_X1 U15810 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n15612) );
  OAI22_X1 U15811 ( .A1(n12740), .A2(n15612), .B1(n12739), .B2(n15999), .ZN(
        n12738) );
  AOI21_X1 U15812 ( .B1(n12742), .B2(P2_REIP_REG_26__SCAN_IN), .A(n12738), 
        .ZN(n15609) );
  INV_X1 U15813 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15603) );
  OAI22_X1 U15814 ( .A1(n12740), .A2(n15603), .B1(n12739), .B2(n15970), .ZN(
        n12741) );
  AOI21_X1 U15815 ( .B1(n12742), .B2(P2_REIP_REG_27__SCAN_IN), .A(n12741), 
        .ZN(n15392) );
  INV_X1 U15816 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20552) );
  OR2_X1 U15817 ( .A1(n14464), .A2(n20552), .ZN(n12744) );
  AOI22_X1 U15818 ( .A1(n12639), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12743) );
  NAND2_X1 U15819 ( .A1(n12744), .A2(n12743), .ZN(n15380) );
  OR2_X1 U15820 ( .A1(n14464), .A2(n20554), .ZN(n12746) );
  AOI22_X1 U15821 ( .A1(n12639), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12745) );
  NAND2_X1 U15822 ( .A1(n12746), .A2(n12745), .ZN(n15363) );
  NOR2_X2 U15823 ( .A1(n15365), .A2(n12747), .ZN(n14466) );
  AOI21_X1 U15824 ( .B1(n12747), .B2(n15365), .A(n14466), .ZN(n15938) );
  NAND2_X1 U15825 ( .A1(n15938), .A2(n19859), .ZN(n12767) );
  NOR2_X1 U15826 ( .A1(n12748), .A2(n19962), .ZN(n12749) );
  NAND2_X1 U15827 ( .A1(n19834), .A2(n12749), .ZN(n13007) );
  NOR4_X1 U15828 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12753) );
  NOR4_X1 U15829 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12752) );
  NOR4_X1 U15830 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12751) );
  NOR4_X1 U15831 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12750) );
  NAND4_X1 U15832 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n12758) );
  NOR4_X1 U15833 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12756) );
  NOR4_X1 U15834 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12755) );
  NOR4_X1 U15835 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n12754) );
  INV_X1 U15836 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20521) );
  NAND4_X1 U15837 ( .A1(n12756), .A2(n12755), .A3(n12754), .A4(n20521), .ZN(
        n12757) );
  NOR2_X2 U15838 ( .A1(n13007), .A2(n13860), .ZN(n19804) );
  NOR2_X2 U15839 ( .A1(n13007), .A2(n13858), .ZN(n19803) );
  AOI22_X1 U15840 ( .A1(n19804), .A2(BUF2_REG_30__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12760) );
  INV_X1 U15841 ( .A(n12761), .ZN(n12762) );
  MUX2_X1 U15842 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n13858), .Z(n19813) );
  AOI22_X1 U15843 ( .A1(n19802), .A2(n19813), .B1(n19858), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n12763) );
  INV_X1 U15844 ( .A(n12763), .ZN(n12764) );
  NOR2_X1 U15845 ( .A1(n12765), .A2(n12764), .ZN(n12766) );
  NAND2_X1 U15846 ( .A1(n12769), .A2(n12768), .ZN(P2_U2889) );
  AND2_X1 U15847 ( .A1(n12770), .A2(n12771), .ZN(n13746) );
  NAND2_X1 U15848 ( .A1(n17055), .A2(n13746), .ZN(n12869) );
  NAND2_X1 U15849 ( .A1(n12869), .A2(n12772), .ZN(n12773) );
  NAND2_X1 U15850 ( .A1(n12774), .A2(n19793), .ZN(n12782) );
  INV_X1 U15851 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n15352) );
  AOI22_X1 U15852 ( .A1(n10882), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12775) );
  OAI21_X1 U15853 ( .B1(n9591), .B2(n15352), .A(n12775), .ZN(n12777) );
  AOI21_X1 U15854 ( .B1(n12778), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12777), .ZN(n14420) );
  NAND2_X1 U15855 ( .A1(n19796), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12779) );
  INV_X1 U15856 ( .A(n12780), .ZN(n12781) );
  NAND2_X1 U15857 ( .A1(n12782), .A2(n12781), .ZN(P2_U2857) );
  NOR2_X1 U15858 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12784) );
  NOR4_X1 U15859 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12783) );
  NAND4_X1 U15860 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12784), .A4(n12783), .ZN(n12797) );
  NOR4_X1 U15861 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12788) );
  NOR4_X1 U15862 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12787) );
  NOR4_X1 U15863 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12786) );
  NOR4_X1 U15864 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12785) );
  AND4_X1 U15865 ( .A1(n12788), .A2(n12787), .A3(n12786), .A4(n12785), .ZN(
        n12793) );
  NOR4_X1 U15866 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n12791) );
  NOR4_X1 U15867 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12790) );
  NOR4_X1 U15868 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12789) );
  INV_X1 U15869 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20985) );
  AND4_X1 U15870 ( .A1(n12791), .A2(n12790), .A3(n12789), .A4(n20985), .ZN(
        n12792) );
  NAND2_X1 U15871 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  INV_X1 U15872 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21047) );
  NOR3_X1 U15873 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21047), .ZN(n12796) );
  NOR4_X1 U15874 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12795) );
  NAND4_X1 U15875 ( .A1(n14738), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12796), .A4(
        n12795), .ZN(U214) );
  NOR2_X1 U15876 ( .A1(n13858), .A2(n12797), .ZN(n17168) );
  NAND2_X1 U15877 ( .A1(n17168), .A2(U214), .ZN(U212) );
  OR2_X1 U15878 ( .A1(n12823), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12799) );
  NAND2_X1 U15879 ( .A1(n12798), .A2(n12799), .ZN(n15857) );
  INV_X1 U15880 ( .A(n15857), .ZN(n12833) );
  INV_X1 U15881 ( .A(n12804), .ZN(n12802) );
  INV_X1 U15882 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12800) );
  NAND2_X1 U15883 ( .A1(n14076), .A2(n12800), .ZN(n12801) );
  NAND2_X1 U15884 ( .A1(n12802), .A2(n12801), .ZN(n14132) );
  INV_X1 U15885 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15514) );
  AOI22_X1 U15886 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12803), .B1(n15514), 
        .B2(n19598), .ZN(n15518) );
  AOI22_X1 U15887 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14480), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19598), .ZN(n14073) );
  NOR2_X1 U15888 ( .A1(n15518), .A2(n14073), .ZN(n14127) );
  AND2_X1 U15889 ( .A1(n14132), .A2(n14127), .ZN(n14114) );
  OAI21_X1 U15890 ( .B1(n12804), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n12805), .ZN(n14120) );
  AND2_X1 U15891 ( .A1(n14114), .A2(n14120), .ZN(n19751) );
  AND2_X1 U15892 ( .A1(n12805), .A2(n14004), .ZN(n12806) );
  OR2_X1 U15893 ( .A1(n12806), .A2(n12807), .ZN(n19752) );
  NAND2_X1 U15894 ( .A1(n19751), .A2(n19752), .ZN(n19756) );
  OR2_X1 U15895 ( .A1(n12807), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12808) );
  AND2_X1 U15896 ( .A1(n12810), .A2(n12808), .ZN(n19720) );
  NOR2_X1 U15897 ( .A1(n19756), .A2(n19720), .ZN(n19707) );
  NAND2_X1 U15898 ( .A1(n12810), .A2(n12809), .ZN(n12811) );
  NAND2_X1 U15899 ( .A1(n12812), .A2(n12811), .ZN(n19709) );
  AND2_X1 U15900 ( .A1(n19707), .A2(n19709), .ZN(n19710) );
  AND2_X1 U15901 ( .A1(n12812), .A2(n15909), .ZN(n12813) );
  OR2_X1 U15902 ( .A1(n12813), .A2(n12814), .ZN(n19697) );
  AND2_X1 U15903 ( .A1(n19710), .A2(n19697), .ZN(n19698) );
  NOR2_X1 U15904 ( .A1(n12814), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12815) );
  OR2_X1 U15905 ( .A1(n12816), .A2(n12815), .ZN(n15902) );
  NAND2_X1 U15906 ( .A1(n19698), .A2(n15902), .ZN(n19688) );
  OR2_X1 U15907 ( .A1(n12816), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12817) );
  AND2_X1 U15908 ( .A1(n12818), .A2(n12817), .ZN(n19689) );
  NOR2_X1 U15909 ( .A1(n19688), .A2(n19689), .ZN(n19670) );
  NAND2_X1 U15910 ( .A1(n12818), .A2(n15880), .ZN(n12819) );
  NAND2_X1 U15911 ( .A1(n12820), .A2(n12819), .ZN(n19672) );
  AND2_X1 U15912 ( .A1(n19670), .A2(n19672), .ZN(n19673) );
  NAND2_X1 U15913 ( .A1(n12820), .A2(n16941), .ZN(n12821) );
  NAND2_X1 U15914 ( .A1(n12822), .A2(n12821), .ZN(n14036) );
  AND2_X1 U15915 ( .A1(n19673), .A2(n14036), .ZN(n14035) );
  AND2_X1 U15916 ( .A1(n12822), .A2(n15865), .ZN(n12824) );
  OR2_X1 U15917 ( .A1(n12824), .A2(n12823), .ZN(n15491) );
  AND2_X1 U15918 ( .A1(n14035), .A2(n15491), .ZN(n12831) );
  INV_X1 U15919 ( .A(n12831), .ZN(n12832) );
  INV_X1 U15920 ( .A(n14430), .ZN(n12827) );
  NAND2_X1 U15921 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12826) );
  INV_X1 U15922 ( .A(n12828), .ZN(n12830) );
  NAND2_X1 U15923 ( .A1(n12830), .A2(n12829), .ZN(n19730) );
  INV_X1 U15924 ( .A(n19730), .ZN(n19757) );
  NAND2_X1 U15925 ( .A1(n12831), .A2(n15857), .ZN(n15479) );
  NAND2_X1 U15926 ( .A1(n15517), .A2(n15479), .ZN(n15490) );
  AOI21_X1 U15927 ( .B1(n12833), .B2(n12832), .A(n15490), .ZN(n12854) );
  INV_X1 U15928 ( .A(n17073), .ZN(n12859) );
  NAND2_X1 U15929 ( .A1(n17069), .A2(n21109), .ZN(n12849) );
  NAND2_X1 U15930 ( .A1(n12849), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12834) );
  NOR2_X1 U15931 ( .A1(n13721), .A2(n12834), .ZN(n12835) );
  NOR2_X1 U15932 ( .A1(n21204), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20489) );
  INV_X1 U15933 ( .A(n20489), .ZN(n12836) );
  NOR2_X1 U15934 ( .A1(n20494), .A2(n12836), .ZN(n17071) );
  NAND2_X1 U15935 ( .A1(n19736), .A2(n19730), .ZN(n12837) );
  OR2_X1 U15936 ( .A1(n17071), .A2(n12837), .ZN(n12838) );
  NAND2_X1 U15937 ( .A1(n19737), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19654) );
  AOI22_X1 U15938 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19732), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19652), .ZN(n12839) );
  OAI211_X1 U15939 ( .C1(n12840), .C2(n19684), .A(n12839), .B(n19736), .ZN(
        n12853) );
  NOR2_X1 U15940 ( .A1(n12881), .A2(n12841), .ZN(n12855) );
  INV_X1 U15941 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19595) );
  NOR2_X1 U15942 ( .A1(n19595), .A2(n20517), .ZN(n20510) );
  NOR2_X1 U15943 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20498) );
  NOR3_X1 U15944 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20510), .A3(n20498), 
        .ZN(n20503) );
  AND2_X1 U15945 ( .A1(n20503), .A2(n17069), .ZN(n13706) );
  AND2_X1 U15946 ( .A1(n13706), .A2(n21109), .ZN(n17075) );
  INV_X1 U15947 ( .A(n17075), .ZN(n12842) );
  NAND2_X1 U15948 ( .A1(n15341), .A2(n12842), .ZN(n12844) );
  INV_X1 U15949 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16898) );
  NAND3_X1 U15950 ( .A1(n12855), .A2(n16898), .A3(n12849), .ZN(n12843) );
  OAI22_X1 U15951 ( .A1(n19665), .A2(n15857), .B1(n19683), .B2(n10884), .ZN(
        n12852) );
  OR2_X1 U15952 ( .A1(n12846), .A2(n12845), .ZN(n12847) );
  NAND2_X1 U15953 ( .A1(n12847), .A2(n15480), .ZN(n19817) );
  AOI21_X1 U15954 ( .B1(n12848), .B2(n15495), .A(n9685), .ZN(n13851) );
  INV_X1 U15955 ( .A(n13851), .ZN(n16125) );
  NOR2_X1 U15956 ( .A1(n13721), .A2(n12849), .ZN(n12850) );
  OAI22_X1 U15957 ( .A1(n19817), .A2(n19726), .B1(n16125), .B2(n19748), .ZN(
        n12851) );
  OR4_X1 U15958 ( .A1(n12854), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        P2_U2842) );
  NOR2_X1 U15959 ( .A1(n12881), .A2(n12623), .ZN(n15511) );
  INV_X1 U15960 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12857) );
  INV_X1 U15961 ( .A(n12855), .ZN(n12856) );
  NAND2_X1 U15962 ( .A1(n20585), .A2(n20495), .ZN(n19597) );
  OAI211_X1 U15963 ( .C1(n15511), .C2(n12857), .A(n12856), .B(n19597), .ZN(
        P2_U2814) );
  NOR4_X1 U15964 ( .A1(n17050), .A2(n12630), .A3(n12858), .A4(n13706), .ZN(
        n17058) );
  NOR2_X1 U15965 ( .A1(n17058), .A2(n12859), .ZN(n20625) );
  OAI21_X1 U15966 ( .B1(n20625), .B2(n12874), .A(n12860), .ZN(P2_U2819) );
  INV_X1 U15967 ( .A(n12861), .ZN(n15299) );
  INV_X1 U15968 ( .A(n19599), .ZN(n12864) );
  INV_X1 U15969 ( .A(n19597), .ZN(n12862) );
  OAI21_X1 U15970 ( .B1(n12862), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n12864), 
        .ZN(n12863) );
  OAI21_X1 U15971 ( .B1(n15299), .B2(n12864), .A(n12863), .ZN(P2_U3612) );
  NAND2_X1 U15972 ( .A1(n10442), .A2(n13706), .ZN(n12865) );
  OR2_X1 U15973 ( .A1(n17050), .A2(n12865), .ZN(n12867) );
  NAND2_X1 U15974 ( .A1(n12867), .A2(n12866), .ZN(n13711) );
  INV_X1 U15975 ( .A(n13711), .ZN(n12868) );
  NAND2_X1 U15976 ( .A1(n12869), .A2(n12868), .ZN(n12870) );
  NOR2_X1 U15977 ( .A1(n12871), .A2(n12870), .ZN(n12873) );
  INV_X1 U15978 ( .A(n12623), .ZN(n12973) );
  NAND3_X1 U15979 ( .A1(n13707), .A2(n12973), .A3(n13706), .ZN(n12872) );
  NAND2_X1 U15980 ( .A1(n12873), .A2(n12872), .ZN(n17064) );
  NAND2_X1 U15981 ( .A1(n17064), .A2(n17073), .ZN(n12877) );
  NOR2_X1 U15982 ( .A1(n19598), .A2(n20606), .ZN(n16556) );
  INV_X1 U15983 ( .A(n16556), .ZN(n17087) );
  OAI22_X1 U15984 ( .A1(n17087), .A2(n12874), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n21204), .ZN(n12875) );
  INV_X1 U15985 ( .A(n12875), .ZN(n12876) );
  NAND2_X1 U15986 ( .A1(n12877), .A2(n12876), .ZN(n20573) );
  INV_X1 U15987 ( .A(n20573), .ZN(n20571) );
  NAND2_X1 U15988 ( .A1(n12973), .A2(n12878), .ZN(n17048) );
  OR4_X1 U15989 ( .A1(n20571), .A2(n20568), .A3(n17047), .A4(n17048), .ZN(
        n12879) );
  OAI21_X1 U15990 ( .B1(n17060), .B2(n20573), .A(n12879), .ZN(P2_U3595) );
  INV_X1 U15991 ( .A(n17069), .ZN(n20509) );
  NOR2_X1 U15992 ( .A1(n12881), .A2(n20509), .ZN(n13718) );
  AND2_X1 U15993 ( .A1(n12880), .A2(n13718), .ZN(n12882) );
  AOI22_X1 U15994 ( .A1(n12913), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12888) );
  INV_X1 U15995 ( .A(n12882), .ZN(n12883) );
  NOR2_X2 U15996 ( .A1(n12883), .A2(n17076), .ZN(n12954) );
  INV_X1 U15997 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12884) );
  OR2_X1 U15998 ( .A1(n13858), .A2(n12884), .ZN(n12886) );
  NAND2_X1 U15999 ( .A1(n13858), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12885) );
  AND2_X1 U16000 ( .A1(n12886), .A2(n12885), .ZN(n19826) );
  INV_X1 U16001 ( .A(n19826), .ZN(n12887) );
  NAND2_X1 U16002 ( .A1(n12954), .A2(n12887), .ZN(n12930) );
  NAND2_X1 U16003 ( .A1(n12888), .A2(n12930), .ZN(P2_U2976) );
  AOI22_X1 U16004 ( .A1(n12913), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16005 ( .A1(n13860), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13858), .ZN(n19957) );
  INV_X1 U16006 ( .A(n19957), .ZN(n19837) );
  NAND2_X1 U16007 ( .A1(n12954), .A2(n19837), .ZN(n12938) );
  NAND2_X1 U16008 ( .A1(n12889), .A2(n12938), .ZN(P2_U2972) );
  AOI22_X1 U16009 ( .A1(n12913), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16010 ( .A1(n13860), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13858), .ZN(n19868) );
  INV_X1 U16011 ( .A(n19868), .ZN(n14101) );
  NAND2_X1 U16012 ( .A1(n12954), .A2(n14101), .ZN(n12942) );
  NAND2_X1 U16013 ( .A1(n12890), .A2(n12942), .ZN(P2_U2953) );
  AOI22_X1 U16014 ( .A1(n12913), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U16015 ( .A1(n13860), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13858), .ZN(n19947) );
  INV_X1 U16016 ( .A(n19947), .ZN(n15654) );
  NAND2_X1 U16017 ( .A1(n12954), .A2(n15654), .ZN(n12944) );
  NAND2_X1 U16018 ( .A1(n12891), .A2(n12944), .ZN(P2_U2970) );
  AOI22_X1 U16019 ( .A1(n12913), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U16020 ( .A1(n13860), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13858), .ZN(n19831) );
  INV_X1 U16021 ( .A(n19831), .ZN(n12892) );
  NAND2_X1 U16022 ( .A1(n12954), .A2(n12892), .ZN(n12936) );
  NAND2_X1 U16023 ( .A1(n12893), .A2(n12936), .ZN(P2_U2974) );
  AOI22_X1 U16024 ( .A1(n12913), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12897) );
  INV_X1 U16025 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14147) );
  OR2_X1 U16026 ( .A1(n13858), .A2(n14147), .ZN(n12895) );
  NAND2_X1 U16027 ( .A1(n13858), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12894) );
  AND2_X1 U16028 ( .A1(n12895), .A2(n12894), .ZN(n19821) );
  INV_X1 U16029 ( .A(n19821), .ZN(n12896) );
  NAND2_X1 U16030 ( .A1(n12954), .A2(n12896), .ZN(n12928) );
  NAND2_X1 U16031 ( .A1(n12897), .A2(n12928), .ZN(P2_U2978) );
  AOI22_X1 U16032 ( .A1(n12913), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12898) );
  INV_X1 U16033 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n17209) );
  INV_X1 U16034 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21197) );
  AOI22_X1 U16035 ( .A1(n13860), .A2(n17209), .B1(n21197), .B2(n13858), .ZN(
        n19833) );
  NAND2_X1 U16036 ( .A1(n12954), .A2(n19833), .ZN(n12914) );
  NAND2_X1 U16037 ( .A1(n12898), .A2(n12914), .ZN(P2_U2973) );
  AOI22_X1 U16038 ( .A1(n12913), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12899) );
  INV_X1 U16039 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n17213) );
  INV_X1 U16040 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18937) );
  AOI22_X1 U16041 ( .A1(n13860), .A2(n17213), .B1(n18937), .B2(n13858), .ZN(
        n19845) );
  NAND2_X1 U16042 ( .A1(n12954), .A2(n19845), .ZN(n12926) );
  NAND2_X1 U16043 ( .A1(n12899), .A2(n12926), .ZN(P2_U2971) );
  NAND3_X1 U16044 ( .A1(n12902), .A2(n12901), .A3(n12900), .ZN(n12903) );
  NAND2_X1 U16045 ( .A1(n12904), .A2(n12903), .ZN(n12906) );
  INV_X1 U16046 ( .A(n14955), .ZN(n12907) );
  NAND2_X1 U16047 ( .A1(n13116), .A2(n12907), .ZN(n12959) );
  NOR2_X1 U16048 ( .A1(n20893), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12993) );
  INV_X1 U16049 ( .A(n13199), .ZN(n12909) );
  AOI211_X1 U16050 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n12992), .A(n12993), 
        .B(n12909), .ZN(n12910) );
  INV_X1 U16051 ( .A(n12910), .ZN(P1_U2801) );
  INV_X1 U16052 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19879) );
  NAND2_X1 U16053 ( .A1(n12913), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12911) );
  MUX2_X1 U16054 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n13858), .Z(n19823) );
  NAND2_X1 U16055 ( .A1(n12954), .A2(n19823), .ZN(n12946) );
  OAI211_X1 U16056 ( .C1(n19879), .C2(n12986), .A(n12911), .B(n12946), .ZN(
        P2_U2977) );
  INV_X1 U16057 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19872) );
  NAND2_X1 U16058 ( .A1(n12913), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12912) );
  NAND2_X1 U16059 ( .A1(n12954), .A2(n19813), .ZN(n12952) );
  OAI211_X1 U16060 ( .C1(n19872), .C2(n12986), .A(n12912), .B(n12952), .ZN(
        P2_U2981) );
  INV_X1 U16061 ( .A(n12913), .ZN(n12987) );
  AOI22_X1 U16062 ( .A1(n12951), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n15341), .ZN(n12915) );
  NAND2_X1 U16063 ( .A1(n12915), .A2(n12914), .ZN(P2_U2958) );
  AOI22_X1 U16064 ( .A1(n12951), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n15341), .ZN(n12920) );
  INV_X1 U16065 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n12916) );
  OR2_X1 U16066 ( .A1(n13858), .A2(n12916), .ZN(n12918) );
  NAND2_X1 U16067 ( .A1(n13858), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12917) );
  AND2_X1 U16068 ( .A1(n12918), .A2(n12917), .ZN(n19829) );
  INV_X1 U16069 ( .A(n19829), .ZN(n12919) );
  NAND2_X1 U16070 ( .A1(n12954), .A2(n12919), .ZN(n12934) );
  NAND2_X1 U16071 ( .A1(n12920), .A2(n12934), .ZN(P2_U2960) );
  AOI22_X1 U16072 ( .A1(n12951), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n15341), .ZN(n12924) );
  INV_X1 U16073 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14373) );
  OR2_X1 U16074 ( .A1(n13858), .A2(n14373), .ZN(n12922) );
  NAND2_X1 U16075 ( .A1(n13858), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12921) );
  AND2_X1 U16076 ( .A1(n12922), .A2(n12921), .ZN(n19816) );
  INV_X1 U16077 ( .A(n19816), .ZN(n12923) );
  NAND2_X1 U16078 ( .A1(n12954), .A2(n12923), .ZN(n12932) );
  NAND2_X1 U16079 ( .A1(n12924), .A2(n12932), .ZN(P2_U2965) );
  AOI22_X1 U16080 ( .A1(n12951), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n15341), .ZN(n12925) );
  OAI22_X1 U16081 ( .A1(n13858), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13860), .ZN(n19942) );
  INV_X1 U16082 ( .A(n19942), .ZN(n16928) );
  NAND2_X1 U16083 ( .A1(n12954), .A2(n16928), .ZN(n12940) );
  NAND2_X1 U16084 ( .A1(n12925), .A2(n12940), .ZN(P2_U2954) );
  AOI22_X1 U16085 ( .A1(n12951), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n15341), .ZN(n12927) );
  NAND2_X1 U16086 ( .A1(n12927), .A2(n12926), .ZN(P2_U2956) );
  AOI22_X1 U16087 ( .A1(n12951), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n15341), .ZN(n12929) );
  NAND2_X1 U16088 ( .A1(n12929), .A2(n12928), .ZN(P2_U2963) );
  AOI22_X1 U16089 ( .A1(n12951), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n15341), .ZN(n12931) );
  NAND2_X1 U16090 ( .A1(n12931), .A2(n12930), .ZN(P2_U2961) );
  AOI22_X1 U16091 ( .A1(n12951), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n15341), .ZN(n12933) );
  NAND2_X1 U16092 ( .A1(n12933), .A2(n12932), .ZN(P2_U2980) );
  AOI22_X1 U16093 ( .A1(n12951), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U16094 ( .A1(n12935), .A2(n12934), .ZN(P2_U2975) );
  AOI22_X1 U16095 ( .A1(n12951), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12937) );
  NAND2_X1 U16096 ( .A1(n12937), .A2(n12936), .ZN(P2_U2959) );
  AOI22_X1 U16097 ( .A1(n12951), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12939) );
  NAND2_X1 U16098 ( .A1(n12939), .A2(n12938), .ZN(P2_U2957) );
  AOI22_X1 U16099 ( .A1(n12951), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12941) );
  NAND2_X1 U16100 ( .A1(n12941), .A2(n12940), .ZN(P2_U2969) );
  AOI22_X1 U16101 ( .A1(n12951), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12943) );
  NAND2_X1 U16102 ( .A1(n12943), .A2(n12942), .ZN(P2_U2968) );
  AOI22_X1 U16103 ( .A1(n12951), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n15341), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U16104 ( .A1(n12945), .A2(n12944), .ZN(P2_U2955) );
  NAND2_X1 U16105 ( .A1(n12951), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12947) );
  OAI211_X1 U16106 ( .C1(n15612), .C2(n12986), .A(n12947), .B(n12946), .ZN(
        P2_U2962) );
  INV_X1 U16107 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n12982) );
  NAND2_X1 U16108 ( .A1(n12951), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12948) );
  MUX2_X1 U16109 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n13858), .Z(n19818) );
  NAND2_X1 U16110 ( .A1(n12954), .A2(n19818), .ZN(n12949) );
  OAI211_X1 U16111 ( .C1(n12982), .C2(n12986), .A(n12948), .B(n12949), .ZN(
        P2_U2964) );
  INV_X1 U16112 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19876) );
  NAND2_X1 U16113 ( .A1(n12951), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12950) );
  OAI211_X1 U16114 ( .C1(n19876), .C2(n12986), .A(n12950), .B(n12949), .ZN(
        P2_U2979) );
  NAND2_X1 U16115 ( .A1(n12951), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12953) );
  OAI211_X1 U16116 ( .C1(n12637), .C2(n12986), .A(n12953), .B(n12952), .ZN(
        P2_U2966) );
  INV_X1 U16117 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12956) );
  INV_X1 U16118 ( .A(n12954), .ZN(n12985) );
  AOI22_X1 U16119 ( .A1(n13860), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13858), .ZN(n19811) );
  INV_X1 U16120 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12955) );
  OAI222_X1 U16121 ( .A1(n12956), .A2(n12987), .B1(n12985), .B2(n19811), .C1(
        n12986), .C2(n12955), .ZN(P2_U2982) );
  INV_X1 U16122 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12958) );
  OAI22_X1 U16123 ( .A1(n13858), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13860), .ZN(n19937) );
  OAI222_X1 U16124 ( .A1(n12958), .A2(n12987), .B1(n12985), .B2(n19937), .C1(
        n12986), .C2(n12957), .ZN(P2_U2967) );
  NAND2_X1 U16125 ( .A1(n12908), .A2(n12959), .ZN(n12961) );
  NAND2_X1 U16126 ( .A1(n14963), .A2(n13576), .ZN(n12960) );
  NAND2_X1 U16127 ( .A1(n12961), .A2(n12960), .ZN(n20634) );
  NAND2_X1 U16128 ( .A1(n13578), .A2(n16528), .ZN(n12964) );
  INV_X1 U16129 ( .A(n12962), .ZN(n12963) );
  NAND2_X1 U16130 ( .A1(n12963), .A2(n20972), .ZN(n16554) );
  NAND2_X1 U16131 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21051) );
  AOI21_X1 U16132 ( .B1(n12964), .B2(n16554), .A(n20973), .ZN(n21053) );
  OR2_X1 U16133 ( .A1(n20634), .A2(n21053), .ZN(n16522) );
  AND2_X1 U16134 ( .A1(n16522), .A2(n14967), .ZN(n20642) );
  INV_X1 U16135 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12972) );
  NOR2_X1 U16136 ( .A1(n13576), .A2(n12965), .ZN(n12966) );
  NAND2_X1 U16137 ( .A1(n11532), .A2(n12966), .ZN(n14969) );
  NAND3_X1 U16138 ( .A1(n12908), .A2(n16520), .A3(n14969), .ZN(n12967) );
  MUX2_X1 U16139 ( .A(n12967), .B(n14981), .S(n14959), .Z(n12968) );
  INV_X1 U16140 ( .A(n12968), .ZN(n12970) );
  NAND2_X1 U16141 ( .A1(n13116), .A2(n14955), .ZN(n12969) );
  NAND2_X1 U16142 ( .A1(n12970), .A2(n12969), .ZN(n16523) );
  NAND2_X1 U16143 ( .A1(n20642), .A2(n16523), .ZN(n12971) );
  OAI21_X1 U16144 ( .B1(n20642), .B2(n12972), .A(n12971), .ZN(P1_U3484) );
  NAND3_X1 U16145 ( .A1(n13707), .A2(n12973), .A3(n17073), .ZN(n12974) );
  NAND2_X1 U16146 ( .A1(n12974), .A2(n12986), .ZN(n12975) );
  NAND2_X1 U16147 ( .A1(n19869), .A2(n12976), .ZN(n13028) );
  NOR2_X1 U16148 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20606), .ZN(n19892) );
  AOI22_X1 U16149 ( .A1(n19900), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12977) );
  OAI21_X1 U16150 ( .B1(n15631), .B2(n13028), .A(n12977), .ZN(P2_U2927) );
  INV_X1 U16151 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15593) );
  AOI22_X1 U16152 ( .A1(n19900), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12978) );
  OAI21_X1 U16153 ( .B1(n15593), .B2(n13028), .A(n12978), .ZN(P2_U2922) );
  INV_X1 U16154 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15620) );
  AOI22_X1 U16155 ( .A1(n19900), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12979) );
  OAI21_X1 U16156 ( .B1(n15620), .B2(n13028), .A(n12979), .ZN(P2_U2926) );
  AOI22_X1 U16157 ( .A1(n19900), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12980) );
  OAI21_X1 U16158 ( .B1(n12637), .B2(n13028), .A(n12980), .ZN(P2_U2921) );
  AOI22_X1 U16159 ( .A1(n19900), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12981) );
  OAI21_X1 U16160 ( .B1(n12982), .B2(n13028), .A(n12981), .ZN(P2_U2923) );
  AOI22_X1 U16161 ( .A1(n19900), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12983) );
  OAI21_X1 U16162 ( .B1(n15612), .B2(n13028), .A(n12983), .ZN(P2_U2925) );
  AOI22_X1 U16163 ( .A1(n19900), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12984) );
  OAI21_X1 U16164 ( .B1(n15603), .B2(n13028), .A(n12984), .ZN(P2_U2924) );
  INV_X1 U16165 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12988) );
  INV_X1 U16166 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13023) );
  OAI222_X1 U16167 ( .A1(n12988), .A2(n12987), .B1(n12986), .B2(n13023), .C1(
        n12985), .C2(n19937), .ZN(P2_U2952) );
  INV_X1 U16168 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19941) );
  NAND2_X1 U16169 ( .A1(n17047), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12989) );
  AND4_X1 U16170 ( .A1(n12989), .A2(n19962), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n21204), .ZN(n12990) );
  MUX2_X1 U16171 ( .A(n15507), .B(n17014), .S(n19784), .Z(n12991) );
  OAI21_X1 U16172 ( .B1(n20609), .B2(n19788), .A(n12991), .ZN(P2_U2887) );
  OAI21_X1 U16173 ( .B1(n12993), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13574), 
        .ZN(n12994) );
  OAI21_X1 U16174 ( .B1(n12995), .B2(n13574), .A(n12994), .ZN(P1_U3487) );
  OAI21_X1 U16175 ( .B1(n12997), .B2(n14078), .A(n12996), .ZN(n12998) );
  XOR2_X1 U16176 ( .A(n12998), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n16204) );
  INV_X1 U16177 ( .A(n16204), .ZN(n13005) );
  INV_X1 U16178 ( .A(n16957), .ZN(n15927) );
  OAI21_X1 U16179 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13000), .A(
        n12999), .ZN(n16205) );
  INV_X1 U16180 ( .A(n16205), .ZN(n13001) );
  AND2_X1 U16181 ( .A1(n19903), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n16207) );
  AOI21_X1 U16182 ( .B1(n15933), .B2(n13001), .A(n16207), .ZN(n13003) );
  NAND2_X1 U16183 ( .A1(n16942), .A2(n14076), .ZN(n13002) );
  OAI211_X1 U16184 ( .C1(n14076), .C2(n16950), .A(n13003), .B(n13002), .ZN(
        n13004) );
  AOI21_X1 U16185 ( .B1(n13005), .B2(n15927), .A(n13004), .ZN(n13006) );
  OAI21_X1 U16186 ( .B1(n16217), .B2(n13859), .A(n13006), .ZN(P2_U3013) );
  NOR2_X1 U16187 ( .A1(n13009), .A2(n13008), .ZN(n13010) );
  NOR2_X1 U16188 ( .A1(n13011), .A2(n13010), .ZN(n15510) );
  INV_X1 U16189 ( .A(n15510), .ZN(n17015) );
  NOR2_X1 U16190 ( .A1(n20609), .A2(n17015), .ZN(n19862) );
  INV_X1 U16191 ( .A(n19862), .ZN(n13012) );
  OAI211_X1 U16192 ( .C1(n16222), .C2(n15510), .A(n13012), .B(n19848), .ZN(
        n13014) );
  AOI22_X1 U16193 ( .A1(n19859), .A2(n15510), .B1(n19858), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13013) );
  OAI211_X1 U16194 ( .C1(n19867), .C2(n19937), .A(n13014), .B(n13013), .ZN(
        P2_U2919) );
  INV_X1 U16195 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13016) );
  AOI22_X1 U16196 ( .A1(n19900), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13015) );
  OAI21_X1 U16197 ( .B1(n13016), .B2(n13028), .A(n13015), .ZN(P2_U2932) );
  AOI22_X1 U16198 ( .A1(n19900), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13017) );
  OAI21_X1 U16199 ( .B1(n15639), .B2(n13028), .A(n13017), .ZN(P2_U2928) );
  INV_X1 U16200 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13019) );
  AOI22_X1 U16201 ( .A1(n19900), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13018) );
  OAI21_X1 U16202 ( .B1(n13019), .B2(n13028), .A(n13018), .ZN(P2_U2930) );
  INV_X1 U16203 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U16204 ( .A1(n19900), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13020) );
  OAI21_X1 U16205 ( .B1(n13021), .B2(n13028), .A(n13020), .ZN(P2_U2933) );
  AOI22_X1 U16206 ( .A1(n19900), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13022) );
  OAI21_X1 U16207 ( .B1(n13023), .B2(n13028), .A(n13022), .ZN(P2_U2935) );
  INV_X1 U16208 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U16209 ( .A1(n19900), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13024) );
  OAI21_X1 U16210 ( .B1(n13025), .B2(n13028), .A(n13024), .ZN(P2_U2931) );
  INV_X1 U16211 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n21115) );
  AOI22_X1 U16212 ( .A1(n19900), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13026) );
  OAI21_X1 U16213 ( .B1(n21115), .B2(n13028), .A(n13026), .ZN(P2_U2934) );
  INV_X1 U16214 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13029) );
  AOI22_X1 U16215 ( .A1(n19900), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13027) );
  OAI21_X1 U16216 ( .B1(n13029), .B2(n13028), .A(n13027), .ZN(P2_U2929) );
  INV_X1 U16217 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20852) );
  INV_X1 U16218 ( .A(n13030), .ZN(n13031) );
  AOI21_X1 U16219 ( .B1(n13032), .B2(n20852), .A(n13031), .ZN(n20848) );
  INV_X1 U16220 ( .A(n20848), .ZN(n13039) );
  INV_X1 U16221 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13038) );
  INV_X1 U16222 ( .A(n13033), .ZN(n13037) );
  INV_X1 U16223 ( .A(n13034), .ZN(n13036) );
  OAI21_X1 U16224 ( .B1(n13037), .B2(n13036), .A(n13035), .ZN(n13705) );
  OAI222_X1 U16225 ( .A1(n13039), .A2(n14730), .B1(n13038), .B2(n20721), .C1(
        n13705), .C2(n14731), .ZN(P1_U2872) );
  AND2_X1 U16226 ( .A1(n13116), .A2(n14978), .ZN(n16508) );
  NAND3_X1 U16227 ( .A1(n16508), .A2(n14967), .A3(n14959), .ZN(n13040) );
  OAI21_X1 U16228 ( .B1(n13199), .B2(n14978), .A(n13040), .ZN(n13041) );
  INV_X1 U16229 ( .A(n16554), .ZN(n14953) );
  NAND2_X1 U16230 ( .A1(n20724), .A2(n14957), .ZN(n13241) );
  NAND2_X1 U16231 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n16848) );
  NAND2_X1 U16232 ( .A1(n20963), .A2(n13181), .ZN(n20726) );
  INV_X2 U16233 ( .A(n20726), .ZN(n20736) );
  NOR2_X4 U16234 ( .A1(n20724), .A2(n20736), .ZN(n20737) );
  AOI22_X1 U16235 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13042) );
  OAI21_X1 U16236 ( .B1(n11802), .B2(n13241), .A(n13042), .ZN(P1_U2909) );
  INV_X1 U16237 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13044) );
  AOI22_X1 U16238 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13043) );
  OAI21_X1 U16239 ( .B1(n13044), .B2(n13241), .A(n13043), .ZN(P1_U2912) );
  INV_X1 U16240 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U16241 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13045) );
  OAI21_X1 U16242 ( .B1(n13046), .B2(n13241), .A(n13045), .ZN(P1_U2910) );
  AOI22_X1 U16243 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13047) );
  OAI21_X1 U16244 ( .B1(n11755), .B2(n13241), .A(n13047), .ZN(P1_U2911) );
  INV_X1 U16245 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U16246 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13048) );
  OAI21_X1 U16247 ( .B1(n13049), .B2(n13241), .A(n13048), .ZN(P1_U2908) );
  INV_X1 U16248 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13051) );
  AOI22_X1 U16249 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13050) );
  OAI21_X1 U16250 ( .B1(n13051), .B2(n13241), .A(n13050), .ZN(P1_U2907) );
  INV_X1 U16251 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U16252 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13052) );
  OAI21_X1 U16253 ( .B1(n13053), .B2(n13241), .A(n13052), .ZN(P1_U2906) );
  NOR2_X1 U16254 ( .A1(n19796), .A2(n16217), .ZN(n13056) );
  AOI21_X1 U16255 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n19796), .A(n13056), .ZN(
        n13057) );
  OAI21_X1 U16256 ( .B1(n16223), .B2(n19788), .A(n13057), .ZN(P2_U2886) );
  NAND2_X1 U16257 ( .A1(n13059), .A2(n13058), .ZN(n13060) );
  MUX2_X1 U16258 ( .A(n13062), .B(n14126), .S(n19796), .Z(n13063) );
  OAI21_X1 U16259 ( .B1(n20054), .B2(n19788), .A(n13063), .ZN(P2_U2885) );
  OAI21_X1 U16260 ( .B1(n13065), .B2(n13064), .A(n13269), .ZN(n13601) );
  OR2_X1 U16261 ( .A1(n13067), .A2(n13066), .ZN(n13069) );
  AND2_X1 U16262 ( .A1(n13069), .A2(n13068), .ZN(n20837) );
  INV_X1 U16263 ( .A(n20837), .ZN(n13595) );
  AOI22_X1 U16264 ( .A1(n13595), .A2(n20717), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14715), .ZN(n13070) );
  OAI21_X1 U16265 ( .B1(n13601), .B2(n14731), .A(n13070), .ZN(P1_U2871) );
  OAI21_X1 U16266 ( .B1(n13071), .B2(n20973), .A(n14969), .ZN(n13072) );
  NAND2_X1 U16267 ( .A1(n13074), .A2(n13073), .ZN(n13075) );
  NAND2_X1 U16268 ( .A1(n9614), .A2(n13297), .ZN(n13080) );
  INV_X1 U16269 ( .A(n13080), .ZN(n13078) );
  INV_X1 U16270 ( .A(n14378), .ZN(n13081) );
  INV_X1 U16271 ( .A(n14738), .ZN(n14377) );
  NAND2_X1 U16272 ( .A1(n14377), .A2(DATAI_0_), .ZN(n13083) );
  NAND2_X1 U16273 ( .A1(n14738), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13082) );
  AND2_X1 U16274 ( .A1(n13083), .A2(n13082), .ZN(n13305) );
  INV_X1 U16275 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20749) );
  OAI222_X1 U16276 ( .A1(n14805), .A2(n13705), .B1(n14804), .B2(n13305), .C1(
        n14802), .C2(n20749), .ZN(P1_U2904) );
  NAND2_X1 U16277 ( .A1(n14377), .A2(DATAI_1_), .ZN(n13085) );
  NAND2_X1 U16278 ( .A1(n14738), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13084) );
  AND2_X1 U16279 ( .A1(n13085), .A2(n13084), .ZN(n14789) );
  INV_X1 U16280 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20746) );
  OAI222_X1 U16281 ( .A1(n14805), .A2(n13601), .B1(n14789), .B2(n14804), .C1(
        n14802), .C2(n20746), .ZN(P1_U2903) );
  INV_X1 U16282 ( .A(n13087), .ZN(n13088) );
  NAND2_X1 U16283 ( .A1(n12171), .A2(n13088), .ZN(n13089) );
  NOR2_X1 U16284 ( .A1(n14113), .A2(n19796), .ZN(n13091) );
  AOI21_X1 U16285 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n19796), .A(n13091), .ZN(
        n13092) );
  OAI21_X1 U16286 ( .B1(n20570), .B2(n19788), .A(n13092), .ZN(P2_U2884) );
  INV_X1 U16287 ( .A(n13093), .ZN(n13095) );
  AOI21_X1 U16288 ( .B1(n13095), .B2(n20852), .A(n13094), .ZN(n20840) );
  INV_X1 U16289 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13096) );
  NOR2_X1 U16290 ( .A1(n16817), .A2(n13096), .ZN(n20841) );
  INV_X1 U16291 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13700) );
  AOI21_X1 U16292 ( .B1(n14947), .B2(n13097), .A(n13700), .ZN(n13098) );
  AOI211_X1 U16293 ( .C1(n20840), .C2(n20792), .A(n20841), .B(n13098), .ZN(
        n13099) );
  OAI21_X1 U16294 ( .B1(n21063), .B2(n13705), .A(n13099), .ZN(P1_U2999) );
  XOR2_X1 U16295 ( .A(n13100), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13105)
         );
  AOI21_X1 U16296 ( .B1(n13102), .B2(n13101), .A(n13191), .ZN(n15921) );
  INV_X1 U16297 ( .A(n15921), .ZN(n19725) );
  NOR2_X1 U16298 ( .A1(n19796), .A2(n19725), .ZN(n13103) );
  AOI21_X1 U16299 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n19796), .A(n13103), .ZN(
        n13104) );
  OAI21_X1 U16300 ( .B1(n13105), .B2(n19788), .A(n13104), .ZN(P2_U2882) );
  NOR2_X1 U16301 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20962), .ZN(n13167) );
  OR2_X1 U16302 ( .A1(n16554), .A2(n20973), .ZN(n13106) );
  OR2_X1 U16303 ( .A1(n14963), .A2(n13106), .ZN(n16529) );
  NAND2_X1 U16304 ( .A1(n13107), .A2(n16529), .ZN(n13109) );
  INV_X1 U16305 ( .A(n14969), .ZN(n13144) );
  OR3_X1 U16306 ( .A1(n16508), .A2(n13134), .A3(n13144), .ZN(n13108) );
  NAND2_X1 U16307 ( .A1(n13109), .A2(n13108), .ZN(n13123) );
  NAND2_X1 U16308 ( .A1(n13110), .A2(n14970), .ZN(n13111) );
  NAND2_X1 U16309 ( .A1(n13111), .A2(n14957), .ZN(n13114) );
  AOI21_X1 U16310 ( .B1(n13114), .B2(n13113), .A(n13112), .ZN(n13131) );
  OR2_X1 U16311 ( .A1(n13115), .A2(n13131), .ZN(n13118) );
  INV_X1 U16312 ( .A(n13116), .ZN(n13117) );
  NAND2_X1 U16313 ( .A1(n13118), .A2(n13117), .ZN(n14965) );
  OR2_X1 U16314 ( .A1(n13578), .A2(n13309), .ZN(n13119) );
  AND4_X1 U16315 ( .A1(n13121), .A2(n14965), .A3(n13120), .A4(n13119), .ZN(
        n13122) );
  INV_X1 U16316 ( .A(n15162), .ZN(n14656) );
  INV_X1 U16317 ( .A(n13578), .ZN(n13125) );
  OAI21_X1 U16318 ( .B1(n13127), .B2(n13126), .A(n13125), .ZN(n13129) );
  NAND2_X1 U16319 ( .A1(n13129), .A2(n13128), .ZN(n13130) );
  NOR2_X1 U16320 ( .A1(n13131), .A2(n13130), .ZN(n13132) );
  AND2_X1 U16321 ( .A1(n13133), .A2(n13132), .ZN(n14985) );
  INV_X1 U16322 ( .A(n13134), .ZN(n13135) );
  AND4_X1 U16323 ( .A1(n13135), .A2(n13173), .A3(n13137), .A4(n13136), .ZN(
        n13138) );
  NAND2_X1 U16324 ( .A1(n14985), .A2(n13138), .ZN(n15169) );
  INV_X1 U16325 ( .A(n13139), .ZN(n13143) );
  INV_X1 U16326 ( .A(n13140), .ZN(n15170) );
  NAND2_X1 U16327 ( .A1(n15170), .A2(n13141), .ZN(n13142) );
  NAND2_X1 U16328 ( .A1(n13143), .A2(n13142), .ZN(n13145) );
  NOR3_X1 U16329 ( .A1(n15169), .A2(n13155), .A3(n13145), .ZN(n13148) );
  INV_X1 U16330 ( .A(n16508), .ZN(n15173) );
  XNOR2_X1 U16331 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13146) );
  NOR2_X1 U16332 ( .A1(n13144), .A2(n14981), .ZN(n13159) );
  INV_X1 U16333 ( .A(n13145), .ZN(n15182) );
  OAI22_X1 U16334 ( .A1(n15173), .A2(n13146), .B1(n13159), .B2(n15182), .ZN(
        n13147) );
  AOI211_X1 U16335 ( .C1(n14656), .C2(n15169), .A(n13148), .B(n13147), .ZN(
        n15184) );
  NAND2_X1 U16336 ( .A1(n13175), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13149) );
  OAI21_X1 U16337 ( .B1(n13175), .B2(n15184), .A(n13149), .ZN(n16512) );
  AOI22_X1 U16338 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13167), .B1(
        n20962), .B2(n16512), .ZN(n13169) );
  INV_X1 U16339 ( .A(n13152), .ZN(n13151) );
  MUX2_X1 U16340 ( .A(n13152), .B(n13151), .S(n13164), .Z(n13162) );
  OAI21_X1 U16341 ( .B1(n13139), .B2(n13164), .A(n13153), .ZN(n13154) );
  INV_X1 U16342 ( .A(n13154), .ZN(n15187) );
  OR3_X1 U16343 ( .A1(n15169), .A2(n15187), .A3(n13155), .ZN(n13161) );
  MUX2_X1 U16344 ( .A(n13156), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13140), .Z(n13157) );
  OR3_X1 U16345 ( .A1(n13159), .A2(n13158), .A3(n13157), .ZN(n13160) );
  OAI211_X1 U16346 ( .C1(n13162), .C2(n15173), .A(n13161), .B(n13160), .ZN(
        n13163) );
  AOI21_X1 U16347 ( .B1(n13150), .B2(n15169), .A(n13163), .ZN(n15188) );
  NAND2_X1 U16348 ( .A1(n15188), .A2(n16503), .ZN(n13166) );
  NAND2_X1 U16349 ( .A1(n13175), .A2(n13164), .ZN(n13165) );
  AOI22_X1 U16350 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13167), .B1(
        n16514), .B2(n20962), .ZN(n13168) );
  NOR2_X1 U16351 ( .A1(n13169), .A2(n13168), .ZN(n16517) );
  INV_X1 U16352 ( .A(n13170), .ZN(n15174) );
  INV_X1 U16353 ( .A(n13420), .ZN(n13326) );
  OR2_X1 U16354 ( .A1(n13171), .A2(n13326), .ZN(n13172) );
  XNOR2_X1 U16355 ( .A(n13172), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20699) );
  INV_X1 U16356 ( .A(n13173), .ZN(n13174) );
  NAND2_X1 U16357 ( .A1(n20699), .A2(n13174), .ZN(n16840) );
  NOR2_X1 U16358 ( .A1(n13175), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13176) );
  NAND2_X1 U16359 ( .A1(n16840), .A2(n13176), .ZN(n13179) );
  INV_X1 U16360 ( .A(n13176), .ZN(n13177) );
  AOI22_X1 U16361 ( .A1(n13177), .A2(n11894), .B1(P1_STATE2_REG_1__SCAN_IN), 
        .B2(P1_FLUSH_REG_SCAN_IN), .ZN(n13178) );
  AOI21_X1 U16362 ( .B1(n16517), .B2(n15174), .A(n16518), .ZN(n13182) );
  NOR2_X1 U16363 ( .A1(n20963), .A2(n16848), .ZN(n16851) );
  INV_X1 U16364 ( .A(n16851), .ZN(n13180) );
  NOR2_X1 U16365 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21054) );
  NAND2_X1 U16366 ( .A1(n16851), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n14447) );
  OAI211_X1 U16367 ( .C1(n13182), .C2(n13180), .A(n13768), .B(n14447), .ZN(
        n20853) );
  NAND2_X1 U16368 ( .A1(n13182), .A2(n13181), .ZN(n16535) );
  INV_X1 U16369 ( .A(n16535), .ZN(n13185) );
  AND2_X1 U16370 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20905), .ZN(n15166) );
  OAI22_X1 U16371 ( .A1(n9606), .A2(n20893), .B1(n14445), .B2(n15166), .ZN(
        n13184) );
  OAI21_X1 U16372 ( .B1(n13185), .B2(n13184), .A(n20853), .ZN(n13186) );
  OAI21_X1 U16373 ( .B1(n20853), .B2(n20864), .A(n13186), .ZN(P1_U3478) );
  NOR2_X1 U16374 ( .A1(n13100), .A2(n19960), .ZN(n13188) );
  OR2_X1 U16375 ( .A1(n13100), .A2(n13187), .ZN(n13242) );
  OAI211_X1 U16376 ( .C1(n13188), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19793), .B(n13242), .ZN(n13197) );
  INV_X1 U16377 ( .A(n13189), .ZN(n13195) );
  INV_X1 U16378 ( .A(n13190), .ZN(n13193) );
  INV_X1 U16379 ( .A(n13191), .ZN(n13192) );
  NAND2_X1 U16380 ( .A1(n13193), .A2(n13192), .ZN(n13194) );
  NAND2_X1 U16381 ( .A1(n13195), .A2(n13194), .ZN(n19715) );
  INV_X1 U16382 ( .A(n19715), .ZN(n16195) );
  NAND2_X1 U16383 ( .A1(n19784), .A2(n16195), .ZN(n13196) );
  OAI211_X1 U16384 ( .C1(n19784), .C2(n10329), .A(n13197), .B(n13196), .ZN(
        P2_U2881) );
  AND2_X1 U16385 ( .A1(n16528), .A2(n20973), .ZN(n13198) );
  NAND2_X1 U16386 ( .A1(n14377), .A2(DATAI_2_), .ZN(n13201) );
  NAND2_X1 U16387 ( .A1(n14738), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13200) );
  AND2_X1 U16388 ( .A1(n13201), .A2(n13200), .ZN(n14782) );
  INV_X1 U16389 ( .A(n14782), .ZN(n13202) );
  NAND2_X1 U16390 ( .A1(n9720), .A2(n13202), .ZN(n13260) );
  AOI22_X1 U16391 ( .A1(n20778), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20783), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13203) );
  NAND2_X1 U16392 ( .A1(n13260), .A2(n13203), .ZN(P1_U2954) );
  INV_X1 U16393 ( .A(DATAI_6_), .ZN(n13205) );
  NAND2_X1 U16394 ( .A1(n14738), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13204) );
  OAI21_X1 U16395 ( .B1(n14738), .B2(n13205), .A(n13204), .ZN(n14767) );
  NAND2_X1 U16396 ( .A1(n9720), .A2(n14767), .ZN(n13256) );
  AOI22_X1 U16397 ( .A1(n20778), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20783), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13206) );
  NAND2_X1 U16398 ( .A1(n13256), .A2(n13206), .ZN(P1_U2958) );
  NAND2_X1 U16399 ( .A1(n14377), .A2(DATAI_4_), .ZN(n13208) );
  NAND2_X1 U16400 ( .A1(n14738), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13207) );
  AND2_X1 U16401 ( .A1(n13208), .A2(n13207), .ZN(n13494) );
  INV_X1 U16402 ( .A(n13494), .ZN(n16641) );
  NAND2_X1 U16403 ( .A1(n9720), .A2(n16641), .ZN(n13252) );
  AOI22_X1 U16404 ( .A1(n20778), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20783), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13209) );
  NAND2_X1 U16405 ( .A1(n13252), .A2(n13209), .ZN(P1_U2956) );
  INV_X1 U16406 ( .A(DATAI_7_), .ZN(n13211) );
  NAND2_X1 U16407 ( .A1(n14738), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13210) );
  OAI21_X1 U16408 ( .B1(n14738), .B2(n13211), .A(n13210), .ZN(n14762) );
  NAND2_X1 U16409 ( .A1(n9720), .A2(n14762), .ZN(n13264) );
  AOI22_X1 U16410 ( .A1(n20778), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20783), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13212) );
  NAND2_X1 U16411 ( .A1(n13264), .A2(n13212), .ZN(P1_U2959) );
  NAND2_X1 U16412 ( .A1(n14377), .A2(DATAI_3_), .ZN(n13214) );
  NAND2_X1 U16413 ( .A1(n14738), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13213) );
  AND2_X1 U16414 ( .A1(n13214), .A2(n13213), .ZN(n14777) );
  INV_X1 U16415 ( .A(n14777), .ZN(n13215) );
  NAND2_X1 U16416 ( .A1(n9720), .A2(n13215), .ZN(n13262) );
  AOI22_X1 U16417 ( .A1(n20778), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20783), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13216) );
  NAND2_X1 U16418 ( .A1(n13262), .A2(n13216), .ZN(P1_U2955) );
  NAND2_X1 U16419 ( .A1(n14377), .A2(DATAI_5_), .ZN(n13218) );
  NAND2_X1 U16420 ( .A1(n14738), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13217) );
  AND2_X1 U16421 ( .A1(n13218), .A2(n13217), .ZN(n14772) );
  INV_X1 U16422 ( .A(n14772), .ZN(n13219) );
  NAND2_X1 U16423 ( .A1(n9720), .A2(n13219), .ZN(n13258) );
  AOI22_X1 U16424 ( .A1(n20778), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20783), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13220) );
  NAND2_X1 U16425 ( .A1(n13258), .A2(n13220), .ZN(P1_U2957) );
  INV_X1 U16426 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13226) );
  INV_X1 U16427 ( .A(n9720), .ZN(n13225) );
  INV_X1 U16428 ( .A(DATAI_15_), .ZN(n13222) );
  INV_X1 U16429 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13221) );
  MUX2_X1 U16430 ( .A(n13222), .B(n13221), .S(n14738), .Z(n14795) );
  INV_X1 U16431 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13224) );
  OAI222_X1 U16432 ( .A1(n13247), .A2(n13226), .B1(n13225), .B2(n14795), .C1(
        n13224), .C2(n13223), .ZN(P1_U2967) );
  INV_X1 U16433 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13228) );
  AOI22_X1 U16434 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13227) );
  OAI21_X1 U16435 ( .B1(n13228), .B2(n13241), .A(n13227), .ZN(P1_U2914) );
  INV_X1 U16436 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13230) );
  AOI22_X1 U16437 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13229) );
  OAI21_X1 U16438 ( .B1(n13230), .B2(n13241), .A(n13229), .ZN(P1_U2917) );
  INV_X1 U16439 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13232) );
  AOI22_X1 U16440 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13231) );
  OAI21_X1 U16441 ( .B1(n13232), .B2(n13241), .A(n13231), .ZN(P1_U2920) );
  INV_X1 U16442 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13234) );
  AOI22_X1 U16443 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13233) );
  OAI21_X1 U16444 ( .B1(n13234), .B2(n13241), .A(n13233), .ZN(P1_U2913) );
  INV_X1 U16445 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U16446 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13235) );
  OAI21_X1 U16447 ( .B1(n13236), .B2(n13241), .A(n13235), .ZN(P1_U2916) );
  INV_X1 U16448 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21114) );
  AOI22_X1 U16449 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13237) );
  OAI21_X1 U16450 ( .B1(n21114), .B2(n13241), .A(n13237), .ZN(P1_U2915) );
  INV_X1 U16451 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13239) );
  AOI22_X1 U16452 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13238) );
  OAI21_X1 U16453 ( .B1(n13239), .B2(n13241), .A(n13238), .ZN(P1_U2918) );
  AOI22_X1 U16454 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13240) );
  OAI21_X1 U16455 ( .B1(n14787), .B2(n13241), .A(n13240), .ZN(P1_U2919) );
  XOR2_X1 U16456 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13242), .Z(n13246)
         );
  NOR2_X1 U16457 ( .A1(n13189), .A2(n13243), .ZN(n13244) );
  NOR2_X1 U16458 ( .A1(n14052), .A2(n13244), .ZN(n16182) );
  INV_X1 U16459 ( .A(n16182), .ZN(n19702) );
  MUX2_X1 U16460 ( .A(n10349), .B(n19702), .S(n19784), .Z(n13245) );
  OAI21_X1 U16461 ( .B1(n13246), .B2(n19788), .A(n13245), .ZN(P2_U2880) );
  INV_X1 U16462 ( .A(n13305), .ZN(n16646) );
  NAND2_X1 U16463 ( .A1(n9720), .A2(n16646), .ZN(n13250) );
  AOI22_X1 U16464 ( .A1(n20778), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20783), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13248) );
  NAND2_X1 U16465 ( .A1(n13250), .A2(n13248), .ZN(P1_U2952) );
  AOI22_X1 U16466 ( .A1(n20778), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13249) );
  NAND2_X1 U16467 ( .A1(n13250), .A2(n13249), .ZN(P1_U2937) );
  AOI22_X1 U16468 ( .A1(n20778), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13251) );
  NAND2_X1 U16469 ( .A1(n13252), .A2(n13251), .ZN(P1_U2941) );
  INV_X1 U16470 ( .A(n14789), .ZN(n13253) );
  NAND2_X1 U16471 ( .A1(n9720), .A2(n13253), .ZN(n13266) );
  AOI22_X1 U16472 ( .A1(n20778), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20783), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13254) );
  NAND2_X1 U16473 ( .A1(n13266), .A2(n13254), .ZN(P1_U2953) );
  AOI22_X1 U16474 ( .A1(n20778), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13255) );
  NAND2_X1 U16475 ( .A1(n13256), .A2(n13255), .ZN(P1_U2943) );
  AOI22_X1 U16476 ( .A1(n20778), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13257) );
  NAND2_X1 U16477 ( .A1(n13258), .A2(n13257), .ZN(P1_U2942) );
  AOI22_X1 U16478 ( .A1(n20778), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13259) );
  NAND2_X1 U16479 ( .A1(n13260), .A2(n13259), .ZN(P1_U2939) );
  AOI22_X1 U16480 ( .A1(n20778), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13261) );
  NAND2_X1 U16481 ( .A1(n13262), .A2(n13261), .ZN(P1_U2940) );
  AOI22_X1 U16482 ( .A1(n20778), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13263) );
  NAND2_X1 U16483 ( .A1(n13264), .A2(n13263), .ZN(P1_U2944) );
  AOI22_X1 U16484 ( .A1(n20778), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13265) );
  NAND2_X1 U16485 ( .A1(n13266), .A2(n13265), .ZN(P1_U2938) );
  INV_X1 U16486 ( .A(n13267), .ZN(n13268) );
  AOI21_X1 U16487 ( .B1(n13270), .B2(n13269), .A(n13268), .ZN(n14666) );
  INV_X1 U16488 ( .A(n14731), .ZN(n20718) );
  AND2_X1 U16489 ( .A1(n13272), .A2(n13271), .ZN(n13273) );
  OR2_X1 U16490 ( .A1(n13282), .A2(n13273), .ZN(n20815) );
  INV_X1 U16491 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13274) );
  OAI22_X1 U16492 ( .A1(n20815), .A2(n14730), .B1(n13274), .B2(n20721), .ZN(
        n13275) );
  AOI21_X1 U16493 ( .B1(n14666), .B2(n20718), .A(n13275), .ZN(n13276) );
  INV_X1 U16494 ( .A(n13276), .ZN(P1_U2870) );
  OR2_X1 U16495 ( .A1(n13278), .A2(n13277), .ZN(n13280) );
  NAND2_X1 U16496 ( .A1(n13280), .A2(n13279), .ZN(n13960) );
  INV_X1 U16497 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20742) );
  OAI222_X1 U16498 ( .A1(n14805), .A2(n13960), .B1(n14777), .B2(n14804), .C1(
        n14802), .C2(n20742), .ZN(P1_U2901) );
  OAI21_X1 U16499 ( .B1(n13282), .B2(n13281), .A(n20697), .ZN(n13945) );
  INV_X1 U16500 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13949) );
  OAI222_X1 U16501 ( .A1(n13945), .A2(n14730), .B1(n20721), .B2(n13949), .C1(
        n13960), .C2(n14731), .ZN(P1_U2869) );
  NOR2_X2 U16502 ( .A1(n21063), .A2(n14377), .ZN(n13317) );
  NOR2_X2 U16503 ( .A1(n14738), .A2(n21063), .ZN(n13318) );
  AOI22_X1 U16504 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n13317), .B1(DATAI_27_), 
        .B2(n13318), .ZN(n15215) );
  NAND2_X1 U16505 ( .A1(n12060), .A2(n13531), .ZN(n13283) );
  INV_X1 U16506 ( .A(n13286), .ZN(n13284) );
  NOR3_X1 U16507 ( .A1(n13284), .A2(n20640), .A3(n20893), .ZN(n13285) );
  NOR3_X1 U16508 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15192) );
  NAND2_X1 U16509 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13293) );
  NAND2_X1 U16510 ( .A1(n13286), .A2(n13663), .ZN(n13786) );
  AOI22_X1 U16511 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n13317), .B1(DATAI_19_), 
        .B2(n13318), .ZN(n15268) );
  INV_X1 U16512 ( .A(n15268), .ZN(n20929) );
  NAND2_X1 U16513 ( .A1(n13319), .A2(n13288), .ZN(n15269) );
  INV_X1 U16514 ( .A(n15192), .ZN(n13289) );
  OR2_X1 U16515 ( .A1(n20864), .A2(n13289), .ZN(n13321) );
  OR2_X1 U16516 ( .A1(n13150), .A2(n14656), .ZN(n15191) );
  OAI21_X1 U16517 ( .B1(n15191), .B2(n13653), .A(n13321), .ZN(n13290) );
  AOI22_X1 U16518 ( .A1(n13290), .A2(n13770), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15192), .ZN(n13320) );
  OAI22_X1 U16519 ( .A1(n15269), .A2(n13321), .B1(n13320), .B2(n20933), .ZN(
        n13291) );
  AOI21_X1 U16520 ( .B1(n13819), .B2(n20929), .A(n13291), .ZN(n13292) );
  OAI211_X1 U16521 ( .C1(n15215), .C2(n15238), .A(n13293), .B(n13292), .ZN(
        P1_U3044) );
  AOI22_X1 U16522 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n13317), .B1(DATAI_28_), 
        .B2(n13318), .ZN(n15220) );
  NAND2_X1 U16523 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13296) );
  AOI22_X1 U16524 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n13317), .B1(DATAI_20_), 
        .B2(n13318), .ZN(n15273) );
  INV_X1 U16525 ( .A(n15273), .ZN(n20935) );
  NAND2_X1 U16526 ( .A1(n13319), .A2(n14977), .ZN(n15274) );
  OAI22_X1 U16527 ( .A1(n15274), .A2(n13321), .B1(n13320), .B2(n20939), .ZN(
        n13294) );
  AOI21_X1 U16528 ( .B1(n13819), .B2(n20935), .A(n13294), .ZN(n13295) );
  OAI211_X1 U16529 ( .C1(n15220), .C2(n15238), .A(n13296), .B(n13295), .ZN(
        P1_U3045) );
  AOI22_X1 U16530 ( .A1(DATAI_31_), .A2(n13318), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n13317), .ZN(n15236) );
  NAND2_X1 U16531 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13300) );
  AOI22_X1 U16532 ( .A1(DATAI_23_), .A2(n13318), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n13317), .ZN(n15289) );
  INV_X1 U16533 ( .A(n15289), .ZN(n20954) );
  INV_X1 U16534 ( .A(n14762), .ZN(n13914) );
  NAND2_X1 U16535 ( .A1(n13319), .A2(n13297), .ZN(n15292) );
  OAI22_X1 U16536 ( .A1(n20960), .A2(n13320), .B1(n15292), .B2(n13321), .ZN(
        n13298) );
  AOI21_X1 U16537 ( .B1(n13819), .B2(n20954), .A(n13298), .ZN(n13299) );
  OAI211_X1 U16538 ( .C1(n15236), .C2(n15238), .A(n13300), .B(n13299), .ZN(
        P1_U3048) );
  AOI22_X1 U16539 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n13317), .B1(DATAI_30_), 
        .B2(n13318), .ZN(n15230) );
  NAND2_X1 U16540 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n13304) );
  AOI22_X1 U16541 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n13317), .B1(DATAI_22_), 
        .B2(n13318), .ZN(n15283) );
  INV_X1 U16542 ( .A(n15283), .ZN(n20947) );
  INV_X1 U16543 ( .A(n14767), .ZN(n13697) );
  NAND2_X1 U16544 ( .A1(n13319), .A2(n13301), .ZN(n15284) );
  OAI22_X1 U16545 ( .A1(n20951), .A2(n13320), .B1(n15284), .B2(n13321), .ZN(
        n13302) );
  AOI21_X1 U16546 ( .B1(n13819), .B2(n20947), .A(n13302), .ZN(n13303) );
  OAI211_X1 U16547 ( .C1(n15230), .C2(n15238), .A(n13304), .B(n13303), .ZN(
        P1_U3047) );
  AOI22_X1 U16548 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n13317), .B1(DATAI_24_), 
        .B2(n13318), .ZN(n15201) );
  NAND2_X1 U16549 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13308) );
  AOI22_X1 U16550 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n13317), .B1(DATAI_16_), 
        .B2(n13318), .ZN(n15253) );
  INV_X1 U16551 ( .A(n15253), .ZN(n20903) );
  NAND2_X1 U16552 ( .A1(n13319), .A2(n14957), .ZN(n15254) );
  OAI22_X1 U16553 ( .A1(n15254), .A2(n13321), .B1(n13320), .B2(n20915), .ZN(
        n13306) );
  AOI21_X1 U16554 ( .B1(n13819), .B2(n20903), .A(n13306), .ZN(n13307) );
  OAI211_X1 U16555 ( .C1(n15201), .C2(n15238), .A(n13308), .B(n13307), .ZN(
        P1_U3041) );
  AOI22_X1 U16556 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n13317), .B1(DATAI_26_), 
        .B2(n13318), .ZN(n15211) );
  NAND2_X1 U16557 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13312) );
  AOI22_X1 U16558 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n13317), .B1(DATAI_18_), 
        .B2(n13318), .ZN(n15263) );
  INV_X1 U16559 ( .A(n15263), .ZN(n20923) );
  NAND2_X1 U16560 ( .A1(n13319), .A2(n13309), .ZN(n15264) );
  OAI22_X1 U16561 ( .A1(n15264), .A2(n13321), .B1(n13320), .B2(n20927), .ZN(
        n13310) );
  AOI21_X1 U16562 ( .B1(n13819), .B2(n20923), .A(n13310), .ZN(n13311) );
  OAI211_X1 U16563 ( .C1(n15211), .C2(n15238), .A(n13312), .B(n13311), .ZN(
        P1_U3043) );
  AOI22_X1 U16564 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n13317), .B1(DATAI_25_), 
        .B2(n13318), .ZN(n15206) );
  NAND2_X1 U16565 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13315) );
  AOI22_X1 U16566 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n13317), .B1(DATAI_17_), 
        .B2(n13318), .ZN(n15258) );
  INV_X1 U16567 ( .A(n15258), .ZN(n20917) );
  NAND2_X1 U16568 ( .A1(n13319), .A2(n14978), .ZN(n15259) );
  OAI22_X1 U16569 ( .A1(n15259), .A2(n13321), .B1(n13320), .B2(n20921), .ZN(
        n13313) );
  AOI21_X1 U16570 ( .B1(n13819), .B2(n20917), .A(n13313), .ZN(n13314) );
  OAI211_X1 U16571 ( .C1(n15206), .C2(n15238), .A(n13315), .B(n13314), .ZN(
        P1_U3042) );
  AOI22_X1 U16572 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n13317), .B1(DATAI_29_), 
        .B2(n13318), .ZN(n15225) );
  NAND2_X1 U16573 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13324) );
  AOI22_X1 U16574 ( .A1(DATAI_21_), .A2(n13318), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n13317), .ZN(n15278) );
  INV_X1 U16575 ( .A(n15278), .ZN(n20941) );
  NAND2_X1 U16576 ( .A1(n13319), .A2(n11116), .ZN(n15279) );
  OAI22_X1 U16577 ( .A1(n15279), .A2(n13321), .B1(n13320), .B2(n20945), .ZN(
        n13322) );
  AOI21_X1 U16578 ( .B1(n13819), .B2(n20941), .A(n13322), .ZN(n13323) );
  OAI211_X1 U16579 ( .C1(n15225), .C2(n15238), .A(n13324), .B(n13323), .ZN(
        P1_U3046) );
  INV_X1 U16580 ( .A(n14666), .ZN(n13325) );
  INV_X1 U16581 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20744) );
  OAI222_X1 U16582 ( .A1(n14805), .A2(n13325), .B1(n14782), .B2(n14804), .C1(
        n14802), .C2(n20744), .ZN(P1_U2902) );
  NOR2_X1 U16583 ( .A1(n15162), .A2(n13326), .ZN(n20897) );
  INV_X1 U16584 ( .A(n14445), .ZN(n13699) );
  AND2_X1 U16585 ( .A1(n13327), .A2(n13699), .ZN(n13534) );
  INV_X1 U16586 ( .A(n13362), .ZN(n13354) );
  AOI21_X1 U16587 ( .B1(n20897), .B2(n13534), .A(n13354), .ZN(n13331) );
  INV_X1 U16588 ( .A(n13331), .ZN(n13328) );
  NAND2_X1 U16589 ( .A1(n13328), .A2(n15157), .ZN(n13330) );
  NAND2_X1 U16590 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13333), .ZN(n13329) );
  AND2_X1 U16591 ( .A1(n13330), .A2(n13329), .ZN(n13358) );
  OR2_X1 U16592 ( .A1(n13531), .A2(n20640), .ZN(n15161) );
  NOR2_X1 U16593 ( .A1(n12060), .A2(n15161), .ZN(n13416) );
  AOI21_X1 U16594 ( .B1(n13416), .B2(n13651), .A(n20893), .ZN(n13415) );
  NAND2_X1 U16595 ( .A1(n13415), .A2(n13331), .ZN(n13332) );
  OAI211_X1 U16596 ( .C1(n13770), .C2(n13333), .A(n13332), .B(n13536), .ZN(
        n13357) );
  NAND2_X1 U16597 ( .A1(n13357), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n13337) );
  NAND4_X1 U16598 ( .A1(n13334), .A2(n15158), .A3(n13663), .A4(n13651), .ZN(
        n15237) );
  NAND4_X1 U16599 ( .A1(n13334), .A2(n15158), .A3(n13651), .A4(n9606), .ZN(
        n13891) );
  OAI22_X1 U16600 ( .A1(n15289), .A2(n15237), .B1(n13891), .B2(n15236), .ZN(
        n13335) );
  AOI21_X1 U16601 ( .B1(n20952), .B2(n13354), .A(n13335), .ZN(n13336) );
  OAI211_X1 U16602 ( .C1(n13358), .C2(n20960), .A(n13337), .B(n13336), .ZN(
        P1_U3160) );
  NAND2_X1 U16603 ( .A1(n13357), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13340) );
  INV_X1 U16604 ( .A(n13891), .ZN(n13902) );
  INV_X1 U16605 ( .A(n15225), .ZN(n20942) );
  OAI22_X1 U16606 ( .A1(n13358), .A2(n20945), .B1(n15237), .B2(n15278), .ZN(
        n13338) );
  AOI21_X1 U16607 ( .B1(n13902), .B2(n20942), .A(n13338), .ZN(n13339) );
  OAI211_X1 U16608 ( .C1(n15279), .C2(n13362), .A(n13340), .B(n13339), .ZN(
        P1_U3158) );
  NAND2_X1 U16609 ( .A1(n13357), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13343) );
  INV_X1 U16610 ( .A(n15215), .ZN(n20930) );
  OAI22_X1 U16611 ( .A1(n13358), .A2(n20933), .B1(n15237), .B2(n15268), .ZN(
        n13341) );
  AOI21_X1 U16612 ( .B1(n13902), .B2(n20930), .A(n13341), .ZN(n13342) );
  OAI211_X1 U16613 ( .C1(n15269), .C2(n13362), .A(n13343), .B(n13342), .ZN(
        P1_U3156) );
  NAND2_X1 U16614 ( .A1(n13357), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13346) );
  INV_X1 U16615 ( .A(n15211), .ZN(n20924) );
  OAI22_X1 U16616 ( .A1(n13358), .A2(n20927), .B1(n15237), .B2(n15263), .ZN(
        n13344) );
  AOI21_X1 U16617 ( .B1(n13902), .B2(n20924), .A(n13344), .ZN(n13345) );
  OAI211_X1 U16618 ( .C1(n15264), .C2(n13362), .A(n13346), .B(n13345), .ZN(
        P1_U3155) );
  NAND2_X1 U16619 ( .A1(n13357), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13349) );
  INV_X1 U16620 ( .A(n15206), .ZN(n20918) );
  OAI22_X1 U16621 ( .A1(n13358), .A2(n20921), .B1(n15237), .B2(n15258), .ZN(
        n13347) );
  AOI21_X1 U16622 ( .B1(n13902), .B2(n20918), .A(n13347), .ZN(n13348) );
  OAI211_X1 U16623 ( .C1(n15259), .C2(n13362), .A(n13349), .B(n13348), .ZN(
        P1_U3154) );
  NAND2_X1 U16624 ( .A1(n13357), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13352) );
  INV_X1 U16625 ( .A(n15220), .ZN(n20936) );
  OAI22_X1 U16626 ( .A1(n13358), .A2(n20939), .B1(n15237), .B2(n15273), .ZN(
        n13350) );
  AOI21_X1 U16627 ( .B1(n13902), .B2(n20936), .A(n13350), .ZN(n13351) );
  OAI211_X1 U16628 ( .C1(n15274), .C2(n13362), .A(n13352), .B(n13351), .ZN(
        P1_U3157) );
  NAND2_X1 U16629 ( .A1(n13357), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n13356) );
  OAI22_X1 U16630 ( .A1(n15283), .A2(n15237), .B1(n13891), .B2(n15230), .ZN(
        n13353) );
  AOI21_X1 U16631 ( .B1(n20946), .B2(n13354), .A(n13353), .ZN(n13355) );
  OAI211_X1 U16632 ( .C1(n13358), .C2(n20951), .A(n13356), .B(n13355), .ZN(
        P1_U3159) );
  NAND2_X1 U16633 ( .A1(n13357), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13361) );
  INV_X1 U16634 ( .A(n15201), .ZN(n20912) );
  OAI22_X1 U16635 ( .A1(n13358), .A2(n20915), .B1(n15237), .B2(n15253), .ZN(
        n13359) );
  AOI21_X1 U16636 ( .B1(n13902), .B2(n20912), .A(n13359), .ZN(n13360) );
  OAI211_X1 U16637 ( .C1(n15254), .C2(n13362), .A(n13361), .B(n13360), .ZN(
        P1_U3153) );
  INV_X1 U16638 ( .A(n13363), .ZN(n19787) );
  OAI211_X1 U16639 ( .C1(n19787), .C2(n12216), .A(n19793), .B(n19779), .ZN(
        n13367) );
  AOI21_X1 U16640 ( .B1(n13365), .B2(n14050), .A(n15884), .ZN(n19691) );
  NAND2_X1 U16641 ( .A1(n19691), .A2(n19784), .ZN(n13366) );
  OAI211_X1 U16642 ( .C1(n19784), .C2(n10351), .A(n13367), .B(n13366), .ZN(
        P2_U2878) );
  AOI21_X1 U16643 ( .B1(n13370), .B2(n13369), .A(n13368), .ZN(n20590) );
  XNOR2_X1 U16644 ( .A(n20054), .B(n20590), .ZN(n13377) );
  XNOR2_X1 U16645 ( .A(n13372), .B(n13371), .ZN(n20603) );
  INV_X1 U16646 ( .A(n20603), .ZN(n13373) );
  NAND2_X1 U16647 ( .A1(n16223), .A2(n13373), .ZN(n13374) );
  OAI21_X1 U16648 ( .B1(n16223), .B2(n13373), .A(n13374), .ZN(n19861) );
  NOR2_X1 U16649 ( .A1(n19861), .A2(n19862), .ZN(n19860) );
  INV_X1 U16650 ( .A(n13374), .ZN(n13375) );
  NOR2_X1 U16651 ( .A1(n19860), .A2(n13375), .ZN(n13376) );
  NOR2_X1 U16652 ( .A1(n13376), .A2(n13377), .ZN(n19838) );
  AOI21_X1 U16653 ( .B1(n13377), .B2(n13376), .A(n19838), .ZN(n13381) );
  AOI22_X1 U16654 ( .A1(n19836), .A2(n16928), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19858), .ZN(n13380) );
  INV_X1 U16655 ( .A(n20590), .ZN(n13378) );
  NAND2_X1 U16656 ( .A1(n13378), .A2(n19859), .ZN(n13379) );
  OAI211_X1 U16657 ( .C1(n13381), .C2(n19863), .A(n13380), .B(n13379), .ZN(
        P2_U2917) );
  INV_X1 U16658 ( .A(n20893), .ZN(n15157) );
  NOR3_X1 U16659 ( .A1(n16513), .A2(n13870), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13384) );
  NAND2_X1 U16660 ( .A1(n13662), .A2(n13651), .ZN(n13387) );
  INV_X1 U16661 ( .A(n13653), .ZN(n13382) );
  INV_X1 U16662 ( .A(n13384), .ZN(n20901) );
  NOR2_X1 U16663 ( .A1(n20864), .A2(n20901), .ZN(n13410) );
  AOI21_X1 U16664 ( .B1(n20897), .B2(n13382), .A(n13410), .ZN(n13386) );
  OAI211_X1 U16665 ( .C1(n13387), .C2(n20640), .A(n13770), .B(n13386), .ZN(
        n13383) );
  OAI211_X1 U16666 ( .C1(n15157), .C2(n13384), .A(n13383), .B(n13536), .ZN(
        n13385) );
  INV_X1 U16667 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13390) );
  OAI22_X1 U16668 ( .A1(n13386), .A2(n20893), .B1(n20901), .B2(n13658), .ZN(
        n13409) );
  AOI22_X1 U16669 ( .A1(n20902), .A2(n13410), .B1(n13660), .B2(n13409), .ZN(
        n13389) );
  AOI22_X1 U16670 ( .A1(n13906), .A2(n20903), .B1(n10195), .B2(n20912), .ZN(
        n13388) );
  OAI211_X1 U16671 ( .C1(n13414), .C2(n13390), .A(n13389), .B(n13388), .ZN(
        P1_U3137) );
  INV_X1 U16672 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13393) );
  AOI22_X1 U16673 ( .A1(n20922), .A2(n13410), .B1(n13682), .B2(n13409), .ZN(
        n13392) );
  AOI22_X1 U16674 ( .A1(n13906), .A2(n20923), .B1(n10195), .B2(n20924), .ZN(
        n13391) );
  OAI211_X1 U16675 ( .C1(n13414), .C2(n13393), .A(n13392), .B(n13391), .ZN(
        P1_U3139) );
  INV_X1 U16676 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13396) );
  AOI22_X1 U16677 ( .A1(n20916), .A2(n13410), .B1(n13678), .B2(n13409), .ZN(
        n13395) );
  AOI22_X1 U16678 ( .A1(n13906), .A2(n20917), .B1(n10195), .B2(n20918), .ZN(
        n13394) );
  OAI211_X1 U16679 ( .C1(n13414), .C2(n13396), .A(n13395), .B(n13394), .ZN(
        P1_U3138) );
  INV_X1 U16680 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13399) );
  AOI22_X1 U16681 ( .A1(n20952), .A2(n13410), .B1(n13898), .B2(n13409), .ZN(
        n13398) );
  INV_X1 U16682 ( .A(n15236), .ZN(n20955) );
  AOI22_X1 U16683 ( .A1(n13906), .A2(n20954), .B1(n10195), .B2(n20955), .ZN(
        n13397) );
  OAI211_X1 U16684 ( .C1(n13414), .C2(n13399), .A(n13398), .B(n13397), .ZN(
        P1_U3144) );
  AOI22_X1 U16685 ( .A1(n20946), .A2(n13410), .B1(n13905), .B2(n13409), .ZN(
        n13401) );
  INV_X1 U16686 ( .A(n15230), .ZN(n20948) );
  AOI22_X1 U16687 ( .A1(n13906), .A2(n20947), .B1(n10195), .B2(n20948), .ZN(
        n13400) );
  OAI211_X1 U16688 ( .C1(n13414), .C2(n13402), .A(n13401), .B(n13400), .ZN(
        P1_U3143) );
  INV_X1 U16689 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13405) );
  AOI22_X1 U16690 ( .A1(n20940), .A2(n13410), .B1(n13691), .B2(n13409), .ZN(
        n13404) );
  AOI22_X1 U16691 ( .A1(n13906), .A2(n20941), .B1(n10195), .B2(n20942), .ZN(
        n13403) );
  OAI211_X1 U16692 ( .C1(n13414), .C2(n13405), .A(n13404), .B(n13403), .ZN(
        P1_U3142) );
  INV_X1 U16693 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13408) );
  AOI22_X1 U16694 ( .A1(n20934), .A2(n13410), .B1(n13668), .B2(n13409), .ZN(
        n13407) );
  AOI22_X1 U16695 ( .A1(n13906), .A2(n20935), .B1(n10195), .B2(n20936), .ZN(
        n13406) );
  OAI211_X1 U16696 ( .C1(n13414), .C2(n13408), .A(n13407), .B(n13406), .ZN(
        P1_U3141) );
  INV_X1 U16697 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U16698 ( .A1(n20928), .A2(n13410), .B1(n13686), .B2(n13409), .ZN(
        n13412) );
  AOI22_X1 U16699 ( .A1(n13906), .A2(n20929), .B1(n10195), .B2(n20930), .ZN(
        n13411) );
  OAI211_X1 U16700 ( .C1(n13414), .C2(n13413), .A(n13412), .B(n13411), .ZN(
        P1_U3140) );
  INV_X1 U16701 ( .A(n15165), .ZN(n13417) );
  INV_X1 U16702 ( .A(n13651), .ZN(n13661) );
  AOI21_X1 U16703 ( .B1(n13417), .B2(n13423), .A(n15248), .ZN(n13418) );
  INV_X1 U16704 ( .A(n13536), .ZN(n13656) );
  INV_X1 U16705 ( .A(n13419), .ZN(n13445) );
  OR2_X1 U16706 ( .A1(n15162), .A2(n13420), .ZN(n15245) );
  INV_X1 U16707 ( .A(n15245), .ZN(n13772) );
  AOI21_X1 U16708 ( .B1(n13772), .B2(n13534), .A(n13445), .ZN(n13422) );
  OAI22_X1 U16709 ( .A1(n13422), .A2(n20893), .B1(n13421), .B2(n13658), .ZN(
        n13444) );
  AOI22_X1 U16710 ( .A1(n20946), .A2(n13445), .B1(n13905), .B2(n13444), .ZN(
        n13425) );
  NAND2_X1 U16711 ( .A1(n13423), .A2(n9606), .ZN(n15290) );
  AOI22_X1 U16712 ( .A1(n13446), .A2(n20948), .B1(n13637), .B2(n20947), .ZN(
        n13424) );
  OAI211_X1 U16713 ( .C1(n13450), .C2(n13426), .A(n13425), .B(n13424), .ZN(
        P1_U3095) );
  AOI22_X1 U16714 ( .A1(n20916), .A2(n13445), .B1(n13678), .B2(n13444), .ZN(
        n13428) );
  AOI22_X1 U16715 ( .A1(n13446), .A2(n20918), .B1(n13637), .B2(n20917), .ZN(
        n13427) );
  OAI211_X1 U16716 ( .C1(n13450), .C2(n13429), .A(n13428), .B(n13427), .ZN(
        P1_U3090) );
  AOI22_X1 U16717 ( .A1(n20952), .A2(n13445), .B1(n13898), .B2(n13444), .ZN(
        n13431) );
  AOI22_X1 U16718 ( .A1(n13446), .A2(n20955), .B1(n13637), .B2(n20954), .ZN(
        n13430) );
  OAI211_X1 U16719 ( .C1(n13450), .C2(n13432), .A(n13431), .B(n13430), .ZN(
        P1_U3096) );
  AOI22_X1 U16720 ( .A1(n20934), .A2(n13445), .B1(n13668), .B2(n13444), .ZN(
        n13434) );
  AOI22_X1 U16721 ( .A1(n13446), .A2(n20936), .B1(n13637), .B2(n20935), .ZN(
        n13433) );
  OAI211_X1 U16722 ( .C1(n13450), .C2(n13435), .A(n13434), .B(n13433), .ZN(
        P1_U3093) );
  AOI22_X1 U16723 ( .A1(n20928), .A2(n13445), .B1(n13686), .B2(n13444), .ZN(
        n13437) );
  AOI22_X1 U16724 ( .A1(n13446), .A2(n20930), .B1(n13637), .B2(n20929), .ZN(
        n13436) );
  OAI211_X1 U16725 ( .C1(n13450), .C2(n13438), .A(n13437), .B(n13436), .ZN(
        P1_U3092) );
  AOI22_X1 U16726 ( .A1(n20940), .A2(n13445), .B1(n13691), .B2(n13444), .ZN(
        n13440) );
  AOI22_X1 U16727 ( .A1(n13446), .A2(n20942), .B1(n13637), .B2(n20941), .ZN(
        n13439) );
  OAI211_X1 U16728 ( .C1(n13450), .C2(n10994), .A(n13440), .B(n13439), .ZN(
        P1_U3094) );
  AOI22_X1 U16729 ( .A1(n20902), .A2(n13445), .B1(n13660), .B2(n13444), .ZN(
        n13442) );
  AOI22_X1 U16730 ( .A1(n13446), .A2(n20912), .B1(n13637), .B2(n20903), .ZN(
        n13441) );
  OAI211_X1 U16731 ( .C1(n13450), .C2(n13443), .A(n13442), .B(n13441), .ZN(
        P1_U3089) );
  AOI22_X1 U16732 ( .A1(n20922), .A2(n13445), .B1(n13682), .B2(n13444), .ZN(
        n13448) );
  AOI22_X1 U16733 ( .A1(n13446), .A2(n20924), .B1(n13637), .B2(n20923), .ZN(
        n13447) );
  OAI211_X1 U16734 ( .C1(n13450), .C2(n13449), .A(n13448), .B(n13447), .ZN(
        P1_U3091) );
  NOR3_X2 U16735 ( .A1(n13535), .A2(n15158), .A3(n13663), .ZN(n13642) );
  AND2_X1 U16736 ( .A1(n13531), .A2(n13663), .ZN(n13451) );
  AND2_X1 U16737 ( .A1(n13150), .A2(n15162), .ZN(n20859) );
  INV_X1 U16738 ( .A(n20859), .ZN(n13453) );
  NOR3_X1 U16739 ( .A1(n13870), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13458) );
  INV_X1 U16740 ( .A(n13458), .ZN(n13602) );
  OR2_X1 U16741 ( .A1(n20864), .A2(n13602), .ZN(n13479) );
  OAI21_X1 U16742 ( .B1(n13453), .B2(n13653), .A(n13479), .ZN(n13455) );
  AOI22_X1 U16743 ( .A1(n13455), .A2(n15157), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13458), .ZN(n13480) );
  OAI22_X1 U16744 ( .A1(n13480), .A2(n20945), .B1(n15279), .B2(n13479), .ZN(
        n13454) );
  AOI21_X1 U16745 ( .B1(n20887), .B2(n20941), .A(n13454), .ZN(n13460) );
  INV_X1 U16746 ( .A(n13455), .ZN(n13456) );
  OAI211_X1 U16747 ( .C1(n13535), .C2(n20640), .A(n13770), .B(n13456), .ZN(
        n13457) );
  OAI211_X1 U16748 ( .C1(n13770), .C2(n13458), .A(n13457), .B(n13536), .ZN(
        n13482) );
  NAND2_X1 U16749 ( .A1(n13482), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n13459) );
  OAI211_X1 U16750 ( .C1(n13485), .C2(n15225), .A(n13460), .B(n13459), .ZN(
        P1_U3110) );
  OAI22_X1 U16751 ( .A1(n20960), .A2(n13480), .B1(n15292), .B2(n13479), .ZN(
        n13461) );
  AOI21_X1 U16752 ( .B1(n20887), .B2(n20954), .A(n13461), .ZN(n13463) );
  NAND2_X1 U16753 ( .A1(n13482), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n13462) );
  OAI211_X1 U16754 ( .C1(n13485), .C2(n15236), .A(n13463), .B(n13462), .ZN(
        P1_U3112) );
  OAI22_X1 U16755 ( .A1(n13480), .A2(n20939), .B1(n15274), .B2(n13479), .ZN(
        n13464) );
  AOI21_X1 U16756 ( .B1(n20887), .B2(n20935), .A(n13464), .ZN(n13466) );
  NAND2_X1 U16757 ( .A1(n13482), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n13465) );
  OAI211_X1 U16758 ( .C1(n13485), .C2(n15220), .A(n13466), .B(n13465), .ZN(
        P1_U3109) );
  OAI22_X1 U16759 ( .A1(n13480), .A2(n20933), .B1(n15269), .B2(n13479), .ZN(
        n13467) );
  AOI21_X1 U16760 ( .B1(n20887), .B2(n20929), .A(n13467), .ZN(n13469) );
  NAND2_X1 U16761 ( .A1(n13482), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n13468) );
  OAI211_X1 U16762 ( .C1(n13485), .C2(n15215), .A(n13469), .B(n13468), .ZN(
        P1_U3108) );
  OAI22_X1 U16763 ( .A1(n13480), .A2(n20927), .B1(n15264), .B2(n13479), .ZN(
        n13470) );
  AOI21_X1 U16764 ( .B1(n20887), .B2(n20923), .A(n13470), .ZN(n13472) );
  NAND2_X1 U16765 ( .A1(n13482), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13471) );
  OAI211_X1 U16766 ( .C1(n13485), .C2(n15211), .A(n13472), .B(n13471), .ZN(
        P1_U3107) );
  OAI22_X1 U16767 ( .A1(n13480), .A2(n20921), .B1(n15259), .B2(n13479), .ZN(
        n13473) );
  AOI21_X1 U16768 ( .B1(n20887), .B2(n20917), .A(n13473), .ZN(n13475) );
  NAND2_X1 U16769 ( .A1(n13482), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13474) );
  OAI211_X1 U16770 ( .C1(n13485), .C2(n15206), .A(n13475), .B(n13474), .ZN(
        P1_U3106) );
  OAI22_X1 U16771 ( .A1(n13480), .A2(n20915), .B1(n15254), .B2(n13479), .ZN(
        n13476) );
  AOI21_X1 U16772 ( .B1(n20887), .B2(n20903), .A(n13476), .ZN(n13478) );
  NAND2_X1 U16773 ( .A1(n13482), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13477) );
  OAI211_X1 U16774 ( .C1(n13485), .C2(n15201), .A(n13478), .B(n13477), .ZN(
        P1_U3105) );
  OAI22_X1 U16775 ( .A1(n20951), .A2(n13480), .B1(n15284), .B2(n13479), .ZN(
        n13481) );
  AOI21_X1 U16776 ( .B1(n20887), .B2(n20947), .A(n13481), .ZN(n13484) );
  NAND2_X1 U16777 ( .A1(n13482), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13483) );
  OAI211_X1 U16778 ( .C1(n13485), .C2(n15230), .A(n13484), .B(n13483), .ZN(
        P1_U3111) );
  NOR2_X1 U16779 ( .A1(n13486), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20824) );
  INV_X1 U16780 ( .A(n20824), .ZN(n13487) );
  NAND3_X1 U16781 ( .A1(n13487), .A2(n20792), .A3(n20832), .ZN(n13491) );
  INV_X2 U16782 ( .A(n16817), .ZN(n21060) );
  AOI22_X1 U16783 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13488) );
  OAI21_X1 U16784 ( .B1(n16695), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13488), .ZN(n13489) );
  INV_X1 U16785 ( .A(n13489), .ZN(n13490) );
  OAI211_X1 U16786 ( .C1(n21063), .C2(n13601), .A(n13491), .B(n13490), .ZN(
        P1_U2998) );
  INV_X1 U16787 ( .A(n13492), .ZN(n13493) );
  XNOR2_X1 U16788 ( .A(n13279), .B(n13493), .ZN(n20790) );
  INV_X1 U16789 ( .A(n20790), .ZN(n13495) );
  INV_X1 U16790 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20740) );
  OAI222_X1 U16791 ( .A1(n14805), .A2(n13495), .B1(n14802), .B2(n20740), .C1(
        n13494), .C2(n14804), .ZN(P1_U2900) );
  NAND2_X1 U16792 ( .A1(n12060), .A2(n15158), .ZN(n13496) );
  INV_X1 U16793 ( .A(n15191), .ZN(n13497) );
  NOR2_X1 U16794 ( .A1(n13533), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13521) );
  AOI21_X1 U16795 ( .B1(n13497), .B2(n13534), .A(n13521), .ZN(n13503) );
  INV_X1 U16796 ( .A(n15161), .ZN(n13498) );
  AND2_X1 U16797 ( .A1(n13499), .A2(n15157), .ZN(n13501) );
  NAND3_X1 U16798 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n13870), .A3(
        n16513), .ZN(n13789) );
  AOI22_X1 U16799 ( .A1(n13503), .A2(n13501), .B1(n20893), .B2(n13789), .ZN(
        n13500) );
  NAND2_X1 U16800 ( .A1(n13536), .A2(n13500), .ZN(n13520) );
  INV_X1 U16801 ( .A(n13501), .ZN(n13502) );
  OAI22_X1 U16802 ( .A1(n13503), .A2(n13502), .B1(n13658), .B2(n13789), .ZN(
        n13519) );
  AOI22_X1 U16803 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13520), .B1(
        n13668), .B2(n13519), .ZN(n13506) );
  NAND2_X1 U16804 ( .A1(n13504), .A2(n9606), .ZN(n13817) );
  AOI22_X1 U16805 ( .A1(n13522), .A2(n20936), .B1(n20934), .B2(n13521), .ZN(
        n13505) );
  OAI211_X1 U16806 ( .C1(n15273), .C2(n13846), .A(n13506), .B(n13505), .ZN(
        P1_U3061) );
  AOI22_X1 U16807 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13520), .B1(
        n13686), .B2(n13519), .ZN(n13508) );
  AOI22_X1 U16808 ( .A1(n13522), .A2(n20930), .B1(n20928), .B2(n13521), .ZN(
        n13507) );
  OAI211_X1 U16809 ( .C1(n15268), .C2(n13846), .A(n13508), .B(n13507), .ZN(
        P1_U3060) );
  AOI22_X1 U16810 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13520), .B1(
        n13682), .B2(n13519), .ZN(n13510) );
  AOI22_X1 U16811 ( .A1(n13522), .A2(n20924), .B1(n20922), .B2(n13521), .ZN(
        n13509) );
  OAI211_X1 U16812 ( .C1(n15263), .C2(n13846), .A(n13510), .B(n13509), .ZN(
        P1_U3059) );
  AOI22_X1 U16813 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13520), .B1(
        n13678), .B2(n13519), .ZN(n13512) );
  AOI22_X1 U16814 ( .A1(n13522), .A2(n20918), .B1(n20916), .B2(n13521), .ZN(
        n13511) );
  OAI211_X1 U16815 ( .C1(n15258), .C2(n13846), .A(n13512), .B(n13511), .ZN(
        P1_U3058) );
  AOI22_X1 U16816 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13520), .B1(
        n13660), .B2(n13519), .ZN(n13514) );
  AOI22_X1 U16817 ( .A1(n13522), .A2(n20912), .B1(n20902), .B2(n13521), .ZN(
        n13513) );
  OAI211_X1 U16818 ( .C1(n15253), .C2(n13846), .A(n13514), .B(n13513), .ZN(
        P1_U3057) );
  AOI22_X1 U16819 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n13520), .B1(
        n13691), .B2(n13519), .ZN(n13516) );
  AOI22_X1 U16820 ( .A1(n13522), .A2(n20942), .B1(n20940), .B2(n13521), .ZN(
        n13515) );
  OAI211_X1 U16821 ( .C1(n15278), .C2(n13846), .A(n13516), .B(n13515), .ZN(
        P1_U3062) );
  AOI22_X1 U16822 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13520), .B1(
        n13905), .B2(n13519), .ZN(n13518) );
  AOI22_X1 U16823 ( .A1(n13522), .A2(n20948), .B1(n20946), .B2(n13521), .ZN(
        n13517) );
  OAI211_X1 U16824 ( .C1(n15283), .C2(n13846), .A(n13518), .B(n13517), .ZN(
        P1_U3063) );
  AOI22_X1 U16825 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13520), .B1(
        n13898), .B2(n13519), .ZN(n13524) );
  AOI22_X1 U16826 ( .A1(n13522), .A2(n20955), .B1(n20952), .B2(n13521), .ZN(
        n13523) );
  OAI211_X1 U16827 ( .C1(n15289), .C2(n13846), .A(n13524), .B(n13523), .ZN(
        P1_U3064) );
  OR2_X1 U16828 ( .A1(n13527), .A2(n13526), .ZN(n13528) );
  AND2_X1 U16829 ( .A1(n13525), .A2(n13528), .ZN(n20714) );
  INV_X1 U16830 ( .A(n20714), .ZN(n13530) );
  INV_X1 U16831 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13529) );
  OAI222_X1 U16832 ( .A1(n13530), .A2(n14805), .B1(n14772), .B2(n14804), .C1(
        n13529), .C2(n14802), .ZN(P1_U2899) );
  NOR3_X1 U16833 ( .A1(n13870), .A2(n13532), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20863) );
  NOR2_X1 U16834 ( .A1(n13533), .A2(n13870), .ZN(n13557) );
  AOI21_X1 U16835 ( .B1(n20859), .B2(n13534), .A(n13557), .ZN(n13540) );
  OAI211_X1 U16836 ( .C1(n13535), .C2(n15161), .A(n13770), .B(n13540), .ZN(
        n13537) );
  OAI211_X1 U16837 ( .C1(n15157), .C2(n20863), .A(n13537), .B(n13536), .ZN(
        n13555) );
  AOI22_X1 U16838 ( .A1(n13555), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n20888), .B2(n20948), .ZN(n13542) );
  INV_X1 U16839 ( .A(n20863), .ZN(n13539) );
  OAI22_X1 U16840 ( .A1(n13540), .A2(n20893), .B1(n13539), .B2(n13658), .ZN(
        n13556) );
  AOI22_X1 U16841 ( .A1(n20946), .A2(n13557), .B1(n13905), .B2(n13556), .ZN(
        n13541) );
  OAI211_X1 U16842 ( .C1(n15283), .C2(n20911), .A(n13542), .B(n13541), .ZN(
        P1_U3127) );
  AOI22_X1 U16843 ( .A1(n13555), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n20888), .B2(n20912), .ZN(n13544) );
  AOI22_X1 U16844 ( .A1(n20902), .A2(n13557), .B1(n13660), .B2(n13556), .ZN(
        n13543) );
  OAI211_X1 U16845 ( .C1(n15253), .C2(n20911), .A(n13544), .B(n13543), .ZN(
        P1_U3121) );
  AOI22_X1 U16846 ( .A1(n13555), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n20888), .B2(n20942), .ZN(n13546) );
  AOI22_X1 U16847 ( .A1(n20940), .A2(n13557), .B1(n13691), .B2(n13556), .ZN(
        n13545) );
  OAI211_X1 U16848 ( .C1(n15278), .C2(n20911), .A(n13546), .B(n13545), .ZN(
        P1_U3126) );
  AOI22_X1 U16849 ( .A1(n13555), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n20888), .B2(n20924), .ZN(n13548) );
  AOI22_X1 U16850 ( .A1(n20922), .A2(n13557), .B1(n13682), .B2(n13556), .ZN(
        n13547) );
  OAI211_X1 U16851 ( .C1(n15263), .C2(n20911), .A(n13548), .B(n13547), .ZN(
        P1_U3123) );
  AOI22_X1 U16852 ( .A1(n13555), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n20888), .B2(n20918), .ZN(n13550) );
  AOI22_X1 U16853 ( .A1(n20916), .A2(n13557), .B1(n13678), .B2(n13556), .ZN(
        n13549) );
  OAI211_X1 U16854 ( .C1(n15258), .C2(n20911), .A(n13550), .B(n13549), .ZN(
        P1_U3122) );
  AOI22_X1 U16855 ( .A1(n13555), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n20888), .B2(n20955), .ZN(n13552) );
  AOI22_X1 U16856 ( .A1(n20952), .A2(n13557), .B1(n13898), .B2(n13556), .ZN(
        n13551) );
  OAI211_X1 U16857 ( .C1(n15289), .C2(n20911), .A(n13552), .B(n13551), .ZN(
        P1_U3128) );
  AOI22_X1 U16858 ( .A1(n13555), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n20888), .B2(n20930), .ZN(n13554) );
  AOI22_X1 U16859 ( .A1(n20928), .A2(n13557), .B1(n13686), .B2(n13556), .ZN(
        n13553) );
  OAI211_X1 U16860 ( .C1(n15268), .C2(n20911), .A(n13554), .B(n13553), .ZN(
        P1_U3124) );
  AOI22_X1 U16861 ( .A1(n13555), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n20888), .B2(n20936), .ZN(n13559) );
  AOI22_X1 U16862 ( .A1(n20934), .A2(n13557), .B1(n13668), .B2(n13556), .ZN(
        n13558) );
  OAI211_X1 U16863 ( .C1(n15273), .C2(n20911), .A(n13559), .B(n13558), .ZN(
        P1_U3125) );
  INV_X1 U16864 ( .A(n19774), .ZN(n13563) );
  OAI21_X1 U16865 ( .B1(n19779), .B2(n13561), .A(n13560), .ZN(n13562) );
  NAND3_X1 U16866 ( .A1(n13563), .A2(n19793), .A3(n13562), .ZN(n13568) );
  NAND2_X1 U16867 ( .A1(n13564), .A2(n15886), .ZN(n13566) );
  INV_X1 U16868 ( .A(n15496), .ZN(n13565) );
  NAND2_X1 U16869 ( .A1(n19784), .A2(n16938), .ZN(n13567) );
  OAI211_X1 U16870 ( .C1(n19784), .C2(n9920), .A(n13568), .B(n13567), .ZN(
        P2_U2876) );
  AND2_X1 U16871 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20963), .ZN(n13570) );
  NAND2_X1 U16872 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21054), .ZN(n16534) );
  INV_X1 U16873 ( .A(n16534), .ZN(n13569) );
  AOI22_X1 U16874 ( .A1(n13571), .A2(n13570), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n13569), .ZN(n13572) );
  AND2_X1 U16875 ( .A1(n16817), .A2(n13572), .ZN(n13573) );
  OR2_X1 U16876 ( .A1(n13579), .A2(n13576), .ZN(n13577) );
  NOR2_X1 U16877 ( .A1(n13579), .A2(n13578), .ZN(n20698) );
  INV_X1 U16878 ( .A(n20698), .ZN(n13598) );
  INV_X1 U16879 ( .A(n13594), .ZN(n13583) );
  NAND2_X1 U16880 ( .A1(n21051), .A2(n20640), .ZN(n13590) );
  INV_X1 U16881 ( .A(n13590), .ZN(n13580) );
  NAND2_X1 U16882 ( .A1(n14956), .A2(n13580), .ZN(n13593) );
  INV_X1 U16883 ( .A(n13593), .ZN(n13581) );
  INV_X1 U16884 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14668) );
  NOR2_X1 U16885 ( .A1(n13581), .A2(n13591), .ZN(n13582) );
  INV_X1 U16886 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21039) );
  NAND2_X1 U16887 ( .A1(n20705), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13588) );
  NOR2_X1 U16888 ( .A1(n13584), .A2(n20962), .ZN(n13585) );
  INV_X1 U16889 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13586) );
  NAND2_X1 U16890 ( .A1(n20687), .A2(n13586), .ZN(n13587) );
  OAI211_X1 U16891 ( .C1(n21039), .C2(n13928), .A(n13588), .B(n13587), .ZN(
        n13589) );
  AOI21_X1 U16892 ( .B1(n20684), .B2(P1_EBX_REG_1__SCAN_IN), .A(n13589), .ZN(
        n13597) );
  NAND2_X1 U16893 ( .A1(n13591), .A2(n13590), .ZN(n13592) );
  NOR2_X2 U16894 ( .A1(n13594), .A2(n13592), .ZN(n20700) );
  AOI22_X1 U16895 ( .A1(n20700), .A2(n13595), .B1(n13944), .B2(n21039), .ZN(
        n13596) );
  OAI211_X1 U16896 ( .C1(n20896), .C2(n13598), .A(n13597), .B(n13596), .ZN(
        n13599) );
  INV_X1 U16897 ( .A(n13599), .ZN(n13600) );
  OAI21_X1 U16898 ( .B1(n13601), .B2(n14655), .A(n13600), .ZN(P1_U2839) );
  OAI21_X1 U16899 ( .B1(n13642), .B2(n13637), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13604) );
  NOR2_X1 U16900 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13602), .ZN(
        n13638) );
  AOI21_X1 U16901 ( .B1(n20859), .B2(n20896), .A(n13638), .ZN(n13605) );
  AND2_X1 U16902 ( .A1(n13606), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20899) );
  OAI21_X1 U16903 ( .B1(n13638), .B2(n20905), .A(n20869), .ZN(n13603) );
  INV_X1 U16904 ( .A(n13605), .ZN(n13608) );
  NOR2_X1 U16905 ( .A1(n13606), .A2(n13658), .ZN(n20861) );
  INV_X1 U16906 ( .A(n13773), .ZN(n13607) );
  NAND2_X1 U16907 ( .A1(n13607), .A2(n13871), .ZN(n20907) );
  INV_X1 U16908 ( .A(n20907), .ZN(n20898) );
  AOI22_X1 U16909 ( .A1(n13608), .A2(n15157), .B1(n20861), .B2(n20898), .ZN(
        n13640) );
  AOI22_X1 U16910 ( .A1(n20934), .A2(n13638), .B1(n13637), .B2(n20936), .ZN(
        n13609) );
  OAI21_X1 U16911 ( .B1(n13640), .B2(n20939), .A(n13609), .ZN(n13610) );
  AOI21_X1 U16912 ( .B1(n13642), .B2(n20935), .A(n13610), .ZN(n13611) );
  OAI21_X1 U16913 ( .B1(n13645), .B2(n13612), .A(n13611), .ZN(P1_U3101) );
  AOI22_X1 U16914 ( .A1(n20940), .A2(n13638), .B1(n13637), .B2(n20942), .ZN(
        n13613) );
  OAI21_X1 U16915 ( .B1(n13640), .B2(n20945), .A(n13613), .ZN(n13614) );
  AOI21_X1 U16916 ( .B1(n13642), .B2(n20941), .A(n13614), .ZN(n13615) );
  OAI21_X1 U16917 ( .B1(n13645), .B2(n13616), .A(n13615), .ZN(P1_U3102) );
  AOI22_X1 U16918 ( .A1(n20946), .A2(n13638), .B1(n13637), .B2(n20948), .ZN(
        n13617) );
  OAI21_X1 U16919 ( .B1(n13640), .B2(n20951), .A(n13617), .ZN(n13618) );
  AOI21_X1 U16920 ( .B1(n13642), .B2(n20947), .A(n13618), .ZN(n13619) );
  OAI21_X1 U16921 ( .B1(n13645), .B2(n13620), .A(n13619), .ZN(P1_U3103) );
  AOI22_X1 U16922 ( .A1(n20952), .A2(n13638), .B1(n13637), .B2(n20955), .ZN(
        n13621) );
  OAI21_X1 U16923 ( .B1(n13640), .B2(n20960), .A(n13621), .ZN(n13622) );
  AOI21_X1 U16924 ( .B1(n13642), .B2(n20954), .A(n13622), .ZN(n13623) );
  OAI21_X1 U16925 ( .B1(n13645), .B2(n13624), .A(n13623), .ZN(P1_U3104) );
  AOI22_X1 U16926 ( .A1(n20916), .A2(n13638), .B1(n13637), .B2(n20918), .ZN(
        n13625) );
  OAI21_X1 U16927 ( .B1(n13640), .B2(n20921), .A(n13625), .ZN(n13626) );
  AOI21_X1 U16928 ( .B1(n13642), .B2(n20917), .A(n13626), .ZN(n13627) );
  OAI21_X1 U16929 ( .B1(n13645), .B2(n13628), .A(n13627), .ZN(P1_U3098) );
  AOI22_X1 U16930 ( .A1(n20902), .A2(n13638), .B1(n13637), .B2(n20912), .ZN(
        n13629) );
  OAI21_X1 U16931 ( .B1(n13640), .B2(n20915), .A(n13629), .ZN(n13630) );
  AOI21_X1 U16932 ( .B1(n13642), .B2(n20903), .A(n13630), .ZN(n13631) );
  OAI21_X1 U16933 ( .B1(n13645), .B2(n13632), .A(n13631), .ZN(P1_U3097) );
  AOI22_X1 U16934 ( .A1(n20922), .A2(n13638), .B1(n13637), .B2(n20924), .ZN(
        n13633) );
  OAI21_X1 U16935 ( .B1(n13640), .B2(n20927), .A(n13633), .ZN(n13634) );
  AOI21_X1 U16936 ( .B1(n13642), .B2(n20923), .A(n13634), .ZN(n13635) );
  OAI21_X1 U16937 ( .B1(n13645), .B2(n13636), .A(n13635), .ZN(P1_U3099) );
  AOI22_X1 U16938 ( .A1(n20928), .A2(n13638), .B1(n13637), .B2(n20930), .ZN(
        n13639) );
  OAI21_X1 U16939 ( .B1(n13640), .B2(n20933), .A(n13639), .ZN(n13641) );
  AOI21_X1 U16940 ( .B1(n13642), .B2(n20929), .A(n13641), .ZN(n13643) );
  OAI21_X1 U16941 ( .B1(n13645), .B2(n13644), .A(n13643), .ZN(P1_U3100) );
  INV_X1 U16942 ( .A(n13646), .ZN(n13647) );
  AOI21_X1 U16943 ( .B1(n13648), .B2(n13525), .A(n13647), .ZN(n20677) );
  INV_X1 U16944 ( .A(n20677), .ZN(n13698) );
  XOR2_X1 U16945 ( .A(n13649), .B(n16831), .Z(n20671) );
  AOI22_X1 U16946 ( .A1(n20671), .A2(n20717), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14715), .ZN(n13650) );
  OAI21_X1 U16947 ( .B1(n13698), .B2(n14731), .A(n13650), .ZN(P1_U2866) );
  OR3_X1 U16948 ( .A1(n16513), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13767) );
  NOR2_X1 U16949 ( .A1(n13651), .A2(n20640), .ZN(n13654) );
  NOR2_X1 U16950 ( .A1(n20864), .A2(n13767), .ZN(n13692) );
  INV_X1 U16951 ( .A(n13692), .ZN(n13652) );
  OAI21_X1 U16952 ( .B1(n15245), .B2(n13653), .A(n13652), .ZN(n13657) );
  AOI211_X1 U16953 ( .C1(n13662), .C2(n13654), .A(n20893), .B(n13657), .ZN(
        n13655) );
  AOI211_X2 U16954 ( .C1(n20893), .C2(n13767), .A(n13656), .B(n13655), .ZN(
        n13696) );
  INV_X1 U16955 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13667) );
  INV_X1 U16956 ( .A(n13657), .ZN(n13659) );
  OAI22_X1 U16957 ( .A1(n13659), .A2(n20893), .B1(n13767), .B2(n13658), .ZN(
        n13690) );
  AOI22_X1 U16958 ( .A1(n20902), .A2(n13692), .B1(n13660), .B2(n13690), .ZN(
        n13666) );
  NAND2_X1 U16959 ( .A1(n13662), .A2(n13661), .ZN(n13664) );
  NOR2_X2 U16960 ( .A1(n13664), .A2(n9606), .ZN(n15294) );
  OR2_X1 U16961 ( .A1(n13664), .A2(n13663), .ZN(n13781) );
  AOI22_X1 U16962 ( .A1(n15294), .A2(n20903), .B1(n13843), .B2(n20912), .ZN(
        n13665) );
  OAI211_X1 U16963 ( .C1(n13696), .C2(n13667), .A(n13666), .B(n13665), .ZN(
        P1_U3073) );
  INV_X1 U16964 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13671) );
  AOI22_X1 U16965 ( .A1(n20934), .A2(n13692), .B1(n13668), .B2(n13690), .ZN(
        n13670) );
  AOI22_X1 U16966 ( .A1(n15294), .A2(n20935), .B1(n13843), .B2(n20936), .ZN(
        n13669) );
  OAI211_X1 U16967 ( .C1(n13696), .C2(n13671), .A(n13670), .B(n13669), .ZN(
        P1_U3077) );
  INV_X1 U16968 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U16969 ( .A1(n20952), .A2(n13692), .B1(n13898), .B2(n13690), .ZN(
        n13673) );
  AOI22_X1 U16970 ( .A1(n15294), .A2(n20954), .B1(n13843), .B2(n20955), .ZN(
        n13672) );
  OAI211_X1 U16971 ( .C1(n13696), .C2(n13674), .A(n13673), .B(n13672), .ZN(
        P1_U3080) );
  INV_X1 U16972 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U16973 ( .A1(n20946), .A2(n13692), .B1(n13905), .B2(n13690), .ZN(
        n13676) );
  AOI22_X1 U16974 ( .A1(n15294), .A2(n20947), .B1(n13843), .B2(n20948), .ZN(
        n13675) );
  OAI211_X1 U16975 ( .C1(n13696), .C2(n13677), .A(n13676), .B(n13675), .ZN(
        P1_U3079) );
  INV_X1 U16976 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13681) );
  AOI22_X1 U16977 ( .A1(n20916), .A2(n13692), .B1(n13678), .B2(n13690), .ZN(
        n13680) );
  AOI22_X1 U16978 ( .A1(n15294), .A2(n20917), .B1(n13843), .B2(n20918), .ZN(
        n13679) );
  OAI211_X1 U16979 ( .C1(n13696), .C2(n13681), .A(n13680), .B(n13679), .ZN(
        P1_U3074) );
  AOI22_X1 U16980 ( .A1(n20922), .A2(n13692), .B1(n13682), .B2(n13690), .ZN(
        n13684) );
  AOI22_X1 U16981 ( .A1(n15294), .A2(n20923), .B1(n13843), .B2(n20924), .ZN(
        n13683) );
  OAI211_X1 U16982 ( .C1(n13696), .C2(n13685), .A(n13684), .B(n13683), .ZN(
        P1_U3075) );
  INV_X1 U16983 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13689) );
  AOI22_X1 U16984 ( .A1(n20928), .A2(n13692), .B1(n13686), .B2(n13690), .ZN(
        n13688) );
  AOI22_X1 U16985 ( .A1(n15294), .A2(n20929), .B1(n13843), .B2(n20930), .ZN(
        n13687) );
  OAI211_X1 U16986 ( .C1(n13696), .C2(n13689), .A(n13688), .B(n13687), .ZN(
        P1_U3076) );
  INV_X1 U16987 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13695) );
  AOI22_X1 U16988 ( .A1(n20940), .A2(n13692), .B1(n13691), .B2(n13690), .ZN(
        n13694) );
  AOI22_X1 U16989 ( .A1(n15294), .A2(n20941), .B1(n13843), .B2(n20942), .ZN(
        n13693) );
  OAI211_X1 U16990 ( .C1(n13696), .C2(n13695), .A(n13694), .B(n13693), .ZN(
        P1_U3078) );
  OAI222_X1 U16991 ( .A1(n14805), .A2(n13698), .B1(n13697), .B2(n14804), .C1(
        n14802), .C2(n11370), .ZN(P1_U2898) );
  AOI22_X1 U16992 ( .A1(n13699), .A2(n20698), .B1(n20700), .B2(n20848), .ZN(
        n13704) );
  AOI21_X1 U16993 ( .B1(n16596), .B2(n20703), .A(n13700), .ZN(n13702) );
  INV_X1 U16994 ( .A(n13928), .ZN(n13952) );
  NOR2_X1 U16995 ( .A1(n16587), .A2(n13096), .ZN(n13701) );
  AOI211_X1 U16996 ( .C1(n20684), .C2(P1_EBX_REG_0__SCAN_IN), .A(n13702), .B(
        n13701), .ZN(n13703) );
  OAI211_X1 U16997 ( .C1(n13705), .C2(n14655), .A(n13704), .B(n13703), .ZN(
        P1_U2840) );
  NAND3_X1 U16998 ( .A1(n13707), .A2(n13706), .A3(n13728), .ZN(n13715) );
  INV_X1 U16999 ( .A(n13707), .ZN(n13710) );
  AOI21_X1 U17000 ( .B1(n13708), .B2(n10451), .A(n10435), .ZN(n13709) );
  NAND2_X1 U17001 ( .A1(n13710), .A2(n13709), .ZN(n13714) );
  NOR2_X1 U17002 ( .A1(n13712), .A2(n13711), .ZN(n13713) );
  NAND3_X1 U17003 ( .A1(n13715), .A2(n13714), .A3(n13713), .ZN(n13716) );
  NAND2_X1 U17004 ( .A1(n13716), .A2(n17073), .ZN(n13720) );
  MUX2_X1 U17005 ( .A(n10442), .B(n13728), .S(n17076), .Z(n13717) );
  NAND2_X1 U17006 ( .A1(n13718), .A2(n13717), .ZN(n13719) );
  NOR2_X1 U17007 ( .A1(n17046), .A2(n13721), .ZN(n20620) );
  XNOR2_X1 U17008 ( .A(n13722), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13723) );
  XNOR2_X1 U17009 ( .A(n13724), .B(n13723), .ZN(n13764) );
  XOR2_X1 U17010 ( .A(n13725), .B(n13726), .Z(n13762) );
  INV_X1 U17011 ( .A(n13727), .ZN(n20621) );
  INV_X1 U17012 ( .A(n14487), .ZN(n17051) );
  NAND2_X1 U17013 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16208) );
  NAND2_X1 U17014 ( .A1(n19925), .A2(n16208), .ZN(n19919) );
  INV_X1 U17015 ( .A(n19919), .ZN(n13741) );
  NAND2_X1 U17016 ( .A1(n13738), .A2(n10435), .ZN(n13729) );
  AOI22_X1 U17017 ( .A1(n15299), .A2(n13729), .B1(n19936), .B2(n13728), .ZN(
        n13730) );
  AND2_X1 U17018 ( .A1(n13731), .A2(n13730), .ZN(n13737) );
  OR2_X1 U17019 ( .A1(n13732), .A2(n17076), .ZN(n14086) );
  NAND2_X1 U17020 ( .A1(n14086), .A2(n13733), .ZN(n13735) );
  AOI21_X1 U17021 ( .B1(n13735), .B2(n19946), .A(n13734), .ZN(n13736) );
  OAI211_X1 U17022 ( .C1(n13739), .C2(n13738), .A(n13737), .B(n13736), .ZN(
        n17032) );
  INV_X1 U17023 ( .A(n17032), .ZN(n16216) );
  NAND2_X1 U17024 ( .A1(n16216), .A2(n12772), .ZN(n13740) );
  NAND2_X1 U17025 ( .A1(n13750), .A2(n13740), .ZN(n19935) );
  INV_X1 U17026 ( .A(n19935), .ZN(n13754) );
  OR2_X1 U17027 ( .A1(n19925), .A2(n16208), .ZN(n19918) );
  AOI22_X1 U17028 ( .A1(n19932), .A2(n13741), .B1(n13754), .B2(n19918), .ZN(
        n13742) );
  NOR2_X1 U17029 ( .A1(n13750), .A2(n19903), .ZN(n17011) );
  INV_X1 U17030 ( .A(n17011), .ZN(n19924) );
  NAND2_X1 U17031 ( .A1(n13742), .A2(n19924), .ZN(n14022) );
  NAND2_X1 U17032 ( .A1(n14022), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13753) );
  OR2_X1 U17033 ( .A1(n13744), .A2(n13743), .ZN(n13745) );
  NAND2_X1 U17034 ( .A1(n13745), .A2(n19739), .ZN(n19839) );
  INV_X1 U17035 ( .A(n19839), .ZN(n20584) );
  INV_X1 U17036 ( .A(n13746), .ZN(n17054) );
  OAI21_X1 U17037 ( .B1(n17076), .B2(n12630), .A(n17054), .ZN(n13747) );
  NAND2_X1 U17038 ( .A1(n17033), .A2(n17076), .ZN(n13748) );
  NAND2_X1 U17039 ( .A1(n13748), .A2(n14484), .ZN(n13749) );
  NAND2_X1 U17040 ( .A1(n19903), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13758) );
  OAI21_X1 U17041 ( .B1(n19911), .B2(n14113), .A(n13758), .ZN(n13751) );
  AOI21_X1 U17042 ( .B1(n20584), .B2(n19909), .A(n13751), .ZN(n13752) );
  NAND2_X1 U17043 ( .A1(n13753), .A2(n13752), .ZN(n13756) );
  NAND2_X1 U17044 ( .A1(n19932), .A2(n19919), .ZN(n14019) );
  AOI211_X1 U17045 ( .C1(n14019), .C2(n19918), .A(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n17022), .ZN(n13755) );
  AOI211_X1 U17046 ( .C1(n13762), .C2(n17013), .A(n13756), .B(n13755), .ZN(
        n13757) );
  OAI21_X1 U17047 ( .B1(n17009), .B2(n13764), .A(n13757), .ZN(P2_U3043) );
  INV_X1 U17048 ( .A(n14120), .ZN(n14115) );
  INV_X1 U17049 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14108) );
  OAI21_X1 U17050 ( .B1(n16950), .B2(n14108), .A(n13758), .ZN(n13759) );
  AOI21_X1 U17051 ( .B1(n16942), .B2(n14115), .A(n13759), .ZN(n13760) );
  OAI21_X1 U17052 ( .B1(n14113), .B2(n13859), .A(n13760), .ZN(n13761) );
  AOI21_X1 U17053 ( .B1(n13762), .B2(n15933), .A(n13761), .ZN(n13763) );
  OAI21_X1 U17054 ( .B1(n16957), .B2(n13764), .A(n13763), .ZN(P2_U3011) );
  AOI21_X1 U17055 ( .B1(n13846), .B2(n13781), .A(n20640), .ZN(n13765) );
  AOI21_X1 U17056 ( .B1(n13772), .B2(n20896), .A(n13765), .ZN(n13766) );
  NOR2_X1 U17057 ( .A1(n13766), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13769) );
  NOR2_X1 U17058 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13767), .ZN(
        n13823) );
  AND2_X1 U17059 ( .A1(n20896), .A2(n13770), .ZN(n13771) );
  NAND2_X1 U17060 ( .A1(n13772), .A2(n13771), .ZN(n13775) );
  AND2_X1 U17061 ( .A1(n13773), .A2(n13871), .ZN(n15198) );
  NAND2_X1 U17062 ( .A1(n20899), .A2(n15198), .ZN(n13774) );
  INV_X1 U17063 ( .A(n13840), .ZN(n13780) );
  AOI22_X1 U17064 ( .A1(n20946), .A2(n13823), .B1(n13905), .B2(n13780), .ZN(
        n13777) );
  OR2_X1 U17065 ( .A1(n13781), .A2(n15283), .ZN(n13776) );
  OAI211_X1 U17066 ( .C1(n15230), .C2(n13846), .A(n13777), .B(n13776), .ZN(
        n13778) );
  AOI21_X1 U17067 ( .B1(n13839), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n13778), .ZN(n13779) );
  INV_X1 U17068 ( .A(n13779), .ZN(P1_U3071) );
  AOI22_X1 U17069 ( .A1(n20952), .A2(n13823), .B1(n13898), .B2(n13780), .ZN(
        n13783) );
  OR2_X1 U17070 ( .A1(n13781), .A2(n15289), .ZN(n13782) );
  OAI211_X1 U17071 ( .C1(n15236), .C2(n13846), .A(n13783), .B(n13782), .ZN(
        n13784) );
  AOI21_X1 U17072 ( .B1(n13839), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n13784), .ZN(n13785) );
  INV_X1 U17073 ( .A(n13785), .ZN(P1_U3072) );
  NAND3_X1 U17074 ( .A1(n13786), .A2(n13817), .A3(n15157), .ZN(n13787) );
  NAND2_X1 U17075 ( .A1(n15157), .A2(n20640), .ZN(n20855) );
  NAND2_X1 U17076 ( .A1(n13787), .A2(n20855), .ZN(n13791) );
  NOR2_X1 U17077 ( .A1(n15191), .A2(n20896), .ZN(n13788) );
  OR2_X1 U17078 ( .A1(n13871), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13792) );
  INV_X1 U17079 ( .A(n13792), .ZN(n15246) );
  INV_X1 U17080 ( .A(n13788), .ZN(n13790) );
  OR2_X1 U17081 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13789), .ZN(
        n13816) );
  AOI22_X1 U17082 ( .A1(n13791), .A2(n13790), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n13816), .ZN(n13793) );
  NAND2_X1 U17083 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13792), .ZN(n15251) );
  NAND3_X1 U17084 ( .A1(n20869), .A2(n13793), .A3(n15251), .ZN(n13815) );
  NAND2_X1 U17085 ( .A1(n13815), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13796) );
  OAI22_X1 U17086 ( .A1(n13817), .A2(n15268), .B1(n13816), .B2(n15269), .ZN(
        n13794) );
  AOI21_X1 U17087 ( .B1(n13819), .B2(n20930), .A(n13794), .ZN(n13795) );
  OAI211_X1 U17088 ( .C1(n13822), .C2(n20933), .A(n13796), .B(n13795), .ZN(
        P1_U3052) );
  NAND2_X1 U17089 ( .A1(n13815), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13799) );
  OAI22_X1 U17090 ( .A1(n13817), .A2(n15273), .B1(n13816), .B2(n15274), .ZN(
        n13797) );
  AOI21_X1 U17091 ( .B1(n13819), .B2(n20936), .A(n13797), .ZN(n13798) );
  OAI211_X1 U17092 ( .C1(n13822), .C2(n20939), .A(n13799), .B(n13798), .ZN(
        P1_U3053) );
  NAND2_X1 U17093 ( .A1(n13815), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13802) );
  OAI22_X1 U17094 ( .A1(n13817), .A2(n15253), .B1(n15254), .B2(n13816), .ZN(
        n13800) );
  AOI21_X1 U17095 ( .B1(n13819), .B2(n20912), .A(n13800), .ZN(n13801) );
  OAI211_X1 U17096 ( .C1(n13822), .C2(n20915), .A(n13802), .B(n13801), .ZN(
        P1_U3049) );
  NAND2_X1 U17097 ( .A1(n13815), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13805) );
  OAI22_X1 U17098 ( .A1(n13817), .A2(n15263), .B1(n13816), .B2(n15264), .ZN(
        n13803) );
  AOI21_X1 U17099 ( .B1(n13819), .B2(n20924), .A(n13803), .ZN(n13804) );
  OAI211_X1 U17100 ( .C1(n13822), .C2(n20927), .A(n13805), .B(n13804), .ZN(
        P1_U3051) );
  NAND2_X1 U17101 ( .A1(n13815), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13808) );
  OAI22_X1 U17102 ( .A1(n13817), .A2(n15283), .B1(n13816), .B2(n15284), .ZN(
        n13806) );
  AOI21_X1 U17103 ( .B1(n13819), .B2(n20948), .A(n13806), .ZN(n13807) );
  OAI211_X1 U17104 ( .C1(n13822), .C2(n20951), .A(n13808), .B(n13807), .ZN(
        P1_U3055) );
  NAND2_X1 U17105 ( .A1(n13815), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13811) );
  OAI22_X1 U17106 ( .A1(n13817), .A2(n15258), .B1(n13816), .B2(n15259), .ZN(
        n13809) );
  AOI21_X1 U17107 ( .B1(n13819), .B2(n20918), .A(n13809), .ZN(n13810) );
  OAI211_X1 U17108 ( .C1(n13822), .C2(n20921), .A(n13811), .B(n13810), .ZN(
        P1_U3050) );
  NAND2_X1 U17109 ( .A1(n13815), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13814) );
  OAI22_X1 U17110 ( .A1(n13817), .A2(n15289), .B1(n13816), .B2(n15292), .ZN(
        n13812) );
  AOI21_X1 U17111 ( .B1(n13819), .B2(n20955), .A(n13812), .ZN(n13813) );
  OAI211_X1 U17112 ( .C1(n13822), .C2(n20960), .A(n13814), .B(n13813), .ZN(
        P1_U3056) );
  NAND2_X1 U17113 ( .A1(n13815), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13821) );
  OAI22_X1 U17114 ( .A1(n13817), .A2(n15278), .B1(n13816), .B2(n15279), .ZN(
        n13818) );
  AOI21_X1 U17115 ( .B1(n13819), .B2(n20942), .A(n13818), .ZN(n13820) );
  OAI211_X1 U17116 ( .C1(n13822), .C2(n20945), .A(n13821), .B(n13820), .ZN(
        P1_U3054) );
  NAND2_X1 U17117 ( .A1(n13839), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13826) );
  INV_X1 U17118 ( .A(n13823), .ZN(n13841) );
  OAI22_X1 U17119 ( .A1(n15264), .A2(n13841), .B1(n13840), .B2(n20927), .ZN(
        n13824) );
  AOI21_X1 U17120 ( .B1(n13843), .B2(n20923), .A(n13824), .ZN(n13825) );
  OAI211_X1 U17121 ( .C1(n15211), .C2(n13846), .A(n13826), .B(n13825), .ZN(
        P1_U3067) );
  NAND2_X1 U17122 ( .A1(n13839), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n13829) );
  OAI22_X1 U17123 ( .A1(n15279), .A2(n13841), .B1(n13840), .B2(n20945), .ZN(
        n13827) );
  AOI21_X1 U17124 ( .B1(n13843), .B2(n20941), .A(n13827), .ZN(n13828) );
  OAI211_X1 U17125 ( .C1(n15225), .C2(n13846), .A(n13829), .B(n13828), .ZN(
        P1_U3070) );
  NAND2_X1 U17126 ( .A1(n13839), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13832) );
  OAI22_X1 U17127 ( .A1(n15254), .A2(n13841), .B1(n13840), .B2(n20915), .ZN(
        n13830) );
  AOI21_X1 U17128 ( .B1(n13843), .B2(n20903), .A(n13830), .ZN(n13831) );
  OAI211_X1 U17129 ( .C1(n15201), .C2(n13846), .A(n13832), .B(n13831), .ZN(
        P1_U3065) );
  NAND2_X1 U17130 ( .A1(n13839), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n13835) );
  OAI22_X1 U17131 ( .A1(n15269), .A2(n13841), .B1(n13840), .B2(n20933), .ZN(
        n13833) );
  AOI21_X1 U17132 ( .B1(n13843), .B2(n20929), .A(n13833), .ZN(n13834) );
  OAI211_X1 U17133 ( .C1(n15215), .C2(n13846), .A(n13835), .B(n13834), .ZN(
        P1_U3068) );
  NAND2_X1 U17134 ( .A1(n13839), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13838) );
  OAI22_X1 U17135 ( .A1(n15259), .A2(n13841), .B1(n13840), .B2(n20921), .ZN(
        n13836) );
  AOI21_X1 U17136 ( .B1(n13843), .B2(n20917), .A(n13836), .ZN(n13837) );
  OAI211_X1 U17137 ( .C1(n15206), .C2(n13846), .A(n13838), .B(n13837), .ZN(
        P1_U3066) );
  NAND2_X1 U17138 ( .A1(n13839), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n13845) );
  OAI22_X1 U17139 ( .A1(n15274), .A2(n13841), .B1(n13840), .B2(n20939), .ZN(
        n13842) );
  AOI21_X1 U17140 ( .B1(n13843), .B2(n20935), .A(n13842), .ZN(n13844) );
  OAI211_X1 U17141 ( .C1(n15220), .C2(n13846), .A(n13845), .B(n13844), .ZN(
        P1_U3069) );
  NAND2_X1 U17142 ( .A1(n19774), .A2(n13847), .ZN(n13849) );
  INV_X1 U17143 ( .A(n13849), .ZN(n15586) );
  INV_X1 U17144 ( .A(n13848), .ZN(n13850) );
  OR2_X1 U17145 ( .A1(n13849), .A2(n13848), .ZN(n19768) );
  OAI211_X1 U17146 ( .C1(n15586), .C2(n13850), .A(n19793), .B(n19768), .ZN(
        n13853) );
  NAND2_X1 U17147 ( .A1(n19784), .A2(n13851), .ZN(n13852) );
  OAI211_X1 U17148 ( .C1(n19784), .C2(n10884), .A(n13853), .B(n13852), .ZN(
        P2_U2874) );
  NAND2_X1 U17149 ( .A1(n20588), .A2(n20597), .ZN(n20021) );
  NOR2_X1 U17150 ( .A1(n20262), .A2(n20021), .ZN(n13854) );
  AOI221_X1 U17151 ( .B1(n20042), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20016), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n13854), .ZN(n13857) );
  AOI21_X1 U17152 ( .B1(n10593), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13855) );
  NOR2_X1 U17153 ( .A1(n20257), .A2(n20021), .ZN(n20014) );
  OAI21_X1 U17154 ( .B1(n13855), .B2(n20014), .A(n20425), .ZN(n13856) );
  AOI22_X1 U17155 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19965), .ZN(n20367) );
  AOI22_X1 U17156 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19965), .ZN(n20329) );
  INV_X1 U17157 ( .A(n20329), .ZN(n20440) );
  AOI22_X1 U17158 ( .A1(n20016), .A2(n20441), .B1(n20042), .B2(n20440), .ZN(
        n13865) );
  OAI21_X1 U17159 ( .B1(n13861), .B2(n20014), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13862) );
  OAI21_X1 U17160 ( .B1(n20021), .B2(n20262), .A(n13862), .ZN(n20015) );
  AND2_X1 U17161 ( .A1(n17047), .A2(n19951), .ZN(n20439) );
  AOI22_X1 U17162 ( .A1(n20015), .A2(n13863), .B1(n20439), .B2(n20014), .ZN(
        n13864) );
  OAI211_X1 U17163 ( .C1(n20020), .C2(n13866), .A(n13865), .B(n13864), .ZN(
        P2_U3065) );
  INV_X1 U17164 ( .A(n20896), .ZN(n20858) );
  AOI21_X1 U17165 ( .B1(n13895), .B2(n13891), .A(n20640), .ZN(n13867) );
  AOI21_X1 U17166 ( .B1(n20897), .B2(n20858), .A(n13867), .ZN(n13868) );
  NOR2_X1 U17167 ( .A1(n13868), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13872) );
  NOR2_X1 U17168 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13869), .ZN(
        n13903) );
  OR2_X1 U17169 ( .A1(n13871), .A2(n13870), .ZN(n13873) );
  NAND2_X1 U17170 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13873), .ZN(n20865) );
  NAND2_X1 U17171 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13878) );
  NAND3_X1 U17172 ( .A1(n20897), .A2(n20858), .A3(n15157), .ZN(n13875) );
  INV_X1 U17173 ( .A(n13873), .ZN(n20860) );
  NAND2_X1 U17174 ( .A1(n20899), .A2(n20860), .ZN(n13874) );
  AND2_X1 U17175 ( .A1(n13875), .A2(n13874), .ZN(n13897) );
  OAI22_X1 U17176 ( .A1(n13891), .A2(n15258), .B1(n13897), .B2(n20921), .ZN(
        n13876) );
  AOI21_X1 U17177 ( .B1(n20916), .B2(n13903), .A(n13876), .ZN(n13877) );
  OAI211_X1 U17178 ( .C1(n15206), .C2(n13895), .A(n13878), .B(n13877), .ZN(
        P1_U3146) );
  NAND2_X1 U17179 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13881) );
  OAI22_X1 U17180 ( .A1(n13891), .A2(n15273), .B1(n13897), .B2(n20939), .ZN(
        n13879) );
  AOI21_X1 U17181 ( .B1(n20934), .B2(n13903), .A(n13879), .ZN(n13880) );
  OAI211_X1 U17182 ( .C1(n15220), .C2(n13895), .A(n13881), .B(n13880), .ZN(
        P1_U3149) );
  NAND2_X1 U17183 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13884) );
  OAI22_X1 U17184 ( .A1(n13891), .A2(n15268), .B1(n13897), .B2(n20933), .ZN(
        n13882) );
  AOI21_X1 U17185 ( .B1(n20928), .B2(n13903), .A(n13882), .ZN(n13883) );
  OAI211_X1 U17186 ( .C1(n15215), .C2(n13895), .A(n13884), .B(n13883), .ZN(
        P1_U3148) );
  NAND2_X1 U17187 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13887) );
  OAI22_X1 U17188 ( .A1(n13891), .A2(n15253), .B1(n13897), .B2(n20915), .ZN(
        n13885) );
  AOI21_X1 U17189 ( .B1(n20902), .B2(n13903), .A(n13885), .ZN(n13886) );
  OAI211_X1 U17190 ( .C1(n15201), .C2(n13895), .A(n13887), .B(n13886), .ZN(
        P1_U3145) );
  NAND2_X1 U17191 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13890) );
  OAI22_X1 U17192 ( .A1(n13891), .A2(n15263), .B1(n13897), .B2(n20927), .ZN(
        n13888) );
  AOI21_X1 U17193 ( .B1(n20922), .B2(n13903), .A(n13888), .ZN(n13889) );
  OAI211_X1 U17194 ( .C1(n15211), .C2(n13895), .A(n13890), .B(n13889), .ZN(
        P1_U3147) );
  NAND2_X1 U17195 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13894) );
  OAI22_X1 U17196 ( .A1(n13891), .A2(n15278), .B1(n13897), .B2(n20945), .ZN(
        n13892) );
  AOI21_X1 U17197 ( .B1(n20940), .B2(n13903), .A(n13892), .ZN(n13893) );
  OAI211_X1 U17198 ( .C1(n15225), .C2(n13895), .A(n13894), .B(n13893), .ZN(
        P1_U3150) );
  INV_X1 U17199 ( .A(n13896), .ZN(n13910) );
  INV_X1 U17200 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U17201 ( .A1(n20952), .A2(n13903), .B1(n13902), .B2(n20954), .ZN(
        n13900) );
  INV_X1 U17202 ( .A(n13897), .ZN(n13904) );
  AOI22_X1 U17203 ( .A1(n13906), .A2(n20955), .B1(n13898), .B2(n13904), .ZN(
        n13899) );
  OAI211_X1 U17204 ( .C1(n13910), .C2(n13901), .A(n13900), .B(n13899), .ZN(
        P1_U3152) );
  INV_X1 U17205 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U17206 ( .A1(n20946), .A2(n13903), .B1(n13902), .B2(n20947), .ZN(
        n13908) );
  AOI22_X1 U17207 ( .A1(n13906), .A2(n20948), .B1(n13905), .B2(n13904), .ZN(
        n13907) );
  OAI211_X1 U17208 ( .C1(n13910), .C2(n13909), .A(n13908), .B(n13907), .ZN(
        P1_U3151) );
  NAND2_X1 U17209 ( .A1(n13646), .A2(n13912), .ZN(n13913) );
  AND2_X1 U17210 ( .A1(n13923), .A2(n13913), .ZN(n20668) );
  INV_X1 U17211 ( .A(n20668), .ZN(n13915) );
  OAI222_X1 U17212 ( .A1(n14805), .A2(n13915), .B1(n13914), .B2(n14804), .C1(
        n14802), .C2(n11386), .ZN(P1_U2897) );
  OR2_X1 U17213 ( .A1(n13917), .A2(n13916), .ZN(n13918) );
  NAND2_X1 U17214 ( .A1(n13937), .A2(n13918), .ZN(n20665) );
  OAI22_X1 U17215 ( .A1(n20665), .A2(n14730), .B1(n13919), .B2(n20721), .ZN(
        n13920) );
  AOI21_X1 U17216 ( .B1(n20668), .B2(n20718), .A(n13920), .ZN(n13921) );
  INV_X1 U17217 ( .A(n13921), .ZN(P1_U2865) );
  AOI21_X1 U17218 ( .B1(n13924), .B2(n13923), .A(n13922), .ZN(n14140) );
  INV_X1 U17219 ( .A(n14140), .ZN(n13943) );
  INV_X1 U17220 ( .A(n14804), .ZN(n13977) );
  INV_X1 U17221 ( .A(DATAI_8_), .ZN(n13926) );
  NAND2_X1 U17222 ( .A1(n14738), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13925) );
  OAI21_X1 U17223 ( .B1(n14738), .B2(n13926), .A(n13925), .ZN(n20750) );
  AOI22_X1 U17224 ( .A1(n13977), .A2(n20750), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n16645), .ZN(n13927) );
  OAI21_X1 U17225 ( .B1(n13943), .B2(n14805), .A(n13927), .ZN(P1_U2896) );
  NAND4_X1 U17226 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n13983)
         );
  INV_X1 U17227 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20987) );
  INV_X1 U17228 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20986) );
  INV_X1 U17229 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20814) );
  NOR4_X1 U17230 ( .A1(n21039), .A2(n20987), .A3(n20986), .A4(n20814), .ZN(
        n13929) );
  NAND2_X1 U17231 ( .A1(n13929), .A2(n13928), .ZN(n20682) );
  NOR2_X1 U17232 ( .A1(n13983), .A2(n20682), .ZN(n14385) );
  NOR2_X1 U17233 ( .A1(n16587), .A2(n14385), .ZN(n13985) );
  NAND3_X1 U17234 ( .A1(n20962), .A2(n13928), .A3(n15157), .ZN(n20702) );
  AOI22_X1 U17235 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20705), .B1(
        n14139), .B2(n20687), .ZN(n13934) );
  INV_X1 U17236 ( .A(n20688), .ZN(n13932) );
  INV_X1 U17237 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13931) );
  AND3_X1 U17238 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n13930) );
  NAND3_X1 U17239 ( .A1(n13932), .A2(n13931), .A3(n13930), .ZN(n13933) );
  NAND2_X1 U17240 ( .A1(n13934), .A2(n13933), .ZN(n13935) );
  AOI211_X1 U17241 ( .C1(P1_REIP_REG_8__SCAN_IN), .C2(n13985), .A(n20660), .B(
        n13935), .ZN(n13941) );
  NAND2_X1 U17242 ( .A1(n13937), .A2(n13936), .ZN(n13938) );
  NAND2_X1 U17243 ( .A1(n13981), .A2(n13938), .ZN(n16810) );
  INV_X1 U17244 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13942) );
  OAI22_X1 U17245 ( .A1(n16810), .A2(n20666), .B1(n13942), .B2(n20707), .ZN(
        n13939) );
  INV_X1 U17246 ( .A(n13939), .ZN(n13940) );
  OAI211_X1 U17247 ( .C1(n13943), .C2(n16601), .A(n13941), .B(n13940), .ZN(
        P1_U2832) );
  OAI222_X1 U17248 ( .A1(n13943), .A2(n14699), .B1(n20721), .B2(n13942), .C1(
        n16810), .C2(n14730), .ZN(P1_U2864) );
  NAND2_X1 U17249 ( .A1(n13944), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14663) );
  NOR2_X1 U17250 ( .A1(n20814), .A2(n14663), .ZN(n20695) );
  INV_X1 U17251 ( .A(n20695), .ZN(n13956) );
  INV_X1 U17252 ( .A(n13945), .ZN(n20803) );
  NAND2_X1 U17253 ( .A1(n20700), .A2(n20803), .ZN(n13948) );
  INV_X1 U17254 ( .A(n13962), .ZN(n13946) );
  AOI22_X1 U17255 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n20705), .B1(
        n20687), .B2(n13946), .ZN(n13947) );
  OAI211_X1 U17256 ( .C1(n13949), .C2(n20707), .A(n13948), .B(n13947), .ZN(
        n13951) );
  NOR2_X1 U17257 ( .A1(n13960), .A2(n14655), .ZN(n13950) );
  AOI211_X1 U17258 ( .C1(n20698), .C2(n13150), .A(n13951), .B(n13950), .ZN(
        n13955) );
  OAI21_X1 U17259 ( .B1(n13952), .B2(n21039), .A(n20683), .ZN(n14662) );
  OAI21_X1 U17260 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n14663), .A(n14662), .ZN(
        n13953) );
  NAND2_X1 U17261 ( .A1(n13953), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13954) );
  OAI211_X1 U17262 ( .C1(n13956), .C2(P1_REIP_REG_3__SCAN_IN), .A(n13955), .B(
        n13954), .ZN(P1_U2837) );
  OAI21_X1 U17263 ( .B1(n13959), .B2(n13958), .A(n13957), .ZN(n20804) );
  INV_X1 U17264 ( .A(n13960), .ZN(n13964) );
  AOI22_X1 U17265 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13961) );
  OAI21_X1 U17266 ( .B1(n16695), .B2(n13962), .A(n13961), .ZN(n13963) );
  AOI21_X1 U17267 ( .B1(n13964), .B2(n20791), .A(n13963), .ZN(n13965) );
  OAI21_X1 U17268 ( .B1(n20804), .B2(n21068), .A(n13965), .ZN(P1_U2996) );
  OAI21_X1 U17269 ( .B1(n13968), .B2(n13967), .A(n13966), .ZN(n20816) );
  AOI22_X1 U17270 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13969) );
  OAI21_X1 U17271 ( .B1(n16695), .B2(n14657), .A(n13969), .ZN(n13970) );
  AOI21_X1 U17272 ( .B1(n14666), .B2(n20791), .A(n13970), .ZN(n13971) );
  OAI21_X1 U17273 ( .B1(n21068), .B2(n20816), .A(n13971), .ZN(P1_U2997) );
  NOR2_X1 U17274 ( .A1(n13922), .A2(n13973), .ZN(n13974) );
  OR2_X1 U17275 ( .A1(n13972), .A2(n13974), .ZN(n14152) );
  INV_X1 U17276 ( .A(DATAI_9_), .ZN(n13976) );
  NAND2_X1 U17277 ( .A1(n14738), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13975) );
  OAI21_X1 U17278 ( .B1(n14738), .B2(n13976), .A(n13975), .ZN(n20752) );
  AOI22_X1 U17279 ( .A1(n13977), .A2(n20752), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n16645), .ZN(n13978) );
  OAI21_X1 U17280 ( .B1(n14152), .B2(n14805), .A(n13978), .ZN(P1_U2895) );
  INV_X1 U17281 ( .A(n14032), .ZN(n13979) );
  AOI21_X1 U17282 ( .B1(n13981), .B2(n13980), .A(n13979), .ZN(n16791) );
  AOI22_X1 U17283 ( .A1(n16791), .A2(n20717), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14715), .ZN(n13982) );
  OAI21_X1 U17284 ( .B1(n14152), .B2(n14699), .A(n13982), .ZN(P1_U2863) );
  NOR2_X2 U17285 ( .A1(n20688), .A2(n13983), .ZN(n16630) );
  INV_X1 U17286 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14063) );
  INV_X1 U17287 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13990) );
  NAND2_X1 U17288 ( .A1(n16791), .A2(n20700), .ZN(n13989) );
  INV_X1 U17289 ( .A(n13984), .ZN(n14154) );
  AOI21_X1 U17290 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n13985), .A(n20660), .ZN(
        n13986) );
  OAI21_X1 U17291 ( .B1(n20703), .B2(n14154), .A(n13986), .ZN(n13987) );
  AOI21_X1 U17292 ( .B1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20705), .A(
        n13987), .ZN(n13988) );
  OAI211_X1 U17293 ( .C1(n13990), .C2(n20707), .A(n13989), .B(n13988), .ZN(
        n13991) );
  AOI21_X1 U17294 ( .B1(n16630), .B2(n14063), .A(n13991), .ZN(n13992) );
  OAI21_X1 U17295 ( .B1(n14152), .B2(n16601), .A(n13992), .ZN(P1_U2831) );
  XNOR2_X1 U17296 ( .A(n13993), .B(n19906), .ZN(n13995) );
  XNOR2_X1 U17297 ( .A(n13995), .B(n13994), .ZN(n19917) );
  NAND2_X1 U17298 ( .A1(n13997), .A2(n13996), .ZN(n13998) );
  AND2_X1 U17299 ( .A1(n13999), .A2(n13998), .ZN(n19914) );
  OR2_X1 U17300 ( .A1(n14001), .A2(n14000), .ZN(n14002) );
  NAND2_X1 U17301 ( .A1(n14002), .A2(n13101), .ZN(n19912) );
  INV_X1 U17302 ( .A(n19752), .ZN(n19755) );
  OAI22_X1 U17303 ( .A1(n16950), .A2(n14004), .B1(n19736), .B2(n14003), .ZN(
        n14005) );
  AOI21_X1 U17304 ( .B1(n16942), .B2(n19755), .A(n14005), .ZN(n14006) );
  OAI21_X1 U17305 ( .B1(n19912), .B2(n13859), .A(n14006), .ZN(n14007) );
  AOI21_X1 U17306 ( .B1(n19914), .B2(n15927), .A(n14007), .ZN(n14008) );
  OAI21_X1 U17307 ( .B1(n16955), .B2(n19917), .A(n14008), .ZN(P2_U3010) );
  OAI21_X1 U17308 ( .B1(n14011), .B2(n14010), .A(n14009), .ZN(n15917) );
  INV_X1 U17309 ( .A(n14012), .ZN(n14018) );
  NAND2_X1 U17310 ( .A1(n14017), .A2(n14013), .ZN(n14016) );
  INV_X1 U17311 ( .A(n14014), .ZN(n14015) );
  AOI22_X1 U17312 ( .A1(n14018), .A2(n14017), .B1(n14016), .B2(n14015), .ZN(
        n15920) );
  NOR2_X1 U17313 ( .A1(n14023), .A2(n19906), .ZN(n14455) );
  AOI221_X1 U17314 ( .B1(n19935), .B2(n14019), .C1(n19918), .C2(n14019), .A(
        n10049), .ZN(n14454) );
  INV_X1 U17315 ( .A(n14454), .ZN(n19907) );
  AOI211_X1 U17316 ( .C1(n14023), .C2(n19906), .A(n14455), .B(n19907), .ZN(
        n14028) );
  OAI21_X1 U17317 ( .B1(n19741), .B2(n14021), .A(n14020), .ZN(n19843) );
  AOI21_X1 U17318 ( .B1(n10049), .B2(n16497), .A(n14022), .ZN(n19905) );
  OAI22_X1 U17319 ( .A1(n19736), .A2(n14024), .B1(n19905), .B2(n14023), .ZN(
        n14025) );
  AOI21_X1 U17320 ( .B1(n19931), .B2(n15921), .A(n14025), .ZN(n14026) );
  OAI21_X1 U17321 ( .B1(n19843), .B2(n19928), .A(n14026), .ZN(n14027) );
  AOI211_X1 U17322 ( .C1(n15920), .C2(n17013), .A(n14028), .B(n14027), .ZN(
        n14029) );
  OAI21_X1 U17323 ( .B1(n17009), .B2(n15917), .A(n14029), .ZN(P2_U3041) );
  OAI21_X1 U17324 ( .B1(n13972), .B2(n14031), .A(n14030), .ZN(n14952) );
  AOI21_X1 U17325 ( .B1(n14033), .B2(n14032), .A(n14159), .ZN(n16780) );
  AOI22_X1 U17326 ( .A1(n16780), .A2(n20717), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14715), .ZN(n14034) );
  OAI21_X1 U17327 ( .B1(n14952), .B2(n14731), .A(n14034), .ZN(P1_U2862) );
  INV_X1 U17328 ( .A(n14035), .ZN(n15492) );
  NAND2_X1 U17329 ( .A1(n15517), .A2(n15492), .ZN(n15506) );
  NOR2_X1 U17330 ( .A1(n19673), .A2(n14036), .ZN(n14048) );
  INV_X1 U17331 ( .A(n14036), .ZN(n16934) );
  OR2_X1 U17332 ( .A1(n14038), .A2(n14037), .ZN(n14039) );
  NAND2_X1 U17333 ( .A1(n14039), .A2(n15493), .ZN(n19822) );
  INV_X1 U17334 ( .A(n19822), .ZN(n16154) );
  NAND2_X1 U17335 ( .A1(n19743), .A2(n16154), .ZN(n14042) );
  AOI22_X1 U17336 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19732), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19652), .ZN(n14041) );
  NAND2_X1 U17337 ( .A1(n19692), .A2(n16938), .ZN(n14040) );
  AND4_X1 U17338 ( .A1(n14042), .A2(n14041), .A3(n19736), .A4(n14040), .ZN(
        n14044) );
  NAND2_X1 U17339 ( .A1(n19744), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n14043) );
  OAI211_X1 U17340 ( .C1(n19684), .C2(n14045), .A(n14044), .B(n14043), .ZN(
        n14046) );
  AOI21_X1 U17341 ( .B1(n15465), .B2(n16934), .A(n14046), .ZN(n14047) );
  OAI21_X1 U17342 ( .B1(n15506), .B2(n14048), .A(n14047), .ZN(P2_U2844) );
  AOI21_X1 U17343 ( .B1(n19757), .B2(n19698), .A(n15465), .ZN(n14062) );
  INV_X1 U17344 ( .A(n15902), .ZN(n14049) );
  NOR3_X1 U17345 ( .A1(n14128), .A2(n14049), .A3(n19698), .ZN(n14060) );
  OAI21_X1 U17346 ( .B1(n14052), .B2(n14051), .A(n14050), .ZN(n19792) );
  AOI22_X1 U17347 ( .A1(n14053), .A2(n19734), .B1(n19744), .B2(
        P2_EBX_REG_8__SCAN_IN), .ZN(n14054) );
  OAI211_X1 U17348 ( .C1(n12689), .C2(n19737), .A(n14054), .B(n19736), .ZN(
        n14055) );
  AOI21_X1 U17349 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19732), .A(
        n14055), .ZN(n14058) );
  AOI21_X1 U17350 ( .B1(n14056), .B2(n16177), .A(n16163), .ZN(n19828) );
  NAND2_X1 U17351 ( .A1(n19743), .A2(n19828), .ZN(n14057) );
  OAI211_X1 U17352 ( .C1(n19792), .C2(n19748), .A(n14058), .B(n14057), .ZN(
        n14059) );
  NOR2_X1 U17353 ( .A1(n14060), .A2(n14059), .ZN(n14061) );
  OAI21_X1 U17354 ( .B1(n14062), .B2(n15902), .A(n14061), .ZN(P2_U2847) );
  INV_X1 U17355 ( .A(n16630), .ZN(n16623) );
  INV_X1 U17356 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20996) );
  OAI21_X1 U17357 ( .B1(n16623), .B2(n14063), .A(n20996), .ZN(n14065) );
  NOR2_X1 U17358 ( .A1(n20996), .A2(n14063), .ZN(n14064) );
  AOI21_X1 U17359 ( .B1(n14385), .B2(n14064), .A(n16587), .ZN(n16634) );
  NAND2_X1 U17360 ( .A1(n14065), .A2(n16634), .ZN(n14072) );
  INV_X1 U17361 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14069) );
  INV_X1 U17362 ( .A(n14066), .ZN(n14949) );
  OAI21_X1 U17363 ( .B1(n16596), .B2(n14946), .A(n20702), .ZN(n14067) );
  AOI21_X1 U17364 ( .B1(n20687), .B2(n14949), .A(n14067), .ZN(n14068) );
  OAI21_X1 U17365 ( .B1(n14069), .B2(n20707), .A(n14068), .ZN(n14070) );
  AOI21_X1 U17366 ( .B1(n16780), .B2(n20700), .A(n14070), .ZN(n14071) );
  OAI211_X1 U17367 ( .C1(n14952), .C2(n16601), .A(n14072), .B(n14071), .ZN(
        P1_U2830) );
  INV_X1 U17368 ( .A(n15511), .ZN(n19749) );
  AOI21_X1 U17369 ( .B1(n14073), .B2(n15518), .A(n14127), .ZN(n14074) );
  NAND2_X1 U17370 ( .A1(n19753), .A2(n14074), .ZN(n14479) );
  INV_X1 U17371 ( .A(n14479), .ZN(n14075) );
  AOI22_X1 U17372 ( .A1(n15465), .A2(n14076), .B1(n14075), .B2(n19757), .ZN(
        n14085) );
  NAND2_X1 U17373 ( .A1(n19744), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n14080) );
  NOR2_X1 U17374 ( .A1(n19654), .A2(n14076), .ZN(n14077) );
  AOI21_X1 U17375 ( .B1(n19734), .B2(n14078), .A(n14077), .ZN(n14079) );
  OAI211_X1 U17376 ( .C1(n19737), .C2(n14081), .A(n14080), .B(n14079), .ZN(
        n14083) );
  NOR2_X1 U17377 ( .A1(n16217), .A2(n19748), .ZN(n14082) );
  AOI211_X1 U17378 ( .C1(n20603), .C2(n19743), .A(n14083), .B(n14082), .ZN(
        n14084) );
  OAI211_X1 U17379 ( .C1(n16223), .C2(n19749), .A(n14085), .B(n14084), .ZN(
        P2_U2854) );
  MUX2_X1 U17380 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n15518), .S(
        n19753), .Z(n14478) );
  INV_X1 U17381 ( .A(n14478), .ZN(n14092) );
  OR2_X1 U17382 ( .A1(n17014), .A2(n16216), .ZN(n14089) );
  INV_X1 U17383 ( .A(n12770), .ZN(n14087) );
  NAND2_X1 U17384 ( .A1(n14087), .A2(n14086), .ZN(n16214) );
  NAND2_X1 U17385 ( .A1(n16214), .A2(n17035), .ZN(n14088) );
  AND2_X1 U17386 ( .A1(n14089), .A2(n14088), .ZN(n17034) );
  OAI22_X1 U17387 ( .A1(n17034), .A2(n20568), .B1(n14090), .B2(n20569), .ZN(
        n14091) );
  AOI21_X1 U17388 ( .B1(n14092), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n14091), 
        .ZN(n14094) );
  AOI21_X1 U17389 ( .B1(n17033), .B2(n20579), .A(n20571), .ZN(n14093) );
  OAI22_X1 U17390 ( .A1(n14094), .A2(n20571), .B1(n14093), .B2(n17035), .ZN(
        P2_U3601) );
  INV_X1 U17391 ( .A(n16911), .ZN(n14096) );
  AOI21_X1 U17392 ( .B1(n14097), .B2(n14095), .A(n14096), .ZN(n15579) );
  INV_X1 U17393 ( .A(n19859), .ZN(n15657) );
  OR2_X1 U17394 ( .A1(n14099), .A2(n14098), .ZN(n14100) );
  NAND2_X1 U17395 ( .A1(n15453), .A2(n14100), .ZN(n19651) );
  AOI22_X1 U17396 ( .A1(n19804), .A2(BUF2_REG_17__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14103) );
  AOI22_X1 U17397 ( .A1(n19802), .A2(n14101), .B1(n19858), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n14102) );
  OAI211_X1 U17398 ( .C1(n15657), .C2(n19651), .A(n14103), .B(n14102), .ZN(
        n14104) );
  AOI21_X1 U17399 ( .B1(n15579), .B2(n19848), .A(n14104), .ZN(n14105) );
  INV_X1 U17400 ( .A(n14105), .ZN(P2_U2902) );
  INV_X1 U17401 ( .A(DATAI_10_), .ZN(n14106) );
  INV_X1 U17402 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17203) );
  MUX2_X1 U17403 ( .A(n14106), .B(n17203), .S(n14738), .Z(n20754) );
  INV_X1 U17404 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14107) );
  OAI222_X1 U17405 ( .A1(n14952), .A2(n14805), .B1(n20754), .B2(n14804), .C1(
        n14107), .C2(n14802), .ZN(P1_U2894) );
  AOI21_X1 U17406 ( .B1(n19757), .B2(n14114), .A(n15465), .ZN(n14121) );
  NOR2_X1 U17407 ( .A1(n19737), .A2(n12673), .ZN(n14111) );
  OAI22_X1 U17408 ( .A1(n19684), .A2(n14109), .B1(n19654), .B2(n14108), .ZN(
        n14110) );
  AOI211_X1 U17409 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19744), .A(n14111), .B(
        n14110), .ZN(n14112) );
  OAI21_X1 U17410 ( .B1(n14113), .B2(n19748), .A(n14112), .ZN(n14117) );
  NOR3_X1 U17411 ( .A1(n14128), .A2(n14115), .A3(n14114), .ZN(n14116) );
  AOI211_X1 U17412 ( .C1(n20584), .C2(n19743), .A(n14117), .B(n14116), .ZN(
        n14119) );
  NAND2_X1 U17413 ( .A1(n20582), .A2(n15511), .ZN(n14118) );
  OAI211_X1 U17414 ( .C1(n14121), .C2(n14120), .A(n14119), .B(n14118), .ZN(
        P2_U2852) );
  AOI21_X1 U17415 ( .B1(n19757), .B2(n14127), .A(n15465), .ZN(n14133) );
  OAI22_X1 U17416 ( .A1(n20590), .A2(n19726), .B1(n12800), .B2(n19654), .ZN(
        n14124) );
  NOR2_X1 U17417 ( .A1(n19684), .A2(n14122), .ZN(n14123) );
  AOI211_X1 U17418 ( .C1(n19652), .C2(P2_REIP_REG_2__SCAN_IN), .A(n14124), .B(
        n14123), .ZN(n14125) );
  OAI21_X1 U17419 ( .B1(n19683), .B2(n14126), .A(n14125), .ZN(n14130) );
  INV_X1 U17420 ( .A(n14132), .ZN(n14439) );
  NOR3_X1 U17421 ( .A1(n14128), .A2(n14439), .A3(n14127), .ZN(n14129) );
  INV_X1 U17422 ( .A(n20054), .ZN(n20595) );
  NAND2_X1 U17423 ( .A1(n20595), .A2(n15511), .ZN(n14131) );
  OAI211_X1 U17424 ( .C1(n14133), .C2(n14132), .A(n9707), .B(n14131), .ZN(
        P2_U2853) );
  OAI21_X1 U17425 ( .B1(n14136), .B2(n14135), .A(n14134), .ZN(n16809) );
  OAI22_X1 U17426 ( .A1(n14947), .A2(n14137), .B1(n16817), .B2(n13931), .ZN(
        n14138) );
  AOI21_X1 U17427 ( .B1(n14139), .B2(n16669), .A(n14138), .ZN(n14142) );
  NAND2_X1 U17428 ( .A1(n14140), .A2(n20791), .ZN(n14141) );
  OAI211_X1 U17429 ( .C1(n16809), .C2(n21068), .A(n14142), .B(n14141), .ZN(
        P1_U2991) );
  OR2_X1 U17430 ( .A1(n14144), .A2(n14143), .ZN(n14145) );
  AND2_X1 U17431 ( .A1(n14146), .A2(n14145), .ZN(n16679) );
  INV_X1 U17432 ( .A(n16679), .ZN(n14160) );
  INV_X1 U17433 ( .A(DATAI_11_), .ZN(n14148) );
  MUX2_X1 U17434 ( .A(n14148), .B(n14147), .S(n14738), .Z(n20757) );
  INV_X1 U17435 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14149) );
  OAI222_X1 U17436 ( .A1(n14160), .A2(n14805), .B1(n20757), .B2(n14804), .C1(
        n14149), .C2(n14802), .ZN(P1_U2893) );
  OAI21_X1 U17437 ( .B1(n14151), .B2(n14150), .A(n16675), .ZN(n16792) );
  INV_X1 U17438 ( .A(n14152), .ZN(n14156) );
  AOI22_X1 U17439 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14153) );
  OAI21_X1 U17440 ( .B1(n16695), .B2(n14154), .A(n14153), .ZN(n14155) );
  AOI21_X1 U17441 ( .B1(n14156), .B2(n20791), .A(n14155), .ZN(n14157) );
  OAI21_X1 U17442 ( .B1(n16792), .B2(n21068), .A(n14157), .ZN(P1_U2990) );
  OAI21_X1 U17443 ( .B1(n14159), .B2(n14158), .A(n14729), .ZN(n16631) );
  INV_X1 U17444 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14161) );
  OAI222_X1 U17445 ( .A1(n16631), .A2(n14730), .B1(n14161), .B2(n20721), .C1(
        n14160), .C2(n14699), .ZN(P1_U2861) );
  INV_X1 U17446 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n14268) );
  NAND2_X1 U17447 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17674) );
  INV_X1 U17448 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17431) );
  INV_X1 U17449 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17479) );
  INV_X1 U17450 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17503) );
  INV_X1 U17451 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17842) );
  INV_X1 U17452 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17860) );
  AOI22_X1 U17453 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14165) );
  INV_X4 U17454 ( .A(n16345), .ZN(n17902) );
  AOI22_X1 U17455 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14164) );
  INV_X2 U17456 ( .A(n10197), .ZN(n17882) );
  AOI22_X1 U17457 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14163) );
  INV_X4 U17458 ( .A(n16247), .ZN(n17894) );
  AOI22_X1 U17459 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14162) );
  NAND4_X1 U17460 ( .A1(n14165), .A2(n14164), .A3(n14163), .A4(n14162), .ZN(
        n14179) );
  INV_X4 U17461 ( .A(n17847), .ZN(n17876) );
  AOI22_X1 U17462 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14177) );
  INV_X2 U17463 ( .A(n17708), .ZN(n17875) );
  AOI22_X1 U17464 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14176) );
  INV_X4 U17465 ( .A(n14256), .ZN(n17862) );
  INV_X4 U17466 ( .A(n16367), .ZN(n17892) );
  AOI22_X1 U17467 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14175) );
  AOI22_X1 U17468 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n17883), .B1(
        n17816), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14174) );
  NAND4_X1 U17469 ( .A1(n14177), .A2(n14176), .A3(n14175), .A4(n14174), .ZN(
        n14178) );
  AOI22_X1 U17470 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14183) );
  AOI22_X1 U17471 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14182) );
  AOI22_X1 U17472 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n17816), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14181) );
  AOI22_X1 U17473 ( .A1(n17883), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14180) );
  NAND4_X1 U17474 ( .A1(n14183), .A2(n14182), .A3(n14181), .A4(n14180), .ZN(
        n14189) );
  AOI22_X1 U17475 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14187) );
  AOI22_X1 U17476 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14186) );
  AOI22_X1 U17477 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n17902), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14185) );
  AOI22_X1 U17478 ( .A1(n16346), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14184) );
  NAND4_X1 U17479 ( .A1(n14187), .A2(n14186), .A3(n14185), .A4(n14184), .ZN(
        n14188) );
  AOI22_X1 U17480 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14201) );
  AOI22_X1 U17481 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n9595), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14200) );
  AOI22_X1 U17482 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14191) );
  OAI21_X1 U17483 ( .B1(n21216), .B2(n14192), .A(n14191), .ZN(n14198) );
  AOI22_X1 U17484 ( .A1(n17883), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14196) );
  AOI22_X1 U17485 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14195) );
  AOI22_X1 U17486 ( .A1(n17902), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14194) );
  AOI22_X1 U17487 ( .A1(n16346), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14193) );
  NAND4_X1 U17488 ( .A1(n14196), .A2(n14195), .A3(n14194), .A4(n14193), .ZN(
        n14197) );
  AOI211_X1 U17489 ( .C1(n17893), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n14198), .B(n14197), .ZN(n14199) );
  NAND3_X1 U17490 ( .A1(n14201), .A2(n14200), .A3(n14199), .ZN(n16416) );
  NAND2_X1 U17491 ( .A1(n18934), .A2(n18930), .ZN(n19368) );
  AOI22_X1 U17492 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14205) );
  AOI22_X1 U17493 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14204) );
  AOI22_X1 U17494 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n14232), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14203) );
  AOI22_X1 U17495 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14202) );
  NAND4_X1 U17496 ( .A1(n14205), .A2(n14204), .A3(n14203), .A4(n14202), .ZN(
        n14211) );
  AOI22_X1 U17497 ( .A1(n17816), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14209) );
  AOI22_X1 U17498 ( .A1(n16346), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14208) );
  AOI22_X1 U17499 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17862), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14207) );
  AOI22_X1 U17500 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14206) );
  NAND4_X1 U17501 ( .A1(n14209), .A2(n14208), .A3(n14207), .A4(n14206), .ZN(
        n14210) );
  AOI22_X1 U17502 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14221) );
  AOI22_X1 U17503 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14220) );
  AOI22_X1 U17504 ( .A1(n17883), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14212) );
  OAI21_X1 U17505 ( .B1(n21139), .B2(n10197), .A(n14212), .ZN(n14218) );
  INV_X2 U17506 ( .A(n10198), .ZN(n17893) );
  AOI22_X1 U17507 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14216) );
  AOI22_X1 U17508 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n14232), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14215) );
  AOI22_X1 U17509 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14214) );
  AOI22_X1 U17510 ( .A1(n16346), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14213) );
  NAND4_X1 U17511 ( .A1(n14216), .A2(n14215), .A3(n14214), .A4(n14213), .ZN(
        n14217) );
  AOI211_X1 U17512 ( .C1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .C2(n17895), .A(
        n14218), .B(n14217), .ZN(n14219) );
  NAND3_X1 U17513 ( .A1(n14221), .A2(n14220), .A3(n14219), .ZN(n16417) );
  NAND2_X1 U17514 ( .A1(n18942), .A2(n16417), .ZN(n16288) );
  AOI22_X1 U17515 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14225) );
  AOI22_X1 U17516 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17892), .ZN(n14224) );
  AOI22_X1 U17517 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n14232), .ZN(n14223) );
  AOI22_X1 U17518 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17894), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17901), .ZN(n14222) );
  NAND4_X1 U17519 ( .A1(n14225), .A2(n14224), .A3(n14223), .A4(n14222), .ZN(
        n14231) );
  AOI22_X1 U17520 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17895), .B1(
        n17862), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14229) );
  AOI22_X1 U17521 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17902), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17882), .ZN(n14228) );
  AOI22_X1 U17522 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17877), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U17523 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17903), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17883), .ZN(n14226) );
  NAND4_X1 U17524 ( .A1(n14229), .A2(n14228), .A3(n14227), .A4(n14226), .ZN(
        n14230) );
  INV_X2 U17525 ( .A(n14343), .ZN(n17895) );
  AOI22_X1 U17526 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14236) );
  AOI22_X1 U17527 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14235) );
  AOI22_X1 U17528 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14234) );
  AOI22_X1 U17529 ( .A1(n17894), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14233) );
  NAND4_X1 U17530 ( .A1(n14236), .A2(n14235), .A3(n14234), .A4(n14233), .ZN(
        n14242) );
  AOI22_X1 U17531 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14240) );
  AOI22_X1 U17532 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17903), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14239) );
  AOI22_X1 U17533 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14238) );
  AOI22_X1 U17534 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14237) );
  NAND4_X1 U17535 ( .A1(n14240), .A2(n14239), .A3(n14238), .A4(n14237), .ZN(
        n14241) );
  NOR2_X1 U17536 ( .A1(n18087), .A2(n16273), .ZN(n14254) );
  OAI22_X1 U17537 ( .A1(n19548), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n19387), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16263) );
  NAND2_X1 U17538 ( .A1(n19385), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16264) );
  NOR2_X1 U17539 ( .A1(n16263), .A2(n16264), .ZN(n14243) );
  AOI22_X1 U17540 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n19403), .B2(n19541), .ZN(
        n14248) );
  NOR2_X1 U17541 ( .A1(n14249), .A2(n14248), .ZN(n14244) );
  AOI22_X1 U17542 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17605), .B1(
        n14245), .B2(n19531), .ZN(n14252) );
  NOR2_X1 U17543 ( .A1(n14245), .A2(n19531), .ZN(n14251) );
  NAND2_X1 U17544 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17605), .ZN(
        n14246) );
  OAI22_X1 U17545 ( .A1(n14252), .A2(n18918), .B1(n14251), .B2(n14246), .ZN(
        n14250) );
  INV_X1 U17546 ( .A(n14250), .ZN(n14247) );
  OAI211_X1 U17547 ( .C1(n19385), .C2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n16264), .B(n14247), .ZN(n16420) );
  XNOR2_X1 U17548 ( .A(n14249), .B(n14248), .ZN(n16421) );
  INV_X1 U17549 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18916) );
  OR2_X1 U17550 ( .A1(n14251), .A2(n18918), .ZN(n14253) );
  OAI211_X1 U17551 ( .C1(n16263), .C2(n16420), .A(n16267), .B(n16265), .ZN(
        n17089) );
  INV_X1 U17552 ( .A(n18934), .ZN(n16274) );
  NAND2_X1 U17553 ( .A1(n16270), .A2(n18930), .ZN(n16271) );
  INV_X2 U17554 ( .A(n16417), .ZN(n18945) );
  NAND2_X1 U17555 ( .A1(n16273), .A2(n18945), .ZN(n19369) );
  NOR2_X2 U17556 ( .A1(n17089), .A2(n16433), .ZN(n16296) );
  INV_X1 U17557 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17937) );
  AOI22_X1 U17558 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14255) );
  OAI21_X1 U17559 ( .B1(n14256), .B2(n17937), .A(n14255), .ZN(n14262) );
  AOI22_X1 U17560 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14260) );
  AOI22_X1 U17561 ( .A1(n17902), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14259) );
  AOI22_X1 U17562 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14258) );
  AOI22_X1 U17563 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14257) );
  NAND4_X1 U17564 ( .A1(n14260), .A2(n14259), .A3(n14258), .A4(n14257), .ZN(
        n14261) );
  AOI211_X1 U17565 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n17883), .A(
        n14262), .B(n14261), .ZN(n14263) );
  NAND2_X1 U17566 ( .A1(n19572), .A2(n19574), .ZN(n17091) );
  INV_X1 U17567 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17914) );
  INV_X1 U17568 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17913) );
  NAND3_X1 U17569 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n17912) );
  NOR4_X1 U17570 ( .A1(n17581), .A2(n17914), .A3(n17913), .A4(n17912), .ZN(
        n14266) );
  AND4_X2 U17571 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(n17938), .A4(n14266), .ZN(n17917) );
  AND2_X2 U17572 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17917), .ZN(n17911) );
  NAND2_X1 U17573 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17829), .ZN(n17812) );
  NAND4_X1 U17574 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(P3_EBX_REG_16__SCAN_IN), .A4(n17788), .ZN(n17758) );
  NAND3_X1 U17575 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(P3_EBX_REG_20__SCAN_IN), 
        .A3(n17744), .ZN(n17732) );
  NAND4_X1 U17576 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(P3_EBX_REG_23__SCAN_IN), .A4(P3_EBX_REG_22__SCAN_IN), .ZN(n14267)
         );
  NAND3_X1 U17577 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(P3_EBX_REG_29__SCAN_IN), 
        .A3(n17670), .ZN(n16245) );
  INV_X1 U17578 ( .A(n16245), .ZN(n16243) );
  AOI21_X1 U17579 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n17670), .A(
        P3_EBX_REG_30__SCAN_IN), .ZN(n14269) );
  NOR2_X1 U17580 ( .A1(n16243), .A2(n14269), .ZN(n14366) );
  AOI22_X1 U17581 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17902), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14273) );
  AOI22_X1 U17582 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17900), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17882), .ZN(n14272) );
  AOI22_X1 U17583 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17883), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n14232), .ZN(n14271) );
  AOI22_X1 U17584 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17876), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17894), .ZN(n14270) );
  NAND4_X1 U17585 ( .A1(n14273), .A2(n14272), .A3(n14271), .A4(n14270), .ZN(
        n14279) );
  AOI22_X1 U17586 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17903), .ZN(n14277) );
  AOI22_X1 U17587 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14276) );
  AOI22_X1 U17588 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14275) );
  AOI22_X1 U17589 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17901), .B1(
        n17816), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14274) );
  NAND4_X1 U17590 ( .A1(n14277), .A2(n14276), .A3(n14275), .A4(n14274), .ZN(
        n14278) );
  NOR2_X1 U17591 ( .A1(n14279), .A2(n14278), .ZN(n14364) );
  AOI22_X1 U17592 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14283) );
  AOI22_X1 U17593 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14282) );
  AOI22_X1 U17594 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14281) );
  AOI22_X1 U17595 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14280) );
  NAND4_X1 U17596 ( .A1(n14283), .A2(n14282), .A3(n14281), .A4(n14280), .ZN(
        n14290) );
  AOI22_X1 U17597 ( .A1(n16346), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14288) );
  AOI22_X1 U17598 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n16368), .B1(
        n17816), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14287) );
  AOI22_X1 U17599 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14286) );
  AOI22_X1 U17600 ( .A1(n17883), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14285) );
  NAND4_X1 U17601 ( .A1(n14288), .A2(n14287), .A3(n14286), .A4(n14285), .ZN(
        n14289) );
  NOR2_X1 U17602 ( .A1(n14290), .A2(n14289), .ZN(n17678) );
  AOI22_X1 U17603 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14294) );
  AOI22_X1 U17604 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14293) );
  AOI22_X1 U17605 ( .A1(n16346), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14292) );
  AOI22_X1 U17606 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n17862), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14291) );
  NAND4_X1 U17607 ( .A1(n14294), .A2(n14293), .A3(n14292), .A4(n14291), .ZN(
        n14300) );
  AOI22_X1 U17608 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n17882), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14298) );
  AOI22_X1 U17609 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14297) );
  AOI22_X1 U17610 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14296) );
  AOI22_X1 U17611 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14295) );
  NAND4_X1 U17612 ( .A1(n14298), .A2(n14297), .A3(n14296), .A4(n14295), .ZN(
        n14299) );
  NOR2_X1 U17613 ( .A1(n14300), .A2(n14299), .ZN(n17688) );
  AOI22_X1 U17614 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14304) );
  AOI22_X1 U17615 ( .A1(n17902), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14303) );
  AOI22_X1 U17616 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17903), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14302) );
  AOI22_X1 U17617 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17894), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14301) );
  NAND4_X1 U17618 ( .A1(n14304), .A2(n14303), .A3(n14302), .A4(n14301), .ZN(
        n14310) );
  AOI22_X1 U17619 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14308) );
  AOI22_X1 U17620 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14307) );
  AOI22_X1 U17621 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14306) );
  AOI22_X1 U17622 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14305) );
  NAND4_X1 U17623 ( .A1(n14308), .A2(n14307), .A3(n14306), .A4(n14305), .ZN(
        n14309) );
  NOR2_X1 U17624 ( .A1(n14310), .A2(n14309), .ZN(n17697) );
  AOI22_X1 U17625 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U17626 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14319) );
  INV_X1 U17627 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n21156) );
  AOI22_X1 U17628 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14311) );
  OAI21_X1 U17629 ( .B1(n21156), .B2(n16247), .A(n14311), .ZN(n14317) );
  AOI22_X1 U17630 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17903), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14315) );
  AOI22_X1 U17631 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U17632 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14313) );
  AOI22_X1 U17633 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14312) );
  NAND4_X1 U17634 ( .A1(n14315), .A2(n14314), .A3(n14313), .A4(n14312), .ZN(
        n14316) );
  AOI211_X1 U17635 ( .C1(n17900), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n14317), .B(n14316), .ZN(n14318) );
  NAND3_X1 U17636 ( .A1(n14320), .A2(n14319), .A3(n14318), .ZN(n17702) );
  AOI22_X1 U17637 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14330) );
  AOI22_X1 U17638 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17877), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14329) );
  INV_X1 U17639 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16303) );
  AOI22_X1 U17640 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17901), .ZN(n14321) );
  OAI21_X1 U17641 ( .B1(n16303), .B2(n10198), .A(n14321), .ZN(n14327) );
  AOI22_X1 U17642 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n9595), .B1(
        n17903), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14325) );
  AOI22_X1 U17643 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17883), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14324) );
  AOI22_X1 U17644 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17894), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U17645 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14232), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17902), .ZN(n14322) );
  NAND4_X1 U17646 ( .A1(n14325), .A2(n14324), .A3(n14323), .A4(n14322), .ZN(
        n14326) );
  AOI211_X1 U17647 ( .C1(n17862), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n14327), .B(n14326), .ZN(n14328) );
  NAND3_X1 U17648 ( .A1(n14330), .A2(n14329), .A3(n14328), .ZN(n17703) );
  NAND2_X1 U17649 ( .A1(n17702), .A2(n17703), .ZN(n17701) );
  NOR2_X1 U17650 ( .A1(n17697), .A2(n17701), .ZN(n17694) );
  AOI22_X1 U17651 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U17652 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U17653 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14331) );
  OAI21_X1 U17654 ( .B1(n21216), .B2(n14332), .A(n14331), .ZN(n14338) );
  AOI22_X1 U17655 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14336) );
  AOI22_X1 U17656 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14335) );
  AOI22_X1 U17657 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14334) );
  AOI22_X1 U17658 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14333) );
  NAND4_X1 U17659 ( .A1(n14336), .A2(n14335), .A3(n14334), .A4(n14333), .ZN(
        n14337) );
  AOI211_X1 U17660 ( .C1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .C2(n17892), .A(
        n14338), .B(n14337), .ZN(n14339) );
  NAND3_X1 U17661 ( .A1(n14341), .A2(n14340), .A3(n14339), .ZN(n17693) );
  NAND2_X1 U17662 ( .A1(n17694), .A2(n17693), .ZN(n17692) );
  NOR2_X1 U17663 ( .A1(n17688), .A2(n17692), .ZN(n17685) );
  AOI22_X1 U17664 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14352) );
  AOI22_X1 U17665 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14351) );
  INV_X1 U17666 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17925) );
  AOI22_X1 U17667 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14342) );
  OAI21_X1 U17668 ( .B1(n14343), .B2(n17925), .A(n14342), .ZN(n14349) );
  AOI22_X1 U17669 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14347) );
  AOI22_X1 U17670 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14346) );
  AOI22_X1 U17671 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14345) );
  AOI22_X1 U17672 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14344) );
  NAND4_X1 U17673 ( .A1(n14347), .A2(n14346), .A3(n14345), .A4(n14344), .ZN(
        n14348) );
  AOI211_X1 U17674 ( .C1(n17816), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n14349), .B(n14348), .ZN(n14350) );
  NAND3_X1 U17675 ( .A1(n14352), .A2(n14351), .A3(n14350), .ZN(n17684) );
  NAND2_X1 U17676 ( .A1(n17685), .A2(n17684), .ZN(n17683) );
  NOR2_X1 U17677 ( .A1(n17678), .A2(n17683), .ZN(n17960) );
  AOI22_X1 U17678 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n16368), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14363) );
  AOI22_X1 U17679 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n17876), .B1(
        n17816), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14362) );
  AOI22_X1 U17680 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14353) );
  OAI21_X1 U17681 ( .B1(n21139), .B2(n14354), .A(n14353), .ZN(n14360) );
  AOI22_X1 U17682 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14358) );
  AOI22_X1 U17683 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14357) );
  AOI22_X1 U17684 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14356) );
  AOI22_X1 U17685 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14355) );
  NAND4_X1 U17686 ( .A1(n14358), .A2(n14357), .A3(n14356), .A4(n14355), .ZN(
        n14359) );
  AOI211_X1 U17687 ( .C1(n17903), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n14360), .B(n14359), .ZN(n14361) );
  NAND3_X1 U17688 ( .A1(n14363), .A2(n14362), .A3(n14361), .ZN(n17959) );
  NAND2_X1 U17689 ( .A1(n17960), .A2(n17959), .ZN(n17958) );
  XNOR2_X1 U17690 ( .A(n14364), .B(n17958), .ZN(n17957) );
  INV_X1 U17691 ( .A(n17957), .ZN(n14365) );
  INV_X1 U17692 ( .A(n17938), .ZN(n17941) );
  MUX2_X1 U17693 ( .A(n14366), .B(n14365), .S(n17942), .Z(P3_U2673) );
  NAND3_X1 U17694 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19523)
         );
  OAI21_X1 U17695 ( .B1(n19391), .B2(n19531), .A(n17605), .ZN(n16299) );
  NOR2_X1 U17696 ( .A1(n17900), .A2(n16299), .ZN(n18907) );
  INV_X1 U17697 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17275) );
  NOR2_X1 U17698 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19580) );
  AOI21_X1 U17699 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n19580), .ZN(n19429) );
  OR2_X1 U17700 ( .A1(n19549), .A2(n19429), .ZN(n18921) );
  OAI221_X1 U17701 ( .B1(n19523), .B2(n18907), .C1(n19523), .C2(n17275), .A(
        n19002), .ZN(n18915) );
  INV_X1 U17702 ( .A(n18915), .ZN(n18910) );
  NAND2_X1 U17703 ( .A1(n19534), .A2(n19524), .ZN(n19526) );
  INV_X1 U17704 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19587) );
  NAND2_X1 U17705 ( .A1(n19587), .A2(n19524), .ZN(n17267) );
  NAND2_X1 U17706 ( .A1(n19526), .A2(n17267), .ZN(n18908) );
  INV_X1 U17707 ( .A(n18908), .ZN(n19571) );
  INV_X1 U17708 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21087) );
  NOR2_X1 U17709 ( .A1(n21087), .A2(n19534), .ZN(n18546) );
  NOR2_X1 U17710 ( .A1(n19571), .A2(n18546), .ZN(n16260) );
  AOI21_X1 U17711 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n16260), .ZN(n16261) );
  NOR2_X1 U17712 ( .A1(n18910), .A2(n16261), .ZN(n14368) );
  NAND3_X1 U17713 ( .A1(n19587), .A2(n19524), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19164) );
  INV_X1 U17714 ( .A(n19164), .ZN(n19265) );
  NAND2_X1 U17715 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19385), .ZN(n18958) );
  NAND2_X1 U17716 ( .A1(n18958), .A2(n18915), .ZN(n16259) );
  OR2_X1 U17717 ( .A1(n19265), .A2(n16259), .ZN(n14367) );
  MUX2_X1 U17718 ( .A(n14368), .B(n14367), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  OR2_X2 U17719 ( .A1(n14369), .A2(n14370), .ZN(n14371) );
  NAND2_X2 U17720 ( .A1(n14372), .A2(n14371), .ZN(n14820) );
  INV_X1 U17721 ( .A(DATAI_13_), .ZN(n14374) );
  MUX2_X1 U17722 ( .A(n14374), .B(n14373), .S(n14738), .Z(n20763) );
  NAND2_X1 U17723 ( .A1(n16645), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n14375) );
  OAI21_X1 U17724 ( .B1(n14788), .B2(n20763), .A(n14375), .ZN(n14376) );
  AOI21_X1 U17725 ( .B1(n16648), .B2(DATAI_29_), .A(n14376), .ZN(n14380) );
  NAND2_X1 U17726 ( .A1(n14791), .A2(BUF1_REG_29__SCAN_IN), .ZN(n14379) );
  OAI211_X1 U17727 ( .C1(n14820), .C2(n14805), .A(n14380), .B(n14379), .ZN(
        P1_U2875) );
  INV_X1 U17728 ( .A(n14525), .ZN(n14383) );
  INV_X1 U17729 ( .A(n14381), .ZN(n14382) );
  OAI21_X1 U17730 ( .B1(n14383), .B2(n14382), .A(n14500), .ZN(n15026) );
  INV_X1 U17731 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14384) );
  OAI222_X1 U17732 ( .A1(n15026), .A2(n14730), .B1(n14384), .B2(n20721), .C1(
        n14820), .C2(n14731), .ZN(P1_U2843) );
  NAND3_X1 U17733 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .ZN(n14386) );
  NAND2_X1 U17734 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14397) );
  INV_X1 U17735 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20998) );
  NAND3_X1 U17736 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .ZN(n16622) );
  NOR2_X1 U17737 ( .A1(n20998), .A2(n16622), .ZN(n14396) );
  NAND2_X1 U17738 ( .A1(n14396), .A2(n14385), .ZN(n16611) );
  NOR2_X1 U17739 ( .A1(n14397), .A2(n16611), .ZN(n16588) );
  NAND4_X1 U17740 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .A4(n16588), .ZN(n14632) );
  NOR2_X1 U17741 ( .A1(n14386), .A2(n14632), .ZN(n14604) );
  NAND3_X1 U17742 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(P1_REIP_REG_21__SCAN_IN), .ZN(n14557) );
  AND3_X1 U17743 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(P1_REIP_REG_26__SCAN_IN), .ZN(n14399) );
  INV_X1 U17744 ( .A(n14399), .ZN(n14544) );
  NOR2_X1 U17745 ( .A1(n14557), .A2(n14544), .ZN(n14387) );
  NAND2_X1 U17746 ( .A1(n14604), .A2(n14387), .ZN(n14388) );
  NAND2_X1 U17747 ( .A1(n14388), .A2(n20683), .ZN(n14559) );
  AND2_X1 U17748 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14389) );
  NAND2_X1 U17749 ( .A1(n14559), .A2(n14389), .ZN(n14390) );
  NAND2_X1 U17750 ( .A1(n14390), .A2(n20683), .ZN(n14508) );
  INV_X1 U17751 ( .A(n14508), .ZN(n14531) );
  INV_X1 U17752 ( .A(n14391), .ZN(n14822) );
  OAI22_X1 U17753 ( .A1(n14392), .A2(n16596), .B1(n20703), .B2(n14822), .ZN(
        n14393) );
  AOI21_X1 U17754 ( .B1(n20684), .B2(P1_EBX_REG_29__SCAN_IN), .A(n14393), .ZN(
        n14394) );
  OAI21_X1 U17755 ( .B1(n15026), .B2(n20666), .A(n14394), .ZN(n14395) );
  AOI21_X1 U17756 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14531), .A(n14395), 
        .ZN(n14402) );
  INV_X1 U17757 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21005) );
  NAND3_X1 U17758 ( .A1(n16593), .A2(P1_REIP_REG_15__SCAN_IN), .A3(
        P1_REIP_REG_16__SCAN_IN), .ZN(n14651) );
  NOR2_X2 U17759 ( .A1(n21005), .A2(n14651), .ZN(n16578) );
  AND3_X1 U17760 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n14398) );
  NAND2_X1 U17761 ( .A1(n14399), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14400) );
  NOR2_X2 U17762 ( .A1(n14563), .A2(n14400), .ZN(n14522) );
  INV_X1 U17763 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21026) );
  NAND3_X1 U17764 ( .A1(n14522), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n21026), 
        .ZN(n14401) );
  OAI211_X1 U17765 ( .C1(n14820), .C2(n16601), .A(n14402), .B(n14401), .ZN(
        P1_U2811) );
  INV_X1 U17766 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17169) );
  NAND3_X1 U17767 ( .A1(n14515), .A2(n14403), .A3(n14802), .ZN(n14405) );
  AOI22_X1 U17768 ( .A1(n16648), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n16645), .ZN(n14404) );
  OAI211_X1 U17769 ( .C1(n16652), .C2(n17169), .A(n14405), .B(n14404), .ZN(
        P1_U2873) );
  INV_X1 U17770 ( .A(n14408), .ZN(n14409) );
  NAND2_X1 U17771 ( .A1(n10773), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14411) );
  XNOR2_X1 U17772 ( .A(n14413), .B(n14411), .ZN(n15355) );
  AOI21_X1 U17773 ( .B1(n15355), .B2(n10350), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15665) );
  AND2_X1 U17774 ( .A1(n10350), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14412) );
  NAND2_X1 U17775 ( .A1(n15355), .A2(n14412), .ZN(n15663) );
  OAI21_X1 U17776 ( .B1(n14413), .B2(P2_EBX_REG_30__SCAN_IN), .A(n10773), .ZN(
        n14415) );
  NAND2_X1 U17777 ( .A1(n14415), .A2(n14414), .ZN(n15339) );
  NOR2_X1 U17778 ( .A1(n15339), .A2(n10362), .ZN(n14416) );
  XOR2_X1 U17779 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n14416), .Z(
        n14417) );
  XNOR2_X1 U17780 ( .A(n14418), .B(n14417), .ZN(n14477) );
  INV_X1 U17781 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n14463) );
  INV_X1 U17782 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14428) );
  OAI22_X1 U17783 ( .A1(n9609), .A2(n14463), .B1(n20495), .B2(n14428), .ZN(
        n14423) );
  AOI21_X1 U17784 ( .B1(n14424), .B2(P2_EBX_REG_31__SCAN_IN), .A(n14423), .ZN(
        n14425) );
  OAI21_X1 U17785 ( .B1(n14426), .B2(n14419), .A(n14425), .ZN(n14427) );
  NAND2_X1 U17786 ( .A1(n19903), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14467) );
  OAI21_X1 U17787 ( .B1(n16950), .B2(n14428), .A(n14467), .ZN(n14429) );
  AOI21_X1 U17788 ( .B1(n14430), .B2(n16942), .A(n14429), .ZN(n14431) );
  OAI21_X1 U17789 ( .B1(n16899), .B2(n13859), .A(n14431), .ZN(n14432) );
  AOI21_X1 U17790 ( .B1(n14475), .B2(n15933), .A(n14432), .ZN(n14433) );
  OAI21_X1 U17791 ( .B1(n14477), .B2(n16957), .A(n14433), .ZN(P2_U2983) );
  NOR2_X1 U17792 ( .A1(n16950), .A2(n12800), .ZN(n14438) );
  OAI21_X1 U17793 ( .B1(n14436), .B2(n14435), .A(n14434), .ZN(n19927) );
  NAND2_X1 U17794 ( .A1(n19903), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19922) );
  OAI21_X1 U17795 ( .B1(n16955), .B2(n19927), .A(n19922), .ZN(n14437) );
  AOI211_X1 U17796 ( .C1(n14439), .C2(n16942), .A(n14438), .B(n14437), .ZN(
        n14443) );
  XOR2_X1 U17797 ( .A(n14441), .B(n14440), .Z(n19921) );
  NAND2_X1 U17798 ( .A1(n19921), .A2(n15927), .ZN(n14442) );
  OAI211_X1 U17799 ( .C1(n13062), .C2(n13859), .A(n14443), .B(n14442), .ZN(
        P2_U3012) );
  INV_X1 U17800 ( .A(n15169), .ZN(n14444) );
  OAI22_X1 U17801 ( .A1(n14445), .A2(n14444), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11531), .ZN(n16507) );
  OAI22_X1 U17802 ( .A1(n20962), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15186), .ZN(n14446) );
  AOI21_X1 U17803 ( .B1(n16507), .B2(n20632), .A(n14446), .ZN(n14452) );
  INV_X1 U17804 ( .A(n14447), .ZN(n14448) );
  AOI21_X1 U17805 ( .B1(n16503), .B2(n14967), .A(n14448), .ZN(n16839) );
  OAI21_X1 U17806 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20905), .A(n16839), 
        .ZN(n16842) );
  INV_X1 U17807 ( .A(n16842), .ZN(n14451) );
  AOI21_X1 U17808 ( .B1(n16508), .B2(n20632), .A(n14451), .ZN(n14450) );
  OAI22_X1 U17809 ( .A1(n14452), .A2(n14451), .B1(n14450), .B2(n14449), .ZN(
        P1_U3474) );
  AND2_X1 U17810 ( .A1(n16497), .A2(n21106), .ZN(n14457) );
  NAND2_X1 U17811 ( .A1(n16497), .A2(n16027), .ZN(n14456) );
  NAND2_X1 U17812 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16056) );
  INV_X1 U17813 ( .A(n16056), .ZN(n16069) );
  AND2_X1 U17814 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n16069), .ZN(
        n14453) );
  NAND2_X1 U17815 ( .A1(n16055), .A2(n14453), .ZN(n14472) );
  NOR2_X1 U17816 ( .A1(n10683), .A2(n10835), .ZN(n17000) );
  NAND2_X1 U17817 ( .A1(n14454), .A2(n14455), .ZN(n14470) );
  NOR2_X1 U17818 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14470), .ZN(
        n16197) );
  OAI21_X1 U17819 ( .B1(n14455), .B2(n17022), .A(n19905), .ZN(n16199) );
  NOR2_X1 U17820 ( .A1(n16197), .A2(n16199), .ZN(n17001) );
  OAI21_X1 U17821 ( .B1(n17022), .B2(n17000), .A(n17001), .ZN(n16166) );
  AOI21_X1 U17822 ( .B1(n16497), .B2(n14472), .A(n16166), .ZN(n16057) );
  NAND2_X1 U17823 ( .A1(n14456), .A2(n16057), .ZN(n16021) );
  NOR2_X1 U17824 ( .A1(n15999), .A2(n15998), .ZN(n15997) );
  INV_X1 U17825 ( .A(n15997), .ZN(n14458) );
  AND2_X1 U17826 ( .A1(n16497), .A2(n14458), .ZN(n14459) );
  NOR2_X1 U17827 ( .A1(n16007), .A2(n14459), .ZN(n15979) );
  NAND3_X1 U17828 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15943) );
  NAND2_X1 U17829 ( .A1(n16497), .A2(n15943), .ZN(n14460) );
  AND2_X1 U17830 ( .A1(n15979), .A2(n14460), .ZN(n15942) );
  OAI21_X1 U17831 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17022), .A(
        n15942), .ZN(n14469) );
  AOI22_X1 U17832 ( .A1(n14461), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12652), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14462) );
  OAI21_X1 U17833 ( .B1(n14464), .B2(n14463), .A(n14462), .ZN(n14465) );
  XNOR2_X1 U17834 ( .A(n14466), .B(n14465), .ZN(n19797) );
  OAI21_X1 U17835 ( .B1(n19797), .B2(n19928), .A(n14467), .ZN(n14468) );
  AOI21_X1 U17836 ( .B1(n14469), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14468), .ZN(n14473) );
  NAND2_X1 U17837 ( .A1(n16998), .A2(n17000), .ZN(n16149) );
  NOR3_X1 U17838 ( .A1(n16026), .A2(n21106), .A3(n16027), .ZN(n15996) );
  NAND2_X1 U17839 ( .A1(n15996), .A2(n15997), .ZN(n15971) );
  OAI21_X1 U17840 ( .B1(n14477), .B2(n17009), .A(n14476), .ZN(P2_U3015) );
  NAND2_X1 U17841 ( .A1(n14478), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16220) );
  OAI21_X1 U17842 ( .B1(n19753), .B2(n14480), .A(n14479), .ZN(n16219) );
  INV_X1 U17843 ( .A(n16219), .ZN(n14481) );
  NOR2_X1 U17844 ( .A1(n16220), .A2(n14481), .ZN(n14497) );
  NOR2_X1 U17845 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14494) );
  INV_X1 U17846 ( .A(n14482), .ZN(n14483) );
  NAND2_X1 U17847 ( .A1(n17033), .A2(n14483), .ZN(n17026) );
  NAND2_X1 U17848 ( .A1(n14484), .A2(n12772), .ZN(n14485) );
  NAND2_X1 U17849 ( .A1(n14485), .A2(n14489), .ZN(n17028) );
  NOR2_X1 U17850 ( .A1(n14486), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14488) );
  NOR2_X1 U17851 ( .A1(n17028), .A2(n14488), .ZN(n14492) );
  NAND2_X1 U17852 ( .A1(n14487), .A2(n17054), .ZN(n17023) );
  INV_X1 U17853 ( .A(n17028), .ZN(n14491) );
  INV_X1 U17854 ( .A(n14488), .ZN(n17027) );
  NAND2_X1 U17855 ( .A1(n14489), .A2(n17027), .ZN(n14490) );
  OAI22_X1 U17856 ( .A1(n14492), .A2(n17023), .B1(n14491), .B2(n14490), .ZN(
        n14493) );
  OAI21_X1 U17857 ( .B1(n14494), .B2(n17026), .A(n14493), .ZN(n14495) );
  OAI22_X1 U17858 ( .A1(n20054), .A2(n20569), .B1(n20568), .B2(n17042), .ZN(
        n14496) );
  OAI21_X1 U17859 ( .B1(n14497), .B2(n14496), .A(n20573), .ZN(n14498) );
  OAI21_X1 U17860 ( .B1(n20573), .B2(n14499), .A(n14498), .ZN(P2_U3599) );
  MUX2_X1 U17861 ( .A(n14502), .B(n14501), .S(n14500), .Z(n14505) );
  AOI22_X1 U17862 ( .A1(n14503), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n9612), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14504) );
  NAND2_X1 U17863 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14506) );
  NAND2_X1 U17864 ( .A1(n20683), .A2(n14506), .ZN(n14507) );
  NAND2_X1 U17865 ( .A1(n14508), .A2(n14507), .ZN(n14519) );
  OAI22_X1 U17866 ( .A1(n20707), .A2(n14668), .B1(n14509), .B2(n16596), .ZN(
        n14510) );
  AOI21_X1 U17867 ( .B1(n14519), .B2(P1_REIP_REG_31__SCAN_IN), .A(n14510), 
        .ZN(n14513) );
  AND2_X1 U17868 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14511) );
  AND2_X1 U17869 ( .A1(n14522), .A2(n14511), .ZN(n14520) );
  NAND3_X1 U17870 ( .A1(n14520), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n21030), 
        .ZN(n14512) );
  OAI211_X1 U17871 ( .C1(n14975), .C2(n20666), .A(n14513), .B(n14512), .ZN(
        n14514) );
  AOI21_X1 U17872 ( .B1(n14515), .B2(n20676), .A(n14514), .ZN(n14516) );
  INV_X1 U17873 ( .A(n14516), .ZN(P1_U2809) );
  OAI22_X1 U17874 ( .A1(n14517), .A2(n16596), .B1(n20703), .B2(n14812), .ZN(
        n14518) );
  OAI21_X1 U17875 ( .B1(n14520), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14519), 
        .ZN(n14521) );
  INV_X1 U17876 ( .A(n14522), .ZN(n14534) );
  AOI21_X1 U17877 ( .B1(n14524), .B2(n14523), .A(n14369), .ZN(n14834) );
  NAND2_X1 U17878 ( .A1(n14834), .A2(n20676), .ZN(n14533) );
  OAI21_X1 U17879 ( .B1(n14539), .B2(n14526), .A(n14525), .ZN(n15036) );
  OAI22_X1 U17880 ( .A1(n14527), .A2(n16596), .B1(n20703), .B2(n14832), .ZN(
        n14528) );
  AOI21_X1 U17881 ( .B1(n20684), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14528), .ZN(
        n14529) );
  OAI21_X1 U17882 ( .B1(n15036), .B2(n20666), .A(n14529), .ZN(n14530) );
  AOI21_X1 U17883 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14531), .A(n14530), 
        .ZN(n14532) );
  OAI211_X1 U17884 ( .C1(P1_REIP_REG_28__SCAN_IN), .C2(n14534), .A(n14533), 
        .B(n14532), .ZN(P1_U2812) );
  OAI21_X1 U17885 ( .B1(n14535), .B2(n14536), .A(n14523), .ZN(n14840) );
  AND2_X1 U17886 ( .A1(n14551), .A2(n14537), .ZN(n14538) );
  NOR2_X1 U17887 ( .A1(n14539), .A2(n14538), .ZN(n15053) );
  INV_X1 U17888 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21019) );
  NOR2_X1 U17889 ( .A1(n14559), .A2(n21019), .ZN(n14543) );
  INV_X1 U17890 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14541) );
  AOI22_X1 U17891 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20705), .B1(
        n20687), .B2(n14841), .ZN(n14540) );
  OAI21_X1 U17892 ( .B1(n20707), .B2(n14541), .A(n14540), .ZN(n14542) );
  AOI211_X1 U17893 ( .C1(n15053), .C2(n20700), .A(n14543), .B(n14542), .ZN(
        n14546) );
  OAI211_X1 U17894 ( .C1(n14840), .C2(n16601), .A(n14546), .B(n14545), .ZN(
        P1_U2813) );
  AOI21_X1 U17896 ( .B1(n14549), .B2(n14548), .A(n14535), .ZN(n14855) );
  INV_X1 U17897 ( .A(n14855), .ZN(n14752) );
  OAI22_X1 U17898 ( .A1(n14550), .A2(n16596), .B1(n20703), .B2(n14853), .ZN(
        n14556) );
  INV_X1 U17899 ( .A(n14551), .ZN(n14552) );
  AOI21_X1 U17900 ( .B1(n14553), .B2(n14569), .A(n14552), .ZN(n15063) );
  INV_X1 U17901 ( .A(n15063), .ZN(n14554) );
  NOR2_X1 U17902 ( .A1(n14554), .A2(n20666), .ZN(n14555) );
  AOI211_X1 U17903 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n20684), .A(n14556), .B(
        n14555), .ZN(n14562) );
  NOR2_X1 U17904 ( .A1(n14563), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14585) );
  INV_X1 U17905 ( .A(n14557), .ZN(n14558) );
  AOI21_X1 U17906 ( .B1(n14604), .B2(n14558), .A(n16587), .ZN(n14598) );
  INV_X1 U17907 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14859) );
  NOR3_X1 U17908 ( .A1(n14585), .A2(n14598), .A3(n14859), .ZN(n14576) );
  INV_X1 U17909 ( .A(n14559), .ZN(n14560) );
  OAI21_X1 U17910 ( .B1(n14576), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14560), 
        .ZN(n14561) );
  OAI211_X1 U17911 ( .C1(n14752), .C2(n16601), .A(n14562), .B(n14561), .ZN(
        P1_U2814) );
  INV_X1 U17912 ( .A(n14563), .ZN(n14564) );
  AOI21_X1 U17913 ( .B1(n14564), .B2(P1_REIP_REG_24__SCAN_IN), .A(
        P1_REIP_REG_25__SCAN_IN), .ZN(n14575) );
  OAI21_X1 U17914 ( .B1(n14565), .B2(n14566), .A(n14548), .ZN(n14673) );
  INV_X1 U17915 ( .A(n14673), .ZN(n14863) );
  NAND2_X1 U17916 ( .A1(n14863), .A2(n20676), .ZN(n14574) );
  INV_X1 U17917 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14568) );
  INV_X1 U17918 ( .A(n14567), .ZN(n14861) );
  OAI22_X1 U17919 ( .A1(n14568), .A2(n16596), .B1(n20703), .B2(n14861), .ZN(
        n14572) );
  OAI21_X1 U17920 ( .B1(n14579), .B2(n14570), .A(n14569), .ZN(n15066) );
  NOR2_X1 U17921 ( .A1(n15066), .A2(n20666), .ZN(n14571) );
  AOI211_X1 U17922 ( .C1(n20684), .C2(P1_EBX_REG_25__SCAN_IN), .A(n14572), .B(
        n14571), .ZN(n14573) );
  OAI211_X1 U17923 ( .C1(n14576), .C2(n14575), .A(n14574), .B(n14573), .ZN(
        P1_U2815) );
  AOI21_X1 U17924 ( .B1(n14578), .B2(n14577), .A(n14565), .ZN(n14872) );
  INV_X1 U17925 ( .A(n14872), .ZN(n14675) );
  INV_X1 U17926 ( .A(n14579), .ZN(n14580) );
  OAI21_X1 U17927 ( .B1(n14592), .B2(n14581), .A(n14580), .ZN(n15075) );
  OAI22_X1 U17928 ( .A1(n14582), .A2(n16596), .B1(n20703), .B2(n14870), .ZN(
        n14583) );
  AOI21_X1 U17929 ( .B1(n20684), .B2(P1_EBX_REG_24__SCAN_IN), .A(n14583), .ZN(
        n14584) );
  OAI21_X1 U17930 ( .B1(n15075), .B2(n20666), .A(n14584), .ZN(n14586) );
  AOI211_X1 U17931 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n14598), .A(n14586), 
        .B(n14585), .ZN(n14587) );
  OAI21_X1 U17932 ( .B1(n14675), .B2(n16601), .A(n14587), .ZN(P1_U2816) );
  OAI21_X1 U17933 ( .B1(n14588), .B2(n14589), .A(n14577), .ZN(n14761) );
  INV_X1 U17934 ( .A(n14590), .ZN(n14878) );
  OAI22_X1 U17935 ( .A1(n14591), .A2(n16596), .B1(n20703), .B2(n14878), .ZN(
        n14596) );
  AOI21_X1 U17936 ( .B1(n14593), .B2(n9652), .A(n14592), .ZN(n15092) );
  INV_X1 U17937 ( .A(n15092), .ZN(n14594) );
  NOR2_X1 U17938 ( .A1(n14594), .A2(n20666), .ZN(n14595) );
  AOI211_X1 U17939 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n20684), .A(n14596), .B(
        n14595), .ZN(n14601) );
  NAND2_X1 U17940 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14597) );
  NOR2_X1 U17941 ( .A1(n14623), .A2(n14597), .ZN(n14599) );
  OAI21_X1 U17942 ( .B1(n14599), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14598), 
        .ZN(n14600) );
  OAI211_X1 U17943 ( .C1(n14761), .C2(n16601), .A(n14601), .B(n14600), .ZN(
        P1_U2817) );
  XNOR2_X1 U17944 ( .A(P1_REIP_REG_21__SCAN_IN), .B(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14613) );
  INV_X1 U17945 ( .A(n14602), .ZN(n14615) );
  AOI21_X1 U17946 ( .B1(n14603), .B2(n14615), .A(n14588), .ZN(n14888) );
  NAND2_X1 U17947 ( .A1(n14888), .A2(n20676), .ZN(n14612) );
  OR2_X1 U17948 ( .A1(n14604), .A2(n16587), .ZN(n16568) );
  INV_X1 U17949 ( .A(n16568), .ZN(n14626) );
  NAND2_X1 U17950 ( .A1(n14617), .A2(n14605), .ZN(n14606) );
  NAND2_X1 U17951 ( .A1(n9652), .A2(n14606), .ZN(n16704) );
  INV_X1 U17952 ( .A(n14886), .ZN(n14607) );
  AOI22_X1 U17953 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20705), .B1(
        n20687), .B2(n14607), .ZN(n14609) );
  NAND2_X1 U17954 ( .A1(n20684), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n14608) );
  OAI211_X1 U17955 ( .C1(n16704), .C2(n20666), .A(n14609), .B(n14608), .ZN(
        n14610) );
  AOI21_X1 U17956 ( .B1(n14626), .B2(P1_REIP_REG_22__SCAN_IN), .A(n14610), 
        .ZN(n14611) );
  OAI211_X1 U17957 ( .C1(n14623), .C2(n14613), .A(n14612), .B(n14611), .ZN(
        P1_U2818) );
  AOI21_X1 U17958 ( .B1(n14616), .B2(n14614), .A(n14602), .ZN(n14896) );
  INV_X1 U17959 ( .A(n14896), .ZN(n14776) );
  OAI21_X1 U17960 ( .B1(n14684), .B2(n14618), .A(n14617), .ZN(n15095) );
  INV_X1 U17961 ( .A(n14619), .ZN(n14894) );
  OAI22_X1 U17962 ( .A1(n14620), .A2(n16596), .B1(n20703), .B2(n14894), .ZN(
        n14621) );
  AOI21_X1 U17963 ( .B1(n20684), .B2(P1_EBX_REG_21__SCAN_IN), .A(n14621), .ZN(
        n14622) );
  OAI21_X1 U17964 ( .B1(n15095), .B2(n20666), .A(n14622), .ZN(n14625) );
  NOR2_X1 U17965 ( .A1(n14623), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14624) );
  AOI211_X1 U17966 ( .C1(n14626), .C2(P1_REIP_REG_21__SCAN_IN), .A(n14625), 
        .B(n14624), .ZN(n14627) );
  OAI21_X1 U17967 ( .B1(n14776), .B2(n16601), .A(n14627), .ZN(P1_U2819) );
  AOI21_X1 U17969 ( .B1(n14631), .B2(n14628), .A(n14630), .ZN(n14911) );
  INV_X1 U17970 ( .A(n14911), .ZN(n14781) );
  INV_X1 U17971 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21009) );
  INV_X1 U17972 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21007) );
  NOR2_X1 U17973 ( .A1(n21009), .A2(n21007), .ZN(n16566) );
  AOI21_X1 U17974 ( .B1(n21009), .B2(n21007), .A(n16566), .ZN(n14640) );
  NAND2_X1 U17975 ( .A1(n20683), .A2(n14632), .ZN(n16582) );
  AOI22_X1 U17976 ( .A1(n20684), .A2(P1_EBX_REG_19__SCAN_IN), .B1(n20687), 
        .B2(n14907), .ZN(n14633) );
  OAI21_X1 U17977 ( .B1(n21009), .B2(n16582), .A(n14633), .ZN(n14639) );
  INV_X1 U17978 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14637) );
  INV_X1 U17979 ( .A(n14683), .ZN(n14634) );
  AOI21_X1 U17980 ( .B1(n14635), .B2(n14694), .A(n14634), .ZN(n16713) );
  NAND2_X1 U17981 ( .A1(n16713), .A2(n20700), .ZN(n14636) );
  OAI211_X1 U17982 ( .C1(n16596), .C2(n14637), .A(n14636), .B(n20702), .ZN(
        n14638) );
  AOI211_X1 U17983 ( .C1(n16578), .C2(n14640), .A(n14639), .B(n14638), .ZN(
        n14641) );
  OAI21_X1 U17984 ( .B1(n14781), .B2(n16601), .A(n14641), .ZN(P1_U2821) );
  AOI21_X1 U17985 ( .B1(n14644), .B2(n14642), .A(n14643), .ZN(n14932) );
  INV_X1 U17986 ( .A(n14932), .ZN(n14794) );
  OR2_X1 U17987 ( .A1(n14704), .A2(n14645), .ZN(n14646) );
  AND2_X1 U17988 ( .A1(n14692), .A2(n14646), .ZN(n16732) );
  INV_X1 U17989 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14647) );
  OAI22_X1 U17990 ( .A1(n20707), .A2(n14647), .B1(n14930), .B2(n20703), .ZN(
        n14648) );
  INV_X1 U17991 ( .A(n14648), .ZN(n14649) );
  OAI211_X1 U17992 ( .C1(n16596), .C2(n14650), .A(n14649), .B(n20702), .ZN(
        n14653) );
  AOI21_X1 U17993 ( .B1(n21005), .B2(n14651), .A(n16582), .ZN(n14652) );
  AOI211_X1 U17994 ( .C1(n16732), .C2(n20700), .A(n14653), .B(n14652), .ZN(
        n14654) );
  OAI21_X1 U17995 ( .B1(n14794), .B2(n16601), .A(n14654), .ZN(P1_U2823) );
  INV_X1 U17996 ( .A(n14655), .ZN(n20709) );
  NAND2_X1 U17997 ( .A1(n14656), .A2(n20698), .ZN(n14661) );
  INV_X1 U17998 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14658) );
  OAI22_X1 U17999 ( .A1(n14658), .A2(n16596), .B1(n20703), .B2(n14657), .ZN(
        n14659) );
  AOI21_X1 U18000 ( .B1(n20684), .B2(P1_EBX_REG_2__SCAN_IN), .A(n14659), .ZN(
        n14660) );
  OAI211_X1 U18001 ( .C1(n20814), .C2(n14662), .A(n14661), .B(n14660), .ZN(
        n14665) );
  OAI22_X1 U18002 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n14663), .B1(n20666), 
        .B2(n20815), .ZN(n14664) );
  AOI211_X1 U18003 ( .C1(n14666), .C2(n20709), .A(n14665), .B(n14664), .ZN(
        n14667) );
  INV_X1 U18004 ( .A(n14667), .ZN(P1_U2838) );
  OAI22_X1 U18005 ( .A1(n14975), .A2(n14730), .B1(n20721), .B2(n14668), .ZN(
        P1_U2841) );
  INV_X1 U18006 ( .A(n14834), .ZN(n14743) );
  INV_X1 U18007 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14669) );
  OAI222_X1 U18008 ( .A1(n14743), .A2(n14731), .B1(n14669), .B2(n20721), .C1(
        n15036), .C2(n14730), .ZN(P1_U2844) );
  AOI22_X1 U18009 ( .A1(n15053), .A2(n20717), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14715), .ZN(n14670) );
  OAI21_X1 U18010 ( .B1(n14840), .B2(n14731), .A(n14670), .ZN(P1_U2845) );
  AOI22_X1 U18011 ( .A1(n15063), .A2(n20717), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14715), .ZN(n14671) );
  OAI21_X1 U18012 ( .B1(n14752), .B2(n14731), .A(n14671), .ZN(P1_U2846) );
  INV_X1 U18013 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14672) );
  OAI222_X1 U18014 ( .A1(n14673), .A2(n14731), .B1(n14672), .B2(n20721), .C1(
        n15066), .C2(n14730), .ZN(P1_U2847) );
  INV_X1 U18015 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14674) );
  OAI222_X1 U18016 ( .A1(n14675), .A2(n14731), .B1(n14674), .B2(n20721), .C1(
        n15075), .C2(n14730), .ZN(P1_U2848) );
  AOI22_X1 U18017 ( .A1(n15092), .A2(n20717), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14715), .ZN(n14676) );
  OAI21_X1 U18018 ( .B1(n14761), .B2(n14731), .A(n14676), .ZN(P1_U2849) );
  INV_X1 U18019 ( .A(n14888), .ZN(n14678) );
  INV_X1 U18020 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14677) );
  OAI222_X1 U18021 ( .A1(n14678), .A2(n14731), .B1(n14677), .B2(n20721), .C1(
        n16704), .C2(n14730), .ZN(P1_U2850) );
  INV_X1 U18022 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14679) );
  OAI222_X1 U18023 ( .A1(n14776), .A2(n14731), .B1(n14679), .B2(n20721), .C1(
        n15095), .C2(n14730), .ZN(P1_U2851) );
  OR2_X1 U18024 ( .A1(n14630), .A2(n14680), .ZN(n14681) );
  AND2_X1 U18025 ( .A1(n14681), .A2(n14614), .ZN(n16642) );
  INV_X1 U18026 ( .A(n16642), .ZN(n14687) );
  INV_X1 U18027 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14686) );
  AND2_X1 U18028 ( .A1(n14683), .A2(n14682), .ZN(n14685) );
  OR2_X1 U18029 ( .A1(n14685), .A2(n14684), .ZN(n16567) );
  OAI222_X1 U18030 ( .A1(n14687), .A2(n14699), .B1(n14686), .B2(n20721), .C1(
        n16567), .C2(n14730), .ZN(P1_U2852) );
  AOI22_X1 U18031 ( .A1(n16713), .A2(n20717), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14715), .ZN(n14688) );
  OAI21_X1 U18032 ( .B1(n14781), .B2(n14699), .A(n14688), .ZN(P1_U2853) );
  NAND2_X1 U18033 ( .A1(n10107), .A2(n14689), .ZN(n14690) );
  AND2_X1 U18034 ( .A1(n14628), .A2(n14690), .ZN(n16579) );
  INV_X1 U18035 ( .A(n16579), .ZN(n14920) );
  NAND2_X1 U18036 ( .A1(n14692), .A2(n14691), .ZN(n14693) );
  NAND2_X1 U18037 ( .A1(n14694), .A2(n14693), .ZN(n16724) );
  INV_X1 U18038 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14695) );
  OAI22_X1 U18039 ( .A1(n16724), .A2(n14730), .B1(n14695), .B2(n20721), .ZN(
        n14696) );
  INV_X1 U18040 ( .A(n14696), .ZN(n14697) );
  OAI21_X1 U18041 ( .B1(n14920), .B2(n14699), .A(n14697), .ZN(P1_U2854) );
  AOI22_X1 U18042 ( .A1(n16732), .A2(n20717), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14715), .ZN(n14698) );
  OAI21_X1 U18043 ( .B1(n14794), .B2(n14699), .A(n14698), .ZN(P1_U2855) );
  OAI21_X1 U18044 ( .B1(n14700), .B2(n14701), .A(n14642), .ZN(n16586) );
  NOR2_X1 U18045 ( .A1(n14713), .A2(n14702), .ZN(n14703) );
  OR2_X1 U18046 ( .A1(n14704), .A2(n14703), .ZN(n16748) );
  INV_X1 U18047 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14705) );
  OAI22_X1 U18048 ( .A1(n16748), .A2(n14730), .B1(n14705), .B2(n20721), .ZN(
        n14706) );
  INV_X1 U18049 ( .A(n14706), .ZN(n14707) );
  OAI21_X1 U18050 ( .B1(n16586), .B2(n14731), .A(n14707), .ZN(P1_U2856) );
  AND2_X1 U18051 ( .A1(n14796), .A2(n14709), .ZN(n14710) );
  OR2_X1 U18052 ( .A1(n14710), .A2(n14700), .ZN(n21064) );
  INV_X1 U18053 ( .A(n15128), .ZN(n14712) );
  AOI21_X1 U18054 ( .B1(n14712), .B2(n15127), .A(n14711), .ZN(n14714) );
  NOR2_X1 U18055 ( .A1(n14714), .A2(n14713), .ZN(n16749) );
  AOI22_X1 U18056 ( .A1(n16749), .A2(n20717), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14715), .ZN(n14716) );
  OAI21_X1 U18057 ( .B1(n21064), .B2(n14731), .A(n14716), .ZN(P1_U2857) );
  INV_X1 U18058 ( .A(n14718), .ZN(n14719) );
  AOI21_X1 U18059 ( .B1(n14720), .B2(n14717), .A(n14719), .ZN(n16617) );
  INV_X1 U18060 ( .A(n16617), .ZN(n14801) );
  INV_X1 U18061 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14725) );
  INV_X1 U18062 ( .A(n14721), .ZN(n14728) );
  INV_X1 U18063 ( .A(n14722), .ZN(n14723) );
  OAI21_X1 U18064 ( .B1(n14729), .B2(n14728), .A(n14723), .ZN(n14724) );
  NAND2_X1 U18065 ( .A1(n14724), .A2(n15128), .ZN(n16758) );
  OAI222_X1 U18066 ( .A1(n14801), .A2(n14731), .B1(n20721), .B2(n14725), .C1(
        n16758), .C2(n14730), .ZN(P1_U2859) );
  OAI21_X1 U18067 ( .B1(n14727), .B2(n14726), .A(n14717), .ZN(n16620) );
  INV_X1 U18068 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16624) );
  XNOR2_X1 U18069 ( .A(n14729), .B(n14728), .ZN(n16625) );
  OAI222_X1 U18070 ( .A1(n14731), .A2(n16620), .B1(n20721), .B2(n16624), .C1(
        n14730), .C2(n16625), .ZN(P1_U2860) );
  INV_X1 U18071 ( .A(DATAI_14_), .ZN(n14733) );
  INV_X1 U18072 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14732) );
  MUX2_X1 U18073 ( .A(n14733), .B(n14732), .S(n14738), .Z(n20766) );
  NAND2_X1 U18074 ( .A1(n16645), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n14734) );
  OAI21_X1 U18075 ( .B1(n14788), .B2(n20766), .A(n14734), .ZN(n14735) );
  AOI21_X1 U18076 ( .B1(n16648), .B2(DATAI_30_), .A(n14735), .ZN(n14737) );
  NAND2_X1 U18077 ( .A1(n14791), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14736) );
  OAI211_X1 U18078 ( .C1(n14815), .C2(n14805), .A(n14737), .B(n14736), .ZN(
        P1_U2874) );
  INV_X1 U18079 ( .A(DATAI_12_), .ZN(n21158) );
  INV_X1 U18080 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n17200) );
  MUX2_X1 U18081 ( .A(n21158), .B(n17200), .S(n14738), .Z(n20760) );
  NAND2_X1 U18082 ( .A1(n16645), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n14739) );
  OAI21_X1 U18083 ( .B1(n14788), .B2(n20760), .A(n14739), .ZN(n14740) );
  AOI21_X1 U18084 ( .B1(n16648), .B2(DATAI_28_), .A(n14740), .ZN(n14742) );
  NAND2_X1 U18085 ( .A1(n14791), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14741) );
  OAI211_X1 U18086 ( .C1(n14743), .C2(n14805), .A(n14742), .B(n14741), .ZN(
        P1_U2876) );
  NAND2_X1 U18087 ( .A1(n16645), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n14744) );
  OAI21_X1 U18088 ( .B1(n14788), .B2(n20757), .A(n14744), .ZN(n14745) );
  AOI21_X1 U18089 ( .B1(n16648), .B2(DATAI_27_), .A(n14745), .ZN(n14747) );
  NAND2_X1 U18090 ( .A1(n14791), .A2(BUF1_REG_27__SCAN_IN), .ZN(n14746) );
  OAI211_X1 U18091 ( .C1(n14840), .C2(n14805), .A(n14747), .B(n14746), .ZN(
        P1_U2877) );
  NAND2_X1 U18092 ( .A1(n16645), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n14748) );
  OAI21_X1 U18093 ( .B1(n14788), .B2(n20754), .A(n14748), .ZN(n14749) );
  AOI21_X1 U18094 ( .B1(n16648), .B2(DATAI_26_), .A(n14749), .ZN(n14751) );
  NAND2_X1 U18095 ( .A1(n14791), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14750) );
  OAI211_X1 U18096 ( .C1(n14752), .C2(n14805), .A(n14751), .B(n14750), .ZN(
        P1_U2878) );
  INV_X1 U18097 ( .A(n14805), .ZN(n16649) );
  NAND2_X1 U18098 ( .A1(n14863), .A2(n16649), .ZN(n14756) );
  AOI22_X1 U18099 ( .A1(n16647), .A2(n20752), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n16645), .ZN(n14755) );
  NAND2_X1 U18100 ( .A1(n14791), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14754) );
  NAND2_X1 U18101 ( .A1(n16648), .A2(DATAI_25_), .ZN(n14753) );
  NAND4_X1 U18102 ( .A1(n14756), .A2(n14755), .A3(n14754), .A4(n14753), .ZN(
        P1_U2879) );
  NAND2_X1 U18103 ( .A1(n14872), .A2(n16649), .ZN(n14760) );
  AOI22_X1 U18104 ( .A1(n16647), .A2(n20750), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n16645), .ZN(n14759) );
  NAND2_X1 U18105 ( .A1(n14791), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14758) );
  NAND2_X1 U18106 ( .A1(n16648), .A2(DATAI_24_), .ZN(n14757) );
  NAND4_X1 U18107 ( .A1(n14760), .A2(n14759), .A3(n14758), .A4(n14757), .ZN(
        P1_U2880) );
  INV_X1 U18108 ( .A(n14761), .ZN(n14880) );
  NAND2_X1 U18109 ( .A1(n14880), .A2(n16649), .ZN(n14766) );
  AOI22_X1 U18110 ( .A1(n16647), .A2(n14762), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n16645), .ZN(n14765) );
  NAND2_X1 U18111 ( .A1(n14791), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14764) );
  NAND2_X1 U18112 ( .A1(n16648), .A2(DATAI_23_), .ZN(n14763) );
  NAND4_X1 U18113 ( .A1(n14766), .A2(n14765), .A3(n14764), .A4(n14763), .ZN(
        P1_U2881) );
  NAND2_X1 U18114 ( .A1(n14888), .A2(n16649), .ZN(n14771) );
  AOI22_X1 U18115 ( .A1(n16647), .A2(n14767), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n16645), .ZN(n14770) );
  NAND2_X1 U18116 ( .A1(n14791), .A2(BUF1_REG_22__SCAN_IN), .ZN(n14769) );
  NAND2_X1 U18117 ( .A1(n16648), .A2(DATAI_22_), .ZN(n14768) );
  NAND4_X1 U18118 ( .A1(n14771), .A2(n14770), .A3(n14769), .A4(n14768), .ZN(
        P1_U2882) );
  OAI22_X1 U18119 ( .A1(n14772), .A2(n14788), .B1(n14802), .B2(n21114), .ZN(
        n14773) );
  AOI21_X1 U18120 ( .B1(n16648), .B2(DATAI_21_), .A(n14773), .ZN(n14775) );
  NAND2_X1 U18121 ( .A1(n14791), .A2(BUF1_REG_21__SCAN_IN), .ZN(n14774) );
  OAI211_X1 U18122 ( .C1(n14776), .C2(n14805), .A(n14775), .B(n14774), .ZN(
        P1_U2883) );
  OAI22_X1 U18123 ( .A1(n14777), .A2(n14788), .B1(n14802), .B2(n13230), .ZN(
        n14778) );
  AOI21_X1 U18124 ( .B1(n16648), .B2(DATAI_19_), .A(n14778), .ZN(n14780) );
  NAND2_X1 U18125 ( .A1(n14791), .A2(BUF1_REG_19__SCAN_IN), .ZN(n14779) );
  OAI211_X1 U18126 ( .C1(n14781), .C2(n14805), .A(n14780), .B(n14779), .ZN(
        P1_U2885) );
  INV_X1 U18127 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14786) );
  NAND2_X1 U18128 ( .A1(n16579), .A2(n16649), .ZN(n14785) );
  OAI22_X1 U18129 ( .A1(n14782), .A2(n14788), .B1(n14802), .B2(n13239), .ZN(
        n14783) );
  AOI21_X1 U18130 ( .B1(n16648), .B2(DATAI_18_), .A(n14783), .ZN(n14784) );
  OAI211_X1 U18131 ( .C1(n16652), .C2(n14786), .A(n14785), .B(n14784), .ZN(
        P1_U2886) );
  OAI22_X1 U18132 ( .A1(n14789), .A2(n14788), .B1(n14802), .B2(n14787), .ZN(
        n14790) );
  AOI21_X1 U18133 ( .B1(n16648), .B2(DATAI_17_), .A(n14790), .ZN(n14793) );
  NAND2_X1 U18134 ( .A1(n14791), .A2(BUF1_REG_17__SCAN_IN), .ZN(n14792) );
  OAI211_X1 U18135 ( .C1(n14794), .C2(n14805), .A(n14793), .B(n14792), .ZN(
        P1_U2887) );
  OAI222_X1 U18136 ( .A1(n21064), .A2(n14805), .B1(n14802), .B2(n13226), .C1(
        n14795), .C2(n14804), .ZN(P1_U2889) );
  INV_X1 U18137 ( .A(n14796), .ZN(n14797) );
  AOI21_X1 U18138 ( .B1(n9722), .B2(n14718), .A(n14797), .ZN(n16665) );
  INV_X1 U18139 ( .A(n16665), .ZN(n14799) );
  INV_X1 U18140 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14798) );
  OAI222_X1 U18141 ( .A1(n14799), .A2(n14805), .B1(n20766), .B2(n14804), .C1(
        n14798), .C2(n14802), .ZN(P1_U2890) );
  INV_X1 U18142 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14800) );
  OAI222_X1 U18143 ( .A1(n14801), .A2(n14805), .B1(n20763), .B2(n14804), .C1(
        n14800), .C2(n14802), .ZN(P1_U2891) );
  INV_X1 U18144 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14803) );
  OAI222_X1 U18145 ( .A1(n16620), .A2(n14805), .B1(n20760), .B2(n14804), .C1(
        n14803), .C2(n14802), .ZN(P1_U2892) );
  INV_X1 U18146 ( .A(n14816), .ZN(n14806) );
  NAND3_X1 U18147 ( .A1(n14838), .A2(n15038), .A3(n14806), .ZN(n14807) );
  OAI21_X1 U18148 ( .B1(n14808), .B2(n14817), .A(n14807), .ZN(n14809) );
  XNOR2_X1 U18149 ( .A(n14809), .B(n15000), .ZN(n15018) );
  INV_X1 U18150 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14810) );
  NOR2_X1 U18151 ( .A1(n16817), .A2(n14810), .ZN(n15020) );
  AOI21_X1 U18152 ( .B1(n21061), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15020), .ZN(n14811) );
  OAI21_X1 U18153 ( .B1(n16695), .B2(n14812), .A(n14811), .ZN(n14813) );
  AOI21_X1 U18154 ( .B1(n15018), .B2(n20792), .A(n14813), .ZN(n14814) );
  OAI21_X1 U18155 ( .B1(n14815), .B2(n21063), .A(n14814), .ZN(P1_U2969) );
  NAND2_X1 U18156 ( .A1(n14817), .A2(n14816), .ZN(n14819) );
  XOR2_X1 U18157 ( .A(n14819), .B(n14818), .Z(n15035) );
  INV_X1 U18158 ( .A(n14820), .ZN(n14824) );
  NOR2_X1 U18159 ( .A1(n16817), .A2(n21026), .ZN(n15027) );
  AOI21_X1 U18160 ( .B1(n21061), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15027), .ZN(n14821) );
  OAI21_X1 U18161 ( .B1(n16695), .B2(n14822), .A(n14821), .ZN(n14823) );
  AOI21_X1 U18162 ( .B1(n14824), .B2(n20791), .A(n14823), .ZN(n14825) );
  OAI21_X1 U18163 ( .B1(n21068), .B2(n15035), .A(n14825), .ZN(P1_U2970) );
  INV_X1 U18164 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14830) );
  NOR2_X1 U18165 ( .A1(n16817), .A2(n14830), .ZN(n15041) );
  AOI21_X1 U18166 ( .B1(n21061), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15041), .ZN(n14831) );
  OAI21_X1 U18167 ( .B1(n16695), .B2(n14832), .A(n14831), .ZN(n14833) );
  AOI21_X1 U18168 ( .B1(n14834), .B2(n20791), .A(n14833), .ZN(n14835) );
  OAI21_X1 U18169 ( .B1(n21068), .B2(n15045), .A(n14835), .ZN(P1_U2971) );
  AND2_X1 U18170 ( .A1(n14849), .A2(n14836), .ZN(n14837) );
  MUX2_X1 U18171 ( .A(n14838), .B(n14837), .S(n15123), .Z(n14839) );
  XNOR2_X1 U18172 ( .A(n14839), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15055) );
  INV_X1 U18173 ( .A(n14840), .ZN(n14845) );
  INV_X1 U18174 ( .A(n14841), .ZN(n14843) );
  NOR2_X1 U18175 ( .A1(n16817), .A2(n21019), .ZN(n15047) );
  AOI21_X1 U18176 ( .B1(n21061), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15047), .ZN(n14842) );
  OAI21_X1 U18177 ( .B1(n16695), .B2(n14843), .A(n14842), .ZN(n14844) );
  AOI21_X1 U18178 ( .B1(n14845), .B2(n20791), .A(n14844), .ZN(n14846) );
  OAI21_X1 U18179 ( .B1(n21068), .B2(n15055), .A(n14846), .ZN(P1_U2972) );
  NOR2_X1 U18180 ( .A1(n15123), .A2(n15009), .ZN(n14848) );
  OAI21_X1 U18181 ( .B1(n14849), .B2(n14848), .A(n14847), .ZN(n14851) );
  XNOR2_X1 U18182 ( .A(n14851), .B(n14850), .ZN(n15065) );
  INV_X1 U18183 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21020) );
  NOR2_X1 U18184 ( .A1(n16817), .A2(n21020), .ZN(n15058) );
  AOI21_X1 U18185 ( .B1(n21061), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15058), .ZN(n14852) );
  OAI21_X1 U18186 ( .B1(n16695), .B2(n14853), .A(n14852), .ZN(n14854) );
  AOI21_X1 U18187 ( .B1(n14855), .B2(n20791), .A(n14854), .ZN(n14856) );
  OAI21_X1 U18188 ( .B1(n21068), .B2(n15065), .A(n14856), .ZN(P1_U2973) );
  XNOR2_X1 U18189 ( .A(n16656), .B(n15089), .ZN(n14874) );
  AOI21_X1 U18190 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15123), .A(
        n14874), .ZN(n14857) );
  OAI211_X1 U18191 ( .C1(n14875), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14857), .B(n14847), .ZN(n14858) );
  XNOR2_X1 U18192 ( .A(n14858), .B(n15067), .ZN(n15074) );
  NOR2_X1 U18193 ( .A1(n16817), .A2(n14859), .ZN(n15069) );
  AOI21_X1 U18194 ( .B1(n21061), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15069), .ZN(n14860) );
  OAI21_X1 U18195 ( .B1(n16695), .B2(n14861), .A(n14860), .ZN(n14862) );
  AOI21_X1 U18196 ( .B1(n14863), .B2(n20791), .A(n14862), .ZN(n14864) );
  OAI21_X1 U18197 ( .B1(n21068), .B2(n15074), .A(n14864), .ZN(P1_U2974) );
  AOI21_X1 U18198 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15123), .A(
        n14865), .ZN(n14866) );
  AOI21_X1 U18199 ( .B1(n15089), .B2(n16656), .A(n14866), .ZN(n14868) );
  XNOR2_X1 U18200 ( .A(n16656), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14867) );
  XNOR2_X1 U18201 ( .A(n14868), .B(n14867), .ZN(n15085) );
  INV_X1 U18202 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21017) );
  NOR2_X1 U18203 ( .A1(n16817), .A2(n21017), .ZN(n15082) );
  AOI21_X1 U18204 ( .B1(n21061), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15082), .ZN(n14869) );
  OAI21_X1 U18205 ( .B1(n16695), .B2(n14870), .A(n14869), .ZN(n14871) );
  AOI21_X1 U18206 ( .B1(n14872), .B2(n20791), .A(n14871), .ZN(n14873) );
  OAI21_X1 U18207 ( .B1(n21068), .B2(n15085), .A(n14873), .ZN(P1_U2975) );
  XNOR2_X1 U18208 ( .A(n14875), .B(n14874), .ZN(n15094) );
  INV_X1 U18209 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14876) );
  NOR2_X1 U18210 ( .A1(n16817), .A2(n14876), .ZN(n15086) );
  AOI21_X1 U18211 ( .B1(n21061), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15086), .ZN(n14877) );
  OAI21_X1 U18212 ( .B1(n16695), .B2(n14878), .A(n14877), .ZN(n14879) );
  AOI21_X1 U18213 ( .B1(n14880), .B2(n20791), .A(n14879), .ZN(n14881) );
  OAI21_X1 U18214 ( .B1(n15094), .B2(n21068), .A(n14881), .ZN(P1_U2976) );
  NAND2_X1 U18215 ( .A1(n14883), .A2(n14882), .ZN(n14884) );
  XOR2_X1 U18216 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14884), .Z(
        n16702) );
  AOI22_X1 U18217 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14885) );
  OAI21_X1 U18218 ( .B1(n16695), .B2(n14886), .A(n14885), .ZN(n14887) );
  AOI21_X1 U18219 ( .B1(n14888), .B2(n20791), .A(n14887), .ZN(n14889) );
  OAI21_X1 U18220 ( .B1(n21068), .B2(n16702), .A(n14889), .ZN(P1_U2977) );
  NOR2_X1 U18221 ( .A1(n14890), .A2(n16656), .ZN(n14898) );
  NOR2_X1 U18222 ( .A1(n14891), .A2(n15123), .ZN(n14899) );
  MUX2_X1 U18223 ( .A(n14898), .B(n14899), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n14892) );
  XNOR2_X1 U18224 ( .A(n14892), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15107) );
  INV_X1 U18225 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21011) );
  NOR2_X1 U18226 ( .A1(n16817), .A2(n21011), .ZN(n15101) );
  AOI21_X1 U18227 ( .B1(n21061), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15101), .ZN(n14893) );
  OAI21_X1 U18228 ( .B1(n16695), .B2(n14894), .A(n14893), .ZN(n14895) );
  AOI21_X1 U18229 ( .B1(n14896), .B2(n20791), .A(n14895), .ZN(n14897) );
  OAI21_X1 U18230 ( .B1(n15107), .B2(n21068), .A(n14897), .ZN(P1_U2978) );
  NOR2_X1 U18231 ( .A1(n14899), .A2(n14898), .ZN(n14900) );
  XOR2_X1 U18232 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n14900), .Z(
        n15119) );
  INV_X1 U18233 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14901) );
  NOR2_X1 U18234 ( .A1(n16817), .A2(n14901), .ZN(n15115) );
  AOI21_X1 U18235 ( .B1(n21061), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15115), .ZN(n14902) );
  OAI21_X1 U18236 ( .B1(n16695), .B2(n16573), .A(n14902), .ZN(n14903) );
  AOI21_X1 U18237 ( .B1(n16642), .B2(n20791), .A(n14903), .ZN(n14904) );
  OAI21_X1 U18238 ( .B1(n15119), .B2(n21068), .A(n14904), .ZN(P1_U2979) );
  OAI21_X1 U18239 ( .B1(n16656), .B2(n16729), .A(n14913), .ZN(n14906) );
  XNOR2_X1 U18240 ( .A(n16656), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14905) );
  XNOR2_X1 U18241 ( .A(n14906), .B(n14905), .ZN(n16712) );
  INV_X1 U18242 ( .A(n14907), .ZN(n14909) );
  AOI22_X1 U18243 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14908) );
  OAI21_X1 U18244 ( .B1(n16695), .B2(n14909), .A(n14908), .ZN(n14910) );
  AOI21_X1 U18245 ( .B1(n14911), .B2(n20791), .A(n14910), .ZN(n14912) );
  OAI21_X1 U18246 ( .B1(n16712), .B2(n21068), .A(n14912), .ZN(P1_U2980) );
  OAI21_X1 U18247 ( .B1(n14915), .B2(n14914), .A(n14913), .ZN(n16725) );
  INV_X1 U18248 ( .A(n16725), .ZN(n14918) );
  AOI22_X1 U18249 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14916) );
  OAI21_X1 U18250 ( .B1(n16695), .B2(n16574), .A(n14916), .ZN(n14917) );
  AOI21_X1 U18251 ( .B1(n14918), .B2(n20792), .A(n14917), .ZN(n14919) );
  OAI21_X1 U18252 ( .B1(n14920), .B2(n21063), .A(n14919), .ZN(P1_U2981) );
  NAND2_X1 U18253 ( .A1(n14922), .A2(n15121), .ZN(n14924) );
  OAI21_X1 U18254 ( .B1(n14921), .B2(n14924), .A(n14923), .ZN(n14926) );
  NAND2_X1 U18255 ( .A1(n14926), .A2(n16742), .ZN(n14925) );
  MUX2_X1 U18256 ( .A(n14926), .B(n14925), .S(n15123), .Z(n14928) );
  XNOR2_X1 U18257 ( .A(n14928), .B(n14927), .ZN(n16731) );
  AOI22_X1 U18258 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n14929) );
  OAI21_X1 U18259 ( .B1(n16695), .B2(n14930), .A(n14929), .ZN(n14931) );
  AOI21_X1 U18260 ( .B1(n14932), .B2(n20791), .A(n14931), .ZN(n14933) );
  OAI21_X1 U18261 ( .B1(n21068), .B2(n16731), .A(n14933), .ZN(P1_U2982) );
  INV_X1 U18262 ( .A(n14934), .ZN(n14936) );
  NOR2_X1 U18263 ( .A1(n14921), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16676) );
  AOI21_X1 U18264 ( .B1(n16676), .B2(n16776), .A(n16656), .ZN(n14935) );
  AOI21_X1 U18265 ( .B1(n14936), .B2(n14921), .A(n14935), .ZN(n15145) );
  INV_X1 U18266 ( .A(n14938), .ZN(n14937) );
  AOI21_X1 U18267 ( .B1(n15123), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14937), .ZN(n15144) );
  NAND2_X1 U18268 ( .A1(n15145), .A2(n15144), .ZN(n15143) );
  NAND2_X1 U18269 ( .A1(n15143), .A2(n14938), .ZN(n14940) );
  XNOR2_X1 U18270 ( .A(n14940), .B(n14939), .ZN(n16765) );
  INV_X1 U18271 ( .A(n16765), .ZN(n14944) );
  AOI22_X1 U18272 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14941) );
  OAI21_X1 U18273 ( .B1(n16695), .B2(n16613), .A(n14941), .ZN(n14942) );
  AOI21_X1 U18274 ( .B1(n16617), .B2(n20791), .A(n14942), .ZN(n14943) );
  OAI21_X1 U18275 ( .B1(n14944), .B2(n21068), .A(n14943), .ZN(P1_U2986) );
  MUX2_X1 U18276 ( .A(n16675), .B(n14921), .S(n15123), .Z(n14945) );
  XOR2_X1 U18277 ( .A(n12132), .B(n14945), .Z(n16787) );
  NAND2_X1 U18278 ( .A1(n16787), .A2(n20792), .ZN(n14951) );
  OAI22_X1 U18279 ( .A1(n14947), .A2(n14946), .B1(n16817), .B2(n20996), .ZN(
        n14948) );
  AOI21_X1 U18280 ( .B1(n16669), .B2(n14949), .A(n14948), .ZN(n14950) );
  OAI211_X1 U18281 ( .C1(n21063), .C2(n14952), .A(n14951), .B(n14950), .ZN(
        P1_U2989) );
  OR2_X1 U18282 ( .A1(n14955), .A2(n14954), .ZN(n14962) );
  NAND2_X1 U18283 ( .A1(n14956), .A2(n21051), .ZN(n14958) );
  OAI211_X1 U18284 ( .C1(n13135), .C2(n14958), .A(n14957), .B(n11204), .ZN(
        n14960) );
  NAND2_X1 U18285 ( .A1(n14960), .A2(n14959), .ZN(n14961) );
  MUX2_X1 U18286 ( .A(n14962), .B(n14961), .S(n11128), .Z(n14966) );
  NAND3_X1 U18287 ( .A1(n14963), .A2(n11532), .A3(n14978), .ZN(n14964) );
  NAND3_X1 U18288 ( .A1(n14966), .A2(n14965), .A3(n14964), .ZN(n14968) );
  OAI211_X1 U18289 ( .C1(n14970), .C2(n14976), .A(n16520), .B(n14969), .ZN(
        n14971) );
  INV_X1 U18290 ( .A(n14971), .ZN(n14972) );
  NAND2_X1 U18291 ( .A1(n14973), .A2(n14972), .ZN(n14974) );
  INV_X1 U18292 ( .A(n14975), .ZN(n15016) );
  OAI22_X1 U18293 ( .A1(n12908), .A2(n14978), .B1(n14977), .B2(n14976), .ZN(
        n14979) );
  NOR2_X1 U18294 ( .A1(n12128), .A2(n16742), .ZN(n16738) );
  NAND3_X1 U18295 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n16738), .ZN(n16723) );
  NOR2_X1 U18296 ( .A1(n16729), .A2(n16723), .ZN(n15007) );
  NAND2_X1 U18297 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20796) );
  NOR2_X1 U18298 ( .A1(n14980), .A2(n20796), .ZN(n16798) );
  OAI21_X1 U18299 ( .B1(n20828), .B2(n20852), .A(n20822), .ZN(n20812) );
  NAND2_X1 U18300 ( .A1(n16798), .A2(n20812), .ZN(n16781) );
  NOR3_X1 U18301 ( .A1(n16815), .A2(n16821), .A3(n16808), .ZN(n16785) );
  NAND3_X1 U18302 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16785), .ZN(n14988) );
  NOR2_X1 U18303 ( .A1(n16781), .A2(n14988), .ZN(n16771) );
  NAND2_X1 U18304 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16771), .ZN(
        n15150) );
  NOR2_X1 U18305 ( .A1(n15154), .A2(n15150), .ZN(n15131) );
  AND2_X1 U18306 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15131), .ZN(
        n16722) );
  AND2_X1 U18307 ( .A1(n15007), .A2(n16722), .ZN(n14991) );
  NAND2_X1 U18308 ( .A1(n14983), .A2(n14982), .ZN(n14984) );
  NAND2_X1 U18309 ( .A1(n14985), .A2(n14984), .ZN(n14986) );
  NAND2_X1 U18310 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20813) );
  INV_X1 U18311 ( .A(n20813), .ZN(n14987) );
  NAND2_X1 U18312 ( .A1(n16798), .A2(n14987), .ZN(n16782) );
  NOR2_X1 U18313 ( .A1(n14988), .A2(n16782), .ZN(n15147) );
  NAND3_X1 U18314 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n15147), .ZN(n16762) );
  INV_X1 U18315 ( .A(n16762), .ZN(n15133) );
  INV_X1 U18316 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16768) );
  INV_X1 U18317 ( .A(n15007), .ZN(n14989) );
  NOR2_X1 U18318 ( .A1(n16768), .A2(n14989), .ZN(n15098) );
  NAND2_X1 U18319 ( .A1(n15133), .A2(n15098), .ZN(n15099) );
  NAND2_X1 U18320 ( .A1(n16801), .A2(n15099), .ZN(n14990) );
  OAI21_X1 U18321 ( .B1(n14991), .B2(n16799), .A(n14990), .ZN(n14993) );
  NOR2_X1 U18322 ( .A1(n21060), .A2(n14992), .ZN(n20839) );
  OR2_X1 U18323 ( .A1(n14993), .A2(n16800), .ZN(n16718) );
  NOR2_X1 U18324 ( .A1(n16717), .A2(n15110), .ZN(n15100) );
  INV_X1 U18325 ( .A(n15100), .ZN(n14994) );
  INV_X1 U18326 ( .A(n16800), .ZN(n20829) );
  INV_X1 U18327 ( .A(n16807), .ZN(n20826) );
  NAND2_X1 U18328 ( .A1(n20829), .A2(n20826), .ZN(n16783) );
  OAI21_X1 U18329 ( .B1(n16718), .B2(n14994), .A(n16783), .ZN(n16703) );
  NAND2_X1 U18330 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16708) );
  NAND2_X1 U18331 ( .A1(n16807), .A2(n16708), .ZN(n14995) );
  AND2_X1 U18332 ( .A1(n16703), .A2(n14995), .ZN(n15090) );
  INV_X1 U18333 ( .A(n14996), .ZN(n15077) );
  NAND2_X1 U18334 ( .A1(n16807), .A2(n15077), .ZN(n15068) );
  AND2_X1 U18335 ( .A1(n15068), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14997) );
  AND2_X1 U18336 ( .A1(n15090), .A2(n14997), .ZN(n15061) );
  NAND2_X1 U18337 ( .A1(n15061), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15046) );
  INV_X1 U18338 ( .A(n15038), .ZN(n14998) );
  OR2_X1 U18339 ( .A1(n15046), .A2(n14998), .ZN(n14999) );
  NAND2_X1 U18340 ( .A1(n14999), .A2(n16783), .ZN(n15031) );
  INV_X1 U18341 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15030) );
  AOI21_X1 U18342 ( .B1(n16807), .B2(n15030), .A(n15000), .ZN(n15001) );
  NAND2_X1 U18343 ( .A1(n15031), .A2(n15001), .ZN(n15022) );
  NAND3_X1 U18344 ( .A1(n15022), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16783), .ZN(n15014) );
  INV_X1 U18345 ( .A(n15002), .ZN(n15013) );
  NOR2_X1 U18346 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20838), .ZN(
        n20825) );
  INV_X1 U18347 ( .A(n20825), .ZN(n15003) );
  NAND2_X1 U18348 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15133), .ZN(
        n16759) );
  INV_X1 U18349 ( .A(n16759), .ZN(n15135) );
  NAND2_X1 U18350 ( .A1(n20811), .A2(n15135), .ZN(n15076) );
  NAND2_X1 U18351 ( .A1(n20827), .A2(n15131), .ZN(n15096) );
  INV_X1 U18352 ( .A(n15096), .ZN(n15004) );
  NAND2_X1 U18353 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15004), .ZN(
        n15005) );
  INV_X1 U18354 ( .A(n16708), .ZN(n15006) );
  NAND4_X1 U18355 ( .A1(n15007), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(n15006), .ZN(n15008) );
  INV_X1 U18356 ( .A(n15009), .ZN(n15056) );
  NAND2_X1 U18357 ( .A1(n15056), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15010) );
  NOR2_X1 U18358 ( .A1(n15057), .A2(n15010), .ZN(n15049) );
  AND2_X1 U18359 ( .A1(n15038), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15011) );
  AND2_X1 U18360 ( .A1(n15049), .A2(n15011), .ZN(n15019) );
  INV_X1 U18361 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21093) );
  NAND3_X1 U18362 ( .A1(n15019), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n21093), .ZN(n15012) );
  NAND3_X1 U18363 ( .A1(n15014), .A2(n15013), .A3(n15012), .ZN(n15015) );
  AOI21_X1 U18364 ( .B1(n15016), .B2(n20849), .A(n15015), .ZN(n15017) );
  OAI21_X1 U18365 ( .B1(n9682), .B2(n20844), .A(n15017), .ZN(P1_U3000) );
  NAND2_X1 U18366 ( .A1(n15018), .A2(n20806), .ZN(n15024) );
  OR2_X1 U18367 ( .A1(n15019), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15021) );
  AOI21_X1 U18368 ( .B1(n15022), .B2(n15021), .A(n15020), .ZN(n15023) );
  OAI211_X1 U18369 ( .C1(n20836), .C2(n15025), .A(n15024), .B(n15023), .ZN(
        P1_U3001) );
  INV_X1 U18370 ( .A(n15026), .ZN(n15033) );
  INV_X1 U18371 ( .A(n15027), .ZN(n15029) );
  NAND3_X1 U18372 ( .A1(n15049), .A2(n15038), .A3(n15030), .ZN(n15028) );
  OAI211_X1 U18373 ( .C1(n15031), .C2(n15030), .A(n15029), .B(n15028), .ZN(
        n15032) );
  AOI21_X1 U18374 ( .B1(n15033), .B2(n20849), .A(n15032), .ZN(n15034) );
  OAI21_X1 U18375 ( .B1(n15035), .B2(n20844), .A(n15034), .ZN(P1_U3002) );
  NOR2_X1 U18376 ( .A1(n15036), .A2(n20836), .ZN(n15043) );
  AND3_X1 U18377 ( .A1(n15046), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16783), .ZN(n15042) );
  INV_X1 U18378 ( .A(n15049), .ZN(n15039) );
  NOR3_X1 U18379 ( .A1(n15039), .A2(n15038), .A3(n15037), .ZN(n15040) );
  NOR4_X1 U18380 ( .A1(n15043), .A2(n15042), .A3(n15041), .A4(n15040), .ZN(
        n15044) );
  OAI21_X1 U18381 ( .B1(n15045), .B2(n20844), .A(n15044), .ZN(P1_U3003) );
  NAND3_X1 U18382 ( .A1(n15046), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16783), .ZN(n15051) );
  AOI21_X1 U18383 ( .B1(n15049), .B2(n15048), .A(n15047), .ZN(n15050) );
  NAND2_X1 U18384 ( .A1(n15051), .A2(n15050), .ZN(n15052) );
  AOI21_X1 U18385 ( .B1(n15053), .B2(n20849), .A(n15052), .ZN(n15054) );
  OAI21_X1 U18386 ( .B1(n15055), .B2(n20844), .A(n15054), .ZN(P1_U3004) );
  INV_X1 U18387 ( .A(n15057), .ZN(n15087) );
  AOI21_X1 U18388 ( .B1(n15087), .B2(n15056), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15060) );
  NOR3_X1 U18389 ( .A1(n15057), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15077), .ZN(n15071) );
  AOI21_X1 U18390 ( .B1(n15071), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15058), .ZN(n15059) );
  OAI21_X1 U18391 ( .B1(n15061), .B2(n15060), .A(n15059), .ZN(n15062) );
  AOI21_X1 U18392 ( .B1(n15063), .B2(n20849), .A(n15062), .ZN(n15064) );
  OAI21_X1 U18393 ( .B1(n15065), .B2(n20844), .A(n15064), .ZN(P1_U3005) );
  NOR2_X1 U18394 ( .A1(n15066), .A2(n20836), .ZN(n15072) );
  AOI21_X1 U18395 ( .B1(n15090), .B2(n15068), .A(n15067), .ZN(n15070) );
  NOR4_X1 U18396 ( .A1(n15072), .A2(n15071), .A3(n15070), .A4(n15069), .ZN(
        n15073) );
  OAI21_X1 U18397 ( .B1(n15074), .B2(n20844), .A(n15073), .ZN(P1_U3006) );
  INV_X1 U18398 ( .A(n15075), .ZN(n15083) );
  INV_X1 U18399 ( .A(n15076), .ZN(n15078) );
  OAI21_X1 U18400 ( .B1(n15078), .B2(n20827), .A(n15077), .ZN(n15080) );
  AOI21_X1 U18401 ( .B1(n15087), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15079) );
  AOI21_X1 U18402 ( .B1(n15090), .B2(n15080), .A(n15079), .ZN(n15081) );
  AOI211_X1 U18403 ( .C1(n15083), .C2(n20849), .A(n15082), .B(n15081), .ZN(
        n15084) );
  OAI21_X1 U18404 ( .B1(n15085), .B2(n20844), .A(n15084), .ZN(P1_U3007) );
  AOI21_X1 U18405 ( .B1(n15087), .B2(n15089), .A(n15086), .ZN(n15088) );
  OAI21_X1 U18406 ( .B1(n15090), .B2(n15089), .A(n15088), .ZN(n15091) );
  AOI21_X1 U18407 ( .B1(n15092), .B2(n20849), .A(n15091), .ZN(n15093) );
  OAI21_X1 U18408 ( .B1(n15094), .B2(n20844), .A(n15093), .ZN(P1_U3008) );
  INV_X1 U18409 ( .A(n15095), .ZN(n15105) );
  INV_X1 U18410 ( .A(n20838), .ZN(n15136) );
  NAND3_X1 U18411 ( .A1(n15132), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n15133), .ZN(n15097) );
  NAND2_X1 U18412 ( .A1(n15097), .A2(n15096), .ZN(n15139) );
  NAND2_X1 U18413 ( .A1(n15139), .A2(n15098), .ZN(n15108) );
  OAI21_X1 U18414 ( .B1(n15099), .B2(n15136), .A(n15108), .ZN(n16716) );
  AND2_X1 U18415 ( .A1(n15100), .A2(n16716), .ZN(n16709) );
  AOI21_X1 U18416 ( .B1(n16709), .B2(n15103), .A(n15101), .ZN(n15102) );
  OAI21_X1 U18417 ( .B1(n16703), .B2(n15103), .A(n15102), .ZN(n15104) );
  AOI21_X1 U18418 ( .B1(n15105), .B2(n20849), .A(n15104), .ZN(n15106) );
  OAI21_X1 U18419 ( .B1(n15107), .B2(n20844), .A(n15106), .ZN(P1_U3010) );
  NOR2_X1 U18420 ( .A1(n16567), .A2(n20836), .ZN(n15117) );
  INV_X1 U18421 ( .A(n16718), .ZN(n15112) );
  INV_X1 U18422 ( .A(n15108), .ZN(n15109) );
  OAI21_X1 U18423 ( .B1(n15109), .B2(n20838), .A(n16717), .ZN(n15111) );
  AOI21_X1 U18424 ( .B1(n15112), .B2(n15111), .A(n15110), .ZN(n15116) );
  INV_X1 U18425 ( .A(n16716), .ZN(n15113) );
  NOR3_X1 U18426 ( .A1(n15113), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n16717), .ZN(n15114) );
  NOR4_X1 U18427 ( .A1(n15117), .A2(n15116), .A3(n15115), .A4(n15114), .ZN(
        n15118) );
  OAI21_X1 U18428 ( .B1(n15119), .B2(n20844), .A(n15118), .ZN(P1_U3011) );
  INV_X1 U18429 ( .A(n14921), .ZN(n15122) );
  AOI21_X1 U18430 ( .B1(n15122), .B2(n15121), .A(n15120), .ZN(n15125) );
  NOR2_X1 U18431 ( .A1(n15125), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15124) );
  MUX2_X1 U18432 ( .A(n15125), .B(n15124), .S(n15123), .Z(n15126) );
  XNOR2_X1 U18433 ( .A(n15126), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16668) );
  XNOR2_X1 U18434 ( .A(n15128), .B(n15127), .ZN(n16638) );
  INV_X1 U18435 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21002) );
  OR2_X1 U18436 ( .A1(n16817), .A2(n21002), .ZN(n15130) );
  NAND3_X1 U18437 ( .A1(n16722), .A2(n16741), .A3(n16829), .ZN(n15129) );
  NAND2_X1 U18438 ( .A1(n15130), .A2(n15129), .ZN(n15141) );
  INV_X1 U18439 ( .A(n15131), .ZN(n15138) );
  INV_X1 U18440 ( .A(n15132), .ZN(n15134) );
  OAI22_X1 U18441 ( .A1(n15136), .A2(n15135), .B1(n15134), .B2(n15133), .ZN(
        n15137) );
  AOI211_X1 U18442 ( .C1(n20827), .C2(n15138), .A(n16800), .B(n15137), .ZN(
        n16769) );
  NAND2_X1 U18443 ( .A1(n16768), .A2(n15139), .ZN(n16766) );
  AOI21_X1 U18444 ( .B1(n16769), .B2(n16766), .A(n16741), .ZN(n15140) );
  AOI211_X1 U18445 ( .C1(n20849), .C2(n16638), .A(n15141), .B(n15140), .ZN(
        n15142) );
  OAI21_X1 U18446 ( .B1(n16668), .B2(n20844), .A(n15142), .ZN(P1_U3017) );
  OAI21_X1 U18447 ( .B1(n15145), .B2(n15144), .A(n15143), .ZN(n15146) );
  INV_X1 U18448 ( .A(n15146), .ZN(n16674) );
  NOR2_X1 U18449 ( .A1(n16778), .A2(n15150), .ZN(n15155) );
  INV_X1 U18450 ( .A(n16801), .ZN(n15148) );
  OAI21_X1 U18451 ( .B1(n15148), .B2(n15147), .A(n20829), .ZN(n15149) );
  AOI21_X1 U18452 ( .B1(n20827), .B2(n15150), .A(n15149), .ZN(n16777) );
  OAI21_X1 U18453 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15151), .A(
        n16777), .ZN(n15153) );
  OAI22_X1 U18454 ( .A1(n16817), .A2(n20998), .B1(n20836), .B2(n16625), .ZN(
        n15152) );
  AOI221_X1 U18455 ( .B1(n15155), .B2(n15154), .C1(n15153), .C2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n15152), .ZN(n15156) );
  OAI21_X1 U18456 ( .B1(n16674), .B2(n20844), .A(n15156), .ZN(P1_U3019) );
  OAI211_X1 U18457 ( .C1(n15158), .C2(P1_STATEBS16_REG_SCAN_IN), .A(n15157), 
        .B(n15161), .ZN(n15159) );
  OAI21_X1 U18458 ( .B1(n15166), .B2(n20896), .A(n15159), .ZN(n15160) );
  MUX2_X1 U18459 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15160), .S(
        n20853), .Z(P1_U3477) );
  XNOR2_X1 U18460 ( .A(n12060), .B(n15161), .ZN(n15163) );
  OAI22_X1 U18461 ( .A1(n15163), .A2(n20893), .B1(n15162), .B2(n15166), .ZN(
        n15164) );
  MUX2_X1 U18462 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15164), .S(
        n20853), .Z(P1_U3476) );
  INV_X1 U18463 ( .A(n13150), .ZN(n15167) );
  OAI21_X1 U18464 ( .B1(n15167), .B2(n15166), .A(n15165), .ZN(n15168) );
  MUX2_X1 U18465 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15168), .S(
        n20853), .Z(P1_U3475) );
  NAND2_X1 U18466 ( .A1(n20858), .A2(n15169), .ZN(n15172) );
  NAND3_X1 U18467 ( .A1(n11532), .A2(n15174), .A3(n15170), .ZN(n15171) );
  OAI211_X1 U18468 ( .C1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n15173), .A(
        n15172), .B(n15171), .ZN(n16504) );
  INV_X1 U18469 ( .A(n16504), .ZN(n15177) );
  INV_X1 U18470 ( .A(n20632), .ZN(n16838) );
  OAI22_X1 U18471 ( .A1(n21093), .A2(n20828), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15179) );
  NOR2_X1 U18472 ( .A1(n20962), .A2(n20852), .ZN(n15181) );
  NOR3_X1 U18473 ( .A1(n13170), .A2(n13140), .A3(n15186), .ZN(n15175) );
  AOI21_X1 U18474 ( .B1(n15179), .B2(n15181), .A(n15175), .ZN(n15176) );
  OAI21_X1 U18475 ( .B1(n15177), .B2(n16838), .A(n15176), .ZN(n15178) );
  MUX2_X1 U18476 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15178), .S(
        n16842), .Z(P1_U3473) );
  INV_X1 U18477 ( .A(n15179), .ZN(n15180) );
  AOI22_X1 U18478 ( .A1(n15182), .A2(n16539), .B1(n15181), .B2(n15180), .ZN(
        n15183) );
  OAI21_X1 U18479 ( .B1(n15184), .B2(n16838), .A(n15183), .ZN(n15185) );
  MUX2_X1 U18480 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15185), .S(
        n16842), .Z(P1_U3472) );
  OAI22_X1 U18481 ( .A1(n15188), .A2(n16838), .B1(n15187), .B2(n15186), .ZN(
        n15189) );
  MUX2_X1 U18482 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15189), .S(
        n16842), .Z(P1_U3469) );
  NAND3_X1 U18483 ( .A1(n15238), .A2(n15157), .A3(n15237), .ZN(n15190) );
  NAND2_X1 U18484 ( .A1(n15190), .A2(n20855), .ZN(n15195) );
  NOR2_X1 U18485 ( .A1(n15191), .A2(n20858), .ZN(n15193) );
  NAND2_X1 U18486 ( .A1(n20864), .A2(n15192), .ZN(n15196) );
  INV_X1 U18487 ( .A(n15196), .ZN(n15241) );
  INV_X1 U18488 ( .A(n15193), .ZN(n15194) );
  AOI22_X1 U18489 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15196), .B1(n15195), 
        .B2(n15194), .ZN(n15197) );
  OAI211_X1 U18490 ( .C1(n15198), .C2(n13658), .A(n20869), .B(n15197), .ZN(
        n15199) );
  OAI22_X1 U18491 ( .A1(n15237), .A2(n15201), .B1(n15200), .B2(n15234), .ZN(
        n15203) );
  NOR2_X1 U18492 ( .A1(n15238), .A2(n15253), .ZN(n15202) );
  AOI211_X1 U18493 ( .C1(n20902), .C2(n15241), .A(n15203), .B(n15202), .ZN(
        n15204) );
  OAI21_X1 U18494 ( .B1(n15243), .B2(n20915), .A(n15204), .ZN(P1_U3033) );
  OAI22_X1 U18495 ( .A1(n15237), .A2(n15206), .B1(n15205), .B2(n15234), .ZN(
        n15208) );
  NOR2_X1 U18496 ( .A1(n15238), .A2(n15258), .ZN(n15207) );
  AOI211_X1 U18497 ( .C1(n15241), .C2(n20916), .A(n15208), .B(n15207), .ZN(
        n15209) );
  OAI21_X1 U18498 ( .B1(n15243), .B2(n20921), .A(n15209), .ZN(P1_U3034) );
  OAI22_X1 U18499 ( .A1(n15237), .A2(n15211), .B1(n15210), .B2(n15234), .ZN(
        n15213) );
  NOR2_X1 U18500 ( .A1(n15238), .A2(n15263), .ZN(n15212) );
  AOI211_X1 U18501 ( .C1(n15241), .C2(n20922), .A(n15213), .B(n15212), .ZN(
        n15214) );
  OAI21_X1 U18502 ( .B1(n15243), .B2(n20927), .A(n15214), .ZN(P1_U3035) );
  OAI22_X1 U18503 ( .A1(n15237), .A2(n15215), .B1(n9837), .B2(n15234), .ZN(
        n15217) );
  NOR2_X1 U18504 ( .A1(n15238), .A2(n15268), .ZN(n15216) );
  AOI211_X1 U18505 ( .C1(n15241), .C2(n20928), .A(n15217), .B(n15216), .ZN(
        n15218) );
  OAI21_X1 U18506 ( .B1(n15243), .B2(n20933), .A(n15218), .ZN(P1_U3036) );
  OAI22_X1 U18507 ( .A1(n15237), .A2(n15220), .B1(n15219), .B2(n15234), .ZN(
        n15222) );
  NOR2_X1 U18508 ( .A1(n15238), .A2(n15273), .ZN(n15221) );
  AOI211_X1 U18509 ( .C1(n15241), .C2(n20934), .A(n15222), .B(n15221), .ZN(
        n15223) );
  OAI21_X1 U18510 ( .B1(n15243), .B2(n20939), .A(n15223), .ZN(P1_U3037) );
  INV_X1 U18511 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15224) );
  OAI22_X1 U18512 ( .A1(n15237), .A2(n15225), .B1(n15224), .B2(n15234), .ZN(
        n15227) );
  NOR2_X1 U18513 ( .A1(n15238), .A2(n15278), .ZN(n15226) );
  AOI211_X1 U18514 ( .C1(n15241), .C2(n20940), .A(n15227), .B(n15226), .ZN(
        n15228) );
  OAI21_X1 U18515 ( .B1(n15243), .B2(n20945), .A(n15228), .ZN(P1_U3038) );
  INV_X1 U18516 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15229) );
  OAI22_X1 U18517 ( .A1(n15237), .A2(n15230), .B1(n15229), .B2(n15234), .ZN(
        n15232) );
  NOR2_X1 U18518 ( .A1(n15238), .A2(n15283), .ZN(n15231) );
  AOI211_X1 U18519 ( .C1(n15241), .C2(n20946), .A(n15232), .B(n15231), .ZN(
        n15233) );
  OAI21_X1 U18520 ( .B1(n15243), .B2(n20951), .A(n15233), .ZN(P1_U3039) );
  OAI22_X1 U18521 ( .A1(n15237), .A2(n15236), .B1(n15235), .B2(n15234), .ZN(
        n15240) );
  NOR2_X1 U18522 ( .A1(n15238), .A2(n15289), .ZN(n15239) );
  AOI211_X1 U18523 ( .C1(n15241), .C2(n20952), .A(n15240), .B(n15239), .ZN(
        n15242) );
  OAI21_X1 U18524 ( .B1(n15243), .B2(n20960), .A(n15242), .ZN(P1_U3040) );
  NAND2_X1 U18525 ( .A1(n15290), .A2(n15157), .ZN(n15244) );
  OAI21_X1 U18526 ( .B1(n15294), .B2(n15244), .A(n20855), .ZN(n15250) );
  NOR2_X1 U18527 ( .A1(n15245), .A2(n20896), .ZN(n15247) );
  INV_X1 U18528 ( .A(n15247), .ZN(n15249) );
  NAND2_X1 U18529 ( .A1(n20864), .A2(n15248), .ZN(n15291) );
  AOI22_X1 U18530 ( .A1(n15250), .A2(n15249), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n15291), .ZN(n15252) );
  NAND3_X1 U18531 ( .A1(n20904), .A2(n15252), .A3(n15251), .ZN(n15288) );
  NAND2_X1 U18532 ( .A1(n15288), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n15257) );
  OAI22_X1 U18533 ( .A1(n15254), .A2(n15291), .B1(n15290), .B2(n15253), .ZN(
        n15255) );
  AOI21_X1 U18534 ( .B1(n15294), .B2(n20912), .A(n15255), .ZN(n15256) );
  OAI211_X1 U18535 ( .C1(n15297), .C2(n20915), .A(n15257), .B(n15256), .ZN(
        P1_U3081) );
  NAND2_X1 U18536 ( .A1(n15288), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n15262) );
  OAI22_X1 U18537 ( .A1(n15259), .A2(n15291), .B1(n15290), .B2(n15258), .ZN(
        n15260) );
  AOI21_X1 U18538 ( .B1(n15294), .B2(n20918), .A(n15260), .ZN(n15261) );
  OAI211_X1 U18539 ( .C1(n15297), .C2(n20921), .A(n15262), .B(n15261), .ZN(
        P1_U3082) );
  NAND2_X1 U18540 ( .A1(n15288), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n15267) );
  OAI22_X1 U18541 ( .A1(n15264), .A2(n15291), .B1(n15290), .B2(n15263), .ZN(
        n15265) );
  AOI21_X1 U18542 ( .B1(n15294), .B2(n20924), .A(n15265), .ZN(n15266) );
  OAI211_X1 U18543 ( .C1(n15297), .C2(n20927), .A(n15267), .B(n15266), .ZN(
        P1_U3083) );
  NAND2_X1 U18544 ( .A1(n15288), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n15272) );
  OAI22_X1 U18545 ( .A1(n15269), .A2(n15291), .B1(n15290), .B2(n15268), .ZN(
        n15270) );
  AOI21_X1 U18546 ( .B1(n15294), .B2(n20930), .A(n15270), .ZN(n15271) );
  OAI211_X1 U18547 ( .C1(n15297), .C2(n20933), .A(n15272), .B(n15271), .ZN(
        P1_U3084) );
  NAND2_X1 U18548 ( .A1(n15288), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n15277) );
  OAI22_X1 U18549 ( .A1(n15274), .A2(n15291), .B1(n15290), .B2(n15273), .ZN(
        n15275) );
  AOI21_X1 U18550 ( .B1(n15294), .B2(n20936), .A(n15275), .ZN(n15276) );
  OAI211_X1 U18551 ( .C1(n15297), .C2(n20939), .A(n15277), .B(n15276), .ZN(
        P1_U3085) );
  NAND2_X1 U18552 ( .A1(n15288), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n15282) );
  OAI22_X1 U18553 ( .A1(n15279), .A2(n15291), .B1(n15290), .B2(n15278), .ZN(
        n15280) );
  AOI21_X1 U18554 ( .B1(n15294), .B2(n20942), .A(n15280), .ZN(n15281) );
  OAI211_X1 U18555 ( .C1(n15297), .C2(n20945), .A(n15282), .B(n15281), .ZN(
        P1_U3086) );
  NAND2_X1 U18556 ( .A1(n15288), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n15287) );
  OAI22_X1 U18557 ( .A1(n15284), .A2(n15291), .B1(n15290), .B2(n15283), .ZN(
        n15285) );
  AOI21_X1 U18558 ( .B1(n15294), .B2(n20948), .A(n15285), .ZN(n15286) );
  OAI211_X1 U18559 ( .C1(n15297), .C2(n20951), .A(n15287), .B(n15286), .ZN(
        P1_U3087) );
  NAND2_X1 U18560 ( .A1(n15288), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n15296) );
  OAI22_X1 U18561 ( .A1(n15292), .A2(n15291), .B1(n15290), .B2(n15289), .ZN(
        n15293) );
  AOI21_X1 U18562 ( .B1(n15294), .B2(n20955), .A(n15293), .ZN(n15295) );
  OAI211_X1 U18563 ( .C1(n15297), .C2(n20960), .A(n15296), .B(n15295), .ZN(
        P1_U3088) );
  OAI21_X1 U18564 ( .B1(n10451), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20503), 
        .ZN(n15298) );
  NAND3_X1 U18565 ( .A1(n15299), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n15298), 
        .ZN(n15301) );
  OAI22_X1 U18566 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17082), .B1(n20509), 
        .B2(n20491), .ZN(n15300) );
  NAND2_X1 U18567 ( .A1(n15301), .A2(n15300), .ZN(n15304) );
  AOI21_X1 U18568 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n17077), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n15302) );
  AOI211_X1 U18569 ( .C1(n17069), .C2(n19900), .A(n15302), .B(n19599), .ZN(
        n15303) );
  MUX2_X1 U18570 ( .A(n15304), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n15303), 
        .Z(P2_U3610) );
  NAND2_X1 U18571 ( .A1(n12798), .A2(n15843), .ZN(n15306) );
  AND2_X1 U18572 ( .A1(n15307), .A2(n15306), .ZN(n15845) );
  NOR2_X1 U18573 ( .A1(n15479), .A2(n15845), .ZN(n19661) );
  AND2_X1 U18574 ( .A1(n15307), .A2(n19655), .ZN(n15308) );
  OR2_X1 U18575 ( .A1(n15308), .A2(n15310), .ZN(n19660) );
  NOR2_X1 U18576 ( .A1(n15310), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15311) );
  OR2_X1 U18577 ( .A1(n15309), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15312) );
  NAND2_X1 U18578 ( .A1(n15314), .A2(n15312), .ZN(n19642) );
  NAND2_X1 U18579 ( .A1(n15314), .A2(n15313), .ZN(n15315) );
  NAND2_X1 U18580 ( .A1(n15316), .A2(n15315), .ZN(n15793) );
  INV_X1 U18581 ( .A(n15793), .ZN(n15447) );
  AND2_X1 U18582 ( .A1(n15316), .A2(n15779), .ZN(n15317) );
  NOR2_X1 U18583 ( .A1(n15318), .A2(n15317), .ZN(n15782) );
  INV_X1 U18584 ( .A(n15782), .ZN(n19628) );
  OAI21_X1 U18585 ( .B1(n19629), .B2(n9934), .A(n19628), .ZN(n15431) );
  NOR2_X1 U18586 ( .A1(n15318), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15319) );
  OR2_X1 U18587 ( .A1(n15320), .A2(n15319), .ZN(n15769) );
  INV_X1 U18588 ( .A(n15769), .ZN(n15432) );
  AOI21_X1 U18589 ( .B1(n15431), .B2(n19753), .A(n15432), .ZN(n15415) );
  OR2_X1 U18590 ( .A1(n15320), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15321) );
  NAND2_X1 U18591 ( .A1(n15322), .A2(n15321), .ZN(n15757) );
  OAI21_X1 U18592 ( .B1(n15415), .B2(n9934), .A(n15757), .ZN(n15417) );
  NAND2_X1 U18593 ( .A1(n15322), .A2(n15734), .ZN(n15323) );
  AND2_X1 U18594 ( .A1(n15324), .A2(n15323), .ZN(n16479) );
  AOI21_X1 U18595 ( .B1(n15417), .B2(n19753), .A(n16479), .ZN(n16482) );
  NAND2_X1 U18596 ( .A1(n15324), .A2(n15408), .ZN(n15325) );
  NAND2_X1 U18597 ( .A1(n15326), .A2(n15325), .ZN(n15724) );
  OAI21_X1 U18598 ( .B1(n16482), .B2(n9934), .A(n15724), .ZN(n15403) );
  AND2_X1 U18599 ( .A1(n15326), .A2(n15716), .ZN(n15327) );
  NOR2_X1 U18600 ( .A1(n15329), .A2(n15327), .ZN(n16889) );
  AOI21_X1 U18601 ( .B1(n15403), .B2(n19753), .A(n16889), .ZN(n16868) );
  OR2_X1 U18602 ( .A1(n15329), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15330) );
  NAND2_X1 U18603 ( .A1(n15328), .A2(n15330), .ZN(n16869) );
  OAI21_X1 U18604 ( .B1(n16868), .B2(n9934), .A(n16869), .ZN(n16860) );
  NAND2_X1 U18605 ( .A1(n15328), .A2(n15700), .ZN(n15331) );
  AND2_X1 U18606 ( .A1(n15332), .A2(n15331), .ZN(n16861) );
  AND2_X1 U18607 ( .A1(n15332), .A2(n15690), .ZN(n15333) );
  NOR2_X1 U18608 ( .A1(n15335), .A2(n15333), .ZN(n15693) );
  INV_X1 U18609 ( .A(n15693), .ZN(n15334) );
  NOR2_X1 U18610 ( .A1(n15335), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15336) );
  OR2_X1 U18611 ( .A1(n10957), .A2(n15336), .ZN(n15684) );
  INV_X1 U18612 ( .A(n15684), .ZN(n15377) );
  XNOR2_X1 U18613 ( .A(n15337), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15670) );
  INV_X1 U18614 ( .A(n15670), .ZN(n15338) );
  NAND2_X1 U18615 ( .A1(n15517), .A2(n15338), .ZN(n15358) );
  INV_X1 U18616 ( .A(n15339), .ZN(n15345) );
  NOR2_X1 U18617 ( .A1(n17075), .A2(n16898), .ZN(n15340) );
  AOI22_X1 U18618 ( .A1(n15341), .A2(n15340), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19732), .ZN(n15343) );
  NAND2_X1 U18619 ( .A1(n19652), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15342) );
  OAI211_X1 U18620 ( .C1(n19797), .C2(n19726), .A(n15343), .B(n15342), .ZN(
        n15344) );
  AOI21_X1 U18621 ( .B1(n15345), .B2(n19734), .A(n15344), .ZN(n15347) );
  OR2_X1 U18622 ( .A1(n16899), .A2(n19748), .ZN(n15346) );
  OAI211_X1 U18623 ( .C1(n15348), .C2(n15358), .A(n15347), .B(n15346), .ZN(
        P2_U2824) );
  INV_X1 U18624 ( .A(n15348), .ZN(n15359) );
  NOR2_X1 U18625 ( .A1(n15348), .A2(n19730), .ZN(n15349) );
  OAI21_X1 U18626 ( .B1(n15349), .B2(n15465), .A(n15670), .ZN(n15357) );
  NAND2_X1 U18627 ( .A1(n15938), .A2(n19743), .ZN(n15351) );
  AOI22_X1 U18628 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19732), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19652), .ZN(n15350) );
  OAI211_X1 U18629 ( .C1(n19683), .C2(n15352), .A(n15351), .B(n15350), .ZN(
        n15354) );
  NOR2_X1 U18630 ( .A1(n15937), .A2(n19748), .ZN(n15353) );
  AOI211_X1 U18631 ( .C1(n19734), .C2(n15355), .A(n15354), .B(n15353), .ZN(
        n15356) );
  OAI211_X1 U18632 ( .C1(n15359), .C2(n15358), .A(n15357), .B(n15356), .ZN(
        P2_U2825) );
  AOI21_X1 U18633 ( .B1(n9931), .B2(n9928), .A(n19730), .ZN(n15361) );
  OAI21_X1 U18634 ( .B1(n15361), .B2(n15465), .A(n15348), .ZN(n15372) );
  OR2_X1 U18635 ( .A1(n15362), .A2(n15363), .ZN(n15364) );
  NAND2_X1 U18636 ( .A1(n15957), .A2(n19743), .ZN(n15367) );
  AOI22_X1 U18637 ( .A1(n19652), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19732), .ZN(n15366) );
  OAI211_X1 U18638 ( .C1(n19683), .C2(n15368), .A(n15367), .B(n15366), .ZN(
        n15369) );
  AOI21_X1 U18639 ( .B1(n15370), .B2(n19734), .A(n15369), .ZN(n15371) );
  OAI211_X1 U18640 ( .C1(n19748), .C2(n15960), .A(n15372), .B(n15371), .ZN(
        P2_U2826) );
  INV_X1 U18641 ( .A(n9661), .ZN(n15375) );
  INV_X1 U18642 ( .A(n15373), .ZN(n15374) );
  AOI21_X1 U18643 ( .B1(n15376), .B2(n15377), .A(n19730), .ZN(n15378) );
  OAI21_X1 U18644 ( .B1(n15465), .B2(n15378), .A(n9931), .ZN(n15387) );
  NOR2_X1 U18645 ( .A1(n15379), .A2(n15380), .ZN(n15381) );
  OR2_X1 U18646 ( .A1(n15362), .A2(n15381), .ZN(n15965) );
  AOI22_X1 U18647 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19732), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19652), .ZN(n15382) );
  OAI21_X1 U18648 ( .B1(n19726), .B2(n15965), .A(n15382), .ZN(n15385) );
  NOR2_X1 U18649 ( .A1(n15383), .A2(n19684), .ZN(n15384) );
  AOI211_X1 U18650 ( .C1(P2_EBX_REG_28__SCAN_IN), .C2(n19744), .A(n15385), .B(
        n15384), .ZN(n15386) );
  OAI211_X1 U18651 ( .C1(n19748), .C2(n15969), .A(n15387), .B(n15386), .ZN(
        P2_U2827) );
  OAI21_X1 U18652 ( .B1(n15540), .B2(n15388), .A(n9661), .ZN(n15983) );
  INV_X1 U18653 ( .A(n15389), .ZN(n16863) );
  AOI21_X1 U18654 ( .B1(n16863), .B2(n15693), .A(n19730), .ZN(n15390) );
  OAI21_X1 U18655 ( .B1(n15390), .B2(n15465), .A(n15376), .ZN(n15400) );
  INV_X1 U18656 ( .A(n15391), .ZN(n15398) );
  INV_X1 U18657 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n15396) );
  AND2_X1 U18658 ( .A1(n15611), .A2(n15392), .ZN(n15393) );
  NOR2_X1 U18659 ( .A1(n15379), .A2(n15393), .ZN(n15980) );
  OAI22_X1 U18660 ( .A1(n15690), .A2(n19654), .B1(n20551), .B2(n19737), .ZN(
        n15394) );
  AOI21_X1 U18661 ( .B1(n15980), .B2(n19743), .A(n15394), .ZN(n15395) );
  OAI21_X1 U18662 ( .B1(n19683), .B2(n15396), .A(n15395), .ZN(n15397) );
  AOI21_X1 U18663 ( .B1(n15398), .B2(n19734), .A(n15397), .ZN(n15399) );
  OAI211_X1 U18664 ( .C1(n19748), .C2(n15983), .A(n15400), .B(n15399), .ZN(
        P2_U2828) );
  INV_X1 U18665 ( .A(n16482), .ZN(n15402) );
  INV_X1 U18666 ( .A(n15724), .ZN(n15401) );
  AOI21_X1 U18667 ( .B1(n15402), .B2(n15401), .A(n19730), .ZN(n15404) );
  OAI21_X1 U18668 ( .B1(n15404), .B2(n15465), .A(n15403), .ZN(n15413) );
  OR2_X1 U18669 ( .A1(n9687), .A2(n15405), .ZN(n15406) );
  AND2_X1 U18670 ( .A1(n15556), .A2(n15406), .ZN(n16900) );
  INV_X1 U18671 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16903) );
  AOI21_X1 U18672 ( .B1(n15407), .B2(n16041), .A(n10161), .ZN(n16031) );
  OAI22_X1 U18673 ( .A1(n19737), .A2(n20542), .B1(n19654), .B2(n15408), .ZN(
        n15409) );
  AOI21_X1 U18674 ( .B1(n16031), .B2(n19743), .A(n15409), .ZN(n15410) );
  OAI21_X1 U18675 ( .B1(n19683), .B2(n16903), .A(n15410), .ZN(n15411) );
  AOI21_X1 U18676 ( .B1(n16900), .B2(n19692), .A(n15411), .ZN(n15412) );
  OAI211_X1 U18677 ( .C1(n19684), .C2(n15414), .A(n15413), .B(n15412), .ZN(
        P2_U2832) );
  INV_X1 U18678 ( .A(n15415), .ZN(n15433) );
  INV_X1 U18679 ( .A(n15757), .ZN(n15416) );
  AOI21_X1 U18680 ( .B1(n15433), .B2(n15416), .A(n19730), .ZN(n15418) );
  OAI21_X1 U18681 ( .B1(n15418), .B2(n15465), .A(n15417), .ZN(n15429) );
  NAND2_X1 U18682 ( .A1(n15419), .A2(n15420), .ZN(n15421) );
  AND2_X1 U18683 ( .A1(n15736), .A2(n15421), .ZN(n16061) );
  OR2_X1 U18684 ( .A1(n15439), .A2(n15422), .ZN(n15424) );
  NAND2_X1 U18685 ( .A1(n15424), .A2(n15423), .ZN(n16063) );
  AOI22_X1 U18686 ( .A1(n19652), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19732), .ZN(n15426) );
  NAND2_X1 U18687 ( .A1(n19744), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15425) );
  OAI211_X1 U18688 ( .C1(n19726), .C2(n16063), .A(n15426), .B(n15425), .ZN(
        n15427) );
  AOI21_X1 U18689 ( .B1(n16061), .B2(n19692), .A(n15427), .ZN(n15428) );
  OAI211_X1 U18690 ( .C1(n19684), .C2(n15430), .A(n15429), .B(n15428), .ZN(
        P2_U2834) );
  AOI21_X1 U18691 ( .B1(n15431), .B2(n15432), .A(n19730), .ZN(n15434) );
  OAI21_X1 U18692 ( .B1(n15465), .B2(n15434), .A(n15433), .ZN(n15444) );
  OR2_X1 U18693 ( .A1(n15569), .A2(n15435), .ZN(n15436) );
  NAND2_X1 U18694 ( .A1(n15419), .A2(n15436), .ZN(n16909) );
  INV_X1 U18695 ( .A(n16909), .ZN(n16073) );
  NOR2_X1 U18696 ( .A1(n15652), .A2(n15437), .ZN(n15438) );
  OR2_X1 U18697 ( .A1(n15439), .A2(n15438), .ZN(n16922) );
  AOI22_X1 U18698 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19732), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19652), .ZN(n15441) );
  NAND2_X1 U18699 ( .A1(n19744), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15440) );
  OAI211_X1 U18700 ( .C1(n19726), .C2(n16922), .A(n15441), .B(n15440), .ZN(
        n15442) );
  AOI21_X1 U18701 ( .B1(n16073), .B2(n19692), .A(n15442), .ZN(n15443) );
  OAI211_X1 U18702 ( .C1(n19684), .C2(n15445), .A(n15444), .B(n15443), .ZN(
        P2_U2835) );
  INV_X1 U18703 ( .A(n15446), .ZN(n15461) );
  AOI21_X1 U18704 ( .B1(n19644), .B2(n15447), .A(n19730), .ZN(n15449) );
  INV_X1 U18705 ( .A(n19629), .ZN(n15448) );
  OAI21_X1 U18706 ( .B1(n15465), .B2(n15449), .A(n15448), .ZN(n15460) );
  NAND2_X1 U18707 ( .A1(n15578), .A2(n15450), .ZN(n15451) );
  NAND2_X1 U18708 ( .A1(n15571), .A2(n15451), .ZN(n16916) );
  INV_X1 U18709 ( .A(n16916), .ZN(n16099) );
  NAND2_X1 U18710 ( .A1(n15453), .A2(n15452), .ZN(n15454) );
  NAND2_X1 U18711 ( .A1(n15651), .A2(n15454), .ZN(n16102) );
  INV_X1 U18712 ( .A(n16102), .ZN(n16929) );
  AOI21_X1 U18713 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19732), .A(
        n19903), .ZN(n15455) );
  OAI21_X1 U18714 ( .B1(n19737), .B2(n15792), .A(n15455), .ZN(n15456) );
  AOI21_X1 U18715 ( .B1(n16929), .B2(n19743), .A(n15456), .ZN(n15457) );
  OAI21_X1 U18716 ( .B1(n19683), .B2(n16913), .A(n15457), .ZN(n15458) );
  AOI21_X1 U18717 ( .B1(n16099), .B2(n19692), .A(n15458), .ZN(n15459) );
  OAI211_X1 U18718 ( .C1(n19684), .C2(n15461), .A(n15460), .B(n15459), .ZN(
        P2_U2837) );
  INV_X1 U18719 ( .A(n15462), .ZN(n15478) );
  AOI21_X1 U18720 ( .B1(n19662), .B2(n10193), .A(n19730), .ZN(n15464) );
  INV_X1 U18721 ( .A(n19643), .ZN(n15463) );
  OAI21_X1 U18722 ( .B1(n15465), .B2(n15464), .A(n15463), .ZN(n15477) );
  OR2_X1 U18723 ( .A1(n15467), .A2(n15468), .ZN(n15469) );
  NAND2_X1 U18724 ( .A1(n15466), .A2(n15469), .ZN(n19767) );
  NOR2_X1 U18725 ( .A1(n19767), .A2(n19748), .ZN(n15475) );
  NAND2_X1 U18726 ( .A1(n15470), .A2(n16962), .ZN(n15471) );
  NAND2_X1 U18727 ( .A1(n15471), .A2(n10156), .ZN(n19805) );
  OAI21_X1 U18728 ( .B1(n19654), .B2(n15819), .A(n19736), .ZN(n15472) );
  AOI21_X1 U18729 ( .B1(n19652), .B2(P2_REIP_REG_16__SCAN_IN), .A(n15472), 
        .ZN(n15473) );
  OAI21_X1 U18730 ( .B1(n19726), .B2(n19805), .A(n15473), .ZN(n15474) );
  AOI211_X1 U18731 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19744), .A(n15475), .B(
        n15474), .ZN(n15476) );
  OAI211_X1 U18732 ( .C1(n19684), .C2(n15478), .A(n15477), .B(n15476), .ZN(
        P2_U2839) );
  OAI21_X1 U18733 ( .B1(n19730), .B2(n15479), .A(n19665), .ZN(n15484) );
  AOI21_X1 U18734 ( .B1(n15481), .B2(n15480), .A(n16963), .ZN(n16981) );
  INV_X1 U18735 ( .A(n16981), .ZN(n19815) );
  OAI21_X1 U18736 ( .B1(n15482), .B2(n9685), .A(n15583), .ZN(n19772) );
  OAI22_X1 U18737 ( .A1(n19726), .A2(n19815), .B1(n19772), .B2(n19748), .ZN(
        n15483) );
  AOI21_X1 U18738 ( .B1(n15484), .B2(n15845), .A(n15483), .ZN(n15489) );
  AOI22_X1 U18739 ( .A1(n15485), .A2(n19734), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19744), .ZN(n15486) );
  OAI211_X1 U18740 ( .C1(n15842), .C2(n19737), .A(n15486), .B(n19736), .ZN(
        n15487) );
  AOI21_X1 U18741 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19732), .A(
        n15487), .ZN(n15488) );
  OAI211_X1 U18742 ( .C1(n15845), .C2(n15490), .A(n15489), .B(n15488), .ZN(
        P2_U2841) );
  INV_X1 U18743 ( .A(n15491), .ZN(n15867) );
  OAI21_X1 U18744 ( .B1(n19730), .B2(n15492), .A(n19665), .ZN(n15504) );
  AOI21_X1 U18745 ( .B1(n15494), .B2(n15493), .A(n12845), .ZN(n16134) );
  OAI21_X1 U18746 ( .B1(n15497), .B2(n15496), .A(n15495), .ZN(n19777) );
  AOI22_X1 U18747 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19732), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19652), .ZN(n15498) );
  OAI211_X1 U18748 ( .C1(n19777), .C2(n19748), .A(n15498), .B(n19736), .ZN(
        n15499) );
  AOI21_X1 U18749 ( .B1(n19743), .B2(n16134), .A(n15499), .ZN(n15501) );
  NAND2_X1 U18750 ( .A1(n19744), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15500) );
  OAI211_X1 U18751 ( .C1(n19684), .C2(n15502), .A(n15501), .B(n15500), .ZN(
        n15503) );
  AOI21_X1 U18752 ( .B1(n15504), .B2(n15867), .A(n15503), .ZN(n15505) );
  OAI21_X1 U18753 ( .B1(n15867), .B2(n15506), .A(n15505), .ZN(P2_U2843) );
  OAI22_X1 U18754 ( .A1(n19684), .A2(n15926), .B1(n10475), .B2(n19737), .ZN(
        n15509) );
  NOR2_X1 U18755 ( .A1(n19683), .A2(n15507), .ZN(n15508) );
  AOI211_X1 U18756 ( .C1(n15510), .C2(n19743), .A(n15509), .B(n15508), .ZN(
        n15513) );
  NAND2_X1 U18757 ( .A1(n16222), .A2(n15511), .ZN(n15512) );
  OAI211_X1 U18758 ( .C1(n19748), .C2(n17014), .A(n15513), .B(n15512), .ZN(
        n15516) );
  AOI21_X1 U18759 ( .B1(n19665), .B2(n19654), .A(n15514), .ZN(n15515) );
  AOI211_X1 U18760 ( .C1(n15518), .C2(n15517), .A(n15516), .B(n15515), .ZN(
        n15519) );
  INV_X1 U18761 ( .A(n15519), .ZN(P2_U2855) );
  OR2_X1 U18762 ( .A1(n15521), .A2(n15520), .ZN(n15592) );
  NAND3_X1 U18763 ( .A1(n15592), .A2(n15522), .A3(n19793), .ZN(n15524) );
  NAND2_X1 U18764 ( .A1(n19796), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15523) );
  OAI211_X1 U18765 ( .C1(n19796), .C2(n15960), .A(n15524), .B(n15523), .ZN(
        P2_U2858) );
  NOR2_X1 U18766 ( .A1(n15526), .A2(n15525), .ZN(n15528) );
  XNOR2_X1 U18767 ( .A(n15528), .B(n15527), .ZN(n15601) );
  NAND2_X1 U18768 ( .A1(n15601), .A2(n19793), .ZN(n15530) );
  NAND2_X1 U18769 ( .A1(n19796), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15529) );
  OAI211_X1 U18770 ( .C1(n19796), .C2(n15969), .A(n15530), .B(n15529), .ZN(
        P2_U2859) );
  OAI21_X1 U18771 ( .B1(n9655), .B2(n15532), .A(n15531), .ZN(n15607) );
  NOR2_X1 U18772 ( .A1(n15983), .A2(n19796), .ZN(n15533) );
  AOI21_X1 U18773 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19796), .A(n15533), .ZN(
        n15534) );
  OAI21_X1 U18774 ( .B1(n15607), .B2(n19788), .A(n15534), .ZN(P2_U2860) );
  OAI21_X1 U18775 ( .B1(n15535), .B2(n15537), .A(n15536), .ZN(n15617) );
  NOR2_X1 U18776 ( .A1(n15548), .A2(n15538), .ZN(n15539) );
  OR2_X1 U18777 ( .A1(n15540), .A2(n15539), .ZN(n16858) );
  NOR2_X1 U18778 ( .A1(n16858), .A2(n19796), .ZN(n15541) );
  AOI21_X1 U18779 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n19796), .A(n15541), .ZN(
        n15542) );
  OAI21_X1 U18780 ( .B1(n15617), .B2(n19788), .A(n15542), .ZN(P2_U2861) );
  OAI21_X1 U18781 ( .B1(n15543), .B2(n15545), .A(n15544), .ZN(n15625) );
  NAND2_X1 U18782 ( .A1(n19796), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15550) );
  AND2_X1 U18783 ( .A1(n15558), .A2(n15546), .ZN(n15547) );
  NOR2_X1 U18784 ( .A1(n15548), .A2(n15547), .ZN(n16874) );
  NAND2_X1 U18785 ( .A1(n16874), .A2(n19784), .ZN(n15549) );
  OAI211_X1 U18786 ( .C1(n15625), .C2(n19788), .A(n15550), .B(n15549), .ZN(
        P2_U2862) );
  AOI21_X1 U18787 ( .B1(n9695), .B2(n15552), .A(n15551), .ZN(n15553) );
  XOR2_X1 U18788 ( .A(n15554), .B(n15553), .Z(n15635) );
  NAND2_X1 U18789 ( .A1(n15556), .A2(n15555), .ZN(n15557) );
  NAND2_X1 U18790 ( .A1(n15558), .A2(n15557), .ZN(n16888) );
  NOR2_X1 U18791 ( .A1(n16888), .A2(n19796), .ZN(n15559) );
  AOI21_X1 U18792 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n19796), .A(n15559), .ZN(
        n15560) );
  OAI21_X1 U18793 ( .B1(n15635), .B2(n19788), .A(n15560), .ZN(P2_U2863) );
  OAI21_X1 U18794 ( .B1(n15561), .B2(n15563), .A(n15562), .ZN(n15649) );
  NOR2_X1 U18795 ( .A1(n19784), .A2(n15564), .ZN(n15565) );
  AOI21_X1 U18796 ( .B1(n16061), .B2(n19784), .A(n15565), .ZN(n15566) );
  OAI21_X1 U18797 ( .B1(n15649), .B2(n19788), .A(n15566), .ZN(P2_U2866) );
  OAI21_X1 U18798 ( .B1(n9689), .B2(n15568), .A(n15567), .ZN(n15660) );
  INV_X1 U18799 ( .A(n15569), .ZN(n15573) );
  NAND2_X1 U18800 ( .A1(n15571), .A2(n15570), .ZN(n15572) );
  NAND2_X1 U18801 ( .A1(n15573), .A2(n15572), .ZN(n19627) );
  NOR2_X1 U18802 ( .A1(n19627), .A2(n19796), .ZN(n15574) );
  AOI21_X1 U18803 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19796), .A(n15574), .ZN(
        n15575) );
  OAI21_X1 U18804 ( .B1(n15660), .B2(n19788), .A(n15575), .ZN(P2_U2868) );
  NAND2_X1 U18805 ( .A1(n15466), .A2(n15576), .ZN(n15577) );
  AND2_X1 U18806 ( .A1(n15578), .A2(n15577), .ZN(n15812) );
  INV_X1 U18807 ( .A(n15812), .ZN(n19641) );
  NAND2_X1 U18808 ( .A1(n15579), .A2(n19793), .ZN(n15581) );
  NAND2_X1 U18809 ( .A1(n19796), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15580) );
  OAI211_X1 U18810 ( .C1(n19641), .C2(n19796), .A(n15581), .B(n15580), .ZN(
        P2_U2870) );
  AND2_X1 U18811 ( .A1(n15583), .A2(n15582), .ZN(n15584) );
  NOR2_X1 U18812 ( .A1(n15467), .A2(n15584), .ZN(n19657) );
  INV_X1 U18813 ( .A(n19657), .ZN(n16970) );
  NOR2_X1 U18814 ( .A1(n19796), .A2(n16970), .ZN(n15590) );
  OR2_X1 U18815 ( .A1(n19768), .A2(n19769), .ZN(n15587) );
  AND2_X1 U18816 ( .A1(n15586), .A2(n15585), .ZN(n19764) );
  AOI211_X1 U18817 ( .C1(n15588), .C2(n15587), .A(n19788), .B(n19764), .ZN(
        n15589) );
  AOI211_X1 U18818 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19796), .A(n15590), .B(
        n15589), .ZN(n15591) );
  INV_X1 U18819 ( .A(n15591), .ZN(P2_U2872) );
  NAND3_X1 U18820 ( .A1(n15592), .A2(n15522), .A3(n19848), .ZN(n15597) );
  OAI22_X1 U18821 ( .A1(n15640), .A2(n19816), .B1(n19834), .B2(n15593), .ZN(
        n15594) );
  AOI21_X1 U18822 ( .B1(n19859), .B2(n15957), .A(n15594), .ZN(n15596) );
  AOI22_X1 U18823 ( .A1(n19804), .A2(BUF2_REG_29__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15595) );
  NAND3_X1 U18824 ( .A1(n15597), .A2(n15596), .A3(n15595), .ZN(P2_U2890) );
  AOI22_X1 U18825 ( .A1(n19804), .A2(BUF2_REG_28__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15599) );
  AOI22_X1 U18826 ( .A1(n19802), .A2(n19818), .B1(n19858), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15598) );
  OAI211_X1 U18827 ( .C1(n15657), .C2(n15965), .A(n15599), .B(n15598), .ZN(
        n15600) );
  AOI21_X1 U18828 ( .B1(n15601), .B2(n19848), .A(n15600), .ZN(n15602) );
  INV_X1 U18829 ( .A(n15602), .ZN(P2_U2891) );
  OAI22_X1 U18830 ( .A1(n15640), .A2(n19821), .B1(n19834), .B2(n15603), .ZN(
        n15604) );
  AOI21_X1 U18831 ( .B1(n19859), .B2(n15980), .A(n15604), .ZN(n15606) );
  AOI22_X1 U18832 ( .A1(n19804), .A2(BUF2_REG_27__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15605) );
  OAI211_X1 U18833 ( .C1(n15607), .C2(n19863), .A(n15606), .B(n15605), .ZN(
        P2_U2892) );
  NAND2_X1 U18834 ( .A1(n15608), .A2(n15609), .ZN(n15610) );
  AND2_X1 U18835 ( .A1(n15611), .A2(n15610), .ZN(n16856) );
  INV_X1 U18836 ( .A(n19823), .ZN(n15613) );
  OAI22_X1 U18837 ( .A1(n15640), .A2(n15613), .B1(n19834), .B2(n15612), .ZN(
        n15614) );
  AOI21_X1 U18838 ( .B1(n19859), .B2(n16856), .A(n15614), .ZN(n15616) );
  AOI22_X1 U18839 ( .A1(n19804), .A2(BUF2_REG_26__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15615) );
  OAI211_X1 U18840 ( .C1(n15617), .C2(n19863), .A(n15616), .B(n15615), .ZN(
        P2_U2893) );
  OR2_X1 U18841 ( .A1(n15626), .A2(n15618), .ZN(n15619) );
  NAND2_X1 U18842 ( .A1(n15608), .A2(n15619), .ZN(n16882) );
  INV_X1 U18843 ( .A(n16882), .ZN(n15622) );
  OAI22_X1 U18844 ( .A1(n15640), .A2(n19826), .B1(n19834), .B2(n15620), .ZN(
        n15621) );
  AOI21_X1 U18845 ( .B1(n19859), .B2(n15622), .A(n15621), .ZN(n15624) );
  AOI22_X1 U18846 ( .A1(n19804), .A2(BUF2_REG_25__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15623) );
  OAI211_X1 U18847 ( .C1(n15625), .C2(n19863), .A(n15624), .B(n15623), .ZN(
        P2_U2894) );
  INV_X1 U18848 ( .A(n15626), .ZN(n15630) );
  NAND2_X1 U18849 ( .A1(n15628), .A2(n15627), .ZN(n15629) );
  NAND2_X1 U18850 ( .A1(n15630), .A2(n15629), .ZN(n16897) );
  INV_X1 U18851 ( .A(n16897), .ZN(n16016) );
  OAI22_X1 U18852 ( .A1(n15640), .A2(n19829), .B1(n19834), .B2(n15631), .ZN(
        n15632) );
  AOI21_X1 U18853 ( .B1(n19859), .B2(n16016), .A(n15632), .ZN(n15634) );
  AOI22_X1 U18854 ( .A1(n19804), .A2(BUF2_REG_24__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15633) );
  OAI211_X1 U18855 ( .C1(n15635), .C2(n19863), .A(n15634), .B(n15633), .ZN(
        P2_U2895) );
  AOI21_X1 U18856 ( .B1(n15638), .B2(n15637), .A(n15636), .ZN(n16901) );
  INV_X1 U18857 ( .A(n16901), .ZN(n15644) );
  OAI22_X1 U18858 ( .A1(n15640), .A2(n19831), .B1(n19834), .B2(n15639), .ZN(
        n15641) );
  AOI21_X1 U18859 ( .B1(n19859), .B2(n16031), .A(n15641), .ZN(n15643) );
  AOI22_X1 U18860 ( .A1(n19804), .A2(BUF2_REG_23__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15642) );
  OAI211_X1 U18861 ( .C1(n15644), .C2(n19863), .A(n15643), .B(n15642), .ZN(
        P2_U2896) );
  AOI22_X1 U18862 ( .A1(n19804), .A2(BUF2_REG_21__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15646) );
  AOI22_X1 U18863 ( .A1(n19802), .A2(n19837), .B1(n19858), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15645) );
  OAI211_X1 U18864 ( .C1(n15657), .C2(n16063), .A(n15646), .B(n15645), .ZN(
        n15647) );
  INV_X1 U18865 ( .A(n15647), .ZN(n15648) );
  OAI21_X1 U18866 ( .B1(n15649), .B2(n19863), .A(n15648), .ZN(P2_U2898) );
  AND2_X1 U18867 ( .A1(n15651), .A2(n15650), .ZN(n15653) );
  OR2_X1 U18868 ( .A1(n15653), .A2(n15652), .ZN(n19636) );
  AOI22_X1 U18869 ( .A1(n19804), .A2(BUF2_REG_19__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U18870 ( .A1(n19802), .A2(n15654), .B1(n19858), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15655) );
  OAI211_X1 U18871 ( .C1(n15657), .C2(n19636), .A(n15656), .B(n15655), .ZN(
        n15658) );
  INV_X1 U18872 ( .A(n15658), .ZN(n15659) );
  OAI21_X1 U18873 ( .B1(n15660), .B2(n19863), .A(n15659), .ZN(P2_U2900) );
  NAND2_X1 U18874 ( .A1(n15662), .A2(n15661), .ZN(n15667) );
  INV_X1 U18875 ( .A(n15663), .ZN(n15664) );
  NOR2_X1 U18876 ( .A1(n15665), .A2(n15664), .ZN(n15666) );
  XNOR2_X1 U18877 ( .A(n15667), .B(n15666), .ZN(n15950) );
  XNOR2_X1 U18878 ( .A(n15668), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15947) );
  NAND2_X1 U18879 ( .A1(n19903), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15940) );
  OAI21_X1 U18880 ( .B1(n16950), .B2(n9938), .A(n15940), .ZN(n15669) );
  AOI21_X1 U18881 ( .B1(n15670), .B2(n16942), .A(n15669), .ZN(n15671) );
  OAI21_X1 U18882 ( .B1(n15937), .B2(n13859), .A(n15671), .ZN(n15672) );
  AOI21_X1 U18883 ( .B1(n15947), .B2(n15933), .A(n15672), .ZN(n15673) );
  OAI21_X1 U18884 ( .B1(n15950), .B2(n16957), .A(n15673), .ZN(P2_U2984) );
  INV_X1 U18885 ( .A(n15676), .ZN(n15678) );
  OAI22_X1 U18886 ( .A1(n15689), .A2(n15970), .B1(n15678), .B2(n15677), .ZN(
        n15681) );
  XNOR2_X1 U18887 ( .A(n15679), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15680) );
  XNOR2_X1 U18888 ( .A(n15681), .B(n15680), .ZN(n15978) );
  AOI21_X1 U18889 ( .B1(n15954), .B2(n15989), .A(n15683), .ZN(n15975) );
  NOR2_X1 U18890 ( .A1(n19736), .A2(n20552), .ZN(n15966) );
  NOR2_X1 U18891 ( .A1(n15684), .A2(n16952), .ZN(n15685) );
  AOI211_X1 U18892 ( .C1(n16954), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15966), .B(n15685), .ZN(n15686) );
  OAI21_X1 U18893 ( .B1(n15969), .B2(n13859), .A(n15686), .ZN(n15687) );
  AOI21_X1 U18894 ( .B1(n15975), .B2(n15933), .A(n15687), .ZN(n15688) );
  OAI21_X1 U18895 ( .B1(n15978), .B2(n16957), .A(n15688), .ZN(P2_U2986) );
  XNOR2_X1 U18896 ( .A(n15689), .B(n15970), .ZN(n15992) );
  NAND2_X1 U18897 ( .A1(n19903), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15982) );
  OAI21_X1 U18898 ( .B1(n16950), .B2(n15690), .A(n15982), .ZN(n15692) );
  NOR2_X1 U18899 ( .A1(n15983), .A2(n13859), .ZN(n15691) );
  AOI211_X1 U18900 ( .C1(n16942), .C2(n15693), .A(n15692), .B(n15691), .ZN(
        n15695) );
  NAND2_X1 U18901 ( .A1(n15697), .A2(n15970), .ZN(n15988) );
  NAND3_X1 U18902 ( .A1(n15989), .A2(n15933), .A3(n15988), .ZN(n15694) );
  OAI211_X1 U18903 ( .C1(n15992), .C2(n16957), .A(n15695), .B(n15694), .ZN(
        P2_U2987) );
  OR2_X1 U18904 ( .A1(n9675), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15696) );
  NAND2_X1 U18905 ( .A1(n15697), .A2(n15696), .ZN(n16004) );
  OAI21_X1 U18906 ( .B1(n15698), .B2(n15706), .A(n15705), .ZN(n15699) );
  XNOR2_X1 U18907 ( .A(n15699), .B(n9662), .ZN(n15993) );
  NAND2_X1 U18908 ( .A1(n15993), .A2(n15927), .ZN(n15704) );
  NAND2_X1 U18909 ( .A1(n19903), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15995) );
  OAI21_X1 U18910 ( .B1(n16950), .B2(n15700), .A(n15995), .ZN(n15702) );
  NOR2_X1 U18911 ( .A1(n16858), .A2(n13859), .ZN(n15701) );
  AOI211_X1 U18912 ( .C1(n16942), .C2(n16861), .A(n15702), .B(n15701), .ZN(
        n15703) );
  OAI211_X1 U18913 ( .C1(n16955), .C2(n16004), .A(n15704), .B(n15703), .ZN(
        P2_U2988) );
  NOR2_X1 U18914 ( .A1(n15706), .A2(n10066), .ZN(n15707) );
  XNOR2_X1 U18915 ( .A(n15698), .B(n15707), .ZN(n16014) );
  AOI21_X1 U18916 ( .B1(n15998), .B2(n15713), .A(n9675), .ZN(n16012) );
  NAND2_X1 U18917 ( .A1(n16874), .A2(n16946), .ZN(n15709) );
  NOR2_X1 U18918 ( .A1(n19736), .A2(n20546), .ZN(n16006) );
  AOI21_X1 U18919 ( .B1(n16954), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16006), .ZN(n15708) );
  OAI211_X1 U18920 ( .C1(n16952), .C2(n16869), .A(n15709), .B(n15708), .ZN(
        n15710) );
  AOI21_X1 U18921 ( .B1(n16012), .B2(n15933), .A(n15710), .ZN(n15711) );
  OAI21_X1 U18922 ( .B1(n16014), .B2(n16957), .A(n15711), .ZN(P2_U2989) );
  NAND2_X1 U18923 ( .A1(n15726), .A2(n21106), .ZN(n15712) );
  NAND2_X1 U18924 ( .A1(n15713), .A2(n15712), .ZN(n16024) );
  XNOR2_X1 U18925 ( .A(n15714), .B(n21106), .ZN(n15715) );
  XNOR2_X1 U18926 ( .A(n9680), .B(n15715), .ZN(n16015) );
  NAND2_X1 U18927 ( .A1(n16015), .A2(n15927), .ZN(n15720) );
  NAND2_X1 U18928 ( .A1(n19903), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16018) );
  OAI21_X1 U18929 ( .B1(n16950), .B2(n15716), .A(n16018), .ZN(n15718) );
  NOR2_X1 U18930 ( .A1(n16888), .A2(n13859), .ZN(n15717) );
  AOI211_X1 U18931 ( .C1(n16942), .C2(n16889), .A(n15718), .B(n15717), .ZN(
        n15719) );
  OAI211_X1 U18932 ( .C1(n16955), .C2(n16024), .A(n15720), .B(n15719), .ZN(
        P2_U2990) );
  XNOR2_X1 U18933 ( .A(n15721), .B(n15722), .ZN(n16038) );
  NOR2_X1 U18934 ( .A1(n19736), .A2(n20542), .ZN(n16030) );
  AOI21_X1 U18935 ( .B1(n16954), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16030), .ZN(n15723) );
  OAI21_X1 U18936 ( .B1(n15724), .B2(n16952), .A(n15723), .ZN(n15728) );
  INV_X1 U18937 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16050) );
  NOR2_X1 U18938 ( .A1(n15758), .A2(n16050), .ZN(n16046) );
  OAI21_X1 U18939 ( .B1(n16046), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15726), .ZN(n16025) );
  NOR2_X1 U18940 ( .A1(n16025), .A2(n16955), .ZN(n15727) );
  AOI211_X1 U18941 ( .C1(n16946), .C2(n16900), .A(n15728), .B(n15727), .ZN(
        n15729) );
  OAI21_X1 U18942 ( .B1(n16038), .B2(n16957), .A(n15729), .ZN(P2_U2991) );
  NAND2_X1 U18943 ( .A1(n9789), .A2(n15731), .ZN(n15732) );
  XNOR2_X1 U18944 ( .A(n9663), .B(n15732), .ZN(n16053) );
  OAI22_X1 U18945 ( .A1(n16950), .A2(n15734), .B1(n15733), .B2(n19736), .ZN(
        n15739) );
  AND2_X1 U18946 ( .A1(n15736), .A2(n15735), .ZN(n15737) );
  OR2_X1 U18947 ( .A1(n15737), .A2(n9687), .ZN(n16906) );
  NOR2_X1 U18948 ( .A1(n16906), .A2(n13859), .ZN(n15738) );
  AOI211_X1 U18949 ( .C1(n16942), .C2(n16479), .A(n15739), .B(n15738), .ZN(
        n15741) );
  NOR2_X1 U18950 ( .A1(n10844), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16047) );
  OR3_X1 U18951 ( .A1(n16047), .A2(n16046), .A3(n16955), .ZN(n15740) );
  OAI211_X1 U18952 ( .C1(n16053), .C2(n16957), .A(n15741), .B(n15740), .ZN(
        P2_U2992) );
  INV_X1 U18953 ( .A(n15743), .ZN(n15744) );
  INV_X1 U18954 ( .A(n15851), .ZN(n15745) );
  INV_X1 U18955 ( .A(n15825), .ZN(n15746) );
  INV_X1 U18956 ( .A(n15817), .ZN(n15747) );
  NOR2_X2 U18957 ( .A1(n15814), .A2(n15747), .ZN(n15800) );
  INV_X1 U18958 ( .A(n15776), .ZN(n15749) );
  NOR2_X1 U18959 ( .A1(n15753), .A2(n15752), .ZN(n15754) );
  XNOR2_X1 U18960 ( .A(n15755), .B(n15754), .ZN(n16068) );
  NOR2_X1 U18961 ( .A1(n19736), .A2(n20540), .ZN(n16060) );
  AOI21_X1 U18962 ( .B1(n16954), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16060), .ZN(n15756) );
  OAI21_X1 U18963 ( .B1(n15757), .B2(n16952), .A(n15756), .ZN(n15760) );
  OAI21_X1 U18964 ( .B1(n15767), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15758), .ZN(n16054) );
  NOR2_X1 U18965 ( .A1(n16054), .A2(n16955), .ZN(n15759) );
  AOI211_X1 U18966 ( .C1(n16946), .C2(n16061), .A(n15760), .B(n15759), .ZN(
        n15761) );
  OAI21_X1 U18967 ( .B1(n16068), .B2(n16957), .A(n15761), .ZN(P2_U2993) );
  NAND2_X1 U18968 ( .A1(n9677), .A2(n15762), .ZN(n15766) );
  NAND2_X1 U18969 ( .A1(n15764), .A2(n15763), .ZN(n15765) );
  XNOR2_X1 U18970 ( .A(n15766), .B(n15765), .ZN(n16080) );
  AOI21_X1 U18971 ( .B1(n16075), .B2(n16090), .A(n15767), .ZN(n16078) );
  NOR2_X1 U18972 ( .A1(n19736), .A2(n15768), .ZN(n16072) );
  NOR2_X1 U18973 ( .A1(n15769), .A2(n16952), .ZN(n15770) );
  AOI211_X1 U18974 ( .C1(n16954), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16072), .B(n15770), .ZN(n15771) );
  OAI21_X1 U18975 ( .B1(n13859), .B2(n16909), .A(n15771), .ZN(n15772) );
  AOI21_X1 U18976 ( .B1(n16078), .B2(n15933), .A(n15772), .ZN(n15773) );
  OAI21_X1 U18977 ( .B1(n16080), .B2(n16957), .A(n15773), .ZN(P2_U2994) );
  NAND2_X1 U18978 ( .A1(n15774), .A2(n15787), .ZN(n15778) );
  NAND2_X1 U18979 ( .A1(n15776), .A2(n15775), .ZN(n15777) );
  XNOR2_X1 U18980 ( .A(n15778), .B(n15777), .ZN(n16094) );
  NAND2_X1 U18981 ( .A1(n19903), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16082) );
  OAI21_X1 U18982 ( .B1(n16950), .B2(n15779), .A(n16082), .ZN(n15781) );
  NOR2_X1 U18983 ( .A1(n19627), .A2(n13859), .ZN(n15780) );
  AOI211_X1 U18984 ( .C1(n16942), .C2(n15782), .A(n15781), .B(n15780), .ZN(
        n15785) );
  INV_X1 U18985 ( .A(n15790), .ZN(n15783) );
  NAND2_X1 U18986 ( .A1(n15783), .A2(n16088), .ZN(n16091) );
  NAND3_X1 U18987 ( .A1(n16091), .A2(n15933), .A3(n16090), .ZN(n15784) );
  OAI211_X1 U18988 ( .C1(n16094), .C2(n16957), .A(n15785), .B(n15784), .ZN(
        P2_U2995) );
  NAND2_X1 U18989 ( .A1(n15787), .A2(n15786), .ZN(n15788) );
  XNOR2_X1 U18990 ( .A(n15789), .B(n15788), .ZN(n16107) );
  NAND2_X1 U18991 ( .A1(n16171), .A2(n16096), .ZN(n15807) );
  AOI21_X1 U18992 ( .B1(n15791), .B2(n15807), .A(n15790), .ZN(n16105) );
  NOR2_X1 U18993 ( .A1(n19736), .A2(n15792), .ZN(n16098) );
  NOR2_X1 U18994 ( .A1(n16952), .A2(n15793), .ZN(n15794) );
  AOI211_X1 U18995 ( .C1(n16954), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16098), .B(n15794), .ZN(n15795) );
  OAI21_X1 U18996 ( .B1(n13859), .B2(n16916), .A(n15795), .ZN(n15796) );
  AOI21_X1 U18997 ( .B1(n16105), .B2(n15933), .A(n15796), .ZN(n15797) );
  OAI21_X1 U18998 ( .B1(n16107), .B2(n16957), .A(n15797), .ZN(P2_U2996) );
  NAND2_X1 U18999 ( .A1(n15799), .A2(n15798), .ZN(n15803) );
  INV_X1 U19000 ( .A(n15800), .ZN(n15815) );
  NAND2_X1 U19001 ( .A1(n15815), .A2(n15801), .ZN(n15802) );
  XOR2_X1 U19002 ( .A(n15803), .B(n15802), .Z(n16502) );
  NOR2_X1 U19003 ( .A1(n20534), .A2(n19736), .ZN(n15804) );
  AOI21_X1 U19004 ( .B1(n16954), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15804), .ZN(n15805) );
  OAI21_X1 U19005 ( .B1(n16952), .B2(n19642), .A(n15805), .ZN(n15811) );
  NAND2_X1 U19006 ( .A1(n16171), .A2(n15806), .ZN(n16111) );
  NOR2_X1 U19007 ( .A1(n16111), .A2(n16968), .ZN(n15829) );
  NAND2_X1 U19008 ( .A1(n15829), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16109) );
  INV_X1 U19009 ( .A(n15807), .ZN(n15808) );
  AOI211_X1 U19010 ( .C1(n16109), .C2(n15809), .A(n15808), .B(n16955), .ZN(
        n15810) );
  AOI211_X1 U19011 ( .C1(n16946), .C2(n15812), .A(n15811), .B(n15810), .ZN(
        n15813) );
  OAI21_X1 U19012 ( .B1(n16502), .B2(n16957), .A(n15813), .ZN(P2_U2997) );
  INV_X1 U19013 ( .A(n15814), .ZN(n15816) );
  OAI21_X1 U19014 ( .B1(n15817), .B2(n15816), .A(n15815), .ZN(n16119) );
  XNOR2_X1 U19015 ( .A(n15829), .B(n16498), .ZN(n15823) );
  NAND2_X1 U19016 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n19903), .ZN(n15818) );
  OAI21_X1 U19017 ( .B1(n16950), .B2(n15819), .A(n15818), .ZN(n15820) );
  AOI21_X1 U19018 ( .B1(n16942), .B2(n10193), .A(n15820), .ZN(n15821) );
  OAI21_X1 U19019 ( .B1(n13859), .B2(n19767), .A(n15821), .ZN(n15822) );
  AOI21_X1 U19020 ( .B1(n15823), .B2(n15933), .A(n15822), .ZN(n15824) );
  OAI21_X1 U19021 ( .B1(n16119), .B2(n16957), .A(n15824), .ZN(P2_U2998) );
  NAND2_X1 U19022 ( .A1(n15826), .A2(n15825), .ZN(n15828) );
  XOR2_X1 U19023 ( .A(n15828), .B(n15827), .Z(n16975) );
  AND2_X1 U19024 ( .A1(n16111), .A2(n16968), .ZN(n15830) );
  OR2_X1 U19025 ( .A1(n15830), .A2(n15829), .ZN(n16971) );
  INV_X1 U19026 ( .A(n19660), .ZN(n15832) );
  OAI22_X1 U19027 ( .A1(n16950), .A2(n19655), .B1(n10889), .B2(n19736), .ZN(
        n15831) );
  AOI21_X1 U19028 ( .B1(n16942), .B2(n15832), .A(n15831), .ZN(n15834) );
  NAND2_X1 U19029 ( .A1(n16946), .A2(n19657), .ZN(n15833) );
  OAI211_X1 U19030 ( .C1(n16971), .C2(n16955), .A(n15834), .B(n15833), .ZN(
        n15835) );
  INV_X1 U19031 ( .A(n15835), .ZN(n15836) );
  OAI21_X1 U19032 ( .B1(n16975), .B2(n16957), .A(n15836), .ZN(P2_U2999) );
  NAND2_X1 U19033 ( .A1(n15838), .A2(n15837), .ZN(n15840) );
  XOR2_X1 U19034 ( .A(n15840), .B(n15839), .Z(n16984) );
  AND2_X2 U19035 ( .A1(n16169), .A2(n16150), .ZN(n16145) );
  INV_X1 U19036 ( .A(n16978), .ZN(n15841) );
  AND2_X1 U19037 ( .A1(n16145), .A2(n15841), .ZN(n15855) );
  OAI21_X1 U19038 ( .B1(n15855), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16111), .ZN(n16982) );
  OAI22_X1 U19039 ( .A1(n16950), .A2(n15843), .B1(n15842), .B2(n19736), .ZN(
        n15844) );
  AOI21_X1 U19040 ( .B1(n16942), .B2(n15845), .A(n15844), .ZN(n15848) );
  INV_X1 U19041 ( .A(n19772), .ZN(n15846) );
  NAND2_X1 U19042 ( .A1(n16946), .A2(n15846), .ZN(n15847) );
  OAI211_X1 U19043 ( .C1(n16982), .C2(n16955), .A(n15848), .B(n15847), .ZN(
        n15849) );
  AOI21_X1 U19044 ( .B1(n16984), .B2(n15927), .A(n15849), .ZN(n15850) );
  INV_X1 U19045 ( .A(n15850), .ZN(P2_U3000) );
  NAND2_X1 U19046 ( .A1(n15852), .A2(n15851), .ZN(n15854) );
  XOR2_X1 U19047 ( .A(n15854), .B(n15853), .Z(n16131) );
  NAND2_X1 U19048 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16145), .ZN(
        n15864) );
  AOI21_X1 U19049 ( .B1(n10734), .B2(n15864), .A(n15855), .ZN(n16124) );
  NAND2_X1 U19050 ( .A1(n15933), .A2(n16124), .ZN(n15856) );
  NAND2_X1 U19051 ( .A1(n19903), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16123) );
  NAND2_X1 U19052 ( .A1(n15856), .A2(n16123), .ZN(n15859) );
  OAI22_X1 U19053 ( .A1(n13859), .A2(n16125), .B1(n16952), .B2(n15857), .ZN(
        n15858) );
  OAI21_X1 U19054 ( .B1(n16131), .B2(n16957), .A(n15860), .ZN(P2_U3001) );
  AOI21_X1 U19055 ( .B1(n15863), .B2(n15862), .A(n15861), .ZN(n16140) );
  OAI21_X1 U19056 ( .B1(n16145), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15864), .ZN(n16137) );
  OAI22_X1 U19057 ( .A1(n16950), .A2(n15865), .B1(n12705), .B2(n19736), .ZN(
        n15866) );
  AOI21_X1 U19058 ( .B1(n16942), .B2(n15867), .A(n15866), .ZN(n15870) );
  INV_X1 U19059 ( .A(n19777), .ZN(n15868) );
  NAND2_X1 U19060 ( .A1(n16946), .A2(n15868), .ZN(n15869) );
  OAI211_X1 U19061 ( .C1(n16137), .C2(n16955), .A(n15870), .B(n15869), .ZN(
        n15871) );
  INV_X1 U19062 ( .A(n15871), .ZN(n15872) );
  OAI21_X1 U19063 ( .B1(n16140), .B2(n16957), .A(n15872), .ZN(P2_U3002) );
  NOR2_X1 U19064 ( .A1(n15873), .A2(n16161), .ZN(n15878) );
  INV_X1 U19065 ( .A(n15874), .ZN(n15876) );
  NAND2_X1 U19066 ( .A1(n15876), .A2(n15875), .ZN(n15877) );
  XNOR2_X1 U19067 ( .A(n15878), .B(n15877), .ZN(n16997) );
  OR2_X1 U19068 ( .A1(n16997), .A2(n16957), .ZN(n15891) );
  INV_X1 U19069 ( .A(n19672), .ZN(n15882) );
  OAI22_X1 U19070 ( .A1(n16950), .A2(n15880), .B1(n19736), .B2(n15879), .ZN(
        n15881) );
  AOI21_X1 U19071 ( .B1(n16942), .B2(n15882), .A(n15881), .ZN(n15890) );
  AND2_X1 U19072 ( .A1(n16169), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16147) );
  NOR2_X1 U19073 ( .A1(n16169), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15883) );
  NOR2_X1 U19074 ( .A1(n16147), .A2(n15883), .ZN(n16994) );
  NAND2_X1 U19075 ( .A1(n16994), .A2(n15933), .ZN(n15889) );
  INV_X1 U19076 ( .A(n15884), .ZN(n15885) );
  NAND2_X1 U19077 ( .A1(n9714), .A2(n15885), .ZN(n15887) );
  AND2_X1 U19078 ( .A1(n15887), .A2(n15886), .ZN(n19780) );
  NAND2_X1 U19079 ( .A1(n16946), .A2(n19780), .ZN(n15888) );
  NAND4_X1 U19080 ( .A1(n15891), .A2(n15890), .A3(n15889), .A4(n15888), .ZN(
        P2_U3004) );
  NAND2_X1 U19081 ( .A1(n15892), .A2(n15905), .ZN(n15895) );
  XNOR2_X1 U19082 ( .A(n15893), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15894) );
  XNOR2_X1 U19083 ( .A(n15895), .B(n15894), .ZN(n17008) );
  INV_X1 U19084 ( .A(n15896), .ZN(n15897) );
  AOI21_X1 U19085 ( .B1(n15899), .B2(n15898), .A(n15897), .ZN(n17005) );
  INV_X1 U19086 ( .A(n19792), .ZN(n17004) );
  NAND2_X1 U19087 ( .A1(n17004), .A2(n16946), .ZN(n15901) );
  AOI22_X1 U19088 ( .A1(n16954), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19903), .B2(P2_REIP_REG_8__SCAN_IN), .ZN(n15900) );
  OAI211_X1 U19089 ( .C1(n15902), .C2(n16952), .A(n15901), .B(n15900), .ZN(
        n15903) );
  AOI21_X1 U19090 ( .B1(n17005), .B2(n15933), .A(n15903), .ZN(n15904) );
  OAI21_X1 U19091 ( .B1(n16957), .B2(n17008), .A(n15904), .ZN(P2_U3006) );
  NOR2_X1 U19092 ( .A1(n10682), .A2(n15906), .ZN(n15907) );
  XNOR2_X1 U19093 ( .A(n15908), .B(n15907), .ZN(n16188) );
  OAI22_X1 U19094 ( .A1(n16950), .A2(n15909), .B1(n10865), .B2(n19736), .ZN(
        n15911) );
  NOR2_X1 U19095 ( .A1(n16952), .A2(n19697), .ZN(n15910) );
  AOI211_X1 U19096 ( .C1(n16182), .C2(n16946), .A(n15911), .B(n15910), .ZN(
        n15916) );
  XNOR2_X1 U19097 ( .A(n15912), .B(n10835), .ZN(n15913) );
  XNOR2_X1 U19098 ( .A(n15914), .B(n15913), .ZN(n16185) );
  NAND2_X1 U19099 ( .A1(n16185), .A2(n15933), .ZN(n15915) );
  OAI211_X1 U19100 ( .C1(n16188), .C2(n16957), .A(n15916), .B(n15915), .ZN(
        P2_U3007) );
  OR2_X1 U19101 ( .A1(n15917), .A2(n16957), .ZN(n15925) );
  OAI22_X1 U19102 ( .A1(n16950), .A2(n15918), .B1(n14024), .B2(n19736), .ZN(
        n15919) );
  AOI21_X1 U19103 ( .B1(n16942), .B2(n19720), .A(n15919), .ZN(n15924) );
  NAND2_X1 U19104 ( .A1(n15920), .A2(n15933), .ZN(n15923) );
  NAND2_X1 U19105 ( .A1(n16946), .A2(n15921), .ZN(n15922) );
  NAND4_X1 U19106 ( .A1(n15925), .A2(n15924), .A3(n15923), .A4(n15922), .ZN(
        P2_U3009) );
  XNOR2_X1 U19107 ( .A(n15926), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17010) );
  AOI22_X1 U19108 ( .A1(n16946), .A2(n15928), .B1(n15927), .B2(n17010), .ZN(
        n15936) );
  NAND2_X1 U19109 ( .A1(n19903), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n17017) );
  OAI21_X1 U19110 ( .B1(n16954), .B2(n15929), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15935) );
  NOR2_X1 U19111 ( .A1(n15930), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15931) );
  NOR2_X1 U19112 ( .A1(n15932), .A2(n15931), .ZN(n17012) );
  NAND2_X1 U19113 ( .A1(n15933), .A2(n17012), .ZN(n15934) );
  NAND4_X1 U19114 ( .A1(n15936), .A2(n17017), .A3(n15935), .A4(n15934), .ZN(
        P2_U3014) );
  INV_X1 U19115 ( .A(n15937), .ZN(n15946) );
  NAND2_X1 U19116 ( .A1(n19909), .A2(n15938), .ZN(n15939) );
  OAI211_X1 U19117 ( .C1(n15942), .C2(n15941), .A(n15940), .B(n15939), .ZN(
        n15945) );
  NOR3_X1 U19118 ( .A1(n15971), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15943), .ZN(n15944) );
  AOI211_X1 U19119 ( .C1(n19931), .C2(n15946), .A(n15945), .B(n15944), .ZN(
        n15949) );
  NAND2_X1 U19120 ( .A1(n15947), .A2(n17013), .ZN(n15948) );
  OAI211_X1 U19121 ( .C1(n15950), .C2(n17009), .A(n15949), .B(n15948), .ZN(
        P2_U3016) );
  INV_X1 U19122 ( .A(n15951), .ZN(n15962) );
  INV_X1 U19123 ( .A(n15971), .ZN(n15952) );
  NAND2_X1 U19124 ( .A1(n15952), .A2(n15970), .ZN(n15984) );
  NAND2_X1 U19125 ( .A1(n15984), .A2(n15979), .ZN(n15974) );
  NOR2_X1 U19126 ( .A1(n15971), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15953) );
  OAI21_X1 U19127 ( .B1(n15974), .B2(n15953), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15959) );
  NOR4_X1 U19128 ( .A1(n15954), .A2(n15970), .A3(n15971), .A4(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15955) );
  AOI211_X1 U19129 ( .C1(n19909), .C2(n15957), .A(n15956), .B(n15955), .ZN(
        n15958) );
  OAI211_X1 U19130 ( .C1(n19911), .C2(n15960), .A(n15959), .B(n15958), .ZN(
        n15961) );
  AOI21_X1 U19131 ( .B1(n15962), .B2(n17013), .A(n15961), .ZN(n15963) );
  OAI21_X1 U19132 ( .B1(n15964), .B2(n17009), .A(n15963), .ZN(P2_U3017) );
  INV_X1 U19133 ( .A(n15965), .ZN(n15967) );
  AOI21_X1 U19134 ( .B1(n19909), .B2(n15967), .A(n15966), .ZN(n15968) );
  OAI21_X1 U19135 ( .B1(n15969), .B2(n19911), .A(n15968), .ZN(n15973) );
  NOR3_X1 U19136 ( .A1(n15971), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15970), .ZN(n15972) );
  AOI211_X1 U19137 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15974), .A(
        n15973), .B(n15972), .ZN(n15977) );
  NAND2_X1 U19138 ( .A1(n15975), .A2(n17013), .ZN(n15976) );
  OAI211_X1 U19139 ( .C1(n15978), .C2(n17009), .A(n15977), .B(n15976), .ZN(
        P2_U3018) );
  INV_X1 U19140 ( .A(n15979), .ZN(n15987) );
  NAND2_X1 U19141 ( .A1(n19909), .A2(n15980), .ZN(n15981) );
  OAI211_X1 U19142 ( .C1(n15983), .C2(n19911), .A(n15982), .B(n15981), .ZN(
        n15986) );
  INV_X1 U19143 ( .A(n15984), .ZN(n15985) );
  AOI211_X1 U19144 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15987), .A(
        n15986), .B(n15985), .ZN(n15991) );
  NAND3_X1 U19145 ( .A1(n15989), .A2(n17013), .A3(n15988), .ZN(n15990) );
  OAI211_X1 U19146 ( .C1(n15992), .C2(n17009), .A(n15991), .B(n15990), .ZN(
        P2_U3019) );
  NAND2_X1 U19147 ( .A1(n15993), .A2(n19920), .ZN(n16003) );
  NAND2_X1 U19148 ( .A1(n19909), .A2(n16856), .ZN(n15994) );
  OAI211_X1 U19149 ( .C1(n16858), .C2(n19911), .A(n15995), .B(n15994), .ZN(
        n16001) );
  INV_X1 U19150 ( .A(n15996), .ZN(n16010) );
  AOI211_X1 U19151 ( .C1(n15999), .C2(n15998), .A(n15997), .B(n16010), .ZN(
        n16000) );
  AOI211_X1 U19152 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n16007), .A(
        n16001), .B(n16000), .ZN(n16002) );
  OAI211_X1 U19153 ( .C1(n16004), .C2(n19926), .A(n16003), .B(n16002), .ZN(
        P2_U3020) );
  NOR2_X1 U19154 ( .A1(n19928), .A2(n16882), .ZN(n16005) );
  AOI211_X1 U19155 ( .C1(n16874), .C2(n19931), .A(n16006), .B(n16005), .ZN(
        n16009) );
  NAND2_X1 U19156 ( .A1(n16007), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16008) );
  OAI211_X1 U19157 ( .C1(n16010), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16009), .B(n16008), .ZN(n16011) );
  AOI21_X1 U19158 ( .B1(n16012), .B2(n17013), .A(n16011), .ZN(n16013) );
  OAI21_X1 U19159 ( .B1(n16014), .B2(n17009), .A(n16013), .ZN(P2_U3021) );
  NAND2_X1 U19160 ( .A1(n16015), .A2(n19920), .ZN(n16023) );
  NAND2_X1 U19161 ( .A1(n19909), .A2(n16016), .ZN(n16017) );
  OAI211_X1 U19162 ( .C1(n16888), .C2(n19911), .A(n16018), .B(n16017), .ZN(
        n16020) );
  NOR3_X1 U19163 ( .A1(n16026), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16027), .ZN(n16019) );
  AOI211_X1 U19164 ( .C1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n16021), .A(
        n16020), .B(n16019), .ZN(n16022) );
  OAI211_X1 U19165 ( .C1(n16024), .C2(n19926), .A(n16023), .B(n16022), .ZN(
        P2_U3022) );
  INV_X1 U19166 ( .A(n16025), .ZN(n16036) );
  INV_X1 U19167 ( .A(n16900), .ZN(n16034) );
  INV_X1 U19168 ( .A(n16026), .ZN(n16051) );
  OAI211_X1 U19169 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16051), .B(n16027), .ZN(
        n16033) );
  NOR2_X1 U19170 ( .A1(n16028), .A2(n16057), .ZN(n16029) );
  AOI211_X1 U19171 ( .C1(n19909), .C2(n16031), .A(n16030), .B(n16029), .ZN(
        n16032) );
  OAI211_X1 U19172 ( .C1(n16034), .C2(n19911), .A(n16033), .B(n16032), .ZN(
        n16035) );
  AOI21_X1 U19173 ( .B1(n16036), .B2(n17013), .A(n16035), .ZN(n16037) );
  OAI21_X1 U19174 ( .B1(n16038), .B2(n17009), .A(n16037), .ZN(P2_U3023) );
  OR2_X1 U19175 ( .A1(n16040), .A2(n16039), .ZN(n16042) );
  AND2_X1 U19176 ( .A1(n16042), .A2(n16041), .ZN(n16917) );
  NAND2_X1 U19177 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19903), .ZN(n16043) );
  OAI21_X1 U19178 ( .B1(n16050), .B2(n16057), .A(n16043), .ZN(n16044) );
  AOI21_X1 U19179 ( .B1(n19909), .B2(n16917), .A(n16044), .ZN(n16045) );
  OAI21_X1 U19180 ( .B1(n16906), .B2(n19911), .A(n16045), .ZN(n16049) );
  NOR3_X1 U19181 ( .A1(n16047), .A2(n16046), .A3(n19926), .ZN(n16048) );
  AOI211_X1 U19182 ( .C1(n16051), .C2(n16050), .A(n16049), .B(n16048), .ZN(
        n16052) );
  OAI21_X1 U19183 ( .B1(n16053), .B2(n17009), .A(n16052), .ZN(P2_U3024) );
  INV_X1 U19184 ( .A(n16054), .ZN(n16066) );
  INV_X1 U19185 ( .A(n16055), .ZN(n16070) );
  OR2_X1 U19186 ( .A1(n16149), .A2(n16070), .ZN(n16081) );
  NOR3_X1 U19187 ( .A1(n16081), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16056), .ZN(n16065) );
  INV_X1 U19188 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16058) );
  NOR2_X1 U19189 ( .A1(n16058), .A2(n16057), .ZN(n16059) );
  AOI211_X1 U19190 ( .C1(n16061), .C2(n19931), .A(n16060), .B(n16059), .ZN(
        n16062) );
  OAI21_X1 U19191 ( .B1(n19928), .B2(n16063), .A(n16062), .ZN(n16064) );
  AOI211_X1 U19192 ( .C1(n16066), .C2(n17013), .A(n16065), .B(n16064), .ZN(
        n16067) );
  OAI21_X1 U19193 ( .B1(n16068), .B2(n17009), .A(n16067), .ZN(P2_U3025) );
  AOI211_X1 U19194 ( .C1(n16075), .C2(n16088), .A(n16069), .B(n16081), .ZN(
        n16077) );
  AOI21_X1 U19195 ( .B1(n16497), .B2(n16070), .A(n16166), .ZN(n16086) );
  NOR2_X1 U19196 ( .A1(n19928), .A2(n16922), .ZN(n16071) );
  AOI211_X1 U19197 ( .C1(n16073), .C2(n19931), .A(n16072), .B(n16071), .ZN(
        n16074) );
  OAI21_X1 U19198 ( .B1(n16086), .B2(n16075), .A(n16074), .ZN(n16076) );
  AOI211_X1 U19199 ( .C1(n16078), .C2(n17013), .A(n16077), .B(n16076), .ZN(
        n16079) );
  OAI21_X1 U19200 ( .B1(n16080), .B2(n17009), .A(n16079), .ZN(P2_U3026) );
  INV_X1 U19201 ( .A(n16081), .ZN(n16089) );
  INV_X1 U19202 ( .A(n19627), .ZN(n16084) );
  OAI21_X1 U19203 ( .B1(n19928), .B2(n19636), .A(n16082), .ZN(n16083) );
  AOI21_X1 U19204 ( .B1(n16084), .B2(n19931), .A(n16083), .ZN(n16085) );
  OAI21_X1 U19205 ( .B1(n16086), .B2(n16088), .A(n16085), .ZN(n16087) );
  AOI21_X1 U19206 ( .B1(n16089), .B2(n16088), .A(n16087), .ZN(n16093) );
  NAND3_X1 U19207 ( .A1(n16091), .A2(n17013), .A3(n16090), .ZN(n16092) );
  OAI211_X1 U19208 ( .C1(n16094), .C2(n17009), .A(n16093), .B(n16092), .ZN(
        P2_U3027) );
  INV_X1 U19209 ( .A(n16096), .ZN(n16095) );
  NOR3_X1 U19210 ( .A1(n16149), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16095), .ZN(n16104) );
  NOR2_X1 U19211 ( .A1(n17022), .A2(n16096), .ZN(n16097) );
  OAI21_X1 U19212 ( .B1(n16097), .B2(n16166), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16101) );
  AOI21_X1 U19213 ( .B1(n19931), .B2(n16099), .A(n16098), .ZN(n16100) );
  OAI211_X1 U19214 ( .C1(n19928), .C2(n16102), .A(n16101), .B(n16100), .ZN(
        n16103) );
  AOI211_X1 U19215 ( .C1(n16105), .C2(n17013), .A(n16104), .B(n16103), .ZN(
        n16106) );
  OAI21_X1 U19216 ( .B1(n16107), .B2(n17009), .A(n16106), .ZN(P2_U3028) );
  AOI21_X1 U19217 ( .B1(n16108), .B2(n16497), .A(n16166), .ZN(n16965) );
  OAI21_X1 U19218 ( .B1(n17013), .B2(n19932), .A(n16109), .ZN(n16110) );
  OAI211_X1 U19219 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n19935), .A(
        n16965), .B(n16110), .ZN(n16499) );
  NOR2_X1 U19220 ( .A1(n19928), .A2(n19805), .ZN(n16117) );
  INV_X1 U19221 ( .A(n16111), .ZN(n16113) );
  OR2_X1 U19222 ( .A1(n16149), .A2(n16120), .ZN(n16976) );
  INV_X1 U19223 ( .A(n16977), .ZN(n16112) );
  NOR2_X1 U19224 ( .A1(n16976), .A2(n16112), .ZN(n16969) );
  AOI21_X1 U19225 ( .B1(n16113), .B2(n17013), .A(n16969), .ZN(n16492) );
  NOR2_X1 U19226 ( .A1(n16492), .A2(n16968), .ZN(n16114) );
  AOI22_X1 U19227 ( .A1(n19903), .A2(P2_REIP_REG_16__SCAN_IN), .B1(n16114), 
        .B2(n16498), .ZN(n16115) );
  OAI21_X1 U19228 ( .B1(n19911), .B2(n19767), .A(n16115), .ZN(n16116) );
  OAI21_X1 U19229 ( .B1(n16119), .B2(n17009), .A(n16118), .ZN(P2_U3030) );
  AOI21_X1 U19230 ( .B1(n16120), .B2(n16497), .A(n16166), .ZN(n16987) );
  OAI21_X1 U19231 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16976), .A(
        n16987), .ZN(n16129) );
  NOR2_X1 U19232 ( .A1(n16133), .A2(n16976), .ZN(n16121) );
  NAND2_X1 U19233 ( .A1(n10734), .A2(n16121), .ZN(n16122) );
  OAI211_X1 U19234 ( .C1(n19928), .C2(n19817), .A(n16123), .B(n16122), .ZN(
        n16128) );
  INV_X1 U19235 ( .A(n16124), .ZN(n16126) );
  OAI22_X1 U19236 ( .A1(n19926), .A2(n16126), .B1(n19911), .B2(n16125), .ZN(
        n16127) );
  AOI211_X1 U19237 ( .C1(n16129), .C2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16128), .B(n16127), .ZN(n16130) );
  OAI21_X1 U19238 ( .B1(n16131), .B2(n17009), .A(n16130), .ZN(P2_U3033) );
  NAND2_X1 U19239 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19903), .ZN(n16132) );
  OAI221_X1 U19240 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16976), 
        .C1(n16133), .C2(n16987), .A(n16132), .ZN(n16136) );
  INV_X1 U19241 ( .A(n16134), .ZN(n19820) );
  OAI22_X1 U19242 ( .A1(n19911), .A2(n19777), .B1(n19928), .B2(n19820), .ZN(
        n16135) );
  NOR2_X1 U19243 ( .A1(n16136), .A2(n16135), .ZN(n16139) );
  OR2_X1 U19244 ( .A1(n16137), .A2(n19926), .ZN(n16138) );
  OAI211_X1 U19245 ( .C1(n16140), .C2(n17009), .A(n16139), .B(n16138), .ZN(
        P2_U3034) );
  NAND2_X1 U19246 ( .A1(n16142), .A2(n16141), .ZN(n16143) );
  XNOR2_X1 U19247 ( .A(n16144), .B(n16143), .ZN(n16936) );
  INV_X1 U19248 ( .A(n16145), .ZN(n16146) );
  OAI21_X1 U19249 ( .B1(n16147), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16146), .ZN(n16935) );
  INV_X1 U19250 ( .A(n16166), .ZN(n16148) );
  OAI21_X1 U19251 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17022), .A(
        n16148), .ZN(n16993) );
  NOR2_X1 U19252 ( .A1(n12702), .A2(n19736), .ZN(n16153) );
  INV_X1 U19253 ( .A(n16149), .ZN(n16175) );
  NAND2_X1 U19254 ( .A1(n16175), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16990) );
  AOI211_X1 U19255 ( .C1(n16151), .C2(n10736), .A(n16150), .B(n16990), .ZN(
        n16152) );
  AOI211_X1 U19256 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16993), .A(
        n16153), .B(n16152), .ZN(n16156) );
  AOI22_X1 U19257 ( .A1(n19931), .A2(n16938), .B1(n19909), .B2(n16154), .ZN(
        n16155) );
  OAI211_X1 U19258 ( .C1(n16935), .C2(n19926), .A(n16156), .B(n16155), .ZN(
        n16157) );
  INV_X1 U19259 ( .A(n16157), .ZN(n16158) );
  OAI21_X1 U19260 ( .B1(n16936), .B2(n17009), .A(n16158), .ZN(P2_U3035) );
  OR2_X1 U19261 ( .A1(n16161), .A2(n16160), .ZN(n16162) );
  XNOR2_X1 U19262 ( .A(n16159), .B(n16162), .ZN(n16943) );
  OAI21_X1 U19263 ( .B1(n16164), .B2(n16163), .A(n16989), .ZN(n19827) );
  NAND2_X1 U19264 ( .A1(n19931), .A2(n19691), .ZN(n16168) );
  NOR2_X1 U19265 ( .A1(n10846), .A2(n19736), .ZN(n16165) );
  AOI21_X1 U19266 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16166), .A(
        n16165), .ZN(n16167) );
  OAI211_X1 U19267 ( .C1(n19928), .C2(n19827), .A(n16168), .B(n16167), .ZN(
        n16173) );
  INV_X1 U19268 ( .A(n16169), .ZN(n16170) );
  OAI21_X1 U19269 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16171), .A(
        n16170), .ZN(n16944) );
  NOR2_X1 U19270 ( .A1(n16944), .A2(n19926), .ZN(n16172) );
  AOI211_X1 U19271 ( .C1(n16175), .C2(n16174), .A(n16173), .B(n16172), .ZN(
        n16176) );
  OAI21_X1 U19272 ( .B1(n17009), .B2(n16943), .A(n16176), .ZN(P2_U3037) );
  OAI21_X1 U19273 ( .B1(n16179), .B2(n16178), .A(n16177), .ZN(n19832) );
  NOR2_X1 U19274 ( .A1(n10865), .A2(n19736), .ZN(n16181) );
  NOR2_X1 U19275 ( .A1(n10835), .A2(n17001), .ZN(n16180) );
  AOI211_X1 U19276 ( .C1(n19931), .C2(n16182), .A(n16181), .B(n16180), .ZN(
        n16183) );
  OAI21_X1 U19277 ( .B1(n19832), .B2(n19928), .A(n16183), .ZN(n16184) );
  AOI21_X1 U19278 ( .B1(n16998), .B2(n10835), .A(n16184), .ZN(n16187) );
  NAND2_X1 U19279 ( .A1(n16185), .A2(n17013), .ZN(n16186) );
  OAI211_X1 U19280 ( .C1(n16188), .C2(n17009), .A(n16187), .B(n16186), .ZN(
        P2_U3039) );
  OR2_X1 U19281 ( .A1(n16191), .A2(n16190), .ZN(n16192) );
  NAND2_X1 U19282 ( .A1(n16189), .A2(n16192), .ZN(n16958) );
  XNOR2_X1 U19283 ( .A(n16194), .B(n16193), .ZN(n19835) );
  NAND2_X1 U19284 ( .A1(n19903), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n16951) );
  NAND2_X1 U19285 ( .A1(n19931), .A2(n16195), .ZN(n16196) );
  OAI211_X1 U19286 ( .C1(n19835), .C2(n19928), .A(n16951), .B(n16196), .ZN(
        n16198) );
  AOI211_X1 U19287 ( .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16199), .A(
        n16198), .B(n16197), .ZN(n16203) );
  OAI21_X1 U19288 ( .B1(n16201), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16200), .ZN(n16956) );
  OR2_X1 U19289 ( .A1(n16956), .A2(n19926), .ZN(n16202) );
  OAI211_X1 U19290 ( .C1(n16958), .C2(n17009), .A(n16203), .B(n16202), .ZN(
        P2_U3040) );
  OAI22_X1 U19291 ( .A1(n19926), .A2(n16205), .B1(n17009), .B2(n16204), .ZN(
        n16206) );
  AOI211_X1 U19292 ( .C1(n17011), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n16207), .B(n16206), .ZN(n16211) );
  OAI211_X1 U19293 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n16497), .B(n16208), .ZN(n16210) );
  AOI22_X1 U19294 ( .A1(n10533), .A2(n19931), .B1(n19909), .B2(n20603), .ZN(
        n16209) );
  NAND3_X1 U19295 ( .A1(n16211), .A2(n16210), .A3(n16209), .ZN(P2_U3045) );
  INV_X1 U19296 ( .A(n20569), .ZN(n17083) );
  NOR2_X1 U19297 ( .A1(n16212), .A2(n14486), .ZN(n16213) );
  AOI22_X1 U19298 ( .A1(n16214), .A2(n16213), .B1(n17033), .B2(n10201), .ZN(
        n16215) );
  OAI21_X1 U19299 ( .B1(n16217), .B2(n16216), .A(n16215), .ZN(n17037) );
  AOI22_X1 U19300 ( .A1(n20599), .A2(n17083), .B1(n20579), .B2(n17037), .ZN(
        n16218) );
  OAI21_X1 U19301 ( .B1(n16220), .B2(n16219), .A(n16218), .ZN(n16221) );
  MUX2_X1 U19302 ( .A(n16221), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n20571), .Z(P2_U3600) );
  NOR3_X1 U19303 ( .A1(n20481), .A2(n19995), .A3(n20578), .ZN(n16224) );
  AND2_X1 U19304 ( .A1(n20585), .A2(n21109), .ZN(n20580) );
  NOR2_X1 U19305 ( .A1(n16224), .A2(n20580), .ZN(n16227) );
  OR2_X1 U19306 ( .A1(n20021), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19975) );
  NOR2_X1 U19307 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19975), .ZN(
        n19963) );
  INV_X1 U19308 ( .A(n19963), .ZN(n16225) );
  AND2_X1 U19309 ( .A1(n20423), .A2(n16225), .ZN(n16230) );
  OAI21_X1 U19310 ( .B1(n16228), .B2(n19963), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16226) );
  INV_X1 U19311 ( .A(n16227), .ZN(n16231) );
  AOI211_X1 U19312 ( .C1(n16228), .C2(n21204), .A(n19963), .B(n20585), .ZN(
        n16229) );
  AOI22_X1 U19313 ( .A1(n20440), .A2(n19995), .B1(n20439), .B2(n19963), .ZN(
        n16233) );
  NAND2_X1 U19314 ( .A1(n20441), .A2(n20481), .ZN(n16232) );
  OAI211_X1 U19315 ( .C1(n19971), .C2(n16234), .A(n16233), .B(n16232), .ZN(
        n16235) );
  AOI21_X1 U19316 ( .B1(n13863), .B2(n19967), .A(n16235), .ZN(n16236) );
  INV_X1 U19317 ( .A(n16236), .ZN(P2_U3049) );
  NOR2_X2 U19318 ( .A1(n19831), .A2(n20395), .ZN(n20478) );
  AOI22_X1 U19319 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19965), .ZN(n20351) );
  AND2_X1 U19320 ( .A1(n16237), .A2(n19951), .ZN(n20476) );
  AOI22_X1 U19321 ( .A1(n20480), .A2(n19995), .B1(n19963), .B2(n20476), .ZN(
        n16239) );
  AOI22_X1 U19322 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19965), .ZN(n20388) );
  NAND2_X1 U19323 ( .A1(n20482), .A2(n20481), .ZN(n16238) );
  OAI211_X1 U19324 ( .C1(n19971), .C2(n16240), .A(n16239), .B(n16238), .ZN(
        n16241) );
  AOI21_X1 U19325 ( .B1(n20478), .B2(n19967), .A(n16241), .ZN(n16242) );
  INV_X1 U19326 ( .A(n16242), .ZN(P2_U3055) );
  INV_X1 U19327 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16244) );
  OAI33_X1 U19328 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16245), .A3(n18087), 
        .B1(n16244), .B2(n17942), .B3(n16243), .ZN(P3_U2672) );
  AOI22_X1 U19329 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16256) );
  AOI22_X1 U19330 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n17900), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16255) );
  INV_X1 U19331 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17921) );
  AOI22_X1 U19332 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17821), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16246) );
  OAI21_X1 U19333 ( .B1(n16247), .B2(n17921), .A(n16246), .ZN(n16253) );
  AOI22_X1 U19334 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16251) );
  AOI22_X1 U19335 ( .A1(n16346), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16250) );
  AOI22_X1 U19336 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16249) );
  AOI22_X1 U19337 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16248) );
  NAND4_X1 U19338 ( .A1(n16251), .A2(n16250), .A3(n16249), .A4(n16248), .ZN(
        n16252) );
  AOI211_X1 U19339 ( .C1(n17893), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n16253), .B(n16252), .ZN(n16254) );
  NAND3_X1 U19340 ( .A1(n16256), .A2(n16255), .A3(n16254), .ZN(n18039) );
  INV_X1 U19341 ( .A(n18039), .ZN(n16258) );
  AOI21_X1 U19342 ( .B1(n17935), .B2(n17857), .A(n17842), .ZN(n17845) );
  NOR2_X1 U19343 ( .A1(n17942), .A2(n17829), .ZN(n17830) );
  OAI21_X1 U19344 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17845), .A(n17830), .ZN(
        n16257) );
  OAI21_X1 U19345 ( .B1(n16258), .B2(n17935), .A(n16257), .ZN(P3_U2690) );
  NAND2_X1 U19346 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19093) );
  AOI221_X1 U19347 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19093), .C1(n16260), 
        .C2(n19093), .A(n16259), .ZN(n18914) );
  NOR2_X1 U19348 ( .A1(n16261), .A2(n19387), .ZN(n16262) );
  OAI21_X1 U19349 ( .B1(n16262), .B2(n19265), .A(n18915), .ZN(n18912) );
  AOI22_X1 U19350 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18914), .B1(
        n18912), .B2(n19403), .ZN(P3_U2865) );
  NAND2_X1 U19351 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19568) );
  XNOR2_X1 U19352 ( .A(n16264), .B(n16263), .ZN(n16266) );
  NOR2_X1 U19353 ( .A1(n19575), .A2(n17271), .ZN(n16559) );
  NAND3_X1 U19354 ( .A1(n18930), .A2(n18938), .A3(n18945), .ZN(n16272) );
  INV_X1 U19355 ( .A(n18141), .ZN(n16285) );
  NOR2_X1 U19356 ( .A1(n18954), .A2(n18102), .ZN(n16275) );
  NAND3_X1 U19357 ( .A1(n16275), .A2(n16268), .A3(n18926), .ZN(n16269) );
  NOR2_X1 U19358 ( .A1(n18942), .A2(n18945), .ZN(n16277) );
  NAND4_X1 U19359 ( .A1(n18934), .A2(n18938), .A3(n16275), .A4(n16277), .ZN(
        n16283) );
  NAND2_X1 U19360 ( .A1(n18923), .A2(n19574), .ZN(n16432) );
  INV_X1 U19361 ( .A(n16439), .ZN(n16284) );
  NAND2_X1 U19362 ( .A1(n16270), .A2(n18945), .ZN(n16563) );
  NOR2_X1 U19363 ( .A1(n18954), .A2(n19381), .ZN(n16561) );
  NAND2_X1 U19364 ( .A1(n18926), .A2(n18102), .ZN(n16431) );
  AOI21_X1 U19365 ( .B1(n16271), .B2(n16272), .A(n16294), .ZN(n16282) );
  INV_X1 U19366 ( .A(n16271), .ZN(n16424) );
  NAND2_X1 U19367 ( .A1(n16424), .A2(n16417), .ZN(n16425) );
  AOI21_X1 U19368 ( .B1(n16272), .B2(n16425), .A(n18102), .ZN(n16281) );
  OAI22_X1 U19369 ( .A1(n16275), .A2(n16274), .B1(n16273), .B2(n16563), .ZN(
        n16280) );
  NOR2_X1 U19370 ( .A1(n18954), .A2(n16277), .ZN(n16278) );
  NAND2_X1 U19371 ( .A1(n16432), .A2(n18930), .ZN(n16287) );
  INV_X1 U19372 ( .A(n16287), .ZN(n16276) );
  OAI22_X1 U19373 ( .A1(n18938), .A2(n16278), .B1(n16277), .B2(n16276), .ZN(
        n16279) );
  NOR3_X1 U19374 ( .A1(n16281), .A2(n16280), .A3(n16279), .ZN(n16291) );
  OAI21_X1 U19375 ( .B1(n18934), .B2(n16282), .A(n16291), .ZN(n16437) );
  NOR2_X2 U19376 ( .A1(n16283), .A2(n16437), .ZN(n16440) );
  INV_X1 U19377 ( .A(n16558), .ZN(n16286) );
  NAND2_X2 U19378 ( .A1(n19584), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19509) );
  OAI211_X1 U19379 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19448), .B(n19509), .ZN(n19440) );
  INV_X1 U19380 ( .A(n19440), .ZN(n19573) );
  NAND2_X1 U19381 ( .A1(n16286), .A2(n18100), .ZN(n16297) );
  NOR2_X1 U19382 ( .A1(n16434), .A2(n16287), .ZN(n16289) );
  OAI211_X1 U19383 ( .C1(n18938), .C2(n19381), .A(n16289), .B(n16288), .ZN(
        n16418) );
  INV_X1 U19384 ( .A(n16418), .ZN(n16292) );
  AOI21_X1 U19385 ( .B1(n16292), .B2(n16291), .A(n16290), .ZN(n16293) );
  INV_X1 U19386 ( .A(n16430), .ZN(n16295) );
  AOI211_X1 U19387 ( .C1(n16559), .C2(n16297), .A(n16296), .B(n16295), .ZN(
        n19398) );
  INV_X1 U19388 ( .A(n19398), .ZN(n19379) );
  NOR2_X1 U19389 ( .A1(n17275), .A2(n19523), .ZN(n16298) );
  NOR2_X1 U19390 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19524), .ZN(n18922) );
  INV_X1 U19391 ( .A(n19555), .ZN(n19552) );
  INV_X1 U19392 ( .A(n19526), .ZN(n19588) );
  INV_X1 U19393 ( .A(n16299), .ZN(n16300) );
  NOR2_X1 U19394 ( .A1(n16300), .A2(n19357), .ZN(n19366) );
  NAND3_X1 U19395 ( .A1(n19552), .A2(n19588), .A3(n19366), .ZN(n16301) );
  OAI21_X1 U19396 ( .B1(n19552), .B2(n17605), .A(n16301), .ZN(P3_U3284) );
  INV_X1 U19397 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U19398 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17903), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16312) );
  AOI22_X1 U19399 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17862), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16311) );
  AOI22_X1 U19400 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16302) );
  OAI21_X1 U19401 ( .B1(n16303), .B2(n10197), .A(n16302), .ZN(n16309) );
  AOI22_X1 U19402 ( .A1(n17883), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16307) );
  AOI22_X1 U19403 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16306) );
  AOI22_X1 U19404 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16305) );
  AOI22_X1 U19405 ( .A1(n17894), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16304) );
  NAND4_X1 U19406 ( .A1(n16307), .A2(n16306), .A3(n16305), .A4(n16304), .ZN(
        n16308) );
  AOI211_X1 U19407 ( .C1(n17900), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n16309), .B(n16308), .ZN(n16310) );
  NAND3_X1 U19408 ( .A1(n16312), .A2(n16311), .A3(n16310), .ZN(n17156) );
  AOI22_X1 U19409 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16316) );
  AOI22_X1 U19410 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16315) );
  AOI22_X1 U19411 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16314) );
  AOI22_X1 U19412 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n17894), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16313) );
  NAND4_X1 U19413 ( .A1(n16316), .A2(n16315), .A3(n16314), .A4(n16313), .ZN(
        n16322) );
  AOI22_X1 U19414 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16320) );
  AOI22_X1 U19415 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16319) );
  AOI22_X1 U19416 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17903), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16318) );
  AOI22_X1 U19417 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16317) );
  NAND4_X1 U19418 ( .A1(n16320), .A2(n16319), .A3(n16318), .A4(n16317), .ZN(
        n16321) );
  AOI22_X1 U19419 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16326) );
  AOI22_X1 U19420 ( .A1(n16346), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16325) );
  AOI22_X1 U19421 ( .A1(n17883), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16324) );
  AOI22_X1 U19422 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n9595), .B1(
        n17816), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16323) );
  NAND4_X1 U19423 ( .A1(n16326), .A2(n16325), .A3(n16324), .A4(n16323), .ZN(
        n16332) );
  AOI22_X1 U19424 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n17901), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16330) );
  AOI22_X1 U19425 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17862), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16329) );
  AOI22_X1 U19426 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16328) );
  AOI22_X1 U19427 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16327) );
  NAND4_X1 U19428 ( .A1(n16330), .A2(n16329), .A3(n16328), .A4(n16327), .ZN(
        n16331) );
  AOI22_X1 U19429 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16343) );
  AOI22_X1 U19430 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16342) );
  AOI22_X1 U19431 ( .A1(n16386), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14168), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16333) );
  OAI21_X1 U19432 ( .B1(n17790), .B2(n17937), .A(n16333), .ZN(n16340) );
  AOI22_X1 U19433 ( .A1(n17883), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16338) );
  AOI22_X1 U19434 ( .A1(n16387), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16334), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16337) );
  AOI22_X1 U19435 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n16346), .B1(
        n16368), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16336) );
  AOI22_X1 U19436 ( .A1(n14170), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16335) );
  NAND4_X1 U19437 ( .A1(n16338), .A2(n16337), .A3(n16336), .A4(n16335), .ZN(
        n16339) );
  AOI22_X1 U19438 ( .A1(n16387), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16355) );
  AOI22_X1 U19439 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16354) );
  AOI22_X1 U19440 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16344) );
  OAI21_X1 U19441 ( .B1(n21216), .B2(n16345), .A(n16344), .ZN(n16352) );
  AOI22_X1 U19442 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n16386), .B1(
        n17816), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16350) );
  AOI22_X1 U19443 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16349) );
  AOI22_X1 U19444 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16346), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16348) );
  AOI22_X1 U19445 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16347) );
  NAND4_X1 U19446 ( .A1(n16350), .A2(n16349), .A3(n16348), .A4(n16347), .ZN(
        n16351) );
  AOI211_X1 U19447 ( .C1(n14170), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n16352), .B(n16351), .ZN(n16353) );
  NAND3_X1 U19448 ( .A1(n16355), .A2(n16354), .A3(n16353), .ZN(n16445) );
  AOI22_X1 U19449 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16365) );
  AOI22_X1 U19450 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17821), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16364) );
  AOI22_X1 U19451 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16356) );
  OAI21_X1 U19452 ( .B1(n17790), .B2(n17925), .A(n16356), .ZN(n16362) );
  AOI22_X1 U19453 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16360) );
  AOI22_X1 U19454 ( .A1(n17883), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16359) );
  AOI22_X1 U19455 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16358) );
  AOI22_X1 U19456 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16357) );
  NAND4_X1 U19457 ( .A1(n16360), .A2(n16359), .A3(n16358), .A4(n16357), .ZN(
        n16361) );
  AOI211_X1 U19458 ( .C1(n17903), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n16362), .B(n16361), .ZN(n16363) );
  NAND3_X1 U19459 ( .A1(n16365), .A2(n16364), .A3(n16363), .ZN(n18080) );
  AOI22_X1 U19460 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16377) );
  AOI22_X1 U19461 ( .A1(n16346), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16376) );
  AOI22_X1 U19462 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16366) );
  OAI21_X1 U19463 ( .B1(n21139), .B2(n16367), .A(n16366), .ZN(n16374) );
  AOI22_X1 U19464 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16372) );
  AOI22_X1 U19465 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16371) );
  AOI22_X1 U19466 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16370) );
  AOI22_X1 U19467 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n16368), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16369) );
  NAND4_X1 U19468 ( .A1(n16372), .A2(n16371), .A3(n16370), .A4(n16369), .ZN(
        n16373) );
  AOI211_X1 U19469 ( .C1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .C2(n17894), .A(
        n16374), .B(n16373), .ZN(n16375) );
  NAND3_X1 U19470 ( .A1(n16377), .A2(n16376), .A3(n16375), .ZN(n18072) );
  NOR2_X4 U19471 ( .A1(n18068), .A2(n17158), .ZN(n18496) );
  INV_X1 U19472 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18217) );
  NAND2_X1 U19473 ( .A1(n18404), .A2(n18217), .ZN(n17155) );
  INV_X1 U19474 ( .A(n17155), .ZN(n16544) );
  INV_X1 U19475 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18612) );
  NOR2_X1 U19476 ( .A1(n18496), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18355) );
  INV_X1 U19477 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18683) );
  NAND2_X1 U19478 ( .A1(n18355), .A2(n18683), .ZN(n16378) );
  NOR2_X1 U19479 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16378), .ZN(
        n18316) );
  INV_X1 U19480 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18318) );
  NAND2_X1 U19481 ( .A1(n18316), .A2(n18318), .ZN(n18292) );
  AOI21_X1 U19482 ( .B1(n18068), .B2(n17158), .A(n18496), .ZN(n16404) );
  XOR2_X1 U19483 ( .A(n16379), .B(n18072), .Z(n16402) );
  INV_X1 U19484 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18850) );
  XOR2_X1 U19485 ( .A(n16380), .B(n18076), .Z(n18529) );
  INV_X1 U19486 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18856) );
  INV_X1 U19487 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16395) );
  NAND2_X1 U19488 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n16381), .ZN(
        n16394) );
  INV_X1 U19489 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19535) );
  AOI22_X1 U19490 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n16346), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16385) );
  AOI22_X1 U19491 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16384) );
  AOI22_X1 U19492 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16383) );
  AOI22_X1 U19493 ( .A1(n14170), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16382) );
  NAND4_X1 U19494 ( .A1(n16385), .A2(n16384), .A3(n16383), .A4(n16382), .ZN(
        n16393) );
  AOI22_X1 U19495 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16391) );
  AOI22_X1 U19496 ( .A1(n17883), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16390) );
  AOI22_X1 U19497 ( .A1(n16387), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16386), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16389) );
  AOI22_X1 U19498 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16388) );
  NAND4_X1 U19499 ( .A1(n16391), .A2(n16390), .A3(n16389), .A4(n16388), .ZN(
        n16392) );
  INV_X1 U19500 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19551) );
  NOR2_X1 U19501 ( .A1(n16564), .A2(n19551), .ZN(n18584) );
  NAND2_X1 U19502 ( .A1(n18584), .A2(n18578), .ZN(n18577) );
  OAI21_X1 U19503 ( .B1(n19535), .B2(n16455), .A(n18577), .ZN(n18565) );
  XNOR2_X1 U19504 ( .A(n16395), .B(n16397), .ZN(n18554) );
  XOR2_X1 U19505 ( .A(n16396), .B(n18084), .Z(n18555) );
  NAND2_X1 U19506 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16397), .ZN(
        n16398) );
  XNOR2_X1 U19507 ( .A(n18856), .B(n16400), .ZN(n18539) );
  XOR2_X1 U19508 ( .A(n16399), .B(n18080), .Z(n18538) );
  NAND2_X1 U19509 ( .A1(n18539), .A2(n18538), .ZN(n18537) );
  NAND2_X1 U19510 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n16400), .ZN(
        n16401) );
  XOR2_X1 U19511 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16402), .Z(
        n18515) );
  NAND2_X1 U19512 ( .A1(n16404), .A2(n16403), .ZN(n16405) );
  INV_X1 U19513 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18769) );
  INV_X1 U19514 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18808) );
  INV_X1 U19515 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18465) );
  NOR2_X1 U19516 ( .A1(n18808), .A2(n18465), .ZN(n18748) );
  NAND2_X1 U19517 ( .A1(n18748), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18770) );
  NAND3_X1 U19518 ( .A1(n18751), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18395) );
  NOR2_X1 U19519 ( .A1(n18769), .A2(n18395), .ZN(n18719) );
  INV_X1 U19520 ( .A(n18719), .ZN(n18708) );
  INV_X1 U19521 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18730) );
  NOR2_X1 U19522 ( .A1(n18708), .A2(n18730), .ZN(n16473) );
  INV_X1 U19523 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18632) );
  INV_X1 U19524 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18711) );
  INV_X1 U19525 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18700) );
  NOR2_X1 U19526 ( .A1(n18711), .A2(n18700), .ZN(n18348) );
  NAND2_X1 U19527 ( .A1(n18348), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18322) );
  INV_X1 U19528 ( .A(n18322), .ZN(n18661) );
  INV_X1 U19529 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18326) );
  NOR2_X1 U19530 ( .A1(n18683), .A2(n18326), .ZN(n18664) );
  NAND2_X1 U19531 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18664), .ZN(
        n18652) );
  INV_X1 U19532 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18650) );
  NOR2_X1 U19533 ( .A1(n18652), .A2(n18650), .ZN(n18631) );
  NAND2_X1 U19534 ( .A1(n18661), .A2(n18631), .ZN(n18638) );
  NOR2_X1 U19535 ( .A1(n18632), .A2(n18638), .ZN(n18272) );
  NOR4_X1 U19536 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16408) );
  AOI21_X1 U19537 ( .B1(n16408), .B2(n16407), .A(n18496), .ZN(n18373) );
  NAND2_X1 U19538 ( .A1(n18348), .A2(n18293), .ZN(n18314) );
  NAND2_X1 U19539 ( .A1(n18324), .A2(n18314), .ZN(n18315) );
  NAND3_X1 U19540 ( .A1(n18631), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18315), .ZN(n18276) );
  NAND2_X1 U19541 ( .A1(n18404), .A2(n18260), .ZN(n16411) );
  OAI221_X1 U19542 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18404), 
        .C1(n18612), .C2(n16412), .A(n16411), .ZN(n18241) );
  NOR2_X1 U19543 ( .A1(n16412), .A2(n18404), .ZN(n18259) );
  NAND2_X1 U19544 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18598) );
  NAND2_X1 U19545 ( .A1(n18496), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17154) );
  AOI21_X1 U19546 ( .B1(n16544), .B2(n18227), .A(n16543), .ZN(n16415) );
  XNOR2_X1 U19547 ( .A(n17128), .B(n16415), .ZN(n17141) );
  NOR2_X1 U19548 ( .A1(n18926), .A2(n16416), .ZN(n16423) );
  NAND2_X1 U19549 ( .A1(n16423), .A2(n16417), .ZN(n16419) );
  INV_X1 U19550 ( .A(n16419), .ZN(n16428) );
  INV_X1 U19551 ( .A(n17271), .ZN(n19356) );
  OAI21_X1 U19552 ( .B1(n16421), .B2(n16420), .A(n19356), .ZN(n19363) );
  INV_X1 U19553 ( .A(n19363), .ZN(n17090) );
  OAI21_X1 U19554 ( .B1(n18930), .B2(n19574), .A(n19440), .ZN(n16422) );
  OAI21_X1 U19555 ( .B1(n16423), .B2(n16422), .A(n19568), .ZN(n17270) );
  NOR3_X1 U19556 ( .A1(n16424), .A2(n17271), .A3(n17270), .ZN(n16427) );
  AOI21_X1 U19557 ( .B1(n18938), .B2(n16425), .A(n17089), .ZN(n16426) );
  AOI211_X1 U19558 ( .C1(n16428), .C2(n17090), .A(n16427), .B(n16426), .ZN(
        n16429) );
  NAND3_X1 U19559 ( .A1(n19364), .A2(n18898), .A3(n17156), .ZN(n18799) );
  OR3_X2 U19560 ( .A1(n19526), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18890) );
  INV_X2 U19561 ( .A(n18890), .ZN(n18902) );
  NAND2_X1 U19562 ( .A1(n16432), .A2(n16431), .ZN(n19589) );
  INV_X1 U19563 ( .A(n16434), .ZN(n16435) );
  NOR3_X1 U19564 ( .A1(n16436), .A2(n16435), .A3(n18926), .ZN(n16438) );
  NOR2_X1 U19565 ( .A1(n16438), .A2(n16437), .ZN(n19367) );
  NAND2_X1 U19566 ( .A1(n19397), .A2(n19382), .ZN(n18707) );
  INV_X1 U19567 ( .A(n18707), .ZN(n18794) );
  NAND2_X1 U19568 ( .A1(n18272), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18614) );
  NOR2_X1 U19569 ( .A1(n18614), .A2(n18598), .ZN(n17114) );
  INV_X1 U19570 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18819) );
  INV_X1 U19571 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18832) );
  INV_X1 U19572 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18831) );
  NOR3_X1 U19573 ( .A1(n18819), .A2(n18832), .A3(n18831), .ZN(n16442) );
  INV_X1 U19574 ( .A(n16442), .ZN(n18692) );
  NAND3_X1 U19575 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16441) );
  INV_X1 U19576 ( .A(n16441), .ZN(n18810) );
  NAND3_X1 U19577 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18810), .ZN(n18811) );
  NOR2_X1 U19578 ( .A1(n18692), .A2(n18811), .ZN(n18792) );
  INV_X1 U19579 ( .A(n18792), .ZN(n18749) );
  NOR2_X1 U19580 ( .A1(n18693), .A2(n18749), .ZN(n18599) );
  INV_X1 U19581 ( .A(n18599), .ZN(n18647) );
  NOR2_X1 U19582 ( .A1(n19551), .A2(n18647), .ZN(n18704) );
  NAND3_X1 U19583 ( .A1(n17114), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n18704), .ZN(n16444) );
  AOI21_X1 U19584 ( .B1(n17114), .B2(n18599), .A(n19382), .ZN(n16443) );
  AOI21_X1 U19585 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18880) );
  NOR2_X1 U19586 ( .A1(n18880), .A2(n16441), .ZN(n18813) );
  NAND2_X1 U19587 ( .A1(n18813), .A2(n16442), .ZN(n18705) );
  NOR2_X1 U19588 ( .A1(n18693), .A2(n18705), .ZN(n18685) );
  AOI21_X1 U19589 ( .B1(n17114), .B2(n18685), .A(n19397), .ZN(n18597) );
  AOI211_X1 U19590 ( .C1(n19380), .C2(n16444), .A(n16443), .B(n18597), .ZN(
        n16546) );
  NAND2_X1 U19591 ( .A1(n18890), .A2(n18887), .ZN(n18815) );
  OAI211_X1 U19592 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n18794), .A(
        n16546), .B(n18815), .ZN(n17161) );
  AOI21_X1 U19593 ( .B1(n18814), .B2(n18217), .A(n17161), .ZN(n16472) );
  NAND2_X1 U19594 ( .A1(n18753), .A2(n18898), .ZN(n18896) );
  NAND2_X1 U19595 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17126) );
  NOR2_X1 U19596 ( .A1(n17126), .A2(n17128), .ZN(n17108) );
  INV_X1 U19597 ( .A(n17114), .ZN(n17153) );
  NOR2_X1 U19598 ( .A1(n18099), .A2(n16564), .ZN(n16456) );
  NOR2_X1 U19599 ( .A1(n16456), .A2(n16445), .ZN(n16451) );
  NOR2_X1 U19600 ( .A1(n18084), .A2(n16451), .ZN(n16449) );
  NAND2_X1 U19601 ( .A1(n16449), .A2(n18080), .ZN(n16448) );
  NOR2_X1 U19602 ( .A1(n18076), .A2(n16448), .ZN(n16447) );
  NAND2_X1 U19603 ( .A1(n16447), .A2(n18072), .ZN(n16446) );
  NOR2_X1 U19604 ( .A1(n18068), .A2(n16446), .ZN(n16470) );
  XNOR2_X1 U19605 ( .A(n17156), .B(n16446), .ZN(n18507) );
  XOR2_X1 U19606 ( .A(n18072), .B(n16447), .Z(n16463) );
  XOR2_X1 U19607 ( .A(n18076), .B(n16448), .Z(n16461) );
  NAND2_X1 U19608 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16461), .ZN(
        n16462) );
  XOR2_X1 U19609 ( .A(n18080), .B(n16449), .Z(n18543) );
  XOR2_X1 U19610 ( .A(n16451), .B(n18084), .Z(n16450) );
  NAND2_X1 U19611 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16450), .ZN(
        n16459) );
  XOR2_X1 U19612 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n16450), .Z(
        n18558) );
  INV_X1 U19613 ( .A(n16564), .ZN(n16453) );
  AOI21_X1 U19614 ( .B1(n16453), .B2(n16452), .A(n16451), .ZN(n16454) );
  OR2_X1 U19615 ( .A1(n9990), .A2(n16454), .ZN(n16458) );
  XOR2_X1 U19616 ( .A(n9990), .B(n16454), .Z(n18569) );
  NOR2_X1 U19617 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16455), .ZN(
        n16457) );
  NAND2_X1 U19618 ( .A1(n16564), .A2(n19551), .ZN(n18585) );
  NOR2_X1 U19619 ( .A1(n18578), .A2(n18585), .ZN(n18576) );
  NOR3_X1 U19620 ( .A1(n16457), .A2(n16456), .A3(n18576), .ZN(n18568) );
  NAND2_X1 U19621 ( .A1(n18569), .A2(n18568), .ZN(n18567) );
  NAND2_X1 U19622 ( .A1(n16458), .A2(n18567), .ZN(n18557) );
  NAND2_X1 U19623 ( .A1(n18558), .A2(n18557), .ZN(n18556) );
  NAND2_X1 U19624 ( .A1(n16459), .A2(n18556), .ZN(n18542) );
  NAND2_X1 U19625 ( .A1(n18543), .A2(n18542), .ZN(n16460) );
  NOR2_X1 U19626 ( .A1(n18543), .A2(n18542), .ZN(n18541) );
  AOI21_X1 U19627 ( .B1(n18856), .B2(n16460), .A(n18541), .ZN(n18526) );
  XOR2_X1 U19628 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n16461), .Z(
        n18525) );
  NAND2_X1 U19629 ( .A1(n18526), .A2(n18525), .ZN(n18524) );
  NAND2_X1 U19630 ( .A1(n16462), .A2(n18524), .ZN(n16464) );
  NAND2_X1 U19631 ( .A1(n16463), .A2(n16464), .ZN(n16465) );
  XOR2_X1 U19632 ( .A(n16464), .B(n16463), .Z(n18513) );
  NAND2_X1 U19633 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18513), .ZN(
        n18512) );
  NAND2_X1 U19634 ( .A1(n16470), .A2(n16466), .ZN(n16471) );
  INV_X1 U19635 ( .A(n16466), .ZN(n16469) );
  NAND2_X1 U19636 ( .A1(n18507), .A2(n18506), .ZN(n16468) );
  NAND2_X1 U19637 ( .A1(n16470), .A2(n16469), .ZN(n16467) );
  OAI211_X1 U19638 ( .C1(n16470), .C2(n16469), .A(n16468), .B(n16467), .ZN(
        n18484) );
  NAND2_X1 U19639 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18484), .ZN(
        n18483) );
  NOR2_X1 U19640 ( .A1(n17153), .A2(n18717), .ZN(n18594) );
  NAND2_X1 U19641 ( .A1(n17108), .A2(n18594), .ZN(n17119) );
  NAND2_X1 U19642 ( .A1(n18068), .A2(n19364), .ZN(n18755) );
  NOR2_X1 U19643 ( .A1(n18887), .A2(n18755), .ZN(n18823) );
  NAND2_X1 U19644 ( .A1(n18403), .A2(n18459), .ZN(n18495) );
  NAND2_X1 U19645 ( .A1(n18412), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18718) );
  NOR2_X1 U19646 ( .A1(n18718), .A2(n17153), .ZN(n18595) );
  NAND2_X1 U19647 ( .A1(n18595), .A2(n17108), .ZN(n17130) );
  AOI22_X1 U19648 ( .A1(n18901), .A2(n17119), .B1(n18823), .B2(n17130), .ZN(
        n16548) );
  OAI21_X1 U19649 ( .B1(n18902), .B2(n16472), .A(n16548), .ZN(n16475) );
  OAI22_X1 U19650 ( .A1(n18454), .A2(n19360), .B1(n18779), .B2(n18755), .ZN(
        n18767) );
  INV_X1 U19651 ( .A(n18685), .ZN(n18611) );
  AOI21_X1 U19652 ( .B1(n19380), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19371), .ZN(n18876) );
  OAI22_X1 U19653 ( .A1(n19397), .A2(n18611), .B1(n18647), .B2(n18876), .ZN(
        n17143) );
  AOI21_X1 U19654 ( .B1(n16473), .B2(n18767), .A(n17143), .ZN(n18639) );
  NAND2_X1 U19655 ( .A1(n17114), .A2(n18660), .ZN(n18601) );
  NOR3_X1 U19656 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17126), .A3(
        n18601), .ZN(n16474) );
  AOI21_X1 U19657 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16475), .A(
        n16474), .ZN(n16476) );
  NAND2_X1 U19658 ( .A1(n18902), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17137) );
  OAI211_X1 U19659 ( .C1(n17141), .C2(n18799), .A(n16476), .B(n17137), .ZN(
        P3_U2833) );
  AOI22_X1 U19660 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19732), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19652), .ZN(n16477) );
  OAI21_X1 U19661 ( .B1(n19683), .B2(n16478), .A(n16477), .ZN(n16485) );
  INV_X1 U19662 ( .A(n15417), .ZN(n16481) );
  INV_X1 U19663 ( .A(n16479), .ZN(n16480) );
  OAI21_X1 U19664 ( .B1(n16481), .B2(n16480), .A(n19757), .ZN(n16483) );
  AOI21_X1 U19665 ( .B1(n19665), .B2(n16483), .A(n16482), .ZN(n16484) );
  AOI211_X1 U19666 ( .C1(n19734), .C2(n16486), .A(n16485), .B(n16484), .ZN(
        n16490) );
  INV_X1 U19667 ( .A(n16917), .ZN(n16487) );
  OAI22_X1 U19668 ( .A1(n16906), .A2(n19748), .B1(n16487), .B2(n19726), .ZN(
        n16488) );
  INV_X1 U19669 ( .A(n16488), .ZN(n16489) );
  NAND2_X1 U19670 ( .A1(n16490), .A2(n16489), .ZN(P2_U2833) );
  OR3_X1 U19671 ( .A1(n16492), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n16491), .ZN(n16496) );
  OAI22_X1 U19672 ( .A1(n19911), .A2(n19641), .B1(n20534), .B2(n19736), .ZN(
        n16494) );
  NOR2_X1 U19673 ( .A1(n19928), .A2(n19651), .ZN(n16493) );
  NOR2_X1 U19674 ( .A1(n16494), .A2(n16493), .ZN(n16495) );
  AND2_X1 U19675 ( .A1(n16496), .A2(n16495), .ZN(n16501) );
  OAI221_X1 U19676 ( .B1(n16499), .B2(n16498), .C1(n16499), .C2(n16497), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16500) );
  OAI211_X1 U19677 ( .C1(n16502), .C2(n17009), .A(n16501), .B(n16500), .ZN(
        P2_U3029) );
  NAND2_X1 U19678 ( .A1(n16504), .A2(n16503), .ZN(n16510) );
  AOI21_X1 U19679 ( .B1(n16510), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n16505), .ZN(n16506) );
  AOI211_X1 U19680 ( .C1(n16508), .C2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n16507), .B(n16506), .ZN(n16509) );
  AOI21_X1 U19681 ( .B1(n16510), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16509), .ZN(n16511) );
  AOI222_X1 U19682 ( .A1(n16513), .A2(n16512), .B1(n16513), .B2(n16511), .C1(
        n16512), .C2(n16511), .ZN(n16516) );
  INV_X1 U19683 ( .A(n16514), .ZN(n16515) );
  AOI222_X1 U19684 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16516), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16515), .C1(n16516), 
        .C2(n16515), .ZN(n16519) );
  AOI211_X1 U19685 ( .C1(n16519), .C2(n20854), .A(n16518), .B(n16517), .ZN(
        n16526) );
  NOR2_X1 U19686 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n16521) );
  OAI211_X1 U19687 ( .C1(n16522), .C2(n16521), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n16520), .ZN(n16524) );
  NOR2_X1 U19688 ( .A1(n16524), .A2(n16523), .ZN(n16525) );
  AND2_X1 U19689 ( .A1(n16526), .A2(n16525), .ZN(n16533) );
  INV_X1 U19690 ( .A(n16537), .ZN(n16532) );
  OR2_X1 U19691 ( .A1(n21051), .A2(n16527), .ZN(n16531) );
  OR2_X1 U19692 ( .A1(n16528), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21052) );
  NOR3_X1 U19693 ( .A1(n13135), .A2(n16529), .A3(n21052), .ZN(n16530) );
  AOI21_X1 U19694 ( .B1(n16532), .B2(n16531), .A(n16530), .ZN(n16847) );
  OAI21_X1 U19695 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n16533), .A(n16847), 
        .ZN(n16843) );
  INV_X1 U19696 ( .A(n16533), .ZN(n16538) );
  OAI211_X1 U19697 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21051), .A(n16535), 
        .B(n16534), .ZN(n16536) );
  AOI211_X1 U19698 ( .C1(n16538), .C2(n16537), .A(n16536), .B(n20963), .ZN(
        n16542) );
  NAND2_X1 U19699 ( .A1(n21054), .A2(n16539), .ZN(n16540) );
  AOI21_X1 U19700 ( .B1(n16540), .B2(n16843), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n16541) );
  AOI21_X1 U19701 ( .B1(n16843), .B2(n16542), .A(n16541), .ZN(P1_U3161) );
  INV_X1 U19702 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17109) );
  NAND2_X1 U19703 ( .A1(n17108), .A2(n17109), .ZN(n17125) );
  NAND2_X1 U19704 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16543), .ZN(
        n17094) );
  NAND2_X1 U19705 ( .A1(n18227), .A2(n16544), .ZN(n16545) );
  NOR2_X1 U19706 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16545), .ZN(
        n17092) );
  NOR2_X1 U19707 ( .A1(n18887), .A2(n18710), .ZN(n18893) );
  INV_X1 U19708 ( .A(n18893), .ZN(n18816) );
  OAI22_X1 U19709 ( .A1(n17108), .A2(n18816), .B1(n16546), .B2(n18887), .ZN(
        n16547) );
  NOR2_X1 U19710 ( .A1(n18892), .A2(n16547), .ZN(n17142) );
  AOI21_X1 U19711 ( .B1(n17142), .B2(n16548), .A(n17109), .ZN(n16549) );
  AOI21_X1 U19712 ( .B1(n18822), .B2(n17121), .A(n16549), .ZN(n16550) );
  NAND2_X1 U19713 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18902), .ZN(n17115) );
  OAI211_X1 U19714 ( .C1(n18601), .C2(n17125), .A(n16550), .B(n17115), .ZN(
        P3_U2832) );
  NAND2_X1 U19715 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20973), .ZN(n16553) );
  INV_X1 U19716 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20969) );
  NOR2_X1 U19717 ( .A1(n20972), .A2(n20969), .ZN(n20974) );
  INV_X1 U19718 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20630) );
  INV_X1 U19719 ( .A(HOLD), .ZN(n20971) );
  NOR2_X1 U19720 ( .A1(n20630), .A2(n20971), .ZN(n16551) );
  INV_X1 U19721 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20982) );
  OAI22_X1 U19722 ( .A1(n20974), .A2(n16551), .B1(n20982), .B2(n20971), .ZN(
        n16552) );
  NAND3_X1 U19723 ( .A1(n16554), .A2(n16553), .A3(n16552), .ZN(P1_U3195) );
  AND2_X1 U19724 ( .A1(n20737), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AOI221_X1 U19725 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n17069), .C1(n19598), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(P2_STATE2_REG_2__SCAN_IN), .ZN(
        n20488) );
  NOR3_X1 U19726 ( .A1(n17082), .A2(n16556), .A3(n20488), .ZN(P2_U3178) );
  INV_X1 U19727 ( .A(n16555), .ZN(n20619) );
  AOI221_X1 U19728 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16556), .C1(n20619), .C2(
        n16556), .A(n20425), .ZN(n20616) );
  INV_X1 U19729 ( .A(n20616), .ZN(n20613) );
  NOR2_X1 U19730 ( .A1(n17068), .A2(n20613), .ZN(P2_U3047) );
  INV_X1 U19731 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18917) );
  INV_X1 U19732 ( .A(n16562), .ZN(n17950) );
  NAND2_X1 U19733 ( .A1(n16561), .A2(n17950), .ZN(n18091) );
  INV_X1 U19734 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18173) );
  AOI21_X1 U19735 ( .B1(n17950), .B2(n18954), .A(P3_EAX_REG_0__SCAN_IN), .ZN(
        n16565) );
  OAI222_X1 U19736 ( .A1(n18917), .A2(n18091), .B1(n17945), .B2(n16565), .C1(
        n18098), .C2(n16564), .ZN(P3_U2735) );
  AOI22_X1 U19737 ( .A1(n20684), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20705), .ZN(n16572) );
  AOI21_X1 U19738 ( .B1(n16578), .B2(n16566), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n16569) );
  OAI22_X1 U19739 ( .A1(n16569), .A2(n16568), .B1(n20666), .B2(n16567), .ZN(
        n16570) );
  AOI21_X1 U19740 ( .B1(n16642), .B2(n20676), .A(n16570), .ZN(n16571) );
  OAI211_X1 U19741 ( .C1(n16573), .C2(n20703), .A(n16572), .B(n16571), .ZN(
        P1_U2820) );
  OAI22_X1 U19742 ( .A1(n20707), .A2(n14695), .B1(n16574), .B2(n20703), .ZN(
        n16575) );
  INV_X1 U19743 ( .A(n16575), .ZN(n16576) );
  OAI21_X1 U19744 ( .B1(n20666), .B2(n16724), .A(n16576), .ZN(n16577) );
  AOI211_X1 U19745 ( .C1(n20705), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20660), .B(n16577), .ZN(n16581) );
  AOI22_X1 U19746 ( .A1(n16579), .A2(n20676), .B1(n16578), .B2(n21007), .ZN(
        n16580) );
  OAI211_X1 U19747 ( .C1(n21007), .C2(n16582), .A(n16581), .B(n16580), .ZN(
        P1_U2822) );
  INV_X1 U19748 ( .A(n16583), .ZN(n16660) );
  AOI22_X1 U19749 ( .A1(n20684), .A2(P1_EBX_REG_16__SCAN_IN), .B1(n16660), 
        .B2(n20687), .ZN(n16584) );
  OAI21_X1 U19750 ( .B1(n20666), .B2(n16748), .A(n16584), .ZN(n16585) );
  AOI211_X1 U19751 ( .C1(n20705), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20660), .B(n16585), .ZN(n16592) );
  INV_X1 U19752 ( .A(n16586), .ZN(n16661) );
  OR2_X1 U19753 ( .A1(n16588), .A2(n16587), .ZN(n16600) );
  INV_X1 U19754 ( .A(n16600), .ZN(n16607) );
  AOI22_X1 U19755 ( .A1(n16661), .A2(n20676), .B1(n16607), .B2(
        P1_REIP_REG_16__SCAN_IN), .ZN(n16591) );
  NAND2_X1 U19756 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n16589) );
  OAI211_X1 U19757 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(P1_REIP_REG_16__SCAN_IN), .A(n16593), .B(n16589), .ZN(n16590) );
  NAND3_X1 U19758 ( .A1(n16592), .A2(n16591), .A3(n16590), .ZN(P1_U2824) );
  INV_X1 U19759 ( .A(n16593), .ZN(n16605) );
  AOI22_X1 U19760 ( .A1(n16749), .A2(n20700), .B1(n20684), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n16594) );
  OAI211_X1 U19761 ( .C1(n16596), .C2(n16595), .A(n16594), .B(n20702), .ZN(
        n16597) );
  AOI21_X1 U19762 ( .B1(n16598), .B2(n20687), .A(n16597), .ZN(n16604) );
  INV_X1 U19763 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n16599) );
  OAI22_X1 U19764 ( .A1(n21064), .A2(n16601), .B1(n16600), .B2(n16599), .ZN(
        n16602) );
  INV_X1 U19765 ( .A(n16602), .ZN(n16603) );
  OAI211_X1 U19766 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n16605), .A(n16604), 
        .B(n16603), .ZN(P1_U2825) );
  AOI22_X1 U19767 ( .A1(n16638), .A2(n20700), .B1(n20684), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n16610) );
  AOI22_X1 U19768 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20705), .B1(
        n16664), .B2(n20687), .ZN(n16609) );
  INV_X1 U19769 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n16760) );
  OAI21_X1 U19770 ( .B1(n16619), .B2(n16760), .A(n21002), .ZN(n16606) );
  AOI22_X1 U19771 ( .A1(n16665), .A2(n20676), .B1(n16607), .B2(n16606), .ZN(
        n16608) );
  NAND4_X1 U19772 ( .A1(n16610), .A2(n16609), .A3(n16608), .A4(n20702), .ZN(
        P1_U2826) );
  NAND2_X1 U19773 ( .A1(n20683), .A2(n16611), .ZN(n16621) );
  AOI21_X1 U19774 ( .B1(n20705), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20660), .ZN(n16612) );
  OAI21_X1 U19775 ( .B1(n20703), .B2(n16613), .A(n16612), .ZN(n16614) );
  AOI21_X1 U19776 ( .B1(n20684), .B2(P1_EBX_REG_13__SCAN_IN), .A(n16614), .ZN(
        n16615) );
  OAI21_X1 U19777 ( .B1(n16758), .B2(n20666), .A(n16615), .ZN(n16616) );
  AOI21_X1 U19778 ( .B1(n16617), .B2(n20676), .A(n16616), .ZN(n16618) );
  OAI221_X1 U19779 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n16619), .C1(n16760), 
        .C2(n16621), .A(n16618), .ZN(P1_U2827) );
  AOI22_X1 U19780 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20705), .B1(
        n16670), .B2(n20687), .ZN(n16629) );
  INV_X1 U19781 ( .A(n16620), .ZN(n16671) );
  AOI221_X1 U19782 ( .B1(n16623), .B2(n20998), .C1(n16622), .C2(n20998), .A(
        n16621), .ZN(n16627) );
  OAI22_X1 U19783 ( .A1(n16625), .A2(n20666), .B1(n16624), .B2(n20707), .ZN(
        n16626) );
  AOI211_X1 U19784 ( .C1(n16671), .C2(n20676), .A(n16627), .B(n16626), .ZN(
        n16628) );
  NAND3_X1 U19785 ( .A1(n16629), .A2(n16628), .A3(n20702), .ZN(P1_U2828) );
  NAND3_X1 U19786 ( .A1(n16630), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .ZN(n16637) );
  INV_X1 U19787 ( .A(n16631), .ZN(n16770) );
  AOI22_X1 U19788 ( .A1(n16770), .A2(n20700), .B1(n20684), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n16632) );
  OAI21_X1 U19789 ( .B1(n16682), .B2(n20703), .A(n16632), .ZN(n16633) );
  AOI211_X1 U19790 ( .C1(n20705), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20660), .B(n16633), .ZN(n16636) );
  AOI22_X1 U19791 ( .A1(n16679), .A2(n20676), .B1(n16634), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16635) );
  OAI211_X1 U19792 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n16637), .A(n16636), 
        .B(n16635), .ZN(P1_U2829) );
  INV_X1 U19793 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n16640) );
  AOI22_X1 U19794 ( .A1(n16665), .A2(n20718), .B1(n20717), .B2(n16638), .ZN(
        n16639) );
  OAI21_X1 U19795 ( .B1(n20721), .B2(n16640), .A(n16639), .ZN(P1_U2858) );
  INV_X1 U19796 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U19797 ( .A1(n16647), .A2(n16641), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16645), .ZN(n16644) );
  AOI22_X1 U19798 ( .A1(n16642), .A2(n16649), .B1(n16648), .B2(DATAI_20_), 
        .ZN(n16643) );
  OAI211_X1 U19799 ( .C1(n16652), .C2(n17189), .A(n16644), .B(n16643), .ZN(
        P1_U2884) );
  INV_X1 U19800 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n21081) );
  AOI22_X1 U19801 ( .A1(n16647), .A2(n16646), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16645), .ZN(n16651) );
  AOI22_X1 U19802 ( .A1(n16661), .A2(n16649), .B1(n16648), .B2(DATAI_16_), 
        .ZN(n16650) );
  OAI211_X1 U19803 ( .C1(n16652), .C2(n21081), .A(n16651), .B(n16650), .ZN(
        P1_U2888) );
  INV_X1 U19804 ( .A(n16653), .ZN(n16655) );
  AOI21_X1 U19805 ( .B1(n14921), .B2(n16655), .A(n16654), .ZN(n16751) );
  MUX2_X1 U19806 ( .A(n12128), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .S(
        n16656), .Z(n16750) );
  NOR2_X1 U19807 ( .A1(n16753), .A2(n16739), .ZN(n16659) );
  OAI22_X1 U19808 ( .A1(n16659), .A2(n16658), .B1(n16753), .B2(n16657), .ZN(
        n16743) );
  AOI22_X1 U19809 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16663) );
  AOI22_X1 U19810 ( .A1(n16661), .A2(n20791), .B1(n16660), .B2(n16669), .ZN(
        n16662) );
  OAI211_X1 U19811 ( .C1(n21068), .C2(n16743), .A(n16663), .B(n16662), .ZN(
        P1_U2983) );
  AOI22_X1 U19812 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16667) );
  AOI22_X1 U19813 ( .A1(n16665), .A2(n20791), .B1(n16664), .B2(n16669), .ZN(
        n16666) );
  OAI211_X1 U19814 ( .C1(n16668), .C2(n21068), .A(n16667), .B(n16666), .ZN(
        P1_U2985) );
  AOI22_X1 U19815 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16673) );
  AOI22_X1 U19816 ( .A1(n16671), .A2(n20791), .B1(n16670), .B2(n16669), .ZN(
        n16672) );
  OAI211_X1 U19817 ( .C1(n16674), .C2(n21068), .A(n16673), .B(n16672), .ZN(
        P1_U2987) );
  AOI22_X1 U19818 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16681) );
  NOR2_X1 U19819 ( .A1(n16675), .A2(n12132), .ZN(n16677) );
  MUX2_X1 U19820 ( .A(n16677), .B(n16676), .S(n15123), .Z(n16678) );
  XNOR2_X1 U19821 ( .A(n16678), .B(n16776), .ZN(n16773) );
  AOI22_X1 U19822 ( .A1(n16773), .A2(n20792), .B1(n20791), .B2(n16679), .ZN(
        n16680) );
  OAI211_X1 U19823 ( .C1(n16695), .C2(n16682), .A(n16681), .B(n16680), .ZN(
        P1_U2988) );
  AOI22_X1 U19824 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16688) );
  OAI21_X1 U19825 ( .B1(n16685), .B2(n16684), .A(n16683), .ZN(n16816) );
  INV_X1 U19826 ( .A(n16816), .ZN(n16686) );
  AOI22_X1 U19827 ( .A1(n16686), .A2(n20792), .B1(n20791), .B2(n20668), .ZN(
        n16687) );
  OAI211_X1 U19828 ( .C1(n16695), .C2(n20661), .A(n16688), .B(n16687), .ZN(
        P1_U2992) );
  AOI22_X1 U19829 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16694) );
  OAI21_X1 U19830 ( .B1(n16691), .B2(n16690), .A(n16689), .ZN(n16692) );
  INV_X1 U19831 ( .A(n16692), .ZN(n16825) );
  AOI22_X1 U19832 ( .A1(n16825), .A2(n20792), .B1(n20791), .B2(n20677), .ZN(
        n16693) );
  OAI211_X1 U19833 ( .C1(n16695), .C2(n20674), .A(n16694), .B(n16693), .ZN(
        P1_U2993) );
  AOI22_X1 U19834 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16701) );
  OAI21_X1 U19835 ( .B1(n16698), .B2(n16697), .A(n16696), .ZN(n16699) );
  INV_X1 U19836 ( .A(n16699), .ZN(n16834) );
  AOI22_X1 U19837 ( .A1(n16834), .A2(n20792), .B1(n20791), .B2(n20714), .ZN(
        n16700) );
  OAI211_X1 U19838 ( .C1(n16695), .C2(n20685), .A(n16701), .B(n16700), .ZN(
        P1_U2994) );
  INV_X1 U19839 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21014) );
  INV_X1 U19840 ( .A(n16702), .ZN(n16707) );
  INV_X1 U19841 ( .A(n16703), .ZN(n16706) );
  INV_X1 U19842 ( .A(n16704), .ZN(n16705) );
  AOI222_X1 U19843 ( .A1(n16707), .A2(n20806), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16706), .C1(n20849), .C2(
        n16705), .ZN(n16711) );
  OAI211_X1 U19844 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16709), .B(n16708), .ZN(
        n16710) );
  OAI211_X1 U19845 ( .C1(n21014), .C2(n16817), .A(n16711), .B(n16710), .ZN(
        P1_U3009) );
  INV_X1 U19846 ( .A(n16712), .ZN(n16714) );
  AOI22_X1 U19847 ( .A1(n16714), .A2(n20806), .B1(n20849), .B2(n16713), .ZN(
        n16720) );
  NOR2_X1 U19848 ( .A1(n16817), .A2(n21009), .ZN(n16715) );
  AOI221_X1 U19849 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16718), 
        .C1(n16717), .C2(n16716), .A(n16715), .ZN(n16719) );
  NAND2_X1 U19850 ( .A1(n16720), .A2(n16719), .ZN(P1_U3012) );
  AOI21_X1 U19851 ( .B1(n16801), .B2(n16759), .A(n16800), .ZN(n16721) );
  OAI21_X1 U19852 ( .B1(n16722), .B2(n16799), .A(n16721), .ZN(n16740) );
  AOI21_X1 U19853 ( .B1(n16807), .B2(n16723), .A(n16740), .ZN(n16737) );
  NOR3_X1 U19854 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16730), .A3(
        n16723), .ZN(n16727) );
  OAI22_X1 U19855 ( .A1(n16725), .A2(n20844), .B1(n20836), .B2(n16724), .ZN(
        n16726) );
  AOI211_X1 U19856 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n21060), .A(n16727), 
        .B(n16726), .ZN(n16728) );
  OAI21_X1 U19857 ( .B1(n16737), .B2(n16729), .A(n16728), .ZN(P1_U3013) );
  NOR2_X1 U19858 ( .A1(n16730), .A2(n16741), .ZN(n16754) );
  AOI21_X1 U19859 ( .B1(n16738), .B2(n16754), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16736) );
  INV_X1 U19860 ( .A(n16731), .ZN(n16733) );
  AOI22_X1 U19861 ( .A1(n16733), .A2(n20806), .B1(n20849), .B2(n16732), .ZN(
        n16735) );
  NAND2_X1 U19862 ( .A1(n21060), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16734) );
  OAI211_X1 U19863 ( .C1(n16737), .C2(n16736), .A(n16735), .B(n16734), .ZN(
        P1_U3014) );
  NOR2_X1 U19864 ( .A1(n16739), .A2(n16738), .ZN(n16745) );
  AOI21_X1 U19865 ( .B1(n16741), .B2(n16807), .A(n16740), .ZN(n16757) );
  OAI22_X1 U19866 ( .A1(n16743), .A2(n20844), .B1(n16757), .B2(n16742), .ZN(
        n16744) );
  AOI21_X1 U19867 ( .B1(n16745), .B2(n16754), .A(n16744), .ZN(n16747) );
  NAND2_X1 U19868 ( .A1(n21060), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16746) );
  OAI211_X1 U19869 ( .C1(n20836), .C2(n16748), .A(n16747), .B(n16746), .ZN(
        P1_U3015) );
  AOI22_X1 U19870 ( .A1(n21060), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n20849), 
        .B2(n16749), .ZN(n16756) );
  NOR2_X1 U19871 ( .A1(n16751), .A2(n16750), .ZN(n16752) );
  AOI22_X1 U19872 ( .A1(n21059), .A2(n20806), .B1(n12128), .B2(n16754), .ZN(
        n16755) );
  OAI211_X1 U19873 ( .C1(n16757), .C2(n12128), .A(n16756), .B(n16755), .ZN(
        P1_U3016) );
  NOR2_X1 U19874 ( .A1(n16758), .A2(n20836), .ZN(n16764) );
  NAND2_X1 U19875 ( .A1(n20838), .A2(n16759), .ZN(n16761) );
  OAI22_X1 U19876 ( .A1(n16762), .A2(n16761), .B1(n16760), .B2(n16817), .ZN(
        n16763) );
  AOI211_X1 U19877 ( .C1(n16765), .C2(n20806), .A(n16764), .B(n16763), .ZN(
        n16767) );
  OAI211_X1 U19878 ( .C1(n16769), .C2(n16768), .A(n16767), .B(n16766), .ZN(
        P1_U3018) );
  INV_X1 U19879 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16776) );
  AOI22_X1 U19880 ( .A1(n21060), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20849), 
        .B2(n16770), .ZN(n16775) );
  NOR2_X1 U19881 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16778), .ZN(
        n16772) );
  AOI22_X1 U19882 ( .A1(n16773), .A2(n20806), .B1(n16772), .B2(n16771), .ZN(
        n16774) );
  OAI211_X1 U19883 ( .C1(n16777), .C2(n16776), .A(n16775), .B(n16774), .ZN(
        P1_U3020) );
  NAND2_X1 U19884 ( .A1(n16785), .A2(n16823), .ZN(n16797) );
  AOI22_X1 U19885 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16779), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n12132), .ZN(n16790) );
  AOI22_X1 U19886 ( .A1(n21060), .A2(P1_REIP_REG_10__SCAN_IN), .B1(n20849), 
        .B2(n16780), .ZN(n16789) );
  AOI211_X1 U19887 ( .C1(n16782), .C2(n16801), .A(n16781), .B(n16800), .ZN(
        n16786) );
  INV_X1 U19888 ( .A(n16783), .ZN(n16784) );
  AOI21_X1 U19889 ( .B1(n16786), .B2(n16785), .A(n16784), .ZN(n16793) );
  AOI22_X1 U19890 ( .A1(n16787), .A2(n20806), .B1(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16793), .ZN(n16788) );
  OAI211_X1 U19891 ( .C1(n16797), .C2(n16790), .A(n16789), .B(n16788), .ZN(
        P1_U3021) );
  AOI22_X1 U19892 ( .A1(n21060), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n20849), 
        .B2(n16791), .ZN(n16796) );
  INV_X1 U19893 ( .A(n16792), .ZN(n16794) );
  AOI22_X1 U19894 ( .A1(n16794), .A2(n20806), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16793), .ZN(n16795) );
  OAI211_X1 U19895 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16797), .A(
        n16796), .B(n16795), .ZN(P1_U3022) );
  OR2_X1 U19896 ( .A1(n20796), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16837) );
  NOR2_X1 U19897 ( .A1(n16798), .A2(n16799), .ZN(n16805) );
  NAND2_X1 U19898 ( .A1(n16801), .A2(n20796), .ZN(n16803) );
  OR2_X1 U19899 ( .A1(n16799), .A2(n20812), .ZN(n16802) );
  AOI21_X1 U19900 ( .B1(n16801), .B2(n20813), .A(n16800), .ZN(n20821) );
  AND2_X1 U19901 ( .A1(n16802), .A2(n20821), .ZN(n20798) );
  NAND2_X1 U19902 ( .A1(n16803), .A2(n20798), .ZN(n16804) );
  INV_X1 U19903 ( .A(n16833), .ZN(n16806) );
  OAI21_X1 U19904 ( .B1(n15151), .B2(n16837), .A(n16806), .ZN(n16824) );
  AOI21_X1 U19905 ( .B1(n16808), .B2(n16807), .A(n16824), .ZN(n16820) );
  INV_X1 U19906 ( .A(n16809), .ZN(n16813) );
  OAI22_X1 U19907 ( .A1(n16810), .A2(n20836), .B1(n13931), .B2(n16817), .ZN(
        n16812) );
  NAND2_X1 U19908 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16823), .ZN(
        n16822) );
  AOI221_X1 U19909 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16815), .C2(n16821), .A(
        n16822), .ZN(n16811) );
  AOI211_X1 U19910 ( .C1(n16813), .C2(n20806), .A(n16812), .B(n16811), .ZN(
        n16814) );
  OAI21_X1 U19911 ( .B1(n16820), .B2(n16815), .A(n16814), .ZN(P1_U3023) );
  INV_X1 U19912 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20670) );
  OAI222_X1 U19913 ( .A1(n20665), .A2(n20836), .B1(n16817), .B2(n20670), .C1(
        n20844), .C2(n16816), .ZN(n16818) );
  INV_X1 U19914 ( .A(n16818), .ZN(n16819) );
  OAI221_X1 U19915 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16822), .C1(
        n16821), .C2(n16820), .A(n16819), .ZN(P1_U3024) );
  INV_X1 U19916 ( .A(n16823), .ZN(n16828) );
  AOI22_X1 U19917 ( .A1(n21060), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20849), 
        .B2(n20671), .ZN(n16827) );
  AOI22_X1 U19918 ( .A1(n16825), .A2(n20806), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16824), .ZN(n16826) );
  OAI211_X1 U19919 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16828), .A(
        n16827), .B(n16826), .ZN(P1_U3025) );
  NAND2_X1 U19920 ( .A1(n20812), .A2(n16829), .ZN(n20810) );
  OAI21_X1 U19921 ( .B1(n20697), .B2(n20696), .A(n16830), .ZN(n16832) );
  AND2_X1 U19922 ( .A1(n16832), .A2(n16831), .ZN(n20713) );
  AOI22_X1 U19923 ( .A1(n21060), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20849), 
        .B2(n20713), .ZN(n16836) );
  AOI22_X1 U19924 ( .A1(n16834), .A2(n20806), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16833), .ZN(n16835) );
  OAI211_X1 U19925 ( .C1(n16837), .C2(n20810), .A(n16836), .B(n16835), .ZN(
        P1_U3026) );
  OR3_X1 U19926 ( .A1(n16840), .A2(n16839), .A3(n16838), .ZN(n16841) );
  OAI21_X1 U19927 ( .B1(n16842), .B2(n11894), .A(n16841), .ZN(P1_U3468) );
  NAND2_X1 U19928 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16843), .ZN(n16852) );
  INV_X1 U19929 ( .A(n21054), .ZN(n16844) );
  AOI21_X1 U19930 ( .B1(n20905), .B2(n21051), .A(n16844), .ZN(n16850) );
  NAND4_X1 U19931 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n13658), .A4(n21051), .ZN(n16845) );
  AND2_X1 U19932 ( .A1(n16846), .A2(n16845), .ZN(n20964) );
  AOI21_X1 U19933 ( .B1(n20964), .B2(n16848), .A(n16847), .ZN(n16849) );
  AOI211_X1 U19934 ( .C1(n20962), .C2(n16852), .A(n16850), .B(n16849), .ZN(
        P1_U3162) );
  AOI21_X1 U19935 ( .B1(n16852), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n16851), 
        .ZN(n16853) );
  INV_X1 U19936 ( .A(n16853), .ZN(P1_U3466) );
  OAI22_X1 U19937 ( .A1(n16854), .A2(n19684), .B1(n20548), .B2(n19737), .ZN(
        n16855) );
  INV_X1 U19938 ( .A(n16855), .ZN(n16867) );
  AOI22_X1 U19939 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19744), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19732), .ZN(n16866) );
  INV_X1 U19940 ( .A(n16856), .ZN(n16857) );
  OAI22_X1 U19941 ( .A1(n16858), .A2(n19748), .B1(n16857), .B2(n19726), .ZN(
        n16859) );
  INV_X1 U19942 ( .A(n16859), .ZN(n16865) );
  NAND3_X1 U19943 ( .A1(n16860), .A2(n19753), .A3(n16861), .ZN(n16862) );
  NAND3_X1 U19944 ( .A1(n16863), .A2(n19757), .A3(n16862), .ZN(n16864) );
  NAND4_X1 U19945 ( .A1(n16867), .A2(n16866), .A3(n16865), .A4(n16864), .ZN(
        P2_U2829) );
  OAI21_X1 U19946 ( .B1(n16868), .B2(n16869), .A(n19757), .ZN(n16870) );
  NAND2_X1 U19947 ( .A1(n16870), .A2(n19665), .ZN(n16880) );
  INV_X1 U19948 ( .A(n16883), .ZN(n16873) );
  INV_X1 U19949 ( .A(n16871), .ZN(n16872) );
  AOI211_X1 U19950 ( .C1(n16873), .C2(P2_EBX_REG_25__SCAN_IN), .A(n16872), .B(
        n19684), .ZN(n16879) );
  NAND2_X1 U19951 ( .A1(n16874), .A2(n19692), .ZN(n16876) );
  AOI22_X1 U19952 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19732), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19652), .ZN(n16875) );
  OAI211_X1 U19953 ( .C1(n19683), .C2(n16877), .A(n16876), .B(n16875), .ZN(
        n16878) );
  AOI211_X1 U19954 ( .C1(n16860), .C2(n16880), .A(n16879), .B(n16878), .ZN(
        n16881) );
  OAI21_X1 U19955 ( .B1(n16882), .B2(n19726), .A(n16881), .ZN(P2_U2830) );
  AOI211_X1 U19956 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n16884), .A(n19684), .B(
        n16883), .ZN(n16887) );
  AOI22_X1 U19957 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19732), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19652), .ZN(n16885) );
  INV_X1 U19958 ( .A(n16885), .ZN(n16886) );
  AOI211_X1 U19959 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n19744), .A(n16887), .B(
        n16886), .ZN(n16896) );
  INV_X1 U19960 ( .A(n16888), .ZN(n16894) );
  INV_X1 U19961 ( .A(n16889), .ZN(n16890) );
  NOR2_X1 U19962 ( .A1(n9934), .A2(n16890), .ZN(n16892) );
  AOI211_X1 U19963 ( .C1(n16892), .C2(n15403), .A(n19730), .B(n16868), .ZN(
        n16893) );
  AOI21_X1 U19964 ( .B1(n19692), .B2(n16894), .A(n16893), .ZN(n16895) );
  OAI211_X1 U19965 ( .C1(n16897), .C2(n19726), .A(n16896), .B(n16895), .ZN(
        P2_U2831) );
  AOI22_X1 U19966 ( .A1(n19784), .A2(n16899), .B1(n16898), .B2(n19796), .ZN(
        P2_U2856) );
  AOI22_X1 U19967 ( .A1(n16901), .A2(n19793), .B1(n19784), .B2(n16900), .ZN(
        n16902) );
  OAI21_X1 U19968 ( .B1(n19784), .B2(n16903), .A(n16902), .ZN(P2_U2864) );
  AOI21_X1 U19969 ( .B1(n16904), .B2(n15562), .A(n9651), .ZN(n16918) );
  AOI22_X1 U19970 ( .A1(n16918), .A2(n19793), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n19796), .ZN(n16905) );
  OAI21_X1 U19971 ( .B1(n19796), .B2(n16906), .A(n16905), .ZN(P2_U2865) );
  AOI21_X1 U19972 ( .B1(n16907), .B2(n15567), .A(n15561), .ZN(n16924) );
  AOI22_X1 U19973 ( .A1(n16924), .A2(n19793), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n19796), .ZN(n16908) );
  OAI21_X1 U19974 ( .B1(n19796), .B2(n16909), .A(n16908), .ZN(P2_U2867) );
  AND2_X1 U19975 ( .A1(n16911), .A2(n16910), .ZN(n16912) );
  NOR2_X1 U19976 ( .A1(n9689), .A2(n16912), .ZN(n16930) );
  NOR2_X1 U19977 ( .A1(n19784), .A2(n16913), .ZN(n16914) );
  AOI21_X1 U19978 ( .B1(n16930), .B2(n19793), .A(n16914), .ZN(n16915) );
  OAI21_X1 U19979 ( .B1(n19796), .B2(n16916), .A(n16915), .ZN(P2_U2869) );
  AOI22_X1 U19980 ( .A1(n19802), .A2(n19833), .B1(n19858), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16921) );
  AOI22_X1 U19981 ( .A1(n19804), .A2(BUF2_REG_22__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16920) );
  AOI22_X1 U19982 ( .A1(n16918), .A2(n19848), .B1(n19859), .B2(n16917), .ZN(
        n16919) );
  NAND3_X1 U19983 ( .A1(n16921), .A2(n16920), .A3(n16919), .ZN(P2_U2897) );
  AOI22_X1 U19984 ( .A1(n19802), .A2(n19845), .B1(n19858), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16927) );
  AOI22_X1 U19985 ( .A1(n19804), .A2(BUF2_REG_20__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16926) );
  INV_X1 U19986 ( .A(n16922), .ZN(n16923) );
  AOI22_X1 U19987 ( .A1(n16924), .A2(n19848), .B1(n19859), .B2(n16923), .ZN(
        n16925) );
  NAND3_X1 U19988 ( .A1(n16927), .A2(n16926), .A3(n16925), .ZN(P2_U2899) );
  AOI22_X1 U19989 ( .A1(n19802), .A2(n16928), .B1(n19858), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U19990 ( .A1(n19804), .A2(BUF2_REG_18__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U19991 ( .A1(n16930), .A2(n19848), .B1(n19859), .B2(n16929), .ZN(
        n16931) );
  NAND3_X1 U19992 ( .A1(n16933), .A2(n16932), .A3(n16931), .ZN(P2_U2901) );
  AOI22_X1 U19993 ( .A1(n16942), .A2(n16934), .B1(n19903), .B2(
        P2_REIP_REG_11__SCAN_IN), .ZN(n16940) );
  OAI22_X1 U19994 ( .A1(n16936), .A2(n16957), .B1(n16955), .B2(n16935), .ZN(
        n16937) );
  AOI21_X1 U19995 ( .B1(n16946), .B2(n16938), .A(n16937), .ZN(n16939) );
  OAI211_X1 U19996 ( .C1(n16950), .C2(n16941), .A(n16940), .B(n16939), .ZN(
        P2_U3003) );
  AOI22_X1 U19997 ( .A1(n16942), .A2(n19689), .B1(n19903), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n16948) );
  OAI22_X1 U19998 ( .A1(n16944), .A2(n16955), .B1(n16957), .B2(n16943), .ZN(
        n16945) );
  AOI21_X1 U19999 ( .B1(n16946), .B2(n19691), .A(n16945), .ZN(n16947) );
  OAI211_X1 U20000 ( .C1(n16950), .C2(n16949), .A(n16948), .B(n16947), .ZN(
        P2_U3005) );
  OAI21_X1 U20001 ( .B1(n16952), .B2(n19709), .A(n16951), .ZN(n16953) );
  AOI21_X1 U20002 ( .B1(n16954), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16953), .ZN(n16961) );
  OAI22_X1 U20003 ( .A1(n16958), .A2(n16957), .B1(n16956), .B2(n16955), .ZN(
        n16959) );
  INV_X1 U20004 ( .A(n16959), .ZN(n16960) );
  OAI211_X1 U20005 ( .C1(n13859), .C2(n19715), .A(n16961), .B(n16960), .ZN(
        P2_U3008) );
  NOR2_X1 U20006 ( .A1(n10889), .A2(n19736), .ZN(n16967) );
  OAI21_X1 U20007 ( .B1(n16964), .B2(n16963), .A(n16962), .ZN(n19812) );
  OAI22_X1 U20008 ( .A1(n19928), .A2(n19812), .B1(n16965), .B2(n16968), .ZN(
        n16966) );
  AOI211_X1 U20009 ( .C1(n16969), .C2(n16968), .A(n16967), .B(n16966), .ZN(
        n16974) );
  OAI22_X1 U20010 ( .A1(n16971), .A2(n19926), .B1(n19911), .B2(n16970), .ZN(
        n16972) );
  INV_X1 U20011 ( .A(n16972), .ZN(n16973) );
  OAI211_X1 U20012 ( .C1(n16975), .C2(n17009), .A(n16974), .B(n16973), .ZN(
        P2_U3031) );
  AOI211_X1 U20013 ( .C1(n21218), .C2(n16978), .A(n16977), .B(n16976), .ZN(
        n16980) );
  NOR2_X1 U20014 ( .A1(n19736), .A2(n15842), .ZN(n16979) );
  AOI211_X1 U20015 ( .C1(n19909), .C2(n16981), .A(n16980), .B(n16979), .ZN(
        n16986) );
  OAI22_X1 U20016 ( .A1(n16982), .A2(n19926), .B1(n19911), .B2(n19772), .ZN(
        n16983) );
  AOI21_X1 U20017 ( .B1(n16984), .B2(n19920), .A(n16983), .ZN(n16985) );
  OAI211_X1 U20018 ( .C1(n16987), .C2(n21218), .A(n16986), .B(n16985), .ZN(
        P2_U3032) );
  NOR2_X1 U20019 ( .A1(n15879), .A2(n19736), .ZN(n16992) );
  XNOR2_X1 U20020 ( .A(n16989), .B(n16988), .ZN(n19825) );
  OAI22_X1 U20021 ( .A1(n16990), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n19825), .B2(n19928), .ZN(n16991) );
  AOI211_X1 U20022 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16993), .A(
        n16992), .B(n16991), .ZN(n16996) );
  AOI22_X1 U20023 ( .A1(n16994), .A2(n17013), .B1(n19931), .B2(n19780), .ZN(
        n16995) );
  OAI211_X1 U20024 ( .C1(n16997), .C2(n17009), .A(n16996), .B(n16995), .ZN(
        P2_U3036) );
  NOR2_X1 U20025 ( .A1(n19736), .A2(n12689), .ZN(n17003) );
  OAI21_X1 U20026 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16998), .ZN(n16999) );
  OAI22_X1 U20027 ( .A1(n17001), .A2(n10683), .B1(n17000), .B2(n16999), .ZN(
        n17002) );
  AOI211_X1 U20028 ( .C1(n19909), .C2(n19828), .A(n17003), .B(n17002), .ZN(
        n17007) );
  AOI22_X1 U20029 ( .A1(n17005), .A2(n17013), .B1(n19931), .B2(n17004), .ZN(
        n17006) );
  OAI211_X1 U20030 ( .C1(n17009), .C2(n17008), .A(n17007), .B(n17006), .ZN(
        P2_U3038) );
  AOI22_X1 U20031 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17011), .B1(
        n19920), .B2(n17010), .ZN(n17021) );
  NAND2_X1 U20032 ( .A1(n17013), .A2(n17012), .ZN(n17019) );
  OR2_X1 U20033 ( .A1(n19911), .A2(n17014), .ZN(n17018) );
  OR2_X1 U20034 ( .A1(n19928), .A2(n17015), .ZN(n17016) );
  AND4_X1 U20035 ( .A1(n17019), .A2(n17018), .A3(n17017), .A4(n17016), .ZN(
        n17020) );
  OAI211_X1 U20036 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n17022), .A(
        n17021), .B(n17020), .ZN(P2_U3046) );
  NAND2_X1 U20037 ( .A1(n17023), .A2(n17027), .ZN(n17025) );
  AOI21_X1 U20038 ( .B1(n17033), .B2(n14482), .A(n10419), .ZN(n17024) );
  NAND2_X1 U20039 ( .A1(n17025), .A2(n17024), .ZN(n17030) );
  NAND3_X1 U20040 ( .A1(n17028), .A2(n17027), .A3(n17026), .ZN(n17029) );
  MUX2_X1 U20041 ( .A(n17030), .B(n17029), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n17031) );
  AOI21_X1 U20042 ( .B1(n10549), .B2(n17032), .A(n17031), .ZN(n20567) );
  INV_X1 U20043 ( .A(n17033), .ZN(n17036) );
  OAI211_X1 U20044 ( .C1(n17036), .C2(n17035), .A(n17034), .B(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17038) );
  OAI21_X1 U20045 ( .B1(n17038), .B2(n20605), .A(n17064), .ZN(n17040) );
  AOI21_X1 U20046 ( .B1(n20605), .B2(n17038), .A(n17037), .ZN(n17039) );
  AOI211_X1 U20047 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n20567), .A(
        n17040), .B(n17039), .ZN(n17043) );
  INV_X1 U20048 ( .A(n17043), .ZN(n17045) );
  NOR2_X1 U20049 ( .A1(n17064), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17041) );
  AOI21_X1 U20050 ( .B1(n17042), .B2(n17064), .A(n17041), .ZN(n17061) );
  OAI211_X1 U20051 ( .C1(n17043), .C2(n20597), .A(n17061), .B(n20588), .ZN(
        n17044) );
  OAI21_X1 U20052 ( .B1(n17045), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n17044), .ZN(n17067) );
  OR2_X1 U20053 ( .A1(P2_MORE_REG_SCAN_IN), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(
        n17057) );
  OAI22_X1 U20054 ( .A1(n17048), .A2(n17047), .B1(n10451), .B2(n17046), .ZN(
        n17056) );
  NAND2_X1 U20055 ( .A1(n17050), .A2(n17049), .ZN(n17053) );
  NAND2_X1 U20056 ( .A1(n17055), .A2(n17051), .ZN(n17052) );
  OAI211_X1 U20057 ( .C1(n17055), .C2(n17054), .A(n17053), .B(n17052), .ZN(
        n20618) );
  AOI211_X1 U20058 ( .C1(n17058), .C2(n17057), .A(n17056), .B(n20618), .ZN(
        n17059) );
  OAI21_X1 U20059 ( .B1(n17060), .B2(n17064), .A(n17059), .ZN(n17066) );
  NOR2_X1 U20060 ( .A1(n17064), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17063) );
  AOI21_X1 U20061 ( .B1(n17068), .B2(n20588), .A(n17061), .ZN(n17062) );
  AOI211_X1 U20062 ( .C1(n20567), .C2(n17064), .A(n17063), .B(n17062), .ZN(
        n17065) );
  AOI211_X1 U20063 ( .C1(n17068), .C2(n17067), .A(n17066), .B(n17065), .ZN(
        n17074) );
  INV_X1 U20064 ( .A(n17074), .ZN(n17072) );
  NOR3_X1 U20065 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19598), .A3(n17069), 
        .ZN(n17070) );
  AOI211_X1 U20066 ( .C1(n17073), .C2(n17072), .A(n17071), .B(n17070), .ZN(
        n17086) );
  AOI21_X1 U20067 ( .B1(n17074), .B2(n20495), .A(n19598), .ZN(n17079) );
  NAND3_X1 U20068 ( .A1(n12880), .A2(n17076), .A3(n17075), .ZN(n17078) );
  NAND3_X1 U20069 ( .A1(n17078), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n17077), 
        .ZN(n17080) );
  INV_X1 U20070 ( .A(n17080), .ZN(n17081) );
  AOI22_X1 U20071 ( .A1(n17083), .A2(n17082), .B1(n17081), .B2(n20509), .ZN(
        n17084) );
  AOI22_X1 U20072 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20490), .B1(n17084), 
        .B2(n19598), .ZN(n17085) );
  OAI211_X1 U20073 ( .C1(n20619), .C2(n17087), .A(n17086), .B(n17085), .ZN(
        P2_U3176) );
  NOR2_X1 U20074 ( .A1(n20490), .A2(n19598), .ZN(n17088) );
  OAI21_X1 U20075 ( .B1(n17088), .B2(n21204), .A(n17087), .ZN(P2_U3593) );
  INV_X1 U20076 ( .A(n17089), .ZN(n19359) );
  NOR2_X1 U20077 ( .A1(n17101), .A2(n17091), .ZN(n17106) );
  NOR2_X1 U20078 ( .A1(n18496), .A2(n17092), .ZN(n17100) );
  OAI21_X1 U20079 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18496), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17093) );
  OAI221_X1 U20080 ( .B1(n17109), .B2(n17094), .C1(n18496), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n17093), .ZN(n17099) );
  OAI21_X1 U20081 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17109), .A(
        n17094), .ZN(n17097) );
  NAND2_X1 U20082 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18496), .ZN(
        n17095) );
  OAI22_X1 U20083 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18496), .B1(
        n17095), .B2(n17109), .ZN(n17096) );
  OAI21_X1 U20084 ( .B1(n17100), .B2(n17097), .A(n17096), .ZN(n17098) );
  OAI21_X1 U20085 ( .B1(n17100), .B2(n17099), .A(n17098), .ZN(n17152) );
  INV_X1 U20086 ( .A(n18546), .ZN(n18489) );
  INV_X1 U20087 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17317) );
  INV_X1 U20088 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18213) );
  NAND2_X1 U20089 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18545) );
  NAND2_X1 U20090 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17492) );
  NAND2_X1 U20091 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18421) );
  NAND2_X1 U20092 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18381) );
  NAND3_X1 U20093 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17303) );
  INV_X1 U20094 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18242) );
  INV_X1 U20095 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19512) );
  NOR2_X1 U20096 ( .A1(n19512), .A2(n18890), .ZN(n17146) );
  NAND2_X1 U20097 ( .A1(n19577), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19432) );
  AOI21_X1 U20098 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18299), .A(
        n19302), .ZN(n18420) );
  OR2_X1 U20099 ( .A1(n17102), .A2(n18420), .ZN(n17117) );
  XNOR2_X1 U20100 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17104) );
  NOR2_X1 U20101 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18364), .ZN(
        n17131) );
  INV_X1 U20102 ( .A(n19432), .ZN(n18378) );
  NAND2_X1 U20103 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17133), .ZN(
        n17296) );
  AOI22_X1 U20104 ( .A1(n19302), .A2(n17102), .B1(n18378), .B2(n17296), .ZN(
        n17103) );
  NAND2_X1 U20105 ( .A1(n17103), .A2(n18587), .ZN(n17132) );
  NOR2_X1 U20106 ( .A1(n17131), .A2(n17132), .ZN(n17116) );
  OAI22_X1 U20107 ( .A1(n17117), .A2(n17104), .B1(n17116), .B2(n17317), .ZN(
        n17105) );
  AOI211_X1 U20108 ( .C1(n18427), .C2(n17655), .A(n17146), .B(n17105), .ZN(
        n17112) );
  NAND2_X1 U20109 ( .A1(n18068), .A2(n17106), .ZN(n18429) );
  INV_X1 U20110 ( .A(n17130), .ZN(n17120) );
  NAND2_X1 U20111 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17120), .ZN(
        n17107) );
  INV_X1 U20112 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19536) );
  XOR2_X1 U20113 ( .A(n17107), .B(n19536), .Z(n17149) );
  NOR2_X2 U20114 ( .A1(n19574), .A2(n17274), .ZN(n18550) );
  NAND4_X1 U20115 ( .A1(n17114), .A2(n17108), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n19536), .ZN(n17144) );
  OAI21_X1 U20116 ( .B1(n17109), .B2(n17119), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17110) );
  OAI21_X1 U20117 ( .B1(n18717), .B2(n17144), .A(n17110), .ZN(n17148) );
  AOI22_X1 U20118 ( .A1(n18498), .A2(n17149), .B1(n18550), .B2(n17148), .ZN(
        n17111) );
  OAI211_X1 U20119 ( .C1(n18471), .C2(n17152), .A(n17112), .B(n17111), .ZN(
        P3_U2799) );
  NAND2_X1 U20120 ( .A1(n17114), .A2(n18388), .ZN(n18231) );
  XNOR2_X1 U20121 ( .A(n9964), .B(n9698), .ZN(n17319) );
  OAI221_X1 U20122 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17117), .C1(
        n9964), .C2(n17116), .A(n17115), .ZN(n17118) );
  AOI21_X1 U20123 ( .B1(n18427), .B2(n17319), .A(n17118), .ZN(n17124) );
  NAND2_X1 U20124 ( .A1(n18550), .A2(n17119), .ZN(n17127) );
  OAI21_X1 U20125 ( .B1(n17120), .B2(n18429), .A(n17127), .ZN(n17122) );
  OAI211_X1 U20126 ( .C1(n17125), .C2(n18231), .A(n17124), .B(n17123), .ZN(
        P3_U2800) );
  INV_X1 U20127 ( .A(n17126), .ZN(n17129) );
  NAND2_X1 U20128 ( .A1(n17129), .A2(n18594), .ZN(n17162) );
  AOI21_X1 U20129 ( .B1(n17162), .B2(n17128), .A(n17127), .ZN(n17139) );
  AND2_X1 U20130 ( .A1(n18595), .A2(n17129), .ZN(n17160) );
  OAI211_X1 U20131 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n17160), .A(
        n18498), .B(n17130), .ZN(n17136) );
  AOI21_X1 U20132 ( .B1(n9963), .B2(n17296), .A(n9698), .ZN(n17328) );
  OAI21_X1 U20133 ( .B1(n17131), .B2(n18427), .A(n17328), .ZN(n17135) );
  OAI221_X1 U20134 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17133), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n19302), .A(n17132), .ZN(
        n17134) );
  NAND4_X1 U20135 ( .A1(n17137), .A2(n17136), .A3(n17135), .A4(n17134), .ZN(
        n17138) );
  NOR2_X1 U20136 ( .A1(n17139), .A2(n17138), .ZN(n17140) );
  OAI21_X1 U20137 ( .B1(n17141), .B2(n18471), .A(n17140), .ZN(P3_U2801) );
  OAI21_X1 U20138 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18816), .A(
        n17142), .ZN(n17147) );
  INV_X1 U20139 ( .A(n17143), .ZN(n18613) );
  NOR3_X1 U20140 ( .A1(n18613), .A2(n18887), .A3(n17144), .ZN(n17145) );
  AOI211_X1 U20141 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17147), .A(
        n17146), .B(n17145), .ZN(n17151) );
  AOI22_X1 U20142 ( .A1(n17149), .A2(n18823), .B1(n18901), .B2(n17148), .ZN(
        n17150) );
  OAI211_X1 U20143 ( .C1(n17152), .C2(n18799), .A(n17151), .B(n17150), .ZN(
        P3_U2831) );
  NAND4_X1 U20144 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18496), .A3(
        n9751), .A4(n18217), .ZN(n17165) );
  NAND2_X1 U20145 ( .A1(n19364), .A2(n18898), .ZN(n18906) );
  NOR3_X1 U20146 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n9988), .A3(
        n17153), .ZN(n18223) );
  NAND2_X1 U20147 ( .A1(n17155), .A2(n17154), .ZN(n18219) );
  AND2_X1 U20148 ( .A1(n19364), .A2(n17156), .ZN(n17157) );
  INV_X1 U20149 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19506) );
  NOR2_X1 U20150 ( .A1(n18890), .A2(n19506), .ZN(n18214) );
  NAND3_X1 U20151 ( .A1(n18822), .A2(n18227), .A3(n18219), .ZN(n17163) );
  OAI211_X1 U20152 ( .C1(n17165), .C2(n18906), .A(n17164), .B(n17163), .ZN(
        P3_U2834) );
  NOR3_X1 U20153 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17167) );
  NOR4_X1 U20154 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17166) );
  INV_X2 U20155 ( .A(n17258), .ZN(U215) );
  NAND4_X1 U20156 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17167), .A3(n17166), .A4(
        U215), .ZN(U213) );
  INV_X1 U20157 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n17260) );
  INV_X2 U20158 ( .A(U214), .ZN(n17221) );
  INV_X1 U20159 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17261) );
  OAI222_X1 U20160 ( .A1(U212), .A2(n17260), .B1(n17223), .B2(n17169), .C1(
        U214), .C2(n17261), .ZN(U216) );
  INV_X1 U20161 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n17171) );
  AOI22_X1 U20162 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n17220), .ZN(n17170) );
  OAI21_X1 U20163 ( .B1(n17171), .B2(n17223), .A(n17170), .ZN(U217) );
  INV_X1 U20164 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U20165 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17220), .ZN(n17172) );
  OAI21_X1 U20166 ( .B1(n17173), .B2(n17223), .A(n17172), .ZN(U218) );
  INV_X1 U20167 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20168 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17220), .ZN(n17174) );
  OAI21_X1 U20169 ( .B1(n17175), .B2(n17223), .A(n17174), .ZN(U219) );
  INV_X1 U20170 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n17177) );
  AOI22_X1 U20171 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17220), .ZN(n17176) );
  OAI21_X1 U20172 ( .B1(n17177), .B2(n17223), .A(n17176), .ZN(U220) );
  INV_X1 U20173 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20174 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17220), .ZN(n17178) );
  OAI21_X1 U20175 ( .B1(n17179), .B2(n17223), .A(n17178), .ZN(U221) );
  INV_X1 U20176 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U20177 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17220), .ZN(n17180) );
  OAI21_X1 U20178 ( .B1(n17181), .B2(n17223), .A(n17180), .ZN(U222) );
  INV_X1 U20179 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n21105) );
  AOI22_X1 U20180 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17220), .ZN(n17182) );
  OAI21_X1 U20181 ( .B1(n21105), .B2(n17223), .A(n17182), .ZN(U223) );
  INV_X1 U20182 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20183 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17220), .ZN(n17183) );
  OAI21_X1 U20184 ( .B1(n17184), .B2(n17223), .A(n17183), .ZN(U224) );
  INV_X1 U20185 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n21122) );
  AOI22_X1 U20186 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17220), .ZN(n17185) );
  OAI21_X1 U20187 ( .B1(n21122), .B2(n17223), .A(n17185), .ZN(U225) );
  INV_X1 U20188 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U20189 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17220), .ZN(n17186) );
  OAI21_X1 U20190 ( .B1(n17187), .B2(n17223), .A(n17186), .ZN(U226) );
  AOI22_X1 U20191 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17220), .ZN(n17188) );
  OAI21_X1 U20192 ( .B1(n17189), .B2(n17223), .A(n17188), .ZN(U227) );
  INV_X1 U20193 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U20194 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17220), .ZN(n17190) );
  OAI21_X1 U20195 ( .B1(n17191), .B2(n17223), .A(n17190), .ZN(U228) );
  AOI22_X1 U20196 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17220), .ZN(n17192) );
  OAI21_X1 U20197 ( .B1(n14786), .B2(n17223), .A(n17192), .ZN(U229) );
  INV_X1 U20198 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20199 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17220), .ZN(n17193) );
  OAI21_X1 U20200 ( .B1(n17194), .B2(n17223), .A(n17193), .ZN(U230) );
  AOI22_X1 U20201 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17220), .ZN(n17195) );
  OAI21_X1 U20202 ( .B1(n21081), .B2(n17223), .A(n17195), .ZN(U231) );
  AOI22_X1 U20203 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17220), .ZN(n17196) );
  OAI21_X1 U20204 ( .B1(n13221), .B2(n17223), .A(n17196), .ZN(U232) );
  AOI22_X1 U20205 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17220), .ZN(n17197) );
  OAI21_X1 U20206 ( .B1(n14732), .B2(n17223), .A(n17197), .ZN(U233) );
  AOI22_X1 U20207 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n17220), .ZN(n17198) );
  OAI21_X1 U20208 ( .B1(n14373), .B2(n17223), .A(n17198), .ZN(U234) );
  AOI22_X1 U20209 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17220), .ZN(n17199) );
  OAI21_X1 U20210 ( .B1(n17200), .B2(n17223), .A(n17199), .ZN(U235) );
  AOI22_X1 U20211 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n17220), .ZN(n17201) );
  OAI21_X1 U20212 ( .B1(n14147), .B2(n17223), .A(n17201), .ZN(U236) );
  AOI22_X1 U20213 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17220), .ZN(n17202) );
  OAI21_X1 U20214 ( .B1(n17203), .B2(n17223), .A(n17202), .ZN(U237) );
  AOI22_X1 U20215 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n17220), .ZN(n17204) );
  OAI21_X1 U20216 ( .B1(n12884), .B2(n17223), .A(n17204), .ZN(U238) );
  AOI22_X1 U20217 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17220), .ZN(n17205) );
  OAI21_X1 U20218 ( .B1(n12916), .B2(n17223), .A(n17205), .ZN(U239) );
  INV_X1 U20219 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n17207) );
  AOI22_X1 U20220 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n17220), .ZN(n17206) );
  OAI21_X1 U20221 ( .B1(n17207), .B2(n17223), .A(n17206), .ZN(U240) );
  AOI22_X1 U20222 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17220), .ZN(n17208) );
  OAI21_X1 U20223 ( .B1(n17209), .B2(n17223), .A(n17208), .ZN(U241) );
  INV_X1 U20224 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20225 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17220), .ZN(n17210) );
  OAI21_X1 U20226 ( .B1(n17211), .B2(n17223), .A(n17210), .ZN(U242) );
  AOI22_X1 U20227 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17220), .ZN(n17212) );
  OAI21_X1 U20228 ( .B1(n17213), .B2(n17223), .A(n17212), .ZN(U243) );
  INV_X1 U20229 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n17215) );
  AOI22_X1 U20230 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n17220), .ZN(n17214) );
  OAI21_X1 U20231 ( .B1(n17215), .B2(n17223), .A(n17214), .ZN(U244) );
  INV_X1 U20232 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20233 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17220), .ZN(n17216) );
  OAI21_X1 U20234 ( .B1(n17217), .B2(n17223), .A(n17216), .ZN(U245) );
  INV_X1 U20235 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n17219) );
  AOI22_X1 U20236 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17220), .ZN(n17218) );
  OAI21_X1 U20237 ( .B1(n17219), .B2(n17223), .A(n17218), .ZN(U246) );
  INV_X1 U20238 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20239 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n17221), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n17220), .ZN(n17222) );
  OAI21_X1 U20240 ( .B1(n17224), .B2(n17223), .A(n17222), .ZN(U247) );
  OAI22_X1 U20241 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n17258), .ZN(n17225) );
  INV_X1 U20242 ( .A(n17225), .ZN(U251) );
  OAI22_X1 U20243 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17258), .ZN(n17226) );
  INV_X1 U20244 ( .A(n17226), .ZN(U252) );
  OAI22_X1 U20245 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n17258), .ZN(n17227) );
  INV_X1 U20246 ( .A(n17227), .ZN(U253) );
  OAI22_X1 U20247 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n17258), .ZN(n17228) );
  INV_X1 U20248 ( .A(n17228), .ZN(U254) );
  OAI22_X1 U20249 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17258), .ZN(n17229) );
  INV_X1 U20250 ( .A(n17229), .ZN(U255) );
  OAI22_X1 U20251 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n17258), .ZN(n17230) );
  INV_X1 U20252 ( .A(n17230), .ZN(U256) );
  OAI22_X1 U20253 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n17258), .ZN(n17231) );
  INV_X1 U20254 ( .A(n17231), .ZN(U257) );
  OAI22_X1 U20255 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n17258), .ZN(n17232) );
  INV_X1 U20256 ( .A(n17232), .ZN(U258) );
  OAI22_X1 U20257 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17258), .ZN(n17233) );
  INV_X1 U20258 ( .A(n17233), .ZN(U259) );
  OAI22_X1 U20259 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n17252), .ZN(n17234) );
  INV_X1 U20260 ( .A(n17234), .ZN(U260) );
  OAI22_X1 U20261 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17252), .ZN(n17235) );
  INV_X1 U20262 ( .A(n17235), .ZN(U261) );
  OAI22_X1 U20263 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n17258), .ZN(n17236) );
  INV_X1 U20264 ( .A(n17236), .ZN(U262) );
  OAI22_X1 U20265 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n17258), .ZN(n17237) );
  INV_X1 U20266 ( .A(n17237), .ZN(U263) );
  OAI22_X1 U20267 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17258), .ZN(n17238) );
  INV_X1 U20268 ( .A(n17238), .ZN(U264) );
  OAI22_X1 U20269 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17258), .ZN(n17239) );
  INV_X1 U20270 ( .A(n17239), .ZN(U265) );
  OAI22_X1 U20271 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17252), .ZN(n17240) );
  INV_X1 U20272 ( .A(n17240), .ZN(U266) );
  OAI22_X1 U20273 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17252), .ZN(n17241) );
  INV_X1 U20274 ( .A(n17241), .ZN(U267) );
  OAI22_X1 U20275 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17252), .ZN(n17242) );
  INV_X1 U20276 ( .A(n17242), .ZN(U268) );
  OAI22_X1 U20277 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17252), .ZN(n17243) );
  INV_X1 U20278 ( .A(n17243), .ZN(U269) );
  OAI22_X1 U20279 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17252), .ZN(n17244) );
  INV_X1 U20280 ( .A(n17244), .ZN(U270) );
  OAI22_X1 U20281 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17252), .ZN(n17245) );
  INV_X1 U20282 ( .A(n17245), .ZN(U271) );
  OAI22_X1 U20283 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17258), .ZN(n17246) );
  INV_X1 U20284 ( .A(n17246), .ZN(U272) );
  OAI22_X1 U20285 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17258), .ZN(n17247) );
  INV_X1 U20286 ( .A(n17247), .ZN(U273) );
  OAI22_X1 U20287 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17252), .ZN(n17248) );
  INV_X1 U20288 ( .A(n17248), .ZN(U274) );
  OAI22_X1 U20289 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17258), .ZN(n17249) );
  INV_X1 U20290 ( .A(n17249), .ZN(U275) );
  OAI22_X1 U20291 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17258), .ZN(n17250) );
  INV_X1 U20292 ( .A(n17250), .ZN(U276) );
  OAI22_X1 U20293 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17258), .ZN(n17251) );
  INV_X1 U20294 ( .A(n17251), .ZN(U277) );
  OAI22_X1 U20295 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17252), .ZN(n17253) );
  INV_X1 U20296 ( .A(n17253), .ZN(U278) );
  OAI22_X1 U20297 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17258), .ZN(n17254) );
  INV_X1 U20298 ( .A(n17254), .ZN(U279) );
  OAI22_X1 U20299 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17258), .ZN(n17255) );
  INV_X1 U20300 ( .A(n17255), .ZN(U280) );
  OAI22_X1 U20301 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17258), .ZN(n17257) );
  INV_X1 U20302 ( .A(n17257), .ZN(U281) );
  INV_X1 U20303 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18948) );
  AOI22_X1 U20304 ( .A1(n17258), .A2(n17260), .B1(n18948), .B2(U215), .ZN(U282) );
  INV_X1 U20305 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17259) );
  AOI222_X1 U20306 ( .A1(n17261), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n17260), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17259), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17262) );
  INV_X2 U20307 ( .A(n17264), .ZN(n17263) );
  INV_X1 U20308 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19470) );
  INV_X1 U20309 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20527) );
  AOI22_X1 U20310 ( .A1(n17263), .A2(n19470), .B1(n20527), .B2(n17264), .ZN(
        U347) );
  INV_X1 U20311 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19468) );
  INV_X1 U20312 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20526) );
  AOI22_X1 U20313 ( .A1(n17263), .A2(n19468), .B1(n20526), .B2(n17264), .ZN(
        U348) );
  INV_X1 U20314 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19466) );
  INV_X1 U20315 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20525) );
  AOI22_X1 U20316 ( .A1(n17263), .A2(n19466), .B1(n20525), .B2(n17264), .ZN(
        U349) );
  INV_X1 U20317 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19464) );
  INV_X1 U20318 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20524) );
  AOI22_X1 U20319 ( .A1(n17263), .A2(n19464), .B1(n20524), .B2(n17264), .ZN(
        U350) );
  INV_X1 U20320 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19462) );
  INV_X1 U20321 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20523) );
  AOI22_X1 U20322 ( .A1(n17263), .A2(n19462), .B1(n20523), .B2(n17264), .ZN(
        U351) );
  INV_X1 U20323 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19460) );
  INV_X1 U20324 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n21125) );
  AOI22_X1 U20325 ( .A1(n17263), .A2(n19460), .B1(n21125), .B2(n17264), .ZN(
        U352) );
  INV_X1 U20326 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19458) );
  INV_X1 U20327 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20522) );
  AOI22_X1 U20328 ( .A1(n17263), .A2(n19458), .B1(n20522), .B2(n17264), .ZN(
        U353) );
  INV_X1 U20329 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19456) );
  AOI22_X1 U20330 ( .A1(n17263), .A2(n19456), .B1(n20521), .B2(n17264), .ZN(
        U354) );
  INV_X1 U20331 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19511) );
  INV_X1 U20332 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20558) );
  AOI22_X1 U20333 ( .A1(n17263), .A2(n19511), .B1(n20558), .B2(n17264), .ZN(
        U355) );
  INV_X1 U20334 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19507) );
  INV_X1 U20335 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20555) );
  AOI22_X1 U20336 ( .A1(n17263), .A2(n19507), .B1(n20555), .B2(n17264), .ZN(
        U356) );
  INV_X1 U20337 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19505) );
  INV_X1 U20338 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20553) );
  AOI22_X1 U20339 ( .A1(n17263), .A2(n19505), .B1(n20553), .B2(n17264), .ZN(
        U357) );
  INV_X1 U20340 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19504) );
  INV_X1 U20341 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20550) );
  AOI22_X1 U20342 ( .A1(n17263), .A2(n19504), .B1(n20550), .B2(n17264), .ZN(
        U358) );
  INV_X1 U20343 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19502) );
  INV_X1 U20344 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20549) );
  AOI22_X1 U20345 ( .A1(n17263), .A2(n19502), .B1(n20549), .B2(n17264), .ZN(
        U359) );
  INV_X1 U20346 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19500) );
  INV_X1 U20347 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20547) );
  AOI22_X1 U20348 ( .A1(n17263), .A2(n19500), .B1(n20547), .B2(n17264), .ZN(
        U360) );
  INV_X1 U20349 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19497) );
  INV_X1 U20350 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20545) );
  AOI22_X1 U20351 ( .A1(n17263), .A2(n19497), .B1(n20545), .B2(n17264), .ZN(
        U361) );
  INV_X1 U20352 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19495) );
  INV_X1 U20353 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20543) );
  AOI22_X1 U20354 ( .A1(n17263), .A2(n19495), .B1(n20543), .B2(n17264), .ZN(
        U362) );
  INV_X1 U20355 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19494) );
  INV_X1 U20356 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20541) );
  AOI22_X1 U20357 ( .A1(n17263), .A2(n19494), .B1(n20541), .B2(n17264), .ZN(
        U363) );
  INV_X1 U20358 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19492) );
  INV_X1 U20359 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n21202) );
  AOI22_X1 U20360 ( .A1(n17263), .A2(n19492), .B1(n21202), .B2(n17264), .ZN(
        U364) );
  INV_X1 U20361 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19454) );
  INV_X1 U20362 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20520) );
  AOI22_X1 U20363 ( .A1(n17263), .A2(n19454), .B1(n20520), .B2(n17264), .ZN(
        U365) );
  INV_X1 U20364 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19489) );
  INV_X1 U20365 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20539) );
  AOI22_X1 U20366 ( .A1(n17263), .A2(n19489), .B1(n20539), .B2(n17264), .ZN(
        U366) );
  INV_X1 U20367 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19488) );
  INV_X1 U20368 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20538) );
  AOI22_X1 U20369 ( .A1(n17263), .A2(n19488), .B1(n20538), .B2(n17264), .ZN(
        U367) );
  INV_X1 U20370 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19486) );
  INV_X1 U20371 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20536) );
  AOI22_X1 U20372 ( .A1(n17263), .A2(n19486), .B1(n20536), .B2(n17264), .ZN(
        U368) );
  INV_X1 U20373 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19483) );
  INV_X1 U20374 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20535) );
  AOI22_X1 U20375 ( .A1(n17263), .A2(n19483), .B1(n20535), .B2(n17264), .ZN(
        U369) );
  INV_X1 U20376 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19482) );
  INV_X1 U20377 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20533) );
  AOI22_X1 U20378 ( .A1(n17263), .A2(n19482), .B1(n20533), .B2(n17264), .ZN(
        U370) );
  INV_X1 U20379 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19480) );
  INV_X1 U20380 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20532) );
  AOI22_X1 U20381 ( .A1(n17263), .A2(n19480), .B1(n20532), .B2(n17264), .ZN(
        U371) );
  INV_X1 U20382 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19477) );
  INV_X1 U20383 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20531) );
  AOI22_X1 U20384 ( .A1(n17263), .A2(n19477), .B1(n20531), .B2(n17264), .ZN(
        U372) );
  INV_X1 U20385 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19476) );
  INV_X1 U20386 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20530) );
  AOI22_X1 U20387 ( .A1(n17263), .A2(n19476), .B1(n20530), .B2(n17264), .ZN(
        U373) );
  INV_X1 U20388 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19473) );
  INV_X1 U20389 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20529) );
  AOI22_X1 U20390 ( .A1(n17263), .A2(n19473), .B1(n20529), .B2(n17264), .ZN(
        U374) );
  INV_X1 U20391 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19472) );
  INV_X1 U20392 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20528) );
  AOI22_X1 U20393 ( .A1(n17263), .A2(n19472), .B1(n20528), .B2(n17264), .ZN(
        U375) );
  INV_X1 U20394 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19451) );
  INV_X1 U20395 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20518) );
  AOI22_X1 U20396 ( .A1(n17263), .A2(n19451), .B1(n20518), .B2(n17264), .ZN(
        U376) );
  INV_X1 U20397 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19450) );
  NAND2_X1 U20398 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19450), .ZN(n19436) );
  AOI22_X1 U20399 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19436), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19448), .ZN(n19521) );
  AOI21_X1 U20400 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19521), .ZN(n17265) );
  INV_X1 U20401 ( .A(n17265), .ZN(P3_U2633) );
  INV_X1 U20402 ( .A(n19424), .ZN(n17291) );
  OAI21_X1 U20403 ( .B1(n17273), .B2(n18101), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17266) );
  OAI21_X1 U20404 ( .B1(n17267), .B2(n17291), .A(n17266), .ZN(P3_U2634) );
  AOI21_X1 U20405 ( .B1(n19448), .B2(n19450), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17268) );
  AOI22_X1 U20406 ( .A1(n19584), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17268), 
        .B2(n19585), .ZN(P3_U2635) );
  NOR2_X1 U20407 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n17269) );
  OAI21_X1 U20408 ( .B1(n17269), .B2(BS16), .A(n19521), .ZN(n19519) );
  OAI21_X1 U20409 ( .B1(n19521), .B2(n21087), .A(n19519), .ZN(P3_U2636) );
  INV_X1 U20410 ( .A(n17270), .ZN(n17272) );
  NOR3_X1 U20411 ( .A1(n17273), .A2(n17272), .A3(n17271), .ZN(n19409) );
  NOR2_X1 U20412 ( .A1(n19409), .A2(n19413), .ZN(n19564) );
  OAI21_X1 U20413 ( .B1(n19564), .B2(n17275), .A(n17274), .ZN(P3_U2637) );
  NOR4_X1 U20414 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n17279) );
  NOR4_X1 U20415 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n17278) );
  NOR4_X1 U20416 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17277) );
  NOR4_X1 U20417 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17276) );
  NAND4_X1 U20418 ( .A1(n17279), .A2(n17278), .A3(n17277), .A4(n17276), .ZN(
        n17285) );
  NOR4_X1 U20419 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n17283) );
  AOI211_X1 U20420 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n17282) );
  NOR4_X1 U20421 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n17281) );
  NOR4_X1 U20422 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n17280) );
  NAND4_X1 U20423 ( .A1(n17283), .A2(n17282), .A3(n17281), .A4(n17280), .ZN(
        n17284) );
  NOR2_X1 U20424 ( .A1(n17285), .A2(n17284), .ZN(n19562) );
  INV_X1 U20425 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17287) );
  NOR3_X1 U20426 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17288) );
  OAI21_X1 U20427 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17288), .A(n19562), .ZN(
        n17286) );
  OAI21_X1 U20428 ( .B1(n19562), .B2(n17287), .A(n17286), .ZN(P3_U2638) );
  INV_X1 U20429 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19452) );
  INV_X1 U20430 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19520) );
  AOI21_X1 U20431 ( .B1(n19452), .B2(n19520), .A(n17288), .ZN(n17290) );
  INV_X1 U20432 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17289) );
  INV_X1 U20433 ( .A(n19562), .ZN(n19559) );
  AOI22_X1 U20434 ( .A1(n19562), .A2(n17290), .B1(n17289), .B2(n19559), .ZN(
        P3_U2639) );
  NOR2_X1 U20435 ( .A1(n19524), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19214) );
  INV_X1 U20436 ( .A(n19214), .ZN(n19422) );
  NOR2_X1 U20437 ( .A1(n17291), .A2(n19422), .ZN(n19418) );
  AOI211_X1 U20438 ( .C1(n18926), .C2(n19440), .A(P3_STATEBS16_REG_SCAN_IN), 
        .B(n19575), .ZN(n19414) );
  NAND2_X1 U20439 ( .A1(n19590), .A2(n18102), .ZN(n17295) );
  INV_X1 U20440 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19510) );
  INV_X1 U20441 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19503) );
  NOR2_X1 U20442 ( .A1(n19506), .A2(n19503), .ZN(n17337) );
  INV_X1 U20443 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19501) );
  INV_X1 U20444 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19499) );
  INV_X1 U20445 ( .A(n17295), .ZN(n17292) );
  INV_X1 U20446 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19493) );
  INV_X1 U20447 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19490) );
  INV_X1 U20448 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19474) );
  INV_X1 U20449 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19467) );
  INV_X1 U20450 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19465) );
  INV_X1 U20451 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19461) );
  INV_X1 U20452 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19455) );
  NAND2_X1 U20453 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17637) );
  NOR2_X1 U20454 ( .A1(n19455), .A2(n17637), .ZN(n17609) );
  NAND3_X1 U20455 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .A3(n17609), .ZN(n17588) );
  NOR2_X1 U20456 ( .A1(n19461), .A2(n17588), .ZN(n17575) );
  NAND2_X1 U20457 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17575), .ZN(n17562) );
  NOR3_X1 U20458 ( .A1(n19467), .A2(n19465), .A3(n17562), .ZN(n17536) );
  NAND3_X1 U20459 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(n17536), .ZN(n17510) );
  NOR2_X1 U20460 ( .A1(n19474), .A2(n17510), .ZN(n17501) );
  NAND3_X1 U20461 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n17501), .ZN(n17424) );
  NAND3_X1 U20462 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n17425) );
  NAND2_X1 U20463 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n17434) );
  NOR4_X1 U20464 ( .A1(n19490), .A2(n17424), .A3(n17425), .A4(n17434), .ZN(
        n17412) );
  NAND2_X1 U20465 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n17412), .ZN(n17396) );
  NOR2_X1 U20466 ( .A1(n19493), .A2(n17396), .ZN(n17387) );
  NAND2_X1 U20467 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17387), .ZN(n17307) );
  NOR2_X1 U20468 ( .A1(n17656), .A2(n17307), .ZN(n17306) );
  NAND2_X1 U20469 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17306), .ZN(n17369) );
  NOR3_X1 U20470 ( .A1(n19501), .A2(n19499), .A3(n17369), .ZN(n17351) );
  NAND3_X1 U20471 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17337), .A3(n17351), 
        .ZN(n17311) );
  NOR3_X1 U20472 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19510), .A3(n17311), 
        .ZN(n17293) );
  AOI21_X1 U20473 ( .B1(n17650), .B2(P3_EBX_REG_31__SCAN_IN), .A(n17293), .ZN(
        n17316) );
  NAND2_X1 U20474 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19574), .ZN(n17294) );
  AOI211_X4 U20475 ( .C1(n21087), .C2(n19568), .A(n17295), .B(n17294), .ZN(
        n17635) );
  NOR3_X1 U20476 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n17633) );
  INV_X1 U20477 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17628) );
  NAND2_X1 U20478 ( .A1(n17633), .A2(n17628), .ZN(n17627) );
  NOR2_X1 U20479 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17627), .ZN(n17604) );
  NAND2_X1 U20480 ( .A1(n17604), .A2(n17914), .ZN(n17600) );
  NAND2_X1 U20481 ( .A1(n17587), .A2(n17581), .ZN(n17580) );
  INV_X1 U20482 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17552) );
  NAND2_X1 U20483 ( .A1(n17561), .A2(n17552), .ZN(n17550) );
  INV_X1 U20484 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17530) );
  NAND2_X1 U20485 ( .A1(n17534), .A2(n17530), .ZN(n17529) );
  NAND2_X1 U20486 ( .A1(n17517), .A2(n17503), .ZN(n17502) );
  NAND2_X1 U20487 ( .A1(n17486), .A2(n17479), .ZN(n17478) );
  INV_X1 U20488 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17761) );
  NAND2_X1 U20489 ( .A1(n17461), .A2(n17761), .ZN(n17453) );
  NAND2_X1 U20490 ( .A1(n17442), .A2(n17431), .ZN(n17429) );
  INV_X1 U20491 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17671) );
  NAND2_X1 U20492 ( .A1(n17415), .A2(n17671), .ZN(n17408) );
  INV_X1 U20493 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17672) );
  NAND2_X1 U20494 ( .A1(n17398), .A2(n17672), .ZN(n17392) );
  INV_X1 U20495 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17673) );
  NAND2_X1 U20496 ( .A1(n17379), .A2(n17673), .ZN(n17372) );
  NOR2_X1 U20497 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17372), .ZN(n17360) );
  INV_X1 U20498 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17353) );
  NAND2_X1 U20499 ( .A1(n17360), .A2(n17353), .ZN(n17352) );
  NOR2_X1 U20500 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17352), .ZN(n17339) );
  INV_X1 U20501 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17676) );
  NAND2_X1 U20502 ( .A1(n17339), .A2(n17676), .ZN(n17318) );
  NOR2_X1 U20503 ( .A1(n17662), .A2(n17318), .ZN(n17323) );
  INV_X1 U20504 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17314) );
  NOR2_X1 U20505 ( .A1(n18581), .A2(n18209), .ZN(n17297) );
  OAI21_X1 U20506 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17297), .A(
        n17296), .ZN(n18226) );
  INV_X1 U20507 ( .A(n18226), .ZN(n17342) );
  INV_X1 U20508 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18238) );
  NAND2_X1 U20509 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18212), .ZN(
        n17298) );
  AOI21_X1 U20510 ( .B1(n18238), .B2(n17298), .A(n17297), .ZN(n18232) );
  NOR2_X1 U20511 ( .A1(n18581), .A2(n18283), .ZN(n18280) );
  INV_X1 U20512 ( .A(n18280), .ZN(n17302) );
  NOR2_X1 U20513 ( .A1(n18254), .A2(n17302), .ZN(n17301) );
  INV_X1 U20514 ( .A(n17301), .ZN(n17300) );
  NOR3_X1 U20515 ( .A1(n9951), .A2(n9952), .A3(n17300), .ZN(n18210) );
  OAI21_X1 U20516 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18210), .A(
        n17298), .ZN(n18244) );
  INV_X1 U20517 ( .A(n18244), .ZN(n17359) );
  NAND2_X1 U20518 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17301), .ZN(
        n17299) );
  AOI21_X1 U20519 ( .B1(n9952), .B2(n17299), .A(n18210), .ZN(n18257) );
  AOI22_X1 U20520 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17301), .B1(
        n17300), .B2(n9951), .ZN(n18270) );
  AOI21_X1 U20521 ( .B1(n18254), .B2(n17302), .A(n17301), .ZN(n18281) );
  INV_X1 U20522 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18302) );
  NOR2_X1 U20523 ( .A1(n18581), .A2(n18336), .ZN(n18335) );
  INV_X1 U20524 ( .A(n18335), .ZN(n17449) );
  NOR2_X1 U20525 ( .A1(n17303), .A2(n17449), .ZN(n17305) );
  NAND2_X1 U20526 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17305), .ZN(
        n17304) );
  AOI21_X1 U20527 ( .B1(n18302), .B2(n17304), .A(n18280), .ZN(n18304) );
  INV_X1 U20528 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18310) );
  XNOR2_X1 U20529 ( .A(n18310), .B(n17305), .ZN(n18313) );
  INV_X1 U20530 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18298) );
  NAND2_X1 U20531 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18335), .ZN(
        n17438) );
  INV_X1 U20532 ( .A(n17438), .ZN(n17426) );
  NAND2_X1 U20533 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17426), .ZN(
        n18296) );
  AOI21_X1 U20534 ( .B1(n18298), .B2(n18296), .A(n17305), .ZN(n18330) );
  INV_X1 U20535 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17456) );
  NAND2_X1 U20536 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18337) );
  NOR2_X1 U20537 ( .A1(n17456), .A2(n18337), .ZN(n18329) );
  NOR2_X1 U20538 ( .A1(n18581), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17644) );
  NAND2_X1 U20539 ( .A1(n18327), .A2(n17644), .ZN(n17439) );
  INV_X1 U20540 ( .A(n17439), .ZN(n17450) );
  AOI21_X1 U20541 ( .B1(n18329), .B2(n17450), .A(n17619), .ZN(n17418) );
  NOR2_X1 U20542 ( .A1(n18330), .A2(n17418), .ZN(n17417) );
  NOR2_X1 U20543 ( .A1(n17417), .A2(n17619), .ZN(n17407) );
  NOR2_X1 U20544 ( .A1(n18281), .A2(n17386), .ZN(n17385) );
  NOR2_X1 U20545 ( .A1(n17385), .A2(n17619), .ZN(n17378) );
  NOR2_X1 U20546 ( .A1(n18270), .A2(n17378), .ZN(n17377) );
  NOR2_X1 U20547 ( .A1(n17377), .A2(n17619), .ZN(n17368) );
  NOR2_X1 U20548 ( .A1(n18257), .A2(n17368), .ZN(n17367) );
  NOR2_X1 U20549 ( .A1(n17367), .A2(n17619), .ZN(n17358) );
  NOR2_X1 U20550 ( .A1(n17359), .A2(n17358), .ZN(n17357) );
  NOR2_X1 U20551 ( .A1(n17357), .A2(n17619), .ZN(n17348) );
  NOR2_X1 U20552 ( .A1(n18232), .A2(n17348), .ZN(n17347) );
  NOR2_X1 U20553 ( .A1(n17347), .A2(n17619), .ZN(n17341) );
  NOR2_X1 U20554 ( .A1(n17342), .A2(n17341), .ZN(n17340) );
  NOR2_X1 U20555 ( .A1(n17340), .A2(n17619), .ZN(n17327) );
  INV_X1 U20556 ( .A(n17651), .ZN(n19428) );
  NAND2_X1 U20557 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17337), .ZN(n17310) );
  INV_X1 U20558 ( .A(n17649), .ZN(n17666) );
  NAND2_X1 U20559 ( .A1(n17666), .A2(n17656), .ZN(n17664) );
  INV_X1 U20560 ( .A(n17664), .ZN(n17309) );
  NOR2_X1 U20561 ( .A1(n19501), .A2(n19499), .ZN(n17308) );
  INV_X1 U20562 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19498) );
  AND2_X1 U20563 ( .A1(n19498), .A2(n17306), .ZN(n17376) );
  NAND2_X1 U20564 ( .A1(n17638), .A2(n17307), .ZN(n17388) );
  NAND2_X1 U20565 ( .A1(n17666), .A2(n17388), .ZN(n17384) );
  NOR2_X1 U20566 ( .A1(n17376), .A2(n17384), .ZN(n17375) );
  OAI21_X1 U20567 ( .B1(n17309), .B2(n17308), .A(n17375), .ZN(n17364) );
  AOI21_X1 U20568 ( .B1(n17638), .B2(n17310), .A(n17364), .ZN(n17336) );
  NOR2_X1 U20569 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17311), .ZN(n17321) );
  INV_X1 U20570 ( .A(n17321), .ZN(n17312) );
  AOI21_X1 U20571 ( .B1(n17336), .B2(n17312), .A(n19512), .ZN(n17313) );
  OAI211_X1 U20572 ( .C1(n17317), .C2(n17652), .A(n17316), .B(n17315), .ZN(
        P3_U2640) );
  NAND2_X1 U20573 ( .A1(n17635), .A2(n17318), .ZN(n17332) );
  XOR2_X1 U20574 ( .A(n17319), .B(n9631), .Z(n17322) );
  OAI22_X1 U20575 ( .A1(n17336), .A2(n19510), .B1(n9964), .B2(n17652), .ZN(
        n17320) );
  AOI211_X1 U20576 ( .C1(n17322), .C2(n17651), .A(n17321), .B(n17320), .ZN(
        n17325) );
  OAI21_X1 U20577 ( .B1(n17650), .B2(n17323), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17324) );
  OAI211_X1 U20578 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17332), .A(n17325), .B(
        n17324), .ZN(P3_U2641) );
  INV_X1 U20579 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19508) );
  AOI211_X1 U20580 ( .C1(n17328), .C2(n17327), .A(n17326), .B(n19428), .ZN(
        n17331) );
  NAND2_X1 U20581 ( .A1(n17337), .A2(n17351), .ZN(n17329) );
  OAI22_X1 U20582 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17329), .B1(n9963), 
        .B2(n17652), .ZN(n17330) );
  AOI211_X1 U20583 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17608), .A(n17331), .B(
        n17330), .ZN(n17335) );
  INV_X1 U20584 ( .A(n17332), .ZN(n17333) );
  OAI21_X1 U20585 ( .B1(n17339), .B2(n17676), .A(n17333), .ZN(n17334) );
  OAI211_X1 U20586 ( .C1(n17336), .C2(n19508), .A(n17335), .B(n17334), .ZN(
        P3_U2642) );
  AOI21_X1 U20587 ( .B1(n19506), .B2(n19503), .A(n17337), .ZN(n17338) );
  AOI22_X1 U20588 ( .A1(n17650), .A2(P3_EBX_REG_28__SCAN_IN), .B1(n17351), 
        .B2(n17338), .ZN(n17346) );
  AOI211_X1 U20589 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17352), .A(n17339), .B(
        n17662), .ZN(n17344) );
  AOI211_X1 U20590 ( .C1(n17342), .C2(n17341), .A(n17340), .B(n19428), .ZN(
        n17343) );
  AOI211_X1 U20591 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17364), .A(n17344), 
        .B(n17343), .ZN(n17345) );
  OAI211_X1 U20592 ( .C1(n18213), .C2(n17652), .A(n17346), .B(n17345), .ZN(
        P3_U2643) );
  INV_X1 U20593 ( .A(n17364), .ZN(n17356) );
  AOI211_X1 U20594 ( .C1(n18232), .C2(n17348), .A(n17347), .B(n19428), .ZN(
        n17350) );
  OAI22_X1 U20595 ( .A1(n18238), .A2(n17652), .B1(n17663), .B2(n17353), .ZN(
        n17349) );
  AOI211_X1 U20596 ( .C1(n17351), .C2(n19503), .A(n17350), .B(n17349), .ZN(
        n17355) );
  OAI211_X1 U20597 ( .C1(n17360), .C2(n17353), .A(n17635), .B(n17352), .ZN(
        n17354) );
  OAI211_X1 U20598 ( .C1(n17356), .C2(n19503), .A(n17355), .B(n17354), .ZN(
        P3_U2644) );
  OAI21_X1 U20599 ( .B1(n19499), .B2(n17369), .A(n19501), .ZN(n17363) );
  AOI211_X1 U20600 ( .C1(n17359), .C2(n17358), .A(n17357), .B(n19428), .ZN(
        n17362) );
  AOI211_X1 U20601 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17372), .A(n17360), .B(
        n17662), .ZN(n17361) );
  AOI211_X1 U20602 ( .C1(n17364), .C2(n17363), .A(n17362), .B(n17361), .ZN(
        n17366) );
  NAND2_X1 U20603 ( .A1(n17650), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n17365) );
  OAI211_X1 U20604 ( .C1(n17652), .C2(n18242), .A(n17366), .B(n17365), .ZN(
        P3_U2645) );
  AOI211_X1 U20605 ( .C1(n18257), .C2(n17368), .A(n17367), .B(n19428), .ZN(
        n17371) );
  OAI22_X1 U20606 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17369), .B1(n9952), 
        .B2(n17652), .ZN(n17370) );
  AOI211_X1 U20607 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n17608), .A(n17371), .B(
        n17370), .ZN(n17374) );
  OAI211_X1 U20608 ( .C1(n17379), .C2(n17673), .A(n17635), .B(n17372), .ZN(
        n17373) );
  OAI211_X1 U20609 ( .C1(n17375), .C2(n19499), .A(n17374), .B(n17373), .ZN(
        P3_U2646) );
  AOI21_X1 U20610 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17650), .A(n17376), .ZN(
        n17383) );
  AOI211_X1 U20611 ( .C1(n18270), .C2(n17378), .A(n17377), .B(n19428), .ZN(
        n17381) );
  AOI211_X1 U20612 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17392), .A(n17379), .B(
        n17662), .ZN(n17380) );
  AOI211_X1 U20613 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n17384), .A(n17381), 
        .B(n17380), .ZN(n17382) );
  OAI211_X1 U20614 ( .C1(n9951), .C2(n17652), .A(n17383), .B(n17382), .ZN(
        P3_U2647) );
  INV_X1 U20615 ( .A(n17384), .ZN(n17395) );
  INV_X1 U20616 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19496) );
  AOI211_X1 U20617 ( .C1(n18281), .C2(n17386), .A(n17385), .B(n19428), .ZN(
        n17391) );
  INV_X1 U20618 ( .A(n17387), .ZN(n17389) );
  OAI22_X1 U20619 ( .A1(n18254), .A2(n17652), .B1(n17389), .B2(n17388), .ZN(
        n17390) );
  AOI211_X1 U20620 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n17608), .A(n17391), .B(
        n17390), .ZN(n17394) );
  OAI211_X1 U20621 ( .C1(n17398), .C2(n17672), .A(n17635), .B(n17392), .ZN(
        n17393) );
  OAI211_X1 U20622 ( .C1(n17395), .C2(n19496), .A(n17394), .B(n17393), .ZN(
        P3_U2648) );
  NOR3_X1 U20623 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17656), .A3(n17396), 
        .ZN(n17397) );
  AOI21_X1 U20624 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17650), .A(n17397), .ZN(
        n17405) );
  OAI221_X1 U20625 ( .B1(n17656), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n17656), 
        .C2(n17412), .A(n17666), .ZN(n17403) );
  AOI211_X1 U20626 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17408), .A(n17398), .B(
        n17662), .ZN(n17402) );
  AOI211_X1 U20627 ( .C1(n18304), .C2(n17400), .A(n17399), .B(n19428), .ZN(
        n17401) );
  AOI211_X1 U20628 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17403), .A(n17402), 
        .B(n17401), .ZN(n17404) );
  OAI211_X1 U20629 ( .C1(n18302), .C2(n17652), .A(n17405), .B(n17404), .ZN(
        P3_U2649) );
  OAI21_X1 U20630 ( .B1(n17412), .B2(n17656), .A(n17666), .ZN(n17421) );
  AOI211_X1 U20631 ( .C1(n18313), .C2(n17407), .A(n17406), .B(n19428), .ZN(
        n17411) );
  OAI211_X1 U20632 ( .C1(n17415), .C2(n17671), .A(n17635), .B(n17408), .ZN(
        n17409) );
  OAI21_X1 U20633 ( .B1(n17652), .B2(n18310), .A(n17409), .ZN(n17410) );
  AOI211_X1 U20634 ( .C1(n17421), .C2(P3_REIP_REG_21__SCAN_IN), .A(n17411), 
        .B(n17410), .ZN(n17414) );
  INV_X1 U20635 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19491) );
  NAND3_X1 U20636 ( .A1(n17638), .A2(n17412), .A3(n19491), .ZN(n17413) );
  OAI211_X1 U20637 ( .C1(n17671), .C2(n17663), .A(n17414), .B(n17413), .ZN(
        P3_U2650) );
  AOI211_X1 U20638 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17429), .A(n17415), .B(
        n17662), .ZN(n17416) );
  AOI21_X1 U20639 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17650), .A(n17416), .ZN(
        n17423) );
  NOR2_X1 U20640 ( .A1(n17656), .A2(n17424), .ZN(n17463) );
  INV_X1 U20641 ( .A(n17463), .ZN(n17481) );
  NOR2_X1 U20642 ( .A1(n17425), .A2(n17481), .ZN(n17435) );
  INV_X1 U20643 ( .A(n17435), .ZN(n17448) );
  NOR2_X1 U20644 ( .A1(n17434), .A2(n17448), .ZN(n17420) );
  AOI211_X1 U20645 ( .C1(n18330), .C2(n17418), .A(n17417), .B(n19428), .ZN(
        n17419) );
  AOI221_X1 U20646 ( .B1(n17421), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n17420), 
        .C2(n19490), .A(n17419), .ZN(n17422) );
  OAI211_X1 U20647 ( .C1(n18298), .C2(n17652), .A(n17423), .B(n17422), .ZN(
        P3_U2651) );
  OR2_X1 U20648 ( .A1(n17424), .A2(n17649), .ZN(n17487) );
  OAI21_X1 U20649 ( .B1(n17425), .B2(n17487), .A(n17664), .ZN(n17460) );
  INV_X1 U20650 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19487) );
  INV_X1 U20651 ( .A(n17644), .ZN(n17541) );
  NOR2_X1 U20652 ( .A1(n18376), .A2(n17541), .ZN(n17475) );
  AOI21_X1 U20653 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17475), .A(
        n17619), .ZN(n17472) );
  AOI21_X1 U20654 ( .B1(n17655), .B2(n17438), .A(n17472), .ZN(n17428) );
  OAI21_X1 U20655 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17426), .A(
        n18296), .ZN(n18340) );
  OAI21_X1 U20656 ( .B1(n17428), .B2(n18340), .A(n17651), .ZN(n17427) );
  AOI21_X1 U20657 ( .B1(n17428), .B2(n18340), .A(n17427), .ZN(n17433) );
  OAI211_X1 U20658 ( .C1(n17442), .C2(n17431), .A(n17635), .B(n17429), .ZN(
        n17430) );
  OAI211_X1 U20659 ( .C1(n17663), .C2(n17431), .A(n18890), .B(n17430), .ZN(
        n17432) );
  AOI211_X1 U20660 ( .C1(n17564), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n17433), .B(n17432), .ZN(n17437) );
  OAI211_X1 U20661 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n17435), .B(n17434), .ZN(n17436) );
  OAI211_X1 U20662 ( .C1(n17460), .C2(n19487), .A(n17437), .B(n17436), .ZN(
        P3_U2652) );
  INV_X1 U20663 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19485) );
  OAI21_X1 U20664 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18335), .A(
        n17438), .ZN(n18350) );
  OAI21_X1 U20665 ( .B1(n17456), .B2(n17439), .A(n17655), .ZN(n17441) );
  OAI21_X1 U20666 ( .B1(n18350), .B2(n17441), .A(n17651), .ZN(n17440) );
  AOI21_X1 U20667 ( .B1(n18350), .B2(n17441), .A(n17440), .ZN(n17446) );
  AOI211_X1 U20668 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17453), .A(n17442), .B(
        n17662), .ZN(n17445) );
  AOI22_X1 U20669 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17564), .B1(
        n17650), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n17443) );
  INV_X1 U20670 ( .A(n17443), .ZN(n17444) );
  NOR4_X1 U20671 ( .A1(n18902), .A2(n17446), .A3(n17445), .A4(n17444), .ZN(
        n17447) );
  OAI221_X1 U20672 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17448), .C1(n19485), 
        .C2(n17460), .A(n17447), .ZN(P3_U2653) );
  INV_X1 U20673 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19484) );
  NOR2_X1 U20674 ( .A1(n18581), .A2(n18376), .ZN(n17476) );
  INV_X1 U20675 ( .A(n17476), .ZN(n18377) );
  NOR2_X1 U20676 ( .A1(n18381), .A2(n18377), .ZN(n17468) );
  OAI21_X1 U20677 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17468), .A(
        n17449), .ZN(n18367) );
  NOR2_X1 U20678 ( .A1(n17450), .A2(n17619), .ZN(n17451) );
  XNOR2_X1 U20679 ( .A(n18367), .B(n17451), .ZN(n17458) );
  NAND2_X1 U20680 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17462) );
  NOR3_X1 U20681 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17462), .A3(n17481), 
        .ZN(n17452) );
  AOI211_X1 U20682 ( .C1(n17650), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18902), .B(
        n17452), .ZN(n17455) );
  OAI211_X1 U20683 ( .C1(n17461), .C2(n17761), .A(n17635), .B(n17453), .ZN(
        n17454) );
  OAI211_X1 U20684 ( .C1(n17652), .C2(n17456), .A(n17455), .B(n17454), .ZN(
        n17457) );
  AOI21_X1 U20685 ( .B1(n17458), .B2(n17651), .A(n17457), .ZN(n17459) );
  OAI21_X1 U20686 ( .B1(n19484), .B2(n17460), .A(n17459), .ZN(P3_U2654) );
  NAND2_X1 U20687 ( .A1(n17664), .A2(n17487), .ZN(n17499) );
  INV_X1 U20688 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19481) );
  AOI211_X1 U20689 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17478), .A(n17461), .B(
        n17662), .ZN(n17467) );
  INV_X1 U20690 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17465) );
  OAI211_X1 U20691 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n17463), .B(n17462), .ZN(n17464) );
  OAI211_X1 U20692 ( .C1(n17663), .C2(n17465), .A(n18890), .B(n17464), .ZN(
        n17466) );
  AOI211_X1 U20693 ( .C1(n17564), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17467), .B(n17466), .ZN(n17474) );
  INV_X1 U20694 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18385) );
  NAND2_X1 U20695 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17476), .ZN(
        n17469) );
  AOI21_X1 U20696 ( .B1(n18385), .B2(n17469), .A(n17468), .ZN(n18383) );
  INV_X1 U20697 ( .A(n18383), .ZN(n17471) );
  INV_X1 U20698 ( .A(n17472), .ZN(n17470) );
  OAI221_X1 U20699 ( .B1(n18383), .B2(n17472), .C1(n17471), .C2(n17470), .A(
        n17651), .ZN(n17473) );
  OAI211_X1 U20700 ( .C1(n17499), .C2(n19481), .A(n17474), .B(n17473), .ZN(
        P3_U2655) );
  INV_X1 U20701 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19479) );
  AOI22_X1 U20702 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17564), .B1(
        n17650), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n17485) );
  NOR2_X1 U20703 ( .A1(n17475), .A2(n17619), .ZN(n17477) );
  INV_X1 U20704 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18391) );
  AOI22_X1 U20705 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17476), .B1(
        n18377), .B2(n18391), .ZN(n18394) );
  XOR2_X1 U20706 ( .A(n17477), .B(n18394), .Z(n17483) );
  OAI211_X1 U20707 ( .C1(n17486), .C2(n17479), .A(n17635), .B(n17478), .ZN(
        n17480) );
  OAI211_X1 U20708 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n17481), .A(n18890), 
        .B(n17480), .ZN(n17482) );
  AOI21_X1 U20709 ( .B1(n17483), .B2(n17651), .A(n17482), .ZN(n17484) );
  OAI211_X1 U20710 ( .C1(n19479), .C2(n17499), .A(n17485), .B(n17484), .ZN(
        P3_U2656) );
  INV_X1 U20711 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19478) );
  AOI211_X1 U20712 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17502), .A(n17486), .B(
        n17662), .ZN(n17491) );
  INV_X1 U20713 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17489) );
  NAND4_X1 U20714 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17638), .A3(n17501), 
        .A4(n17487), .ZN(n17488) );
  OAI211_X1 U20715 ( .C1(n17489), .C2(n17652), .A(n18890), .B(n17488), .ZN(
        n17490) );
  AOI211_X1 U20716 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17608), .A(n17491), .B(
        n17490), .ZN(n17498) );
  INV_X1 U20717 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18424) );
  NAND2_X1 U20718 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17493) );
  NOR2_X1 U20719 ( .A1(n18581), .A2(n18487), .ZN(n17571) );
  INV_X1 U20720 ( .A(n17571), .ZN(n17559) );
  NOR2_X1 U20721 ( .A1(n17492), .A2(n17559), .ZN(n17540) );
  INV_X1 U20722 ( .A(n17540), .ZN(n17547) );
  NOR2_X1 U20723 ( .A1(n17493), .A2(n17547), .ZN(n18417) );
  NAND2_X1 U20724 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18417), .ZN(
        n17513) );
  NOR2_X1 U20725 ( .A1(n18424), .A2(n17513), .ZN(n17500) );
  OAI21_X1 U20726 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17500), .A(
        n18377), .ZN(n18410) );
  INV_X1 U20727 ( .A(n18408), .ZN(n17494) );
  OAI21_X1 U20728 ( .B1(n17494), .B2(n17541), .A(n17655), .ZN(n17496) );
  AOI21_X1 U20729 ( .B1(n18410), .B2(n17496), .A(n19428), .ZN(n17495) );
  OAI21_X1 U20730 ( .B1(n18410), .B2(n17496), .A(n17495), .ZN(n17497) );
  OAI211_X1 U20731 ( .C1(n17499), .C2(n19478), .A(n17498), .B(n17497), .ZN(
        P3_U2657) );
  AOI21_X1 U20732 ( .B1(n18424), .B2(n17513), .A(n17500), .ZN(n18426) );
  OAI21_X1 U20733 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17513), .A(
        n17655), .ZN(n17516) );
  XOR2_X1 U20734 ( .A(n18426), .B(n17516), .Z(n17509) );
  AOI22_X1 U20735 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17564), .B1(
        n17650), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n17508) );
  NOR2_X1 U20736 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17656), .ZN(n17511) );
  AOI21_X1 U20737 ( .B1(n17510), .B2(n17638), .A(n17649), .ZN(n17527) );
  INV_X1 U20738 ( .A(n17527), .ZN(n17520) );
  NAND2_X1 U20739 ( .A1(n17638), .A2(n17501), .ZN(n17505) );
  OAI211_X1 U20740 ( .C1(n17517), .C2(n17503), .A(n17635), .B(n17502), .ZN(
        n17504) );
  OAI211_X1 U20741 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17505), .A(n18890), 
        .B(n17504), .ZN(n17506) );
  AOI221_X1 U20742 ( .B1(n17511), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n17520), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n17506), .ZN(n17507) );
  OAI211_X1 U20743 ( .C1(n19428), .C2(n17509), .A(n17508), .B(n17507), .ZN(
        P3_U2658) );
  INV_X1 U20744 ( .A(n17510), .ZN(n17512) );
  AOI22_X1 U20745 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17564), .B1(
        n17512), .B2(n17511), .ZN(n17523) );
  OAI21_X1 U20746 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18417), .A(
        n17513), .ZN(n18435) );
  NAND2_X1 U20747 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17540), .ZN(
        n17539) );
  NOR2_X1 U20748 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17539), .ZN(
        n17514) );
  AOI211_X1 U20749 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17514), .A(
        n17619), .B(n18435), .ZN(n17515) );
  AOI211_X1 U20750 ( .C1(n18435), .C2(n17516), .A(n17515), .B(n19428), .ZN(
        n17519) );
  AOI211_X1 U20751 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17529), .A(n17517), .B(
        n17662), .ZN(n17518) );
  AOI211_X1 U20752 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17650), .A(n17519), .B(
        n17518), .ZN(n17522) );
  NAND2_X1 U20753 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17520), .ZN(n17521) );
  NAND4_X1 U20754 ( .A1(n17523), .A2(n17522), .A3(n18890), .A4(n17521), .ZN(
        P3_U2659) );
  INV_X1 U20755 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17533) );
  AND2_X1 U20756 ( .A1(n17638), .A2(n17536), .ZN(n17538) );
  AOI21_X1 U20757 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n17538), .A(
        P3_REIP_REG_11__SCAN_IN), .ZN(n17526) );
  AOI21_X1 U20758 ( .B1(n17533), .B2(n17539), .A(n18417), .ZN(n18453) );
  OAI21_X1 U20759 ( .B1(n17539), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n17655), .ZN(n17524) );
  INV_X1 U20760 ( .A(n17524), .ZN(n17543) );
  XNOR2_X1 U20761 ( .A(n18453), .B(n17543), .ZN(n17525) );
  OAI22_X1 U20762 ( .A1(n17527), .A2(n17526), .B1(n19428), .B2(n17525), .ZN(
        n17528) );
  AOI211_X1 U20763 ( .C1(n17650), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18902), .B(
        n17528), .ZN(n17532) );
  OAI211_X1 U20764 ( .C1(n17534), .C2(n17530), .A(n17635), .B(n17529), .ZN(
        n17531) );
  OAI211_X1 U20765 ( .C1(n17652), .C2(n17533), .A(n17532), .B(n17531), .ZN(
        P3_U2660) );
  AOI211_X1 U20766 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17550), .A(n17534), .B(
        n17662), .ZN(n17535) );
  AOI21_X1 U20767 ( .B1(n17564), .B2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17535), .ZN(n17546) );
  OAI21_X1 U20768 ( .B1(n17536), .B2(n17656), .A(n17666), .ZN(n17555) );
  INV_X1 U20769 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19469) );
  OAI21_X1 U20770 ( .B1(n17663), .B2(n17860), .A(n18890), .ZN(n17537) );
  AOI221_X1 U20771 ( .B1(n17555), .B2(P3_REIP_REG_10__SCAN_IN), .C1(n17538), 
        .C2(n19469), .A(n17537), .ZN(n17545) );
  OAI21_X1 U20772 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17540), .A(
        n17539), .ZN(n17542) );
  INV_X1 U20773 ( .A(n17542), .ZN(n18468) );
  INV_X1 U20774 ( .A(n18449), .ZN(n18461) );
  OAI21_X1 U20775 ( .B1(n18461), .B2(n17541), .A(n17655), .ZN(n17548) );
  OAI221_X1 U20776 ( .B1(n18468), .B2(n17543), .C1(n17542), .C2(n17548), .A(
        n17651), .ZN(n17544) );
  NAND3_X1 U20777 ( .A1(n17546), .A2(n17545), .A3(n17544), .ZN(P3_U2661) );
  NAND2_X1 U20778 ( .A1(n17651), .A2(n17619), .ZN(n17647) );
  INV_X1 U20779 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18486) );
  NOR2_X1 U20780 ( .A1(n18486), .A2(n17559), .ZN(n17558) );
  OAI21_X1 U20781 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17558), .A(
        n17547), .ZN(n18475) );
  NOR2_X1 U20782 ( .A1(n9956), .A2(n18486), .ZN(n18485) );
  AND2_X1 U20783 ( .A1(n18488), .A2(n17644), .ZN(n17572) );
  AOI21_X1 U20784 ( .B1(n18485), .B2(n17572), .A(n18475), .ZN(n17549) );
  NOR3_X1 U20785 ( .A1(n17549), .A2(n17548), .A3(n19428), .ZN(n17554) );
  OAI211_X1 U20786 ( .C1(n17561), .C2(n17552), .A(n17635), .B(n17550), .ZN(
        n17551) );
  OAI211_X1 U20787 ( .C1(n17663), .C2(n17552), .A(n18890), .B(n17551), .ZN(
        n17553) );
  AOI211_X1 U20788 ( .C1(n17564), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17554), .B(n17553), .ZN(n17557) );
  NOR2_X1 U20789 ( .A1(n17656), .A2(n17562), .ZN(n17563) );
  OAI221_X1 U20790 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(P3_REIP_REG_8__SCAN_IN), 
        .C1(P3_REIP_REG_9__SCAN_IN), .C2(n17563), .A(n17555), .ZN(n17556) );
  OAI211_X1 U20791 ( .C1(n17647), .C2(n18475), .A(n17557), .B(n17556), .ZN(
        P3_U2662) );
  AOI21_X1 U20792 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17572), .A(
        n17619), .ZN(n17560) );
  AOI21_X1 U20793 ( .B1(n18486), .B2(n17559), .A(n17558), .ZN(n18493) );
  XNOR2_X1 U20794 ( .A(n17560), .B(n18493), .ZN(n17569) );
  AOI211_X1 U20795 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17580), .A(n17561), .B(
        n17662), .ZN(n17567) );
  AOI21_X1 U20796 ( .B1(n17638), .B2(n17562), .A(n17649), .ZN(n17570) );
  AOI22_X1 U20797 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17564), .B1(
        n17563), .B2(n19465), .ZN(n17565) );
  OAI211_X1 U20798 ( .C1(n19465), .C2(n17570), .A(n17565), .B(n18890), .ZN(
        n17566) );
  AOI211_X1 U20799 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17650), .A(n17567), .B(
        n17566), .ZN(n17568) );
  OAI21_X1 U20800 ( .B1(n19428), .B2(n17569), .A(n17568), .ZN(P3_U2663) );
  INV_X1 U20801 ( .A(n17570), .ZN(n17579) );
  NOR2_X1 U20802 ( .A1(n18581), .A2(n18517), .ZN(n17595) );
  NAND2_X1 U20803 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17595), .ZN(
        n17584) );
  AOI21_X1 U20804 ( .B1(n9956), .B2(n17584), .A(n17571), .ZN(n18509) );
  NOR2_X1 U20805 ( .A1(n17572), .A2(n17619), .ZN(n17574) );
  INV_X1 U20806 ( .A(n18509), .ZN(n17573) );
  INV_X1 U20807 ( .A(n17574), .ZN(n17586) );
  AOI221_X1 U20808 ( .B1(n18509), .B2(n17574), .C1(n17573), .C2(n17586), .A(
        n19428), .ZN(n17578) );
  INV_X1 U20809 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19463) );
  NAND3_X1 U20810 ( .A1(n17638), .A2(n17575), .A3(n19463), .ZN(n17576) );
  OAI211_X1 U20811 ( .C1(n17663), .C2(n17581), .A(n18890), .B(n17576), .ZN(
        n17577) );
  AOI211_X1 U20812 ( .C1(n17579), .C2(P3_REIP_REG_7__SCAN_IN), .A(n17578), .B(
        n17577), .ZN(n17583) );
  OAI211_X1 U20813 ( .C1(n17587), .C2(n17581), .A(n17635), .B(n17580), .ZN(
        n17582) );
  OAI211_X1 U20814 ( .C1(n17652), .C2(n9956), .A(n17583), .B(n17582), .ZN(
        P3_U2664) );
  INV_X1 U20815 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17654) );
  OAI221_X1 U20816 ( .B1(n17619), .B2(n17595), .C1(n17619), .C2(n17654), .A(
        n17651), .ZN(n17594) );
  OAI21_X1 U20817 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17595), .A(
        n17584), .ZN(n18523) );
  NOR3_X1 U20818 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17656), .A3(n17588), .ZN(
        n17585) );
  AOI211_X1 U20819 ( .C1(n17650), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18902), .B(
        n17585), .ZN(n17593) );
  NOR2_X1 U20820 ( .A1(n19428), .A2(n17586), .ZN(n17591) );
  AOI211_X1 U20821 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17600), .A(n17587), .B(
        n17662), .ZN(n17590) );
  AOI21_X1 U20822 ( .B1(n17638), .B2(n17588), .A(n17649), .ZN(n17597) );
  OAI22_X1 U20823 ( .A1(n18520), .A2(n17652), .B1(n19461), .B2(n17597), .ZN(
        n17589) );
  AOI211_X1 U20824 ( .C1(n17591), .C2(n18523), .A(n17590), .B(n17589), .ZN(
        n17592) );
  OAI211_X1 U20825 ( .C1(n17594), .C2(n18523), .A(n17593), .B(n17592), .ZN(
        P3_U2665) );
  INV_X1 U20826 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17603) );
  NOR3_X1 U20827 ( .A1(n17656), .A2(n19455), .A3(n17637), .ZN(n17615) );
  AOI21_X1 U20828 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17615), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17598) );
  NAND2_X1 U20829 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18527), .ZN(
        n17611) );
  AOI21_X1 U20830 ( .B1(n17603), .B2(n17611), .A(n17595), .ZN(n18535) );
  OAI21_X1 U20831 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17611), .A(
        n17655), .ZN(n17610) );
  XOR2_X1 U20832 ( .A(n18535), .B(n17610), .Z(n17596) );
  OAI22_X1 U20833 ( .A1(n17598), .A2(n17597), .B1(n19428), .B2(n17596), .ZN(
        n17599) );
  AOI211_X1 U20834 ( .C1(n17650), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18902), .B(
        n17599), .ZN(n17602) );
  OAI211_X1 U20835 ( .C1(n17604), .C2(n17914), .A(n17635), .B(n17600), .ZN(
        n17601) );
  OAI211_X1 U20836 ( .C1(n17652), .C2(n17603), .A(n17602), .B(n17601), .ZN(
        P3_U2666) );
  AOI211_X1 U20837 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17627), .A(n17604), .B(
        n17662), .ZN(n17607) );
  NAND2_X1 U20838 ( .A1(n18923), .A2(n19590), .ZN(n17669) );
  OAI221_X1 U20839 ( .B1(n17669), .B2(n17790), .C1(n17669), .C2(n17605), .A(
        n18890), .ZN(n17606) );
  AOI211_X1 U20840 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17608), .A(n17607), .B(
        n17606), .ZN(n17617) );
  OAI21_X1 U20841 ( .B1(n17609), .B2(n17656), .A(n17666), .ZN(n17626) );
  INV_X1 U20842 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19457) );
  NOR2_X1 U20843 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18545), .ZN(
        n18540) );
  INV_X1 U20844 ( .A(n17610), .ZN(n17612) );
  NOR2_X1 U20845 ( .A1(n18581), .A2(n18545), .ZN(n17618) );
  OAI21_X1 U20846 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17618), .A(
        n17611), .ZN(n18548) );
  AOI22_X1 U20847 ( .A1(n17644), .A2(n18540), .B1(n17612), .B2(n18548), .ZN(
        n17613) );
  OAI22_X1 U20848 ( .A1(n17613), .A2(n19428), .B1(n18548), .B2(n17647), .ZN(
        n17614) );
  AOI221_X1 U20849 ( .B1(n17626), .B2(P3_REIP_REG_4__SCAN_IN), .C1(n17615), 
        .C2(n19457), .A(n17614), .ZN(n17616) );
  OAI211_X1 U20850 ( .C1(n18547), .C2(n17652), .A(n17617), .B(n17616), .ZN(
        P3_U2667) );
  INV_X1 U20851 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17631) );
  OAI21_X1 U20852 ( .B1(n17656), .B2(n17637), .A(n19455), .ZN(n17625) );
  NAND2_X1 U20853 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17632) );
  AOI21_X1 U20854 ( .B1(n17631), .B2(n17632), .A(n17618), .ZN(n18562) );
  INV_X1 U20855 ( .A(n17632), .ZN(n17620) );
  AOI21_X1 U20856 ( .B1(n17620), .B2(n17654), .A(n17619), .ZN(n17643) );
  OAI21_X1 U20857 ( .B1(n18562), .B2(n17643), .A(n17651), .ZN(n17621) );
  AOI21_X1 U20858 ( .B1(n18562), .B2(n17643), .A(n17621), .ZN(n17624) );
  INV_X1 U20859 ( .A(n17669), .ZN(n19592) );
  OR2_X1 U20860 ( .A1(n19554), .A2(n19391), .ZN(n19370) );
  AOI21_X1 U20861 ( .B1(n19531), .B2(n19370), .A(n14232), .ZN(n19529) );
  AOI22_X1 U20862 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17650), .B1(n19592), .B2(
        n19529), .ZN(n17622) );
  INV_X1 U20863 ( .A(n17622), .ZN(n17623) );
  AOI211_X1 U20864 ( .C1(n17626), .C2(n17625), .A(n17624), .B(n17623), .ZN(
        n17630) );
  OAI211_X1 U20865 ( .C1(n17633), .C2(n17628), .A(n17635), .B(n17627), .ZN(
        n17629) );
  OAI211_X1 U20866 ( .C1(n17652), .C2(n17631), .A(n17630), .B(n17629), .ZN(
        P3_U2668) );
  OAI21_X1 U20867 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17632), .ZN(n18570) );
  INV_X1 U20868 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17930) );
  INV_X1 U20869 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18574) );
  OAI22_X1 U20870 ( .A1(n17930), .A2(n17663), .B1(n18574), .B2(n17652), .ZN(
        n17642) );
  OAI21_X1 U20871 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n19372), .A(
        n19370), .ZN(n19390) );
  NOR2_X1 U20872 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17636) );
  INV_X1 U20873 ( .A(n17633), .ZN(n17634) );
  OAI211_X1 U20874 ( .C1(n17636), .C2(n17930), .A(n17635), .B(n17634), .ZN(
        n17640) );
  OAI211_X1 U20875 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17638), .B(n17637), .ZN(n17639) );
  OAI211_X1 U20876 ( .C1(n17669), .C2(n19390), .A(n17640), .B(n17639), .ZN(
        n17641) );
  AOI211_X1 U20877 ( .C1(n17649), .C2(P3_REIP_REG_2__SCAN_IN), .A(n17642), .B(
        n17641), .ZN(n17646) );
  OAI211_X1 U20878 ( .C1(n17644), .C2(n18570), .A(n17651), .B(n17643), .ZN(
        n17645) );
  OAI211_X1 U20879 ( .C1(n17647), .C2(n18570), .A(n17646), .B(n17645), .ZN(
        P3_U2669) );
  NAND2_X1 U20880 ( .A1(n19394), .A2(n17648), .ZN(n19542) );
  AOI22_X1 U20881 ( .A1(n17650), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n17649), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17661) );
  NAND2_X1 U20882 ( .A1(n17655), .A2(n17651), .ZN(n17653) );
  OAI21_X1 U20883 ( .B1(n17654), .B2(n17653), .A(n17652), .ZN(n17659) );
  AOI21_X1 U20884 ( .B1(n17655), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n19428), .ZN(n17658) );
  NAND2_X1 U20885 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17931) );
  OAI21_X1 U20886 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17931), .ZN(n17940) );
  OAI22_X1 U20887 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17656), .B1(n17662), 
        .B2(n17940), .ZN(n17657) );
  AOI221_X1 U20888 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17659), .C1(
        n18581), .C2(n17658), .A(n17657), .ZN(n17660) );
  OAI211_X1 U20889 ( .C1(n19542), .C2(n17669), .A(n17661), .B(n17660), .ZN(
        P3_U2670) );
  NAND2_X1 U20890 ( .A1(n17663), .A2(n17662), .ZN(n17665) );
  AOI22_X1 U20891 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17665), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17664), .ZN(n17668) );
  NAND3_X1 U20892 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19526), .A3(
        n17666), .ZN(n17667) );
  OAI211_X1 U20893 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17669), .A(
        n17668), .B(n17667), .ZN(P3_U2671) );
  NAND2_X1 U20894 ( .A1(n18954), .A2(n17670), .ZN(n17677) );
  INV_X1 U20895 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17745) );
  NAND2_X1 U20896 ( .A1(n18954), .A2(n17744), .ZN(n17731) );
  NOR3_X2 U20897 ( .A1(n17671), .A2(n17745), .A3(n17731), .ZN(n17706) );
  NAND2_X1 U20898 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17706), .ZN(n17700) );
  NOR2_X2 U20899 ( .A1(n17672), .A2(n17700), .ZN(n17705) );
  NAND2_X1 U20900 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17705), .ZN(n17691) );
  NAND2_X1 U20901 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17696), .ZN(n17687) );
  OAI21_X1 U20902 ( .B1(n17687), .B2(n17674), .A(n17935), .ZN(n17680) );
  OAI211_X1 U20903 ( .C1(n17960), .C2(n17959), .A(n17942), .B(n17958), .ZN(
        n17675) );
  OAI221_X1 U20904 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n17677), .C1(n17676), 
        .C2(n17680), .A(n17675), .ZN(P3_U2674) );
  INV_X1 U20905 ( .A(n17687), .ZN(n17690) );
  NAND2_X1 U20906 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17690), .ZN(n17682) );
  INV_X1 U20907 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17681) );
  AOI21_X1 U20908 ( .B1(n17678), .B2(n17683), .A(n17960), .ZN(n17965) );
  NAND2_X1 U20909 ( .A1(n17942), .A2(n17965), .ZN(n17679) );
  OAI221_X1 U20910 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17682), .C1(n17681), 
        .C2(n17680), .A(n17679), .ZN(P3_U2675) );
  OAI21_X1 U20911 ( .B1(n17685), .B2(n17684), .A(n17683), .ZN(n17974) );
  NAND3_X1 U20912 ( .A1(n17687), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17935), 
        .ZN(n17686) );
  OAI221_X1 U20913 ( .B1(n17687), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17935), 
        .C2(n17974), .A(n17686), .ZN(P3_U2676) );
  AOI21_X1 U20914 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17935), .A(n17696), .ZN(
        n17689) );
  XNOR2_X1 U20915 ( .A(n17688), .B(n17692), .ZN(n17979) );
  OAI22_X1 U20916 ( .A1(n17690), .A2(n17689), .B1(n17935), .B2(n17979), .ZN(
        P3_U2677) );
  INV_X1 U20917 ( .A(n17691), .ZN(n17699) );
  AOI21_X1 U20918 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17935), .A(n17699), .ZN(
        n17695) );
  OAI21_X1 U20919 ( .B1(n17694), .B2(n17693), .A(n17692), .ZN(n17984) );
  OAI22_X1 U20920 ( .A1(n17696), .A2(n17695), .B1(n17935), .B2(n17984), .ZN(
        P3_U2678) );
  AOI21_X1 U20921 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17935), .A(n17705), .ZN(
        n17698) );
  XNOR2_X1 U20922 ( .A(n17697), .B(n17701), .ZN(n17989) );
  OAI22_X1 U20923 ( .A1(n17699), .A2(n17698), .B1(n17935), .B2(n17989), .ZN(
        P3_U2679) );
  INV_X1 U20924 ( .A(n17700), .ZN(n17720) );
  AOI21_X1 U20925 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17935), .A(n17720), .ZN(
        n17704) );
  OAI21_X1 U20926 ( .B1(n17703), .B2(n17702), .A(n17701), .ZN(n17994) );
  OAI22_X1 U20927 ( .A1(n17705), .A2(n17704), .B1(n17935), .B2(n17994), .ZN(
        P3_U2680) );
  AOI21_X1 U20928 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17935), .A(n17706), .ZN(
        n17719) );
  AOI22_X1 U20929 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17717) );
  AOI22_X1 U20930 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17716) );
  AOI22_X1 U20931 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17707) );
  OAI21_X1 U20932 ( .B1(n21139), .B2(n17708), .A(n17707), .ZN(n17714) );
  AOI22_X1 U20933 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17712) );
  AOI22_X1 U20934 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17711) );
  AOI22_X1 U20935 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n9595), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17710) );
  AOI22_X1 U20936 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n17895), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17709) );
  NAND4_X1 U20937 ( .A1(n17712), .A2(n17711), .A3(n17710), .A4(n17709), .ZN(
        n17713) );
  AOI211_X1 U20938 ( .C1(n17816), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n17714), .B(n17713), .ZN(n17715) );
  NAND3_X1 U20939 ( .A1(n17717), .A2(n17716), .A3(n17715), .ZN(n17995) );
  INV_X1 U20940 ( .A(n17995), .ZN(n17718) );
  OAI22_X1 U20941 ( .A1(n17720), .A2(n17719), .B1(n17718), .B2(n17935), .ZN(
        P3_U2681) );
  AOI22_X1 U20942 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17724) );
  AOI22_X1 U20943 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17723) );
  AOI22_X1 U20944 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17722) );
  AOI22_X1 U20945 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17721) );
  NAND4_X1 U20946 ( .A1(n17724), .A2(n17723), .A3(n17722), .A4(n17721), .ZN(
        n17730) );
  AOI22_X1 U20947 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17728) );
  AOI22_X1 U20948 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n17895), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17727) );
  AOI22_X1 U20949 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17726) );
  AOI22_X1 U20950 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17725) );
  NAND4_X1 U20951 ( .A1(n17728), .A2(n17727), .A3(n17726), .A4(n17725), .ZN(
        n17729) );
  NOR2_X1 U20952 ( .A1(n17730), .A2(n17729), .ZN(n18003) );
  INV_X1 U20953 ( .A(n17731), .ZN(n17746) );
  OAI221_X1 U20954 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(P3_EBX_REG_20__SCAN_IN), 
        .C1(P3_EBX_REG_21__SCAN_IN), .C2(n17746), .A(n17732), .ZN(n17733) );
  AOI22_X1 U20955 ( .A1(n17942), .A2(n18003), .B1(n17733), .B2(n17935), .ZN(
        P3_U2682) );
  AOI22_X1 U20956 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17737) );
  AOI22_X1 U20957 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17736) );
  AOI22_X1 U20958 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16334), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17735) );
  AOI22_X1 U20959 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17734) );
  NAND4_X1 U20960 ( .A1(n17737), .A2(n17736), .A3(n17735), .A4(n17734), .ZN(
        n17743) );
  AOI22_X1 U20961 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17741) );
  AOI22_X1 U20962 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17740) );
  AOI22_X1 U20963 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17739) );
  AOI22_X1 U20964 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17738) );
  NAND4_X1 U20965 ( .A1(n17741), .A2(n17740), .A3(n17739), .A4(n17738), .ZN(
        n17742) );
  NOR2_X1 U20966 ( .A1(n17743), .A2(n17742), .ZN(n18007) );
  NOR2_X1 U20967 ( .A1(n17942), .A2(n17744), .ZN(n17759) );
  AOI22_X1 U20968 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17759), .B1(n17746), 
        .B2(n17745), .ZN(n17747) );
  OAI21_X1 U20969 ( .B1(n18007), .B2(n17935), .A(n17747), .ZN(P3_U2683) );
  AOI22_X1 U20970 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n17903), .B1(
        n17862), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U20971 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17750) );
  AOI22_X1 U20972 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U20973 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17748) );
  NAND4_X1 U20974 ( .A1(n17751), .A2(n17750), .A3(n17749), .A4(n17748), .ZN(
        n17757) );
  AOI22_X1 U20975 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17755) );
  AOI22_X1 U20976 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17754) );
  AOI22_X1 U20977 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n17877), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17753) );
  AOI22_X1 U20978 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17752) );
  NAND4_X1 U20979 ( .A1(n17755), .A2(n17754), .A3(n17753), .A4(n17752), .ZN(
        n17756) );
  NOR2_X1 U20980 ( .A1(n17757), .A2(n17756), .ZN(n18012) );
  INV_X1 U20981 ( .A(n17758), .ZN(n17775) );
  OAI21_X1 U20982 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17775), .A(n17759), .ZN(
        n17760) );
  OAI21_X1 U20983 ( .B1(n18012), .B2(n17935), .A(n17760), .ZN(P3_U2684) );
  NAND3_X1 U20984 ( .A1(n18954), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17788), 
        .ZN(n17787) );
  NOR2_X1 U20985 ( .A1(n17761), .A2(n17787), .ZN(n17762) );
  AOI21_X1 U20986 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17935), .A(n17762), .ZN(
        n17774) );
  AOI22_X1 U20987 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17767) );
  AOI22_X1 U20988 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17766) );
  AOI22_X1 U20989 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17765) );
  AOI22_X1 U20990 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17764) );
  NAND4_X1 U20991 ( .A1(n17767), .A2(n17766), .A3(n17765), .A4(n17764), .ZN(
        n17773) );
  AOI22_X1 U20992 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17771) );
  AOI22_X1 U20993 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n17882), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17770) );
  AOI22_X1 U20994 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17769) );
  AOI22_X1 U20995 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n17876), .B1(
        n16368), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17768) );
  NAND4_X1 U20996 ( .A1(n17771), .A2(n17770), .A3(n17769), .A4(n17768), .ZN(
        n17772) );
  NOR2_X1 U20997 ( .A1(n17773), .A2(n17772), .ZN(n18017) );
  OAI22_X1 U20998 ( .A1(n17775), .A2(n17774), .B1(n18017), .B2(n17935), .ZN(
        P3_U2685) );
  AOI22_X1 U20999 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14232), .B1(
        n17862), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17779) );
  AOI22_X1 U21000 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17778) );
  AOI22_X1 U21001 ( .A1(n17894), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17777) );
  AOI22_X1 U21002 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17776) );
  NAND4_X1 U21003 ( .A1(n17779), .A2(n17778), .A3(n17777), .A4(n17776), .ZN(
        n17785) );
  AOI22_X1 U21004 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17783) );
  AOI22_X1 U21005 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17782) );
  AOI22_X1 U21006 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17781) );
  AOI22_X1 U21007 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17780) );
  NAND4_X1 U21008 ( .A1(n17783), .A2(n17782), .A3(n17781), .A4(n17780), .ZN(
        n17784) );
  NOR2_X1 U21009 ( .A1(n17785), .A2(n17784), .ZN(n18023) );
  NAND3_X1 U21010 ( .A1(n17787), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n17935), 
        .ZN(n17786) );
  OAI221_X1 U21011 ( .B1(n17787), .B2(P3_EBX_REG_17__SCAN_IN), .C1(n17935), 
        .C2(n18023), .A(n17786), .ZN(P3_U2686) );
  NAND2_X1 U21012 ( .A1(n18954), .A2(n17788), .ZN(n17801) );
  NOR2_X1 U21013 ( .A1(n17942), .A2(n17788), .ZN(n17813) );
  AOI22_X1 U21014 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17799) );
  AOI22_X1 U21015 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17798) );
  AOI22_X1 U21016 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17789) );
  OAI21_X1 U21017 ( .B1(n21156), .B2(n17790), .A(n17789), .ZN(n17796) );
  AOI22_X1 U21018 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17794) );
  AOI22_X1 U21019 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17793) );
  AOI22_X1 U21020 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17903), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17792) );
  AOI22_X1 U21021 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17791) );
  NAND4_X1 U21022 ( .A1(n17794), .A2(n17793), .A3(n17792), .A4(n17791), .ZN(
        n17795) );
  AOI211_X1 U21023 ( .C1(n17893), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n17796), .B(n17795), .ZN(n17797) );
  NAND3_X1 U21024 ( .A1(n17799), .A2(n17798), .A3(n17797), .ZN(n18024) );
  AOI22_X1 U21025 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17813), .B1(n17942), 
        .B2(n18024), .ZN(n17800) );
  OAI21_X1 U21026 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17801), .A(n17800), .ZN(
        P3_U2687) );
  AOI22_X1 U21027 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17805) );
  AOI22_X1 U21028 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14232), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17877), .ZN(n17804) );
  AOI22_X1 U21029 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17876), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17803) );
  AOI22_X1 U21030 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17802) );
  NAND4_X1 U21031 ( .A1(n17805), .A2(n17804), .A3(n17803), .A4(n17802), .ZN(
        n17811) );
  AOI22_X1 U21032 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17809) );
  AOI22_X1 U21033 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17901), .B1(
        n17903), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17808) );
  AOI22_X1 U21034 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17892), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17902), .ZN(n17807) );
  AOI22_X1 U21035 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17895), .ZN(n17806) );
  NAND4_X1 U21036 ( .A1(n17809), .A2(n17808), .A3(n17807), .A4(n17806), .ZN(
        n17810) );
  NOR2_X1 U21037 ( .A1(n17811), .A2(n17810), .ZN(n18033) );
  INV_X1 U21038 ( .A(n17812), .ZN(n17814) );
  OAI21_X1 U21039 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17814), .A(n17813), .ZN(
        n17815) );
  OAI21_X1 U21040 ( .B1(n18033), .B2(n17935), .A(n17815), .ZN(P3_U2688) );
  AOI22_X1 U21041 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17820) );
  AOI22_X1 U21042 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17819) );
  AOI22_X1 U21043 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n17816), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17818) );
  AOI22_X1 U21044 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17817) );
  NAND4_X1 U21045 ( .A1(n17820), .A2(n17819), .A3(n17818), .A4(n17817), .ZN(
        n17827) );
  AOI22_X1 U21046 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17825) );
  AOI22_X1 U21047 ( .A1(n17821), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17824) );
  AOI22_X1 U21048 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n17900), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17823) );
  AOI22_X1 U21049 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n17902), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17822) );
  NAND4_X1 U21050 ( .A1(n17825), .A2(n17824), .A3(n17823), .A4(n17822), .ZN(
        n17826) );
  NOR2_X1 U21051 ( .A1(n17827), .A2(n17826), .ZN(n18038) );
  NOR2_X1 U21052 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18087), .ZN(n17828) );
  AOI22_X1 U21053 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17830), .B1(n17829), 
        .B2(n17828), .ZN(n17831) );
  OAI21_X1 U21054 ( .B1(n18038), .B2(n17935), .A(n17831), .ZN(P3_U2689) );
  AOI22_X1 U21055 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17835) );
  AOI22_X1 U21056 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17834) );
  AOI22_X1 U21057 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17833) );
  AOI22_X1 U21058 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17832) );
  NAND4_X1 U21059 ( .A1(n17835), .A2(n17834), .A3(n17833), .A4(n17832), .ZN(
        n17841) );
  AOI22_X1 U21060 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17839) );
  AOI22_X1 U21061 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17838) );
  AOI22_X1 U21062 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17837) );
  AOI22_X1 U21063 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17836) );
  NAND4_X1 U21064 ( .A1(n17839), .A2(n17838), .A3(n17837), .A4(n17836), .ZN(
        n17840) );
  NOR2_X1 U21065 ( .A1(n17841), .A2(n17840), .ZN(n18044) );
  OAI21_X1 U21066 ( .B1(n18087), .B2(n17857), .A(n17842), .ZN(n17843) );
  INV_X1 U21067 ( .A(n17843), .ZN(n17844) );
  OAI22_X1 U21068 ( .A1(n18044), .A2(n17935), .B1(n17845), .B2(n17844), .ZN(
        P3_U2691) );
  AOI22_X1 U21069 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17856) );
  AOI22_X1 U21070 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n17883), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17855) );
  INV_X1 U21071 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21084) );
  AOI22_X1 U21072 ( .A1(n17894), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17846) );
  OAI21_X1 U21073 ( .B1(n21084), .B2(n17847), .A(n17846), .ZN(n17853) );
  AOI22_X1 U21074 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17851) );
  AOI22_X1 U21075 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17850) );
  AOI22_X1 U21076 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17849) );
  AOI22_X1 U21077 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17903), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17848) );
  NAND4_X1 U21078 ( .A1(n17851), .A2(n17850), .A3(n17849), .A4(n17848), .ZN(
        n17852) );
  AOI211_X1 U21079 ( .C1(n17900), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n17853), .B(n17852), .ZN(n17854) );
  NAND3_X1 U21080 ( .A1(n17856), .A2(n17855), .A3(n17854), .ZN(n18048) );
  INV_X1 U21081 ( .A(n18048), .ZN(n17859) );
  OAI211_X1 U21082 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n17874), .A(n17857), .B(
        n17935), .ZN(n17858) );
  OAI21_X1 U21083 ( .B1(n17859), .B2(n17935), .A(n17858), .ZN(P3_U2692) );
  AOI21_X1 U21084 ( .B1(n17860), .B2(n17890), .A(n17942), .ZN(n17861) );
  INV_X1 U21085 ( .A(n17861), .ZN(n17873) );
  AOI22_X1 U21086 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17895), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17866) );
  AOI22_X1 U21087 ( .A1(n17882), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17865) );
  AOI22_X1 U21088 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n17877), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17864) );
  AOI22_X1 U21089 ( .A1(n17862), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17863) );
  NAND4_X1 U21090 ( .A1(n17866), .A2(n17865), .A3(n17864), .A4(n17863), .ZN(
        n17872) );
  AOI22_X1 U21091 ( .A1(n17892), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17870) );
  AOI22_X1 U21092 ( .A1(n17883), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17869) );
  AOI22_X1 U21093 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n9595), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17868) );
  AOI22_X1 U21094 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17903), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17867) );
  NAND4_X1 U21095 ( .A1(n17870), .A2(n17869), .A3(n17868), .A4(n17867), .ZN(
        n17871) );
  NOR2_X1 U21096 ( .A1(n17872), .A2(n17871), .ZN(n18052) );
  OAI22_X1 U21097 ( .A1(n17874), .A2(n17873), .B1(n18052), .B2(n17935), .ZN(
        P3_U2693) );
  AOI22_X1 U21098 ( .A1(n17876), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17881) );
  AOI22_X1 U21099 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17877), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17880) );
  AOI22_X1 U21100 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17879) );
  AOI22_X1 U21101 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17878) );
  NAND4_X1 U21102 ( .A1(n17881), .A2(n17880), .A3(n17879), .A4(n17878), .ZN(
        n17889) );
  AOI22_X1 U21103 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17887) );
  AOI22_X1 U21104 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17886) );
  AOI22_X1 U21105 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17885) );
  AOI22_X1 U21106 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17862), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17884) );
  NAND4_X1 U21107 ( .A1(n17887), .A2(n17886), .A3(n17885), .A4(n17884), .ZN(
        n17888) );
  NOR2_X1 U21108 ( .A1(n17889), .A2(n17888), .ZN(n18057) );
  OAI21_X1 U21109 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17911), .A(n17890), .ZN(
        n17891) );
  AOI22_X1 U21110 ( .A1(n17942), .A2(n18057), .B1(n17891), .B2(n17935), .ZN(
        P3_U2694) );
  OAI21_X1 U21111 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17917), .A(n17935), .ZN(
        n17910) );
  AOI22_X1 U21112 ( .A1(n17893), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17892), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17899) );
  AOI22_X1 U21113 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n17862), .B1(
        n17821), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17898) );
  AOI22_X1 U21114 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17882), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17897) );
  AOI22_X1 U21115 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17894), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17896) );
  NAND4_X1 U21116 ( .A1(n17899), .A2(n17898), .A3(n17897), .A4(n17896), .ZN(
        n17909) );
  AOI22_X1 U21117 ( .A1(n17900), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17883), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17907) );
  AOI22_X1 U21118 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17906) );
  AOI22_X1 U21119 ( .A1(n16368), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17876), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17905) );
  AOI22_X1 U21120 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17902), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17904) );
  NAND4_X1 U21121 ( .A1(n17907), .A2(n17906), .A3(n17905), .A4(n17904), .ZN(
        n17908) );
  NOR2_X1 U21122 ( .A1(n17909), .A2(n17908), .ZN(n18065) );
  OAI22_X1 U21123 ( .A1(n17911), .A2(n17910), .B1(n18065), .B2(n17935), .ZN(
        P3_U2695) );
  NAND2_X1 U21124 ( .A1(n18954), .A2(n17938), .ZN(n17944) );
  NOR2_X1 U21125 ( .A1(n17912), .A2(n17944), .ZN(n17932) );
  NAND2_X1 U21126 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17932), .ZN(n17926) );
  NOR3_X1 U21127 ( .A1(n17914), .A2(n17913), .A3(n17926), .ZN(n17923) );
  AND2_X1 U21128 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17923), .ZN(n17920) );
  AOI21_X1 U21129 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17935), .A(n17920), .ZN(
        n17916) );
  INV_X1 U21130 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17915) );
  OAI22_X1 U21131 ( .A1(n17917), .A2(n17916), .B1(n17915), .B2(n17935), .ZN(
        P3_U2696) );
  AOI21_X1 U21132 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17935), .A(n17923), .ZN(
        n17919) );
  INV_X1 U21133 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17918) );
  OAI22_X1 U21134 ( .A1(n17920), .A2(n17919), .B1(n17918), .B2(n17935), .ZN(
        P3_U2697) );
  INV_X1 U21135 ( .A(n17926), .ZN(n17929) );
  AOI22_X1 U21136 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17935), .B1(
        P3_EBX_REG_4__SCAN_IN), .B2(n17929), .ZN(n17922) );
  OAI22_X1 U21137 ( .A1(n17923), .A2(n17922), .B1(n17921), .B2(n17935), .ZN(
        P3_U2698) );
  NAND3_X1 U21138 ( .A1(n17926), .A2(P3_EBX_REG_4__SCAN_IN), .A3(n17935), .ZN(
        n17924) );
  OAI221_X1 U21139 ( .B1(n17926), .B2(P3_EBX_REG_4__SCAN_IN), .C1(n17935), 
        .C2(n17925), .A(n17924), .ZN(P3_U2699) );
  AOI21_X1 U21140 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17935), .A(n17932), .ZN(
        n17928) );
  INV_X1 U21141 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17927) );
  OAI22_X1 U21142 ( .A1(n17929), .A2(n17928), .B1(n17927), .B2(n17935), .ZN(
        P3_U2700) );
  OAI221_X1 U21143 ( .B1(n17931), .B2(n17941), .C1(n18954), .C2(n17941), .A(
        n17930), .ZN(n17934) );
  INV_X1 U21144 ( .A(n17932), .ZN(n17933) );
  OAI211_X1 U21145 ( .C1(n17935), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17934), .B(n17933), .ZN(n17936) );
  INV_X1 U21146 ( .A(n17936), .ZN(P3_U2701) );
  INV_X1 U21147 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17939) );
  OAI222_X1 U21148 ( .A1(n17944), .A2(n17940), .B1(n17939), .B2(n17938), .C1(
        n17937), .C2(n17935), .ZN(P3_U2702) );
  AOI22_X1 U21149 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17942), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17941), .ZN(n17943) );
  OAI21_X1 U21150 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17944), .A(n17943), .ZN(
        P3_U2703) );
  INV_X1 U21151 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18167) );
  INV_X1 U21152 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18163) );
  INV_X1 U21153 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18208) );
  NAND2_X1 U21154 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n18066) );
  NAND3_X1 U21155 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .ZN(n18067) );
  NAND3_X1 U21156 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(n17946), .ZN(n18062) );
  NAND4_X1 U21157 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17947)
         );
  NOR2_X1 U21158 ( .A1(n18062), .A2(n17947), .ZN(n17948) );
  NAND4_X1 U21159 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .A4(n17948), .ZN(n18035) );
  INV_X1 U21160 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18155) );
  INV_X1 U21161 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18153) );
  NAND4_X1 U21162 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17949)
         );
  NAND2_X1 U21163 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17991), .ZN(n17990) );
  NAND2_X1 U21164 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17986), .ZN(n17985) );
  NAND2_X1 U21165 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17967), .ZN(n17961) );
  NAND2_X1 U21166 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17954), .ZN(n17953) );
  NAND2_X1 U21167 ( .A1(n17953), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n17952) );
  NOR2_X2 U21168 ( .A1(n18945), .A2(n18095), .ZN(n18025) );
  NAND2_X1 U21169 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18025), .ZN(n17951) );
  OAI221_X1 U21170 ( .B1(n17953), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n17952), 
        .C2(n18061), .A(n17951), .ZN(P3_U2704) );
  NAND2_X1 U21171 ( .A1(n18942), .A2(n18061), .ZN(n18029) );
  AOI22_X1 U21172 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18025), .ZN(n17956) );
  OAI211_X1 U21173 ( .C1(n17954), .C2(P3_EAX_REG_30__SCAN_IN), .A(n18095), .B(
        n17953), .ZN(n17955) );
  OAI211_X1 U21174 ( .C1(n17957), .C2(n18098), .A(n17956), .B(n17955), .ZN(
        P3_U2705) );
  OAI21_X1 U21175 ( .B1(n17960), .B2(n17959), .A(n17958), .ZN(n17964) );
  AOI22_X1 U21176 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18025), .ZN(n17963) );
  OAI211_X1 U21177 ( .C1(n17967), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18095), .B(
        n17961), .ZN(n17962) );
  OAI211_X1 U21178 ( .C1(n17964), .C2(n18098), .A(n17963), .B(n17962), .ZN(
        P3_U2706) );
  INV_X1 U21179 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18047) );
  INV_X1 U21180 ( .A(n17965), .ZN(n17966) );
  OAI22_X1 U21181 ( .A1(n18047), .A2(n18029), .B1(n18098), .B2(n17966), .ZN(
        n17969) );
  AOI211_X1 U21182 ( .C1(n18167), .C2(n17971), .A(n17967), .B(n18061), .ZN(
        n17968) );
  AOI211_X1 U21183 ( .C1(n18025), .C2(BUF2_REG_28__SCAN_IN), .A(n17969), .B(
        n17968), .ZN(n17970) );
  INV_X1 U21184 ( .A(n17970), .ZN(P3_U2707) );
  AOI22_X1 U21185 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18025), .ZN(n17973) );
  OAI211_X1 U21186 ( .C1(n17975), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18095), .B(
        n17971), .ZN(n17972) );
  OAI211_X1 U21187 ( .C1(n17974), .C2(n18098), .A(n17973), .B(n17972), .ZN(
        P3_U2708) );
  AOI22_X1 U21188 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18025), .ZN(n17978) );
  AOI211_X1 U21189 ( .C1(n18163), .C2(n17980), .A(n17975), .B(n18061), .ZN(
        n17976) );
  INV_X1 U21190 ( .A(n17976), .ZN(n17977) );
  OAI211_X1 U21191 ( .C1(n17979), .C2(n18098), .A(n17978), .B(n17977), .ZN(
        P3_U2709) );
  AOI22_X1 U21192 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18025), .ZN(n17983) );
  OAI211_X1 U21193 ( .C1(n17981), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18095), .B(
        n17980), .ZN(n17982) );
  OAI211_X1 U21194 ( .C1(n17984), .C2(n18098), .A(n17983), .B(n17982), .ZN(
        P3_U2710) );
  AOI22_X1 U21195 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18025), .ZN(n17988) );
  OAI211_X1 U21196 ( .C1(n17986), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18095), .B(
        n17985), .ZN(n17987) );
  OAI211_X1 U21197 ( .C1(n17989), .C2(n18098), .A(n17988), .B(n17987), .ZN(
        P3_U2711) );
  AOI22_X1 U21198 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18025), .ZN(n17993) );
  OAI211_X1 U21199 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17991), .A(n18095), .B(
        n17990), .ZN(n17992) );
  OAI211_X1 U21200 ( .C1(n17994), .C2(n18098), .A(n17993), .B(n17992), .ZN(
        P3_U2712) );
  AOI22_X1 U21201 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18025), .B1(n18049), .B2(
        n17995), .ZN(n17998) );
  INV_X1 U21202 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18149) );
  NOR2_X1 U21203 ( .A1(n18087), .A2(n18026), .ZN(n18020) );
  NAND2_X1 U21204 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n18020), .ZN(n18019) );
  NAND2_X1 U21205 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18008), .ZN(n18004) );
  NAND2_X1 U21206 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18000), .ZN(n17999) );
  OAI21_X1 U21207 ( .B1(n18155), .B2(n18061), .A(n17999), .ZN(n17996) );
  OAI21_X1 U21208 ( .B1(n18155), .B2(n17999), .A(n17996), .ZN(n17997) );
  OAI211_X1 U21209 ( .C1(n21197), .C2(n18029), .A(n17998), .B(n17997), .ZN(
        P3_U2713) );
  AOI22_X1 U21210 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18025), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n18018), .ZN(n18002) );
  OAI211_X1 U21211 ( .C1(n18000), .C2(P3_EAX_REG_21__SCAN_IN), .A(n18095), .B(
        n17999), .ZN(n18001) );
  OAI211_X1 U21212 ( .C1(n18003), .C2(n18098), .A(n18002), .B(n18001), .ZN(
        P3_U2714) );
  AOI22_X1 U21213 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18025), .ZN(n18006) );
  OAI211_X1 U21214 ( .C1(n18008), .C2(P3_EAX_REG_20__SCAN_IN), .A(n18095), .B(
        n18004), .ZN(n18005) );
  OAI211_X1 U21215 ( .C1(n18007), .C2(n18098), .A(n18006), .B(n18005), .ZN(
        P3_U2715) );
  AOI22_X1 U21216 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18025), .ZN(n18011) );
  AOI211_X1 U21217 ( .C1(n18149), .C2(n18013), .A(n18008), .B(n18061), .ZN(
        n18009) );
  INV_X1 U21218 ( .A(n18009), .ZN(n18010) );
  OAI211_X1 U21219 ( .C1(n18012), .C2(n18098), .A(n18011), .B(n18010), .ZN(
        P3_U2716) );
  AOI22_X1 U21220 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18025), .ZN(n18016) );
  OAI211_X1 U21221 ( .C1(n18014), .C2(P3_EAX_REG_18__SCAN_IN), .A(n18095), .B(
        n18013), .ZN(n18015) );
  OAI211_X1 U21222 ( .C1(n18017), .C2(n18098), .A(n18016), .B(n18015), .ZN(
        P3_U2717) );
  AOI22_X1 U21223 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18018), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18025), .ZN(n18022) );
  OAI211_X1 U21224 ( .C1(n18020), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18095), .B(
        n18019), .ZN(n18021) );
  OAI211_X1 U21225 ( .C1(n18023), .C2(n18098), .A(n18022), .B(n18021), .ZN(
        P3_U2718) );
  AOI22_X1 U21226 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n18025), .B1(n18049), .B2(
        n18024), .ZN(n18028) );
  OAI211_X1 U21227 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18030), .A(n18095), .B(
        n18026), .ZN(n18027) );
  OAI211_X1 U21228 ( .C1(n18029), .C2(n18917), .A(n18028), .B(n18027), .ZN(
        P3_U2719) );
  INV_X1 U21229 ( .A(n18091), .ZN(n18093) );
  AOI211_X1 U21230 ( .C1(n18208), .C2(n18035), .A(n18061), .B(n18030), .ZN(
        n18031) );
  AOI21_X1 U21231 ( .B1(n18093), .B2(BUF2_REG_15__SCAN_IN), .A(n18031), .ZN(
        n18032) );
  OAI21_X1 U21232 ( .B1(n18033), .B2(n18098), .A(n18032), .ZN(P3_U2720) );
  INV_X1 U21233 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18195) );
  INV_X1 U21234 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18191) );
  NOR2_X1 U21235 ( .A1(n18087), .A2(n18062), .ZN(n18070) );
  NAND2_X1 U21236 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18070), .ZN(n18056) );
  NAND2_X1 U21237 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18059), .ZN(n18051) );
  NOR2_X1 U21238 ( .A1(n18195), .A2(n18051), .ZN(n18043) );
  NAND2_X1 U21239 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18043), .ZN(n18042) );
  NOR2_X1 U21240 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18042), .ZN(n18034) );
  AOI22_X1 U21241 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18093), .B1(
        P3_EAX_REG_13__SCAN_IN), .B2(n18034), .ZN(n18037) );
  NAND3_X1 U21242 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18095), .A3(n18035), 
        .ZN(n18036) );
  OAI211_X1 U21243 ( .C1(n18038), .C2(n18098), .A(n18037), .B(n18036), .ZN(
        P3_U2721) );
  NAND2_X1 U21244 ( .A1(n18042), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n18041) );
  AOI22_X1 U21245 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18093), .B1(n18049), .B2(
        n18039), .ZN(n18040) );
  OAI221_X1 U21246 ( .B1(n18042), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n18041), 
        .C2(n18061), .A(n18040), .ZN(P3_U2722) );
  INV_X1 U21247 ( .A(n18042), .ZN(n18046) );
  AOI21_X1 U21248 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18095), .A(n18043), .ZN(
        n18045) );
  OAI222_X1 U21249 ( .A1(n18091), .A2(n18047), .B1(n18046), .B2(n18045), .C1(
        n18098), .C2(n18044), .ZN(P3_U2723) );
  NAND2_X1 U21250 ( .A1(n18095), .A2(n18051), .ZN(n18054) );
  AOI22_X1 U21251 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18093), .B1(n18049), .B2(
        n18048), .ZN(n18050) );
  OAI221_X1 U21252 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18051), .C1(n18195), 
        .C2(n18054), .A(n18050), .ZN(P3_U2724) );
  INV_X1 U21253 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18055) );
  NOR2_X1 U21254 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18059), .ZN(n18053) );
  OAI222_X1 U21255 ( .A1(n18091), .A2(n18055), .B1(n18054), .B2(n18053), .C1(
        n18098), .C2(n18052), .ZN(P3_U2725) );
  INV_X1 U21256 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21071) );
  INV_X1 U21257 ( .A(n18056), .ZN(n18060) );
  AOI21_X1 U21258 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18095), .A(n18060), .ZN(
        n18058) );
  OAI222_X1 U21259 ( .A1(n18091), .A2(n21071), .B1(n18059), .B2(n18058), .C1(
        n18098), .C2(n18057), .ZN(P3_U2726) );
  INV_X1 U21260 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18189) );
  AOI211_X1 U21261 ( .C1(n18062), .C2(n18189), .A(n18061), .B(n18060), .ZN(
        n18063) );
  AOI21_X1 U21262 ( .B1(n18093), .B2(BUF2_REG_8__SCAN_IN), .A(n18063), .ZN(
        n18064) );
  OAI21_X1 U21263 ( .B1(n18065), .B2(n18098), .A(n18064), .ZN(P3_U2727) );
  INV_X1 U21264 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18951) );
  NOR3_X1 U21265 ( .A1(n18087), .A2(n18094), .A3(n18066), .ZN(n18090) );
  NAND2_X1 U21266 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18090), .ZN(n18079) );
  NOR2_X1 U21267 ( .A1(n18067), .A2(n18079), .ZN(n18074) );
  AOI21_X1 U21268 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18095), .A(n18074), .ZN(
        n18069) );
  OAI222_X1 U21269 ( .A1(n18091), .A2(n18951), .B1(n18070), .B2(n18069), .C1(
        n18098), .C2(n18068), .ZN(P3_U2728) );
  NAND2_X1 U21270 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n18071) );
  NOR2_X1 U21271 ( .A1(n18071), .A2(n18079), .ZN(n18077) );
  AOI21_X1 U21272 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18095), .A(n18077), .ZN(
        n18075) );
  INV_X1 U21273 ( .A(n18072), .ZN(n18073) );
  OAI222_X1 U21274 ( .A1(n18091), .A2(n21197), .B1(n18075), .B2(n18074), .C1(
        n18098), .C2(n18073), .ZN(P3_U2729) );
  INV_X1 U21275 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18941) );
  INV_X1 U21276 ( .A(n18079), .ZN(n18086) );
  AOI22_X1 U21277 ( .A1(n18086), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n18095), .ZN(n18078) );
  OAI222_X1 U21278 ( .A1(n18091), .A2(n18941), .B1(n18078), .B2(n18077), .C1(
        n18098), .C2(n18076), .ZN(P3_U2730) );
  INV_X1 U21279 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18181) );
  NOR2_X1 U21280 ( .A1(n18181), .A2(n18079), .ZN(n18083) );
  AOI21_X1 U21281 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18095), .A(n18086), .ZN(
        n18082) );
  INV_X1 U21282 ( .A(n18080), .ZN(n18081) );
  OAI222_X1 U21283 ( .A1(n18937), .A2(n18091), .B1(n18083), .B2(n18082), .C1(
        n18098), .C2(n18081), .ZN(P3_U2731) );
  INV_X1 U21284 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18933) );
  AOI21_X1 U21285 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18095), .A(n18090), .ZN(
        n18085) );
  OAI222_X1 U21286 ( .A1(n18933), .A2(n18091), .B1(n18086), .B2(n18085), .C1(
        n18098), .C2(n18084), .ZN(P3_U2732) );
  INV_X1 U21287 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18929) );
  NOR2_X1 U21288 ( .A1(n18087), .A2(n18094), .ZN(n18092) );
  AOI22_X1 U21289 ( .A1(n18092), .A2(P3_EAX_REG_1__SCAN_IN), .B1(
        P3_EAX_REG_2__SCAN_IN), .B2(n18095), .ZN(n18089) );
  OAI222_X1 U21290 ( .A1(n18929), .A2(n18091), .B1(n18090), .B2(n18089), .C1(
        n18098), .C2(n18088), .ZN(P3_U2733) );
  INV_X1 U21291 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18175) );
  AOI22_X1 U21292 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18093), .B1(n18092), .B2(
        n18175), .ZN(n18097) );
  NAND3_X1 U21293 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n18095), .A3(n18094), .ZN(
        n18096) );
  OAI211_X1 U21294 ( .C1(n18099), .C2(n18098), .A(n18097), .B(n18096), .ZN(
        P3_U2734) );
  AND2_X1 U21295 ( .A1(n18131), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U21296 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18171) );
  NAND2_X1 U21297 ( .A1(n18119), .A2(n18102), .ZN(n18118) );
  AOI22_X1 U21298 ( .A1(n19569), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18103) );
  OAI21_X1 U21299 ( .B1(n18171), .B2(n18118), .A(n18103), .ZN(P3_U2737) );
  INV_X1 U21300 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18169) );
  AOI22_X1 U21301 ( .A1(n19569), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18104) );
  OAI21_X1 U21302 ( .B1(n18169), .B2(n18118), .A(n18104), .ZN(P3_U2738) );
  AOI22_X1 U21303 ( .A1(n19569), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18131), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18105) );
  OAI21_X1 U21304 ( .B1(n18167), .B2(n18118), .A(n18105), .ZN(P3_U2739) );
  INV_X1 U21305 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18165) );
  AOI22_X1 U21306 ( .A1(n19569), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18131), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18106) );
  OAI21_X1 U21307 ( .B1(n18165), .B2(n18118), .A(n18106), .ZN(P3_U2740) );
  AOI22_X1 U21308 ( .A1(P3_UWORD_REG_10__SCAN_IN), .A2(n19569), .B1(n18137), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18107) );
  OAI21_X1 U21309 ( .B1(n18163), .B2(n18118), .A(n18107), .ZN(P3_U2741) );
  INV_X1 U21310 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18161) );
  AOI22_X1 U21311 ( .A1(n19569), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18131), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18108) );
  OAI21_X1 U21312 ( .B1(n18161), .B2(n18118), .A(n18108), .ZN(P3_U2742) );
  INV_X1 U21313 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18159) );
  AOI22_X1 U21314 ( .A1(n19569), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18131), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18109) );
  OAI21_X1 U21315 ( .B1(n18159), .B2(n18118), .A(n18109), .ZN(P3_U2743) );
  INV_X1 U21316 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18157) );
  AOI22_X1 U21317 ( .A1(n19569), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18110) );
  OAI21_X1 U21318 ( .B1(n18157), .B2(n18118), .A(n18110), .ZN(P3_U2744) );
  AOI22_X1 U21319 ( .A1(n19569), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18111) );
  OAI21_X1 U21320 ( .B1(n18155), .B2(n18118), .A(n18111), .ZN(P3_U2745) );
  AOI22_X1 U21321 ( .A1(n18129), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18112) );
  OAI21_X1 U21322 ( .B1(n18153), .B2(n18118), .A(n18112), .ZN(P3_U2746) );
  INV_X1 U21323 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18151) );
  AOI22_X1 U21324 ( .A1(n18129), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18113) );
  OAI21_X1 U21325 ( .B1(n18151), .B2(n18118), .A(n18113), .ZN(P3_U2747) );
  AOI22_X1 U21326 ( .A1(n18129), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18114) );
  OAI21_X1 U21327 ( .B1(n18149), .B2(n18118), .A(n18114), .ZN(P3_U2748) );
  INV_X1 U21328 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18147) );
  AOI22_X1 U21329 ( .A1(n18129), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18115) );
  OAI21_X1 U21330 ( .B1(n18147), .B2(n18118), .A(n18115), .ZN(P3_U2749) );
  INV_X1 U21331 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18145) );
  AOI22_X1 U21332 ( .A1(n18129), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18116) );
  OAI21_X1 U21333 ( .B1(n18145), .B2(n18118), .A(n18116), .ZN(P3_U2750) );
  INV_X1 U21334 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18143) );
  AOI22_X1 U21335 ( .A1(n18129), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18117) );
  OAI21_X1 U21336 ( .B1(n18143), .B2(n18118), .A(n18117), .ZN(P3_U2751) );
  AOI22_X1 U21337 ( .A1(n18129), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18120) );
  OAI21_X1 U21338 ( .B1(n18208), .B2(n18139), .A(n18120), .ZN(P3_U2752) );
  INV_X1 U21339 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18203) );
  AOI22_X1 U21340 ( .A1(n18129), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18121) );
  OAI21_X1 U21341 ( .B1(n18203), .B2(n18139), .A(n18121), .ZN(P3_U2753) );
  INV_X1 U21342 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18201) );
  AOI22_X1 U21343 ( .A1(n18129), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18122) );
  OAI21_X1 U21344 ( .B1(n18201), .B2(n18139), .A(n18122), .ZN(P3_U2754) );
  INV_X1 U21345 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18198) );
  AOI22_X1 U21346 ( .A1(n18129), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18123) );
  OAI21_X1 U21347 ( .B1(n18198), .B2(n18139), .A(n18123), .ZN(P3_U2755) );
  AOI22_X1 U21348 ( .A1(n19569), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18131), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18124) );
  OAI21_X1 U21349 ( .B1(n18195), .B2(n18139), .A(n18124), .ZN(P3_U2756) );
  INV_X1 U21350 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18193) );
  AOI22_X1 U21351 ( .A1(n19569), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18131), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18125) );
  OAI21_X1 U21352 ( .B1(n18193), .B2(n18139), .A(n18125), .ZN(P3_U2757) );
  AOI22_X1 U21353 ( .A1(n19569), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18131), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18126) );
  OAI21_X1 U21354 ( .B1(n18191), .B2(n18139), .A(n18126), .ZN(P3_U2758) );
  AOI22_X1 U21355 ( .A1(n19569), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18131), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18127) );
  OAI21_X1 U21356 ( .B1(n18189), .B2(n18139), .A(n18127), .ZN(P3_U2759) );
  INV_X1 U21357 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18187) );
  AOI22_X1 U21358 ( .A1(n19569), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18131), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18128) );
  OAI21_X1 U21359 ( .B1(n18187), .B2(n18139), .A(n18128), .ZN(P3_U2760) );
  INV_X1 U21360 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18185) );
  AOI22_X1 U21361 ( .A1(n18129), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18130) );
  OAI21_X1 U21362 ( .B1(n18185), .B2(n18139), .A(n18130), .ZN(P3_U2761) );
  INV_X1 U21363 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18183) );
  AOI22_X1 U21364 ( .A1(n19569), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18131), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18132) );
  OAI21_X1 U21365 ( .B1(n18183), .B2(n18139), .A(n18132), .ZN(P3_U2762) );
  AOI22_X1 U21366 ( .A1(n19569), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18133) );
  OAI21_X1 U21367 ( .B1(n18181), .B2(n18139), .A(n18133), .ZN(P3_U2763) );
  INV_X1 U21368 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18179) );
  AOI22_X1 U21369 ( .A1(n19569), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18134) );
  OAI21_X1 U21370 ( .B1(n18179), .B2(n18139), .A(n18134), .ZN(P3_U2764) );
  INV_X1 U21371 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18177) );
  AOI22_X1 U21372 ( .A1(n19569), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18135) );
  OAI21_X1 U21373 ( .B1(n18177), .B2(n18139), .A(n18135), .ZN(P3_U2765) );
  AOI22_X1 U21374 ( .A1(n19569), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18136) );
  OAI21_X1 U21375 ( .B1(n18175), .B2(n18139), .A(n18136), .ZN(P3_U2766) );
  AOI22_X1 U21376 ( .A1(n19569), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18137), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18138) );
  OAI21_X1 U21377 ( .B1(n18173), .B2(n18139), .A(n18138), .ZN(P3_U2767) );
  NAND2_X2 U21378 ( .A1(n18140), .A2(n19415), .ZN(n18207) );
  AOI22_X1 U21379 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18205), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18204), .ZN(n18142) );
  OAI21_X1 U21380 ( .B1(n18143), .B2(n18207), .A(n18142), .ZN(P3_U2768) );
  AOI22_X1 U21381 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18205), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18204), .ZN(n18144) );
  OAI21_X1 U21382 ( .B1(n18145), .B2(n18207), .A(n18144), .ZN(P3_U2769) );
  AOI22_X1 U21383 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18205), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18204), .ZN(n18146) );
  OAI21_X1 U21384 ( .B1(n18147), .B2(n18207), .A(n18146), .ZN(P3_U2770) );
  AOI22_X1 U21385 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18196), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18204), .ZN(n18148) );
  OAI21_X1 U21386 ( .B1(n18149), .B2(n18207), .A(n18148), .ZN(P3_U2771) );
  AOI22_X1 U21387 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18196), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18204), .ZN(n18150) );
  OAI21_X1 U21388 ( .B1(n18151), .B2(n18207), .A(n18150), .ZN(P3_U2772) );
  AOI22_X1 U21389 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18196), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18204), .ZN(n18152) );
  OAI21_X1 U21390 ( .B1(n18153), .B2(n18207), .A(n18152), .ZN(P3_U2773) );
  AOI22_X1 U21391 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18196), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18204), .ZN(n18154) );
  OAI21_X1 U21392 ( .B1(n18155), .B2(n18207), .A(n18154), .ZN(P3_U2774) );
  AOI22_X1 U21393 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18196), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18204), .ZN(n18156) );
  OAI21_X1 U21394 ( .B1(n18157), .B2(n18207), .A(n18156), .ZN(P3_U2775) );
  AOI22_X1 U21395 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18196), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18204), .ZN(n18158) );
  OAI21_X1 U21396 ( .B1(n18159), .B2(n18207), .A(n18158), .ZN(P3_U2776) );
  AOI22_X1 U21397 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18196), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18204), .ZN(n18160) );
  OAI21_X1 U21398 ( .B1(n18161), .B2(n18207), .A(n18160), .ZN(P3_U2777) );
  AOI22_X1 U21399 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18196), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18204), .ZN(n18162) );
  OAI21_X1 U21400 ( .B1(n18163), .B2(n18207), .A(n18162), .ZN(P3_U2778) );
  AOI22_X1 U21401 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18196), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18204), .ZN(n18164) );
  OAI21_X1 U21402 ( .B1(n18165), .B2(n18207), .A(n18164), .ZN(P3_U2779) );
  AOI22_X1 U21403 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18205), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18204), .ZN(n18166) );
  OAI21_X1 U21404 ( .B1(n18167), .B2(n18207), .A(n18166), .ZN(P3_U2780) );
  AOI22_X1 U21405 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18205), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18204), .ZN(n18168) );
  OAI21_X1 U21406 ( .B1(n18169), .B2(n18207), .A(n18168), .ZN(P3_U2781) );
  AOI22_X1 U21407 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18205), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18204), .ZN(n18170) );
  OAI21_X1 U21408 ( .B1(n18171), .B2(n18207), .A(n18170), .ZN(P3_U2782) );
  AOI22_X1 U21409 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18204), .ZN(n18172) );
  OAI21_X1 U21410 ( .B1(n18173), .B2(n18207), .A(n18172), .ZN(P3_U2783) );
  AOI22_X1 U21411 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18204), .ZN(n18174) );
  OAI21_X1 U21412 ( .B1(n18175), .B2(n18207), .A(n18174), .ZN(P3_U2784) );
  AOI22_X1 U21413 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18199), .ZN(n18176) );
  OAI21_X1 U21414 ( .B1(n18177), .B2(n18207), .A(n18176), .ZN(P3_U2785) );
  AOI22_X1 U21415 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18199), .ZN(n18178) );
  OAI21_X1 U21416 ( .B1(n18179), .B2(n18207), .A(n18178), .ZN(P3_U2786) );
  AOI22_X1 U21417 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18199), .ZN(n18180) );
  OAI21_X1 U21418 ( .B1(n18181), .B2(n18207), .A(n18180), .ZN(P3_U2787) );
  AOI22_X1 U21419 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18199), .ZN(n18182) );
  OAI21_X1 U21420 ( .B1(n18183), .B2(n18207), .A(n18182), .ZN(P3_U2788) );
  AOI22_X1 U21421 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18199), .ZN(n18184) );
  OAI21_X1 U21422 ( .B1(n18185), .B2(n18207), .A(n18184), .ZN(P3_U2789) );
  AOI22_X1 U21423 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18199), .ZN(n18186) );
  OAI21_X1 U21424 ( .B1(n18187), .B2(n18207), .A(n18186), .ZN(P3_U2790) );
  AOI22_X1 U21425 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18199), .ZN(n18188) );
  OAI21_X1 U21426 ( .B1(n18189), .B2(n18207), .A(n18188), .ZN(P3_U2791) );
  AOI22_X1 U21427 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18199), .ZN(n18190) );
  OAI21_X1 U21428 ( .B1(n18191), .B2(n18207), .A(n18190), .ZN(P3_U2792) );
  AOI22_X1 U21429 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18196), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18204), .ZN(n18192) );
  OAI21_X1 U21430 ( .B1(n18193), .B2(n18207), .A(n18192), .ZN(P3_U2793) );
  AOI22_X1 U21431 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18199), .ZN(n18194) );
  OAI21_X1 U21432 ( .B1(n18195), .B2(n18207), .A(n18194), .ZN(P3_U2794) );
  AOI22_X1 U21433 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18196), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18204), .ZN(n18197) );
  OAI21_X1 U21434 ( .B1(n18198), .B2(n18207), .A(n18197), .ZN(P3_U2795) );
  AOI22_X1 U21435 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18199), .ZN(n18200) );
  OAI21_X1 U21436 ( .B1(n18201), .B2(n18207), .A(n18200), .ZN(P3_U2796) );
  AOI22_X1 U21437 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18204), .ZN(n18202) );
  OAI21_X1 U21438 ( .B1(n18203), .B2(n18207), .A(n18202), .ZN(P3_U2797) );
  AOI22_X1 U21439 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18205), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18204), .ZN(n18206) );
  OAI21_X1 U21440 ( .B1(n18208), .B2(n18207), .A(n18206), .ZN(P3_U2798) );
  NOR2_X1 U21441 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18209), .ZN(
        n18216) );
  INV_X1 U21442 ( .A(n18420), .ZN(n18379) );
  OR2_X1 U21443 ( .A1(n19432), .A2(n18210), .ZN(n18211) );
  OAI211_X1 U21444 ( .C1(n18212), .C2(n18489), .A(n18587), .B(n18211), .ZN(
        n18247) );
  AOI21_X1 U21445 ( .B1(n18299), .B2(n18242), .A(n18247), .ZN(n18239) );
  NAND3_X1 U21446 ( .A1(n18212), .A2(n18379), .A3(n18238), .ZN(n18236) );
  AOI21_X1 U21447 ( .B1(n18239), .B2(n18236), .A(n18213), .ZN(n18215) );
  AOI211_X1 U21448 ( .C1(n18216), .C2(n18379), .A(n18215), .B(n18214), .ZN(
        n18225) );
  NOR2_X1 U21449 ( .A1(n18498), .A2(n18550), .ZN(n18323) );
  OAI22_X1 U21450 ( .A1(n18595), .A2(n18429), .B1(n18594), .B2(n18591), .ZN(
        n18248) );
  NOR2_X1 U21451 ( .A1(n9988), .A2(n18248), .ZN(n18230) );
  NOR3_X1 U21452 ( .A1(n18323), .A2(n18230), .A3(n18217), .ZN(n18222) );
  AOI211_X1 U21453 ( .C1(n18220), .C2(n18219), .A(n18218), .B(n18471), .ZN(
        n18221) );
  AOI211_X1 U21454 ( .C1(n18223), .C2(n18388), .A(n18222), .B(n18221), .ZN(
        n18224) );
  OAI211_X1 U21455 ( .C1(n18436), .C2(n18226), .A(n18225), .B(n18224), .ZN(
        P3_U2802) );
  NAND2_X1 U21456 ( .A1(n9986), .A2(n18228), .ZN(n18229) );
  XOR2_X1 U21457 ( .A(n18496), .B(n18229), .Z(n18593) );
  AOI21_X1 U21458 ( .B1(n9988), .B2(n18231), .A(n18230), .ZN(n18235) );
  AOI22_X1 U21459 ( .A1(n18902), .A2(P3_REIP_REG_27__SCAN_IN), .B1(n18427), 
        .B2(n18232), .ZN(n18233) );
  INV_X1 U21460 ( .A(n18233), .ZN(n18234) );
  AOI211_X1 U21461 ( .C1(n18497), .C2(n18593), .A(n18235), .B(n18234), .ZN(
        n18237) );
  OAI211_X1 U21462 ( .C1(n18239), .C2(n18238), .A(n18237), .B(n18236), .ZN(
        P3_U2803) );
  AOI21_X1 U21463 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18241), .A(
        n18240), .ZN(n18610) );
  OAI21_X1 U21464 ( .B1(n18243), .B2(n18949), .A(n18242), .ZN(n18246) );
  AOI21_X1 U21465 ( .B1(n18436), .B2(n18364), .A(n18244), .ZN(n18245) );
  NOR2_X1 U21466 ( .A1(n18890), .A2(n19501), .ZN(n18605) );
  AOI211_X1 U21467 ( .C1(n18247), .C2(n18246), .A(n18245), .B(n18605), .ZN(
        n18250) );
  NOR3_X1 U21468 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18612), .A3(
        n18614), .ZN(n18606) );
  AOI22_X1 U21469 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18248), .B1(
        n18388), .B2(n18606), .ZN(n18249) );
  OAI211_X1 U21470 ( .C1(n18610), .C2(n18471), .A(n18250), .B(n18249), .ZN(
        P3_U2804) );
  NAND2_X1 U21471 ( .A1(n18272), .A2(n18251), .ZN(n18628) );
  INV_X1 U21472 ( .A(n18628), .ZN(n18252) );
  NAND2_X1 U21473 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18252), .ZN(
        n18253) );
  XOR2_X1 U21474 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18253), .Z(
        n18625) );
  NAND2_X1 U21475 ( .A1(n9713), .A2(n18379), .ZN(n18268) );
  AOI221_X1 U21476 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C1(n9951), .C2(n9952), .A(n18268), 
        .ZN(n18256) );
  OR2_X1 U21477 ( .A1(n18949), .A2(n9713), .ZN(n18284) );
  OAI211_X1 U21478 ( .C1(n18280), .C2(n19432), .A(n18587), .B(n18284), .ZN(
        n18290) );
  AOI21_X1 U21479 ( .B1(n18299), .B2(n18254), .A(n18290), .ZN(n18267) );
  OAI22_X1 U21480 ( .A1(n18267), .A2(n9952), .B1(n18890), .B2(n19499), .ZN(
        n18255) );
  AOI211_X1 U21481 ( .C1(n18257), .C2(n18427), .A(n18256), .B(n18255), .ZN(
        n18263) );
  INV_X1 U21482 ( .A(n18718), .ZN(n18305) );
  NAND3_X1 U21483 ( .A1(n18305), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n18272), .ZN(n18258) );
  XOR2_X1 U21484 ( .A(n18258), .B(n18612), .Z(n18622) );
  AOI21_X1 U21485 ( .B1(n18260), .B2(n18404), .A(n18259), .ZN(n18261) );
  XOR2_X1 U21486 ( .A(n18261), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18621) );
  AOI22_X1 U21487 ( .A1(n18498), .A2(n18622), .B1(n18497), .B2(n18621), .ZN(
        n18262) );
  OAI211_X1 U21488 ( .C1(n18591), .C2(n18625), .A(n18263), .B(n18262), .ZN(
        P3_U2805) );
  AOI21_X1 U21489 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18265), .A(
        n18264), .ZN(n18637) );
  NAND2_X1 U21490 ( .A1(n18902), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18266) );
  OAI221_X1 U21491 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18268), .C1(
        n9951), .C2(n18267), .A(n18266), .ZN(n18269) );
  AOI21_X1 U21492 ( .B1(n18427), .B2(n18270), .A(n18269), .ZN(n18275) );
  NAND2_X1 U21493 ( .A1(n18305), .A2(n18272), .ZN(n18627) );
  AOI22_X1 U21494 ( .A1(n18498), .A2(n18627), .B1(n18550), .B2(n18628), .ZN(
        n18271) );
  INV_X1 U21495 ( .A(n18271), .ZN(n18286) );
  INV_X1 U21496 ( .A(n18272), .ZN(n18273) );
  NOR2_X1 U21497 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18273), .ZN(
        n18626) );
  AOI22_X1 U21498 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18286), .B1(
        n18388), .B2(n18626), .ZN(n18274) );
  OAI211_X1 U21499 ( .C1(n18637), .C2(n18471), .A(n18275), .B(n18274), .ZN(
        P3_U2806) );
  AOI22_X1 U21500 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18404), .B1(
        n18276), .B2(n18292), .ZN(n18277) );
  NAND2_X1 U21501 ( .A1(n18324), .A2(n18277), .ZN(n18278) );
  XOR2_X1 U21502 ( .A(n18278), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n18644) );
  NOR2_X1 U21503 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18364), .ZN(
        n18279) );
  AOI22_X1 U21504 ( .A1(n18427), .A2(n18281), .B1(n18280), .B2(n18279), .ZN(
        n18282) );
  NAND2_X1 U21505 ( .A1(n18902), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18643) );
  OAI211_X1 U21506 ( .C1(n18284), .C2(n18283), .A(n18282), .B(n18643), .ZN(
        n18289) );
  INV_X1 U21507 ( .A(n18388), .ZN(n18285) );
  NOR2_X1 U21508 ( .A1(n18638), .A2(n18285), .ZN(n18287) );
  MUX2_X1 U21509 ( .A(n18287), .B(n18286), .S(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n18288) );
  AOI211_X1 U21510 ( .C1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n18290), .A(
        n18289), .B(n18288), .ZN(n18291) );
  OAI21_X1 U21511 ( .B1(n18471), .B2(n18644), .A(n18291), .ZN(P3_U2807) );
  INV_X1 U21512 ( .A(n18292), .ZN(n18294) );
  NOR2_X1 U21513 ( .A1(n18322), .A2(n18652), .ZN(n18653) );
  OAI221_X1 U21514 ( .B1(n18294), .B2(n18293), .C1(n18294), .C2(n18653), .A(
        n18324), .ZN(n18295) );
  XOR2_X1 U21515 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18295), .Z(
        n18659) );
  NOR2_X1 U21516 ( .A1(n18890), .A2(n19493), .ZN(n18657) );
  NAND2_X1 U21517 ( .A1(n18378), .A2(n18296), .ZN(n18297) );
  OAI211_X1 U21518 ( .C1(n18300), .C2(n18489), .A(n18587), .B(n18297), .ZN(
        n18328) );
  AOI21_X1 U21519 ( .B1(n18299), .B2(n18298), .A(n18328), .ZN(n18309) );
  NAND2_X1 U21520 ( .A1(n18300), .A2(n18379), .ZN(n18311) );
  AOI22_X1 U21521 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18302), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18310), .ZN(n18301) );
  OAI22_X1 U21522 ( .A1(n18309), .A2(n18302), .B1(n18311), .B2(n18301), .ZN(
        n18303) );
  AOI211_X1 U21523 ( .C1(n18304), .C2(n18427), .A(n18657), .B(n18303), .ZN(
        n18307) );
  NOR2_X1 U21524 ( .A1(n18305), .A2(n18429), .ZN(n18399) );
  AOI21_X1 U21525 ( .B1(n18550), .B2(n18717), .A(n18399), .ZN(n18349) );
  OAI21_X1 U21526 ( .B1(n18323), .B2(n18653), .A(n18349), .ZN(n18319) );
  OAI222_X1 U21527 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18388), 
        .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18653), .C1(n18650), 
        .C2(n18319), .ZN(n18306) );
  OAI211_X1 U21528 ( .C1(n18471), .C2(n18659), .A(n18307), .B(n18306), .ZN(
        P3_U2808) );
  NAND2_X1 U21529 ( .A1(n18664), .A2(n18318), .ZN(n18668) );
  NAND2_X1 U21530 ( .A1(n18661), .A2(n18388), .ZN(n18347) );
  NAND2_X1 U21531 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n18902), .ZN(n18308) );
  OAI221_X1 U21532 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18311), .C1(
        n18310), .C2(n18309), .A(n18308), .ZN(n18312) );
  AOI21_X1 U21533 ( .B1(n18427), .B2(n18313), .A(n18312), .ZN(n18321) );
  INV_X1 U21534 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18360) );
  NOR3_X1 U21535 ( .A1(n18404), .A2(n18360), .A3(n18314), .ZN(n18342) );
  INV_X1 U21536 ( .A(n18315), .ZN(n18356) );
  AOI22_X1 U21537 ( .A1(n18664), .A2(n18342), .B1(n18356), .B2(n18316), .ZN(
        n18317) );
  XOR2_X1 U21538 ( .A(n18318), .B(n18317), .Z(n18662) );
  AOI22_X1 U21539 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18319), .B1(
        n18497), .B2(n18662), .ZN(n18320) );
  OAI211_X1 U21540 ( .C1(n18668), .C2(n18347), .A(n18321), .B(n18320), .ZN(
        P3_U2809) );
  NAND2_X1 U21541 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18326), .ZN(
        n18679) );
  NOR2_X1 U21542 ( .A1(n18322), .A2(n18683), .ZN(n18670) );
  OAI21_X1 U21543 ( .B1(n18323), .B2(n18670), .A(n18349), .ZN(n18344) );
  OAI221_X1 U21544 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18355), 
        .C1(n18683), .C2(n18342), .A(n18324), .ZN(n18325) );
  XOR2_X1 U21545 ( .A(n18326), .B(n18325), .Z(n18675) );
  AOI22_X1 U21546 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18344), .B1(
        n18497), .B2(n18675), .ZN(n18333) );
  NAND2_X1 U21547 ( .A1(n18902), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18677) );
  AND2_X1 U21548 ( .A1(n18950), .A2(n18327), .ZN(n18361) );
  OAI221_X1 U21549 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18329), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18361), .A(n18328), .ZN(
        n18332) );
  OAI21_X1 U21550 ( .B1(n18427), .B2(n18299), .A(n18330), .ZN(n18331) );
  AND4_X1 U21551 ( .A1(n18333), .A2(n18677), .A3(n18332), .A4(n18331), .ZN(
        n18334) );
  OAI21_X1 U21552 ( .B1(n18679), .B2(n18347), .A(n18334), .ZN(P3_U2810) );
  OAI21_X1 U21553 ( .B1(n18573), .B2(n18336), .A(n18582), .ZN(n18371) );
  OAI21_X1 U21554 ( .B1(n18335), .B2(n19432), .A(n18371), .ZN(n18352) );
  NOR2_X1 U21555 ( .A1(n18420), .A2(n18336), .ZN(n18354) );
  OAI211_X1 U21556 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18354), .B(n18337), .ZN(n18339) );
  NAND2_X1 U21557 ( .A1(n18902), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18338) );
  OAI211_X1 U21558 ( .C1(n18436), .C2(n18340), .A(n18339), .B(n18338), .ZN(
        n18341) );
  AOI21_X1 U21559 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18352), .A(
        n18341), .ZN(n18346) );
  AOI21_X1 U21560 ( .B1(n18355), .B2(n18356), .A(n18342), .ZN(n18343) );
  XOR2_X1 U21561 ( .A(n18683), .B(n18343), .Z(n18680) );
  AOI22_X1 U21562 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18344), .B1(
        n18497), .B2(n18680), .ZN(n18345) );
  OAI211_X1 U21563 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18347), .A(
        n18346), .B(n18345), .ZN(P3_U2811) );
  INV_X1 U21564 ( .A(n18348), .ZN(n18686) );
  INV_X1 U21565 ( .A(n18349), .ZN(n18387) );
  AOI21_X1 U21566 ( .B1(n18388), .B2(n18686), .A(n18387), .ZN(n18366) );
  INV_X1 U21567 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18353) );
  OAI22_X1 U21568 ( .A1(n18890), .A2(n19485), .B1(n18436), .B2(n18350), .ZN(
        n18351) );
  AOI221_X1 U21569 ( .B1(n18354), .B2(n18353), .C1(n18352), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18351), .ZN(n18359) );
  AOI21_X1 U21570 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18496), .A(
        n18355), .ZN(n18357) );
  XOR2_X1 U21571 ( .A(n18357), .B(n18356), .Z(n18695) );
  NOR2_X1 U21572 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18686), .ZN(
        n18694) );
  AOI22_X1 U21573 ( .A1(n18497), .A2(n18695), .B1(n18388), .B2(n18694), .ZN(
        n18358) );
  OAI211_X1 U21574 ( .C1(n18366), .C2(n18360), .A(n18359), .B(n18358), .ZN(
        P3_U2812) );
  NOR2_X1 U21575 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18361), .ZN(
        n18372) );
  OAI21_X1 U21576 ( .B1(n18363), .B2(n18700), .A(n18362), .ZN(n18698) );
  AOI21_X1 U21577 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18388), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18365) );
  OAI22_X1 U21578 ( .A1(n18571), .A2(n18367), .B1(n18366), .B2(n18365), .ZN(
        n18368) );
  AOI21_X1 U21579 ( .B1(n18497), .B2(n18698), .A(n18368), .ZN(n18370) );
  NAND2_X1 U21580 ( .A1(n18902), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18369) );
  OAI211_X1 U21581 ( .C1(n18372), .C2(n18371), .A(n18370), .B(n18369), .ZN(
        P3_U2813) );
  AOI21_X1 U21582 ( .B1(n18496), .B2(n18374), .A(n18373), .ZN(n18375) );
  XOR2_X1 U21583 ( .A(n18711), .B(n18375), .Z(n18716) );
  INV_X1 U21584 ( .A(n18376), .ZN(n18380) );
  OAI21_X1 U21585 ( .B1(n18380), .B2(n18489), .A(n18587), .ZN(n18407) );
  AOI21_X1 U21586 ( .B1(n18378), .B2(n18377), .A(n18407), .ZN(n18390) );
  NAND2_X1 U21587 ( .A1(n18380), .A2(n18379), .ZN(n18392) );
  AOI21_X1 U21588 ( .B1(n18391), .B2(n18385), .A(n18392), .ZN(n18382) );
  AOI22_X1 U21589 ( .A1(n18383), .A2(n18427), .B1(n18382), .B2(n18381), .ZN(
        n18384) );
  NAND2_X1 U21590 ( .A1(n18902), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18714) );
  OAI211_X1 U21591 ( .C1(n18390), .C2(n18385), .A(n18384), .B(n18714), .ZN(
        n18386) );
  AOI221_X1 U21592 ( .B1(n18388), .B2(n18711), .C1(n18387), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n18386), .ZN(n18389) );
  OAI21_X1 U21593 ( .B1(n18471), .B2(n18716), .A(n18389), .ZN(P3_U2814) );
  INV_X1 U21594 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18416) );
  INV_X1 U21595 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18740) );
  NAND2_X1 U21596 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18751), .ZN(
        n18428) );
  NOR2_X1 U21597 ( .A1(n18428), .A2(n18454), .ZN(n18430) );
  INV_X1 U21598 ( .A(n18430), .ZN(n18752) );
  NOR3_X1 U21599 ( .A1(n18416), .A2(n18740), .A3(n18752), .ZN(n18413) );
  NOR2_X1 U21600 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18413), .ZN(
        n18724) );
  NAND2_X1 U21601 ( .A1(n18550), .A2(n18717), .ZN(n18402) );
  NAND2_X1 U21602 ( .A1(n18902), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18728) );
  OAI221_X1 U21603 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18392), .C1(
        n18391), .C2(n18390), .A(n18728), .ZN(n18393) );
  AOI21_X1 U21604 ( .B1(n18427), .B2(n18394), .A(n18393), .ZN(n18401) );
  NOR4_X1 U21605 ( .A1(n18496), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A4(n18459), .ZN(n18455) );
  INV_X1 U21606 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18757) );
  NAND2_X1 U21607 ( .A1(n18455), .A2(n18757), .ZN(n18442) );
  OAI22_X1 U21608 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18442), .B1(
        n18403), .B2(n18395), .ZN(n18396) );
  OAI221_X1 U21609 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18740), 
        .C1(n18769), .C2(n18496), .A(n18396), .ZN(n18397) );
  XOR2_X1 U21610 ( .A(n18730), .B(n18397), .Z(n18726) );
  NOR2_X1 U21611 ( .A1(n18412), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18722) );
  INV_X1 U21612 ( .A(n18722), .ZN(n18398) );
  AOI22_X1 U21613 ( .A1(n18497), .A2(n18726), .B1(n18399), .B2(n18398), .ZN(
        n18400) );
  OAI211_X1 U21614 ( .C1(n18724), .C2(n18402), .A(n18401), .B(n18400), .ZN(
        P3_U2815) );
  INV_X1 U21615 ( .A(n18428), .ZN(n18733) );
  NOR2_X1 U21616 ( .A1(n18404), .A2(n18403), .ZN(n18473) );
  NAND2_X1 U21617 ( .A1(n18733), .A2(n18473), .ZN(n18431) );
  NAND2_X1 U21618 ( .A1(n18769), .A2(n18416), .ZN(n18405) );
  OAI22_X1 U21619 ( .A1(n18416), .A2(n18431), .B1(n18405), .B2(n18442), .ZN(
        n18406) );
  XOR2_X1 U21620 ( .A(n18740), .B(n18406), .Z(n18746) );
  OAI221_X1 U21621 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19302), .C1(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n18408), .A(n18407), .ZN(
        n18409) );
  OAI21_X1 U21622 ( .B1(n18571), .B2(n18410), .A(n18409), .ZN(n18411) );
  AOI21_X1 U21623 ( .B1(n18902), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18411), 
        .ZN(n18415) );
  NOR2_X1 U21624 ( .A1(n18416), .A2(n18428), .ZN(n18737) );
  INV_X1 U21625 ( .A(n18737), .ZN(n18732) );
  AOI221_X1 U21626 ( .B1(n18779), .B2(n18740), .C1(n18732), .C2(n18740), .A(
        n18412), .ZN(n18743) );
  AOI221_X1 U21627 ( .B1(n18416), .B2(n18740), .C1(n18752), .C2(n18740), .A(
        n18413), .ZN(n18742) );
  AOI22_X1 U21628 ( .A1(n18498), .A2(n18743), .B1(n18550), .B2(n18742), .ZN(
        n18414) );
  OAI211_X1 U21629 ( .C1(n18746), .C2(n18471), .A(n18415), .B(n18414), .ZN(
        P3_U2816) );
  NAND2_X1 U21630 ( .A1(n18733), .A2(n18416), .ZN(n18762) );
  OAI21_X1 U21631 ( .B1(n18417), .B2(n19432), .A(n18587), .ZN(n18418) );
  AOI21_X1 U21632 ( .B1(n18546), .B2(n18419), .A(n18418), .ZN(n18437) );
  NOR2_X1 U21633 ( .A1(n18420), .A2(n18419), .ZN(n18441) );
  OAI211_X1 U21634 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18441), .B(n18421), .ZN(n18423) );
  NAND2_X1 U21635 ( .A1(n18902), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18422) );
  OAI211_X1 U21636 ( .C1(n18437), .C2(n18424), .A(n18423), .B(n18422), .ZN(
        n18425) );
  AOI21_X1 U21637 ( .B1(n18427), .B2(n18426), .A(n18425), .ZN(n18434) );
  NOR2_X1 U21638 ( .A1(n18779), .A2(n18428), .ZN(n18756) );
  OAI22_X1 U21639 ( .A1(n18430), .A2(n18591), .B1(n18756), .B2(n18429), .ZN(
        n18445) );
  OAI21_X1 U21640 ( .B1(n18442), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18431), .ZN(n18432) );
  XOR2_X1 U21641 ( .A(n18432), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18747) );
  AOI22_X1 U21642 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18445), .B1(
        n18497), .B2(n18747), .ZN(n18433) );
  OAI211_X1 U21643 ( .C1(n18482), .C2(n18762), .A(n18434), .B(n18433), .ZN(
        P3_U2817) );
  NAND2_X1 U21644 ( .A1(n18751), .A2(n18769), .ZN(n18448) );
  INV_X1 U21645 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18440) );
  NOR2_X1 U21646 ( .A1(n18890), .A2(n19474), .ZN(n18439) );
  OAI22_X1 U21647 ( .A1(n18437), .A2(n18440), .B1(n18436), .B2(n18435), .ZN(
        n18438) );
  AOI211_X1 U21648 ( .C1(n18441), .C2(n18440), .A(n18439), .B(n18438), .ZN(
        n18447) );
  INV_X1 U21649 ( .A(n18473), .ZN(n18443) );
  OAI21_X1 U21650 ( .B1(n18770), .B2(n18443), .A(n18442), .ZN(n18444) );
  XOR2_X1 U21651 ( .A(n18444), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18763) );
  AOI22_X1 U21652 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18445), .B1(
        n18497), .B2(n18763), .ZN(n18446) );
  OAI211_X1 U21653 ( .C1(n18482), .C2(n18448), .A(n18447), .B(n18446), .ZN(
        P3_U2818) );
  NAND2_X1 U21654 ( .A1(n18748), .A2(n18757), .ZN(n18790) );
  NAND3_X1 U21655 ( .A1(n18950), .A2(n18449), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18464) );
  NAND3_X1 U21656 ( .A1(n18582), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n18464), .ZN(n18451) );
  NAND2_X1 U21657 ( .A1(n18902), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18450) );
  OAI211_X1 U21658 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18464), .A(
        n18451), .B(n18450), .ZN(n18452) );
  AOI21_X1 U21659 ( .B1(n18453), .B2(n18580), .A(n18452), .ZN(n18458) );
  AOI22_X1 U21660 ( .A1(n18498), .A2(n18779), .B1(n18550), .B2(n18454), .ZN(
        n18481) );
  OAI21_X1 U21661 ( .B1(n18748), .B2(n18482), .A(n18481), .ZN(n18467) );
  AOI21_X1 U21662 ( .B1(n18748), .B2(n18473), .A(n18455), .ZN(n18456) );
  XOR2_X1 U21663 ( .A(n18757), .B(n18456), .Z(n18777) );
  AOI22_X1 U21664 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18467), .B1(
        n18497), .B2(n18777), .ZN(n18457) );
  OAI211_X1 U21665 ( .C1(n18482), .C2(n18790), .A(n18458), .B(n18457), .ZN(
        P3_U2819) );
  NOR2_X1 U21666 ( .A1(n18496), .A2(n18459), .ZN(n18472) );
  AOI22_X1 U21667 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18473), .B1(
        n18472), .B2(n18808), .ZN(n18460) );
  XNOR2_X1 U21668 ( .A(n18465), .B(n18460), .ZN(n18800) );
  NOR2_X1 U21669 ( .A1(n18949), .A2(n18461), .ZN(n18477) );
  AOI21_X1 U21670 ( .B1(n18582), .B2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18477), .ZN(n18462) );
  INV_X1 U21671 ( .A(n18462), .ZN(n18463) );
  AOI22_X1 U21672 ( .A1(n18902), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18464), 
        .B2(n18463), .ZN(n18470) );
  OAI21_X1 U21673 ( .B1(n18482), .B2(n18808), .A(n18465), .ZN(n18466) );
  AOI22_X1 U21674 ( .A1(n18468), .A2(n18580), .B1(n18467), .B2(n18466), .ZN(
        n18469) );
  OAI211_X1 U21675 ( .C1(n18800), .C2(n18471), .A(n18470), .B(n18469), .ZN(
        P3_U2820) );
  NOR2_X1 U21676 ( .A1(n18473), .A2(n18472), .ZN(n18474) );
  XOR2_X1 U21677 ( .A(n18474), .B(n18808), .Z(n18805) );
  NOR2_X1 U21678 ( .A1(n18890), .A2(n19467), .ZN(n18479) );
  NOR3_X1 U21679 ( .A1(n18949), .A2(n18517), .A3(n18520), .ZN(n18504) );
  AOI22_X1 U21680 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18582), .B1(
        n18504), .B2(n18485), .ZN(n18476) );
  OAI22_X1 U21681 ( .A1(n18477), .A2(n18476), .B1(n18571), .B2(n18475), .ZN(
        n18478) );
  AOI211_X1 U21682 ( .C1(n18497), .C2(n18805), .A(n18479), .B(n18478), .ZN(
        n18480) );
  OAI221_X1 U21683 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18482), .C1(
        n18808), .C2(n18481), .A(n18480), .ZN(P3_U2821) );
  OAI21_X1 U21684 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18484), .A(
        n18483), .ZN(n18827) );
  AOI211_X1 U21685 ( .C1(n18487), .C2(n18486), .A(n18485), .B(n18949), .ZN(
        n18492) );
  OAI21_X1 U21686 ( .B1(n18489), .B2(n18488), .A(n18587), .ZN(n18503) );
  AOI22_X1 U21687 ( .A1(n18503), .A2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n18902), .B2(P3_REIP_REG_8__SCAN_IN), .ZN(n18490) );
  INV_X1 U21688 ( .A(n18490), .ZN(n18491) );
  AOI211_X1 U21689 ( .C1(n18493), .C2(n18580), .A(n18492), .B(n18491), .ZN(
        n18500) );
  INV_X1 U21690 ( .A(n18495), .ZN(n18824) );
  AOI21_X1 U21691 ( .B1(n18496), .B2(n18495), .A(n18494), .ZN(n18821) );
  AOI22_X1 U21692 ( .A1(n18498), .A2(n18824), .B1(n18497), .B2(n18821), .ZN(
        n18499) );
  OAI211_X1 U21693 ( .C1(n18591), .C2(n18827), .A(n18500), .B(n18499), .ZN(
        P3_U2822) );
  OAI21_X1 U21694 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18502), .A(
        n18501), .ZN(n18837) );
  NOR2_X1 U21695 ( .A1(n18890), .A2(n19463), .ZN(n18828) );
  AOI221_X1 U21696 ( .B1(n18504), .B2(n9956), .C1(n18503), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18828), .ZN(n18511) );
  AOI21_X1 U21697 ( .B1(n18507), .B2(n18506), .A(n18505), .ZN(n18508) );
  XOR2_X1 U21698 ( .A(n18508), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18833) );
  AOI22_X1 U21699 ( .A1(n18550), .A2(n18833), .B1(n18509), .B2(n18580), .ZN(
        n18510) );
  OAI211_X1 U21700 ( .C1(n18590), .C2(n18837), .A(n18511), .B(n18510), .ZN(
        P3_U2823) );
  NOR2_X1 U21701 ( .A1(n18949), .A2(n18517), .ZN(n18521) );
  OAI21_X1 U21702 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18513), .A(
        n18512), .ZN(n18840) );
  OAI22_X1 U21703 ( .A1(n18591), .A2(n18840), .B1(n18890), .B2(n19461), .ZN(
        n18519) );
  OAI21_X1 U21704 ( .B1(n18516), .B2(n18515), .A(n18514), .ZN(n18845) );
  OAI21_X1 U21705 ( .B1(n18517), .B2(n18949), .A(n18582), .ZN(n18532) );
  OAI22_X1 U21706 ( .A1(n18590), .A2(n18845), .B1(n18520), .B2(n18532), .ZN(
        n18518) );
  AOI211_X1 U21707 ( .C1(n18521), .C2(n18520), .A(n18519), .B(n18518), .ZN(
        n18522) );
  OAI21_X1 U21708 ( .B1(n18571), .B2(n18523), .A(n18522), .ZN(P3_U2824) );
  OAI21_X1 U21709 ( .B1(n18526), .B2(n18525), .A(n18524), .ZN(n18847) );
  AOI21_X1 U21710 ( .B1(n18527), .B2(n18587), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18533) );
  OAI21_X1 U21711 ( .B1(n18530), .B2(n18529), .A(n18528), .ZN(n18531) );
  XOR2_X1 U21712 ( .A(n18531), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18853) );
  OAI22_X1 U21713 ( .A1(n18533), .A2(n18532), .B1(n18590), .B2(n18853), .ZN(
        n18534) );
  AOI21_X1 U21714 ( .B1(n18535), .B2(n18580), .A(n18534), .ZN(n18536) );
  NAND2_X1 U21715 ( .A1(n18902), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18846) );
  OAI211_X1 U21716 ( .C1(n18591), .C2(n18847), .A(n18536), .B(n18846), .ZN(
        P3_U2825) );
  OAI21_X1 U21717 ( .B1(n18539), .B2(n18538), .A(n18537), .ZN(n18863) );
  AOI22_X1 U21718 ( .A1(n18902), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n19302), 
        .B2(n18540), .ZN(n18552) );
  AOI21_X1 U21719 ( .B1(n18543), .B2(n18542), .A(n18541), .ZN(n18544) );
  XOR2_X1 U21720 ( .A(n18544), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18861) );
  AOI21_X1 U21721 ( .B1(n18546), .B2(n18545), .A(n18573), .ZN(n18559) );
  OAI22_X1 U21722 ( .A1(n18571), .A2(n18548), .B1(n18547), .B2(n18559), .ZN(
        n18549) );
  AOI21_X1 U21723 ( .B1(n18550), .B2(n18861), .A(n18549), .ZN(n18551) );
  OAI211_X1 U21724 ( .C1(n18590), .C2(n18863), .A(n18552), .B(n18551), .ZN(
        P3_U2826) );
  OAI21_X1 U21725 ( .B1(n18555), .B2(n18554), .A(n18553), .ZN(n18868) );
  AOI21_X1 U21726 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18587), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18560) );
  OAI21_X1 U21727 ( .B1(n18558), .B2(n18557), .A(n18556), .ZN(n18871) );
  OAI22_X1 U21728 ( .A1(n18560), .A2(n18559), .B1(n18591), .B2(n18871), .ZN(
        n18561) );
  AOI21_X1 U21729 ( .B1(n18562), .B2(n18580), .A(n18561), .ZN(n18563) );
  NAND2_X1 U21730 ( .A1(n18902), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18867) );
  OAI211_X1 U21731 ( .C1(n18590), .C2(n18868), .A(n18563), .B(n18867), .ZN(
        P3_U2827) );
  OAI21_X1 U21732 ( .B1(n18566), .B2(n18565), .A(n18564), .ZN(n18886) );
  OAI21_X1 U21733 ( .B1(n18569), .B2(n18568), .A(n18567), .ZN(n18881) );
  OAI22_X1 U21734 ( .A1(n18571), .A2(n18570), .B1(n18591), .B2(n18881), .ZN(
        n18572) );
  AOI221_X1 U21735 ( .B1(n19302), .B2(n18574), .C1(n18573), .C2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n18572), .ZN(n18575) );
  NAND2_X1 U21736 ( .A1(n18902), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18884) );
  OAI211_X1 U21737 ( .C1(n18590), .C2(n18886), .A(n18575), .B(n18884), .ZN(
        P3_U2828) );
  AOI21_X1 U21738 ( .B1(n18578), .B2(n18585), .A(n18576), .ZN(n18897) );
  OAI21_X1 U21739 ( .B1(n18584), .B2(n18578), .A(n18577), .ZN(n18889) );
  OAI22_X1 U21740 ( .A1(n18590), .A2(n18889), .B1(n18890), .B2(n19452), .ZN(
        n18579) );
  AOI221_X1 U21741 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18582), .C1(
        n18581), .C2(n18580), .A(n18579), .ZN(n18583) );
  OAI21_X1 U21742 ( .B1(n18897), .B2(n18591), .A(n18583), .ZN(P3_U2829) );
  INV_X1 U21743 ( .A(n18584), .ZN(n18586) );
  NAND2_X1 U21744 ( .A1(n18586), .A2(n18585), .ZN(n18905) );
  INV_X1 U21745 ( .A(n18905), .ZN(n18592) );
  NAND3_X1 U21746 ( .A1(n19534), .A2(n19432), .A3(n18587), .ZN(n18588) );
  AOI22_X1 U21747 ( .A1(n18902), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18588), .ZN(n18589) );
  OAI221_X1 U21748 ( .B1(n18592), .B2(n18591), .C1(n18905), .C2(n18590), .A(
        n18589), .ZN(P3_U2830) );
  AOI22_X1 U21749 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18892), .B1(
        n18822), .B2(n18593), .ZN(n18604) );
  INV_X1 U21750 ( .A(n19380), .ZN(n19375) );
  NAND2_X1 U21751 ( .A1(n19375), .A2(n19382), .ZN(n18872) );
  OAI22_X1 U21752 ( .A1(n18595), .A2(n18755), .B1(n18594), .B2(n19360), .ZN(
        n18596) );
  AOI211_X1 U21753 ( .C1(n18598), .C2(n18872), .A(n18597), .B(n18596), .ZN(
        n18600) );
  NAND2_X1 U21754 ( .A1(n19380), .A2(n19551), .ZN(n18874) );
  NAND2_X1 U21755 ( .A1(n18599), .A2(n18874), .ZN(n18688) );
  OAI21_X1 U21756 ( .B1(n18614), .B2(n18688), .A(n18872), .ZN(n18617) );
  NAND2_X1 U21757 ( .A1(n18600), .A2(n18617), .ZN(n18607) );
  OAI21_X1 U21758 ( .B1(n9988), .B2(n18887), .A(n18601), .ZN(n18602) );
  OAI21_X1 U21759 ( .B1(n9988), .B2(n18607), .A(n18602), .ZN(n18603) );
  OAI211_X1 U21760 ( .C1(n19503), .C2(n18890), .A(n18604), .B(n18603), .ZN(
        P3_U2835) );
  AOI21_X1 U21761 ( .B1(n18606), .B2(n18660), .A(n18605), .ZN(n18609) );
  OAI211_X1 U21762 ( .C1(n18887), .C2(n18607), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n18890), .ZN(n18608) );
  OAI211_X1 U21763 ( .C1(n18610), .C2(n18799), .A(n18609), .B(n18608), .ZN(
        P3_U2836) );
  NOR2_X1 U21764 ( .A1(n18890), .A2(n19499), .ZN(n18620) );
  AOI221_X1 U21765 ( .B1(n18614), .B2(n18879), .C1(n18611), .C2(n18879), .A(
        n18612), .ZN(n18618) );
  OAI21_X1 U21766 ( .B1(n18614), .B2(n18613), .A(n18612), .ZN(n18615) );
  INV_X1 U21767 ( .A(n18615), .ZN(n18616) );
  AOI211_X1 U21768 ( .C1(n18618), .C2(n18617), .A(n18616), .B(n18887), .ZN(
        n18619) );
  AOI211_X1 U21769 ( .C1(n18892), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18620), .B(n18619), .ZN(n18624) );
  AOI22_X1 U21770 ( .A1(n18823), .A2(n18622), .B1(n18822), .B2(n18621), .ZN(
        n18623) );
  OAI211_X1 U21771 ( .C1(n18896), .C2(n18625), .A(n18624), .B(n18623), .ZN(
        P3_U2837) );
  AOI22_X1 U21772 ( .A1(n18902), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18660), 
        .B2(n18626), .ZN(n18636) );
  INV_X1 U21773 ( .A(n18755), .ZN(n18780) );
  AOI22_X1 U21774 ( .A1(n18753), .A2(n18628), .B1(n18780), .B2(n18627), .ZN(
        n18630) );
  OAI21_X1 U21775 ( .B1(n18638), .B2(n18688), .A(n18872), .ZN(n18629) );
  NAND3_X1 U21776 ( .A1(n18630), .A2(n18815), .A3(n18629), .ZN(n18634) );
  NOR2_X1 U21777 ( .A1(n18631), .A2(n19397), .ZN(n18651) );
  AOI21_X1 U21778 ( .B1(n18661), .B2(n18685), .A(n19397), .ZN(n18645) );
  NOR4_X1 U21779 ( .A1(n18651), .A2(n18645), .A3(n18632), .A4(n18634), .ZN(
        n18633) );
  NOR2_X1 U21780 ( .A1(n18902), .A2(n18633), .ZN(n18640) );
  OAI211_X1 U21781 ( .C1(n18814), .C2(n18634), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18640), .ZN(n18635) );
  OAI211_X1 U21782 ( .C1(n18637), .C2(n18799), .A(n18636), .B(n18635), .ZN(
        P3_U2838) );
  NOR3_X1 U21783 ( .A1(n18892), .A2(n18639), .A3(n18638), .ZN(n18641) );
  OAI21_X1 U21784 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18641), .A(
        n18640), .ZN(n18642) );
  OAI211_X1 U21785 ( .C1(n18644), .C2(n18799), .A(n18643), .B(n18642), .ZN(
        P3_U2839) );
  AOI22_X1 U21786 ( .A1(n18718), .A2(n18780), .B1(n18717), .B2(n18753), .ZN(
        n18691) );
  INV_X1 U21787 ( .A(n18691), .ZN(n18669) );
  INV_X1 U21788 ( .A(n18670), .ZN(n18646) );
  AOI221_X1 U21789 ( .B1(n18647), .B2(n19371), .C1(n18646), .C2(n19371), .A(
        n18645), .ZN(n18648) );
  OAI221_X1 U21790 ( .B1(n19375), .B2(n18661), .C1(n19375), .C2(n18704), .A(
        n18648), .ZN(n18673) );
  NAND2_X1 U21791 ( .A1(n19360), .A2(n18755), .ZN(n18784) );
  INV_X1 U21792 ( .A(n18784), .ZN(n18671) );
  OAI22_X1 U21793 ( .A1(n19382), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18671), .B2(n18653), .ZN(n18649) );
  NOR3_X1 U21794 ( .A1(n18669), .A2(n18673), .A3(n18649), .ZN(n18663) );
  AOI211_X1 U21795 ( .C1(n18652), .C2(n18872), .A(n18651), .B(n18650), .ZN(
        n18655) );
  AOI22_X1 U21796 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18898), .B1(
        n18660), .B2(n18653), .ZN(n18654) );
  AOI21_X1 U21797 ( .B1(n18663), .B2(n18655), .A(n18654), .ZN(n18656) );
  AOI211_X1 U21798 ( .C1(n18892), .C2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n18657), .B(n18656), .ZN(n18658) );
  OAI21_X1 U21799 ( .B1(n18799), .B2(n18659), .A(n18658), .ZN(P3_U2840) );
  NAND2_X1 U21800 ( .A1(n18661), .A2(n18660), .ZN(n18684) );
  AOI22_X1 U21801 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n18902), .B1(n18822), 
        .B2(n18662), .ZN(n18667) );
  OAI211_X1 U21802 ( .C1(n18888), .C2(n18664), .A(n18898), .B(n18663), .ZN(
        n18665) );
  NAND3_X1 U21803 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18890), .A3(
        n18665), .ZN(n18666) );
  OAI211_X1 U21804 ( .C1(n18684), .C2(n18668), .A(n18667), .B(n18666), .ZN(
        P3_U2841) );
  NAND2_X1 U21805 ( .A1(n18683), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18674) );
  NOR2_X1 U21806 ( .A1(n18892), .A2(n18669), .ZN(n18709) );
  OAI21_X1 U21807 ( .B1(n18671), .B2(n18670), .A(n18709), .ZN(n18672) );
  OAI21_X1 U21808 ( .B1(n18673), .B2(n18672), .A(n18890), .ZN(n18682) );
  OAI21_X1 U21809 ( .B1(n18888), .B2(n18674), .A(n18682), .ZN(n18676) );
  AOI22_X1 U21810 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18676), .B1(
        n18822), .B2(n18675), .ZN(n18678) );
  OAI211_X1 U21811 ( .C1(n18684), .C2(n18679), .A(n18678), .B(n18677), .ZN(
        P3_U2842) );
  AOI22_X1 U21812 ( .A1(n18902), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n18822), 
        .B2(n18680), .ZN(n18681) );
  OAI221_X1 U21813 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18684), 
        .C1(n18683), .C2(n18682), .A(n18681), .ZN(P3_U2843) );
  NOR2_X1 U21814 ( .A1(n18685), .A2(n19397), .ZN(n18687) );
  OAI22_X1 U21815 ( .A1(n18879), .A2(n18784), .B1(n18687), .B2(n18686), .ZN(
        n18690) );
  OAI21_X1 U21816 ( .B1(n18711), .B2(n18688), .A(n18872), .ZN(n18689) );
  NAND4_X1 U21817 ( .A1(n18691), .A2(n18898), .A3(n18690), .A4(n18689), .ZN(
        n18699) );
  OAI221_X1 U21818 ( .B1(n18699), .B2(n18700), .C1(n18699), .C2(n18872), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18697) );
  NAND2_X1 U21819 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18854) );
  OAI22_X1 U21820 ( .A1(n18880), .A2(n19397), .B1(n18854), .B2(n18876), .ZN(
        n18865) );
  NAND2_X1 U21821 ( .A1(n18810), .A2(n18865), .ZN(n18830) );
  NOR2_X1 U21822 ( .A1(n18692), .A2(n18830), .ZN(n18768) );
  OAI21_X1 U21823 ( .B1(n18768), .B2(n18767), .A(n18898), .ZN(n18809) );
  NOR2_X1 U21824 ( .A1(n18693), .A2(n18809), .ZN(n18712) );
  AOI22_X1 U21825 ( .A1(n18822), .A2(n18695), .B1(n18712), .B2(n18694), .ZN(
        n18696) );
  OAI221_X1 U21826 ( .B1(n18902), .B2(n18697), .C1(n18890), .C2(n19485), .A(
        n18696), .ZN(P3_U2844) );
  AOI22_X1 U21827 ( .A1(n18902), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18822), 
        .B2(n18698), .ZN(n18703) );
  NAND3_X1 U21828 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18890), .A3(
        n18699), .ZN(n18702) );
  NAND3_X1 U21829 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18712), .A3(
        n18700), .ZN(n18701) );
  NAND3_X1 U21830 ( .A1(n18703), .A2(n18702), .A3(n18701), .ZN(P3_U2845) );
  AOI21_X1 U21831 ( .B1(n19371), .B2(n18749), .A(n19380), .ZN(n18802) );
  AOI21_X1 U21832 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18802), .A(
        n18704), .ZN(n18706) );
  NAND2_X1 U21833 ( .A1(n18879), .A2(n18705), .ZN(n18731) );
  INV_X1 U21834 ( .A(n18731), .ZN(n18778) );
  AOI211_X1 U21835 ( .C1(n18708), .C2(n18707), .A(n18706), .B(n18778), .ZN(
        n18720) );
  AOI221_X1 U21836 ( .B1(n18710), .B2(n18709), .C1(n18720), .C2(n18709), .A(
        n18902), .ZN(n18713) );
  AOI22_X1 U21837 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18713), .B1(
        n18712), .B2(n18711), .ZN(n18715) );
  OAI211_X1 U21838 ( .C1(n18716), .C2(n18799), .A(n18715), .B(n18714), .ZN(
        P3_U2846) );
  NAND2_X1 U21839 ( .A1(n18753), .A2(n18717), .ZN(n18725) );
  NAND2_X1 U21840 ( .A1(n18780), .A2(n18718), .ZN(n18723) );
  AOI21_X1 U21841 ( .B1(n18719), .B2(n18768), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18721) );
  OAI222_X1 U21842 ( .A1(n18725), .A2(n18724), .B1(n18723), .B2(n18722), .C1(
        n18721), .C2(n18720), .ZN(n18727) );
  AOI22_X1 U21843 ( .A1(n18898), .A2(n18727), .B1(n18822), .B2(n18726), .ZN(
        n18729) );
  OAI211_X1 U21844 ( .C1(n18815), .C2(n18730), .A(n18729), .B(n18728), .ZN(
        P3_U2847) );
  OAI211_X1 U21845 ( .C1(n18733), .C2(n19397), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18731), .ZN(n18736) );
  OAI21_X1 U21846 ( .B1(n18749), .B2(n18732), .A(n19371), .ZN(n18734) );
  NOR2_X1 U21847 ( .A1(n19551), .A2(n18749), .ZN(n18801) );
  NAND2_X1 U21848 ( .A1(n18733), .A2(n18801), .ZN(n18764) );
  NAND2_X1 U21849 ( .A1(n19380), .A2(n18764), .ZN(n18758) );
  OAI211_X1 U21850 ( .C1(n18888), .C2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n18734), .B(n18758), .ZN(n18735) );
  OAI21_X1 U21851 ( .B1(n18736), .B2(n18735), .A(n18898), .ZN(n18739) );
  NAND2_X1 U21852 ( .A1(n18768), .A2(n18737), .ZN(n18738) );
  AOI222_X1 U21853 ( .A1(n18740), .A2(n18739), .B1(n18740), .B2(n18738), .C1(
        n18739), .C2(n18815), .ZN(n18741) );
  AOI21_X1 U21854 ( .B1(n18902), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18741), 
        .ZN(n18745) );
  AOI22_X1 U21855 ( .A1(n18823), .A2(n18743), .B1(n18901), .B2(n18742), .ZN(
        n18744) );
  OAI211_X1 U21856 ( .C1(n18746), .C2(n18799), .A(n18745), .B(n18744), .ZN(
        P3_U2848) );
  AOI22_X1 U21857 ( .A1(n18902), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18822), 
        .B2(n18747), .ZN(n18761) );
  INV_X1 U21858 ( .A(n18748), .ZN(n18785) );
  OAI21_X1 U21859 ( .B1(n18785), .B2(n18749), .A(n19371), .ZN(n18750) );
  OAI21_X1 U21860 ( .B1(n18751), .B2(n19397), .A(n18750), .ZN(n18787) );
  AOI211_X1 U21861 ( .C1(n18753), .C2(n18752), .A(n18778), .B(n18787), .ZN(
        n18754) );
  OAI21_X1 U21862 ( .B1(n18756), .B2(n18755), .A(n18754), .ZN(n18773) );
  AOI21_X1 U21863 ( .B1(n19371), .B2(n18757), .A(n18769), .ZN(n18766) );
  OAI211_X1 U21864 ( .C1(n18794), .C2(n18766), .A(n18898), .B(n18758), .ZN(
        n18759) );
  OAI211_X1 U21865 ( .C1(n18773), .C2(n18759), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18890), .ZN(n18760) );
  OAI211_X1 U21866 ( .C1(n18809), .C2(n18762), .A(n18761), .B(n18760), .ZN(
        P3_U2849) );
  AOI22_X1 U21867 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18892), .B1(
        n18822), .B2(n18763), .ZN(n18776) );
  INV_X1 U21868 ( .A(n18764), .ZN(n18765) );
  AOI21_X1 U21869 ( .B1(n18766), .B2(n19375), .A(n18765), .ZN(n18774) );
  NOR2_X1 U21870 ( .A1(n18768), .A2(n18767), .ZN(n18771) );
  OAI21_X1 U21871 ( .B1(n18771), .B2(n18770), .A(n18769), .ZN(n18772) );
  OAI211_X1 U21872 ( .C1(n18774), .C2(n18773), .A(n18898), .B(n18772), .ZN(
        n18775) );
  OAI211_X1 U21873 ( .C1(n19474), .C2(n18890), .A(n18776), .B(n18775), .ZN(
        P3_U2850) );
  AOI22_X1 U21874 ( .A1(n18902), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18822), 
        .B2(n18777), .ZN(n18789) );
  AOI21_X1 U21875 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18801), .A(
        n19375), .ZN(n18783) );
  AOI211_X1 U21876 ( .C1(n18780), .C2(n18779), .A(n18778), .B(n18887), .ZN(
        n18781) );
  OAI21_X1 U21877 ( .B1(n19360), .B2(n18782), .A(n18781), .ZN(n18804) );
  AOI211_X1 U21878 ( .C1(n18785), .C2(n18784), .A(n18783), .B(n18804), .ZN(
        n18793) );
  OAI21_X1 U21879 ( .B1(n19375), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18793), .ZN(n18786) );
  OAI211_X1 U21880 ( .C1(n18787), .C2(n18786), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18890), .ZN(n18788) );
  OAI211_X1 U21881 ( .C1(n18809), .C2(n18790), .A(n18789), .B(n18788), .ZN(
        P3_U2851) );
  NOR2_X1 U21882 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18809), .ZN(
        n18791) );
  AOI22_X1 U21883 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18791), .B1(
        n18902), .B2(P3_REIP_REG_10__SCAN_IN), .ZN(n18798) );
  NOR2_X1 U21884 ( .A1(n19382), .A2(n18792), .ZN(n18796) );
  OAI21_X1 U21885 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18794), .A(
        n18793), .ZN(n18795) );
  OAI211_X1 U21886 ( .C1(n18796), .C2(n18795), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18890), .ZN(n18797) );
  OAI211_X1 U21887 ( .C1(n18800), .C2(n18799), .A(n18798), .B(n18797), .ZN(
        P3_U2852) );
  NOR2_X1 U21888 ( .A1(n18802), .A2(n18801), .ZN(n18803) );
  OAI21_X1 U21889 ( .B1(n18804), .B2(n18803), .A(n18890), .ZN(n18807) );
  AOI22_X1 U21890 ( .A1(n18902), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18822), 
        .B2(n18805), .ZN(n18806) );
  OAI221_X1 U21891 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18809), .C1(
        n18808), .C2(n18807), .A(n18806), .ZN(P3_U2853) );
  NAND3_X1 U21892 ( .A1(n18810), .A2(n18898), .A3(n18865), .ZN(n18841) );
  NOR3_X1 U21893 ( .A1(n18832), .A2(n18831), .A3(n18841), .ZN(n18820) );
  NAND2_X1 U21894 ( .A1(n18811), .A2(n18872), .ZN(n18812) );
  OAI211_X1 U21895 ( .C1(n18813), .C2(n19397), .A(n18874), .B(n18812), .ZN(
        n18838) );
  AOI211_X1 U21896 ( .C1(n18814), .C2(n18832), .A(n18831), .B(n18838), .ZN(
        n18829) );
  OAI21_X1 U21897 ( .B1(n18829), .B2(n18816), .A(n18815), .ZN(n18818) );
  NOR2_X1 U21898 ( .A1(n18890), .A2(n19465), .ZN(n18817) );
  AOI221_X1 U21899 ( .B1(n18820), .B2(n18819), .C1(n18818), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18817), .ZN(n18826) );
  AOI22_X1 U21900 ( .A1(n18824), .A2(n18823), .B1(n18822), .B2(n18821), .ZN(
        n18825) );
  OAI211_X1 U21901 ( .C1(n18896), .C2(n18827), .A(n18826), .B(n18825), .ZN(
        P3_U2854) );
  AOI21_X1 U21902 ( .B1(n18892), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18828), .ZN(n18836) );
  AOI221_X1 U21903 ( .B1(n18832), .B2(n18831), .C1(n18830), .C2(n18831), .A(
        n18829), .ZN(n18834) );
  AOI22_X1 U21904 ( .A1(n18898), .A2(n18834), .B1(n18901), .B2(n18833), .ZN(
        n18835) );
  OAI211_X1 U21905 ( .C1(n18906), .C2(n18837), .A(n18836), .B(n18835), .ZN(
        P3_U2855) );
  AOI21_X1 U21906 ( .B1(n18838), .B2(n18898), .A(n18892), .ZN(n18839) );
  INV_X1 U21907 ( .A(n18839), .ZN(n18849) );
  NOR2_X1 U21908 ( .A1(n18890), .A2(n19461), .ZN(n18843) );
  OAI22_X1 U21909 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18841), .B1(
        n18840), .B2(n18896), .ZN(n18842) );
  AOI211_X1 U21910 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18849), .A(
        n18843), .B(n18842), .ZN(n18844) );
  OAI21_X1 U21911 ( .B1(n18906), .B2(n18845), .A(n18844), .ZN(P3_U2856) );
  NAND3_X1 U21912 ( .A1(n18898), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18865), .ZN(n18857) );
  NOR2_X1 U21913 ( .A1(n18856), .A2(n18857), .ZN(n18851) );
  OAI21_X1 U21914 ( .B1(n18896), .B2(n18847), .A(n18846), .ZN(n18848) );
  AOI221_X1 U21915 ( .B1(n18851), .B2(n18850), .C1(n18849), .C2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n18848), .ZN(n18852) );
  OAI21_X1 U21916 ( .B1(n18906), .B2(n18853), .A(n18852), .ZN(P3_U2857) );
  NOR2_X1 U21917 ( .A1(n18890), .A2(n19457), .ZN(n18860) );
  AOI22_X1 U21918 ( .A1(n18879), .A2(n18880), .B1(n18854), .B2(n18872), .ZN(
        n18855) );
  NAND3_X1 U21919 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18855), .A3(
        n18874), .ZN(n18864) );
  AOI21_X1 U21920 ( .B1(n18893), .B2(n18864), .A(n18892), .ZN(n18858) );
  AOI22_X1 U21921 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18858), .B1(
        n18857), .B2(n18856), .ZN(n18859) );
  AOI211_X1 U21922 ( .C1(n18861), .C2(n18901), .A(n18860), .B(n18859), .ZN(
        n18862) );
  OAI21_X1 U21923 ( .B1(n18906), .B2(n18863), .A(n18862), .ZN(P3_U2858) );
  OAI211_X1 U21924 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18865), .A(
        n18898), .B(n18864), .ZN(n18866) );
  OAI211_X1 U21925 ( .C1(n18906), .C2(n18868), .A(n18867), .B(n18866), .ZN(
        n18869) );
  AOI21_X1 U21926 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18892), .A(
        n18869), .ZN(n18870) );
  OAI21_X1 U21927 ( .B1(n18896), .B2(n18871), .A(n18870), .ZN(P3_U2859) );
  NOR2_X1 U21928 ( .A1(n19551), .A2(n19535), .ZN(n18873) );
  AOI22_X1 U21929 ( .A1(n18879), .A2(n18873), .B1(n19535), .B2(n18872), .ZN(
        n18875) );
  AOI21_X1 U21930 ( .B1(n18875), .B2(n18874), .A(n9990), .ZN(n18878) );
  NOR3_X1 U21931 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19535), .A3(
        n18876), .ZN(n18877) );
  AOI211_X1 U21932 ( .C1(n18880), .C2(n18879), .A(n18878), .B(n18877), .ZN(
        n18882) );
  OAI22_X1 U21933 ( .A1(n18882), .A2(n18887), .B1(n18896), .B2(n18881), .ZN(
        n18883) );
  AOI21_X1 U21934 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18892), .A(
        n18883), .ZN(n18885) );
  OAI211_X1 U21935 ( .C1(n18906), .C2(n18886), .A(n18885), .B(n18884), .ZN(
        P3_U2860) );
  NOR3_X1 U21936 ( .A1(n18888), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18887), .ZN(n18900) );
  OAI22_X1 U21937 ( .A1(n18890), .A2(n19452), .B1(n18906), .B2(n18889), .ZN(
        n18891) );
  AOI221_X1 U21938 ( .B1(n18892), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18900), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n18891), .ZN(
        n18895) );
  OAI211_X1 U21939 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19371), .A(
        n18893), .B(n19535), .ZN(n18894) );
  OAI211_X1 U21940 ( .C1(n18897), .C2(n18896), .A(n18895), .B(n18894), .ZN(
        P3_U2861) );
  AOI211_X1 U21941 ( .C1(n19382), .C2(n18898), .A(n18902), .B(n19551), .ZN(
        n18899) );
  AOI211_X1 U21942 ( .C1(n18901), .C2(n18905), .A(n18900), .B(n18899), .ZN(
        n18904) );
  NAND2_X1 U21943 ( .A1(n18902), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18903) );
  OAI211_X1 U21944 ( .C1(n18906), .C2(n18905), .A(n18904), .B(n18903), .ZN(
        P3_U2862) );
  OAI211_X1 U21945 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18907), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n19421)
         );
  OAI21_X1 U21946 ( .B1(n18910), .B2(n18908), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18909) );
  OAI221_X1 U21947 ( .B1(n18910), .B2(n19421), .C1(n18910), .C2(n18958), .A(
        n18909), .ZN(P3_U2863) );
  NOR2_X1 U21948 ( .A1(n19403), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19094) );
  INV_X1 U21949 ( .A(n19094), .ZN(n19048) );
  NAND2_X1 U21950 ( .A1(n19403), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19187) );
  INV_X1 U21951 ( .A(n19187), .ZN(n18911) );
  NAND2_X1 U21952 ( .A1(n19265), .A2(n18911), .ZN(n19209) );
  AND2_X1 U21953 ( .A1(n19048), .A2(n19209), .ZN(n18913) );
  OAI22_X1 U21954 ( .A1(n18914), .A2(n18918), .B1(n18913), .B2(n18912), .ZN(
        P3_U2866) );
  NOR2_X1 U21955 ( .A1(n18916), .A2(n18915), .ZN(P3_U2867) );
  NAND2_X1 U21956 ( .A1(n19302), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19269) );
  NAND2_X1 U21957 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18919) );
  NAND2_X1 U21958 ( .A1(n19385), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19163) );
  NOR2_X2 U21959 ( .A1(n18919), .A2(n19163), .ZN(n19293) );
  INV_X1 U21960 ( .A(n19293), .ZN(n18973) );
  NOR2_X1 U21961 ( .A1(n18919), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19301) );
  NAND2_X1 U21962 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19301), .ZN(
        n19355) );
  INV_X1 U21963 ( .A(n19355), .ZN(n19339) );
  NAND2_X1 U21964 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19302), .ZN(n19306) );
  INV_X1 U21965 ( .A(n19306), .ZN(n19262) );
  NOR2_X2 U21966 ( .A1(n19002), .A2(n18917), .ZN(n19297) );
  NOR2_X1 U21967 ( .A1(n18918), .A2(n19093), .ZN(n19300) );
  NAND2_X1 U21968 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19300), .ZN(
        n19000) );
  NOR2_X1 U21969 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19116) );
  NOR2_X1 U21970 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19003) );
  NAND2_X1 U21971 ( .A1(n19116), .A2(n19003), .ZN(n19018) );
  NAND2_X1 U21972 ( .A1(n19000), .A2(n19018), .ZN(n18920) );
  INV_X1 U21973 ( .A(n18920), .ZN(n18978) );
  NOR2_X1 U21974 ( .A1(n19214), .A2(n18978), .ZN(n18952) );
  AOI22_X1 U21975 ( .A1(n19339), .A2(n19262), .B1(n19297), .B2(n18952), .ZN(
        n18925) );
  NAND2_X1 U21976 ( .A1(n19387), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19142) );
  AND2_X1 U21977 ( .A1(n19163), .A2(n19142), .ZN(n19210) );
  NOR2_X1 U21978 ( .A1(n19210), .A2(n18919), .ZN(n19266) );
  AOI21_X1 U21979 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n19002), .ZN(n19263) );
  AOI22_X1 U21980 ( .A1(n19302), .A2(n19266), .B1(n19263), .B2(n18920), .ZN(
        n18955) );
  INV_X1 U21981 ( .A(n19018), .ZN(n19020) );
  NAND2_X1 U21982 ( .A1(n18922), .A2(n18921), .ZN(n18953) );
  NOR2_X2 U21983 ( .A1(n18923), .A2(n18953), .ZN(n19303) );
  AOI22_X1 U21984 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18955), .B1(
        n19020), .B2(n19303), .ZN(n18924) );
  OAI211_X1 U21985 ( .C1(n19269), .C2(n18973), .A(n18925), .B(n18924), .ZN(
        P3_U2868) );
  NAND2_X1 U21986 ( .A1(n18950), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19273) );
  NAND2_X1 U21987 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19302), .ZN(n19312) );
  INV_X1 U21988 ( .A(n19312), .ZN(n19270) );
  INV_X1 U21989 ( .A(n19002), .ZN(n19212) );
  AND2_X1 U21990 ( .A1(n19212), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19307) );
  AOI22_X1 U21991 ( .A1(n19339), .A2(n19270), .B1(n18952), .B2(n19307), .ZN(
        n18928) );
  NOR2_X2 U21992 ( .A1(n18926), .A2(n18953), .ZN(n19309) );
  AOI22_X1 U21993 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18955), .B1(
        n19020), .B2(n19309), .ZN(n18927) );
  OAI211_X1 U21994 ( .C1(n18973), .C2(n19273), .A(n18928), .B(n18927), .ZN(
        P3_U2869) );
  NAND2_X1 U21995 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19302), .ZN(n19245) );
  NAND2_X1 U21996 ( .A1(n18950), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19318) );
  INV_X1 U21997 ( .A(n19318), .ZN(n19242) );
  NOR2_X2 U21998 ( .A1(n19002), .A2(n18929), .ZN(n19313) );
  AOI22_X1 U21999 ( .A1(n19293), .A2(n19242), .B1(n18952), .B2(n19313), .ZN(
        n18932) );
  NOR2_X2 U22000 ( .A1(n18930), .A2(n18953), .ZN(n19315) );
  AOI22_X1 U22001 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18955), .B1(
        n19020), .B2(n19315), .ZN(n18931) );
  OAI211_X1 U22002 ( .C1(n19355), .C2(n19245), .A(n18932), .B(n18931), .ZN(
        P3_U2870) );
  NAND2_X1 U22003 ( .A1(n19302), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19324) );
  NAND2_X1 U22004 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18950), .ZN(n19224) );
  INV_X1 U22005 ( .A(n19224), .ZN(n19320) );
  NOR2_X2 U22006 ( .A1(n19002), .A2(n18933), .ZN(n19319) );
  AOI22_X1 U22007 ( .A1(n19339), .A2(n19320), .B1(n18952), .B2(n19319), .ZN(
        n18936) );
  NOR2_X2 U22008 ( .A1(n18934), .A2(n18953), .ZN(n19321) );
  AOI22_X1 U22009 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18955), .B1(
        n19020), .B2(n19321), .ZN(n18935) );
  OAI211_X1 U22010 ( .C1(n18973), .C2(n19324), .A(n18936), .B(n18935), .ZN(
        P3_U2871) );
  NAND2_X1 U22011 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19302), .ZN(n19282) );
  NAND2_X1 U22012 ( .A1(n18950), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19330) );
  INV_X1 U22013 ( .A(n19330), .ZN(n19278) );
  NOR2_X2 U22014 ( .A1(n19002), .A2(n18937), .ZN(n19325) );
  AOI22_X1 U22015 ( .A1(n19293), .A2(n19278), .B1(n18952), .B2(n19325), .ZN(
        n18940) );
  NOR2_X2 U22016 ( .A1(n18938), .A2(n18953), .ZN(n19327) );
  AOI22_X1 U22017 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18955), .B1(
        n19020), .B2(n19327), .ZN(n18939) );
  OAI211_X1 U22018 ( .C1(n19355), .C2(n19282), .A(n18940), .B(n18939), .ZN(
        P3_U2872) );
  NAND2_X1 U22019 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18950), .ZN(n19286) );
  NAND2_X1 U22020 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18950), .ZN(n19336) );
  INV_X1 U22021 ( .A(n19336), .ZN(n19283) );
  NOR2_X2 U22022 ( .A1(n18941), .A2(n19002), .ZN(n19331) );
  AOI22_X1 U22023 ( .A1(n19339), .A2(n19283), .B1(n18952), .B2(n19331), .ZN(
        n18944) );
  NOR2_X2 U22024 ( .A1(n18942), .A2(n18953), .ZN(n19333) );
  AOI22_X1 U22025 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18955), .B1(
        n19020), .B2(n19333), .ZN(n18943) );
  OAI211_X1 U22026 ( .C1(n18973), .C2(n19286), .A(n18944), .B(n18943), .ZN(
        P3_U2873) );
  NAND2_X1 U22027 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19302), .ZN(n19290) );
  NAND2_X1 U22028 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19302), .ZN(n19344) );
  INV_X1 U22029 ( .A(n19344), .ZN(n19287) );
  NOR2_X2 U22030 ( .A1(n21197), .A2(n19002), .ZN(n19337) );
  AOI22_X1 U22031 ( .A1(n19339), .A2(n19287), .B1(n18952), .B2(n19337), .ZN(
        n18947) );
  NOR2_X2 U22032 ( .A1(n18945), .A2(n18953), .ZN(n19340) );
  AOI22_X1 U22033 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18955), .B1(
        n19020), .B2(n19340), .ZN(n18946) );
  OAI211_X1 U22034 ( .C1(n18973), .C2(n19290), .A(n18947), .B(n18946), .ZN(
        P3_U2874) );
  NOR2_X1 U22035 ( .A1(n18949), .A2(n18948), .ZN(n19348) );
  INV_X1 U22036 ( .A(n19348), .ZN(n19261) );
  NAND2_X1 U22037 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18950), .ZN(n19354) );
  INV_X1 U22038 ( .A(n19354), .ZN(n19255) );
  NOR2_X2 U22039 ( .A1(n18951), .A2(n19002), .ZN(n19346) );
  AOI22_X1 U22040 ( .A1(n19293), .A2(n19255), .B1(n18952), .B2(n19346), .ZN(
        n18957) );
  NOR2_X2 U22041 ( .A1(n18954), .A2(n18953), .ZN(n19349) );
  AOI22_X1 U22042 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18955), .B1(
        n19020), .B2(n19349), .ZN(n18956) );
  OAI211_X1 U22043 ( .C1(n19355), .C2(n19261), .A(n18957), .B(n18956), .ZN(
        P3_U2875) );
  INV_X1 U22044 ( .A(n19003), .ZN(n19001) );
  NAND2_X1 U22045 ( .A1(n19387), .A2(n19422), .ZN(n19139) );
  NOR2_X1 U22046 ( .A1(n19001), .A2(n19139), .ZN(n18974) );
  AOI22_X1 U22047 ( .A1(n19293), .A2(n19262), .B1(n19297), .B2(n18974), .ZN(
        n18960) );
  NAND2_X1 U22048 ( .A1(n19212), .A2(n18958), .ZN(n19140) );
  NOR2_X1 U22049 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19140), .ZN(
        n19046) );
  AOI22_X1 U22050 ( .A1(n19302), .A2(n19300), .B1(n19003), .B2(n19046), .ZN(
        n18975) );
  NOR2_X2 U22051 ( .A1(n19001), .A2(n19142), .ZN(n19042) );
  AOI22_X1 U22052 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18975), .B1(
        n19303), .B2(n19042), .ZN(n18959) );
  OAI211_X1 U22053 ( .C1(n19269), .C2(n19000), .A(n18960), .B(n18959), .ZN(
        P3_U2876) );
  AOI22_X1 U22054 ( .A1(n19293), .A2(n19270), .B1(n19307), .B2(n18974), .ZN(
        n18962) );
  AOI22_X1 U22055 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18975), .B1(
        n19309), .B2(n19042), .ZN(n18961) );
  OAI211_X1 U22056 ( .C1(n19000), .C2(n19273), .A(n18962), .B(n18961), .ZN(
        P3_U2877) );
  INV_X1 U22057 ( .A(n19000), .ZN(n19350) );
  AOI22_X1 U22058 ( .A1(n19350), .A2(n19242), .B1(n19313), .B2(n18974), .ZN(
        n18964) );
  AOI22_X1 U22059 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18975), .B1(
        n19315), .B2(n19042), .ZN(n18963) );
  OAI211_X1 U22060 ( .C1(n18973), .C2(n19245), .A(n18964), .B(n18963), .ZN(
        P3_U2878) );
  INV_X1 U22061 ( .A(n19324), .ZN(n19221) );
  AOI22_X1 U22062 ( .A1(n19350), .A2(n19221), .B1(n19319), .B2(n18974), .ZN(
        n18966) );
  AOI22_X1 U22063 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18975), .B1(
        n19321), .B2(n19042), .ZN(n18965) );
  OAI211_X1 U22064 ( .C1(n18973), .C2(n19224), .A(n18966), .B(n18965), .ZN(
        P3_U2879) );
  AOI22_X1 U22065 ( .A1(n19350), .A2(n19278), .B1(n19325), .B2(n18974), .ZN(
        n18968) );
  AOI22_X1 U22066 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18975), .B1(
        n19327), .B2(n19042), .ZN(n18967) );
  OAI211_X1 U22067 ( .C1(n18973), .C2(n19282), .A(n18968), .B(n18967), .ZN(
        P3_U2880) );
  INV_X1 U22068 ( .A(n19286), .ZN(n19332) );
  AOI22_X1 U22069 ( .A1(n19350), .A2(n19332), .B1(n19331), .B2(n18974), .ZN(
        n18970) );
  AOI22_X1 U22070 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18975), .B1(
        n19333), .B2(n19042), .ZN(n18969) );
  OAI211_X1 U22071 ( .C1(n18973), .C2(n19336), .A(n18970), .B(n18969), .ZN(
        P3_U2881) );
  INV_X1 U22072 ( .A(n19290), .ZN(n19338) );
  AOI22_X1 U22073 ( .A1(n19350), .A2(n19338), .B1(n19337), .B2(n18974), .ZN(
        n18972) );
  AOI22_X1 U22074 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18975), .B1(
        n19340), .B2(n19042), .ZN(n18971) );
  OAI211_X1 U22075 ( .C1(n18973), .C2(n19344), .A(n18972), .B(n18971), .ZN(
        P3_U2882) );
  AOI22_X1 U22076 ( .A1(n19293), .A2(n19348), .B1(n19346), .B2(n18974), .ZN(
        n18977) );
  AOI22_X1 U22077 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18975), .B1(
        n19349), .B2(n19042), .ZN(n18976) );
  OAI211_X1 U22078 ( .C1(n19000), .C2(n19354), .A(n18977), .B(n18976), .ZN(
        P3_U2883) );
  NOR2_X2 U22079 ( .A1(n19163), .A2(n19001), .ZN(n19065) );
  NOR2_X1 U22080 ( .A1(n19042), .A2(n19065), .ZN(n19024) );
  OAI21_X1 U22081 ( .B1(n19164), .B2(n18978), .A(n19024), .ZN(n18979) );
  OAI211_X1 U22082 ( .C1(n19524), .C2(n19065), .A(n18979), .B(n19212), .ZN(
        n18997) );
  INV_X1 U22083 ( .A(n18997), .ZN(n18985) );
  INV_X1 U22084 ( .A(n19269), .ZN(n19298) );
  NOR2_X1 U22085 ( .A1(n19214), .A2(n19024), .ZN(n18996) );
  AOI22_X1 U22086 ( .A1(n19298), .A2(n19020), .B1(n19297), .B2(n18996), .ZN(
        n18981) );
  AOI22_X1 U22087 ( .A1(n19350), .A2(n19262), .B1(n19303), .B2(n19065), .ZN(
        n18980) );
  OAI211_X1 U22088 ( .C1(n18985), .C2(n21156), .A(n18981), .B(n18980), .ZN(
        P3_U2884) );
  INV_X1 U22089 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18984) );
  INV_X1 U22090 ( .A(n19273), .ZN(n19308) );
  AOI22_X1 U22091 ( .A1(n19020), .A2(n19308), .B1(n19307), .B2(n18996), .ZN(
        n18983) );
  AOI22_X1 U22092 ( .A1(n19350), .A2(n19270), .B1(n19309), .B2(n19065), .ZN(
        n18982) );
  OAI211_X1 U22093 ( .C1(n18985), .C2(n18984), .A(n18983), .B(n18982), .ZN(
        P3_U2885) );
  AOI22_X1 U22094 ( .A1(n19020), .A2(n19242), .B1(n19313), .B2(n18996), .ZN(
        n18987) );
  AOI22_X1 U22095 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18997), .B1(
        n19315), .B2(n19065), .ZN(n18986) );
  OAI211_X1 U22096 ( .C1(n19000), .C2(n19245), .A(n18987), .B(n18986), .ZN(
        P3_U2886) );
  AOI22_X1 U22097 ( .A1(n19350), .A2(n19320), .B1(n19319), .B2(n18996), .ZN(
        n18989) );
  AOI22_X1 U22098 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18997), .B1(
        n19321), .B2(n19065), .ZN(n18988) );
  OAI211_X1 U22099 ( .C1(n19018), .C2(n19324), .A(n18989), .B(n18988), .ZN(
        P3_U2887) );
  AOI22_X1 U22100 ( .A1(n19020), .A2(n19278), .B1(n19325), .B2(n18996), .ZN(
        n18991) );
  AOI22_X1 U22101 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18997), .B1(
        n19327), .B2(n19065), .ZN(n18990) );
  OAI211_X1 U22102 ( .C1(n19000), .C2(n19282), .A(n18991), .B(n18990), .ZN(
        P3_U2888) );
  AOI22_X1 U22103 ( .A1(n19020), .A2(n19332), .B1(n19331), .B2(n18996), .ZN(
        n18993) );
  AOI22_X1 U22104 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18997), .B1(
        n19333), .B2(n19065), .ZN(n18992) );
  OAI211_X1 U22105 ( .C1(n19000), .C2(n19336), .A(n18993), .B(n18992), .ZN(
        P3_U2889) );
  AOI22_X1 U22106 ( .A1(n19350), .A2(n19287), .B1(n19337), .B2(n18996), .ZN(
        n18995) );
  AOI22_X1 U22107 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18997), .B1(
        n19340), .B2(n19065), .ZN(n18994) );
  OAI211_X1 U22108 ( .C1(n19018), .C2(n19290), .A(n18995), .B(n18994), .ZN(
        P3_U2890) );
  AOI22_X1 U22109 ( .A1(n19020), .A2(n19255), .B1(n19346), .B2(n18996), .ZN(
        n18999) );
  AOI22_X1 U22110 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18997), .B1(
        n19349), .B2(n19065), .ZN(n18998) );
  OAI211_X1 U22111 ( .C1(n19000), .C2(n19261), .A(n18999), .B(n18998), .ZN(
        P3_U2891) );
  NOR2_X1 U22112 ( .A1(n19387), .A2(n19001), .ZN(n19047) );
  AND2_X1 U22113 ( .A1(n19422), .A2(n19047), .ZN(n19019) );
  AOI22_X1 U22114 ( .A1(n19298), .A2(n19042), .B1(n19297), .B2(n19019), .ZN(
        n19005) );
  NAND2_X1 U22115 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19047), .ZN(
        n19069) );
  AOI21_X1 U22116 ( .B1(n19387), .B2(n19164), .A(n19002), .ZN(n19095) );
  OAI211_X1 U22117 ( .C1(n19089), .C2(n19524), .A(n19003), .B(n19095), .ZN(
        n19021) );
  AOI22_X1 U22118 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19021), .B1(
        n19303), .B2(n19089), .ZN(n19004) );
  OAI211_X1 U22119 ( .C1(n19018), .C2(n19306), .A(n19005), .B(n19004), .ZN(
        P3_U2892) );
  INV_X1 U22120 ( .A(n19042), .ZN(n19040) );
  AOI22_X1 U22121 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19021), .B1(
        n19307), .B2(n19019), .ZN(n19007) );
  AOI22_X1 U22122 ( .A1(n19020), .A2(n19270), .B1(n19309), .B2(n19089), .ZN(
        n19006) );
  OAI211_X1 U22123 ( .C1(n19273), .C2(n19040), .A(n19007), .B(n19006), .ZN(
        P3_U2893) );
  AOI22_X1 U22124 ( .A1(n19242), .A2(n19042), .B1(n19313), .B2(n19019), .ZN(
        n19009) );
  AOI22_X1 U22125 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19021), .B1(
        n19315), .B2(n19089), .ZN(n19008) );
  OAI211_X1 U22126 ( .C1(n19018), .C2(n19245), .A(n19009), .B(n19008), .ZN(
        P3_U2894) );
  AOI22_X1 U22127 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19021), .B1(
        n19319), .B2(n19019), .ZN(n19011) );
  AOI22_X1 U22128 ( .A1(n19221), .A2(n19042), .B1(n19321), .B2(n19089), .ZN(
        n19010) );
  OAI211_X1 U22129 ( .C1(n19018), .C2(n19224), .A(n19011), .B(n19010), .ZN(
        P3_U2895) );
  AOI22_X1 U22130 ( .A1(n19278), .A2(n19042), .B1(n19325), .B2(n19019), .ZN(
        n19013) );
  AOI22_X1 U22131 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19021), .B1(
        n19327), .B2(n19089), .ZN(n19012) );
  OAI211_X1 U22132 ( .C1(n19018), .C2(n19282), .A(n19013), .B(n19012), .ZN(
        P3_U2896) );
  AOI22_X1 U22133 ( .A1(n19332), .A2(n19042), .B1(n19331), .B2(n19019), .ZN(
        n19015) );
  AOI22_X1 U22134 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19021), .B1(
        n19333), .B2(n19089), .ZN(n19014) );
  OAI211_X1 U22135 ( .C1(n19018), .C2(n19336), .A(n19015), .B(n19014), .ZN(
        P3_U2897) );
  AOI22_X1 U22136 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19021), .B1(
        n19337), .B2(n19019), .ZN(n19017) );
  AOI22_X1 U22137 ( .A1(n19338), .A2(n19042), .B1(n19340), .B2(n19089), .ZN(
        n19016) );
  OAI211_X1 U22138 ( .C1(n19018), .C2(n19344), .A(n19017), .B(n19016), .ZN(
        P3_U2898) );
  AOI22_X1 U22139 ( .A1(n19020), .A2(n19348), .B1(n19346), .B2(n19019), .ZN(
        n19023) );
  AOI22_X1 U22140 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19021), .B1(
        n19349), .B2(n19089), .ZN(n19022) );
  OAI211_X1 U22141 ( .C1(n19354), .C2(n19040), .A(n19023), .B(n19022), .ZN(
        P3_U2899) );
  NAND2_X1 U22142 ( .A1(n19116), .A2(n19094), .ZN(n19115) );
  INV_X1 U22143 ( .A(n19115), .ZN(n19108) );
  NOR2_X1 U22144 ( .A1(n19089), .A2(n19108), .ZN(n19072) );
  NOR2_X1 U22145 ( .A1(n19214), .A2(n19072), .ZN(n19041) );
  AOI22_X1 U22146 ( .A1(n19298), .A2(n19065), .B1(n19297), .B2(n19041), .ZN(
        n19027) );
  OAI21_X1 U22147 ( .B1(n19024), .B2(n19164), .A(n19072), .ZN(n19025) );
  OAI211_X1 U22148 ( .C1(n19108), .C2(n19524), .A(n19212), .B(n19025), .ZN(
        n19043) );
  AOI22_X1 U22149 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19043), .B1(
        n19303), .B2(n19108), .ZN(n19026) );
  OAI211_X1 U22150 ( .C1(n19306), .C2(n19040), .A(n19027), .B(n19026), .ZN(
        P3_U2900) );
  AOI22_X1 U22151 ( .A1(n19308), .A2(n19065), .B1(n19307), .B2(n19041), .ZN(
        n19029) );
  AOI22_X1 U22152 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19043), .B1(
        n19309), .B2(n19108), .ZN(n19028) );
  OAI211_X1 U22153 ( .C1(n19312), .C2(n19040), .A(n19029), .B(n19028), .ZN(
        P3_U2901) );
  AOI22_X1 U22154 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19043), .B1(
        n19313), .B2(n19041), .ZN(n19031) );
  AOI22_X1 U22155 ( .A1(n19315), .A2(n19108), .B1(n19242), .B2(n19065), .ZN(
        n19030) );
  OAI211_X1 U22156 ( .C1(n19245), .C2(n19040), .A(n19031), .B(n19030), .ZN(
        P3_U2902) );
  INV_X1 U22157 ( .A(n19065), .ZN(n19063) );
  AOI22_X1 U22158 ( .A1(n19320), .A2(n19042), .B1(n19319), .B2(n19041), .ZN(
        n19033) );
  AOI22_X1 U22159 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19043), .B1(
        n19321), .B2(n19108), .ZN(n19032) );
  OAI211_X1 U22160 ( .C1(n19324), .C2(n19063), .A(n19033), .B(n19032), .ZN(
        P3_U2903) );
  AOI22_X1 U22161 ( .A1(n19278), .A2(n19065), .B1(n19325), .B2(n19041), .ZN(
        n19035) );
  AOI22_X1 U22162 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19043), .B1(
        n19327), .B2(n19108), .ZN(n19034) );
  OAI211_X1 U22163 ( .C1(n19282), .C2(n19040), .A(n19035), .B(n19034), .ZN(
        P3_U2904) );
  AOI22_X1 U22164 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19043), .B1(
        n19331), .B2(n19041), .ZN(n19037) );
  AOI22_X1 U22165 ( .A1(n19333), .A2(n19108), .B1(n19283), .B2(n19042), .ZN(
        n19036) );
  OAI211_X1 U22166 ( .C1(n19286), .C2(n19063), .A(n19037), .B(n19036), .ZN(
        P3_U2905) );
  AOI22_X1 U22167 ( .A1(n19338), .A2(n19065), .B1(n19337), .B2(n19041), .ZN(
        n19039) );
  AOI22_X1 U22168 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19043), .B1(
        n19340), .B2(n19108), .ZN(n19038) );
  OAI211_X1 U22169 ( .C1(n19344), .C2(n19040), .A(n19039), .B(n19038), .ZN(
        P3_U2906) );
  AOI22_X1 U22170 ( .A1(n19348), .A2(n19042), .B1(n19346), .B2(n19041), .ZN(
        n19045) );
  AOI22_X1 U22171 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19043), .B1(
        n19349), .B2(n19108), .ZN(n19044) );
  OAI211_X1 U22172 ( .C1(n19354), .C2(n19063), .A(n19045), .B(n19044), .ZN(
        P3_U2907) );
  NOR2_X1 U22173 ( .A1(n19139), .A2(n19048), .ZN(n19064) );
  AOI22_X1 U22174 ( .A1(n19298), .A2(n19089), .B1(n19297), .B2(n19064), .ZN(
        n19050) );
  AOI22_X1 U22175 ( .A1(n19302), .A2(n19047), .B1(n19046), .B2(n19094), .ZN(
        n19066) );
  NOR2_X2 U22176 ( .A1(n19142), .A2(n19048), .ZN(n19135) );
  AOI22_X1 U22177 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19066), .B1(
        n19303), .B2(n19135), .ZN(n19049) );
  OAI211_X1 U22178 ( .C1(n19306), .C2(n19063), .A(n19050), .B(n19049), .ZN(
        P3_U2908) );
  AOI22_X1 U22179 ( .A1(n19308), .A2(n19089), .B1(n19307), .B2(n19064), .ZN(
        n19052) );
  AOI22_X1 U22180 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19066), .B1(
        n19309), .B2(n19135), .ZN(n19051) );
  OAI211_X1 U22181 ( .C1(n19312), .C2(n19063), .A(n19052), .B(n19051), .ZN(
        P3_U2909) );
  AOI22_X1 U22182 ( .A1(n19242), .A2(n19089), .B1(n19313), .B2(n19064), .ZN(
        n19054) );
  AOI22_X1 U22183 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19066), .B1(
        n19315), .B2(n19135), .ZN(n19053) );
  OAI211_X1 U22184 ( .C1(n19245), .C2(n19063), .A(n19054), .B(n19053), .ZN(
        P3_U2910) );
  AOI22_X1 U22185 ( .A1(n19221), .A2(n19089), .B1(n19319), .B2(n19064), .ZN(
        n19056) );
  AOI22_X1 U22186 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19066), .B1(
        n19321), .B2(n19135), .ZN(n19055) );
  OAI211_X1 U22187 ( .C1(n19224), .C2(n19063), .A(n19056), .B(n19055), .ZN(
        P3_U2911) );
  INV_X1 U22188 ( .A(n19282), .ZN(n19326) );
  AOI22_X1 U22189 ( .A1(n19326), .A2(n19065), .B1(n19325), .B2(n19064), .ZN(
        n19058) );
  AOI22_X1 U22190 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19066), .B1(
        n19327), .B2(n19135), .ZN(n19057) );
  OAI211_X1 U22191 ( .C1(n19330), .C2(n19069), .A(n19058), .B(n19057), .ZN(
        P3_U2912) );
  AOI22_X1 U22192 ( .A1(n19332), .A2(n19089), .B1(n19331), .B2(n19064), .ZN(
        n19060) );
  AOI22_X1 U22193 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19066), .B1(
        n19333), .B2(n19135), .ZN(n19059) );
  OAI211_X1 U22194 ( .C1(n19336), .C2(n19063), .A(n19060), .B(n19059), .ZN(
        P3_U2913) );
  AOI22_X1 U22195 ( .A1(n19338), .A2(n19089), .B1(n19337), .B2(n19064), .ZN(
        n19062) );
  AOI22_X1 U22196 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19066), .B1(
        n19340), .B2(n19135), .ZN(n19061) );
  OAI211_X1 U22197 ( .C1(n19344), .C2(n19063), .A(n19062), .B(n19061), .ZN(
        P3_U2914) );
  AOI22_X1 U22198 ( .A1(n19348), .A2(n19065), .B1(n19346), .B2(n19064), .ZN(
        n19068) );
  AOI22_X1 U22199 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19066), .B1(
        n19349), .B2(n19135), .ZN(n19067) );
  OAI211_X1 U22200 ( .C1(n19354), .C2(n19069), .A(n19068), .B(n19067), .ZN(
        P3_U2915) );
  INV_X1 U22201 ( .A(n19135), .ZN(n19131) );
  INV_X1 U22202 ( .A(n19163), .ZN(n19070) );
  NAND2_X1 U22203 ( .A1(n19070), .A2(n19094), .ZN(n19157) );
  NAND2_X1 U22204 ( .A1(n19131), .A2(n19157), .ZN(n19117) );
  INV_X1 U22205 ( .A(n19117), .ZN(n19071) );
  NOR2_X1 U22206 ( .A1(n19214), .A2(n19071), .ZN(n19088) );
  AOI22_X1 U22207 ( .A1(n19262), .A2(n19089), .B1(n19297), .B2(n19088), .ZN(
        n19075) );
  OAI21_X1 U22208 ( .B1(n19072), .B2(n19164), .A(n19071), .ZN(n19073) );
  OAI211_X1 U22209 ( .C1(n19159), .C2(n19524), .A(n19212), .B(n19073), .ZN(
        n19090) );
  AOI22_X1 U22210 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19090), .B1(
        n19303), .B2(n19159), .ZN(n19074) );
  OAI211_X1 U22211 ( .C1(n19269), .C2(n19115), .A(n19075), .B(n19074), .ZN(
        P3_U2916) );
  AOI22_X1 U22212 ( .A1(n19270), .A2(n19089), .B1(n19307), .B2(n19088), .ZN(
        n19077) );
  AOI22_X1 U22213 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19090), .B1(
        n19309), .B2(n19159), .ZN(n19076) );
  OAI211_X1 U22214 ( .C1(n19273), .C2(n19115), .A(n19077), .B(n19076), .ZN(
        P3_U2917) );
  INV_X1 U22215 ( .A(n19245), .ZN(n19314) );
  AOI22_X1 U22216 ( .A1(n19314), .A2(n19089), .B1(n19313), .B2(n19088), .ZN(
        n19079) );
  AOI22_X1 U22217 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19090), .B1(
        n19315), .B2(n19159), .ZN(n19078) );
  OAI211_X1 U22218 ( .C1(n19318), .C2(n19115), .A(n19079), .B(n19078), .ZN(
        P3_U2918) );
  AOI22_X1 U22219 ( .A1(n19320), .A2(n19089), .B1(n19319), .B2(n19088), .ZN(
        n19081) );
  AOI22_X1 U22220 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19090), .B1(
        n19321), .B2(n19159), .ZN(n19080) );
  OAI211_X1 U22221 ( .C1(n19324), .C2(n19115), .A(n19081), .B(n19080), .ZN(
        P3_U2919) );
  AOI22_X1 U22222 ( .A1(n19326), .A2(n19089), .B1(n19325), .B2(n19088), .ZN(
        n19083) );
  AOI22_X1 U22223 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19090), .B1(
        n19327), .B2(n19159), .ZN(n19082) );
  OAI211_X1 U22224 ( .C1(n19330), .C2(n19115), .A(n19083), .B(n19082), .ZN(
        P3_U2920) );
  AOI22_X1 U22225 ( .A1(n19283), .A2(n19089), .B1(n19331), .B2(n19088), .ZN(
        n19085) );
  AOI22_X1 U22226 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19090), .B1(
        n19333), .B2(n19159), .ZN(n19084) );
  OAI211_X1 U22227 ( .C1(n19286), .C2(n19115), .A(n19085), .B(n19084), .ZN(
        P3_U2921) );
  AOI22_X1 U22228 ( .A1(n19287), .A2(n19089), .B1(n19337), .B2(n19088), .ZN(
        n19087) );
  AOI22_X1 U22229 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19090), .B1(
        n19340), .B2(n19159), .ZN(n19086) );
  OAI211_X1 U22230 ( .C1(n19290), .C2(n19115), .A(n19087), .B(n19086), .ZN(
        P3_U2922) );
  AOI22_X1 U22231 ( .A1(n19348), .A2(n19089), .B1(n19346), .B2(n19088), .ZN(
        n19092) );
  AOI22_X1 U22232 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19090), .B1(
        n19349), .B2(n19159), .ZN(n19091) );
  OAI211_X1 U22233 ( .C1(n19354), .C2(n19115), .A(n19092), .B(n19091), .ZN(
        P3_U2923) );
  NOR2_X1 U22234 ( .A1(n19093), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19141) );
  AND2_X1 U22235 ( .A1(n19422), .A2(n19141), .ZN(n19111) );
  AOI22_X1 U22236 ( .A1(n19298), .A2(n19135), .B1(n19297), .B2(n19111), .ZN(
        n19097) );
  NAND2_X1 U22237 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19141), .ZN(
        n19186) );
  INV_X1 U22238 ( .A(n19186), .ZN(n19179) );
  OAI211_X1 U22239 ( .C1(n19179), .C2(n19524), .A(n19095), .B(n19094), .ZN(
        n19112) );
  AOI22_X1 U22240 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19112), .B1(
        n19303), .B2(n19179), .ZN(n19096) );
  OAI211_X1 U22241 ( .C1(n19306), .C2(n19115), .A(n19097), .B(n19096), .ZN(
        P3_U2924) );
  AOI22_X1 U22242 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19112), .B1(
        n19307), .B2(n19111), .ZN(n19099) );
  AOI22_X1 U22243 ( .A1(n19308), .A2(n19135), .B1(n19309), .B2(n19179), .ZN(
        n19098) );
  OAI211_X1 U22244 ( .C1(n19312), .C2(n19115), .A(n19099), .B(n19098), .ZN(
        P3_U2925) );
  AOI22_X1 U22245 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19112), .B1(
        n19313), .B2(n19111), .ZN(n19101) );
  AOI22_X1 U22246 ( .A1(n19315), .A2(n19179), .B1(n19242), .B2(n19135), .ZN(
        n19100) );
  OAI211_X1 U22247 ( .C1(n19245), .C2(n19115), .A(n19101), .B(n19100), .ZN(
        P3_U2926) );
  AOI22_X1 U22248 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19112), .B1(
        n19319), .B2(n19111), .ZN(n19103) );
  AOI22_X1 U22249 ( .A1(n19221), .A2(n19135), .B1(n19321), .B2(n19179), .ZN(
        n19102) );
  OAI211_X1 U22250 ( .C1(n19224), .C2(n19115), .A(n19103), .B(n19102), .ZN(
        P3_U2927) );
  AOI22_X1 U22251 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19112), .B1(
        n19325), .B2(n19111), .ZN(n19105) );
  AOI22_X1 U22252 ( .A1(n19327), .A2(n19179), .B1(n19278), .B2(n19135), .ZN(
        n19104) );
  OAI211_X1 U22253 ( .C1(n19282), .C2(n19115), .A(n19105), .B(n19104), .ZN(
        P3_U2928) );
  AOI22_X1 U22254 ( .A1(n19332), .A2(n19135), .B1(n19331), .B2(n19111), .ZN(
        n19107) );
  AOI22_X1 U22255 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19112), .B1(
        n19333), .B2(n19179), .ZN(n19106) );
  OAI211_X1 U22256 ( .C1(n19336), .C2(n19115), .A(n19107), .B(n19106), .ZN(
        P3_U2929) );
  AOI22_X1 U22257 ( .A1(n19287), .A2(n19108), .B1(n19337), .B2(n19111), .ZN(
        n19110) );
  AOI22_X1 U22258 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19112), .B1(
        n19340), .B2(n19179), .ZN(n19109) );
  OAI211_X1 U22259 ( .C1(n19290), .C2(n19131), .A(n19110), .B(n19109), .ZN(
        P3_U2930) );
  AOI22_X1 U22260 ( .A1(n19346), .A2(n19111), .B1(n19255), .B2(n19135), .ZN(
        n19114) );
  AOI22_X1 U22261 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19112), .B1(
        n19349), .B2(n19179), .ZN(n19113) );
  OAI211_X1 U22262 ( .C1(n19261), .C2(n19115), .A(n19114), .B(n19113), .ZN(
        P3_U2931) );
  INV_X1 U22263 ( .A(n19116), .ZN(n19388) );
  NOR2_X2 U22264 ( .A1(n19388), .A2(n19187), .ZN(n19205) );
  NOR2_X1 U22265 ( .A1(n19179), .A2(n19205), .ZN(n19165) );
  INV_X1 U22266 ( .A(n19165), .ZN(n19118) );
  OAI221_X1 U22267 ( .B1(n19118), .B2(n19265), .C1(n19118), .C2(n19117), .A(
        n19263), .ZN(n19136) );
  NOR2_X1 U22268 ( .A1(n19214), .A2(n19165), .ZN(n19134) );
  AOI22_X1 U22269 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19136), .B1(
        n19297), .B2(n19134), .ZN(n19120) );
  AOI22_X1 U22270 ( .A1(n19298), .A2(n19159), .B1(n19303), .B2(n19205), .ZN(
        n19119) );
  OAI211_X1 U22271 ( .C1(n19306), .C2(n19131), .A(n19120), .B(n19119), .ZN(
        P3_U2932) );
  AOI22_X1 U22272 ( .A1(n19308), .A2(n19159), .B1(n19307), .B2(n19134), .ZN(
        n19122) );
  AOI22_X1 U22273 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19136), .B1(
        n19309), .B2(n19205), .ZN(n19121) );
  OAI211_X1 U22274 ( .C1(n19312), .C2(n19131), .A(n19122), .B(n19121), .ZN(
        P3_U2933) );
  AOI22_X1 U22275 ( .A1(n19242), .A2(n19159), .B1(n19313), .B2(n19134), .ZN(
        n19124) );
  AOI22_X1 U22276 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19136), .B1(
        n19315), .B2(n19205), .ZN(n19123) );
  OAI211_X1 U22277 ( .C1(n19245), .C2(n19131), .A(n19124), .B(n19123), .ZN(
        P3_U2934) );
  AOI22_X1 U22278 ( .A1(n19320), .A2(n19135), .B1(n19319), .B2(n19134), .ZN(
        n19126) );
  AOI22_X1 U22279 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19136), .B1(
        n19321), .B2(n19205), .ZN(n19125) );
  OAI211_X1 U22280 ( .C1(n19324), .C2(n19157), .A(n19126), .B(n19125), .ZN(
        P3_U2935) );
  AOI22_X1 U22281 ( .A1(n19326), .A2(n19135), .B1(n19325), .B2(n19134), .ZN(
        n19128) );
  AOI22_X1 U22282 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19136), .B1(
        n19327), .B2(n19205), .ZN(n19127) );
  OAI211_X1 U22283 ( .C1(n19330), .C2(n19157), .A(n19128), .B(n19127), .ZN(
        P3_U2936) );
  AOI22_X1 U22284 ( .A1(n19332), .A2(n19159), .B1(n19331), .B2(n19134), .ZN(
        n19130) );
  AOI22_X1 U22285 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19136), .B1(
        n19333), .B2(n19205), .ZN(n19129) );
  OAI211_X1 U22286 ( .C1(n19336), .C2(n19131), .A(n19130), .B(n19129), .ZN(
        P3_U2937) );
  AOI22_X1 U22287 ( .A1(n19287), .A2(n19135), .B1(n19337), .B2(n19134), .ZN(
        n19133) );
  AOI22_X1 U22288 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19136), .B1(
        n19340), .B2(n19205), .ZN(n19132) );
  OAI211_X1 U22289 ( .C1(n19290), .C2(n19157), .A(n19133), .B(n19132), .ZN(
        P3_U2938) );
  AOI22_X1 U22290 ( .A1(n19348), .A2(n19135), .B1(n19346), .B2(n19134), .ZN(
        n19138) );
  AOI22_X1 U22291 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19136), .B1(
        n19349), .B2(n19205), .ZN(n19137) );
  OAI211_X1 U22292 ( .C1(n19354), .C2(n19157), .A(n19138), .B(n19137), .ZN(
        P3_U2939) );
  NOR2_X1 U22293 ( .A1(n19139), .A2(n19187), .ZN(n19158) );
  AOI22_X1 U22294 ( .A1(n19262), .A2(n19159), .B1(n19297), .B2(n19158), .ZN(
        n19144) );
  INV_X1 U22295 ( .A(n19140), .ZN(n19299) );
  NOR2_X1 U22296 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19187), .ZN(
        n19188) );
  AOI22_X1 U22297 ( .A1(n19302), .A2(n19141), .B1(n19299), .B2(n19188), .ZN(
        n19160) );
  NOR2_X2 U22298 ( .A1(n19142), .A2(n19187), .ZN(n19233) );
  AOI22_X1 U22299 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19160), .B1(
        n19303), .B2(n19233), .ZN(n19143) );
  OAI211_X1 U22300 ( .C1(n19269), .C2(n19186), .A(n19144), .B(n19143), .ZN(
        P3_U2940) );
  AOI22_X1 U22301 ( .A1(n19270), .A2(n19159), .B1(n19307), .B2(n19158), .ZN(
        n19146) );
  AOI22_X1 U22302 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19160), .B1(
        n19309), .B2(n19233), .ZN(n19145) );
  OAI211_X1 U22303 ( .C1(n19273), .C2(n19186), .A(n19146), .B(n19145), .ZN(
        P3_U2941) );
  AOI22_X1 U22304 ( .A1(n19242), .A2(n19179), .B1(n19313), .B2(n19158), .ZN(
        n19148) );
  AOI22_X1 U22305 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19160), .B1(
        n19315), .B2(n19233), .ZN(n19147) );
  OAI211_X1 U22306 ( .C1(n19245), .C2(n19157), .A(n19148), .B(n19147), .ZN(
        P3_U2942) );
  AOI22_X1 U22307 ( .A1(n19221), .A2(n19179), .B1(n19319), .B2(n19158), .ZN(
        n19150) );
  AOI22_X1 U22308 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19160), .B1(
        n19321), .B2(n19233), .ZN(n19149) );
  OAI211_X1 U22309 ( .C1(n19224), .C2(n19157), .A(n19150), .B(n19149), .ZN(
        P3_U2943) );
  AOI22_X1 U22310 ( .A1(n19326), .A2(n19159), .B1(n19325), .B2(n19158), .ZN(
        n19152) );
  AOI22_X1 U22311 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19160), .B1(
        n19327), .B2(n19233), .ZN(n19151) );
  OAI211_X1 U22312 ( .C1(n19330), .C2(n19186), .A(n19152), .B(n19151), .ZN(
        P3_U2944) );
  AOI22_X1 U22313 ( .A1(n19283), .A2(n19159), .B1(n19331), .B2(n19158), .ZN(
        n19154) );
  AOI22_X1 U22314 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19160), .B1(
        n19333), .B2(n19233), .ZN(n19153) );
  OAI211_X1 U22315 ( .C1(n19286), .C2(n19186), .A(n19154), .B(n19153), .ZN(
        P3_U2945) );
  AOI22_X1 U22316 ( .A1(n19338), .A2(n19179), .B1(n19337), .B2(n19158), .ZN(
        n19156) );
  AOI22_X1 U22317 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19160), .B1(
        n19340), .B2(n19233), .ZN(n19155) );
  OAI211_X1 U22318 ( .C1(n19344), .C2(n19157), .A(n19156), .B(n19155), .ZN(
        P3_U2946) );
  AOI22_X1 U22319 ( .A1(n19348), .A2(n19159), .B1(n19346), .B2(n19158), .ZN(
        n19162) );
  AOI22_X1 U22320 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19160), .B1(
        n19349), .B2(n19233), .ZN(n19161) );
  OAI211_X1 U22321 ( .C1(n19354), .C2(n19186), .A(n19162), .B(n19161), .ZN(
        P3_U2947) );
  INV_X1 U22322 ( .A(n19205), .ZN(n19199) );
  NOR2_X2 U22323 ( .A1(n19163), .A2(n19187), .ZN(n19246) );
  INV_X1 U22324 ( .A(n19246), .ZN(n19260) );
  AOI21_X1 U22325 ( .B1(n19231), .B2(n19260), .A(n19214), .ZN(n19182) );
  AOI22_X1 U22326 ( .A1(n19262), .A2(n19179), .B1(n19297), .B2(n19182), .ZN(
        n19168) );
  OAI211_X1 U22327 ( .C1(n19165), .C2(n19164), .A(n19231), .B(n19260), .ZN(
        n19166) );
  OAI211_X1 U22328 ( .C1(n19246), .C2(n19524), .A(n19212), .B(n19166), .ZN(
        n19183) );
  AOI22_X1 U22329 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19183), .B1(
        n19303), .B2(n19246), .ZN(n19167) );
  OAI211_X1 U22330 ( .C1(n19269), .C2(n19199), .A(n19168), .B(n19167), .ZN(
        P3_U2948) );
  AOI22_X1 U22331 ( .A1(n19308), .A2(n19205), .B1(n19307), .B2(n19182), .ZN(
        n19170) );
  AOI22_X1 U22332 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19183), .B1(
        n19309), .B2(n19246), .ZN(n19169) );
  OAI211_X1 U22333 ( .C1(n19312), .C2(n19186), .A(n19170), .B(n19169), .ZN(
        P3_U2949) );
  AOI22_X1 U22334 ( .A1(n19242), .A2(n19205), .B1(n19313), .B2(n19182), .ZN(
        n19172) );
  AOI22_X1 U22335 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19183), .B1(
        n19315), .B2(n19246), .ZN(n19171) );
  OAI211_X1 U22336 ( .C1(n19245), .C2(n19186), .A(n19172), .B(n19171), .ZN(
        P3_U2950) );
  AOI22_X1 U22337 ( .A1(n19320), .A2(n19179), .B1(n19319), .B2(n19182), .ZN(
        n19174) );
  AOI22_X1 U22338 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19183), .B1(
        n19321), .B2(n19246), .ZN(n19173) );
  OAI211_X1 U22339 ( .C1(n19324), .C2(n19199), .A(n19174), .B(n19173), .ZN(
        P3_U2951) );
  AOI22_X1 U22340 ( .A1(n19326), .A2(n19179), .B1(n19325), .B2(n19182), .ZN(
        n19176) );
  AOI22_X1 U22341 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19183), .B1(
        n19327), .B2(n19246), .ZN(n19175) );
  OAI211_X1 U22342 ( .C1(n19330), .C2(n19199), .A(n19176), .B(n19175), .ZN(
        P3_U2952) );
  AOI22_X1 U22343 ( .A1(n19332), .A2(n19205), .B1(n19331), .B2(n19182), .ZN(
        n19178) );
  AOI22_X1 U22344 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19183), .B1(
        n19333), .B2(n19246), .ZN(n19177) );
  OAI211_X1 U22345 ( .C1(n19336), .C2(n19186), .A(n19178), .B(n19177), .ZN(
        P3_U2953) );
  AOI22_X1 U22346 ( .A1(n19287), .A2(n19179), .B1(n19337), .B2(n19182), .ZN(
        n19181) );
  AOI22_X1 U22347 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19183), .B1(
        n19340), .B2(n19246), .ZN(n19180) );
  OAI211_X1 U22348 ( .C1(n19290), .C2(n19199), .A(n19181), .B(n19180), .ZN(
        P3_U2954) );
  AOI22_X1 U22349 ( .A1(n19346), .A2(n19182), .B1(n19255), .B2(n19205), .ZN(
        n19185) );
  AOI22_X1 U22350 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19183), .B1(
        n19349), .B2(n19246), .ZN(n19184) );
  OAI211_X1 U22351 ( .C1(n19261), .C2(n19186), .A(n19185), .B(n19184), .ZN(
        P3_U2955) );
  NOR2_X1 U22352 ( .A1(n19387), .A2(n19187), .ZN(n19237) );
  AND2_X1 U22353 ( .A1(n19422), .A2(n19237), .ZN(n19204) );
  AOI22_X1 U22354 ( .A1(n19262), .A2(n19205), .B1(n19297), .B2(n19204), .ZN(
        n19190) );
  AOI22_X1 U22355 ( .A1(n19302), .A2(n19188), .B1(n19299), .B2(n19237), .ZN(
        n19206) );
  NAND2_X1 U22356 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19237), .ZN(
        n19281) );
  INV_X1 U22357 ( .A(n19281), .ZN(n19292) );
  AOI22_X1 U22358 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19206), .B1(
        n19303), .B2(n19292), .ZN(n19189) );
  OAI211_X1 U22359 ( .C1(n19269), .C2(n19231), .A(n19190), .B(n19189), .ZN(
        P3_U2956) );
  AOI22_X1 U22360 ( .A1(n19270), .A2(n19205), .B1(n19307), .B2(n19204), .ZN(
        n19192) );
  AOI22_X1 U22361 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19206), .B1(
        n19309), .B2(n19292), .ZN(n19191) );
  OAI211_X1 U22362 ( .C1(n19273), .C2(n19231), .A(n19192), .B(n19191), .ZN(
        P3_U2957) );
  AOI22_X1 U22363 ( .A1(n19314), .A2(n19205), .B1(n19313), .B2(n19204), .ZN(
        n19194) );
  AOI22_X1 U22364 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19206), .B1(
        n19315), .B2(n19292), .ZN(n19193) );
  OAI211_X1 U22365 ( .C1(n19318), .C2(n19231), .A(n19194), .B(n19193), .ZN(
        P3_U2958) );
  AOI22_X1 U22366 ( .A1(n19221), .A2(n19233), .B1(n19319), .B2(n19204), .ZN(
        n19196) );
  AOI22_X1 U22367 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19206), .B1(
        n19321), .B2(n19292), .ZN(n19195) );
  OAI211_X1 U22368 ( .C1(n19224), .C2(n19199), .A(n19196), .B(n19195), .ZN(
        P3_U2959) );
  AOI22_X1 U22369 ( .A1(n19278), .A2(n19233), .B1(n19325), .B2(n19204), .ZN(
        n19198) );
  AOI22_X1 U22370 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19206), .B1(
        n19327), .B2(n19292), .ZN(n19197) );
  OAI211_X1 U22371 ( .C1(n19282), .C2(n19199), .A(n19198), .B(n19197), .ZN(
        P3_U2960) );
  AOI22_X1 U22372 ( .A1(n19283), .A2(n19205), .B1(n19331), .B2(n19204), .ZN(
        n19201) );
  AOI22_X1 U22373 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19206), .B1(
        n19333), .B2(n19292), .ZN(n19200) );
  OAI211_X1 U22374 ( .C1(n19286), .C2(n19231), .A(n19201), .B(n19200), .ZN(
        P3_U2961) );
  AOI22_X1 U22375 ( .A1(n19287), .A2(n19205), .B1(n19337), .B2(n19204), .ZN(
        n19203) );
  AOI22_X1 U22376 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19206), .B1(
        n19340), .B2(n19292), .ZN(n19202) );
  OAI211_X1 U22377 ( .C1(n19290), .C2(n19231), .A(n19203), .B(n19202), .ZN(
        P3_U2962) );
  AOI22_X1 U22378 ( .A1(n19348), .A2(n19205), .B1(n19346), .B2(n19204), .ZN(
        n19208) );
  AOI22_X1 U22379 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19206), .B1(
        n19349), .B2(n19292), .ZN(n19207) );
  OAI211_X1 U22380 ( .C1(n19354), .C2(n19231), .A(n19208), .B(n19207), .ZN(
        P3_U2963) );
  NAND2_X1 U22381 ( .A1(n19385), .A2(n19301), .ZN(n19343) );
  INV_X1 U22382 ( .A(n19343), .ZN(n19347) );
  NAND2_X1 U22383 ( .A1(n19281), .A2(n19343), .ZN(n19264) );
  INV_X1 U22384 ( .A(n19264), .ZN(n19213) );
  OAI21_X1 U22385 ( .B1(n19210), .B2(n19209), .A(n19213), .ZN(n19211) );
  OAI211_X1 U22386 ( .C1(n19347), .C2(n19524), .A(n19212), .B(n19211), .ZN(
        n19234) );
  NOR2_X1 U22387 ( .A1(n19214), .A2(n19213), .ZN(n19232) );
  AOI22_X1 U22388 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19234), .B1(
        n19297), .B2(n19232), .ZN(n19216) );
  AOI22_X1 U22389 ( .A1(n19298), .A2(n19246), .B1(n19303), .B2(n19347), .ZN(
        n19215) );
  OAI211_X1 U22390 ( .C1(n19306), .C2(n19231), .A(n19216), .B(n19215), .ZN(
        P3_U2964) );
  AOI22_X1 U22391 ( .A1(n19308), .A2(n19246), .B1(n19307), .B2(n19232), .ZN(
        n19218) );
  AOI22_X1 U22392 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19234), .B1(
        n19309), .B2(n19347), .ZN(n19217) );
  OAI211_X1 U22393 ( .C1(n19312), .C2(n19231), .A(n19218), .B(n19217), .ZN(
        P3_U2965) );
  AOI22_X1 U22394 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19234), .B1(
        n19313), .B2(n19232), .ZN(n19220) );
  AOI22_X1 U22395 ( .A1(n19315), .A2(n19347), .B1(n19242), .B2(n19246), .ZN(
        n19219) );
  OAI211_X1 U22396 ( .C1(n19245), .C2(n19231), .A(n19220), .B(n19219), .ZN(
        P3_U2966) );
  AOI22_X1 U22397 ( .A1(n19221), .A2(n19246), .B1(n19319), .B2(n19232), .ZN(
        n19223) );
  AOI22_X1 U22398 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19234), .B1(
        n19321), .B2(n19347), .ZN(n19222) );
  OAI211_X1 U22399 ( .C1(n19224), .C2(n19231), .A(n19223), .B(n19222), .ZN(
        P3_U2967) );
  AOI22_X1 U22400 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19234), .B1(
        n19325), .B2(n19232), .ZN(n19226) );
  AOI22_X1 U22401 ( .A1(n19326), .A2(n19233), .B1(n19327), .B2(n19347), .ZN(
        n19225) );
  OAI211_X1 U22402 ( .C1(n19330), .C2(n19260), .A(n19226), .B(n19225), .ZN(
        P3_U2968) );
  AOI22_X1 U22403 ( .A1(n19332), .A2(n19246), .B1(n19331), .B2(n19232), .ZN(
        n19228) );
  AOI22_X1 U22404 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19234), .B1(
        n19333), .B2(n19347), .ZN(n19227) );
  OAI211_X1 U22405 ( .C1(n19336), .C2(n19231), .A(n19228), .B(n19227), .ZN(
        P3_U2969) );
  AOI22_X1 U22406 ( .A1(n19338), .A2(n19246), .B1(n19337), .B2(n19232), .ZN(
        n19230) );
  AOI22_X1 U22407 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19234), .B1(
        n19340), .B2(n19347), .ZN(n19229) );
  OAI211_X1 U22408 ( .C1(n19344), .C2(n19231), .A(n19230), .B(n19229), .ZN(
        P3_U2970) );
  AOI22_X1 U22409 ( .A1(n19348), .A2(n19233), .B1(n19346), .B2(n19232), .ZN(
        n19236) );
  AOI22_X1 U22410 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19234), .B1(
        n19349), .B2(n19347), .ZN(n19235) );
  OAI211_X1 U22411 ( .C1(n19354), .C2(n19260), .A(n19236), .B(n19235), .ZN(
        P3_U2971) );
  AND2_X1 U22412 ( .A1(n19422), .A2(n19301), .ZN(n19256) );
  AOI22_X1 U22413 ( .A1(n19262), .A2(n19246), .B1(n19297), .B2(n19256), .ZN(
        n19239) );
  AOI22_X1 U22414 ( .A1(n19302), .A2(n19237), .B1(n19301), .B2(n19299), .ZN(
        n19257) );
  AOI22_X1 U22415 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19257), .B1(
        n19303), .B2(n19339), .ZN(n19238) );
  OAI211_X1 U22416 ( .C1(n19269), .C2(n19281), .A(n19239), .B(n19238), .ZN(
        P3_U2972) );
  AOI22_X1 U22417 ( .A1(n19308), .A2(n19292), .B1(n19307), .B2(n19256), .ZN(
        n19241) );
  AOI22_X1 U22418 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19257), .B1(
        n19339), .B2(n19309), .ZN(n19240) );
  OAI211_X1 U22419 ( .C1(n19312), .C2(n19260), .A(n19241), .B(n19240), .ZN(
        P3_U2973) );
  AOI22_X1 U22420 ( .A1(n19242), .A2(n19292), .B1(n19313), .B2(n19256), .ZN(
        n19244) );
  AOI22_X1 U22421 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19257), .B1(
        n19339), .B2(n19315), .ZN(n19243) );
  OAI211_X1 U22422 ( .C1(n19245), .C2(n19260), .A(n19244), .B(n19243), .ZN(
        P3_U2974) );
  AOI22_X1 U22423 ( .A1(n19320), .A2(n19246), .B1(n19319), .B2(n19256), .ZN(
        n19248) );
  AOI22_X1 U22424 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19257), .B1(
        n19339), .B2(n19321), .ZN(n19247) );
  OAI211_X1 U22425 ( .C1(n19324), .C2(n19281), .A(n19248), .B(n19247), .ZN(
        P3_U2975) );
  AOI22_X1 U22426 ( .A1(n19278), .A2(n19292), .B1(n19325), .B2(n19256), .ZN(
        n19250) );
  AOI22_X1 U22427 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19257), .B1(
        n19339), .B2(n19327), .ZN(n19249) );
  OAI211_X1 U22428 ( .C1(n19282), .C2(n19260), .A(n19250), .B(n19249), .ZN(
        P3_U2976) );
  AOI22_X1 U22429 ( .A1(n19332), .A2(n19292), .B1(n19331), .B2(n19256), .ZN(
        n19252) );
  AOI22_X1 U22430 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19257), .B1(
        n19339), .B2(n19333), .ZN(n19251) );
  OAI211_X1 U22431 ( .C1(n19336), .C2(n19260), .A(n19252), .B(n19251), .ZN(
        P3_U2977) );
  AOI22_X1 U22432 ( .A1(n19338), .A2(n19292), .B1(n19337), .B2(n19256), .ZN(
        n19254) );
  AOI22_X1 U22433 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19257), .B1(
        n19339), .B2(n19340), .ZN(n19253) );
  OAI211_X1 U22434 ( .C1(n19344), .C2(n19260), .A(n19254), .B(n19253), .ZN(
        P3_U2978) );
  AOI22_X1 U22435 ( .A1(n19346), .A2(n19256), .B1(n19255), .B2(n19292), .ZN(
        n19259) );
  AOI22_X1 U22436 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19257), .B1(
        n19339), .B2(n19349), .ZN(n19258) );
  OAI211_X1 U22437 ( .C1(n19261), .C2(n19260), .A(n19259), .B(n19258), .ZN(
        P3_U2979) );
  AND2_X1 U22438 ( .A1(n19422), .A2(n19266), .ZN(n19291) );
  AOI22_X1 U22439 ( .A1(n19262), .A2(n19292), .B1(n19297), .B2(n19291), .ZN(
        n19268) );
  OAI221_X1 U22440 ( .B1(n19266), .B2(n19265), .C1(n19266), .C2(n19264), .A(
        n19263), .ZN(n19294) );
  AOI22_X1 U22441 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19294), .B1(
        n19293), .B2(n19303), .ZN(n19267) );
  OAI211_X1 U22442 ( .C1(n19269), .C2(n19343), .A(n19268), .B(n19267), .ZN(
        P3_U2980) );
  AOI22_X1 U22443 ( .A1(n19270), .A2(n19292), .B1(n19307), .B2(n19291), .ZN(
        n19272) );
  AOI22_X1 U22444 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19294), .B1(
        n19293), .B2(n19309), .ZN(n19271) );
  OAI211_X1 U22445 ( .C1(n19273), .C2(n19343), .A(n19272), .B(n19271), .ZN(
        P3_U2981) );
  AOI22_X1 U22446 ( .A1(n19314), .A2(n19292), .B1(n19313), .B2(n19291), .ZN(
        n19275) );
  AOI22_X1 U22447 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19294), .B1(
        n19293), .B2(n19315), .ZN(n19274) );
  OAI211_X1 U22448 ( .C1(n19318), .C2(n19343), .A(n19275), .B(n19274), .ZN(
        P3_U2982) );
  AOI22_X1 U22449 ( .A1(n19320), .A2(n19292), .B1(n19319), .B2(n19291), .ZN(
        n19277) );
  AOI22_X1 U22450 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19294), .B1(
        n19293), .B2(n19321), .ZN(n19276) );
  OAI211_X1 U22451 ( .C1(n19324), .C2(n19343), .A(n19277), .B(n19276), .ZN(
        P3_U2983) );
  AOI22_X1 U22452 ( .A1(n19278), .A2(n19347), .B1(n19325), .B2(n19291), .ZN(
        n19280) );
  AOI22_X1 U22453 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19294), .B1(
        n19293), .B2(n19327), .ZN(n19279) );
  OAI211_X1 U22454 ( .C1(n19282), .C2(n19281), .A(n19280), .B(n19279), .ZN(
        P3_U2984) );
  AOI22_X1 U22455 ( .A1(n19283), .A2(n19292), .B1(n19331), .B2(n19291), .ZN(
        n19285) );
  AOI22_X1 U22456 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19294), .B1(
        n19293), .B2(n19333), .ZN(n19284) );
  OAI211_X1 U22457 ( .C1(n19286), .C2(n19343), .A(n19285), .B(n19284), .ZN(
        P3_U2985) );
  AOI22_X1 U22458 ( .A1(n19287), .A2(n19292), .B1(n19337), .B2(n19291), .ZN(
        n19289) );
  AOI22_X1 U22459 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19294), .B1(
        n19293), .B2(n19340), .ZN(n19288) );
  OAI211_X1 U22460 ( .C1(n19290), .C2(n19343), .A(n19289), .B(n19288), .ZN(
        P3_U2986) );
  AOI22_X1 U22461 ( .A1(n19348), .A2(n19292), .B1(n19346), .B2(n19291), .ZN(
        n19296) );
  AOI22_X1 U22462 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19294), .B1(
        n19293), .B2(n19349), .ZN(n19295) );
  OAI211_X1 U22463 ( .C1(n19354), .C2(n19343), .A(n19296), .B(n19295), .ZN(
        P3_U2987) );
  AND2_X1 U22464 ( .A1(n19422), .A2(n19300), .ZN(n19345) );
  AOI22_X1 U22465 ( .A1(n19298), .A2(n19339), .B1(n19297), .B2(n19345), .ZN(
        n19305) );
  AOI22_X1 U22466 ( .A1(n19302), .A2(n19301), .B1(n19300), .B2(n19299), .ZN(
        n19351) );
  AOI22_X1 U22467 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19303), .ZN(n19304) );
  OAI211_X1 U22468 ( .C1(n19306), .C2(n19343), .A(n19305), .B(n19304), .ZN(
        P3_U2988) );
  AOI22_X1 U22469 ( .A1(n19339), .A2(n19308), .B1(n19307), .B2(n19345), .ZN(
        n19311) );
  AOI22_X1 U22470 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19309), .ZN(n19310) );
  OAI211_X1 U22471 ( .C1(n19312), .C2(n19343), .A(n19311), .B(n19310), .ZN(
        P3_U2989) );
  AOI22_X1 U22472 ( .A1(n19314), .A2(n19347), .B1(n19313), .B2(n19345), .ZN(
        n19317) );
  AOI22_X1 U22473 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19315), .ZN(n19316) );
  OAI211_X1 U22474 ( .C1(n19355), .C2(n19318), .A(n19317), .B(n19316), .ZN(
        P3_U2990) );
  AOI22_X1 U22475 ( .A1(n19320), .A2(n19347), .B1(n19319), .B2(n19345), .ZN(
        n19323) );
  AOI22_X1 U22476 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19321), .ZN(n19322) );
  OAI211_X1 U22477 ( .C1(n19355), .C2(n19324), .A(n19323), .B(n19322), .ZN(
        P3_U2991) );
  AOI22_X1 U22478 ( .A1(n19326), .A2(n19347), .B1(n19325), .B2(n19345), .ZN(
        n19329) );
  AOI22_X1 U22479 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19327), .ZN(n19328) );
  OAI211_X1 U22480 ( .C1(n19355), .C2(n19330), .A(n19329), .B(n19328), .ZN(
        P3_U2992) );
  AOI22_X1 U22481 ( .A1(n19339), .A2(n19332), .B1(n19331), .B2(n19345), .ZN(
        n19335) );
  AOI22_X1 U22482 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19333), .ZN(n19334) );
  OAI211_X1 U22483 ( .C1(n19336), .C2(n19343), .A(n19335), .B(n19334), .ZN(
        P3_U2993) );
  AOI22_X1 U22484 ( .A1(n19339), .A2(n19338), .B1(n19337), .B2(n19345), .ZN(
        n19342) );
  AOI22_X1 U22485 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19340), .ZN(n19341) );
  OAI211_X1 U22486 ( .C1(n19344), .C2(n19343), .A(n19342), .B(n19341), .ZN(
        P3_U2994) );
  AOI22_X1 U22487 ( .A1(n19348), .A2(n19347), .B1(n19346), .B2(n19345), .ZN(
        n19353) );
  AOI22_X1 U22488 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19349), .ZN(n19352) );
  OAI211_X1 U22489 ( .C1(n19355), .C2(n19354), .A(n19353), .B(n19352), .ZN(
        P3_U2995) );
  AOI21_X1 U22490 ( .B1(n19358), .B2(n19357), .A(n19356), .ZN(n19362) );
  AOI21_X1 U22491 ( .B1(n19397), .B2(n19360), .A(n19359), .ZN(n19361) );
  AOI211_X1 U22492 ( .C1(n19364), .C2(n19363), .A(n19362), .B(n19361), .ZN(
        n19566) );
  AOI211_X1 U22493 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n19398), .A(
        n19366), .B(n19365), .ZN(n19412) );
  OAI21_X1 U22494 ( .B1(n19369), .B2(n19368), .A(n19367), .ZN(n19393) );
  AOI22_X1 U22495 ( .A1(n19391), .A2(n19371), .B1(n19370), .B2(n19393), .ZN(
        n19374) );
  NOR2_X1 U22496 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19372), .ZN(
        n19376) );
  INV_X1 U22497 ( .A(n19376), .ZN(n19373) );
  NAND2_X1 U22498 ( .A1(n19374), .A2(n19373), .ZN(n19530) );
  NOR2_X1 U22499 ( .A1(n19531), .A2(n19530), .ZN(n19378) );
  OAI21_X1 U22500 ( .B1(n19554), .B2(n19375), .A(n19382), .ZN(n19392) );
  INV_X1 U22501 ( .A(n19392), .ZN(n19383) );
  OAI22_X1 U22502 ( .A1(n19383), .A2(n19391), .B1(n19376), .B2(n19397), .ZN(
        n19527) );
  AOI21_X1 U22503 ( .B1(n19527), .B2(n19379), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19377) );
  AOI21_X1 U22504 ( .B1(n19379), .B2(n19378), .A(n19377), .ZN(n19408) );
  NOR2_X1 U22505 ( .A1(n19381), .A2(n19380), .ZN(n19384) );
  AOI22_X1 U22506 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19382), .B1(
        n19384), .B2(n19554), .ZN(n19550) );
  OAI22_X1 U22507 ( .A1(n19384), .A2(n19542), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19383), .ZN(n19546) );
  OR3_X1 U22508 ( .A1(n19550), .A2(n19387), .A3(n19385), .ZN(n19386) );
  AOI22_X1 U22509 ( .A1(n19550), .A2(n19387), .B1(n19546), .B2(n19386), .ZN(
        n19389) );
  OAI21_X1 U22510 ( .B1(n19398), .B2(n19389), .A(n19388), .ZN(n19402) );
  NAND2_X1 U22511 ( .A1(n19403), .A2(n19402), .ZN(n19400) );
  INV_X1 U22512 ( .A(n19390), .ZN(n19537) );
  OAI211_X1 U22513 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n19392), .B(n19391), .ZN(
        n19396) );
  NAND3_X1 U22514 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19394), .A3(
        n19393), .ZN(n19395) );
  OAI211_X1 U22515 ( .C1(n19537), .C2(n19397), .A(n19396), .B(n19395), .ZN(
        n19539) );
  MUX2_X1 U22516 ( .A(n19539), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n19398), .Z(n19401) );
  INV_X1 U22517 ( .A(n19401), .ZN(n19399) );
  OAI221_X1 U22518 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n19400), .A(n19399), .ZN(
        n19407) );
  NOR2_X1 U22519 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19406) );
  OAI222_X1 U22520 ( .A1(n19403), .A2(n19402), .B1(n19403), .B2(n19401), .C1(
        n19402), .C2(n19401), .ZN(n19404) );
  INV_X1 U22521 ( .A(n19404), .ZN(n19405) );
  AOI22_X1 U22522 ( .A1(n19408), .A2(n19407), .B1(n19406), .B2(n19405), .ZN(
        n19411) );
  OAI21_X1 U22523 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19409), .ZN(n19410) );
  NAND4_X1 U22524 ( .A1(n19566), .A2(n19412), .A3(n19411), .A4(n19410), .ZN(
        n19419) );
  AOI211_X1 U22525 ( .C1(n19415), .C2(n19414), .A(n19413), .B(n19419), .ZN(
        n19522) );
  AOI21_X1 U22526 ( .B1(n19575), .B2(n19587), .A(n19522), .ZN(n19423) );
  NAND2_X1 U22527 ( .A1(n19575), .A2(n19569), .ZN(n19427) );
  INV_X1 U22528 ( .A(n19427), .ZN(n19416) );
  AOI211_X1 U22529 ( .C1(n19549), .C2(n19580), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n19416), .ZN(n19417) );
  AOI211_X1 U22530 ( .C1(n19572), .C2(n19419), .A(n19418), .B(n19417), .ZN(
        n19420) );
  OAI221_X1 U22531 ( .B1(n19577), .B2(n19423), .C1(n19577), .C2(n19421), .A(
        n19420), .ZN(P3_U2996) );
  NOR4_X1 U22532 ( .A1(n19577), .A2(n19534), .A3(n19568), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19430) );
  INV_X1 U22533 ( .A(n19430), .ZN(n19426) );
  NAND3_X1 U22534 ( .A1(n19424), .A2(n19423), .A3(n19422), .ZN(n19425) );
  NAND4_X1 U22535 ( .A1(n19428), .A2(n19427), .A3(n19426), .A4(n19425), .ZN(
        P3_U2997) );
  OAI21_X1 U22536 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(
        P3_STATE2_REG_0__SCAN_IN), .A(n19429), .ZN(n19431) );
  AOI21_X1 U22537 ( .B1(n19432), .B2(n19431), .A(n19430), .ZN(P3_U2998) );
  AND2_X1 U22538 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19433), .ZN(
        P3_U2999) );
  AND2_X1 U22539 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19433), .ZN(
        P3_U3000) );
  AND2_X1 U22540 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19433), .ZN(
        P3_U3001) );
  AND2_X1 U22541 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19433), .ZN(
        P3_U3002) );
  AND2_X1 U22542 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19433), .ZN(
        P3_U3003) );
  AND2_X1 U22543 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19433), .ZN(
        P3_U3004) );
  AND2_X1 U22544 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19433), .ZN(
        P3_U3005) );
  AND2_X1 U22545 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19433), .ZN(
        P3_U3006) );
  AND2_X1 U22546 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19433), .ZN(
        P3_U3007) );
  AND2_X1 U22547 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19433), .ZN(
        P3_U3008) );
  AND2_X1 U22548 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19433), .ZN(
        P3_U3009) );
  AND2_X1 U22549 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19433), .ZN(
        P3_U3010) );
  AND2_X1 U22550 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19433), .ZN(
        P3_U3011) );
  AND2_X1 U22551 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19433), .ZN(
        P3_U3012) );
  AND2_X1 U22552 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19433), .ZN(
        P3_U3013) );
  AND2_X1 U22553 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19433), .ZN(
        P3_U3014) );
  AND2_X1 U22554 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19433), .ZN(
        P3_U3015) );
  AND2_X1 U22555 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19433), .ZN(
        P3_U3016) );
  AND2_X1 U22556 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19433), .ZN(
        P3_U3017) );
  AND2_X1 U22557 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19433), .ZN(
        P3_U3018) );
  AND2_X1 U22558 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19433), .ZN(
        P3_U3019) );
  AND2_X1 U22559 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19433), .ZN(
        P3_U3020) );
  AND2_X1 U22560 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19433), .ZN(P3_U3021) );
  AND2_X1 U22561 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19433), .ZN(P3_U3022) );
  AND2_X1 U22562 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19433), .ZN(P3_U3023) );
  AND2_X1 U22563 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19433), .ZN(P3_U3024) );
  AND2_X1 U22564 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19433), .ZN(P3_U3025) );
  AND2_X1 U22565 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19433), .ZN(P3_U3026) );
  AND2_X1 U22566 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19433), .ZN(P3_U3027) );
  AND2_X1 U22567 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19433), .ZN(P3_U3028) );
  INV_X1 U22568 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19437) );
  NOR2_X1 U22569 ( .A1(n19450), .A2(n20971), .ZN(n19446) );
  INV_X1 U22570 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19582) );
  NOR2_X1 U22571 ( .A1(n19446), .A2(n19582), .ZN(n19439) );
  OAI21_X1 U22572 ( .B1(n19437), .B2(n20971), .A(n19439), .ZN(n19434) );
  AOI22_X1 U22573 ( .A1(n19448), .A2(n19450), .B1(n19585), .B2(n19434), .ZN(
        n19435) );
  NAND3_X1 U22574 ( .A1(NA), .A2(n19448), .A3(n19437), .ZN(n19443) );
  OAI211_X1 U22575 ( .C1(n19568), .C2(n19436), .A(n19435), .B(n19443), .ZN(
        P3_U3029) );
  NOR2_X1 U22576 ( .A1(n19437), .A2(n20971), .ZN(n19438) );
  AOI22_X1 U22577 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19439), .B1(n19438), 
        .B2(n19450), .ZN(n19441) );
  NAND2_X1 U22578 ( .A1(n19575), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19444) );
  NAND3_X1 U22579 ( .A1(n19441), .A2(n19440), .A3(n19444), .ZN(P3_U3030) );
  INV_X1 U22580 ( .A(n19444), .ZN(n19442) );
  AOI21_X1 U22581 ( .B1(n19448), .B2(n19443), .A(n19442), .ZN(n19449) );
  OAI22_X1 U22582 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19444), .ZN(n19445) );
  OAI22_X1 U22583 ( .A1(n19446), .A2(n19445), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19447) );
  OAI22_X1 U22584 ( .A1(n19449), .A2(n19450), .B1(n19448), .B2(n19447), .ZN(
        P3_U3031) );
  INV_X1 U22585 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19453) );
  OAI222_X1 U22586 ( .A1(n19452), .A2(n19509), .B1(n19451), .B2(n19584), .C1(
        n19453), .C2(n19513), .ZN(P3_U3032) );
  OAI222_X1 U22587 ( .A1(n19513), .A2(n19455), .B1(n19454), .B2(n19584), .C1(
        n19453), .C2(n19509), .ZN(P3_U3033) );
  OAI222_X1 U22588 ( .A1(n19513), .A2(n19457), .B1(n19456), .B2(n19584), .C1(
        n19455), .C2(n19509), .ZN(P3_U3034) );
  INV_X1 U22589 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19459) );
  OAI222_X1 U22590 ( .A1(n19513), .A2(n19459), .B1(n19458), .B2(n19584), .C1(
        n19457), .C2(n19509), .ZN(P3_U3035) );
  OAI222_X1 U22591 ( .A1(n19513), .A2(n19461), .B1(n19460), .B2(n19584), .C1(
        n19459), .C2(n19509), .ZN(P3_U3036) );
  OAI222_X1 U22592 ( .A1(n19513), .A2(n19463), .B1(n19462), .B2(n19584), .C1(
        n19461), .C2(n19509), .ZN(P3_U3037) );
  OAI222_X1 U22593 ( .A1(n19513), .A2(n19465), .B1(n19464), .B2(n19584), .C1(
        n19463), .C2(n19509), .ZN(P3_U3038) );
  OAI222_X1 U22594 ( .A1(n19513), .A2(n19467), .B1(n19466), .B2(n19584), .C1(
        n19465), .C2(n19509), .ZN(P3_U3039) );
  OAI222_X1 U22595 ( .A1(n19513), .A2(n19469), .B1(n19468), .B2(n19584), .C1(
        n19467), .C2(n19509), .ZN(P3_U3040) );
  INV_X1 U22596 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19471) );
  OAI222_X1 U22597 ( .A1(n19513), .A2(n19471), .B1(n19470), .B2(n19584), .C1(
        n19469), .C2(n19509), .ZN(P3_U3041) );
  OAI222_X1 U22598 ( .A1(n19513), .A2(n19474), .B1(n19472), .B2(n19584), .C1(
        n19471), .C2(n19509), .ZN(P3_U3042) );
  INV_X1 U22599 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19475) );
  OAI222_X1 U22600 ( .A1(n19474), .A2(n19509), .B1(n19473), .B2(n19584), .C1(
        n19475), .C2(n19513), .ZN(P3_U3043) );
  OAI222_X1 U22601 ( .A1(n19513), .A2(n19478), .B1(n19476), .B2(n19584), .C1(
        n19475), .C2(n19509), .ZN(P3_U3044) );
  OAI222_X1 U22602 ( .A1(n19478), .A2(n19509), .B1(n19477), .B2(n19584), .C1(
        n19479), .C2(n19513), .ZN(P3_U3045) );
  OAI222_X1 U22603 ( .A1(n19513), .A2(n19481), .B1(n19480), .B2(n19584), .C1(
        n19479), .C2(n19509), .ZN(P3_U3046) );
  OAI222_X1 U22604 ( .A1(n19513), .A2(n19484), .B1(n19482), .B2(n19584), .C1(
        n19481), .C2(n19509), .ZN(P3_U3047) );
  OAI222_X1 U22605 ( .A1(n19484), .A2(n19509), .B1(n19483), .B2(n19584), .C1(
        n19485), .C2(n19513), .ZN(P3_U3048) );
  OAI222_X1 U22606 ( .A1(n19513), .A2(n19487), .B1(n19486), .B2(n19584), .C1(
        n19485), .C2(n19509), .ZN(P3_U3049) );
  OAI222_X1 U22607 ( .A1(n19513), .A2(n19490), .B1(n19488), .B2(n19584), .C1(
        n19487), .C2(n19509), .ZN(P3_U3050) );
  OAI222_X1 U22608 ( .A1(n19509), .A2(n19490), .B1(n19489), .B2(n19584), .C1(
        n19491), .C2(n19513), .ZN(P3_U3051) );
  OAI222_X1 U22609 ( .A1(n19513), .A2(n19493), .B1(n19492), .B2(n19584), .C1(
        n19491), .C2(n19509), .ZN(P3_U3052) );
  OAI222_X1 U22610 ( .A1(n19513), .A2(n19496), .B1(n19494), .B2(n19584), .C1(
        n19493), .C2(n19509), .ZN(P3_U3053) );
  OAI222_X1 U22611 ( .A1(n19496), .A2(n19509), .B1(n19495), .B2(n19584), .C1(
        n19498), .C2(n19513), .ZN(P3_U3054) );
  OAI222_X1 U22612 ( .A1(n19498), .A2(n19509), .B1(n19497), .B2(n19584), .C1(
        n19499), .C2(n19513), .ZN(P3_U3055) );
  OAI222_X1 U22613 ( .A1(n19513), .A2(n19501), .B1(n19500), .B2(n19584), .C1(
        n19499), .C2(n19509), .ZN(P3_U3056) );
  OAI222_X1 U22614 ( .A1(n19513), .A2(n19503), .B1(n19502), .B2(n19584), .C1(
        n19501), .C2(n19509), .ZN(P3_U3057) );
  OAI222_X1 U22615 ( .A1(n19513), .A2(n19506), .B1(n19504), .B2(n19584), .C1(
        n19503), .C2(n19509), .ZN(P3_U3058) );
  OAI222_X1 U22616 ( .A1(n19506), .A2(n19509), .B1(n19505), .B2(n19584), .C1(
        n19508), .C2(n19513), .ZN(P3_U3059) );
  OAI222_X1 U22617 ( .A1(n19509), .A2(n19508), .B1(n19507), .B2(n19584), .C1(
        n19510), .C2(n19513), .ZN(P3_U3060) );
  OAI222_X1 U22618 ( .A1(n19513), .A2(n19512), .B1(n19511), .B2(n19584), .C1(
        n19510), .C2(n19509), .ZN(P3_U3061) );
  OAI22_X1 U22619 ( .A1(n19585), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19584), .ZN(n19514) );
  INV_X1 U22620 ( .A(n19514), .ZN(P3_U3274) );
  OAI22_X1 U22621 ( .A1(n19585), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19584), .ZN(n19515) );
  INV_X1 U22622 ( .A(n19515), .ZN(P3_U3275) );
  OAI22_X1 U22623 ( .A1(n19585), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19584), .ZN(n19516) );
  INV_X1 U22624 ( .A(n19516), .ZN(P3_U3276) );
  OAI22_X1 U22625 ( .A1(n19585), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19584), .ZN(n19517) );
  INV_X1 U22626 ( .A(n19517), .ZN(P3_U3277) );
  OAI21_X1 U22627 ( .B1(n19521), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19519), 
        .ZN(n19518) );
  INV_X1 U22628 ( .A(n19518), .ZN(P3_U3280) );
  OAI21_X1 U22629 ( .B1(n19521), .B2(n19520), .A(n19519), .ZN(P3_U3281) );
  NOR2_X1 U22630 ( .A1(n19522), .A2(n19577), .ZN(n19525) );
  OAI21_X1 U22631 ( .B1(n19525), .B2(n19524), .A(n19523), .ZN(P3_U3282) );
  NOR2_X1 U22632 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19526), .ZN(
        n19528) );
  AOI22_X1 U22633 ( .A1(n19549), .A2(n19529), .B1(n19528), .B2(n19527), .ZN(
        n19533) );
  AOI21_X1 U22634 ( .B1(n19588), .B2(n19530), .A(n19555), .ZN(n19532) );
  OAI22_X1 U22635 ( .A1(n19555), .A2(n19533), .B1(n19532), .B2(n19531), .ZN(
        P3_U3285) );
  NOR2_X1 U22636 ( .A1(n19534), .A2(n19551), .ZN(n19543) );
  OAI22_X1 U22637 ( .A1(n19536), .A2(n19535), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19544) );
  INV_X1 U22638 ( .A(n19544), .ZN(n19538) );
  AOI222_X1 U22639 ( .A1(n19539), .A2(n19588), .B1(n19543), .B2(n19538), .C1(
        n19549), .C2(n19537), .ZN(n19540) );
  AOI22_X1 U22640 ( .A1(n19555), .A2(n19541), .B1(n19540), .B2(n19552), .ZN(
        P3_U3288) );
  INV_X1 U22641 ( .A(n19542), .ZN(n19545) );
  AOI222_X1 U22642 ( .A1(n19546), .A2(n19588), .B1(n19549), .B2(n19545), .C1(
        n19544), .C2(n19543), .ZN(n19547) );
  AOI22_X1 U22643 ( .A1(n19555), .A2(n19548), .B1(n19547), .B2(n19552), .ZN(
        P3_U3289) );
  AOI222_X1 U22644 ( .A1(n19551), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19588), 
        .B2(n19550), .C1(n19554), .C2(n19549), .ZN(n19553) );
  AOI22_X1 U22645 ( .A1(n19555), .A2(n19554), .B1(n19553), .B2(n19552), .ZN(
        P3_U3290) );
  AOI211_X1 U22646 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19556) );
  AOI21_X1 U22647 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19556), .ZN(n19558) );
  INV_X1 U22648 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19557) );
  AOI22_X1 U22649 ( .A1(n19562), .A2(n19558), .B1(n19557), .B2(n19559), .ZN(
        P3_U3292) );
  NOR2_X1 U22650 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n19561) );
  INV_X1 U22651 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19560) );
  AOI22_X1 U22652 ( .A1(n19562), .A2(n19561), .B1(n19560), .B2(n19559), .ZN(
        P3_U3293) );
  INV_X1 U22653 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19591) );
  OAI22_X1 U22654 ( .A1(n19585), .A2(n19591), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n19584), .ZN(n19563) );
  INV_X1 U22655 ( .A(n19563), .ZN(P3_U3294) );
  INV_X1 U22656 ( .A(n19564), .ZN(n19567) );
  NAND2_X1 U22657 ( .A1(n19567), .A2(P3_MORE_REG_SCAN_IN), .ZN(n19565) );
  OAI21_X1 U22658 ( .B1(n19567), .B2(n19566), .A(n19565), .ZN(P3_U3295) );
  AOI21_X1 U22659 ( .B1(n19569), .B2(n19568), .A(n19590), .ZN(n19570) );
  OAI21_X1 U22660 ( .B1(n19572), .B2(n19571), .A(n19570), .ZN(n19583) );
  OAI21_X1 U22661 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n19574), .A(n19573), 
        .ZN(n19576) );
  AOI211_X1 U22662 ( .C1(n19589), .C2(n19576), .A(n19575), .B(n19587), .ZN(
        n19578) );
  NOR2_X1 U22663 ( .A1(n19578), .A2(n19577), .ZN(n19579) );
  OAI21_X1 U22664 ( .B1(n19580), .B2(n19579), .A(n19583), .ZN(n19581) );
  OAI21_X1 U22665 ( .B1(n19583), .B2(n19582), .A(n19581), .ZN(P3_U3296) );
  OAI22_X1 U22666 ( .A1(n19585), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19584), .ZN(n19586) );
  INV_X1 U22667 ( .A(n19586), .ZN(P3_U3297) );
  AOI21_X1 U22668 ( .B1(n19588), .B2(n19587), .A(n19590), .ZN(n19594) );
  AOI22_X1 U22669 ( .A1(n19594), .A2(n19591), .B1(n19590), .B2(n19589), .ZN(
        P3_U3298) );
  INV_X1 U22670 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19593) );
  AOI21_X1 U22671 ( .B1(n19594), .B2(n19593), .A(n19592), .ZN(P3_U3299) );
  NAND2_X1 U22672 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20517), .ZN(n20507) );
  NAND2_X1 U22673 ( .A1(n19600), .A2(n19595), .ZN(n20504) );
  OAI21_X1 U22674 ( .B1(n19600), .B2(n20507), .A(n20504), .ZN(n20566) );
  AOI21_X1 U22675 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20566), .ZN(n19596) );
  INV_X1 U22676 ( .A(n19596), .ZN(P2_U2815) );
  INV_X1 U22677 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19601) );
  OAI22_X1 U22678 ( .A1(n19599), .A2(n19601), .B1(n19598), .B2(n19597), .ZN(
        P2_U2816) );
  INV_X1 U22679 ( .A(n20498), .ZN(n20512) );
  NAND2_X1 U22680 ( .A1(n19600), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20628) );
  INV_X2 U22681 ( .A(n20628), .ZN(n20627) );
  AOI22_X1 U22682 ( .A1(n20627), .A2(n19601), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n20628), .ZN(n19602) );
  OAI21_X1 U22683 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20512), .A(n19602), 
        .ZN(P2_U2817) );
  OAI21_X1 U22684 ( .B1(n20498), .B2(BS16), .A(n20566), .ZN(n20564) );
  OAI21_X1 U22685 ( .B1(n20566), .B2(n21109), .A(n20564), .ZN(P2_U2818) );
  NOR4_X1 U22686 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19606) );
  NOR4_X1 U22687 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19605) );
  NOR4_X1 U22688 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19604) );
  NOR4_X1 U22689 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19603) );
  NAND4_X1 U22690 ( .A1(n19606), .A2(n19605), .A3(n19604), .A4(n19603), .ZN(
        n19612) );
  NOR4_X1 U22691 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19610) );
  AOI211_X1 U22692 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19609) );
  NOR4_X1 U22693 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19608) );
  NOR4_X1 U22694 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19607) );
  NAND4_X1 U22695 ( .A1(n19610), .A2(n19609), .A3(n19608), .A4(n19607), .ZN(
        n19611) );
  NOR2_X1 U22696 ( .A1(n19612), .A2(n19611), .ZN(n19622) );
  INV_X1 U22697 ( .A(n19622), .ZN(n19620) );
  NOR2_X1 U22698 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19620), .ZN(n19615) );
  INV_X1 U22699 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19613) );
  AOI22_X1 U22700 ( .A1(n19615), .A2(n10475), .B1(n19620), .B2(n19613), .ZN(
        P2_U2820) );
  OR3_X1 U22701 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19619) );
  INV_X1 U22702 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19614) );
  AOI22_X1 U22703 ( .A1(n19615), .A2(n19619), .B1(n19620), .B2(n19614), .ZN(
        P2_U2821) );
  INV_X1 U22704 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20565) );
  NAND2_X1 U22705 ( .A1(n19615), .A2(n20565), .ZN(n19618) );
  OAI21_X1 U22706 ( .B1(n14081), .B2(n10475), .A(n19622), .ZN(n19616) );
  OAI21_X1 U22707 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19622), .A(n19616), 
        .ZN(n19617) );
  OAI221_X1 U22708 ( .B1(n19618), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19618), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19617), .ZN(P2_U2822) );
  INV_X1 U22709 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19621) );
  OAI221_X1 U22710 ( .B1(n19622), .B2(n19621), .C1(n19620), .C2(n19619), .A(
        n19618), .ZN(P2_U2823) );
  INV_X1 U22711 ( .A(n19623), .ZN(n19634) );
  AOI21_X1 U22712 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19732), .A(
        n19903), .ZN(n19624) );
  OAI21_X1 U22713 ( .B1(n19737), .B2(n20537), .A(n19624), .ZN(n19625) );
  AOI21_X1 U22714 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19744), .A(n19625), .ZN(
        n19626) );
  OAI21_X1 U22715 ( .B1(n19627), .B2(n19748), .A(n19626), .ZN(n19633) );
  OAI21_X1 U22716 ( .B1(n19629), .B2(n19628), .A(n19757), .ZN(n19631) );
  INV_X1 U22717 ( .A(n15431), .ZN(n19630) );
  AOI21_X1 U22718 ( .B1(n19665), .B2(n19631), .A(n19630), .ZN(n19632) );
  AOI211_X1 U22719 ( .C1(n19734), .C2(n19634), .A(n19633), .B(n19632), .ZN(
        n19635) );
  OAI21_X1 U22720 ( .B1(n19636), .B2(n19726), .A(n19635), .ZN(P2_U2836) );
  INV_X1 U22721 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19638) );
  NAND2_X1 U22722 ( .A1(n19652), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n19637) );
  OAI211_X1 U22723 ( .C1(n19654), .C2(n19638), .A(n19637), .B(n19736), .ZN(
        n19639) );
  AOI21_X1 U22724 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n19744), .A(n19639), .ZN(
        n19640) );
  OAI21_X1 U22725 ( .B1(n19641), .B2(n19748), .A(n19640), .ZN(n19648) );
  OAI21_X1 U22726 ( .B1(n19643), .B2(n19642), .A(n19757), .ZN(n19646) );
  INV_X1 U22727 ( .A(n19644), .ZN(n19645) );
  AOI21_X1 U22728 ( .B1(n19665), .B2(n19646), .A(n19645), .ZN(n19647) );
  AOI211_X1 U22729 ( .C1(n19734), .C2(n19649), .A(n19648), .B(n19647), .ZN(
        n19650) );
  OAI21_X1 U22730 ( .B1(n19651), .B2(n19726), .A(n19650), .ZN(P2_U2838) );
  INV_X1 U22731 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n19659) );
  AOI21_X1 U22732 ( .B1(P2_REIP_REG_15__SCAN_IN), .B2(n19652), .A(n19903), 
        .ZN(n19653) );
  OAI21_X1 U22733 ( .B1(n19655), .B2(n19654), .A(n19653), .ZN(n19656) );
  AOI21_X1 U22734 ( .B1(n19657), .B2(n19692), .A(n19656), .ZN(n19658) );
  OAI21_X1 U22735 ( .B1(n19683), .B2(n19659), .A(n19658), .ZN(n19667) );
  OAI21_X1 U22736 ( .B1(n19661), .B2(n19660), .A(n19757), .ZN(n19664) );
  INV_X1 U22737 ( .A(n19662), .ZN(n19663) );
  AOI21_X1 U22738 ( .B1(n19665), .B2(n19664), .A(n19663), .ZN(n19666) );
  AOI211_X1 U22739 ( .C1(n19734), .C2(n19668), .A(n19667), .B(n19666), .ZN(
        n19669) );
  OAI21_X1 U22740 ( .B1(n19726), .B2(n19812), .A(n19669), .ZN(P2_U2840) );
  NOR2_X1 U22741 ( .A1(n19670), .A2(n19672), .ZN(n19671) );
  MUX2_X1 U22742 ( .A(n19672), .B(n19671), .S(n19753), .Z(n19674) );
  OR2_X1 U22743 ( .A1(n19674), .A2(n19673), .ZN(n19681) );
  AOI22_X1 U22744 ( .A1(n19675), .A2(n19734), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19732), .ZN(n19676) );
  OAI211_X1 U22745 ( .C1(n15879), .C2(n19737), .A(n19676), .B(n19736), .ZN(
        n19679) );
  INV_X1 U22746 ( .A(n19780), .ZN(n19677) );
  OAI22_X1 U22747 ( .A1(n19726), .A2(n19825), .B1(n19748), .B2(n19677), .ZN(
        n19678) );
  AOI211_X1 U22748 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n19744), .A(n19679), .B(
        n19678), .ZN(n19680) );
  OAI21_X1 U22749 ( .B1(n19730), .B2(n19681), .A(n19680), .ZN(P2_U2845) );
  OAI21_X1 U22750 ( .B1(n10846), .B2(n19737), .A(n19736), .ZN(n19687) );
  INV_X1 U22751 ( .A(n19682), .ZN(n19685) );
  OAI22_X1 U22752 ( .A1(n19685), .A2(n19684), .B1(n19683), .B2(n10351), .ZN(
        n19686) );
  AOI211_X1 U22753 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19732), .A(
        n19687), .B(n19686), .ZN(n19695) );
  NAND2_X1 U22754 ( .A1(n19753), .A2(n19688), .ZN(n19690) );
  XNOR2_X1 U22755 ( .A(n19690), .B(n19689), .ZN(n19693) );
  AOI22_X1 U22756 ( .A1(n19693), .A2(n19757), .B1(n19692), .B2(n19691), .ZN(
        n19694) );
  OAI211_X1 U22757 ( .C1(n19726), .C2(n19827), .A(n19695), .B(n19694), .ZN(
        P2_U2846) );
  NOR2_X1 U22758 ( .A1(n19710), .A2(n19697), .ZN(n19696) );
  MUX2_X1 U22759 ( .A(n19697), .B(n19696), .S(n19753), .Z(n19699) );
  OR2_X1 U22760 ( .A1(n19699), .A2(n19698), .ZN(n19706) );
  AOI22_X1 U22761 ( .A1(n19700), .A2(n19734), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19732), .ZN(n19701) );
  OAI211_X1 U22762 ( .C1(n10865), .C2(n19737), .A(n19701), .B(n19736), .ZN(
        n19704) );
  OAI22_X1 U22763 ( .A1(n19832), .A2(n19726), .B1(n19748), .B2(n19702), .ZN(
        n19703) );
  AOI211_X1 U22764 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19744), .A(n19704), .B(
        n19703), .ZN(n19705) );
  OAI21_X1 U22765 ( .B1(n19706), .B2(n19730), .A(n19705), .ZN(P2_U2848) );
  NOR2_X1 U22766 ( .A1(n19707), .A2(n19709), .ZN(n19708) );
  MUX2_X1 U22767 ( .A(n19709), .B(n19708), .S(n19753), .Z(n19711) );
  OR2_X1 U22768 ( .A1(n19711), .A2(n19710), .ZN(n19719) );
  INV_X1 U22769 ( .A(n19712), .ZN(n19713) );
  AOI22_X1 U22770 ( .A1(n19744), .A2(P2_EBX_REG_6__SCAN_IN), .B1(n19713), .B2(
        n19734), .ZN(n19714) );
  OAI211_X1 U22771 ( .C1(n10861), .C2(n19737), .A(n19714), .B(n19736), .ZN(
        n19717) );
  OAI22_X1 U22772 ( .A1(n19835), .A2(n19726), .B1(n19748), .B2(n19715), .ZN(
        n19716) );
  AOI211_X1 U22773 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19732), .A(
        n19717), .B(n19716), .ZN(n19718) );
  OAI21_X1 U22774 ( .B1(n19730), .B2(n19719), .A(n19718), .ZN(P2_U2849) );
  NAND2_X1 U22775 ( .A1(n19753), .A2(n19756), .ZN(n19721) );
  XOR2_X1 U22776 ( .A(n19721), .B(n19720), .Z(n19731) );
  INV_X1 U22777 ( .A(n19722), .ZN(n19723) );
  AOI22_X1 U22778 ( .A1(n19744), .A2(P2_EBX_REG_5__SCAN_IN), .B1(n19734), .B2(
        n19723), .ZN(n19724) );
  OAI211_X1 U22779 ( .C1(n14024), .C2(n19737), .A(n19724), .B(n19736), .ZN(
        n19728) );
  OAI22_X1 U22780 ( .A1(n19843), .A2(n19726), .B1(n19748), .B2(n19725), .ZN(
        n19727) );
  AOI211_X1 U22781 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19732), .A(
        n19728), .B(n19727), .ZN(n19729) );
  OAI21_X1 U22782 ( .B1(n19731), .B2(n19730), .A(n19729), .ZN(P2_U2850) );
  AOI22_X1 U22783 ( .A1(n19734), .A2(n19733), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19732), .ZN(n19735) );
  OAI211_X1 U22784 ( .C1(n14003), .C2(n19737), .A(n19736), .B(n19735), .ZN(
        n19738) );
  INV_X1 U22785 ( .A(n19738), .ZN(n19762) );
  NAND2_X1 U22786 ( .A1(n19740), .A2(n19739), .ZN(n19742) );
  AND2_X1 U22787 ( .A1(n19742), .A2(n10147), .ZN(n19910) );
  AOI22_X1 U22788 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19744), .B1(n19743), .B2(
        n19910), .ZN(n19761) );
  OR2_X1 U22789 ( .A1(n19746), .A2(n19745), .ZN(n19747) );
  NAND2_X1 U22790 ( .A1(n13100), .A2(n19747), .ZN(n19847) );
  OAI22_X1 U22791 ( .A1(n19847), .A2(n19749), .B1(n19748), .B2(n19912), .ZN(
        n19750) );
  INV_X1 U22792 ( .A(n19750), .ZN(n19760) );
  OR2_X1 U22793 ( .A1(n19752), .A2(n19751), .ZN(n19754) );
  MUX2_X1 U22794 ( .A(n19755), .B(n19754), .S(n19753), .Z(n19758) );
  NAND3_X1 U22795 ( .A1(n19758), .A2(n19757), .A3(n19756), .ZN(n19759) );
  NAND4_X1 U22796 ( .A1(n19762), .A2(n19761), .A3(n19760), .A4(n19759), .ZN(
        P2_U2851) );
  OR2_X1 U22797 ( .A1(n19764), .A2(n19763), .ZN(n19765) );
  AND2_X1 U22798 ( .A1(n14095), .A2(n19765), .ZN(n19807) );
  AOI22_X1 U22799 ( .A1(n19807), .A2(n19793), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19796), .ZN(n19766) );
  OAI21_X1 U22800 ( .B1(n19796), .B2(n19767), .A(n19766), .ZN(P2_U2871) );
  XOR2_X1 U22801 ( .A(n19769), .B(n19768), .Z(n19770) );
  AOI22_X1 U22802 ( .A1(n19770), .A2(n19793), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19796), .ZN(n19771) );
  OAI21_X1 U22803 ( .B1(n19772), .B2(n19796), .A(n19771), .ZN(P2_U2873) );
  XNOR2_X1 U22804 ( .A(n19774), .B(n19773), .ZN(n19775) );
  AOI22_X1 U22805 ( .A1(n19775), .A2(n19793), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n19796), .ZN(n19776) );
  OAI21_X1 U22806 ( .B1(n19777), .B2(n19796), .A(n19776), .ZN(P2_U2875) );
  XNOR2_X1 U22807 ( .A(n19779), .B(n19778), .ZN(n19781) );
  AOI22_X1 U22808 ( .A1(n19781), .A2(n19793), .B1(n19784), .B2(n19780), .ZN(
        n19782) );
  OAI21_X1 U22809 ( .B1(n19784), .B2(n19783), .A(n19782), .ZN(P2_U2877) );
  AOI211_X1 U22810 ( .C1(n19789), .C2(n9638), .A(n19788), .B(n19787), .ZN(
        n19790) );
  AOI21_X1 U22811 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19796), .A(n19790), .ZN(
        n19791) );
  OAI21_X1 U22812 ( .B1(n19792), .B2(n19796), .A(n19791), .ZN(P2_U2879) );
  INV_X1 U22813 ( .A(n19847), .ZN(n19794) );
  AOI22_X1 U22814 ( .A1(n19794), .A2(n19793), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n19796), .ZN(n19795) );
  OAI21_X1 U22815 ( .B1(n19796), .B2(n19912), .A(n19795), .ZN(P2_U2883) );
  INV_X1 U22816 ( .A(n19797), .ZN(n19798) );
  AOI22_X1 U22817 ( .A1(n19804), .A2(BUF2_REG_31__SCAN_IN), .B1(n19798), .B2(
        n19859), .ZN(n19800) );
  AOI22_X1 U22818 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19858), .B1(n19803), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19799) );
  NAND2_X1 U22819 ( .A1(n19800), .A2(n19799), .ZN(P2_U2888) );
  INV_X1 U22820 ( .A(n19937), .ZN(n19801) );
  AOI22_X1 U22821 ( .A1(n19802), .A2(n19801), .B1(n19858), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19810) );
  AOI22_X1 U22822 ( .A1(n19804), .A2(BUF2_REG_16__SCAN_IN), .B1(n19803), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19809) );
  INV_X1 U22823 ( .A(n19805), .ZN(n19806) );
  AOI22_X1 U22824 ( .A1(n19807), .A2(n19848), .B1(n19859), .B2(n19806), .ZN(
        n19808) );
  NAND3_X1 U22825 ( .A1(n19810), .A2(n19809), .A3(n19808), .ZN(P2_U2903) );
  OAI222_X1 U22826 ( .A1(n19812), .A2(n19844), .B1(n12955), .B2(n19834), .C1(
        n19811), .C2(n19867), .ZN(P2_U2904) );
  AOI22_X1 U22827 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19858), .B1(n19813), 
        .B2(n19836), .ZN(n19814) );
  OAI21_X1 U22828 ( .B1(n19844), .B2(n19815), .A(n19814), .ZN(P2_U2905) );
  INV_X1 U22829 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19874) );
  OAI222_X1 U22830 ( .A1(n19817), .A2(n19844), .B1(n19874), .B2(n19834), .C1(
        n19867), .C2(n19816), .ZN(P2_U2906) );
  AOI22_X1 U22831 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19858), .B1(n19818), 
        .B2(n19836), .ZN(n19819) );
  OAI21_X1 U22832 ( .B1(n19844), .B2(n19820), .A(n19819), .ZN(P2_U2907) );
  INV_X1 U22833 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n21136) );
  OAI222_X1 U22834 ( .A1(n19822), .A2(n19844), .B1(n21136), .B2(n19834), .C1(
        n19867), .C2(n19821), .ZN(P2_U2908) );
  AOI22_X1 U22835 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19858), .B1(n19823), 
        .B2(n19836), .ZN(n19824) );
  OAI21_X1 U22836 ( .B1(n19844), .B2(n19825), .A(n19824), .ZN(P2_U2909) );
  INV_X1 U22837 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19881) );
  OAI222_X1 U22838 ( .A1(n19827), .A2(n19844), .B1(n19881), .B2(n19834), .C1(
        n19867), .C2(n19826), .ZN(P2_U2910) );
  INV_X1 U22839 ( .A(n19828), .ZN(n19830) );
  INV_X1 U22840 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19883) );
  OAI222_X1 U22841 ( .A1(n19830), .A2(n19844), .B1(n19883), .B2(n19834), .C1(
        n19867), .C2(n19829), .ZN(P2_U2911) );
  OAI222_X1 U22842 ( .A1(n19832), .A2(n19844), .B1(n19885), .B2(n19834), .C1(
        n19867), .C2(n19831), .ZN(P2_U2912) );
  INV_X1 U22843 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19887) );
  INV_X1 U22844 ( .A(n19833), .ZN(n19964) );
  OAI222_X1 U22845 ( .A1(n19835), .A2(n19844), .B1(n19887), .B2(n19834), .C1(
        n19867), .C2(n19964), .ZN(P2_U2913) );
  AOI22_X1 U22846 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19858), .B1(n19837), .B2(
        n19836), .ZN(n19842) );
  AOI21_X1 U22847 ( .B1(n20590), .B2(n20054), .A(n19838), .ZN(n19854) );
  XNOR2_X1 U22848 ( .A(n20582), .B(n20584), .ZN(n19853) );
  NOR2_X1 U22849 ( .A1(n19854), .A2(n19853), .ZN(n19852) );
  AOI21_X1 U22850 ( .B1(n20570), .B2(n19839), .A(n19852), .ZN(n19840) );
  NOR2_X1 U22851 ( .A1(n19840), .A2(n19910), .ZN(n19846) );
  OR3_X1 U22852 ( .A1(n19846), .A2(n19847), .A3(n19863), .ZN(n19841) );
  OAI211_X1 U22853 ( .C1(n19844), .C2(n19843), .A(n19842), .B(n19841), .ZN(
        P2_U2914) );
  INV_X1 U22854 ( .A(n19845), .ZN(n19953) );
  AOI22_X1 U22855 ( .A1(n19859), .A2(n19910), .B1(n19858), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19851) );
  XOR2_X1 U22856 ( .A(n19847), .B(n19846), .Z(n19849) );
  NAND2_X1 U22857 ( .A1(n19849), .A2(n19848), .ZN(n19850) );
  OAI211_X1 U22858 ( .C1(n19953), .C2(n19867), .A(n19851), .B(n19850), .ZN(
        P2_U2915) );
  AOI22_X1 U22859 ( .A1(n20584), .A2(n19859), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19858), .ZN(n19857) );
  AOI21_X1 U22860 ( .B1(n19854), .B2(n19853), .A(n19852), .ZN(n19855) );
  OR2_X1 U22861 ( .A1(n19855), .A2(n19863), .ZN(n19856) );
  OAI211_X1 U22862 ( .C1(n19947), .C2(n19867), .A(n19857), .B(n19856), .ZN(
        P2_U2916) );
  AOI22_X1 U22863 ( .A1(n19859), .A2(n20603), .B1(n19858), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19866) );
  AOI21_X1 U22864 ( .B1(n19862), .B2(n19861), .A(n19860), .ZN(n19864) );
  OR2_X1 U22865 ( .A1(n19864), .A2(n19863), .ZN(n19865) );
  OAI211_X1 U22866 ( .C1(n19868), .C2(n19867), .A(n19866), .B(n19865), .ZN(
        P2_U2918) );
  AND2_X1 U22867 ( .A1(n19889), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22868 ( .A1(n19900), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19870) );
  OAI21_X1 U22869 ( .B1(n12955), .B2(n19902), .A(n19870), .ZN(P2_U2936) );
  AOI22_X1 U22870 ( .A1(n19900), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19871) );
  OAI21_X1 U22871 ( .B1(n19872), .B2(n19902), .A(n19871), .ZN(P2_U2937) );
  AOI22_X1 U22872 ( .A1(n19900), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19873) );
  OAI21_X1 U22873 ( .B1(n19874), .B2(n19902), .A(n19873), .ZN(P2_U2938) );
  AOI22_X1 U22874 ( .A1(n19892), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19875) );
  OAI21_X1 U22875 ( .B1(n19876), .B2(n19902), .A(n19875), .ZN(P2_U2939) );
  AOI22_X1 U22876 ( .A1(n19892), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19877) );
  OAI21_X1 U22877 ( .B1(n21136), .B2(n19902), .A(n19877), .ZN(P2_U2940) );
  AOI22_X1 U22878 ( .A1(n19892), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19878) );
  OAI21_X1 U22879 ( .B1(n19879), .B2(n19902), .A(n19878), .ZN(P2_U2941) );
  AOI22_X1 U22880 ( .A1(n19892), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19880) );
  OAI21_X1 U22881 ( .B1(n19881), .B2(n19902), .A(n19880), .ZN(P2_U2942) );
  AOI22_X1 U22882 ( .A1(n19892), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19882) );
  OAI21_X1 U22883 ( .B1(n19883), .B2(n19902), .A(n19882), .ZN(P2_U2943) );
  AOI22_X1 U22884 ( .A1(n19892), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19884) );
  OAI21_X1 U22885 ( .B1(n19885), .B2(n19902), .A(n19884), .ZN(P2_U2944) );
  AOI22_X1 U22886 ( .A1(n19892), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19886) );
  OAI21_X1 U22887 ( .B1(n19887), .B2(n19902), .A(n19886), .ZN(P2_U2945) );
  INV_X1 U22888 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n21072) );
  AOI22_X1 U22889 ( .A1(n19892), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19888) );
  OAI21_X1 U22890 ( .B1(n21072), .B2(n19902), .A(n19888), .ZN(P2_U2946) );
  INV_X1 U22891 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19891) );
  AOI22_X1 U22892 ( .A1(n19892), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19889), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19890) );
  OAI21_X1 U22893 ( .B1(n19891), .B2(n19902), .A(n19890), .ZN(P2_U2947) );
  INV_X1 U22894 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U22895 ( .A1(n19892), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19893) );
  OAI21_X1 U22896 ( .B1(n19894), .B2(n19902), .A(n19893), .ZN(P2_U2948) );
  AOI22_X1 U22897 ( .A1(n19900), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19895) );
  OAI21_X1 U22898 ( .B1(n19896), .B2(n19902), .A(n19895), .ZN(P2_U2949) );
  INV_X1 U22899 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19898) );
  AOI22_X1 U22900 ( .A1(n19900), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19897) );
  OAI21_X1 U22901 ( .B1(n19898), .B2(n19902), .A(n19897), .ZN(P2_U2950) );
  AOI22_X1 U22902 ( .A1(n19900), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19899), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19901) );
  OAI21_X1 U22903 ( .B1(n12957), .B2(n19902), .A(n19901), .ZN(P2_U2951) );
  NAND2_X1 U22904 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19903), .ZN(n19904) );
  OAI221_X1 U22905 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19907), .C1(
        n19906), .C2(n19905), .A(n19904), .ZN(n19908) );
  AOI21_X1 U22906 ( .B1(n19910), .B2(n19909), .A(n19908), .ZN(n19916) );
  NOR2_X1 U22907 ( .A1(n19912), .A2(n19911), .ZN(n19913) );
  AOI21_X1 U22908 ( .B1(n19914), .B2(n19920), .A(n19913), .ZN(n19915) );
  OAI211_X1 U22909 ( .C1(n19926), .C2(n19917), .A(n19916), .B(n19915), .ZN(
        P2_U3042) );
  NAND2_X1 U22910 ( .A1(n19919), .A2(n19918), .ZN(n19934) );
  NAND2_X1 U22911 ( .A1(n19921), .A2(n19920), .ZN(n19923) );
  OAI211_X1 U22912 ( .C1(n19925), .C2(n19924), .A(n19923), .B(n19922), .ZN(
        n19930) );
  OAI22_X1 U22913 ( .A1(n20590), .A2(n19928), .B1(n19927), .B2(n19926), .ZN(
        n19929) );
  NAND2_X1 U22914 ( .A1(n19932), .A2(n19934), .ZN(n19933) );
  OAI211_X1 U22915 ( .C1(n19935), .C2(n19934), .A(n9708), .B(n19933), .ZN(
        P2_U3044) );
  AOI22_X1 U22916 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19965), .ZN(n20364) );
  INV_X1 U22917 ( .A(n20364), .ZN(n20435) );
  AND2_X1 U22918 ( .A1(n19936), .A2(n19951), .ZN(n20434) );
  AOI22_X1 U22919 ( .A1(n20435), .A2(n20481), .B1(n19963), .B2(n20434), .ZN(
        n19940) );
  AOI22_X1 U22920 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19965), .ZN(n20326) );
  AOI22_X1 U22921 ( .A1(n19938), .A2(n19967), .B1(n19995), .B2(n20436), .ZN(
        n19939) );
  OAI211_X1 U22922 ( .C1(n19971), .C2(n19941), .A(n19940), .B(n19939), .ZN(
        P2_U3048) );
  AOI22_X1 U22923 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19965), .ZN(n20370) );
  INV_X1 U22924 ( .A(n20370), .ZN(n20446) );
  NOR2_X2 U22925 ( .A1(n10444), .A2(n19961), .ZN(n20444) );
  AOI22_X1 U22926 ( .A1(n20446), .A2(n20481), .B1(n19963), .B2(n20444), .ZN(
        n19944) );
  NOR2_X2 U22927 ( .A1(n19942), .A2(n20395), .ZN(n20445) );
  AOI22_X1 U22928 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19965), .ZN(n20332) );
  AOI22_X1 U22929 ( .A1(n20445), .A2(n19967), .B1(n19995), .B2(n20447), .ZN(
        n19943) );
  OAI211_X1 U22930 ( .C1(n19971), .C2(n19945), .A(n19944), .B(n19943), .ZN(
        P2_U3050) );
  AOI22_X1 U22931 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19965), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19966), .ZN(n20373) );
  AOI22_X1 U22932 ( .A1(n20452), .A2(n20481), .B1(n19963), .B2(n20450), .ZN(
        n19949) );
  NOR2_X2 U22933 ( .A1(n19947), .A2(n20395), .ZN(n20451) );
  AOI22_X1 U22934 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19965), .ZN(n20335) );
  AOI22_X1 U22935 ( .A1(n20451), .A2(n19967), .B1(n19995), .B2(n20453), .ZN(
        n19948) );
  OAI211_X1 U22936 ( .C1(n19971), .C2(n19950), .A(n19949), .B(n19948), .ZN(
        P2_U3051) );
  AOI22_X1 U22937 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19965), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19966), .ZN(n20376) );
  AOI22_X1 U22938 ( .A1(n20460), .A2(n20481), .B1(n19963), .B2(n20457), .ZN(
        n19955) );
  NOR2_X2 U22939 ( .A1(n19953), .A2(n20395), .ZN(n20458) );
  AOI22_X1 U22940 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19965), .ZN(n20338) );
  INV_X1 U22941 ( .A(n20338), .ZN(n20459) );
  AOI22_X1 U22942 ( .A1(n20458), .A2(n19967), .B1(n19995), .B2(n20459), .ZN(
        n19954) );
  OAI211_X1 U22943 ( .C1(n19971), .C2(n19956), .A(n19955), .B(n19954), .ZN(
        P2_U3052) );
  AOI22_X1 U22944 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19965), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19966), .ZN(n20379) );
  NOR2_X2 U22945 ( .A1(n10773), .A2(n19961), .ZN(n20464) );
  AOI22_X1 U22946 ( .A1(n20467), .A2(n20481), .B1(n19963), .B2(n20464), .ZN(
        n19959) );
  NOR2_X2 U22947 ( .A1(n19957), .A2(n20395), .ZN(n20465) );
  AOI22_X1 U22948 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19965), .ZN(n20341) );
  AOI22_X1 U22949 ( .A1(n20465), .A2(n19967), .B1(n19995), .B2(n20466), .ZN(
        n19958) );
  OAI211_X1 U22950 ( .C1(n19971), .C2(n19960), .A(n19959), .B(n19958), .ZN(
        P2_U3053) );
  AOI22_X1 U22951 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19965), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19966), .ZN(n20382) );
  NOR2_X2 U22952 ( .A1(n19962), .A2(n19961), .ZN(n20470) );
  AOI22_X1 U22953 ( .A1(n20473), .A2(n20481), .B1(n19963), .B2(n20470), .ZN(
        n19969) );
  NOR2_X2 U22954 ( .A1(n19964), .A2(n20395), .ZN(n20471) );
  AOI22_X1 U22955 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19966), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19965), .ZN(n20344) );
  INV_X1 U22956 ( .A(n20344), .ZN(n20472) );
  AOI22_X1 U22957 ( .A1(n20471), .A2(n19967), .B1(n19995), .B2(n20472), .ZN(
        n19968) );
  OAI211_X1 U22958 ( .C1(n19971), .C2(n19970), .A(n19969), .B(n19968), .ZN(
        P2_U3054) );
  NOR2_X1 U22959 ( .A1(n20221), .A2(n20021), .ZN(n19993) );
  INV_X1 U22960 ( .A(n19993), .ZN(n19972) );
  AND2_X1 U22961 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19972), .ZN(n19973) );
  NAND2_X1 U22962 ( .A1(n10594), .A2(n19973), .ZN(n19976) );
  AOI21_X1 U22963 ( .B1(n20491), .B2(n19975), .A(n20489), .ZN(n19974) );
  AND2_X1 U22964 ( .A1(n19976), .A2(n19974), .ZN(n19994) );
  AOI22_X1 U22965 ( .A1(n19994), .A2(n19938), .B1(n20434), .B2(n19993), .ZN(
        n19980) );
  NAND2_X1 U22966 ( .A1(n20570), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20143) );
  OAI21_X1 U22967 ( .B1(n20143), .B2(n20222), .A(n19975), .ZN(n19977) );
  AND2_X1 U22968 ( .A1(n19977), .A2(n19976), .ZN(n19978) );
  OAI211_X1 U22969 ( .C1(n19993), .C2(n21204), .A(n19978), .B(n20425), .ZN(
        n19996) );
  AOI22_X1 U22970 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19996), .B1(
        n19995), .B2(n20435), .ZN(n19979) );
  OAI211_X1 U22971 ( .C1(n20326), .C2(n19999), .A(n19980), .B(n19979), .ZN(
        P2_U3056) );
  AOI22_X1 U22972 ( .A1(n19994), .A2(n13863), .B1(n20439), .B2(n19993), .ZN(
        n19982) );
  AOI22_X1 U22973 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19996), .B1(
        n19995), .B2(n20441), .ZN(n19981) );
  OAI211_X1 U22974 ( .C1(n20329), .C2(n19999), .A(n19982), .B(n19981), .ZN(
        P2_U3057) );
  AOI22_X1 U22975 ( .A1(n19994), .A2(n20445), .B1(n20444), .B2(n19993), .ZN(
        n19984) );
  AOI22_X1 U22976 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19996), .B1(
        n19995), .B2(n20446), .ZN(n19983) );
  OAI211_X1 U22977 ( .C1(n20332), .C2(n19999), .A(n19984), .B(n19983), .ZN(
        P2_U3058) );
  AOI22_X1 U22978 ( .A1(n19994), .A2(n20451), .B1(n20450), .B2(n19993), .ZN(
        n19986) );
  AOI22_X1 U22979 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19996), .B1(
        n19995), .B2(n20452), .ZN(n19985) );
  OAI211_X1 U22980 ( .C1(n20335), .C2(n19999), .A(n19986), .B(n19985), .ZN(
        P2_U3059) );
  AOI22_X1 U22981 ( .A1(n19994), .A2(n20458), .B1(n20457), .B2(n19993), .ZN(
        n19988) );
  AOI22_X1 U22982 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19996), .B1(
        n19995), .B2(n20460), .ZN(n19987) );
  OAI211_X1 U22983 ( .C1(n20338), .C2(n19999), .A(n19988), .B(n19987), .ZN(
        P2_U3060) );
  AOI22_X1 U22984 ( .A1(n19994), .A2(n20465), .B1(n20464), .B2(n19993), .ZN(
        n19990) );
  AOI22_X1 U22985 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19996), .B1(
        n19995), .B2(n20467), .ZN(n19989) );
  OAI211_X1 U22986 ( .C1(n20341), .C2(n19999), .A(n19990), .B(n19989), .ZN(
        P2_U3061) );
  AOI22_X1 U22987 ( .A1(n19994), .A2(n20471), .B1(n20470), .B2(n19993), .ZN(
        n19992) );
  AOI22_X1 U22988 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19996), .B1(
        n19995), .B2(n20473), .ZN(n19991) );
  OAI211_X1 U22989 ( .C1(n20344), .C2(n19999), .A(n19992), .B(n19991), .ZN(
        P2_U3062) );
  AOI22_X1 U22990 ( .A1(n19994), .A2(n20478), .B1(n20476), .B2(n19993), .ZN(
        n19998) );
  AOI22_X1 U22991 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19996), .B1(
        n19995), .B2(n20482), .ZN(n19997) );
  OAI211_X1 U22992 ( .C1(n20351), .C2(n19999), .A(n19998), .B(n19997), .ZN(
        P2_U3063) );
  AOI22_X1 U22993 ( .A1(n20015), .A2(n19938), .B1(n20014), .B2(n20434), .ZN(
        n20001) );
  AOI22_X1 U22994 ( .A1(n20042), .A2(n20436), .B1(n20016), .B2(n20435), .ZN(
        n20000) );
  OAI211_X1 U22995 ( .C1(n20020), .C2(n12413), .A(n20001), .B(n20000), .ZN(
        P2_U3064) );
  AOI22_X1 U22996 ( .A1(n20015), .A2(n20445), .B1(n20014), .B2(n20444), .ZN(
        n20003) );
  AOI22_X1 U22997 ( .A1(n20042), .A2(n20447), .B1(n20016), .B2(n20446), .ZN(
        n20002) );
  OAI211_X1 U22998 ( .C1(n20020), .C2(n12338), .A(n20003), .B(n20002), .ZN(
        P2_U3066) );
  AOI22_X1 U22999 ( .A1(n20015), .A2(n20451), .B1(n20014), .B2(n20450), .ZN(
        n20005) );
  AOI22_X1 U23000 ( .A1(n20042), .A2(n20453), .B1(n20016), .B2(n20452), .ZN(
        n20004) );
  OAI211_X1 U23001 ( .C1(n20020), .C2(n10579), .A(n20005), .B(n20004), .ZN(
        P2_U3067) );
  INV_X1 U23002 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n20008) );
  AOI22_X1 U23003 ( .A1(n20015), .A2(n20458), .B1(n20014), .B2(n20457), .ZN(
        n20007) );
  AOI22_X1 U23004 ( .A1(n20016), .A2(n20460), .B1(n20042), .B2(n20459), .ZN(
        n20006) );
  OAI211_X1 U23005 ( .C1(n20020), .C2(n20008), .A(n20007), .B(n20006), .ZN(
        P2_U3068) );
  INV_X1 U23006 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n20011) );
  AOI22_X1 U23007 ( .A1(n20015), .A2(n20465), .B1(n20014), .B2(n20464), .ZN(
        n20010) );
  AOI22_X1 U23008 ( .A1(n20016), .A2(n20467), .B1(n20042), .B2(n20466), .ZN(
        n20009) );
  OAI211_X1 U23009 ( .C1(n20020), .C2(n20011), .A(n20010), .B(n20009), .ZN(
        P2_U3069) );
  AOI22_X1 U23010 ( .A1(n20015), .A2(n20471), .B1(n20014), .B2(n20470), .ZN(
        n20013) );
  AOI22_X1 U23011 ( .A1(n20016), .A2(n20473), .B1(n20042), .B2(n20472), .ZN(
        n20012) );
  OAI211_X1 U23012 ( .C1(n20020), .C2(n10646), .A(n20013), .B(n20012), .ZN(
        P2_U3070) );
  AOI22_X1 U23013 ( .A1(n20015), .A2(n20478), .B1(n20014), .B2(n20476), .ZN(
        n20018) );
  AOI22_X1 U23014 ( .A1(n20016), .A2(n20482), .B1(n20042), .B2(n20480), .ZN(
        n20017) );
  OAI211_X1 U23015 ( .C1(n20020), .C2(n20019), .A(n20018), .B(n20017), .ZN(
        P2_U3071) );
  NOR2_X1 U23016 ( .A1(n20286), .A2(n20021), .ZN(n20045) );
  AOI22_X1 U23017 ( .A1(n20436), .A2(n20071), .B1(n20045), .B2(n20434), .ZN(
        n20031) );
  OAI21_X1 U23018 ( .B1(n20143), .B2(n20576), .A(n20585), .ZN(n20029) );
  NOR2_X1 U23019 ( .A1(n20605), .A2(n20021), .ZN(n20025) );
  INV_X1 U23020 ( .A(n20045), .ZN(n20022) );
  OAI211_X1 U23021 ( .C1(n20023), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20022), 
        .B(n20578), .ZN(n20024) );
  OAI211_X1 U23022 ( .C1(n20029), .C2(n20025), .A(n20425), .B(n20024), .ZN(
        n20047) );
  INV_X1 U23023 ( .A(n20025), .ZN(n20028) );
  OAI21_X1 U23024 ( .B1(n20026), .B2(n20045), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20027) );
  AOI22_X1 U23025 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20047), .B1(
        n19938), .B2(n20046), .ZN(n20030) );
  OAI211_X1 U23026 ( .C1(n20364), .C2(n20050), .A(n20031), .B(n20030), .ZN(
        P2_U3072) );
  AOI22_X1 U23027 ( .A1(n20441), .A2(n20042), .B1(n20439), .B2(n20045), .ZN(
        n20033) );
  AOI22_X1 U23028 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20047), .B1(
        n13863), .B2(n20046), .ZN(n20032) );
  OAI211_X1 U23029 ( .C1(n20329), .C2(n20079), .A(n20033), .B(n20032), .ZN(
        P2_U3073) );
  AOI22_X1 U23030 ( .A1(n20447), .A2(n20071), .B1(n20045), .B2(n20444), .ZN(
        n20035) );
  AOI22_X1 U23031 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20047), .B1(
        n20445), .B2(n20046), .ZN(n20034) );
  OAI211_X1 U23032 ( .C1(n20370), .C2(n20050), .A(n20035), .B(n20034), .ZN(
        P2_U3074) );
  AOI22_X1 U23033 ( .A1(n20453), .A2(n20071), .B1(n20045), .B2(n20450), .ZN(
        n20037) );
  AOI22_X1 U23034 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20047), .B1(
        n20451), .B2(n20046), .ZN(n20036) );
  OAI211_X1 U23035 ( .C1(n20373), .C2(n20050), .A(n20037), .B(n20036), .ZN(
        P2_U3075) );
  AOI22_X1 U23036 ( .A1(n20459), .A2(n20071), .B1(n20045), .B2(n20457), .ZN(
        n20039) );
  AOI22_X1 U23037 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20047), .B1(
        n20458), .B2(n20046), .ZN(n20038) );
  OAI211_X1 U23038 ( .C1(n20376), .C2(n20050), .A(n20039), .B(n20038), .ZN(
        P2_U3076) );
  AOI22_X1 U23039 ( .A1(n20466), .A2(n20071), .B1(n20045), .B2(n20464), .ZN(
        n20041) );
  AOI22_X1 U23040 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20047), .B1(
        n20465), .B2(n20046), .ZN(n20040) );
  OAI211_X1 U23041 ( .C1(n20379), .C2(n20050), .A(n20041), .B(n20040), .ZN(
        P2_U3077) );
  AOI22_X1 U23042 ( .A1(n20473), .A2(n20042), .B1(n20045), .B2(n20470), .ZN(
        n20044) );
  AOI22_X1 U23043 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20047), .B1(
        n20471), .B2(n20046), .ZN(n20043) );
  OAI211_X1 U23044 ( .C1(n20344), .C2(n20079), .A(n20044), .B(n20043), .ZN(
        P2_U3078) );
  AOI22_X1 U23045 ( .A1(n20480), .A2(n20071), .B1(n20476), .B2(n20045), .ZN(
        n20049) );
  AOI22_X1 U23046 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20047), .B1(
        n20478), .B2(n20046), .ZN(n20048) );
  OAI211_X1 U23047 ( .C1(n20388), .C2(n20050), .A(n20049), .B(n20048), .ZN(
        P2_U3079) );
  NOR2_X1 U23048 ( .A1(n20052), .A2(n20051), .ZN(n20317) );
  NAND2_X1 U23049 ( .A1(n20317), .A2(n20588), .ZN(n20057) );
  OR2_X1 U23050 ( .A1(n20057), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20053) );
  NAND2_X1 U23051 ( .A1(n20588), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20134) );
  NOR2_X1 U23052 ( .A1(n20134), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20082) );
  INV_X1 U23053 ( .A(n20082), .ZN(n20085) );
  NOR2_X1 U23054 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20085), .ZN(
        n20074) );
  NOR3_X1 U23055 ( .A1(n10598), .A2(n20074), .A3(n20491), .ZN(n20055) );
  AOI21_X1 U23056 ( .B1(n20491), .B2(n20053), .A(n20055), .ZN(n20075) );
  AOI22_X1 U23057 ( .A1(n20075), .A2(n19938), .B1(n20434), .B2(n20074), .ZN(
        n20060) );
  OAI21_X1 U23058 ( .B1(n20071), .B2(n20102), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20056) );
  AOI211_X1 U23059 ( .C1(n20057), .C2(n20056), .A(n20395), .B(n20055), .ZN(
        n20058) );
  AOI22_X1 U23060 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20076), .B1(
        n20102), .B2(n20436), .ZN(n20059) );
  OAI211_X1 U23061 ( .C1(n20364), .C2(n20079), .A(n20060), .B(n20059), .ZN(
        P2_U3080) );
  AOI22_X1 U23062 ( .A1(n20075), .A2(n13863), .B1(n20439), .B2(n20074), .ZN(
        n20062) );
  AOI22_X1 U23063 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20076), .B1(
        n20071), .B2(n20441), .ZN(n20061) );
  OAI211_X1 U23064 ( .C1(n20329), .C2(n20099), .A(n20062), .B(n20061), .ZN(
        P2_U3081) );
  AOI22_X1 U23065 ( .A1(n20075), .A2(n20445), .B1(n20444), .B2(n20074), .ZN(
        n20064) );
  AOI22_X1 U23066 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20076), .B1(
        n20102), .B2(n20447), .ZN(n20063) );
  OAI211_X1 U23067 ( .C1(n20370), .C2(n20079), .A(n20064), .B(n20063), .ZN(
        P2_U3082) );
  AOI22_X1 U23068 ( .A1(n20075), .A2(n20451), .B1(n20450), .B2(n20074), .ZN(
        n20066) );
  AOI22_X1 U23069 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20076), .B1(
        n20102), .B2(n20453), .ZN(n20065) );
  OAI211_X1 U23070 ( .C1(n20373), .C2(n20079), .A(n20066), .B(n20065), .ZN(
        P2_U3083) );
  AOI22_X1 U23071 ( .A1(n20075), .A2(n20458), .B1(n20457), .B2(n20074), .ZN(
        n20068) );
  AOI22_X1 U23072 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20076), .B1(
        n20102), .B2(n20459), .ZN(n20067) );
  OAI211_X1 U23073 ( .C1(n20376), .C2(n20079), .A(n20068), .B(n20067), .ZN(
        P2_U3084) );
  AOI22_X1 U23074 ( .A1(n20075), .A2(n20465), .B1(n20464), .B2(n20074), .ZN(
        n20070) );
  AOI22_X1 U23075 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20076), .B1(
        n20071), .B2(n20467), .ZN(n20069) );
  OAI211_X1 U23076 ( .C1(n20341), .C2(n20099), .A(n20070), .B(n20069), .ZN(
        P2_U3085) );
  AOI22_X1 U23077 ( .A1(n20075), .A2(n20471), .B1(n20470), .B2(n20074), .ZN(
        n20073) );
  AOI22_X1 U23078 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20076), .B1(
        n20071), .B2(n20473), .ZN(n20072) );
  OAI211_X1 U23079 ( .C1(n20344), .C2(n20099), .A(n20073), .B(n20072), .ZN(
        P2_U3086) );
  AOI22_X1 U23080 ( .A1(n20075), .A2(n20478), .B1(n20476), .B2(n20074), .ZN(
        n20078) );
  AOI22_X1 U23081 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20076), .B1(
        n20102), .B2(n20480), .ZN(n20077) );
  OAI211_X1 U23082 ( .C1(n20388), .C2(n20079), .A(n20078), .B(n20077), .ZN(
        P2_U3087) );
  NOR2_X1 U23083 ( .A1(n20221), .A2(n20134), .ZN(n20109) );
  AOI22_X1 U23084 ( .A1(n20435), .A2(n20102), .B1(n20109), .B2(n20434), .ZN(
        n20088) );
  OAI21_X1 U23085 ( .B1(n20143), .B2(n20360), .A(n20585), .ZN(n20086) );
  INV_X1 U23086 ( .A(n20109), .ZN(n20080) );
  OAI211_X1 U23087 ( .C1(n10599), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20080), 
        .B(n20578), .ZN(n20081) );
  OAI211_X1 U23088 ( .C1(n20086), .C2(n20082), .A(n20425), .B(n20081), .ZN(
        n20104) );
  OAI21_X1 U23089 ( .B1(n20083), .B2(n20109), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20084) );
  AOI22_X1 U23090 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20104), .B1(
        n19938), .B2(n20103), .ZN(n20087) );
  OAI211_X1 U23091 ( .C1(n20326), .C2(n20133), .A(n20088), .B(n20087), .ZN(
        P2_U3088) );
  AOI22_X1 U23092 ( .A1(n20440), .A2(n20125), .B1(n20439), .B2(n20109), .ZN(
        n20090) );
  AOI22_X1 U23093 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20104), .B1(
        n13863), .B2(n20103), .ZN(n20089) );
  OAI211_X1 U23094 ( .C1(n20367), .C2(n20099), .A(n20090), .B(n20089), .ZN(
        P2_U3089) );
  AOI22_X1 U23095 ( .A1(n20447), .A2(n20125), .B1(n20109), .B2(n20444), .ZN(
        n20092) );
  AOI22_X1 U23096 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20104), .B1(
        n20445), .B2(n20103), .ZN(n20091) );
  OAI211_X1 U23097 ( .C1(n20370), .C2(n20099), .A(n20092), .B(n20091), .ZN(
        P2_U3090) );
  AOI22_X1 U23098 ( .A1(n20452), .A2(n20102), .B1(n20109), .B2(n20450), .ZN(
        n20094) );
  AOI22_X1 U23099 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20104), .B1(
        n20451), .B2(n20103), .ZN(n20093) );
  OAI211_X1 U23100 ( .C1(n20335), .C2(n20133), .A(n20094), .B(n20093), .ZN(
        P2_U3091) );
  AOI22_X1 U23101 ( .A1(n20460), .A2(n20102), .B1(n20109), .B2(n20457), .ZN(
        n20096) );
  AOI22_X1 U23102 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20104), .B1(
        n20458), .B2(n20103), .ZN(n20095) );
  OAI211_X1 U23103 ( .C1(n20338), .C2(n20133), .A(n20096), .B(n20095), .ZN(
        P2_U3092) );
  AOI22_X1 U23104 ( .A1(n20466), .A2(n20125), .B1(n20109), .B2(n20464), .ZN(
        n20098) );
  AOI22_X1 U23105 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20104), .B1(
        n20465), .B2(n20103), .ZN(n20097) );
  OAI211_X1 U23106 ( .C1(n20379), .C2(n20099), .A(n20098), .B(n20097), .ZN(
        P2_U3093) );
  AOI22_X1 U23107 ( .A1(n20473), .A2(n20102), .B1(n20109), .B2(n20470), .ZN(
        n20101) );
  AOI22_X1 U23108 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20104), .B1(
        n20471), .B2(n20103), .ZN(n20100) );
  OAI211_X1 U23109 ( .C1(n20344), .C2(n20133), .A(n20101), .B(n20100), .ZN(
        P2_U3094) );
  AOI22_X1 U23110 ( .A1(n20482), .A2(n20102), .B1(n20476), .B2(n20109), .ZN(
        n20106) );
  AOI22_X1 U23111 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20104), .B1(
        n20478), .B2(n20103), .ZN(n20105) );
  OAI211_X1 U23112 ( .C1(n20351), .C2(n20133), .A(n20106), .B(n20105), .ZN(
        P2_U3095) );
  NOR2_X1 U23113 ( .A1(n20257), .A2(n20134), .ZN(n20128) );
  OAI21_X1 U23114 ( .B1(n10664), .B2(n20128), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20107) );
  OAI21_X1 U23115 ( .B1(n20134), .B2(n20262), .A(n20107), .ZN(n20129) );
  AOI22_X1 U23116 ( .A1(n20129), .A2(n19938), .B1(n20434), .B2(n20128), .ZN(
        n20114) );
  AOI221_X1 U23117 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20125), .C1(
        P2_STATEBS16_REG_SCAN_IN), .C2(n20187), .A(n20109), .ZN(n20110) );
  AOI211_X1 U23118 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20111), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20110), .ZN(n20112) );
  AOI22_X1 U23119 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20130), .B1(
        n20187), .B2(n20436), .ZN(n20113) );
  OAI211_X1 U23120 ( .C1(n20364), .C2(n20133), .A(n20114), .B(n20113), .ZN(
        P2_U3096) );
  AOI22_X1 U23121 ( .A1(n20129), .A2(n13863), .B1(n20439), .B2(n20128), .ZN(
        n20116) );
  AOI22_X1 U23122 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20130), .B1(
        n20125), .B2(n20441), .ZN(n20115) );
  OAI211_X1 U23123 ( .C1(n20329), .C2(n20177), .A(n20116), .B(n20115), .ZN(
        P2_U3097) );
  AOI22_X1 U23124 ( .A1(n20129), .A2(n20445), .B1(n20444), .B2(n20128), .ZN(
        n20118) );
  AOI22_X1 U23125 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20130), .B1(
        n20187), .B2(n20447), .ZN(n20117) );
  OAI211_X1 U23126 ( .C1(n20370), .C2(n20133), .A(n20118), .B(n20117), .ZN(
        P2_U3098) );
  AOI22_X1 U23127 ( .A1(n20129), .A2(n20451), .B1(n20450), .B2(n20128), .ZN(
        n20120) );
  AOI22_X1 U23128 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20130), .B1(
        n20187), .B2(n20453), .ZN(n20119) );
  OAI211_X1 U23129 ( .C1(n20373), .C2(n20133), .A(n20120), .B(n20119), .ZN(
        P2_U3099) );
  AOI22_X1 U23130 ( .A1(n20129), .A2(n20458), .B1(n20457), .B2(n20128), .ZN(
        n20122) );
  AOI22_X1 U23131 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20130), .B1(
        n20125), .B2(n20460), .ZN(n20121) );
  OAI211_X1 U23132 ( .C1(n20338), .C2(n20177), .A(n20122), .B(n20121), .ZN(
        P2_U3100) );
  AOI22_X1 U23133 ( .A1(n20129), .A2(n20465), .B1(n20464), .B2(n20128), .ZN(
        n20124) );
  AOI22_X1 U23134 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20130), .B1(
        n20187), .B2(n20466), .ZN(n20123) );
  OAI211_X1 U23135 ( .C1(n20379), .C2(n20133), .A(n20124), .B(n20123), .ZN(
        P2_U3101) );
  AOI22_X1 U23136 ( .A1(n20129), .A2(n20471), .B1(n20470), .B2(n20128), .ZN(
        n20127) );
  AOI22_X1 U23137 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20130), .B1(
        n20125), .B2(n20473), .ZN(n20126) );
  OAI211_X1 U23138 ( .C1(n20344), .C2(n20177), .A(n20127), .B(n20126), .ZN(
        P2_U3102) );
  AOI22_X1 U23139 ( .A1(n20129), .A2(n20478), .B1(n20476), .B2(n20128), .ZN(
        n20132) );
  AOI22_X1 U23140 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20130), .B1(
        n20187), .B2(n20480), .ZN(n20131) );
  OAI211_X1 U23141 ( .C1(n20388), .C2(n20133), .A(n20132), .B(n20131), .ZN(
        P2_U3103) );
  INV_X1 U23142 ( .A(n20286), .ZN(n20136) );
  INV_X1 U23143 ( .A(n20134), .ZN(n20135) );
  NAND2_X1 U23144 ( .A1(n20136), .A2(n20135), .ZN(n20194) );
  NAND2_X1 U23145 ( .A1(n20194), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20137) );
  NAND2_X1 U23146 ( .A1(n20393), .A2(n20588), .ZN(n20144) );
  AOI21_X1 U23147 ( .B1(n20491), .B2(n20144), .A(n20489), .ZN(n20139) );
  NAND2_X1 U23148 ( .A1(n20146), .A2(n20139), .ZN(n20185) );
  INV_X1 U23149 ( .A(n19938), .ZN(n20141) );
  INV_X1 U23150 ( .A(n20434), .ZN(n20140) );
  OAI22_X1 U23151 ( .A1(n20185), .A2(n20141), .B1(n20194), .B2(n20140), .ZN(
        n20142) );
  INV_X1 U23152 ( .A(n20142), .ZN(n20151) );
  OR2_X1 U23153 ( .A1(n20429), .A2(n20143), .ZN(n20575) );
  AOI22_X1 U23154 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20194), .B1(n20575), 
        .B2(n20144), .ZN(n20145) );
  NAND3_X1 U23155 ( .A1(n20146), .A2(n20425), .A3(n20145), .ZN(n20188) );
  INV_X1 U23156 ( .A(n20147), .ZN(n20149) );
  INV_X1 U23157 ( .A(n20429), .ZN(n20148) );
  AOI22_X1 U23158 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20188), .B1(
        n20216), .B2(n20436), .ZN(n20150) );
  OAI211_X1 U23159 ( .C1(n20364), .C2(n20177), .A(n20151), .B(n20150), .ZN(
        P2_U3104) );
  INV_X1 U23160 ( .A(n13863), .ZN(n20153) );
  INV_X1 U23161 ( .A(n20439), .ZN(n20152) );
  OAI22_X1 U23162 ( .A1(n20185), .A2(n20153), .B1(n20152), .B2(n20194), .ZN(
        n20154) );
  INV_X1 U23163 ( .A(n20154), .ZN(n20156) );
  AOI22_X1 U23164 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20188), .B1(
        n20187), .B2(n20441), .ZN(n20155) );
  OAI211_X1 U23165 ( .C1(n20329), .C2(n20208), .A(n20156), .B(n20155), .ZN(
        P2_U3105) );
  INV_X1 U23166 ( .A(n20445), .ZN(n20158) );
  INV_X1 U23167 ( .A(n20444), .ZN(n20157) );
  OAI22_X1 U23168 ( .A1(n20185), .A2(n20158), .B1(n20194), .B2(n20157), .ZN(
        n20159) );
  INV_X1 U23169 ( .A(n20159), .ZN(n20161) );
  AOI22_X1 U23170 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20188), .B1(
        n20187), .B2(n20446), .ZN(n20160) );
  OAI211_X1 U23171 ( .C1(n20332), .C2(n20208), .A(n20161), .B(n20160), .ZN(
        P2_U3106) );
  INV_X1 U23172 ( .A(n20451), .ZN(n20163) );
  INV_X1 U23173 ( .A(n20450), .ZN(n20162) );
  OAI22_X1 U23174 ( .A1(n20185), .A2(n20163), .B1(n20194), .B2(n20162), .ZN(
        n20164) );
  INV_X1 U23175 ( .A(n20164), .ZN(n20166) );
  AOI22_X1 U23176 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20188), .B1(
        n20187), .B2(n20452), .ZN(n20165) );
  OAI211_X1 U23177 ( .C1(n20335), .C2(n20208), .A(n20166), .B(n20165), .ZN(
        P2_U3107) );
  INV_X1 U23178 ( .A(n20458), .ZN(n20168) );
  INV_X1 U23179 ( .A(n20457), .ZN(n20167) );
  OAI22_X1 U23180 ( .A1(n20185), .A2(n20168), .B1(n20194), .B2(n20167), .ZN(
        n20169) );
  INV_X1 U23181 ( .A(n20169), .ZN(n20171) );
  AOI22_X1 U23182 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20188), .B1(
        n20187), .B2(n20460), .ZN(n20170) );
  OAI211_X1 U23183 ( .C1(n20338), .C2(n20208), .A(n20171), .B(n20170), .ZN(
        P2_U3108) );
  INV_X1 U23184 ( .A(n20465), .ZN(n20173) );
  INV_X1 U23185 ( .A(n20464), .ZN(n20172) );
  OAI22_X1 U23186 ( .A1(n20185), .A2(n20173), .B1(n20194), .B2(n20172), .ZN(
        n20174) );
  INV_X1 U23187 ( .A(n20174), .ZN(n20176) );
  AOI22_X1 U23188 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20188), .B1(
        n20216), .B2(n20466), .ZN(n20175) );
  OAI211_X1 U23189 ( .C1(n20379), .C2(n20177), .A(n20176), .B(n20175), .ZN(
        P2_U3109) );
  INV_X1 U23190 ( .A(n20471), .ZN(n20179) );
  INV_X1 U23191 ( .A(n20470), .ZN(n20178) );
  OAI22_X1 U23192 ( .A1(n20185), .A2(n20179), .B1(n20194), .B2(n20178), .ZN(
        n20180) );
  INV_X1 U23193 ( .A(n20180), .ZN(n20182) );
  AOI22_X1 U23194 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20188), .B1(
        n20187), .B2(n20473), .ZN(n20181) );
  OAI211_X1 U23195 ( .C1(n20344), .C2(n20208), .A(n20182), .B(n20181), .ZN(
        P2_U3110) );
  INV_X1 U23196 ( .A(n20478), .ZN(n20184) );
  INV_X1 U23197 ( .A(n20476), .ZN(n20183) );
  OAI22_X1 U23198 ( .A1(n20185), .A2(n20184), .B1(n20183), .B2(n20194), .ZN(
        n20186) );
  INV_X1 U23199 ( .A(n20186), .ZN(n20190) );
  AOI22_X1 U23200 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20188), .B1(
        n20187), .B2(n20482), .ZN(n20189) );
  OAI211_X1 U23201 ( .C1(n20351), .C2(n20208), .A(n20190), .B(n20189), .ZN(
        P2_U3111) );
  NAND2_X1 U23202 ( .A1(n20597), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20285) );
  INV_X1 U23203 ( .A(n20285), .ZN(n20287) );
  NAND2_X1 U23204 ( .A1(n20287), .A2(n20605), .ZN(n20230) );
  NOR2_X1 U23205 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20230), .ZN(
        n20215) );
  AOI22_X1 U23206 ( .A1(n20436), .A2(n20242), .B1(n20434), .B2(n20215), .ZN(
        n20201) );
  AOI21_X1 U23207 ( .B1(n20208), .B2(n20251), .A(n21109), .ZN(n20191) );
  NOR2_X1 U23208 ( .A1(n20191), .A2(n20578), .ZN(n20195) );
  OAI21_X1 U23209 ( .B1(n20197), .B2(n20491), .A(n21204), .ZN(n20192) );
  AOI21_X1 U23210 ( .B1(n20195), .B2(n20194), .A(n20192), .ZN(n20193) );
  OAI21_X1 U23211 ( .B1(n20215), .B2(n20193), .A(n20425), .ZN(n20218) );
  INV_X1 U23212 ( .A(n20194), .ZN(n20196) );
  OAI21_X1 U23213 ( .B1(n20196), .B2(n20215), .A(n20195), .ZN(n20199) );
  OAI21_X1 U23214 ( .B1(n20197), .B2(n20215), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20198) );
  AOI22_X1 U23215 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20218), .B1(
        n19938), .B2(n20217), .ZN(n20200) );
  OAI211_X1 U23216 ( .C1(n20364), .C2(n20208), .A(n20201), .B(n20200), .ZN(
        P2_U3112) );
  AOI22_X1 U23217 ( .A1(n20216), .A2(n20441), .B1(n20439), .B2(n20215), .ZN(
        n20203) );
  AOI22_X1 U23218 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20218), .B1(
        n13863), .B2(n20217), .ZN(n20202) );
  OAI211_X1 U23219 ( .C1(n20329), .C2(n20251), .A(n20203), .B(n20202), .ZN(
        P2_U3113) );
  AOI22_X1 U23220 ( .A1(n20447), .A2(n20242), .B1(n20444), .B2(n20215), .ZN(
        n20205) );
  AOI22_X1 U23221 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20218), .B1(
        n20445), .B2(n20217), .ZN(n20204) );
  OAI211_X1 U23222 ( .C1(n20370), .C2(n20208), .A(n20205), .B(n20204), .ZN(
        P2_U3114) );
  AOI22_X1 U23223 ( .A1(n20453), .A2(n20242), .B1(n20450), .B2(n20215), .ZN(
        n20207) );
  AOI22_X1 U23224 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20218), .B1(
        n20451), .B2(n20217), .ZN(n20206) );
  OAI211_X1 U23225 ( .C1(n20373), .C2(n20208), .A(n20207), .B(n20206), .ZN(
        P2_U3115) );
  AOI22_X1 U23226 ( .A1(n20216), .A2(n20460), .B1(n20457), .B2(n20215), .ZN(
        n20210) );
  AOI22_X1 U23227 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20218), .B1(
        n20458), .B2(n20217), .ZN(n20209) );
  OAI211_X1 U23228 ( .C1(n20338), .C2(n20251), .A(n20210), .B(n20209), .ZN(
        P2_U3116) );
  AOI22_X1 U23229 ( .A1(n20467), .A2(n20216), .B1(n20464), .B2(n20215), .ZN(
        n20212) );
  AOI22_X1 U23230 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20218), .B1(
        n20465), .B2(n20217), .ZN(n20211) );
  OAI211_X1 U23231 ( .C1(n20341), .C2(n20251), .A(n20212), .B(n20211), .ZN(
        P2_U3117) );
  AOI22_X1 U23232 ( .A1(n20216), .A2(n20473), .B1(n20470), .B2(n20215), .ZN(
        n20214) );
  AOI22_X1 U23233 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20218), .B1(
        n20471), .B2(n20217), .ZN(n20213) );
  OAI211_X1 U23234 ( .C1(n20344), .C2(n20251), .A(n20214), .B(n20213), .ZN(
        P2_U3118) );
  AOI22_X1 U23235 ( .A1(n20482), .A2(n20216), .B1(n20476), .B2(n20215), .ZN(
        n20220) );
  AOI22_X1 U23236 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20218), .B1(
        n20478), .B2(n20217), .ZN(n20219) );
  OAI211_X1 U23237 ( .C1(n20351), .C2(n20251), .A(n20220), .B(n20219), .ZN(
        P2_U3119) );
  NOR2_X1 U23238 ( .A1(n20221), .A2(n20285), .ZN(n20253) );
  AOI22_X1 U23239 ( .A1(n20436), .A2(n20281), .B1(n20434), .B2(n20253), .ZN(
        n20233) );
  NAND2_X1 U23240 ( .A1(n20582), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20428) );
  OR2_X1 U23241 ( .A1(n20428), .A2(n20222), .ZN(n20223) );
  INV_X1 U23242 ( .A(n20253), .ZN(n20224) );
  NAND2_X1 U23243 ( .A1(n10609), .A2(n20224), .ZN(n20228) );
  NOR2_X1 U23244 ( .A1(n20228), .A2(n20491), .ZN(n20225) );
  AOI21_X1 U23245 ( .B1(n20227), .B2(n20230), .A(n20225), .ZN(n20226) );
  OAI211_X1 U23246 ( .C1(n20253), .C2(n21204), .A(n20226), .B(n20425), .ZN(
        n20248) );
  INV_X1 U23247 ( .A(n20227), .ZN(n20231) );
  INV_X1 U23248 ( .A(n20228), .ZN(n20229) );
  AOI22_X1 U23249 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20248), .B1(
        n19938), .B2(n20247), .ZN(n20232) );
  OAI211_X1 U23250 ( .C1(n20364), .C2(n20251), .A(n20233), .B(n20232), .ZN(
        P2_U3120) );
  AOI22_X1 U23251 ( .A1(n20440), .A2(n20281), .B1(n20439), .B2(n20253), .ZN(
        n20235) );
  AOI22_X1 U23252 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20248), .B1(
        n13863), .B2(n20247), .ZN(n20234) );
  OAI211_X1 U23253 ( .C1(n20367), .C2(n20251), .A(n20235), .B(n20234), .ZN(
        P2_U3121) );
  AOI22_X1 U23254 ( .A1(n20446), .A2(n20242), .B1(n20444), .B2(n20253), .ZN(
        n20237) );
  AOI22_X1 U23255 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20248), .B1(
        n20445), .B2(n20247), .ZN(n20236) );
  OAI211_X1 U23256 ( .C1(n20332), .C2(n20272), .A(n20237), .B(n20236), .ZN(
        P2_U3122) );
  AOI22_X1 U23257 ( .A1(n20452), .A2(n20242), .B1(n20450), .B2(n20253), .ZN(
        n20239) );
  AOI22_X1 U23258 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20248), .B1(
        n20451), .B2(n20247), .ZN(n20238) );
  OAI211_X1 U23259 ( .C1(n20335), .C2(n20272), .A(n20239), .B(n20238), .ZN(
        P2_U3123) );
  AOI22_X1 U23260 ( .A1(n20459), .A2(n20281), .B1(n20457), .B2(n20253), .ZN(
        n20241) );
  AOI22_X1 U23261 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20248), .B1(
        n20458), .B2(n20247), .ZN(n20240) );
  OAI211_X1 U23262 ( .C1(n20376), .C2(n20251), .A(n20241), .B(n20240), .ZN(
        P2_U3124) );
  AOI22_X1 U23263 ( .A1(n20467), .A2(n20242), .B1(n20464), .B2(n20253), .ZN(
        n20244) );
  AOI22_X1 U23264 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20248), .B1(
        n20465), .B2(n20247), .ZN(n20243) );
  OAI211_X1 U23265 ( .C1(n20341), .C2(n20272), .A(n20244), .B(n20243), .ZN(
        P2_U3125) );
  AOI22_X1 U23266 ( .A1(n20472), .A2(n20281), .B1(n20470), .B2(n20253), .ZN(
        n20246) );
  AOI22_X1 U23267 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20248), .B1(
        n20471), .B2(n20247), .ZN(n20245) );
  OAI211_X1 U23268 ( .C1(n20382), .C2(n20251), .A(n20246), .B(n20245), .ZN(
        P2_U3126) );
  AOI22_X1 U23269 ( .A1(n20480), .A2(n20281), .B1(n20476), .B2(n20253), .ZN(
        n20250) );
  AOI22_X1 U23270 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20248), .B1(
        n20478), .B2(n20247), .ZN(n20249) );
  OAI211_X1 U23271 ( .C1(n20388), .C2(n20251), .A(n20250), .B(n20249), .ZN(
        P2_U3127) );
  NAND2_X1 U23272 ( .A1(n10610), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20256) );
  AOI21_X1 U23273 ( .B1(n20315), .B2(n20272), .A(n21109), .ZN(n20252) );
  NOR2_X1 U23274 ( .A1(n20253), .A2(n20252), .ZN(n20254) );
  NOR2_X1 U23275 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20254), .ZN(n20255) );
  NAND2_X1 U23276 ( .A1(n20256), .A2(n20255), .ZN(n20259) );
  NOR2_X1 U23277 ( .A1(n20257), .A2(n20285), .ZN(n20279) );
  INV_X1 U23278 ( .A(n20279), .ZN(n20258) );
  AOI21_X1 U23279 ( .B1(n20259), .B2(n20258), .A(n20395), .ZN(n20265) );
  INV_X1 U23280 ( .A(n10610), .ZN(n20260) );
  OAI21_X1 U23281 ( .B1(n20260), .B2(n20279), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20261) );
  AOI22_X1 U23282 ( .A1(n20280), .A2(n19938), .B1(n20434), .B2(n20279), .ZN(
        n20264) );
  AOI22_X1 U23283 ( .A1(n20297), .A2(n20436), .B1(n20281), .B2(n20435), .ZN(
        n20263) );
  OAI211_X1 U23284 ( .C1(n20265), .C2(n12188), .A(n20264), .B(n20263), .ZN(
        P2_U3128) );
  AOI22_X1 U23285 ( .A1(n20280), .A2(n13863), .B1(n20439), .B2(n20279), .ZN(
        n20267) );
  AOI22_X1 U23286 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20282), .B1(
        n20281), .B2(n20441), .ZN(n20266) );
  OAI211_X1 U23287 ( .C1(n20329), .C2(n20315), .A(n20267), .B(n20266), .ZN(
        P2_U3129) );
  AOI22_X1 U23288 ( .A1(n20280), .A2(n20445), .B1(n20444), .B2(n20279), .ZN(
        n20269) );
  AOI22_X1 U23289 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20282), .B1(
        n20297), .B2(n20447), .ZN(n20268) );
  OAI211_X1 U23290 ( .C1(n20370), .C2(n20272), .A(n20269), .B(n20268), .ZN(
        P2_U3130) );
  AOI22_X1 U23291 ( .A1(n20280), .A2(n20451), .B1(n20450), .B2(n20279), .ZN(
        n20271) );
  AOI22_X1 U23292 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20282), .B1(
        n20297), .B2(n20453), .ZN(n20270) );
  OAI211_X1 U23293 ( .C1(n20373), .C2(n20272), .A(n20271), .B(n20270), .ZN(
        P2_U3131) );
  AOI22_X1 U23294 ( .A1(n20280), .A2(n20458), .B1(n20457), .B2(n20279), .ZN(
        n20274) );
  AOI22_X1 U23295 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20282), .B1(
        n20281), .B2(n20460), .ZN(n20273) );
  OAI211_X1 U23296 ( .C1(n20338), .C2(n20315), .A(n20274), .B(n20273), .ZN(
        P2_U3132) );
  AOI22_X1 U23297 ( .A1(n20280), .A2(n20465), .B1(n20464), .B2(n20279), .ZN(
        n20276) );
  AOI22_X1 U23298 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20282), .B1(
        n20281), .B2(n20467), .ZN(n20275) );
  OAI211_X1 U23299 ( .C1(n20341), .C2(n20315), .A(n20276), .B(n20275), .ZN(
        P2_U3133) );
  AOI22_X1 U23300 ( .A1(n20280), .A2(n20471), .B1(n20470), .B2(n20279), .ZN(
        n20278) );
  AOI22_X1 U23301 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20282), .B1(
        n20281), .B2(n20473), .ZN(n20277) );
  OAI211_X1 U23302 ( .C1(n20344), .C2(n20315), .A(n20278), .B(n20277), .ZN(
        P2_U3134) );
  AOI22_X1 U23303 ( .A1(n20280), .A2(n20478), .B1(n20476), .B2(n20279), .ZN(
        n20284) );
  AOI22_X1 U23304 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20282), .B1(
        n20281), .B2(n20482), .ZN(n20283) );
  OAI211_X1 U23305 ( .C1(n20351), .C2(n20315), .A(n20284), .B(n20283), .ZN(
        P2_U3135) );
  INV_X1 U23306 ( .A(n20347), .ZN(n20318) );
  NOR2_X1 U23307 ( .A1(n20286), .A2(n20285), .ZN(n20310) );
  NOR3_X1 U23308 ( .A1(n10613), .A2(n20310), .A3(n20491), .ZN(n20290) );
  NAND2_X1 U23309 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20287), .ZN(
        n20293) );
  INV_X1 U23310 ( .A(n20293), .ZN(n20288) );
  AOI21_X1 U23311 ( .B1(n20288), .B2(n21204), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20289) );
  AOI22_X1 U23312 ( .A1(n20311), .A2(n19938), .B1(n20434), .B2(n20310), .ZN(
        n20296) );
  INV_X1 U23313 ( .A(n20290), .ZN(n20291) );
  OAI211_X1 U23314 ( .C1(n20310), .C2(n21204), .A(n20291), .B(n20425), .ZN(
        n20292) );
  AOI221_X1 U23315 ( .B1(n20293), .B2(n20576), .C1(n20293), .C2(n20428), .A(
        n20292), .ZN(n20294) );
  AOI22_X1 U23316 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20312), .B1(
        n20297), .B2(n20435), .ZN(n20295) );
  OAI211_X1 U23317 ( .C1(n20326), .C2(n20318), .A(n20296), .B(n20295), .ZN(
        P2_U3136) );
  AOI22_X1 U23318 ( .A1(n20311), .A2(n13863), .B1(n20439), .B2(n20310), .ZN(
        n20299) );
  AOI22_X1 U23319 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20312), .B1(
        n20297), .B2(n20441), .ZN(n20298) );
  OAI211_X1 U23320 ( .C1(n20329), .C2(n20318), .A(n20299), .B(n20298), .ZN(
        P2_U3137) );
  AOI22_X1 U23321 ( .A1(n20311), .A2(n20445), .B1(n20444), .B2(n20310), .ZN(
        n20301) );
  AOI22_X1 U23322 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20312), .B1(
        n20347), .B2(n20447), .ZN(n20300) );
  OAI211_X1 U23323 ( .C1(n20370), .C2(n20315), .A(n20301), .B(n20300), .ZN(
        P2_U3138) );
  AOI22_X1 U23324 ( .A1(n20311), .A2(n20451), .B1(n20450), .B2(n20310), .ZN(
        n20303) );
  AOI22_X1 U23325 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20312), .B1(
        n20347), .B2(n20453), .ZN(n20302) );
  OAI211_X1 U23326 ( .C1(n20373), .C2(n20315), .A(n20303), .B(n20302), .ZN(
        P2_U3139) );
  AOI22_X1 U23327 ( .A1(n20311), .A2(n20458), .B1(n20457), .B2(n20310), .ZN(
        n20305) );
  AOI22_X1 U23328 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20312), .B1(
        n20347), .B2(n20459), .ZN(n20304) );
  OAI211_X1 U23329 ( .C1(n20376), .C2(n20315), .A(n20305), .B(n20304), .ZN(
        P2_U3140) );
  AOI22_X1 U23330 ( .A1(n20311), .A2(n20465), .B1(n20464), .B2(n20310), .ZN(
        n20307) );
  AOI22_X1 U23331 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20312), .B1(
        n20347), .B2(n20466), .ZN(n20306) );
  OAI211_X1 U23332 ( .C1(n20379), .C2(n20315), .A(n20307), .B(n20306), .ZN(
        P2_U3141) );
  AOI22_X1 U23333 ( .A1(n20311), .A2(n20471), .B1(n20470), .B2(n20310), .ZN(
        n20309) );
  AOI22_X1 U23334 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20312), .B1(
        n20347), .B2(n20472), .ZN(n20308) );
  OAI211_X1 U23335 ( .C1(n20382), .C2(n20315), .A(n20309), .B(n20308), .ZN(
        P2_U3142) );
  AOI22_X1 U23336 ( .A1(n20311), .A2(n20478), .B1(n20476), .B2(n20310), .ZN(
        n20314) );
  AOI22_X1 U23337 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20312), .B1(
        n20347), .B2(n20480), .ZN(n20313) );
  OAI211_X1 U23338 ( .C1(n20388), .C2(n20315), .A(n20314), .B(n20313), .ZN(
        P2_U3143) );
  NOR2_X1 U23339 ( .A1(n10597), .A2(n20491), .ZN(n20320) );
  NAND3_X1 U23340 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20605), .ZN(n20358) );
  NOR2_X1 U23341 ( .A1(n20358), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20345) );
  INV_X1 U23342 ( .A(n20345), .ZN(n20319) );
  NAND3_X1 U23343 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20317), .A3(
        n21204), .ZN(n20316) );
  AOI22_X1 U23344 ( .A1(n20320), .A2(n20319), .B1(n20316), .B2(n20491), .ZN(
        n20346) );
  AOI22_X1 U23345 ( .A1(n20346), .A2(n19938), .B1(n20434), .B2(n20345), .ZN(
        n20325) );
  AND2_X1 U23346 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20317), .ZN(
        n20323) );
  AOI21_X1 U23347 ( .B1(n20387), .B2(n20318), .A(n21109), .ZN(n20322) );
  OAI21_X1 U23348 ( .B1(n20320), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20319), 
        .ZN(n20321) );
  OAI211_X1 U23349 ( .C1(n20323), .C2(n20322), .A(n20425), .B(n20321), .ZN(
        n20348) );
  AOI22_X1 U23350 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20435), .ZN(n20324) );
  OAI211_X1 U23351 ( .C1(n20326), .C2(n20387), .A(n20325), .B(n20324), .ZN(
        P2_U3144) );
  AOI22_X1 U23352 ( .A1(n20346), .A2(n13863), .B1(n20439), .B2(n20345), .ZN(
        n20328) );
  AOI22_X1 U23353 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20441), .ZN(n20327) );
  OAI211_X1 U23354 ( .C1(n20329), .C2(n20387), .A(n20328), .B(n20327), .ZN(
        P2_U3145) );
  AOI22_X1 U23355 ( .A1(n20346), .A2(n20445), .B1(n20444), .B2(n20345), .ZN(
        n20331) );
  AOI22_X1 U23356 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20446), .ZN(n20330) );
  OAI211_X1 U23357 ( .C1(n20332), .C2(n20387), .A(n20331), .B(n20330), .ZN(
        P2_U3146) );
  AOI22_X1 U23358 ( .A1(n20346), .A2(n20451), .B1(n20450), .B2(n20345), .ZN(
        n20334) );
  AOI22_X1 U23359 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20452), .ZN(n20333) );
  OAI211_X1 U23360 ( .C1(n20335), .C2(n20387), .A(n20334), .B(n20333), .ZN(
        P2_U3147) );
  AOI22_X1 U23361 ( .A1(n20346), .A2(n20458), .B1(n20457), .B2(n20345), .ZN(
        n20337) );
  AOI22_X1 U23362 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20460), .ZN(n20336) );
  OAI211_X1 U23363 ( .C1(n20338), .C2(n20387), .A(n20337), .B(n20336), .ZN(
        P2_U3148) );
  AOI22_X1 U23364 ( .A1(n20346), .A2(n20465), .B1(n20464), .B2(n20345), .ZN(
        n20340) );
  AOI22_X1 U23365 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20467), .ZN(n20339) );
  OAI211_X1 U23366 ( .C1(n20341), .C2(n20387), .A(n20340), .B(n20339), .ZN(
        P2_U3149) );
  AOI22_X1 U23367 ( .A1(n20346), .A2(n20471), .B1(n20470), .B2(n20345), .ZN(
        n20343) );
  AOI22_X1 U23368 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20473), .ZN(n20342) );
  OAI211_X1 U23369 ( .C1(n20344), .C2(n20387), .A(n20343), .B(n20342), .ZN(
        P2_U3150) );
  AOI22_X1 U23370 ( .A1(n20346), .A2(n20478), .B1(n20476), .B2(n20345), .ZN(
        n20350) );
  AOI22_X1 U23371 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20482), .ZN(n20349) );
  OAI211_X1 U23372 ( .C1(n20351), .C2(n20387), .A(n20350), .B(n20349), .ZN(
        P2_U3151) );
  NOR2_X1 U23373 ( .A1(n20615), .A2(n20358), .ZN(n20394) );
  NOR3_X1 U23374 ( .A1(n20352), .A2(n20394), .A3(n20491), .ZN(n20355) );
  INV_X1 U23375 ( .A(n20358), .ZN(n20353) );
  AOI21_X1 U23376 ( .B1(n21204), .B2(n20353), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20354) );
  NOR2_X1 U23377 ( .A1(n20355), .A2(n20354), .ZN(n20383) );
  AOI22_X1 U23378 ( .A1(n20383), .A2(n19938), .B1(n20434), .B2(n20394), .ZN(
        n20363) );
  INV_X1 U23379 ( .A(n20355), .ZN(n20356) );
  OAI211_X1 U23380 ( .C1(n20394), .C2(n21204), .A(n20356), .B(n20425), .ZN(
        n20357) );
  AOI221_X1 U23381 ( .B1(n20358), .B2(n20360), .C1(n20358), .C2(n20428), .A(
        n20357), .ZN(n20359) );
  AOI22_X1 U23382 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20384), .B1(
        n20418), .B2(n20436), .ZN(n20362) );
  OAI211_X1 U23383 ( .C1(n20364), .C2(n20387), .A(n20363), .B(n20362), .ZN(
        P2_U3152) );
  AOI22_X1 U23384 ( .A1(n20383), .A2(n13863), .B1(n20439), .B2(n20394), .ZN(
        n20366) );
  AOI22_X1 U23385 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20384), .B1(
        n20418), .B2(n20440), .ZN(n20365) );
  OAI211_X1 U23386 ( .C1(n20367), .C2(n20387), .A(n20366), .B(n20365), .ZN(
        P2_U3153) );
  AOI22_X1 U23387 ( .A1(n20383), .A2(n20445), .B1(n20444), .B2(n20394), .ZN(
        n20369) );
  AOI22_X1 U23388 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20384), .B1(
        n20418), .B2(n20447), .ZN(n20368) );
  OAI211_X1 U23389 ( .C1(n20370), .C2(n20387), .A(n20369), .B(n20368), .ZN(
        P2_U3154) );
  AOI22_X1 U23390 ( .A1(n20383), .A2(n20451), .B1(n20450), .B2(n20394), .ZN(
        n20372) );
  AOI22_X1 U23391 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20384), .B1(
        n20418), .B2(n20453), .ZN(n20371) );
  OAI211_X1 U23392 ( .C1(n20373), .C2(n20387), .A(n20372), .B(n20371), .ZN(
        P2_U3155) );
  AOI22_X1 U23393 ( .A1(n20383), .A2(n20458), .B1(n20457), .B2(n20394), .ZN(
        n20375) );
  AOI22_X1 U23394 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20384), .B1(
        n20418), .B2(n20459), .ZN(n20374) );
  OAI211_X1 U23395 ( .C1(n20376), .C2(n20387), .A(n20375), .B(n20374), .ZN(
        P2_U3156) );
  AOI22_X1 U23396 ( .A1(n20383), .A2(n20465), .B1(n20464), .B2(n20394), .ZN(
        n20378) );
  AOI22_X1 U23397 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20384), .B1(
        n20418), .B2(n20466), .ZN(n20377) );
  OAI211_X1 U23398 ( .C1(n20379), .C2(n20387), .A(n20378), .B(n20377), .ZN(
        P2_U3157) );
  AOI22_X1 U23399 ( .A1(n20383), .A2(n20471), .B1(n20470), .B2(n20394), .ZN(
        n20381) );
  AOI22_X1 U23400 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20384), .B1(
        n20418), .B2(n20472), .ZN(n20380) );
  OAI211_X1 U23401 ( .C1(n20382), .C2(n20387), .A(n20381), .B(n20380), .ZN(
        P2_U3158) );
  AOI22_X1 U23402 ( .A1(n20383), .A2(n20478), .B1(n20476), .B2(n20394), .ZN(
        n20386) );
  AOI22_X1 U23403 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20384), .B1(
        n20418), .B2(n20480), .ZN(n20385) );
  OAI211_X1 U23404 ( .C1(n20388), .C2(n20387), .A(n20386), .B(n20385), .ZN(
        P2_U3159) );
  INV_X1 U23405 ( .A(n20418), .ZN(n20389) );
  NAND2_X1 U23406 ( .A1(n20389), .A2(n20585), .ZN(n20392) );
  INV_X1 U23407 ( .A(n20580), .ZN(n20391) );
  OAI21_X1 U23408 ( .B1(n20392), .B2(n20483), .A(n20391), .ZN(n20397) );
  NAND2_X1 U23409 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20393), .ZN(
        n20430) );
  NOR2_X1 U23410 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20430), .ZN(
        n20417) );
  NOR2_X1 U23411 ( .A1(n20417), .A2(n20394), .ZN(n20399) );
  AOI211_X1 U23412 ( .C1(n10665), .C2(n21204), .A(n20417), .B(n20585), .ZN(
        n20396) );
  AOI22_X1 U23413 ( .A1(n20436), .A2(n20483), .B1(n20434), .B2(n20417), .ZN(
        n20402) );
  INV_X1 U23414 ( .A(n20397), .ZN(n20400) );
  OAI21_X1 U23415 ( .B1(n10665), .B2(n20417), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20398) );
  AOI22_X1 U23416 ( .A1(n19938), .A2(n20419), .B1(n20418), .B2(n20435), .ZN(
        n20401) );
  OAI211_X1 U23417 ( .C1(n20422), .C2(n20403), .A(n20402), .B(n20401), .ZN(
        P2_U3160) );
  AOI22_X1 U23418 ( .A1(n20440), .A2(n20483), .B1(n20439), .B2(n20417), .ZN(
        n20405) );
  AOI22_X1 U23419 ( .A1(n13863), .A2(n20419), .B1(n20418), .B2(n20441), .ZN(
        n20404) );
  OAI211_X1 U23420 ( .C1(n20422), .C2(n12452), .A(n20405), .B(n20404), .ZN(
        P2_U3161) );
  AOI22_X1 U23421 ( .A1(n20446), .A2(n20418), .B1(n20444), .B2(n20417), .ZN(
        n20407) );
  AOI22_X1 U23422 ( .A1(n20445), .A2(n20419), .B1(n20483), .B2(n20447), .ZN(
        n20406) );
  OAI211_X1 U23423 ( .C1(n20422), .C2(n12229), .A(n20407), .B(n20406), .ZN(
        P2_U3162) );
  AOI22_X1 U23424 ( .A1(n20452), .A2(n20418), .B1(n20450), .B2(n20417), .ZN(
        n20409) );
  AOI22_X1 U23425 ( .A1(n20451), .A2(n20419), .B1(n20483), .B2(n20453), .ZN(
        n20408) );
  OAI211_X1 U23426 ( .C1(n20422), .C2(n20410), .A(n20409), .B(n20408), .ZN(
        P2_U3163) );
  AOI22_X1 U23427 ( .A1(n20460), .A2(n20418), .B1(n20457), .B2(n20417), .ZN(
        n20412) );
  AOI22_X1 U23428 ( .A1(n20458), .A2(n20419), .B1(n20483), .B2(n20459), .ZN(
        n20411) );
  OAI211_X1 U23429 ( .C1(n20422), .C2(n12530), .A(n20412), .B(n20411), .ZN(
        P2_U3164) );
  AOI22_X1 U23430 ( .A1(n20467), .A2(n20418), .B1(n20464), .B2(n20417), .ZN(
        n20414) );
  AOI22_X1 U23431 ( .A1(n20465), .A2(n20419), .B1(n20483), .B2(n20466), .ZN(
        n20413) );
  OAI211_X1 U23432 ( .C1(n20422), .C2(n12559), .A(n20414), .B(n20413), .ZN(
        P2_U3165) );
  AOI22_X1 U23433 ( .A1(n20473), .A2(n20418), .B1(n20470), .B2(n20417), .ZN(
        n20416) );
  AOI22_X1 U23434 ( .A1(n20471), .A2(n20419), .B1(n20483), .B2(n20472), .ZN(
        n20415) );
  OAI211_X1 U23435 ( .C1(n20422), .C2(n12576), .A(n20416), .B(n20415), .ZN(
        P2_U3166) );
  AOI22_X1 U23436 ( .A1(n20482), .A2(n20418), .B1(n20476), .B2(n20417), .ZN(
        n20421) );
  AOI22_X1 U23437 ( .A1(n20478), .A2(n20419), .B1(n20483), .B2(n20480), .ZN(
        n20420) );
  OAI211_X1 U23438 ( .C1(n20422), .C2(n12256), .A(n20421), .B(n20420), .ZN(
        P2_U3167) );
  INV_X1 U23439 ( .A(n20423), .ZN(n20477) );
  NOR3_X1 U23440 ( .A1(n20424), .A2(n20477), .A3(n20491), .ZN(n20433) );
  INV_X1 U23441 ( .A(n20433), .ZN(n20426) );
  OAI211_X1 U23442 ( .C1(n20477), .C2(n21204), .A(n20426), .B(n20425), .ZN(
        n20427) );
  INV_X1 U23443 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n21219) );
  INV_X1 U23444 ( .A(n20430), .ZN(n20431) );
  AOI21_X1 U23445 ( .B1(n21204), .B2(n20431), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20432) );
  NOR2_X1 U23446 ( .A1(n20433), .A2(n20432), .ZN(n20479) );
  AOI22_X1 U23447 ( .A1(n20479), .A2(n19938), .B1(n20477), .B2(n20434), .ZN(
        n20438) );
  AOI22_X1 U23448 ( .A1(n20481), .A2(n20436), .B1(n20483), .B2(n20435), .ZN(
        n20437) );
  OAI211_X1 U23449 ( .C1(n20487), .C2(n21219), .A(n20438), .B(n20437), .ZN(
        P2_U3168) );
  AOI22_X1 U23450 ( .A1(n20479), .A2(n13863), .B1(n20477), .B2(n20439), .ZN(
        n20443) );
  AOI22_X1 U23451 ( .A1(n20483), .A2(n20441), .B1(n20481), .B2(n20440), .ZN(
        n20442) );
  OAI211_X1 U23452 ( .C1(n20487), .C2(n12314), .A(n20443), .B(n20442), .ZN(
        P2_U3169) );
  AOI22_X1 U23453 ( .A1(n20479), .A2(n20445), .B1(n20477), .B2(n20444), .ZN(
        n20449) );
  AOI22_X1 U23454 ( .A1(n20481), .A2(n20447), .B1(n20483), .B2(n20446), .ZN(
        n20448) );
  OAI211_X1 U23455 ( .C1(n20487), .C2(n12479), .A(n20449), .B(n20448), .ZN(
        P2_U3170) );
  INV_X1 U23456 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20456) );
  AOI22_X1 U23457 ( .A1(n20479), .A2(n20451), .B1(n20477), .B2(n20450), .ZN(
        n20455) );
  AOI22_X1 U23458 ( .A1(n20481), .A2(n20453), .B1(n20483), .B2(n20452), .ZN(
        n20454) );
  OAI211_X1 U23459 ( .C1(n20487), .C2(n20456), .A(n20455), .B(n20454), .ZN(
        P2_U3171) );
  INV_X1 U23460 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n20463) );
  AOI22_X1 U23461 ( .A1(n20479), .A2(n20458), .B1(n20477), .B2(n20457), .ZN(
        n20462) );
  AOI22_X1 U23462 ( .A1(n20483), .A2(n20460), .B1(n20481), .B2(n20459), .ZN(
        n20461) );
  OAI211_X1 U23463 ( .C1(n20487), .C2(n20463), .A(n20462), .B(n20461), .ZN(
        P2_U3172) );
  AOI22_X1 U23464 ( .A1(n20479), .A2(n20465), .B1(n20477), .B2(n20464), .ZN(
        n20469) );
  AOI22_X1 U23465 ( .A1(n20483), .A2(n20467), .B1(n20481), .B2(n20466), .ZN(
        n20468) );
  OAI211_X1 U23466 ( .C1(n20487), .C2(n10601), .A(n20469), .B(n20468), .ZN(
        P2_U3173) );
  AOI22_X1 U23467 ( .A1(n20479), .A2(n20471), .B1(n20477), .B2(n20470), .ZN(
        n20475) );
  AOI22_X1 U23468 ( .A1(n20483), .A2(n20473), .B1(n20481), .B2(n20472), .ZN(
        n20474) );
  OAI211_X1 U23469 ( .C1(n20487), .C2(n10658), .A(n20475), .B(n20474), .ZN(
        P2_U3174) );
  AOI22_X1 U23470 ( .A1(n20479), .A2(n20478), .B1(n20477), .B2(n20476), .ZN(
        n20485) );
  AOI22_X1 U23471 ( .A1(n20483), .A2(n20482), .B1(n20481), .B2(n20480), .ZN(
        n20484) );
  OAI211_X1 U23472 ( .C1(n20487), .C2(n20486), .A(n20485), .B(n20484), .ZN(
        P2_U3175) );
  AOI21_X1 U23473 ( .B1(n20509), .B2(n20490), .A(n20488), .ZN(n20496) );
  AOI211_X1 U23474 ( .C1(n20491), .C2(n20509), .A(n20490), .B(n20489), .ZN(
        n20492) );
  INV_X1 U23475 ( .A(n20492), .ZN(n20493) );
  OAI22_X1 U23476 ( .A1(n20496), .A2(n20495), .B1(n20494), .B2(n20493), .ZN(
        P2_U3177) );
  AND2_X1 U23477 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20497), .ZN(
        P2_U3179) );
  AND2_X1 U23478 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20497), .ZN(
        P2_U3180) );
  AND2_X1 U23479 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20497), .ZN(
        P2_U3181) );
  AND2_X1 U23480 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20497), .ZN(
        P2_U3182) );
  AND2_X1 U23481 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20497), .ZN(
        P2_U3183) );
  AND2_X1 U23482 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20497), .ZN(
        P2_U3184) );
  AND2_X1 U23483 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20497), .ZN(
        P2_U3185) );
  AND2_X1 U23484 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20497), .ZN(
        P2_U3186) );
  AND2_X1 U23485 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20497), .ZN(
        P2_U3187) );
  AND2_X1 U23486 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20497), .ZN(
        P2_U3188) );
  AND2_X1 U23487 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20497), .ZN(
        P2_U3189) );
  AND2_X1 U23488 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20497), .ZN(
        P2_U3190) );
  AND2_X1 U23489 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20497), .ZN(
        P2_U3191) );
  AND2_X1 U23490 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20497), .ZN(
        P2_U3192) );
  AND2_X1 U23491 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20497), .ZN(
        P2_U3193) );
  AND2_X1 U23492 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20497), .ZN(
        P2_U3194) );
  AND2_X1 U23493 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20497), .ZN(
        P2_U3195) );
  AND2_X1 U23494 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20497), .ZN(
        P2_U3196) );
  AND2_X1 U23495 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20497), .ZN(
        P2_U3197) );
  AND2_X1 U23496 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20497), .ZN(
        P2_U3198) );
  AND2_X1 U23497 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20497), .ZN(
        P2_U3199) );
  AND2_X1 U23498 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20497), .ZN(
        P2_U3200) );
  AND2_X1 U23499 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20497), .ZN(P2_U3201) );
  AND2_X1 U23500 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20497), .ZN(P2_U3202) );
  AND2_X1 U23501 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20497), .ZN(P2_U3203) );
  AND2_X1 U23502 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20497), .ZN(P2_U3204) );
  AND2_X1 U23503 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20497), .ZN(P2_U3205) );
  AND2_X1 U23504 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20497), .ZN(P2_U3206) );
  AND2_X1 U23505 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20497), .ZN(P2_U3207) );
  AND2_X1 U23506 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20497), .ZN(P2_U3208) );
  NAND2_X1 U23507 ( .A1(n20509), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20511) );
  NAND3_X1 U23508 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20511), .ZN(n20500) );
  AOI211_X1 U23509 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20971), .A(
        n20498), .B(n20627), .ZN(n20499) );
  INV_X1 U23510 ( .A(NA), .ZN(n20976) );
  NOR2_X1 U23511 ( .A1(n20976), .A2(n20504), .ZN(n20516) );
  AOI211_X1 U23512 ( .C1(n20517), .C2(n20500), .A(n20499), .B(n20516), .ZN(
        n20501) );
  INV_X1 U23513 ( .A(n20501), .ZN(P2_U3209) );
  INV_X1 U23514 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20502) );
  AOI21_X1 U23515 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20971), .A(n20517), 
        .ZN(n20508) );
  NOR2_X1 U23516 ( .A1(n20502), .A2(n20508), .ZN(n20505) );
  AOI21_X1 U23517 ( .B1(n20505), .B2(n20504), .A(n20503), .ZN(n20506) );
  OAI211_X1 U23518 ( .C1(n20971), .C2(n20507), .A(n20506), .B(n20511), .ZN(
        P2_U3210) );
  AOI21_X1 U23519 ( .B1(n20510), .B2(n20509), .A(n20508), .ZN(n20515) );
  OAI22_X1 U23520 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20512), .B1(NA), 
        .B2(n20511), .ZN(n20513) );
  OAI211_X1 U23521 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20513), .ZN(n20514) );
  OAI21_X1 U23522 ( .B1(n20516), .B2(n20515), .A(n20514), .ZN(P2_U3211) );
  OAI222_X1 U23523 ( .A1(n20559), .A2(n20519), .B1(n20518), .B2(n20627), .C1(
        n14081), .C2(n20556), .ZN(P2_U3212) );
  OAI222_X1 U23524 ( .A1(n20559), .A2(n12673), .B1(n20520), .B2(n20627), .C1(
        n20519), .C2(n20556), .ZN(P2_U3213) );
  OAI222_X1 U23525 ( .A1(n20559), .A2(n14003), .B1(n20521), .B2(n20627), .C1(
        n12673), .C2(n20556), .ZN(P2_U3214) );
  OAI222_X1 U23526 ( .A1(n20559), .A2(n14024), .B1(n20522), .B2(n20627), .C1(
        n14003), .C2(n20556), .ZN(P2_U3215) );
  OAI222_X1 U23527 ( .A1(n20559), .A2(n10861), .B1(n21125), .B2(n20627), .C1(
        n14024), .C2(n20556), .ZN(P2_U3216) );
  OAI222_X1 U23528 ( .A1(n20559), .A2(n10865), .B1(n20523), .B2(n20627), .C1(
        n10861), .C2(n20556), .ZN(P2_U3217) );
  OAI222_X1 U23529 ( .A1(n20559), .A2(n12689), .B1(n20524), .B2(n20627), .C1(
        n10865), .C2(n20556), .ZN(P2_U3218) );
  OAI222_X1 U23530 ( .A1(n20559), .A2(n10846), .B1(n20525), .B2(n20627), .C1(
        n12689), .C2(n20556), .ZN(P2_U3219) );
  OAI222_X1 U23531 ( .A1(n20559), .A2(n15879), .B1(n20526), .B2(n20627), .C1(
        n10846), .C2(n20556), .ZN(P2_U3220) );
  OAI222_X1 U23532 ( .A1(n20559), .A2(n12702), .B1(n20527), .B2(n20627), .C1(
        n15879), .C2(n20556), .ZN(P2_U3221) );
  OAI222_X1 U23533 ( .A1(n20559), .A2(n12705), .B1(n20528), .B2(n20627), .C1(
        n12702), .C2(n20556), .ZN(P2_U3222) );
  OAI222_X1 U23534 ( .A1(n20559), .A2(n12710), .B1(n20529), .B2(n20627), .C1(
        n12705), .C2(n20556), .ZN(P2_U3223) );
  OAI222_X1 U23535 ( .A1(n20559), .A2(n15842), .B1(n20530), .B2(n20627), .C1(
        n12710), .C2(n20556), .ZN(P2_U3224) );
  OAI222_X1 U23536 ( .A1(n20559), .A2(n10889), .B1(n20531), .B2(n20627), .C1(
        n15842), .C2(n20556), .ZN(P2_U3225) );
  OAI222_X1 U23537 ( .A1(n20559), .A2(n12720), .B1(n20532), .B2(n20627), .C1(
        n10889), .C2(n20556), .ZN(P2_U3226) );
  OAI222_X1 U23538 ( .A1(n20559), .A2(n20534), .B1(n20533), .B2(n20627), .C1(
        n12720), .C2(n20556), .ZN(P2_U3227) );
  OAI222_X1 U23539 ( .A1(n20559), .A2(n15792), .B1(n20535), .B2(n20627), .C1(
        n20534), .C2(n20556), .ZN(P2_U3228) );
  OAI222_X1 U23540 ( .A1(n20559), .A2(n20537), .B1(n20536), .B2(n20627), .C1(
        n15792), .C2(n20556), .ZN(P2_U3229) );
  OAI222_X1 U23541 ( .A1(n20559), .A2(n15768), .B1(n20538), .B2(n20627), .C1(
        n20537), .C2(n20556), .ZN(P2_U3230) );
  OAI222_X1 U23542 ( .A1(n20559), .A2(n20540), .B1(n20539), .B2(n20627), .C1(
        n15768), .C2(n20556), .ZN(P2_U3231) );
  OAI222_X1 U23543 ( .A1(n20559), .A2(n15733), .B1(n21202), .B2(n20627), .C1(
        n20540), .C2(n20556), .ZN(P2_U3232) );
  OAI222_X1 U23544 ( .A1(n20559), .A2(n20542), .B1(n20541), .B2(n20627), .C1(
        n15733), .C2(n20556), .ZN(P2_U3233) );
  INV_X1 U23545 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20544) );
  OAI222_X1 U23546 ( .A1(n20559), .A2(n20544), .B1(n20543), .B2(n20627), .C1(
        n20542), .C2(n20556), .ZN(P2_U3234) );
  OAI222_X1 U23547 ( .A1(n20559), .A2(n20546), .B1(n20545), .B2(n20627), .C1(
        n20544), .C2(n20556), .ZN(P2_U3235) );
  OAI222_X1 U23548 ( .A1(n20559), .A2(n20548), .B1(n20547), .B2(n20627), .C1(
        n20546), .C2(n20556), .ZN(P2_U3236) );
  OAI222_X1 U23549 ( .A1(n20559), .A2(n20551), .B1(n20549), .B2(n20627), .C1(
        n20548), .C2(n20556), .ZN(P2_U3237) );
  OAI222_X1 U23550 ( .A1(n20556), .A2(n20551), .B1(n20550), .B2(n20627), .C1(
        n20552), .C2(n20559), .ZN(P2_U3238) );
  OAI222_X1 U23551 ( .A1(n20559), .A2(n20554), .B1(n20553), .B2(n20627), .C1(
        n20552), .C2(n20556), .ZN(P2_U3239) );
  INV_X1 U23552 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20557) );
  OAI222_X1 U23553 ( .A1(n20559), .A2(n20557), .B1(n20555), .B2(n20627), .C1(
        n20554), .C2(n20556), .ZN(P2_U3240) );
  OAI222_X1 U23554 ( .A1(n20559), .A2(n14463), .B1(n20558), .B2(n20627), .C1(
        n20557), .C2(n20556), .ZN(P2_U3241) );
  OAI22_X1 U23555 ( .A1(n20628), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20627), .ZN(n20560) );
  INV_X1 U23556 ( .A(n20560), .ZN(P2_U3585) );
  MUX2_X1 U23557 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20628), .Z(P2_U3586) );
  OAI22_X1 U23558 ( .A1(n20628), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20627), .ZN(n20561) );
  INV_X1 U23559 ( .A(n20561), .ZN(P2_U3587) );
  OAI22_X1 U23560 ( .A1(n20628), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20627), .ZN(n20562) );
  INV_X1 U23561 ( .A(n20562), .ZN(P2_U3588) );
  OAI21_X1 U23562 ( .B1(n20566), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20564), 
        .ZN(n20563) );
  INV_X1 U23563 ( .A(n20563), .ZN(P2_U3591) );
  OAI21_X1 U23564 ( .B1(n20566), .B2(n20565), .A(n20564), .ZN(P2_U3592) );
  OAI22_X1 U23565 ( .A1(n20570), .A2(n20569), .B1(n20568), .B2(n20567), .ZN(
        n20572) );
  OAI22_X1 U23566 ( .A1(n20573), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20572), .B2(n20571), .ZN(n20574) );
  INV_X1 U23567 ( .A(n20574), .ZN(P2_U3596) );
  INV_X1 U23568 ( .A(n20575), .ZN(n20586) );
  INV_X1 U23569 ( .A(n20576), .ZN(n20577) );
  AND2_X1 U23570 ( .A1(n20585), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20601) );
  NAND2_X1 U23571 ( .A1(n20577), .A2(n20601), .ZN(n20591) );
  OR2_X1 U23572 ( .A1(n20599), .A2(n20578), .ZN(n20581) );
  NOR2_X1 U23573 ( .A1(n20580), .A2(n20579), .ZN(n20598) );
  AND2_X1 U23574 ( .A1(n20581), .A2(n20598), .ZN(n20589) );
  NAND2_X1 U23575 ( .A1(n20591), .A2(n20589), .ZN(n20583) );
  AOI222_X1 U23576 ( .A1(n20586), .A2(n20585), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20584), .C1(n20583), .C2(n20582), .ZN(n20587) );
  AOI22_X1 U23577 ( .A1(n20616), .A2(n20588), .B1(n20587), .B2(n20613), .ZN(
        P2_U3602) );
  INV_X1 U23578 ( .A(n20589), .ZN(n20594) );
  NOR2_X1 U23579 ( .A1(n20590), .A2(n21204), .ZN(n20593) );
  INV_X1 U23580 ( .A(n20591), .ZN(n20592) );
  AOI211_X1 U23581 ( .C1(n20595), .C2(n20594), .A(n20593), .B(n20592), .ZN(
        n20596) );
  AOI22_X1 U23582 ( .A1(n20616), .A2(n20597), .B1(n20596), .B2(n20613), .ZN(
        P2_U3603) );
  INV_X1 U23583 ( .A(n20598), .ZN(n20600) );
  MUX2_X1 U23584 ( .A(n20601), .B(n20600), .S(n20599), .Z(n20602) );
  AOI21_X1 U23585 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20603), .A(n20602), 
        .ZN(n20604) );
  AOI22_X1 U23586 ( .A1(n20616), .A2(n20605), .B1(n20604), .B2(n20613), .ZN(
        P2_U3604) );
  INV_X1 U23587 ( .A(n20606), .ZN(n20612) );
  INV_X1 U23588 ( .A(n20607), .ZN(n20608) );
  OAI22_X1 U23589 ( .A1(n20609), .A2(n20608), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21204), .ZN(n20610) );
  AOI21_X1 U23590 ( .B1(n20612), .B2(n20611), .A(n20610), .ZN(n20614) );
  AOI22_X1 U23591 ( .A1(n20616), .A2(n20615), .B1(n20614), .B2(n20613), .ZN(
        P2_U3605) );
  INV_X1 U23592 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20617) );
  AOI22_X1 U23593 ( .A1(n20627), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20617), 
        .B2(n20628), .ZN(P2_U3608) );
  INV_X1 U23594 ( .A(n20618), .ZN(n20624) );
  AOI22_X1 U23595 ( .A1(n20622), .A2(n20621), .B1(n20620), .B2(n20619), .ZN(
        n20623) );
  NAND2_X1 U23596 ( .A1(n20624), .A2(n20623), .ZN(n20626) );
  MUX2_X1 U23597 ( .A(P2_MORE_REG_SCAN_IN), .B(n20626), .S(n20625), .Z(
        P2_U3609) );
  OAI22_X1 U23598 ( .A1(n20628), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20627), .ZN(n20629) );
  INV_X1 U23599 ( .A(n20629), .ZN(P2_U3611) );
  NOR2_X1 U23600 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20630), .ZN(n20980) );
  NOR2_X1 U23601 ( .A1(n20980), .A2(n20972), .ZN(n20638) );
  INV_X1 U23602 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20631) );
  AOI21_X1 U23603 ( .B1(n20638), .B2(n20631), .A(n21048), .ZN(P1_U2802) );
  NAND2_X1 U23604 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20632), .ZN(n20636) );
  OAI21_X1 U23605 ( .B1(n20634), .B2(n20633), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20635) );
  OAI21_X1 U23606 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20636), .A(n20635), 
        .ZN(P1_U2803) );
  NOR2_X1 U23607 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20639) );
  OAI21_X1 U23608 ( .B1(n20639), .B2(P1_D_C_N_REG_SCAN_IN), .A(n9598), .ZN(
        n20637) );
  OAI21_X1 U23609 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n9598), .A(n20637), 
        .ZN(P1_U2804) );
  NOR2_X1 U23610 ( .A1(n21048), .A2(n20638), .ZN(n21038) );
  OAI21_X1 U23611 ( .B1(BS16), .B2(n20639), .A(n21038), .ZN(n21036) );
  OAI21_X1 U23612 ( .B1(n21038), .B2(n20640), .A(n21036), .ZN(P1_U2805) );
  INV_X1 U23613 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20641) );
  OAI21_X1 U23614 ( .B1(n20642), .B2(n20641), .A(n21068), .ZN(P1_U2806) );
  NOR4_X1 U23615 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20646) );
  NOR4_X1 U23616 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20645) );
  NOR4_X1 U23617 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20644) );
  NOR4_X1 U23618 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20643) );
  NAND4_X1 U23619 ( .A1(n20646), .A2(n20645), .A3(n20644), .A4(n20643), .ZN(
        n20652) );
  NOR4_X1 U23620 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20650) );
  AOI211_X1 U23621 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_4__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20649) );
  NOR4_X1 U23622 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20648) );
  NOR4_X1 U23623 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20647) );
  NAND4_X1 U23624 ( .A1(n20650), .A2(n20649), .A3(n20648), .A4(n20647), .ZN(
        n20651) );
  NOR2_X1 U23625 ( .A1(n20652), .A2(n20651), .ZN(n21043) );
  INV_X1 U23626 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20654) );
  NOR3_X1 U23627 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20655) );
  OAI21_X1 U23628 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20655), .A(n21043), .ZN(
        n20653) );
  OAI21_X1 U23629 ( .B1(n21043), .B2(n20654), .A(n20653), .ZN(P1_U2807) );
  INV_X1 U23630 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21037) );
  AOI21_X1 U23631 ( .B1(n21039), .B2(n21037), .A(n20655), .ZN(n20657) );
  INV_X1 U23632 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20656) );
  INV_X1 U23633 ( .A(n21043), .ZN(n21045) );
  AOI22_X1 U23634 ( .A1(n21043), .A2(n20657), .B1(n20656), .B2(n21045), .ZN(
        P1_U2808) );
  NAND2_X1 U23635 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20658) );
  OAI21_X1 U23636 ( .B1(n20658), .B2(n20682), .A(n20683), .ZN(n20680) );
  NOR3_X1 U23637 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20688), .A3(n20658), .ZN(
        n20659) );
  AOI211_X1 U23638 ( .C1(n20705), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20660), .B(n20659), .ZN(n20664) );
  INV_X1 U23639 ( .A(n20661), .ZN(n20662) );
  AOI22_X1 U23640 ( .A1(n20684), .A2(P1_EBX_REG_7__SCAN_IN), .B1(n20662), .B2(
        n20687), .ZN(n20663) );
  OAI211_X1 U23641 ( .C1(n20666), .C2(n20665), .A(n20664), .B(n20663), .ZN(
        n20667) );
  AOI21_X1 U23642 ( .B1(n20676), .B2(n20668), .A(n20667), .ZN(n20669) );
  OAI21_X1 U23643 ( .B1(n20670), .B2(n20680), .A(n20669), .ZN(P1_U2833) );
  INV_X1 U23644 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20681) );
  AOI22_X1 U23645 ( .A1(n20671), .A2(n20700), .B1(n20684), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n20679) );
  NOR2_X1 U23646 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20688), .ZN(n20672) );
  AOI22_X1 U23647 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20705), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20672), .ZN(n20673) );
  OAI211_X1 U23648 ( .C1(n20674), .C2(n20703), .A(n20673), .B(n20702), .ZN(
        n20675) );
  AOI21_X1 U23649 ( .B1(n20677), .B2(n20676), .A(n20675), .ZN(n20678) );
  OAI211_X1 U23650 ( .C1(n20681), .C2(n20680), .A(n20679), .B(n20678), .ZN(
        P1_U2834) );
  INV_X1 U23651 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20989) );
  NAND2_X1 U23652 ( .A1(n20683), .A2(n20682), .ZN(n20711) );
  AOI22_X1 U23653 ( .A1(n20684), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n20700), .B2(
        n20713), .ZN(n20694) );
  NAND2_X1 U23654 ( .A1(n20714), .A2(n20709), .ZN(n20692) );
  INV_X1 U23655 ( .A(n20685), .ZN(n20686) );
  AOI22_X1 U23656 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20705), .B1(
        n20687), .B2(n20686), .ZN(n20691) );
  OAI21_X1 U23657 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20688), .A(n20702), .ZN(
        n20689) );
  INV_X1 U23658 ( .A(n20689), .ZN(n20690) );
  AND3_X1 U23659 ( .A1(n20692), .A2(n20691), .A3(n20690), .ZN(n20693) );
  OAI211_X1 U23660 ( .C1(n20989), .C2(n20711), .A(n20694), .B(n20693), .ZN(
        P1_U2835) );
  AOI21_X1 U23661 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n20695), .A(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20712) );
  INV_X1 U23662 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20720) );
  XNOR2_X1 U23663 ( .A(n20697), .B(n9973), .ZN(n20797) );
  AOI22_X1 U23664 ( .A1(n20700), .A2(n20797), .B1(n20699), .B2(n20698), .ZN(
        n20701) );
  OAI211_X1 U23665 ( .C1(n20703), .C2(n20795), .A(n20702), .B(n20701), .ZN(
        n20704) );
  AOI21_X1 U23666 ( .B1(n20705), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20704), .ZN(n20706) );
  OAI21_X1 U23667 ( .B1(n20720), .B2(n20707), .A(n20706), .ZN(n20708) );
  AOI21_X1 U23668 ( .B1(n20790), .B2(n20709), .A(n20708), .ZN(n20710) );
  OAI21_X1 U23669 ( .B1(n20712), .B2(n20711), .A(n20710), .ZN(P1_U2836) );
  INV_X1 U23670 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20716) );
  AOI22_X1 U23671 ( .A1(n20714), .A2(n20718), .B1(n20717), .B2(n20713), .ZN(
        n20715) );
  OAI21_X1 U23672 ( .B1(n20721), .B2(n20716), .A(n20715), .ZN(P1_U2867) );
  AOI22_X1 U23673 ( .A1(n20790), .A2(n20718), .B1(n20717), .B2(n20797), .ZN(
        n20719) );
  OAI21_X1 U23674 ( .B1(n20721), .B2(n20720), .A(n20719), .ZN(P1_U2868) );
  AOI22_X1 U23675 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20722) );
  OAI21_X1 U23676 ( .B1(n13226), .B2(n20748), .A(n20722), .ZN(P1_U2921) );
  AOI22_X1 U23677 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20723) );
  OAI21_X1 U23678 ( .B1(n14798), .B2(n20748), .A(n20723), .ZN(P1_U2922) );
  INV_X1 U23679 ( .A(P1_LWORD_REG_13__SCAN_IN), .ZN(n21128) );
  AOI22_X1 U23680 ( .A1(P1_EAX_REG_13__SCAN_IN), .A2(n20724), .B1(n20737), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20725) );
  OAI21_X1 U23681 ( .B1(n21128), .B2(n20726), .A(n20725), .ZN(P1_U2923) );
  AOI22_X1 U23682 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20727) );
  OAI21_X1 U23683 ( .B1(n14803), .B2(n20748), .A(n20727), .ZN(P1_U2924) );
  AOI22_X1 U23684 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20728) );
  OAI21_X1 U23685 ( .B1(n14149), .B2(n20748), .A(n20728), .ZN(P1_U2925) );
  AOI22_X1 U23686 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20729) );
  OAI21_X1 U23687 ( .B1(n14107), .B2(n20748), .A(n20729), .ZN(P1_U2926) );
  INV_X1 U23688 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20731) );
  AOI22_X1 U23689 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20730) );
  OAI21_X1 U23690 ( .B1(n20731), .B2(n20748), .A(n20730), .ZN(P1_U2927) );
  INV_X1 U23691 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20733) );
  AOI22_X1 U23692 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20732) );
  OAI21_X1 U23693 ( .B1(n20733), .B2(n20748), .A(n20732), .ZN(P1_U2928) );
  AOI22_X1 U23694 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20734) );
  OAI21_X1 U23695 ( .B1(n11386), .B2(n20748), .A(n20734), .ZN(P1_U2929) );
  AOI22_X1 U23696 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20735) );
  OAI21_X1 U23697 ( .B1(n11370), .B2(n20748), .A(n20735), .ZN(P1_U2930) );
  AOI22_X1 U23698 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20737), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20736), .ZN(n20738) );
  OAI21_X1 U23699 ( .B1(n13529), .B2(n20748), .A(n20738), .ZN(P1_U2931) );
  AOI22_X1 U23700 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20739) );
  OAI21_X1 U23701 ( .B1(n20740), .B2(n20748), .A(n20739), .ZN(P1_U2932) );
  AOI22_X1 U23702 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20741) );
  OAI21_X1 U23703 ( .B1(n20742), .B2(n20748), .A(n20741), .ZN(P1_U2933) );
  AOI22_X1 U23704 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20743) );
  OAI21_X1 U23705 ( .B1(n20744), .B2(n20748), .A(n20743), .ZN(P1_U2934) );
  AOI22_X1 U23706 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20745) );
  OAI21_X1 U23707 ( .B1(n20746), .B2(n20748), .A(n20745), .ZN(P1_U2935) );
  AOI22_X1 U23708 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20736), .B1(n20737), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20747) );
  OAI21_X1 U23709 ( .B1(n20749), .B2(n20748), .A(n20747), .ZN(P1_U2936) );
  AOI22_X1 U23710 ( .A1(n20778), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20783), .ZN(n20751) );
  NAND2_X1 U23711 ( .A1(n9720), .A2(n20750), .ZN(n20770) );
  NAND2_X1 U23712 ( .A1(n20751), .A2(n20770), .ZN(P1_U2945) );
  AOI22_X1 U23713 ( .A1(n20778), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20753) );
  NAND2_X1 U23714 ( .A1(n9720), .A2(n20752), .ZN(n20772) );
  NAND2_X1 U23715 ( .A1(n20753), .A2(n20772), .ZN(P1_U2946) );
  AOI22_X1 U23716 ( .A1(n20778), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20756) );
  INV_X1 U23717 ( .A(n20754), .ZN(n20755) );
  NAND2_X1 U23718 ( .A1(n9720), .A2(n20755), .ZN(n20774) );
  NAND2_X1 U23719 ( .A1(n20756), .A2(n20774), .ZN(P1_U2947) );
  AOI22_X1 U23720 ( .A1(n20778), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20759) );
  INV_X1 U23721 ( .A(n20757), .ZN(n20758) );
  NAND2_X1 U23722 ( .A1(n9720), .A2(n20758), .ZN(n20776) );
  NAND2_X1 U23723 ( .A1(n20759), .A2(n20776), .ZN(P1_U2948) );
  AOI22_X1 U23724 ( .A1(n20778), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20762) );
  INV_X1 U23725 ( .A(n20760), .ZN(n20761) );
  NAND2_X1 U23726 ( .A1(n9720), .A2(n20761), .ZN(n20779) );
  NAND2_X1 U23727 ( .A1(n20762), .A2(n20779), .ZN(P1_U2949) );
  AOI22_X1 U23728 ( .A1(n20778), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20765) );
  INV_X1 U23729 ( .A(n20763), .ZN(n20764) );
  NAND2_X1 U23730 ( .A1(n9720), .A2(n20764), .ZN(n20781) );
  NAND2_X1 U23731 ( .A1(n20765), .A2(n20781), .ZN(P1_U2950) );
  AOI22_X1 U23732 ( .A1(n20778), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20783), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20769) );
  INV_X1 U23733 ( .A(n20766), .ZN(n20767) );
  NAND2_X1 U23734 ( .A1(n9720), .A2(n20767), .ZN(n20784) );
  NAND2_X1 U23735 ( .A1(n20769), .A2(n20784), .ZN(P1_U2951) );
  AOI22_X1 U23736 ( .A1(n20778), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20783), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20771) );
  NAND2_X1 U23737 ( .A1(n20771), .A2(n20770), .ZN(P1_U2960) );
  AOI22_X1 U23738 ( .A1(n20778), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20783), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20773) );
  NAND2_X1 U23739 ( .A1(n20773), .A2(n20772), .ZN(P1_U2961) );
  AOI22_X1 U23740 ( .A1(n20778), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20783), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20775) );
  NAND2_X1 U23741 ( .A1(n20775), .A2(n20774), .ZN(P1_U2962) );
  AOI22_X1 U23742 ( .A1(n20778), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20783), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20777) );
  NAND2_X1 U23743 ( .A1(n20777), .A2(n20776), .ZN(P1_U2963) );
  AOI22_X1 U23744 ( .A1(n20778), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20783), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20780) );
  NAND2_X1 U23745 ( .A1(n20780), .A2(n20779), .ZN(P1_U2964) );
  AOI22_X1 U23746 ( .A1(n20778), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20783), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20782) );
  NAND2_X1 U23747 ( .A1(n20782), .A2(n20781), .ZN(P1_U2965) );
  AOI22_X1 U23748 ( .A1(n20778), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20783), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20785) );
  NAND2_X1 U23749 ( .A1(n20785), .A2(n20784), .ZN(P1_U2966) );
  AOI22_X1 U23750 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20794) );
  OAI21_X1 U23751 ( .B1(n20788), .B2(n20787), .A(n20786), .ZN(n20789) );
  INV_X1 U23752 ( .A(n20789), .ZN(n20799) );
  AOI22_X1 U23753 ( .A1(n20799), .A2(n20792), .B1(n20791), .B2(n20790), .ZN(
        n20793) );
  OAI211_X1 U23754 ( .C1(n16695), .C2(n20795), .A(n20794), .B(n20793), .ZN(
        P1_U2995) );
  OAI21_X1 U23755 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20796), .ZN(n20802) );
  AOI22_X1 U23756 ( .A1(n21060), .A2(P1_REIP_REG_4__SCAN_IN), .B1(n20849), 
        .B2(n20797), .ZN(n20801) );
  INV_X1 U23757 ( .A(n20798), .ZN(n20805) );
  AOI22_X1 U23758 ( .A1(n20799), .A2(n20806), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20805), .ZN(n20800) );
  OAI211_X1 U23759 ( .C1(n20810), .C2(n20802), .A(n20801), .B(n20800), .ZN(
        P1_U3027) );
  AOI22_X1 U23760 ( .A1(n21060), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n20849), 
        .B2(n20803), .ZN(n20809) );
  INV_X1 U23761 ( .A(n20804), .ZN(n20807) );
  AOI22_X1 U23762 ( .A1(n20807), .A2(n20806), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20805), .ZN(n20808) );
  OAI211_X1 U23763 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20810), .A(
        n20809), .B(n20808), .ZN(P1_U3028) );
  NAND2_X1 U23764 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20811), .ZN(
        n20823) );
  OAI21_X1 U23765 ( .B1(n20852), .B2(n20813), .A(n20812), .ZN(n20819) );
  OAI22_X1 U23766 ( .A1(n20836), .A2(n20815), .B1(n20814), .B2(n16817), .ZN(
        n20818) );
  NOR2_X1 U23767 ( .A1(n20816), .A2(n20844), .ZN(n20817) );
  AOI211_X1 U23768 ( .C1(n20827), .C2(n20819), .A(n20818), .B(n20817), .ZN(
        n20820) );
  OAI221_X1 U23769 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20823), .C1(
        n20822), .C2(n20821), .A(n20820), .ZN(P1_U3029) );
  NOR2_X1 U23770 ( .A1(n20824), .A2(n20844), .ZN(n20833) );
  NOR3_X1 U23771 ( .A1(n20826), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n20825), .ZN(n20831) );
  NAND2_X1 U23772 ( .A1(n20827), .A2(n20852), .ZN(n20842) );
  AOI21_X1 U23773 ( .B1(n20829), .B2(n20842), .A(n20828), .ZN(n20830) );
  AOI211_X1 U23774 ( .C1(n20833), .C2(n20832), .A(n20831), .B(n20830), .ZN(
        n20835) );
  NAND2_X1 U23775 ( .A1(n21060), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20834) );
  OAI211_X1 U23776 ( .C1(n20837), .C2(n20836), .A(n20835), .B(n20834), .ZN(
        P1_U3030) );
  NOR2_X1 U23777 ( .A1(n20839), .A2(n20838), .ZN(n20851) );
  INV_X1 U23778 ( .A(n20840), .ZN(n20845) );
  INV_X1 U23779 ( .A(n20841), .ZN(n20843) );
  OAI211_X1 U23780 ( .C1(n20845), .C2(n20844), .A(n20843), .B(n20842), .ZN(
        n20846) );
  AOI211_X1 U23781 ( .C1(n20849), .C2(n20848), .A(n20847), .B(n20846), .ZN(
        n20850) );
  OAI21_X1 U23782 ( .B1(n20852), .B2(n20851), .A(n20850), .ZN(P1_U3031) );
  NOR2_X1 U23783 ( .A1(n20854), .A2(n20853), .ZN(P1_U3032) );
  NOR2_X1 U23784 ( .A1(n20887), .A2(n20893), .ZN(n20857) );
  INV_X1 U23785 ( .A(n20855), .ZN(n20894) );
  AOI21_X1 U23786 ( .B1(n20857), .B2(n20856), .A(n20894), .ZN(n20871) );
  INV_X1 U23787 ( .A(n20871), .ZN(n20862) );
  AND2_X1 U23788 ( .A1(n20859), .A2(n20858), .ZN(n20870) );
  NAND2_X1 U23789 ( .A1(n20864), .A2(n20863), .ZN(n20867) );
  INV_X1 U23790 ( .A(n20867), .ZN(n20886) );
  AOI22_X1 U23791 ( .A1(n20888), .A2(n20903), .B1(n20886), .B2(n20902), .ZN(
        n20873) );
  INV_X1 U23792 ( .A(n20865), .ZN(n20866) );
  AOI21_X1 U23793 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20867), .A(n20866), 
        .ZN(n20868) );
  OAI211_X1 U23794 ( .C1(n20871), .C2(n20870), .A(n20869), .B(n20868), .ZN(
        n20889) );
  AOI22_X1 U23795 ( .A1(n20889), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n20887), .B2(n20912), .ZN(n20872) );
  OAI211_X1 U23796 ( .C1(n20892), .C2(n20915), .A(n20873), .B(n20872), .ZN(
        P1_U3113) );
  AOI22_X1 U23797 ( .A1(n20888), .A2(n20917), .B1(n20886), .B2(n20916), .ZN(
        n20875) );
  AOI22_X1 U23798 ( .A1(n20889), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n20887), .B2(n20918), .ZN(n20874) );
  OAI211_X1 U23799 ( .C1(n20892), .C2(n20921), .A(n20875), .B(n20874), .ZN(
        P1_U3114) );
  AOI22_X1 U23800 ( .A1(n20888), .A2(n20923), .B1(n20886), .B2(n20922), .ZN(
        n20877) );
  AOI22_X1 U23801 ( .A1(n20889), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n20887), .B2(n20924), .ZN(n20876) );
  OAI211_X1 U23802 ( .C1(n20892), .C2(n20927), .A(n20877), .B(n20876), .ZN(
        P1_U3115) );
  AOI22_X1 U23803 ( .A1(n20887), .A2(n20930), .B1(n20928), .B2(n20886), .ZN(
        n20879) );
  AOI22_X1 U23804 ( .A1(n20889), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n20888), .B2(n20929), .ZN(n20878) );
  OAI211_X1 U23805 ( .C1(n20892), .C2(n20933), .A(n20879), .B(n20878), .ZN(
        P1_U3116) );
  AOI22_X1 U23806 ( .A1(n20887), .A2(n20936), .B1(n20934), .B2(n20886), .ZN(
        n20881) );
  AOI22_X1 U23807 ( .A1(n20889), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n20888), .B2(n20935), .ZN(n20880) );
  OAI211_X1 U23808 ( .C1(n20892), .C2(n20939), .A(n20881), .B(n20880), .ZN(
        P1_U3117) );
  AOI22_X1 U23809 ( .A1(n20887), .A2(n20942), .B1(n20940), .B2(n20886), .ZN(
        n20883) );
  AOI22_X1 U23810 ( .A1(n20889), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n20888), .B2(n20941), .ZN(n20882) );
  OAI211_X1 U23811 ( .C1(n20892), .C2(n20945), .A(n20883), .B(n20882), .ZN(
        P1_U3118) );
  AOI22_X1 U23812 ( .A1(n20887), .A2(n20948), .B1(n20946), .B2(n20886), .ZN(
        n20885) );
  AOI22_X1 U23813 ( .A1(n20889), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n20888), .B2(n20947), .ZN(n20884) );
  OAI211_X1 U23814 ( .C1(n20892), .C2(n20951), .A(n20885), .B(n20884), .ZN(
        P1_U3119) );
  AOI22_X1 U23815 ( .A1(n20887), .A2(n20955), .B1(n20952), .B2(n20886), .ZN(
        n20891) );
  AOI22_X1 U23816 ( .A1(n20889), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n20888), .B2(n20954), .ZN(n20890) );
  OAI211_X1 U23817 ( .C1(n20892), .C2(n20960), .A(n20891), .B(n20890), .ZN(
        P1_U3120) );
  NOR2_X1 U23818 ( .A1(n10195), .A2(n20893), .ZN(n20895) );
  AOI21_X1 U23819 ( .B1(n20895), .B2(n20911), .A(n20894), .ZN(n20910) );
  INV_X1 U23820 ( .A(n20910), .ZN(n20900) );
  AND2_X1 U23821 ( .A1(n20897), .A2(n20896), .ZN(n20909) );
  NOR2_X1 U23822 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20901), .ZN(
        n20953) );
  AOI22_X1 U23823 ( .A1(n10195), .A2(n20903), .B1(n20953), .B2(n20902), .ZN(
        n20914) );
  OAI21_X1 U23824 ( .B1(n20905), .B2(n20953), .A(n20904), .ZN(n20906) );
  AOI21_X1 U23825 ( .B1(n20907), .B2(P1_STATE2_REG_2__SCAN_IN), .A(n20906), 
        .ZN(n20908) );
  OAI21_X1 U23826 ( .B1(n20910), .B2(n20909), .A(n20908), .ZN(n20957) );
  AOI22_X1 U23827 ( .A1(n20957), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n20956), .B2(n20912), .ZN(n20913) );
  OAI211_X1 U23828 ( .C1(n20961), .C2(n20915), .A(n20914), .B(n20913), .ZN(
        P1_U3129) );
  AOI22_X1 U23829 ( .A1(n10195), .A2(n20917), .B1(n20953), .B2(n20916), .ZN(
        n20920) );
  AOI22_X1 U23830 ( .A1(n20957), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n20956), .B2(n20918), .ZN(n20919) );
  OAI211_X1 U23831 ( .C1(n20961), .C2(n20921), .A(n20920), .B(n20919), .ZN(
        P1_U3130) );
  AOI22_X1 U23832 ( .A1(n10195), .A2(n20923), .B1(n20953), .B2(n20922), .ZN(
        n20926) );
  AOI22_X1 U23833 ( .A1(n20957), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n20956), .B2(n20924), .ZN(n20925) );
  OAI211_X1 U23834 ( .C1(n20961), .C2(n20927), .A(n20926), .B(n20925), .ZN(
        P1_U3131) );
  AOI22_X1 U23835 ( .A1(n10195), .A2(n20929), .B1(n20953), .B2(n20928), .ZN(
        n20932) );
  AOI22_X1 U23836 ( .A1(n20957), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n20956), .B2(n20930), .ZN(n20931) );
  OAI211_X1 U23837 ( .C1(n20961), .C2(n20933), .A(n20932), .B(n20931), .ZN(
        P1_U3132) );
  AOI22_X1 U23838 ( .A1(n10195), .A2(n20935), .B1(n20953), .B2(n20934), .ZN(
        n20938) );
  AOI22_X1 U23839 ( .A1(n20957), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n20956), .B2(n20936), .ZN(n20937) );
  OAI211_X1 U23840 ( .C1(n20961), .C2(n20939), .A(n20938), .B(n20937), .ZN(
        P1_U3133) );
  AOI22_X1 U23841 ( .A1(n10195), .A2(n20941), .B1(n20953), .B2(n20940), .ZN(
        n20944) );
  AOI22_X1 U23842 ( .A1(n20957), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n20956), .B2(n20942), .ZN(n20943) );
  OAI211_X1 U23843 ( .C1(n20961), .C2(n20945), .A(n20944), .B(n20943), .ZN(
        P1_U3134) );
  AOI22_X1 U23844 ( .A1(n10195), .A2(n20947), .B1(n20953), .B2(n20946), .ZN(
        n20950) );
  AOI22_X1 U23845 ( .A1(n20957), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n20956), .B2(n20948), .ZN(n20949) );
  OAI211_X1 U23846 ( .C1(n20961), .C2(n20951), .A(n20950), .B(n20949), .ZN(
        P1_U3135) );
  AOI22_X1 U23847 ( .A1(n10195), .A2(n20954), .B1(n20953), .B2(n20952), .ZN(
        n20959) );
  AOI22_X1 U23848 ( .A1(n20957), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n20956), .B2(n20955), .ZN(n20958) );
  OAI211_X1 U23849 ( .C1(n20961), .C2(n20960), .A(n20959), .B(n20958), .ZN(
        P1_U3136) );
  NOR2_X1 U23850 ( .A1(n20963), .A2(n20962), .ZN(n20965) );
  OAI21_X1 U23851 ( .B1(n20965), .B2(n13658), .A(n20964), .ZN(P1_U3163) );
  AND2_X1 U23852 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20966), .ZN(
        P1_U3164) );
  AND2_X1 U23853 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20966), .ZN(
        P1_U3165) );
  AND2_X1 U23854 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20966), .ZN(
        P1_U3166) );
  AND2_X1 U23855 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20966), .ZN(
        P1_U3167) );
  AND2_X1 U23856 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20966), .ZN(
        P1_U3168) );
  AND2_X1 U23857 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20966), .ZN(
        P1_U3169) );
  AND2_X1 U23858 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20966), .ZN(
        P1_U3170) );
  AND2_X1 U23859 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20966), .ZN(
        P1_U3171) );
  AND2_X1 U23860 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20966), .ZN(
        P1_U3172) );
  AND2_X1 U23861 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20966), .ZN(
        P1_U3173) );
  AND2_X1 U23862 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20966), .ZN(
        P1_U3174) );
  AND2_X1 U23863 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20966), .ZN(
        P1_U3175) );
  AND2_X1 U23864 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20966), .ZN(
        P1_U3176) );
  AND2_X1 U23865 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20966), .ZN(
        P1_U3177) );
  AND2_X1 U23866 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20966), .ZN(
        P1_U3178) );
  AND2_X1 U23867 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20966), .ZN(
        P1_U3179) );
  AND2_X1 U23868 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20966), .ZN(
        P1_U3180) );
  AND2_X1 U23869 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20966), .ZN(
        P1_U3181) );
  AND2_X1 U23870 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20966), .ZN(
        P1_U3182) );
  AND2_X1 U23871 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20966), .ZN(
        P1_U3183) );
  AND2_X1 U23872 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20966), .ZN(
        P1_U3184) );
  AND2_X1 U23873 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20966), .ZN(
        P1_U3185) );
  AND2_X1 U23874 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20966), .ZN(P1_U3186) );
  AND2_X1 U23875 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20966), .ZN(P1_U3187) );
  AND2_X1 U23876 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20966), .ZN(P1_U3188) );
  AND2_X1 U23877 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20966), .ZN(P1_U3189) );
  AND2_X1 U23878 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20966), .ZN(P1_U3190) );
  INV_X1 U23879 ( .A(P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n21153) );
  NOR2_X1 U23880 ( .A1(n21038), .A2(n21153), .ZN(P1_U3191) );
  AND2_X1 U23881 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20966), .ZN(P1_U3192) );
  AND2_X1 U23882 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20966), .ZN(P1_U3193) );
  AOI21_X1 U23883 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20973), .A(n20972), 
        .ZN(n20977) );
  NOR2_X1 U23884 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20967) );
  OAI22_X1 U23885 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20976), .B1(n20967), 
        .B2(n20971), .ZN(n20968) );
  NOR2_X1 U23886 ( .A1(n20969), .A2(n20968), .ZN(n20970) );
  OAI22_X1 U23887 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20977), .B1(n21048), 
        .B2(n20970), .ZN(P1_U3194) );
  AOI211_X1 U23888 ( .C1(n20982), .C2(P1_REQUESTPENDING_REG_SCAN_IN), .A(
        n20972), .B(n20971), .ZN(n20975) );
  INV_X1 U23889 ( .A(n20975), .ZN(n20981) );
  OAI211_X1 U23890 ( .C1(n20975), .C2(n20974), .A(P1_STATE_REG_1__SCAN_IN), 
        .B(n20973), .ZN(n20979) );
  OAI21_X1 U23891 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20976), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n20978) );
  OAI222_X1 U23892 ( .A1(n20981), .A2(n20980), .B1(NA), .B2(n20979), .C1(
        n20978), .C2(n20977), .ZN(P1_U3196) );
  NOR2_X2 U23893 ( .A1(n9598), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21023) );
  NOR2_X2 U23894 ( .A1(n20982), .A2(n9598), .ZN(n21027) );
  AOI222_X1 U23895 ( .A1(n21023), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n21027), .ZN(n20983) );
  INV_X1 U23896 ( .A(n20983), .ZN(P1_U3197) );
  AOI222_X1 U23897 ( .A1(n21027), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n21023), .ZN(n20984) );
  INV_X1 U23898 ( .A(n20984), .ZN(P1_U3198) );
  INV_X1 U23899 ( .A(n21027), .ZN(n21025) );
  INV_X1 U23900 ( .A(n21023), .ZN(n21029) );
  OAI222_X1 U23901 ( .A1(n21025), .A2(n20986), .B1(n20985), .B2(n21048), .C1(
        n20987), .C2(n21029), .ZN(P1_U3199) );
  INV_X1 U23902 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20988) );
  OAI222_X1 U23903 ( .A1(n21029), .A2(n20989), .B1(n20988), .B2(n21048), .C1(
        n20987), .C2(n21025), .ZN(P1_U3200) );
  AOI222_X1 U23904 ( .A1(n21027), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n21023), .ZN(n20990) );
  INV_X1 U23905 ( .A(n20990), .ZN(P1_U3201) );
  AOI222_X1 U23906 ( .A1(n21027), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n21023), .ZN(n20991) );
  INV_X1 U23907 ( .A(n20991), .ZN(P1_U3202) );
  AOI222_X1 U23908 ( .A1(n21027), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21023), .ZN(n20992) );
  INV_X1 U23909 ( .A(n20992), .ZN(P1_U3203) );
  AOI222_X1 U23910 ( .A1(n21023), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21027), .ZN(n20993) );
  INV_X1 U23911 ( .A(n20993), .ZN(P1_U3204) );
  AOI222_X1 U23912 ( .A1(n21027), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21023), .ZN(n20994) );
  INV_X1 U23913 ( .A(n20994), .ZN(P1_U3205) );
  AOI22_X1 U23914 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n21023), .ZN(n20995) );
  OAI21_X1 U23915 ( .B1(n20996), .B2(n21025), .A(n20995), .ZN(P1_U3206) );
  AOI22_X1 U23916 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n21027), .ZN(n20997) );
  OAI21_X1 U23917 ( .B1(n20998), .B2(n21029), .A(n20997), .ZN(P1_U3207) );
  AOI222_X1 U23918 ( .A1(n21023), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21027), .ZN(n20999) );
  INV_X1 U23919 ( .A(n20999), .ZN(P1_U3208) );
  AOI222_X1 U23920 ( .A1(n21027), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21023), .ZN(n21000) );
  INV_X1 U23921 ( .A(n21000), .ZN(P1_U3209) );
  AOI22_X1 U23922 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n21023), .ZN(n21001) );
  OAI21_X1 U23923 ( .B1(n21002), .B2(n21025), .A(n21001), .ZN(P1_U3210) );
  AOI22_X1 U23924 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21023), .ZN(n21003) );
  OAI21_X1 U23925 ( .B1(n16599), .B2(n21025), .A(n21003), .ZN(P1_U3211) );
  AOI22_X1 U23926 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21027), .ZN(n21004) );
  OAI21_X1 U23927 ( .B1(n21005), .B2(n21029), .A(n21004), .ZN(P1_U3212) );
  AOI222_X1 U23928 ( .A1(n21023), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n21027), .ZN(n21006) );
  INV_X1 U23929 ( .A(n21006), .ZN(P1_U3213) );
  INV_X1 U23930 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n21089) );
  OAI222_X1 U23931 ( .A1(n21025), .A2(n21007), .B1(n21089), .B2(n21048), .C1(
        n21009), .C2(n21029), .ZN(P1_U3214) );
  AOI22_X1 U23932 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21023), .ZN(n21008) );
  OAI21_X1 U23933 ( .B1(n21009), .B2(n21025), .A(n21008), .ZN(P1_U3215) );
  AOI22_X1 U23934 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21027), .ZN(n21010) );
  OAI21_X1 U23935 ( .B1(n21011), .B2(n21029), .A(n21010), .ZN(P1_U3216) );
  AOI222_X1 U23936 ( .A1(n21027), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n21023), .ZN(n21012) );
  INV_X1 U23937 ( .A(n21012), .ZN(P1_U3217) );
  AOI22_X1 U23938 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21023), .ZN(n21013) );
  OAI21_X1 U23939 ( .B1(n21014), .B2(n21025), .A(n21013), .ZN(P1_U3218) );
  AOI22_X1 U23940 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21027), .ZN(n21015) );
  OAI21_X1 U23941 ( .B1(n21017), .B2(n21029), .A(n21015), .ZN(P1_U3219) );
  AOI22_X1 U23942 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(n21023), .ZN(n21016) );
  OAI21_X1 U23943 ( .B1(n21017), .B2(n21025), .A(n21016), .ZN(P1_U3220) );
  AOI22_X1 U23944 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(n21027), .ZN(n21018) );
  OAI21_X1 U23945 ( .B1(n21020), .B2(n21029), .A(n21018), .ZN(P1_U3221) );
  INV_X1 U23946 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21078) );
  OAI222_X1 U23947 ( .A1(n21025), .A2(n21020), .B1(n21078), .B2(n21048), .C1(
        n21019), .C2(n21029), .ZN(P1_U3222) );
  AOI222_X1 U23948 ( .A1(n21027), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n21023), .ZN(n21021) );
  INV_X1 U23949 ( .A(n21021), .ZN(P1_U3223) );
  AOI222_X1 U23950 ( .A1(n21027), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n9598), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21023), .ZN(n21022) );
  INV_X1 U23951 ( .A(n21022), .ZN(P1_U3224) );
  AOI22_X1 U23952 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n21023), .ZN(n21024) );
  OAI21_X1 U23953 ( .B1(n21026), .B2(n21025), .A(n21024), .ZN(P1_U3225) );
  AOI22_X1 U23954 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(n9598), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n21027), .ZN(n21028) );
  OAI21_X1 U23955 ( .B1(n21030), .B2(n21029), .A(n21028), .ZN(P1_U3226) );
  OAI22_X1 U23956 ( .A1(n9598), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21048), .ZN(n21031) );
  INV_X1 U23957 ( .A(n21031), .ZN(P1_U3458) );
  OAI22_X1 U23958 ( .A1(n9598), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21048), .ZN(n21032) );
  INV_X1 U23959 ( .A(n21032), .ZN(P1_U3459) );
  OAI22_X1 U23960 ( .A1(n9598), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21048), .ZN(n21033) );
  INV_X1 U23961 ( .A(n21033), .ZN(P1_U3460) );
  OAI22_X1 U23962 ( .A1(n9598), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21048), .ZN(n21034) );
  INV_X1 U23963 ( .A(n21034), .ZN(P1_U3461) );
  OAI21_X1 U23964 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21038), .A(n21036), 
        .ZN(n21035) );
  INV_X1 U23965 ( .A(n21035), .ZN(P1_U3464) );
  OAI21_X1 U23966 ( .B1(n21038), .B2(n21037), .A(n21036), .ZN(P1_U3465) );
  AOI21_X1 U23967 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21040) );
  AOI22_X1 U23968 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21040), .B2(n21039), .ZN(n21042) );
  INV_X1 U23969 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21041) );
  AOI22_X1 U23970 ( .A1(n21043), .A2(n21042), .B1(n21041), .B2(n21045), .ZN(
        P1_U3481) );
  INV_X1 U23971 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21046) );
  NOR2_X1 U23972 ( .A1(n21045), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21044) );
  AOI22_X1 U23973 ( .A1(n21046), .A2(n21045), .B1(n13096), .B2(n21044), .ZN(
        P1_U3482) );
  AOI22_X1 U23974 ( .A1(n21048), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21047), 
        .B2(n9598), .ZN(P1_U3483) );
  AOI211_X1 U23975 ( .C1(n20736), .C2(n21051), .A(n21050), .B(n21049), .ZN(
        n21058) );
  NAND3_X1 U23976 ( .A1(n21053), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n21052), 
        .ZN(n21055) );
  AOI21_X1 U23977 ( .B1(n21055), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n21054), 
        .ZN(n21057) );
  NAND2_X1 U23978 ( .A1(n21058), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21056) );
  OAI21_X1 U23979 ( .B1(n21058), .B2(n21057), .A(n21056), .ZN(P1_U3485) );
  MUX2_X1 U23980 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n9598), .Z(P1_U3486) );
  INV_X1 U23981 ( .A(n21059), .ZN(n21069) );
  AOI22_X1 U23982 ( .A1(n21061), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n21060), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n21067) );
  OAI22_X1 U23983 ( .A1(n21064), .A2(n21063), .B1(n21062), .B2(n16695), .ZN(
        n21065) );
  INV_X1 U23984 ( .A(n21065), .ZN(n21066) );
  OAI211_X1 U23985 ( .C1(n21069), .C2(n21068), .A(n21067), .B(n21066), .ZN(
        n21232) );
  AOI22_X1 U23986 ( .A1(n21072), .A2(keyinput28), .B1(keyinput21), .B2(n21071), 
        .ZN(n21070) );
  OAI221_X1 U23987 ( .B1(n21072), .B2(keyinput28), .C1(n21071), .C2(keyinput21), .A(n21070), .ZN(n21103) );
  INV_X1 U23988 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n21075) );
  INV_X1 U23989 ( .A(keyinput35), .ZN(n21074) );
  AOI22_X1 U23990 ( .A1(n21075), .A2(keyinput3), .B1(
        P3_INSTQUEUE_REG_15__5__SCAN_IN), .B2(n21074), .ZN(n21073) );
  OAI221_X1 U23991 ( .B1(n21075), .B2(keyinput3), .C1(n21074), .C2(
        P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(n21073), .ZN(n21102) );
  INV_X1 U23992 ( .A(keyinput14), .ZN(n21083) );
  INV_X1 U23993 ( .A(keyinput8), .ZN(n21080) );
  INV_X1 U23994 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n21077) );
  AOI22_X1 U23995 ( .A1(n21078), .A2(keyinput56), .B1(n21077), .B2(keyinput44), 
        .ZN(n21076) );
  OAI221_X1 U23996 ( .B1(n21078), .B2(keyinput56), .C1(n21077), .C2(keyinput44), .A(n21076), .ZN(n21079) );
  AOI221_X1 U23997 ( .B1(keyinput8), .B2(n21081), .C1(n21080), .C2(
        BUF1_REG_16__SCAN_IN), .A(n21079), .ZN(n21082) );
  OAI221_X1 U23998 ( .B1(keyinput14), .B2(n21084), .C1(n21083), .C2(
        P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(n21082), .ZN(n21101) );
  INV_X1 U23999 ( .A(keyinput41), .ZN(n21086) );
  OAI22_X1 U24000 ( .A1(keyinput32), .A2(n21087), .B1(n21086), .B2(
        P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n21085) );
  AOI221_X1 U24001 ( .B1(n21087), .B2(keyinput32), .C1(n21086), .C2(
        P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(n21085), .ZN(n21099) );
  OAI22_X1 U24002 ( .A1(n12578), .A2(keyinput40), .B1(n21089), .B2(keyinput43), 
        .ZN(n21088) );
  AOI221_X1 U24003 ( .B1(n12578), .B2(keyinput40), .C1(keyinput43), .C2(n21089), .A(n21088), .ZN(n21098) );
  INV_X1 U24004 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n21092) );
  INV_X1 U24005 ( .A(keyinput33), .ZN(n21091) );
  OAI22_X1 U24006 ( .A1(n21092), .A2(keyinput19), .B1(n21091), .B2(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n21090) );
  AOI221_X1 U24007 ( .B1(n21092), .B2(keyinput19), .C1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .C2(n21091), .A(n21090), .ZN(n21097)
         );
  XOR2_X1 U24008 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B(keyinput5), .Z(
        n21095) );
  XNOR2_X1 U24009 ( .A(n21093), .B(keyinput60), .ZN(n21094) );
  NOR2_X1 U24010 ( .A1(n21095), .A2(n21094), .ZN(n21096) );
  NAND4_X1 U24011 ( .A1(n21099), .A2(n21098), .A3(n21097), .A4(n21096), .ZN(
        n21100) );
  NOR4_X1 U24012 ( .A1(n21103), .A2(n21102), .A3(n21101), .A4(n21100), .ZN(
        n21230) );
  AOI22_X1 U24013 ( .A1(n21106), .A2(keyinput12), .B1(keyinput55), .B2(n21105), 
        .ZN(n21104) );
  OAI221_X1 U24014 ( .B1(n21106), .B2(keyinput12), .C1(n21105), .C2(keyinput55), .A(n21104), .ZN(n21119) );
  INV_X1 U24015 ( .A(keyinput47), .ZN(n21108) );
  AOI22_X1 U24016 ( .A1(n21109), .A2(keyinput34), .B1(P3_EBX_REG_3__SCAN_IN), 
        .B2(n21108), .ZN(n21107) );
  OAI221_X1 U24017 ( .B1(n21109), .B2(keyinput34), .C1(n21108), .C2(
        P3_EBX_REG_3__SCAN_IN), .A(n21107), .ZN(n21118) );
  INV_X1 U24018 ( .A(READY1), .ZN(n21112) );
  INV_X1 U24019 ( .A(keyinput50), .ZN(n21111) );
  AOI22_X1 U24020 ( .A1(n21112), .A2(keyinput1), .B1(P1_DATAO_REG_5__SCAN_IN), 
        .B2(n21111), .ZN(n21110) );
  OAI221_X1 U24021 ( .B1(n21112), .B2(keyinput1), .C1(n21111), .C2(
        P1_DATAO_REG_5__SCAN_IN), .A(n21110), .ZN(n21117) );
  AOI22_X1 U24022 ( .A1(n21115), .A2(keyinput54), .B1(keyinput45), .B2(n21114), 
        .ZN(n21113) );
  OAI221_X1 U24023 ( .B1(n21115), .B2(keyinput54), .C1(n21114), .C2(keyinput45), .A(n21113), .ZN(n21116) );
  NOR4_X1 U24024 ( .A1(n21119), .A2(n21118), .A3(n21117), .A4(n21116), .ZN(
        n21229) );
  INV_X1 U24025 ( .A(keyinput39), .ZN(n21121) );
  OAI22_X1 U24026 ( .A1(n21122), .A2(keyinput59), .B1(n21121), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n21120) );
  AOI221_X1 U24027 ( .B1(n21122), .B2(keyinput59), .C1(BUF2_REG_21__SCAN_IN), 
        .C2(n21121), .A(n21120), .ZN(n21133) );
  INV_X1 U24028 ( .A(keyinput13), .ZN(n21124) );
  OAI22_X1 U24029 ( .A1(n21125), .A2(keyinput29), .B1(n21124), .B2(
        P3_EBX_REG_2__SCAN_IN), .ZN(n21123) );
  AOI221_X1 U24030 ( .B1(n21125), .B2(keyinput29), .C1(P3_EBX_REG_2__SCAN_IN), 
        .C2(n21124), .A(n21123), .ZN(n21132) );
  INV_X1 U24031 ( .A(keyinput30), .ZN(n21127) );
  OAI22_X1 U24032 ( .A1(keyinput4), .A2(n21128), .B1(n21127), .B2(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n21126) );
  AOI221_X1 U24033 ( .B1(n21128), .B2(keyinput4), .C1(n21127), .C2(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(n21126), .ZN(n21131) );
  XOR2_X1 U24034 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B(keyinput0), .Z(
        n21129) );
  AOI21_X1 U24035 ( .B1(keyinput10), .B2(n12673), .A(n21129), .ZN(n21130) );
  NAND4_X1 U24036 ( .A1(n21133), .A2(n21132), .A3(n21131), .A4(n21130), .ZN(
        n21166) );
  INV_X1 U24037 ( .A(keyinput42), .ZN(n21135) );
  OAI22_X1 U24038 ( .A1(n21136), .A2(keyinput2), .B1(n21135), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n21134) );
  AOI221_X1 U24039 ( .B1(n21136), .B2(keyinput2), .C1(P1_LWORD_REG_2__SCAN_IN), 
        .C2(n21135), .A(n21134), .ZN(n21148) );
  INV_X1 U24040 ( .A(keyinput38), .ZN(n21138) );
  OAI22_X1 U24041 ( .A1(keyinput18), .A2(n21139), .B1(n21138), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n21137) );
  AOI221_X1 U24042 ( .B1(n21139), .B2(keyinput18), .C1(n21138), .C2(
        P1_LWORD_REG_0__SCAN_IN), .A(n21137), .ZN(n21147) );
  INV_X1 U24043 ( .A(keyinput62), .ZN(n21141) );
  OAI22_X1 U24044 ( .A1(n13677), .A2(keyinput26), .B1(n21141), .B2(
        P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n21140) );
  AOI221_X1 U24045 ( .B1(n13677), .B2(keyinput26), .C1(
        P3_INSTQUEUE_REG_9__2__SCAN_IN), .C2(n21141), .A(n21140), .ZN(n21146)
         );
  INV_X1 U24046 ( .A(DATAI_30_), .ZN(n21144) );
  INV_X1 U24047 ( .A(keyinput61), .ZN(n21143) );
  OAI22_X1 U24048 ( .A1(n21144), .A2(keyinput24), .B1(n21143), .B2(
        P3_REIP_REG_30__SCAN_IN), .ZN(n21142) );
  AOI221_X1 U24049 ( .B1(n21144), .B2(keyinput24), .C1(P3_REIP_REG_30__SCAN_IN), .C2(n21143), .A(n21142), .ZN(n21145) );
  NAND4_X1 U24050 ( .A1(n21148), .A2(n21147), .A3(n21146), .A4(n21145), .ZN(
        n21165) );
  INV_X1 U24051 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21150) );
  AOI22_X1 U24052 ( .A1(n21150), .A2(keyinput57), .B1(n12413), .B2(keyinput16), 
        .ZN(n21149) );
  OAI221_X1 U24053 ( .B1(n21150), .B2(keyinput57), .C1(n12413), .C2(keyinput16), .A(n21149), .ZN(n21164) );
  INV_X1 U24054 ( .A(keyinput20), .ZN(n21152) );
  OAI22_X1 U24055 ( .A1(keyinput49), .A2(n21153), .B1(n21152), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21151) );
  AOI221_X1 U24056 ( .B1(n21153), .B2(keyinput49), .C1(n21152), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n21151), .ZN(n21162) );
  INV_X1 U24057 ( .A(keyinput36), .ZN(n21155) );
  OAI22_X1 U24058 ( .A1(keyinput58), .A2(n21156), .B1(n21155), .B2(
        P3_REIP_REG_21__SCAN_IN), .ZN(n21154) );
  AOI221_X1 U24059 ( .B1(n21156), .B2(keyinput58), .C1(n21155), .C2(
        P3_REIP_REG_21__SCAN_IN), .A(n21154), .ZN(n21161) );
  INV_X1 U24060 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21159) );
  OAI22_X1 U24061 ( .A1(n21159), .A2(keyinput15), .B1(n21158), .B2(keyinput51), 
        .ZN(n21157) );
  AOI221_X1 U24062 ( .B1(n21159), .B2(keyinput15), .C1(keyinput51), .C2(n21158), .A(n21157), .ZN(n21160) );
  NAND3_X1 U24063 ( .A1(n21162), .A2(n21161), .A3(n21160), .ZN(n21163) );
  NOR4_X1 U24064 ( .A1(n21166), .A2(n21165), .A3(n21164), .A4(n21163), .ZN(
        n21228) );
  NOR2_X1 U24065 ( .A1(keyinput14), .A2(keyinput8), .ZN(n21172) );
  NAND2_X1 U24066 ( .A1(keyinput44), .A2(keyinput5), .ZN(n21170) );
  NOR3_X1 U24067 ( .A1(keyinput45), .A2(keyinput3), .A3(keyinput28), .ZN(
        n21168) );
  NOR3_X1 U24068 ( .A1(keyinput21), .A2(keyinput41), .A3(keyinput19), .ZN(
        n21167) );
  NAND4_X1 U24069 ( .A1(keyinput35), .A2(n21168), .A3(keyinput32), .A4(n21167), 
        .ZN(n21169) );
  NOR4_X1 U24070 ( .A1(keyinput40), .A2(keyinput60), .A3(n21170), .A4(n21169), 
        .ZN(n21171) );
  NAND4_X1 U24071 ( .A1(keyinput33), .A2(keyinput56), .A3(n21172), .A4(n21171), 
        .ZN(n21194) );
  NOR3_X1 U24072 ( .A1(keyinput22), .A2(keyinput53), .A3(keyinput17), .ZN(
        n21192) );
  NOR2_X1 U24073 ( .A1(keyinput43), .A2(keyinput27), .ZN(n21173) );
  NAND3_X1 U24074 ( .A1(keyinput9), .A2(keyinput23), .A3(n21173), .ZN(n21177)
         );
  NAND3_X1 U24075 ( .A1(keyinput7), .A2(keyinput52), .A3(keyinput37), .ZN(
        n21176) );
  NOR2_X1 U24076 ( .A1(keyinput46), .A2(keyinput6), .ZN(n21174) );
  NAND3_X1 U24077 ( .A1(keyinput11), .A2(keyinput25), .A3(n21174), .ZN(n21175)
         );
  NOR4_X1 U24078 ( .A1(keyinput63), .A2(n21177), .A3(n21176), .A4(n21175), 
        .ZN(n21191) );
  NAND4_X1 U24079 ( .A1(keyinput38), .A2(keyinput26), .A3(keyinput62), .A4(
        keyinput61), .ZN(n21189) );
  NAND3_X1 U24080 ( .A1(keyinput13), .A2(keyinput39), .A3(keyinput59), .ZN(
        n21179) );
  NAND3_X1 U24081 ( .A1(keyinput30), .A2(keyinput2), .A3(keyinput42), .ZN(
        n21178) );
  NOR4_X1 U24082 ( .A1(keyinput4), .A2(keyinput18), .A3(n21179), .A4(n21178), 
        .ZN(n21181) );
  INV_X1 U24083 ( .A(keyinput48), .ZN(n21180) );
  NAND4_X1 U24084 ( .A1(keyinput29), .A2(keyinput0), .A3(n21181), .A4(n21180), 
        .ZN(n21188) );
  NOR3_X1 U24085 ( .A1(keyinput58), .A2(keyinput36), .A3(keyinput15), .ZN(
        n21183) );
  NOR3_X1 U24086 ( .A1(keyinput34), .A2(keyinput1), .A3(keyinput54), .ZN(
        n21182) );
  NAND4_X1 U24087 ( .A1(keyinput16), .A2(n21183), .A3(keyinput50), .A4(n21182), 
        .ZN(n21187) );
  NOR2_X1 U24088 ( .A1(keyinput24), .A2(keyinput20), .ZN(n21185) );
  NOR4_X1 U24089 ( .A1(keyinput51), .A2(keyinput12), .A3(keyinput55), .A4(
        keyinput47), .ZN(n21184) );
  NAND4_X1 U24090 ( .A1(keyinput49), .A2(keyinput57), .A3(n21185), .A4(n21184), 
        .ZN(n21186) );
  NOR4_X1 U24091 ( .A1(n21189), .A2(n21188), .A3(n21187), .A4(n21186), .ZN(
        n21190) );
  NAND4_X1 U24092 ( .A1(keyinput31), .A2(n21192), .A3(n21191), .A4(n21190), 
        .ZN(n21193) );
  OAI21_X1 U24093 ( .B1(n21194), .B2(n21193), .A(keyinput10), .ZN(n21226) );
  INV_X1 U24094 ( .A(keyinput25), .ZN(n21196) );
  OAI22_X1 U24095 ( .A1(keyinput53), .A2(n21197), .B1(n21196), .B2(
        P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n21195) );
  AOI221_X1 U24096 ( .B1(n21197), .B2(keyinput53), .C1(n21196), .C2(
        P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(n21195), .ZN(n21208) );
  INV_X1 U24097 ( .A(keyinput22), .ZN(n21199) );
  OAI22_X1 U24098 ( .A1(n10649), .A2(keyinput17), .B1(n21199), .B2(
        P3_ADDRESS_REG_11__SCAN_IN), .ZN(n21198) );
  AOI221_X1 U24099 ( .B1(n10649), .B2(keyinput17), .C1(
        P3_ADDRESS_REG_11__SCAN_IN), .C2(n21199), .A(n21198), .ZN(n21207) );
  INV_X1 U24100 ( .A(keyinput6), .ZN(n21201) );
  OAI22_X1 U24101 ( .A1(n21202), .A2(keyinput48), .B1(n21201), .B2(DATAI_15_), 
        .ZN(n21200) );
  AOI221_X1 U24102 ( .B1(n21202), .B2(keyinput48), .C1(DATAI_15_), .C2(n21201), 
        .A(n21200), .ZN(n21206) );
  OAI22_X1 U24103 ( .A1(n12188), .A2(keyinput11), .B1(n21204), .B2(keyinput46), 
        .ZN(n21203) );
  AOI221_X1 U24104 ( .B1(n12188), .B2(keyinput11), .C1(keyinput46), .C2(n21204), .A(n21203), .ZN(n21205) );
  NAND4_X1 U24105 ( .A1(n21208), .A2(n21207), .A3(n21206), .A4(n21205), .ZN(
        n21225) );
  INV_X1 U24106 ( .A(keyinput23), .ZN(n21210) );
  OAI22_X1 U24107 ( .A1(n10351), .A2(keyinput7), .B1(n21210), .B2(
        P3_UWORD_REG_10__SCAN_IN), .ZN(n21209) );
  AOI221_X1 U24108 ( .B1(n10351), .B2(keyinput7), .C1(P3_UWORD_REG_10__SCAN_IN), .C2(n21210), .A(n21209), .ZN(n21223) );
  INV_X1 U24109 ( .A(keyinput9), .ZN(n21212) );
  OAI22_X1 U24110 ( .A1(n21213), .A2(keyinput27), .B1(n21212), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n21211) );
  AOI221_X1 U24111 ( .B1(n21213), .B2(keyinput27), .C1(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n21212), .A(n21211), .ZN(
        n21222) );
  INV_X1 U24112 ( .A(keyinput31), .ZN(n21215) );
  OAI22_X1 U24113 ( .A1(keyinput37), .A2(n21216), .B1(n21215), .B2(
        P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n21214) );
  AOI221_X1 U24114 ( .B1(n21216), .B2(keyinput37), .C1(n21215), .C2(
        P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(n21214), .ZN(n21221) );
  OAI22_X1 U24115 ( .A1(n21219), .A2(keyinput63), .B1(n21218), .B2(keyinput52), 
        .ZN(n21217) );
  AOI221_X1 U24116 ( .B1(n21219), .B2(keyinput63), .C1(keyinput52), .C2(n21218), .A(n21217), .ZN(n21220) );
  NAND4_X1 U24117 ( .A1(n21223), .A2(n21222), .A3(n21221), .A4(n21220), .ZN(
        n21224) );
  AOI211_X1 U24118 ( .C1(P2_REIP_REG_3__SCAN_IN), .C2(n21226), .A(n21225), .B(
        n21224), .ZN(n21227) );
  NAND4_X1 U24119 ( .A1(n21230), .A2(n21229), .A3(n21228), .A4(n21227), .ZN(
        n21231) );
  XNOR2_X1 U24120 ( .A(n21232), .B(n21231), .ZN(P1_U2984) );
  NAND2_X1 U11387 ( .A1(n11243), .A2(n11242), .ZN(n13334) );
  NOR2_X2 U11044 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10202) );
  CLKBUF_X1 U11097 ( .A(n14422), .Z(n9609) );
  CLKBUF_X1 U11110 ( .A(n14629), .Z(n14630) );
  CLKBUF_X1 U11154 ( .A(n15725), .Z(n15758) );
  CLKBUF_X3 U11311 ( .A(n14284), .Z(n17900) );
  CLKBUF_X1 U11316 ( .A(n14547), .Z(n14548) );
  CLKBUF_X1 U11390 ( .A(n19892), .Z(n19900) );
  CLKBUF_X1 U11987 ( .A(n10450), .Z(n17033) );
  CLKBUF_X1 U12262 ( .A(n19899), .Z(n19889) );
  CLKBUF_X1 U12263 ( .A(n18129), .Z(n19569) );
  CLKBUF_X1 U12357 ( .A(n18196), .Z(n18205) );
endmodule

