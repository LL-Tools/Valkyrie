
module b22_C_2inp_gates_syn ( 
    P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
    SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_,
    SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_,
    SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
    P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
    P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
    P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
    P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
    P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
    P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
    P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
    P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
    P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
    P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
    P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
    P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
    P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
    P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
    P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
    P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
    P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
    P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
    P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
    P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
    P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
    P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
    P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
    P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
    P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
    P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
    P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
    P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
    P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
    P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN,
    P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
    P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
    P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
    P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
    P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
    P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
    P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
    P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
    P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
    P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
    P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
    P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
    P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
    P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
    P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
    P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
    P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
    P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
    P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
    P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
    P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
    P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
    P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
    P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
    P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
    P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
    P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
    P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
    P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
    P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
    P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
    P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
    P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
    P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
    P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
    P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
    P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
    P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
    P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
    P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
    P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
    P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
    P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
    P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
    P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
    P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
    P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
    P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
    P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
    P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
    P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
    P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
    P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
    P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
    P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
    P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
    P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
    P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
    P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
    P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
    P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
    P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
    P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
    P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
    P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
    P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
    P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
    P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
    P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
    P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
    P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
    P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
    P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
    P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
    P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
    P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
    P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
    P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
    P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
    P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
    P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
    P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
    P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
    P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
    P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
    P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
    P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
    P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
    P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
    P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
    P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
    P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
    P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
    P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
    P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
    P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
    P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
    P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
    P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
    P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
    P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
    P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
    P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
    P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
    P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
    P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
    P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
    P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
    P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
    P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
    P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
    P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
    P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
    P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
    P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
    P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
    P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
    P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
    P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
    P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
    P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
    P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
    P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
    P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
    P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
    P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
    P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
    P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
    P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN,
    SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
    SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
    SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
    SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
    U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
    P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
    P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
    P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
    P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
    P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
    P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
    P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
    P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
    P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
    P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
    P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
    P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
    P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
    P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
    P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
    P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
    P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
    P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
    P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
    P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
    P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
    P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
    P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
    P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
    P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
    P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
    P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
    P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
    P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
    P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
    P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
    P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
    P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
    P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
    P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
    P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
    P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
    P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
    P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
    P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
    P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
    P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
    P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
    P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
    P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
    P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
    P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
    P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
    P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
    P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
    P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
    P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
    P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
    P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
    P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
    P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
    P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
    P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
    P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
    P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
    P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
    P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
    P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
    P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
    P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
    P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
    P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
    P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
    P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
    P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
    P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
    P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
    P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
    P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
    P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
    P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
    P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
    P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
    P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
    P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
    P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
    P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
    P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
    P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
    P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
    P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
    P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
    P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
    P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
    P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
    P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
    P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
    P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
    P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
    P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
    P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
    P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
    P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
    P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
    P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
    P3_U3897  );
  input  P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_,
    SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
    SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
    SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
    P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
    P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
    P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
    P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
    P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
    P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
    P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
    P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
    P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
    P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
    P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
    P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
    P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
    P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
    P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
    P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
    P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
    P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
    P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
    P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
    P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
    P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
    P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
    P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
    P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
    P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
    P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
    P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
    P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
    P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN,
    P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
    P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
    P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
    P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
    P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
    P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
    P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
    P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
    P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
    P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
    P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
    P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
    P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
    P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
    P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
    P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
    P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
    P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
    P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
    P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
    P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
    P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
    P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
    P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
    P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
    P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
    P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
    P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
    P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
    P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
    P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
    P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
    P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
    P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
    P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
    P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
    P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
    P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
    P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
    P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
    P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
    P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
    P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
    P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
    P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
    P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
    P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
    P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
    P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
    P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
    P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
    P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
    P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
    P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
    P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
    P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
    P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
    P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
    P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
    P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
    P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
    P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
    P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
    P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
    P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
    P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
    P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
    P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
    P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
    P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
    P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
    P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
    P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
    P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
    P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
    P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
    P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
    P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
    P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
    P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
    P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
    P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
    P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
    P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
    P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
    P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
    P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
    P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
    P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
    P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
    P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
    P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
    P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
    P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
    P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
    P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
    P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
    P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
    P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
    P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
    P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
    P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
    P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
    P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
    P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
    P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
    P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
    P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
    P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
    P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
    P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
    P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
    P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
    P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
    P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
    P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
    P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
    P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
    P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
    P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
    P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
    P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
    P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
    P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
    P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
    P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
    P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
    P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
    P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
    SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
    SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
    SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
    U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
    P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
    P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
    P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
    P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
    P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
    P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
    P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
    P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
    P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
    P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
    P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
    P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
    P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
    P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
    P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
    P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
    P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
    P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
    P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
    P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
    P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
    P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
    P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
    P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
    P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
    P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
    P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
    P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
    P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
    P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
    P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
    P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
    P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
    P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
    P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
    P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
    P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
    P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
    P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
    P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
    P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
    P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
    P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
    P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
    P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
    P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
    P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
    P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
    P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
    P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
    P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
    P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
    P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
    P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
    P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
    P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
    P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
    P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
    P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
    P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
    P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
    P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
    P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
    P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
    P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
    P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
    P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
    P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
    P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
    P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
    P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
    P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
    P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
    P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
    P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
    P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
    P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
    P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
    P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
    P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
    P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
    P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
    P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
    P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
    P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
    P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
    P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
    P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
    P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
    P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
    P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
    P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
    P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
    P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
    P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
    P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
    P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
    P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
    P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
    P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
    P3_U3897;
  wire n25267, n24316, n14111, n13133, n25489, n25214, n21353, n26252,
    n13124, n21402, n26152, n13116, n26459, n16572, n15554, n13134, n19178,
    n14091, n14654, n15113, n13563, n21975, n25264, n17487, n23967, n24190,
    n17312, n13866, n20556, n21598, n25104, n22889, n23906, n22998, n24213,
    n24131, n26205, n25389, n25284, n16928, n13118, n16337, n13119, n13120,
    n14511, n15008, n13987, n18666, n14933, n14923, n13527, n13123, n18563,
    n24449, n21032, n25884, n19816, n19033, n25921, n19985, n15111, n13121,
    n13122, n16232, n24516, n22544, n18026, n19334, n26335, n16343, n14836,
    n20065, n20066, n25800, n13867, n22234, n19176, n18900, n13611, n14630,
    n18805, n21910, n22905, n21932, n22618, n15689, n22041, n15630, n13582,
    n23264, n15133, n18649, n21377, n23818, n21309, n24000, n15647, n23903,
    n25420, n13794, n24319, n15219, n15270, n23132, n18501, n17049, n23905,
    n17036, n13970, n13734, n18497, n18141, n22076, n22458, n22841, n14255,
    n20589, n13872, n13698, n20117, n20110, n18080, n14116, n19630, n18904,
    n13830, n13449, n21676, n22472, n23171, n14848, n23173, n13619, n19003,
    n21333, n22174, n23114, n13668, n19095, n14398, n22132, n13671, n21487,
    n22632, n13787, n13503, n22832, n14631, n13673, n14622, n26030, n23137,
    n20197, n22819, n26005, n19994, n22604, n21921, n13901, n22617, n22495,
    n18020, n21965, n20976, n21954, n21660, n22728, n15637, n22862, n24950,
    n17423, n17691, n15693, n17463, n22746, n13451, n14820, n21986, n21997,
    n20892, n22664, n13714, n17679, n17346, n22029, n20349, n14443, n23015,
    n15629, n22295, n17664, n18041, n14828, n15660, n26182, n14446, n22018,
    n23203, n14163, n24982, n24473, n23740, n22341, n20209, n24308, n24394,
    n23051, n25506, n23831, n13552, n15486, n25067, n24231, n13142, n25479,
    n13125, n14499, n25882, n18877, n19980, n13666, n25454, n15372, n25240,
    n25330, n25150, n25114, n24976, n13196, n23872, n23278, n14032, n25689,
    n26212, n23753, n23825, n23853, n22790, n13583, n13888, n25021, n25049,
    n25126, n25432, n25252, n25254, n25274, n15640, n15046, n15122, n23854,
    n14503, n17357, n14991, n17382, n23993, n26351, n26086, n26085, n26343,
    n26229, n26245, n16941, n15021, n15860, n13614, n13480, n25841, n14500,
    n25771, n14810, n18385, n15859, n26287, n26286, n25399, n19975, n14581,
    n21356, n14109, n13915, n16939, n18547, n22139, n13129, n15559, n16777,
    n16780, n18920, n13525, n15036, n16460, n14175, n14430, n14930, n16851,
    n19868, n14100, n14935, n16484, n15033, n17502, n17657, n15339, n22133,
    n25802, n15309, n19847, n18861, n24333, n20773, n15371, n15175, n14580,
    n15034, n19809, n23156, n15387, n16110, n18854, n17071, n20794, n15206,
    n15078, n15354, n13128, n14938, n20752, n23723, n17632, n16471, n19840,
    n17597, n15452, n16574, n14959, n14960, n14963, n13537, n14922, n14890,
    n14889, n16074, n15962, n15963, n15992, n14891, n14892, n15991, n14962,
    n19806, n15958, n15990, n15988, n14887, n14888, n14886, n14894, n14893,
    n15014, n15668, n15011, n17359, n13126, n13127, n15451, n18512, n15167,
    n15085, n13795, n15865, n13130, n13131, n15421, n22817, n22450, n13132,
    n21460, n17873, n18545, n14983, n14087, n13589, n14444, n14445, n14629,
    n14073, n14450, n14451, n14455, n14663, n13543, n17365, n15450, n13545,
    n14329, n18627, n14162, n21219, n14594, n14596, n14609, n21240, n14565,
    n14837, n19479, n13939, n14710, n14823, n13781, n14456, n14457, n14148,
    n18549, n15719, n16106, n13651, n13652, n20184, n18255, n14310, n14464,
    n14085, n14088, n14387, n13884, n13153, n14279, n14758, n14640, n17814,
    n14074, n14765, n14448, n24997, n17790, n14366, n14041, n14665, n14770,
    n14772, n14512, n14513, n13623, n14783, n18876, n14784, n14096, n15662,
    n15543, n13420, n14338, n14339, n19253, n17198, n19222, n13439, n13440,
    n14745, n14746, n20478, n17152, n14053, n14054, n14055, n13434, n13435,
    n13436, n13703, n17565, n14489, n14490, n14491, n16031, n14121, n21031,
    n13984, n13985, n21619, n21323, n13539, n14628, n21664, n13988, n21744,
    n13677, n13679, n14072, n14453, n13773, n13772, n17954, n17014, n13881,
    n18901, n13721, n13599, n14781, n14393, n22223, n14395, n13916, n13917,
    n18046, n17366, n22457, n23991, n14419, n15546, n16095, n13653, n14187,
    n25995, n14269, n18351, n19228, n16789, n13705, n17058, n13824, n13825,
    n16878, n16587, n17961, n17955, n14164, n15418, n13973, n13609, n15553,
    n18865, n14297, n13889, n15448, n13809, n13810, n23189, n14603, n16548,
    n13483, n13484, n13485, n17881, n19314, n14556, n21071, n14012, n14027,
    n13817, n14025, n14599, n14141, n21218, n19452, n14796, n13469, n13905,
    n14607, n18535, n18537, n14154, n13902, n13940, n14360, n13834, n13833,
    n21328, n21437, n13410, n14460, n18881, n13687, n13688, n13689, n18279,
    n19460, n14853, n19315, n19312, n15983, n14089, n13158, n14760, n14183,
    n14316, n14318, n14768, n19248, n13903, n13862, n13759, n20108, n13441,
    n14832, n14224, n13446, n13922, n18302, n14750, n14751, n14842, n13576,
    n13577, n20374, n14216, n14218, n14841, n14202, n18202, n14821, n13566,
    n14822, n18189, n14220, n19335, n19327, n17140, n14487, n14480, n14302,
    n14812, n14286, n14287, n14611, n14267, n13813, n14171, n21446, n14642,
    n17486, n14755, n14756, n14374, n14375, n14623, n14624, n14639, n14180,
    n14181, n17678, n21681, n17816, n14643, n14646, n14764, n21868, n14637,
    n17564, n25076, n25135, n25155, n14432, n14433, n17508, n13836, n18899,
    n13690, n15697, n14043, n18021, n18045, n13636, n14657, n14123, n14124,
    n14400, n14402, n13800, n13801, n13502, n14785, n23772, n17389, n13629,
    n15751, n14136, n14135, n15805, n14700, n13548, n14493, n14498, n14958,
    n14957, n16094, n16093, n14573, n16314, n13424, n17942, n19493, n19494,
    n14331, n14190, n14334, n14336, n13648, n14002, n19813, n14234, n14241,
    n14242, n14240, n18366, n13842, n20152, n13843, n18339, n13844, n18323,
    n20261, n16414, n26200, n19257, n26282, n18455, n20129, n20185, n18437,
    n13930, n13447, n20333, n14713, n13921, n14736, n18411, n14868, n19346,
    n14732, n14731, n26258, n18448, n13637, n13642, n18306, n18291, n14469,
    n18443, n17143, n17147, n14488, n14808, n14066, n14070, n16024, n17039,
    n14860, n17589, n14863, n21037, n16661, n24927, n13991, n21886, n25025,
    n25083, n21395, n21345, n21445, n21409, n14373, n13591, n13592, n14632,
    n17745, n17708, n21772, n21826, n21841, n24947, n25017, n17863, n15955,
    n16569, n14084, n15968, n15965, n15970, n15966, n15979, n14363, n14365,
    n13604, n23266, n15628, n14997, n15585, n15931, n13473, n14157, n13544,
    n13733, n19084, n13595, n13597, n14523, n14524, n22494, n14514, n22570,
    n14779, n18018, n15609, n18896, n14392, n14394, n22678, n14777, n14520,
    n17375, n23749, n24178, n18843, n15812, n13625, n13626, n13627, n14510,
    n22522, n23765, n23851, n13495, n13496, n14298, n14299, n13462, n15806,
    n13534, n15784, n15749, n14097, n14095, n14372, n14924, n15577, n13879,
    n14496, n14497, n15485, n15315, n15069, n13508, n13523, n14582, n14586,
    n17918, n13427, n19061, n14538, n20141, n14184, n14185, n25638, n25660,
    n20495, n19750, n19766, n14470, n14471, n14715, n19300, n14717, n14718,
    n14719, n18326, n14003, n13875, n13966, n14237, n19990, n13859, n13855,
    n19827, n26046, n14238, n14239, n20034, n20006, n20097, n13955, n13956,
    n13951, n13960, n18492, n20174, n14468, n18321, n18322, n26150, n20528,
    n26303, n18482, n17101, n16338, n14044, n17177, n13575, n14045, n17299,
    n14056, n14058, n14059, n14807, n13704, n16117, n14792, n21586, n14825,
    n14843, n14425, n18915, n14120, n17046, n20863, n14126, n24389, n17525,
    n21845, n21560, n24471, n13829, n24521, n21462, n14168, n17694, n17682,
    n16674, n16590, n18106, n18105, n14816, n22124, n14306, n15836, n15843,
    n25194, n15273, n13661, n15269, n14406, n13610, n22187, n13978, n14691,
    n14678, n14679, n14689, n22702, n15500, n15930, n14690, n22515, n15936,
    n13616, n13481, n13725, n23552, n23623, n14246, n23655, n13729, n23706,
    n22421, n17982, n22422, n22452, n22429, n18070, n13541, n15757, n14035,
    n22952, n14271, n24015, n22414, n22810, n18135, n14653, n24034, n24033,
    n14300, n14293, n14294, n14296, n14295, n17975, n14146, n14587, n14176,
    n16101, n13486, n17315, n23164, n17924, n13516, n13518, n13517, n20656,
    n18223, n26138, n18436, n20665, n18216, n20648, n25964, n18253, n26297,
    n25093, n14602, n14327, n21456, n14112, n23331, n14414, n13684, n14105,
    n14412, n23493, n14243, n14244, n23729, n13553, n13551, n13412, n23166,
    n23192, n19313, n19333, n21070, n13471, n21090, n14368, n14410, n14411,
    n14026, n14548, n18626, n14595, n21168, n14567, n13466, n13464, n14798,
    n14799, n19450, n13822, n13821, n14561, n14791, n14417, n14021, n14153,
    n21259, n19288, n13904, n13411, n13478, n13693, n13694, n13695, n14563,
    n14382, n13590, n14321, n14323, n19160, n14226, n14223, n14833, n14749,
    n13927, n13926, n14214, n14215, n14212, n14213, n14727, n14729, n14730,
    n13569, n13573, n13570, n13571, n13572, n14206, n14207, n14813, n13832,
    n14361, n14877, n13838, n14614, n14358, n21365, n14172, n21441, n21440,
    n14378, n14379, n14380, n14381, n14461, n13549, n14757, n14388, n14466,
    n14385, n14386, n14644, n14766, n14077, n14078, n14459, n13778, n18893,
    n13686, n13691, n13692, n14667, n14659, n14660, n17400, n14572, n19177,
    n14534, n14189, n14335, n14800, n13947, n13770, n13845, n13840, n13841,
    n13851, n13846, n13847, n19364, n13445, n13932, n13931, n13933, n20208,
    n18283, n20282, n13707, n13936, n14723, n14724, n14725, n14722, n14726,
    n14734, n14819, n14854, n19338, n14200, n14705, n14703, n18297, n16954,
    n15987, n14802, n14803, n13452, n14313, n21444, n13674, n17734, n14619,
    n14620, n14625, n14465, n13675, n13676, n13678, n14454, n13682, n14440,
    n14441, n25045, n25120, n14617, n25209, n14081, n14083, n14080, n13774,
    n13775, n13776, n13777, n15961, n14139, n15959, n14282, n16037, n15123,
    n14150, n14407, n14506, n14507, n15851, n13492, n14505, n23777, n13621,
    n13498, n14030, n23926, n15750, n14098, n15716, n14699, n13432, n13429,
    n19138, n14535, n19135, n13641, n14188, n13657, n13658, n13654, n13643,
    n13907, n13877, n14235, n13858, n19822, n25974, n14232, n14233, n13860,
    n13861, n13863, n16063, n13760, n13763, n20082, n13753, n17091, n16899,
    n16798, n16529, n16501, n16491, n13850, n16363, n14198, n16373, n16376,
    n16425, n13852, n26256, n26279, n19503, n18365, n20144, n14831, n19295,
    n20142, n14742, n13562, n14861, n20205, n20233, n20293, n20331, n20352,
    n20385, n20387, n13706, n18425, n14838, n13574, n14740, n14733, n26054,
    n14818, n26076, n26126, n26233, n26273, n14549, n14550, n14330, n14483,
    n14476, n14478, n16039, n16034, n16027, n14793, n14794, n16021, n18939,
    n18937, n13458, n14846, n14847, n14132, n14127, n14128, n14129, n14301,
    n13459, n14849, n14851, n14850, n24489, n24488, n18936, n17533, n14283,
    n14284, n14165, n14166, n14167, n13828, n21455, n21449, n24741, n15957,
    n17758, n21597, n17737, n17722, n17711, n17685, n16751, n17578, n25245,
    n21609, n21631, n21661, n14177, n21694, n21757, n21790, n21843, n13681,
    n14634, n24948, n14449, n25077, n14431, n25219, n25217, n14817, n25241,
    n15830, n14138, n17613, n15267, n17569, n13975, n15730, n14692, n13979,
    n14680, n14677, n14673, n15646, n15654, n15650, n15353, n14697, n15815,
    n15766, n15481, n15758, n15610, n14042, n15939, n14038, n13912, n22705,
    n22729, n13499, n13798, n22753, n14518, n14650, n14350, n22777, n15223,
    n13535, n13536, n13804, n14516, n15020, n13796, n13506, n14122, n13712,
    n22780, n14345, n23751, n23823, n14782, n23849, n23886, n23924, n15777,
    n15828, n15905, n15907, n15446, n14502, n15012, n14574, n13811, n13416,
    n13557, n13555, n13558, n13415, n13556, n13559, n13425, n17940, n13421,
    n13418, n19065, n19064, n25603, n14539, n14540, n14541, n19547, n14196,
    n25616, n25651, n19597, n19413, n20454, n19666, n16452, n16473, n19708,
    n26125, n19703, n19304, n19721, n19735, n13646, n25730, n20165, n13839,
    n20310, n20334, n20398, n25773, n25780, n13745, n14000, n14001, n25783,
    n13876, n13873, n13739, n25839, n25928, n25950, n25949, n25971, n26012,
    n19947, n19269, n14061, n18355, n20220, n18310, n18431, n18273, n20526,
    n26174, n20540, n19501, n18495, n20585, n18288, n13697, n20462, n26158,
    n26391, n17178, n18348, n14063, n16286, n16014, n19308, n17300, n17302,
    n17270, n13437, n16872, n16254, n16043, n14068, n13438, n16203, n16138,
    n14805, n16204, n18169, n16146, n16154, n16082, n16175, n24341, n17621,
    n14383, n21684, n17603, n17641, n14857, n14858, n17651, n25079, n24491,
    n13886, n21478, n16615, n14324, n24796, n21521, n21542, n16676, n16686,
    n16725, n17497, n17494, n25273, n25233, n25277, n18150, n18121, n21477,
    n14390, n14093, n14094, n21541, n14627, n14633, n21618, n14621, n21662,
    n18146, n17059, n14328, n16580, n17033, n22156, n17008, n17015, n15661,
    n21407, n17022, n13584, n13585, n17521, n17503, n22874, n23235, n13601,
    n13600, n13602, n15527, n15386, n14684, n14685, n15323, n14265, n14260,
    n15023, n22293, n13980, n13982, n23332, n17377, n18856, n14156, n14159,
    n13542, n18863, n22516, n22551, n16511, n13731, n23437, n23483, n14245,
    n23516, n23660, n14252, n23721, n14250, n14251, n14522, n22492, n22845,
    n13918, n14668, n22569, n22565, n14786, n22625, n13630, n14519, n14651,
    n22568, n17466, n15252, n15288, n23820, n13605, n13606, n15189, n13618,
    n24027, n22824, n24241, n24123, n15933, n14955, n22150, n15781, n22163,
    n15870, n14934, n14420, n14936, n15664, n13715, n15604, n14107, n14106,
    n13887, n15602, n15344, n13460, n13659, n14276, n16823, n14248, n23350,
    n16239, n16540, n13807, n13507, n16546, n13533, n13560, n16836, n13520,
    n13522, n17316, n17915, n13530, n19581, n20601, n25666, n20632, n18247,
    n20593, n26359, n20560, n19781, n14342, n25725, n14018, n14714, n14720,
    n14721, n26455, n26451, n26448, n26445, n26439, n26436, n20267, n19674,
    n19406, n19552, n26059, n26116, n26189, n16483, n26454, n25765, n25763,
    n25873, n13865, n13740, n26043, n13764, n13950, n13954, n13870, n20535,
    n19230, n18354, n13448, n20369, n14795, n26393, n26224, n26431, n26390,
    n14835, n20759, n20779, n18335, n14062, n20801, n18301, n19306, n17138,
    n17076, n14052, n16053, n18219, n16519, n14479, n18203, n16118, n20806,
    n14133, n14134, n21830, n13455, n24455, n14428, n18916, n20865, n20878,
    n24452, n14815, n24470, n24499, n25580, n25574, n25571, n25568, n25565,
    n25562, n25556, n21436, n21735, n21818, n21413, n21817, n24955, n25000,
    n25022, n24934, n13898, n21461, n13989, n21470, n25105, n25551, n25515,
    n25373, n14438, n23130, n17974, n15845, n22165, n17324, n25297, n25325,
    n15244, n13662, n22172, n22186, n14683, n23311, n15558, n23277, n24320,
    n24311, n24304, n24301, n22999, n23034, n23874, n13615, n13482, n13718,
    n13717, n23583, n13726, n13724, n23629, n13730, n23657, n23707, n22413,
    n22446, n14261, n14405, n22695, n23936, n24284, n13910, n24240, n14292,
    n14291, n23351, n15442, n24053, n24066, n24072, n24078, n24084, n16115,
    n16243, n13909, n13808, n13728, n14571, n17899, n14584, n13532, n19219,
    n14601, n14885, n13911, n14253, n16834, n14598, n15391, n13135, n18829,
    n18159, n13136, n21058, n13137, n21556, n13138, n14597, n13139, n16003,
    n13140, n13141, n19446, n13906, n19427, n13143, n17196, n13144, n13145,
    n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13154, n13155,
    n13156, n13157, n13159, n13160, n24298, n13716, n14752, n13161, n13162,
    n13163, n13164, n13779, n13165, n13166, n13167, n13168, n15518, n23801,
    n13169, n13170, n13171, n13172, n13981, n22589, n24295, n17029, n13173,
    n13174, n13175, n13176, n17897, n14662, n15530, n18050, n13177, n18125,
    n13178, n13179, n13180, n14709, n13181, n24052, n18176, n13182, n13183,
    n23254, n13184, n14289, n18340, n19273, n17704, n26442, n13185, n21359,
    n25697, n13186, n18860, n19545, n13187, n13188, n13189, n13190, n20461,
    n14570, n13191, n13192, n13193, n13194, n13195, n13197, n13198, n13199,
    n13200, n20163, n14834, n13201, n13202, n14577, n17944, n13203, n20539,
    n13596, n18887, n13204, n13205, n13206, n13207, n18544, n14463, n13208,
    n13209, n13210, n13211, n21582, n22264, n20405, n13212, n14462, n14384,
    n13213, n13214, n13215, n13216, n13217, n13218, n21544, n13219, n13220,
    n13221, n13222, n13223, n22491, n13224, n14525, n13225, n13226, n13227,
    n13228, n13229, n16583, n22535, n26383, n13581, n13230, n23769, n14344,
    n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n20881,
    n25577, n13239, n13240, n13786, n14158, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n14266, n25692, n20517, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
    n14515, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n14615,
    n13267, n13268, n19092, n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n14711, n14712, n20160, n14256,
    n13280, n13281, n26316, n14005, n13282, n13283, n20524, n19391, n13284,
    n13285, n16144, n13986, n13683, n13286, n13287, n13914, n19085, n14526,
    n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
    n14257, n18059, n17174, n13423, n17927, n13297, n13298, n13299, n17179,
    n24059, n13300, n13301, n13302, n13303, n13304, n13719, n13720, n22513,
    n14762, n14763, n22488, n13305, n26199, n13306, n13307, n21469, n13990,
    n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n20330, n13319, n13320, n13321, n16345, n13322, n13323,
    n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
    n14956, n15603, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
    n14839, n14840, n13340, n13341, n13342, n13343, n17399, n13344, n13345,
    n13346, n13347, n13348, n13349, n13350, n13351, n13352, n14033, n13353,
    n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
    n13363, n14193, n14194, n13364, n13365, n14790, n13366, n13367, n13368,
    n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
    n20257, n13934, n13378, n13379, n13380, n14701, n14702, n14494, n14495,
    n15904, n14090, n13885, n13381, n13538, n13598, n13493, n22008, n18779,
    n14434, n25673, n22775, n15901, n17631, n20492, n25028, n20452, n22745,
    n23794, n24967, n24365, n25118, n13382, n13383, n13384, n13385, n16076,
    n20376, n13386, n15443, n15445, n13387, n13388, n13723, n13389, n13390,
    n13511, n17037, n13391, n13392, n13393, n26053, n13394, n13874, n13395,
    n13396, n13397, n13398, n15605, n15573, n14688, n14809, n25270, n25246,
    n13399, n13400, n14236, n14137, n13401, n14079, n14521, n13402, n23940,
    n23949, n13403, n13404, n14604, n14173, n14174, n26129, n13405, n14605,
    n13406, n13407, n19835, n13408, n13409, n13793, n24565, n14424, n14568,
    n14004, n25503, n25378, n21916, n13992, n13995, n13413, n14108, n21532,
    n17310, n13711, n13567, n13554, n21432, n14376, n20007, n19819, n13744,
    n13414, n13999, n25779, n13586, n14357, n17259, n16838, n16839, n17934,
    n13417, n13419, n13422, n16926, n13893, n13426, n13428, n13430, n17905,
    n13431, n13433, n16049, n16052, n14484, n16058, n13701, n13919, n13442,
    n13443, n13444, n19013, n19009, n20960, n13454, n13450, n24354, n13453,
    n13789, n13456, n13457, n20849, n15268, n25342, n13461, n13463, n14909,
    n14950, n14527, n13465, n13467, n13470, n13468, n18718, n18551, n13472,
    n18822, n13474, n13475, n18772, n13476, n13477, n13513, n23191, n13479,
    n18599, n13487, n13488, n13489, n13490, n13491, n23878, n13494, n17362,
    n13497, n22652, n13500, n13501, n13504, n13802, n13505, n19078, n13509,
    n23188, n13510, n13512, n16320, n13514, n13561, n13896, n13515, n13519,
    n23198, n13521, n17257, n16937, n13524, n13550, n13529, n13806, n13526,
    n13528, n13531, n17945, n15222, n13540, n15600, n18902, n15631, n13546,
    n13547, n16835, n16316, n13713, n17254, n16073, n14228, n14227, n20206,
    n13564, n13565, n16539, n16543, n13568, n20470, n15998, n16002, n14219,
    n20372, n16114, n13579, n13578, n13580, n13878, n14492, n25302, n14117,
    n15370, n13587, n13588, n21507, n13593, n13594, n13603, n22320, n22221,
    n13607, n23848, n23873, n13608, n15308, n22200, n23307, n13612, n13613,
    n22703, n22633, n13617, n14517, n14788, n22649, n22648, n13622, n13620,
    n13624, n13628, n17384, n13633, n13631, n13632, n13634, n22770, n13635,
    n14530, n13638, n17205, n13639, n13640, n17213, n16000, n14706, n14704,
    n13645, n19130, n17236, n13644, n13650, n19706, n13647, n13649, n19594,
    n13655, n13656, n14588, n14591, n17520, n13660, n13664, n13663, n14439,
    n18477, n13670, n17828, n13667, n14626, n13669, n21584, n13672, n14645,
    n13680, n17811, n13685, n23845, n13696, n16275, n13699, n14475, n13700,
    n16249, n13702, n16050, n16137, n20384, n13708, n13710, n13709, n23181,
    n23183, n14401, n22871, n22904, n23541, n13722, n23596, n23708, n13727,
    n17260, n13732, n23464, n14508, n19100, n13735, n13736, n13737, n13738,
    n13993, n25821, n13996, n26028, n25860, n13741, n13742, n13743, n19967,
    n13746, n13751, n13747, n13748, n13749, n13750, n20105, n13752, n13757,
    n13754, n13755, n13756, n25943, n13758, n13762, n20039, n13761, n13768,
    n13765, n13766, n13767, n25904, n13769, n17611, n13771, n14759, n14075,
    n13780, n21555, n13782, n13783, n13784, n13785, n20988, n20920, n13788,
    n13790, n24377, n13791, n24340, n13792, n21000, n21001, n23941, n17948,
    n22749, n13797, n13799, n22588, n23852, n23829, n13803, n18144, n13805,
    n19060, n16929, n16933, n13908, n16109, n14613, n13812, n13814, n13815,
    n13816, n13818, n21234, n13819, n13820, n21228, n21408, n13823, n21454,
    n13826, n13827, n13831, n14359, n13835, n17023, n13837, n17025, n16852,
    n16374, n13848, n13849, n16386, n13853, n25945, n13854, n13856, n13857,
    n25983, n13864, n20062, n19971, n16089, n16339, n17180, n16958, n16160,
    n16139, n20128, n13868, n13869, n13871, n19977, n15544, n13880, n17834,
    n17872, n15408, n13882, n15375, n13883, n14618, n21640, n21707, n15574,
    n15579, n13890, n16923, n16924, n13891, n13892, n16930, n13894, n13895,
    n14575, n17894, n23178, n17925, n17903, n23167, n19077, n23204, n19106,
    n14016, n14268, n14051, n26255, n18393, n14013, n13920, n13897, n13899,
    n15724, n13900, n21483, n14319, n14047, n19279, n19297, n14332, n14192,
    n14254, n16245, n16564, n14092, n21866, n25467, n14118, n17991, n19049,
    n14830, n14826, n15717, n14125, n13913, n14579, n14104, n14103, n25348,
    n20546, n18464, n18476, n18419, n20672, n13924, n13923, n13925, n13928,
    n20363, n20207, n13929, n20234, n13935, n13937, n13938, n13941, n13942,
    n18421, n20443, n26109, n13943, n13944, n13945, n25863, n13946, n13948,
    n13949, n13952, n13958, n13953, n13957, n20102, n13959, n13961, n13962,
    n13963, n25823, n13964, n13965, n20033, n20029, n20031, n13967, n14895,
    n14921, n23342, n13968, n13969, n22306, n13971, n13972, n13976, n22334,
    n13974, n22219, n13977, n25361, n25088, n13983, n17853, n19811, n19824,
    n19829, n13994, n20127, n13997, n13998, n14006, n14007, n14008, n19344,
    n14009, n14010, n14011, n19492, n14014, n14015, n14019, n14017, n19471,
    n14020, n14022, n14566, n14023, n14024, n14028, n14029, n14547, n18007,
    n23897, n14031, n24158, n23925, n14034, n14036, n14037, n22656, n14039,
    n14040, n22543, n18033, n14348, n19242, n20758, n18363, n20772, n14046,
    n14048, n14049, n14050, n16951, n14057, n20749, n14060, n18337, n14064,
    n14065, n16202, n16223, n14067, n14069, n17456, n14071, n21755, n14767,
    n14076, n14082, n14754, n14086, n14437, n17550, n25051, n14099, n14101,
    n14102, n14110, n14113, n22447, n14114, n14115, n15337, n20931, n14119,
    n20942, n14130, n14131, n14140, n14142, n14143, n14144, n14145, n14147,
    n14149, n18731, n14151, n14416, n14152, n14155, n14160, n18859, n14161,
    n14389, n21371, n14169, n14170, n15444, n17624, n14178, n14179, n14182,
    n17819, n14641, n14186, n19533, n19217, n14191, n19763, n14195, n18208,
    n14197, n18211, n14201, n18399, n14199, n14203, n14204, n14205, n20515,
    n14208, n14209, n14210, n14211, n14217, n18235, n20433, n14222, n14221,
    n26112, n14225, n18333, n20182, n14229, n14230, n19844, n19845, n20076,
    n14231, n19883, n14247, n23726, n14249, n25848, n25934, n20095, n19940,
    n19941, n14855, n20281, n26130, n14259, n14672, n18174, n26161, n15001,
    n14258, n23252, n23124, n19321, n16467, n14696, n14666, n15056, n15070,
    n18022, n22725, n14262, n14263, n23898, n23069, n14264, n17391, n22722,
    n14281, n23336, n15054, n23274, n17886, n14353, n14560, n14554, n22607,
    n14270, n25997, n18039, n19094, n22545, n14272, n14273, n14501, n23250,
    n14274, n14391, n15039, n18810, n20472, n14592, n17352, n14806, n14275,
    n14993, n15652, n15112, n15037, n24970, n14277, n14278, n15302, n15304,
    n14280, n23187, n16108, n23180, n14408, n14285, n14288, n17980, n14290,
    n20818, n14303, n17020, n14304, n14305, n14307, n14308, n19008, n15271,
    n15242, n14309, n14312, n14311, n17799, n14314, n14315, n14317, n24944,
    n14320, n14322, n16778, n16771, n14325, n14326, n18122, n16578, n19174,
    n16956, n17084, n19145, n14333, n14337, n14340, n14341, n14343, n14346,
    n14347, n14349, n14351, n14352, n14354, n14355, n14356, n21072, n21297,
    n14362, n17013, n14364, n17021, n21109, n14367, n14369, n21203, n14370,
    n14371, n23149, n14377, n21492, n15139, n22630, n14396, n14397, n14399,
    n14403, n14404, n14409, n18583, n14413, n18744, n14415, n14421, n14972,
    n14418, n14423, n14422, n14429, n14426, n14427, n25206, n21720, n14435,
    n21774, n14436, n16575, n17532, n14442, n24994, n14447, n21787, n14452,
    n14458, n17703, n14467, n14472, n14473, n14474, n14477, n16322, n14481,
    n16889, n14482, n16871, n14485, n14486, n17280, n14804, n16033, n16029,
    n16131, n16157, n15407, n14504, n22510, n14509, n22548, n23942, n23963,
    n22830, n18069, n16818, n14528, n17134, n14529, n14531, n14532, n19185,
    n19565, n25642, n14533, n14537, n19166, n14536, n14542, n14543, n14544,
    n14545, n14546, n19384, n14552, n14551, n16340, n14555, n14553, n14557,
    n14558, n14559, n14562, n14564, n19423, n14569, n17891, n14576, n16240,
    n16241, n14578, n16544, n14583, n17912, n14585, n23174, n23185, n25661,
    n14589, n14590, n14593, n15138, n14600, n14606, n21250, n14608, n21252,
    n14610, n14612, n17795, n14616, n25042, n25139, n21518, n21559, n14635,
    n14636, n14638, n24996, n21708, n18040, n14647, n14648, n14649, n14652,
    n15077, n15072, n14655, n14656, n22776, n14658, n14664, n14661, n22699,
    n22723, n22676, n22698, n16968, n14669, n14670, n14671, n16969, n14674,
    n14675, n22348, n19101, n14676, n14682, n17994, n14681, n22250, n14686,
    n14687, n14693, n22386, n14698, n14694, n23207, n14695, n23238, n14939,
    n17172, n14707, n14708, n20423, n14716, n14728, n18406, n14739, n20525,
    n14735, n18416, n14737, n14738, n26052, n14741, n14743, n20164, n14744,
    n14747, n14748, n14753, n14761, n21652, n21815, n17044, n14905, n14773,
    n14769, n14771, n14778, n14774, n14775, n17481, n14776, n14780, n22564,
    n14787, n22603, n14789, n14907, n14797, n19510, n19513, n14801, n16520,
    n18161, n26234, n16469, n26306, n25683, n25710, n26253, n14811, n14814,
    n24400, n25279, n25243, n24440, n14824, n24439, n14827, n14829, n20396,
    n20414, n14845, n19042, n14844, n20959, n14856, n14852, n26184, n18927,
    n24424, n14859, n18938, n24504, n14862, n14949, n14981, n15454, n20245,
    n23983, n15866, n25174, n16588, n14864, n24021, n14865, n24012, n14866,
    n14867, n14869, n14870, n14871, n18424, n14872, n14873, n14874, n16051,
    n26315, n23016, n14875, n17017, n14876, n14878, n14879, n14880, n14881,
    n14882, n14883, n14884, n21074, n19441, n19431, n19449, n19465, n15048,
    n15129, n18410, n17040, n15953, n15049, n23737, n26227, n17787, n17634,
    n15352, n14952, n15659, n15999, n26198, n26288, n16326, n15986, n17746,
    n17695, n17768, n16603, n25253, n23222, n15788, n15102, n18062, n22761,
    n15156, n23958, n14926, n15667, n15517, n20354, n20235, n16470, n26280,
    n26137, n16960, n19051, n19029, n17671, n15960, n21352, n21412, n25248,
    n16589, n25509, n22253, n15810, n23796, n23988, n17962, n20416, n25706,
    n20186, n26013, n20501, n20627, n26140, n18307, n16181, n24500, n24475,
    n16779, n17864, n15967, n17345, n23322, n24230, n18060, n15871, n24011,
    n24228, n15867, n14932, n23656, n15338, n15212, n16008, n20552, n25611,
    n16403, n25667, n18487, n18473, n19224, n24511, n21025, n16617, n24916,
    n21828, n25099, n18145, n17006, n23329, n18907, n22847, n23724, n23684,
    n23892, n23944, n17442, n17443, n16313, n25734, n19752, n26027, n26031,
    n26270, n26433, n26398, n17285, n24336, n24508, n24506, n25583, n25559,
    n24875, n25263, n25282, n25553, n25289, n24707, n22164, n23343, n23309,
    n23688, n23722, n22772, n24026, n24019, n24286, n24251, n24113, n24106,
    n17461, n25592, n25368, n14896, n14898, n14897, n14902, n14900, n14899,
    n14901, n14903, n14904, n14906, n14913, n14908, n14915, n14910, n14912,
    n14911, n14914, n23117, n14918, n14917, n14916, n14920, n14919, n14974,
    n14925, n14931, n14928, n14927, n14929, n15911, n14937, n14945, n14940,
    n14943, n14941, n14942, n14944, n18853, n15024, n14948, n14946, n14947,
    n14971, n14951, n14954, n14953, n16809, n14977, n14970, n14965, n14961,
    n14964, n14966, n16176, n14968, n14967, n14989, n16103, n14969, n24122,
    n14973, n14975, n15912, n15925, n24001, n14976, n14979, n14978, n14980,
    n14982, n14986, n14984, n14985, n14987, n15007, n14988, n16078, n15073,
    n17038, n14990, n14992, n14994, n14996, n14995, n14998, n15000, n14999,
    n23316, n15003, n15002, n15004, n15006, n15005, n15074, n15010, n15009,
    n15022, n15018, n15013, n15016, n15015, n15017, n24107, n15019, n24144,
    n15026, n15823, n15025, n15052, n23317, n23221, n15028, n15027, n15032,
    n15030, n15062, n15029, n15031, n18575, n15035, n15038, n15081, n15040,
    n15041, n15044, n15042, n15089, n17949, n15043, n15045, n15047, n15051,
    n15050, n15057, n15053, n23220, n15055, n23225, n15058, n15060, n15059,
    n15068, n15066, n15061, n15063, n15157, n23919, n15064, n15065, n15067,
    n15100, n17207, n15071, n15076, n15075, n15084, n15080, n15079, n15083,
    n15082, n15087, n15086, n15088, n25354, n15099, n15097, n15094, n15090,
    n15093, n15091, n15092, n15095, n15142, n24101, n15096, n15098, n24165,
    n23265, n15130, n23271, n15101, n15103, n23293, n15104, n15128, n15106,
    n15105, n15110, n23867, n15108, n15107, n15109, n15124, n15114, n15116,
    n15115, n15117, n15120, n15118, n15143, n23444, n15119, n15121, n15125,
    n15127, n15126, n15131, n15137, n15135, n15132, n15134, n15136, n15170,
    n15141, n15140, n15176, n15155, n15153, n15144, n15145, n15146, n15149,
    n15147, n15148, n15151, n15150, n24096, n15152, n15154, n15165, n15186,
    n15159, n23842, n15158, n15163, n15669, n15161, n15160, n15162, n23875,
    n15164, n15166, n15171, n15169, n15168, n15172, n15174, n15173, n23337,
    n15177, n15179, n15178, n15207, n15180, n15184, n15182, n23486, n15183,
    n15185, n15195, n15251, n15188, n15187, n15193, n23815, n15191, n15190,
    n15192, n23234, n15194, n15196, n15199, n15198, n15197, n15200, n15204,
    n15202, n15201, n15203, n15205, n15264, n15211, n15209, n15208, n15210,
    n15265, n15238, n25335, n15218, n15216, n15318, n15214, n15213, n24091,
    n15215, n15217, n15231, n15221, n15220, n15229, n15227, n15224, n23805,
    n15225, n15226, n15228, n17396, n15230, n15232, n15236, n15234, n15233,
    n15235, n23237, n15237, n15239, n15241, n15240, n15243, n15247, n15245,
    n15279, n24088, n15246, n15248, n15260, n15250, n15249, n15258, n15256,
    n15253, n23789, n15254, n15255, n15257, n23241, n15259, n15261, n23308,
    n15263, n15262, n22199, n15299, n15266, n15272, n15274, n15276, n15275,
    n15277, n15285, n15283, n15278, n15280, n15281, n24081, n15282, n15284,
    n15295, n15287, n15286, n15293, n15289, n22209, n15291, n15290, n15292,
    n15294, n15296, n22203, n15298, n15297, n22202, n22367, n15300, n15301,
    n15306, n15303, n15305, n15307, n15310, n15312, n15311, n15313, n15314,
    n25320, n15321, n15316, n15317, n15319, n24075, n15320, n15322, n15331,
    n15325, n15324, n15329, n22376, n15327, n15326, n15328, n22207, n15330,
    n15332, n15336, n15334, n15333, n15335, n22371, n15341, n15340, n15342,
    n15343, n15369, n24065, n15349, n15377, n15345, n24069, n15347, n15346,
    n15348, n22257, n15361, n15351, n15350, n15359, n15355, n17414, n22252,
    n15357, n15356, n15358, n15360, n15362, n15365, n15364, n15363, n15366,
    n22247, n15368, n15367, n22248, n15374, n15373, n15405, n25311, n15383,
    n15376, n15378, n15412, n24062, n15381, n15379, n15380, n15382, n15397,
    n15385, n15384, n15395, n15390, n15419, n15389, n15388, n22337, n15393,
    n15392, n15394, n23017, n22754, n15396, n15398, n15401, n15400, n15399,
    n15402, n22333, n15404, n15403, n22332, n15406, n16792, n15440, n15410,
    n21363, n15409, n15411, n15413, n15414, n24056, n15416, n15415, n15417,
    n15429, n15420, n15467, n22756, n15423, n15422, n15427, n15425, n15424,
    n15426, n23035, n22731, n15428, n15433, n15431, n15430, n15432, n15435,
    n22171, n15434, n15437, n15436, n15438, n15439, n15447, n15441, n15449,
    n15465, n16884, n15463, n15453, n15455, n15495, n15461, n15456, n15459,
    n15457, n15458, n15460, n23632, n15462, n15464, n15476, n15466, n15468,
    n22732, n15470, n15469, n15474, n15472, n15471, n15473, n22176, n15475,
    n15477, n15482, n15478, n22399, n18702, n15480, n15479, n22401, n15484,
    n15483, n22400, n22277, n15488, n15487, n15489, n15490, n15516, n16056,
    n15498, n15491, n15493, n15494, n15492, n15496, n15523, n23678, n15497,
    n15499, n15510, n15501, n15502, n22708, n15504, n15503, n15508, n15506,
    n15505, n15507, n15509, n15511, n15515, n15513, n15512, n15514, n22279,
    n15520, n15519, n15521, n15522, n15542, n25296, n15550, n24044, n15525,
    n24041, n15524, n15526, n15536, n22296, n15534, n15529, n15528, n15532,
    n15531, n15533, n22982, n15535, n15537, n15541, n15539, n15538, n15540,
    n22291, n22290, n15545, n18249, n15548, n15547, n25290, n15549, n15552,
    n15551, n23711, n15556, n17077, n15555, n15557, n15567, n22389, n22665,
    n15565, n15561, n15560, n15563, n22660, n15562, n15564, n24289, n15566,
    n15568, n15572, n15570, n15569, n15571, n22387, n15576, n15575, n15578,
    n15583, n17271, n15581, n15580, n15582, n15593, n15584, n22635, n15591,
    n15587, n15586, n15589, n15588, n15590, n24292, n15592, n15597, n15595,
    n15594, n15596, n15598, n22218, n15599, n15601, n15607, n15606, n17294,
    n15608, n15619, n15611, n22612, n15617, n15613, n15612, n15615, n15614,
    n15616, n15618, n15620, n15623, n15622, n15621, n15624, n15626, n15625,
    n15627, n22319, n15632, n15634, n15633, n18271, n15635, n17281, n15636,
    n15639, n15638, n15644, n22590, n15642, n15641, n15643, n15645, n15648,
    n15653, n15649, n22233, n15651, n15656, n15655, n22349, n15657, n18268,
    n15658, n15663, n15666, n15665, n15677, n22356, n15675, n15671, n15670,
    n15673, n15672, n15674, n15676, n15678, n15683, n15681, n15680, n15679,
    n15682, n15684, n22351, n15685, n15687, n15686, n15688, n15691, n15690,
    n15721, n15692, n17718, n15695, n17451, n15694, n15706, n15696, n22550,
    n15698, n15704, n15700, n15699, n15702, n15701, n15703, n15705, n15707,
    n15712, n15709, n15708, n15710, n15711, n15713, n15714, n15715, n15718,
    n15720, n15723, n15722, n15726, n15725, n15748, n15727, n17732, n15729,
    n17331, n15728, n15739, n15731, n22527, n15737, n15733, n15732, n15735,
    n15734, n15736, n15738, n15740, n15743, n15742, n18031, n15741, n15744,
    n22307, n15747, n15745, n15746, n15753, n15752, n15754, n15755, n23159,
    n15756, n15768, n22496, n15759, n15765, n15761, n15760, n15763, n15762,
    n15764, n15767, n15773, n15770, n15769, n15771, n15772, n22265, n15775,
    n15774, n15776, n15779, n15778, n15780, n15804, n15827, n15782, n15786,
    n15783, n15785, n23151, n15787, n15796, n17997, n22474, n15794, n15790,
    n15789, n15792, n15791, n15793, n15795, n15797, n15800, n15799, n15798,
    n15801, n17995, n15803, n15802, n17996, n15833, n15807, n15809, n15808,
    n15837, n23144, n15811, n15822, n15814, n15813, n15820, n15816, n19108,
    n15818, n15817, n15819, n15821, n15915, n15825, n15824, n15826, n15916,
    n19102, n15831, n15829, n15835, n15832, n15834, n15838, n15840, n15839,
    n15841, n15842, n15844, n15846, n15848, n18361, n15847, n15857, n15850,
    n15849, n15855, n15853, n15852, n15854, n15856, n15858, n15864, n15862,
    n15861, n15863, n15921, n15868, n15869, n15877, n15875, n15873, n15872,
    n15874, n15876, n15893, n15879, n15878, n15883, n15881, n15880, n15882,
    n15891, n15885, n15884, n15889, n15887, n15886, n15888, n15890, n15892,
    n15898, n15895, n15894, n15896, n15897, n15899, n15900, n17438, n24117,
    n15902, n17434, n17408, n15903, n15906, n15909, n15908, n15910, n16808,
    n15922, n15913, n23339, n15914, n15919, n15917, n15918, n15920, n15951,
    n23931, n23966, n15924, n15923, n17436, n15949, n15927, n15926, n15928,
    n16972, n15929, n15947, n15932, n23217, n23391, n15935, n15934, n15945,
    n23279, n15938, n15937, n15943, n15941, n22432, n15940, n15942, n15944,
    n15946, n15948, n15950, n15952, n15954, n15956, n17596, n16568, n16565,
    n15964, n15974, n15969, n15971, n15972, n15973, n17011, n15975, n15978,
    n15976, n15977, n15980, n17447, n21339, n15982, n15981, n15985, n15984,
    n16132, n16009, n15997, n15989, n16010, n16012, n15995, n16011, n15993,
    n15994, n15996, n16001, n16007, n16005, n16004, n16006, n16287, n20802,
    n19831, n16016, n16955, n16013, n16015, n16017, n16018, n16020, n16019,
    n16182, n16023, n16022, n16184, n16155, n16026, n16025, n16130, n16028,
    n16145, n16030, n16032, n16035, n16036, n16038, n16040, n16224, n16041,
    n16042, n16250, n16044, n16045, n16276, n16046, n16047, n16323, n16048,
    n16054, n16870, n16055, n16890, n16057, n16059, n18243, n20792, n16070,
    n16324, n16060, n16522, n16062, n16061, n16790, n16891, n16064, n16893,
    n16066, n16065, n20094, n16068, n20796, n20774, n16067, n16069, n16071,
    n16096, n16072, n16075, n16098, n16097, n16077, n16079, n17042, n16081,
    n16080, n16083, n16085, n16084, n17193, n16092, n19964, n16086, n16087,
    n16088, n16090, n16091, n16100, n16099, n16102, n16105, n16104, n16107,
    n16238, n16111, n16112, n16244, n16113, n16116, n16242, n18168, n16129,
    n16119, n16124, n16120, n16123, n16121, n16122, n16125, n25875, n16127,
    n16126, n16128, n17230, n16136, n16147, n19972, n16134, n16133, n16135,
    n18175, n16143, n25893, n16141, n16140, n16142, n18165, n16153, n16148,
    n16149, n25850, n16151, n16150, n16152, n16156, n17218, n16164, n16158,
    n16159, n25811, n16162, n16161, n16163, n25360, n16172, n25337, n16170,
    n16167, n16165, n16166, n16168, n16169, n16171, n16174, n16173, n16180,
    n16178, n16177, n17197, n16179, n16183, n17206, n16188, n16186, n16185,
    n16187, n16189, n16201, n17492, n16190, n16215, n17510, n16191, n17512,
    n17515, n16192, n16195, n16193, n16194, n16197, n16196, n24647, n24631,
    n16199, n16198, n16200, n18182, n16212, n16251, n16205, n16207, n16206,
    n16208, n16225, n25916, n16210, n18183, n16209, n16211, n16213, n16222,
    n16214, n16217, n16216, n16218, n24606, n24576, n16220, n16219, n16221,
    n18190, n16230, n16226, n19984, n16228, n16227, n16229, n16231, n16237,
    n24085, n16233, n16235, n16234, n16236, n16318, n16248, n16246, n16247,
    n18196, n16260, n16252, n16253, n16255, n16256, n19987, n16258, n16257,
    n16259, n16264, n16262, n24110, n16261, n16263, n26311, n17133, n16290,
    n16265, n17106, n16266, n16267, n16268, n16269, n16270, n16274, n16272,
    n16271, n16273, n16285, n16277, n16280, n16278, n16279, n16281, n19989,
    n16283, n16282, n16284, n16289, n20786, n17135, n16288, n26312, n16291,
    n16292, n16293, n16294, n16295, n16296, n17105, n16297, n16298, n16299,
    n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
    n16309, n16310, n16311, n16312, n16315, n16317, n16319, n16321, n16334,
    n16325, n16328, n16327, n16329, n25988, n16330, n16332, n16331, n16333,
    n16336, n16335, n16422, n16342, n20766, n16341, n16349, n16344, n25699,
    n16347, n16463, n18368, n16346, n16348, n16351, n16350, n16353, n16352,
    n16358, n16354, n26151, n16356, n16355, n16357, n16360, n16359, n16362,
    n16361, n16368, n16364, n20485, n16366, n16365, n16367, n16370, n16369,
    n16372, n16371, n16380, n16375, n20508, n16378, n16377, n16379, n16382,
    n16381, n16384, n16383, n16390, n16385, n26175, n16388, n16387, n16389,
    n16392, n16391, n16394, n16393, n16399, n16395, n26067, n16397, n16396,
    n16398, n16401, n16400, n16405, n16402, n26094, n16404, n16409, n16407,
    n16406, n16408, n16411, n16410, n16413, n16412, n16419, n16415, n20463,
    n16417, n16416, n16418, n16421, n16420, n16424, n18380, n16423, n16430,
    n16426, n26141, n16428, n16427, n16429, n19134, n26165, n16432, n16431,
    n16434, n16433, n16438, n16436, n16435, n16437, n16440, n16439, n16442,
    n16441, n16447, n16445, n16443, n16444, n16446, n16449, n16448, n16451,
    n16450, n16457, n16453, n26213, n16455, n16454, n16456, n16459, n16458,
    n16462, n16461, n16465, n16464, n16466, n16468, n16475, n16472, n26101,
    n16474, n16479, n16477, n16476, n16478, n16481, n16480, n16482, n16488,
    n16486, n16485, n16487, n16490, n16489, n16492, n20444, n16494, n16493,
    n16498, n16496, n16495, n16497, n19646, n16500, n16499, n16502, n20425,
    n16508, n16504, n16503, n16506, n16505, n16507, n19795, n16510, n16509,
    n16512, n16514, n16513, n16516, n16515, n16518, n16517, n16521, n18212,
    n16527, n16523, n19993, n16525, n16524, n16526, n16528, n16530, n20407,
    n16536, n16532, n16531, n16534, n16533, n16535, n19771, n16538, n16537,
    n16541, n16542, n16545, n16547, n16549, n16551, n16550, n16553, n16552,
    n16555, n16554, n16557, n16556, n16559, n16558, n16561, n16560, n16563,
    n16562, n16567, n16566, n16571, n16570, n16576, n16573, n16577, n16579,
    n16582, n16581, n16584, n16586, n16781, n16585, n16595, n16593, n16742,
    n16714, n16622, n25033, n16591, n16592, n16594, n16597, n16596, n16599,
    n16598, n16601, n16600, n16608, n16602, n16701, n16604, n16605, n16606,
    n21723, n16607, n21734, n16610, n16609, n16612, n16611, n16613, n16614,
    n16616, n16619, n16618, n16621, n16620, n16630, n16628, n17780, n16624,
    n16623, n16625, n25009, n16626, n16627, n16629, n16632, n16631, n16634,
    n16633, n16638, n21831, n16636, n16635, n16637, n16640, n16639, n16644,
    n16642, n16641, n16643, n21745, n16646, n16645, n16650, n16648, n16647,
    n16649, n16652, n16651, n16654, n16653, n16658, n24390, n24395, n16656,
    n16655, n16657, n16660, n16659, n20824, n16663, n16662, n21805, n16665,
    n16664, n16669, n16667, n16666, n16668, n16671, n16670, n16673, n16672,
    n16681, n16679, n16675, n24941, n16677, n16678, n16680, n16683, n16682,
    n16685, n16684, n16690, n16688, n24964, n16687, n16689, n16692, n16691,
    n16694, n16693, n16698, n16696, n25188, n16695, n16697, n16700, n16699,
    n24474, n16703, n16702, n16707, n16705, n16704, n16706, n16709, n16708,
    n16711, n16710, n16720, n16718, n16713, n16712, n16715, n25059, n16716,
    n16717, n16719, n16722, n16721, n16724, n16723, n16730, n16728, n25073,
    n16726, n16727, n16729, n16732, n16731, n16733, n25106, n16735, n16734,
    n16736, n16738, n16737, n16740, n16739, n16747, n16745, n16741, n16743,
    n24429, n25160, n16744, n16746, n25183, n16749, n16748, n16750, n21778,
    n16753, n16752, n16757, n16755, n16754, n16756, n16759, n16758, n16761,
    n16760, n16763, n16762, n16765, n16764, n16767, n16766, n16769, n16768,
    n16773, n16770, n16772, n16775, n16774, n16776, n16785, n16783, n16782,
    n16784, n16787, n16786, n16788, n16796, n16791, n19997, n26036, n16794,
    n16793, n16795, n16797, n16799, n20381, n16805, n16801, n16800, n16803,
    n20391, n16802, n16804, n16807, n16806, n23219, n18905, n18908, n16817,
    n16810, n16815, n16811, n16831, n23409, n23364, n23363, n23390, n16813,
    n23366, n16812, n23401, n23400, n23399, n23380, n16814, n23410, n16820,
    n16816, n23356, n16819, n23720, n16829, n16821, n23501, n16822, n23372,
    n23371, n23374, n16824, n23382, n23381, n16826, n16825, n23414, n23415,
    n16827, n16828, n16830, n16833, n23416, n16832, n16841, n16837, n16921,
    n16920, n16840, n16919, n16932, n19587, n16842, n16848, n16844, n16843,
    n16846, n20366, n16845, n16847, n16850, n16849, n19583, n16853, n20342,
    n16859, n16855, n16854, n16857, n16856, n16858, n19602, n16861, n16860,
    n16863, n16862, n16865, n16864, n16867, n16866, n16869, n16868, n18228,
    n16877, n16873, n19999, n16875, n16874, n16876, n16883, n16879, n24863,
    n24842, n16881, n17625, n16880, n16882, n16888, n16886, n16885, n16887,
    n18236, n16898, n16892, n16894, n20059, n16896, n18238, n16895, n16897,
    n16900, n20321, n16906, n16902, n16901, n16904, n16903, n16905, n16908,
    n16907, n16938, n16909, n16910, n20273, n16916, n16912, n16911, n16914,
    n16913, n16915, n19692, n16918, n16917, n16922, n16925, n16927, n16931,
    n16936, n16934, n16935, n17256, n16940, n20299, n16947, n16943, n16942,
    n16945, n16944, n16946, n16949, n16948, n16950, n16952, n16953, n18248,
    n16965, n16957, n16959, n16961, n20106, n16963, n16962, n16964, n16967,
    n16966, n16971, n23389, n16970, n16974, n23319, n16973, n16975, n16976,
    n16982, n16980, n16978, n16977, n16979, n16981, n16998, n16984, n16983,
    n16988, n16986, n16985, n16987, n16996, n16990, n16989, n16994, n16992,
    n16991, n16993, n16995, n16997, n17003, n17000, n16999, n17001, n17002,
    n17004, n17005, n17862, n25374, n17007, n25370, n17009, n17010, n17069,
    n17012, n17030, n21030, n17016, n17018, n17019, n17024, n17026, n17027,
    n25441, n17028, n17031, n17032, n17035, n17034, n17041, n17043, n24454,
    n17045, n17047, n17048, n17057, n21401, n17050, n25092, n17051, n17498,
    n17055, n17052, n24484, n17053, n17054, n17056, n17068, n17063, n17061,
    n17860, n17060, n17062, n17066, n17290, n17064, n17065, n24487, n17067,
    n17074, n21417, n25091, n17072, n17070, n17073, n25291, n17075, n17078,
    n17079, n18256, n17090, n17080, n17083, n17081, n17082, n17086, n17085,
    n17137, n20119, n17088, n18257, n17087, n17089, n17092, n20246, n17098,
    n17094, n17093, n17096, n17095, n17097, n20266, n17100, n17099, n26310,
    n17103, n17102, n17104, n17130, n17112, n17110, n17108, n17107, n17109,
    n17111, n17128, n17114, n17113, n17118, n17116, n17115, n17117, n17126,
    n17120, n17119, n17124, n17122, n17121, n17123, n17125, n17127, n17129,
    n17131, n17132, n17155, n18449, n17136, n17171, n18467, n17139, n19522,
    n17190, n17141, n17142, n17145, n17144, n17146, n19301, n17148, n17151,
    n17149, n17150, n17153, n18454, n18468, n17154, n17164, n17156, n18470,
    n17157, n17159, n17158, n17161, n17160, n18457, n18465, n17162, n17163,
    n17166, n18453, n17165, n17167, n17169, n19834, n19524, n17168, n17252,
    n17170, n17238, n17173, n17176, n17175, n17181, n17182, n20000, n18191,
    n18258, n18387, n17183, n25728, n17250, n25819, n17248, n17186, n17184,
    n17185, n17187, n25732, n17188, n17192, n17189, n17191, n17195, n17194,
    n26277, n17200, n17199, n17203, n17201, n17202, n17204, n25659, n25712,
    n17212, n17209, n17208, n17210, n17211, n17214, n17217, n17215, n18158,
    n17216, n25711, n25714, n25629, n17224, n17220, n17219, n17222, n17221,
    n17225, n25630, n17223, n17227, n17226, n17229, n17228, n17232, n17231,
    n17233, n19129, n17234, n17235, n17237, n17246, n17239, n25724, n17244,
    n17240, n17242, n26278, n20673, n17241, n17243, n17245, n17247, n17249,
    n17251, n17253, n17255, n17258, n17309, n17264, n17262, n17261, n17263,
    n17268, n17266, n17665, n17265, n17267, n17269, n17272, n18267, n17276,
    n17274, n17273, n17275, n17680, n17278, n17692, n17277, n17279, n17282,
    n17706, n17457, n17283, n17284, n17455, n18263, n17288, n19305, n19526,
    n17286, n17287, n17292, n25365, n17289, n17291, n17293, n17298, n17296,
    n17295, n17297, n17301, n17304, n17303, n18270, n17308, n17306, n17305,
    n17307, n17311, n17313, n17320, n17314, n17882, n17319, n17318, n17317,
    n17323, n17321, n17322, n17329, n17328, n17326, n18293, n17325, n17327,
    n17335, n17330, n17333, n17332, n17334, n17339, n17337, n17336, n17338,
    n17340, n17344, n17342, n17341, n17343, n17705, n17347, n17351, n17349,
    n17348, n17350, n18868, n17354, n17353, n17386, n18869, n17385, n17355,
    n17356, n17358, n18871, n18866, n23880, n17360, n18872, n17361, n23828,
    n17363, n17364, n17367, n17368, n17395, n23776, n17369, n17372, n17370,
    n17371, n17373, n17374, n17464, n17376, n18885, n17413, n23914, n17381,
    n24014, n17379, n22789, n17378, n17380, n17407, n17383, n23950, n17387,
    n17388, n17390, n17392, n17393, n17394, n17398, n17397, n23739, n22782,
    n22784, n18883, n22783, n17401, n17402, n18882, n17480, n17405, n17404,
    n17403, n17406, n17433, n17409, n22436, n17412, n17410, n17411, n17422,
    n17426, n23970, n17420, n24155, n24242, n17427, n17418, n23980, n17416,
    n17415, n17417, n17419, n17421, n17425, n18909, n17424, n24220, n17431,
    n24216, n17429, n17428, n17430, n17432, n17444, n17435, n17437, n17439,
    n17441, n17440, n17446, n17445, n17450, n21403, n21457, n18292, n17448,
    n17449, n17454, n17452, n17453, n18289, n18285, n17459, n17458, n17460,
    n17462, n22750, n17465, n18006, n23031, n22752, n17479, n23032, n17477,
    n23033, n17475, n22707, n17471, n17469, n24022, n17467, n17468, n17470,
    n17473, n22755, n22713, n17472, n17474, n17476, n17478, n17483, n23044,
    n17482, n17484, n25244, n21061, n17485, n17495, n17488, n17491, n17489,
    n17490, n17493, n24586, n17496, n17500, n17499, n25175, n17501, n17507,
    n17505, n17504, n17506, n25410, n25137, n25111, n25136, n17509, n17518,
    n17511, n17514, n17513, n17516, n24627, n17517, n17519, n17792, n25142,
    n17530, n24482, n25119, n17528, n17523, n17522, n17524, n17526, n17527,
    n17529, n17531, n17538, n17536, n17534, n24668, n17535, n17537, n25090,
    n17793, n17539, n17547, n17540, n17545, n17541, n17542, n17543, n24687,
    n17544, n17546, n17548, n17549, n17561, n25336, n17559, n17551, n17556,
    n17552, n17555, n17553, n17554, n17557, n17558, n17560, n17800, n17562,
    n17563, n17574, n17566, n17568, n17570, n17567, n17572, n17571, n17586,
    n24725, n17573, n17575, n24971, n17576, n17577, n17583, n17581, n17579,
    n24751, n17580, n17582, n24434, n17584, n17585, n17593, n17587, n17588,
    n24765, n17591, n17590, n17592, n17805, n17806, n24349, n17594, n17595,
    n17601, n17598, n17605, n17599, n24779, n17600, n17602, n21415, n17604,
    n21414, n17610, n17608, n17606, n24817, n17607, n17609, n21431, n21430,
    n17612, n17619, n17615, n17614, n17616, n17617, n24832, n17618, n17620,
    n24462, n17622, n17623, n17627, n17626, n21035, n21760, n17628, n21804,
    n17629, n17630, n17639, n17633, n17636, n17635, n17637, n24886, n17638,
    n17640, n21791, n17642, n17644, n17643, n21732, n17649, n17646, n17645,
    n17655, n17647, n24903, n17648, n17650, n21759, n17652, n17654, n17653,
    n21705, n17656, n24928, n17659, n17658, n17660, n17661, n17663, n17662,
    n17667, n17666, n17668, n17670, n17669, n17676, n17672, n21695, n17674,
    n17673, n17675, n21709, n17677, n17681, n17684, n17683, n17690, n17686,
    n21666, n17688, n17687, n17689, n17693, n17696, n21642, n17698, n17697,
    n17702, n17700, n17699, n17701, n20948, n21411, n17707, n17710, n17709,
    n17716, n17712, n21621, n17714, n17713, n17715, n17717, n17720, n17719,
    n17721, n17723, n21599, n17725, n17724, n17729, n17727, n17726, n17728,
    n17730, n17731, n17733, n17736, n17735, n17742, n17738, n21572, n17740,
    n17739, n17741, n21558, n21587, n17743, n22166, n17744, n17747, n21545,
    n17749, n17748, n17753, n17751, n17750, n17752, n17754, n22158, n17755,
    n17757, n17756, n17763, n17759, n21522, n17761, n17760, n17762, n21410,
    n21508, n17764, n22151, n17765, n17767, n17766, n17772, n17777, n20807,
    n17770, n17769, n17771, n17773, n17775, n22145, n17774, n17776, n17778,
    n18126, n17779, n17786, n17782, n17781, n17784, n17783, n17785, n18084,
    n18113, n17789, n21394, n17788, n17848, n25218, n17791, n25040, n25043,
    n17794, n17796, n17797, n25052, n17798, n25029, n17801, n17802, n17803,
    n17804, n21880, n17807, n17808, n17809, n17810, n17812, n17813, n17815,
    n21789, n21758, n17817, n17818, n17820, n21678, n17821, n17822, n20867,
    n17823, n17824, n21617, n17825, n21561, n17826, n21943, n17827, n17829,
    n17830, n21517, n17831, n17832, n17833, n18118, n17835, n17849, n17836,
    n17846, n17842, n17838, n17837, n17840, n17839, n17841, n25586, n21340,
    n17844, n17843, n17845, n17847, n21486, n17858, n21722, n17852, n25156,
    n17850, n17851, n21829, n21802, n21771, n21620, n21497, n17854, n17855,
    n25505, n17856, n17857, n17859, n18147, n17865, n17861, n18109, n17867,
    n17866, n17871, n18088, n17869, n17868, n17870, n21495, n17877, n21496,
    n17875, n17874, n17876, n17878, n17880, n17879, n23532, n17883, n17884,
    n17885, n17895, n17887, n17889, n17888, n17890, n17900, n17892, n17893,
    n17896, n17898, n17902, n17901, n23574, n17904, n17906, n17907, n17916,
    n17908, n17910, n17909, n17911, n17921, n17913, n17914, n17917, n17919,
    n17923, n17920, n17922, n23184, n23606, n17926, n17928, n17929, n17931,
    n17930, n17932, n17935, n17933, n17936, n17937, n17938, n17939, n23645,
    n17943, n17941, n17946, n17947, n17953, n17951, n17950, n17952, n17957,
    n17956, n17958, n17959, n17973, n17960, n17964, n17963, n17965, n17979,
    n17966, n17968, n17967, n17969, n17970, n17972, n23118, n17971, n22730,
    n17976, n17978, n19225, n17977, n23125, n17981, n17983, n17989, n17985,
    n17984, n17987, n17986, n18510, n24330, n18910, n17988, n19086, n22811,
    n17990, n23060, n17993, n17992, n18005, n18003, n18001, n17999, n17998,
    n18000, n18002, n18004, n18864, n22953, n22624, n18008, n18009, n18010,
    n18044, n18011, n18012, n18013, n22680, n18014, n22706, n18015, n22655,
    n18016, n18048, n18017, n22629, n18019, n18052, n18024, n18023, n22585,
    n18025, n18027, n18028, n18029, n18056, n18030, n22514, n18032, n22509,
    n18034, n18035, n18036, n18037, n18038, n18066, n22771, n18042, n18043,
    n18891, n18892, n18047, n18049, n18051, n18053, n18054, n18055, n18057,
    n18058, n18061, n18065, n18064, n18063, n18068, n18067, n18079, n18077,
    n18136, n18075, n18073, n18071, n18072, n18074, n18076, n18078, n18087,
    n18082, n22140, n18081, n21447, n18083, n18104, n18085, n18086, n18102,
    n18123, n18089, n18090, n18100, n18098, n18091, n18092, n21463, n18094,
    n18093, n18096, n18095, n25589, n18097, n18099, n18101, n18103, n18154,
    n18107, n18108, n18110, n18112, n18111, n18134, n18117, n18114, n18116,
    n18115, n18120, n18119, n18124, n18132, n18151, n21803, n18130, n21459,
    n25189, n18128, n18127, n18129, n18131, n18133, n18140, n18138, n18137,
    n18139, n18142, n18143, n25488, n18149, n18148, n25477, n22038, n18153,
    n18152, n18156, n18155, n18157, n18402, n26232, n19322, n19274, n25707,
    n19329, n25626, n18160, n25624, n19340, n18162, n25723, n18164, n18163,
    n18167, n18166, n19345, n26181, n26183, n18227, n18173, n18171, n18170,
    n18172, n18405, n26160, n19357, n26127, n18180, n18178, n18177, n18179,
    n26367, n26106, n25597, n18181, n18187, n18185, n18184, n18186, n19360,
    n26375, n19371, n19363, n18188, n18195, n18193, n18192, n18194, n18200,
    n18198, n18197, n18199, n18201, n18207, n18205, n18204, n18206, n20681,
    n18413, n18414, n18209, n18210, n20507, n18418, n18417, n18214, n18213,
    n18215, n18217, n20484, n18218, n18221, n18220, n18222, n18226, n18224,
    n18225, n18232, n18230, n18229, n18231, n18233, n19415, n18234, n18237,
    n18242, n18240, n18239, n18241, n20424, n19287, n19424, n18245, n18244,
    n18246, n20406, n18251, n18250, n18252, n19430, n18254, n18260, n18259,
    n18261, n19453, n18262, n20280, n18265, n18264, n18266, n18280, n18275,
    n18269, n20306, n18272, n18274, n20283, n18276, n20298, n18278, n18277,
    n20254, n18284, n18282, n18281, n20253, n18286, n18287, n19568, n19466,
    n20287, n19467, n20263, n20228, n18290, n18295, n18294, n18308, n18296,
    n18298, n18299, n18300, n20210, n18303, n18305, n18304, n20229, n18319,
    n18318, n20793, n20795, n18309, n20221, n18316, n18312, n18311, n18314,
    n18313, n18315, n19480, n18317, n18320, n18334, n20785, n20787, n20198,
    n18330, n18325, n18324, n18328, n20193, n18327, n18329, n18331, n18332,
    n18336, n18347, n20780, n18338, n20175, n18346, n18342, n18341, n18344,
    n18343, n18345, n18350, n18349, n18360, n18352, n18353, n18356, n18358,
    n18357, n18359, n18362, n19223, n20765, n20767, n18364, n18367, n19231,
    n18372, n18370, n18369, n18371, n19499, n18374, n18373, n19252, n18375,
    n18376, n18377, n18378, n18391, n18379, n18384, n18382, n18381, n18383,
    n19509, n19520, n19950, n18386, n20130, n18389, n18388, n18390, n18392,
    n18396, n18394, n18395, n18488, n18397, n18447, n19309, n18398, n26248,
    n18400, n18401, n18403, n18404, n26074, n26111, n26075, n19373, n18407,
    n18412, n18409, n26107, n18408, n19372, n19388, n19379, n18415, n20493,
    n19397, n19401, n19400, n19405, n20442, n19417, n18420, n20435, n18422,
    n19442, n18423, n18426, n18427, n18428, n19459, n18429, n19456, n20315,
    n20258, n20260, n19462, n18430, n19461, n18433, n20259, n18432, n18434,
    n18435, n19271, n19473, n19270, n19472, n18438, n18439, n18440, n18441,
    n18442, n18445, n18444, n18452, n20684, n18446, n18451, n18450, n18481,
    n18480, n18461, n18479, n18456, n18458, n18459, n18460, n18462, n18463,
    n18466, n18472, n18469, n18471, n18474, n18475, n18478, n18485, n18483,
    n18484, n18486, n18489, n18491, n18490, n18493, n20131, n18494, n26249,
    n20388, n18496, n18499, n18498, n18500, n18506, n18502, n18511, n18507,
    n18503, n18505, n18504, n18509, n18508, n18522, n18521, n18849, n18735,
    n18520, n18517, n18516, n18514, n18513, n18515, n24327, n18518, n18519,
    n18845, n18526, n18523, n18524, n18525, n18844, n18532, n18528, n24323,
    n18527, n18836, n18530, n18529, n18835, n18531, n18533, n18842, n18534,
    n18763, n18536, n18762, n18761, n18539, n18538, n18757, n18541, n18540,
    n18756, n18755, n18543, n18542, n18559, n18552, n18546, n18548, n18550,
    n18558, n18554, n18553, n18556, n18555, n18557, n18561, n18560, n18562,
    n18569, n18566, n18565, n18564, n18568, n18567, n18571, n18570, n18572,
    n18574, n18573, n18581, n18576, n18578, n18577, n18593, n18580, n18579,
    n18592, n18586, n18582, n18584, n18585, n18587, n18589, n18588, n18605,
    n18591, n18590, n18604, n18597, n18595, n18594, n18596, n18598, n18611,
    n18601, n18600, n18616, n18603, n18602, n18615, n18609, n18607, n18606,
    n18608, n18610, n18612, n18614, n18613, n18625, n18620, n18618, n18617,
    n18619, n18622, n18621, n18637, n18624, n18623, n18636, n18630, n18628,
    n18629, n18631, n18633, n18632, n18644, n18635, n18634, n18643, n18641,
    n18639, n18638, n18640, n18642, n18646, n18645, n18653, n18648, n18647,
    n18660, n18651, n18650, n18659, n18652, n18654, n18656, n18655, n18672,
    n18658, n18657, n18671, n18664, n18662, n18661, n18663, n18665, n18668,
    n18667, n18682, n18670, n18669, n18681, n18676, n18674, n18673, n18675,
    n18678, n18677, n18689, n18680, n18679, n18688, n18686, n18684, n18683,
    n18685, n18687, n18691, n18690, n18692, n18694, n18693, n18699, n18696,
    n18695, n18698, n18697, n18701, n18700, n18704, n18703, n18709, n18706,
    n18705, n18708, n18707, n18711, n18710, n18712, n18714, n18713, n18720,
    n18716, n18715, n18719, n18717, n18724, n18722, n18721, n18723, n18726,
    n18725, n18730, n18728, n18727, n18729, n18732, n18734, n18733, n18740,
    n18737, n18736, n18739, n18738, n18742, n18741, n18743, n18746, n18745,
    n18751, n18748, n18747, n18750, n18749, n18753, n18752, n18754, n18759,
    n18758, n18760, n18765, n18764, n18766, n18768, n18767, n18774, n18770,
    n18769, n18773, n18771, n18778, n18776, n18775, n18777, n18788, n18781,
    n18780, n18789, n18787, n18783, n18782, n18797, n18785, n18784, n18796,
    n18786, n18791, n18790, n18795, n18793, n18792, n18794, n18799, n18798,
    n18800, n18802, n18801, n18809, n18804, n18803, n18815, n18807, n18806,
    n18814, n18808, n18812, n18811, n18813, n18816, n18818, n18817, n18824,
    n18820, n18819, n18823, n18821, n18828, n18826, n18825, n18827, n18834,
    n18831, n18830, n18838, n18833, n18832, n18837, n18840, n18839, n18841,
    n18847, n18846, n18848, n18851, n18850, n18852, n18855, n18857, n18858,
    n18862, n19081, n19098, n18898, n22521, n18867, n23910, n18870, n23990,
    n18875, n23885, n18873, n24121, n18874, n18878, n18879, n18880, n18884,
    n22786, n18886, n18888, n18889, n18890, n22694, n18894, n18895, n18897,
    n18903, n18906, n18913, n18911, n18912, n18914, n18917, n18918, n18919,
    n18921, n18922, n24366, n18924, n18923, n18925, n18926, n24422, n24423,
    n24410, n18928, n18929, n18933, n18931, n18930, n18932, n24411, n18935,
    n24505, n18934, n18940, n18941, n18942, n18944, n18943, n24378, n24379,
    n18945, n18946, n18950, n18948, n18947, n18949, n24438, n18951, n18952,
    n24353, n18953, n18954, n18955, n18956, n20974, n18959, n18958, n18957,
    n20973, n18960, n18961, n24401, n18963, n18962, n24402, n18965, n18964,
    n24467, n24466, n18966, n18967, n18981, n18969, n18968, n18970, n20899,
    n20896, n18977, n18971, n20903, n18973, n18974, n20819, n18972, n18984,
    n18980, n18976, n18975, n21017, n18979, n20894, n18978, n20901, n18982,
    n18983, n20918, n18985, n18986, n18990, n18988, n18987, n18989, n20917,
    n18993, n18992, n20987, n18991, n18994, n18995, n18996, n20851, n18998,
    n18997, n20850, n18999, n19000, n20944, n19002, n19001, n20943, n19005,
    n19004, n19006, n20961, n19010, n19007, n19011, n20834, n20836, n19014,
    n19012, n20835, n19015, n19016, n20930, n19017, n19018, n19021, n19019,
    n20879, n19020, n19022, n19023, n19024, n19026, n19025, n19027, n21002,
    n19028, n19031, n19030, n20805, n19032, n19034, n19043, n19035, n19037,
    n19036, n19038, n19041, n19039, n19040, n19046, n19044, n19045, n19047,
    n19048, n19059, n19050, n19055, n19053, n19052, n19054, n19057, n19056,
    n19058, n19063, n19062, n19067, n23685, n19068, n19066, n23197, n19070,
    n19069, n19072, n19071, n19075, n19073, n19074, n19076, n19080, n19079,
    n19082, n19083, n19091, n19089, n22435, n19087, n19088, n19090, n19093,
    n19097, n19096, n19099, n19104, n19103, n19105, n19107, n19118, n19116,
    n19114, n22463, n19112, n19110, n19109, n19111, n19113, n19115, n19117,
    n19119, n19668, n19120, n19652, n19792, n19121, n19161, n19122, n19128,
    n19123, n19124, n19549, n19737, n19125, n19157, n19126, n19156, n19127,
    n19644, n25672, n19131, n19133, n19132, n25671, n19136, n25731, n19137,
    n25600, n19140, n19139, n19141, n19142, n25643, n19143, n19144, n19146,
    n19149, n19147, n19148, n19704, n19150, n25615, n19151, n19152, n25695,
    n19153, n19154, n19155, n19614, n19546, n19158, n19643, n19159, n19664,
    n19164, n19670, n19162, n19163, n19165, n19167, n19168, n19169, n19765,
    n19170, n19579, n19171, n19719, n19172, n19596, n19173, n19175, n19563,
    n19179, n19183, n19180, n19181, n19688, n19182, n19184, n19186, n19189,
    n19187, n19188, n19629, n19190, n19191, n19194, n19192, n19193, n19195,
    n19201, n19198, n19196, n19197, n19532, n19215, n19199, n19203, n19200,
    n19202, n19214, n19212, n19210, n25654, n19204, n19208, n20147, n19206,
    n19205, n19207, n19209, n19211, n19213, n25684, n19216, n19218, n19220,
    n19221, n19227, n19226, n19240, n20760, n19229, n19238, n19232, n19236,
    n19234, n19233, n19235, n19237, n19255, n19239, n19246, n19241, n19244,
    n19243, n19245, n19516, n19247, n19249, n19256, n19250, n19251, n19263,
    n19511, n19265, n19254, n19261, n19258, n19259, n19260, n19262, n19264,
    n19266, n19267, n19268, n19514, n19299, n20292, n20362, n20477, n20500,
    n19272, n19278, n19275, n26305, n19276, n19277, n19280, n19281, n26081,
    n26078, n19282, n19283, n19284, n19285, n19286, n19289, n19290, n19291,
    n19292, n19293, n19294, n19296, n19298, n19302, n19303, n19307, n19311,
    n19310, n19320, n19318, n19316, n19317, n19319, n19326, n19324, n19323,
    n19325, n19328, n19332, n19330, n19331, n19337, n19336, n19339, n19343,
    n19341, n19342, n19355, n19348, n19347, n19353, n19350, n19349, n19356,
    n19351, n19352, n19354, n19358, n19359, n19362, n19361, n19370, n19369,
    n19365, n19367, n19366, n19368, n19375, n19374, n19376, n20674, n19396,
    n25691, n19377, n19378, n19382, n19380, n19381, n19385, n19383, n19395,
    n19394, n19386, n19387, n19390, n19389, n19392, n19393, n19399, n19398,
    n19403, n19402, n19404, n19409, n19407, n19408, n19410, n20640, n19412,
    n19411, n19425, n19414, n19421, n19416, n19419, n19418, n19420, n19422,
    n19426, n19429, n19428, n19433, n19440, n19432, n19437, n19443, n19434,
    n19435, n19436, n19439, n19438, n20624, n19445, n19444, n19448, n19447,
    n19451, n19454, n20609, n19455, n19458, n19457, n19464, n19463, n19469,
    n19468, n19470, n19477, n19475, n19474, n19476, n19478, n19482, n19481,
    n19483, n19486, n19484, n19485, n19487, n19490, n19488, n19489, n19491,
    n20155, n19498, n19496, n19495, n19497, n19500, n19508, n19502, n19506,
    n19504, n19505, n19507, n19512, n19515, n19518, n19517, n19519, n19521,
    n19832, n19523, n19525, n19529, n19527, n19528, n19530, n19531, n19534,
    n19544, n19542, n19538, n19536, n19535, n19537, n19540, n19539, n19541,
    n19543, n19548, n19550, n19551, n19561, n19559, n19557, n19553, n26035,
    n19555, n19554, n19556, n19558, n19560, n19562, n19685, n19564, n19566,
    n19684, n19567, n19578, n19576, n19572, n19570, n19569, n19571, n19574,
    n19573, n19575, n19577, n19580, n19582, n19593, n20616, n19591, n19586,
    n19584, n20120, n19585, n19589, n20359, n19588, n19590, n19592, n19595,
    n19600, n19598, n19599, n19601, n19612, n19610, n19606, n19604, n19603,
    n19605, n19608, n19607, n19609, n19611, n19736, n19613, n19618, n19616,
    n19615, n19617, n19619, n19628, n19626, n19624, n19620, n25990, n19622,
    n19621, n19623, n19625, n19627, n19631, n19642, n20568, n19640, n19632,
    n19636, n19634, n19633, n19635, n19638, n19637, n19639, n19641, n19645,
    n19647, n19665, n19648, n19649, n19793, n19651, n19650, n19653, n19654,
    n19663, n19661, n19659, n19655, n20022, n19657, n19656, n19658, n19660,
    n19662, n19667, n19669, n19672, n19671, n19673, n19683, n19681, n19679,
    n19675, n20050, n19677, n19676, n19678, n19680, n19682, n19687, n19686,
    n19689, n19690, n19702, n19700, n19698, n19691, n19696, n19694, n19693,
    n19695, n19697, n19699, n19701, n19717, n19715, n19713, n19705, n19707,
    n19711, n25924, n19709, n19710, n19712, n19714, n19716, n19718, n19723,
    n19720, n19722, n19724, n19734, n19732, n19726, n19725, n19728, n19727,
    n19730, n19729, n19731, n19733, n19739, n19738, n19740, n19749, n19747,
    n19745, n19741, n26016, n19743, n19742, n19744, n19746, n19748, n19751,
    n19762, n19760, n19756, n19754, n19753, n19755, n19758, n19757, n19759,
    n19761, n19764, n19769, n19767, n19768, n19770, n19780, n19778, n19774,
    n19772, n20086, n19773, n19776, n19775, n19777, n19779, n19791, n19789,
    n19787, n19783, n19782, n19785, n19784, n19786, n19788, n19790, n19794,
    n19804, n19802, n19800, n19796, n19956, n19798, n19797, n19799, n19801,
    n19803, n19805, n25742, n19807, n25778, n19808, n19970, n19810, n25820,
    n25832, n19812, n19974, n19814, n25859, n19815, n19979, n19817, n25903,
    n19818, n25923, n19820, n25942, n25955, n19821, n25966, n19823, n25986,
    n19825, n25985, n19826, n26017, n19828, n26026, n19830, n19837, n19833,
    n19955, n19836, n19953, n20002, n20078, n25741, n19963, n19839, n19838,
    n19841, n19885, n19843, n26300, n19842, n25751, n25750, n25789, n19849,
    n19846, n19848, n19850, n19853, n19851, n19852, n25790, n19854, n25807,
    n19856, n19855, n19857, n19860, n19858, n19859, n25806, n25809, n25829,
    n19862, n26216, n19861, n19863, n19866, n19864, n19865, n25830, n19867,
    n19870, n19869, n19871, n25846, n19873, n26178, n19872, n19874, n25845,
    n19876, n26155, n19875, n19877, n25870, n19878, n19880, n19879, n19882,
    n19881, n25869, n25889, n19887, n19884, n19886, n19888, n19891, n19889,
    n19890, n25888, n25891, n25913, n19894, n19892, n19893, n19896, n19895,
    n19899, n19897, n19898, n25914, n19900, n19901, n19903, n19902, n19904,
    n25931, n19906, n26093, n19905, n19907, n25930, n19909, n26066, n19908,
    n19910, n19913, n19911, n19912, n25948, n19916, n19914, n19915, n19917,
    n25973, n19920, n19918, n19919, n19921, n19923, n20504, n25982, n19922,
    n25996, n19925, n19924, n19926, n19927, n19929, n26007, n19928, n19930,
    n26011, n19931, n19932, n26029, n19934, n19933, n26042, n19937, n19935,
    n19936, n19938, n19939, n20010, n20030, n19942, n19945, n19943, n19944,
    n19946, n19948, n19949, n19961, n19952, n19951, n25894, n26037, n19959,
    n19954, n26033, n19957, n19958, n19960, n19962, n20005, n25746, n19965,
    n19966, n25782, n19969, n19968, n25822, n19973, n19976, n25862, n19978,
    n19982, n19981, n25907, n25906, n19983, n19986, n25946, n19988, n19991,
    n19992, n26008, n19996, n19995, n19998, n20003, n20001, n20004, n20038,
    n20008, n20009, n20028, n20013, n20011, n20012, n20014, n20046, n20015,
    n20017, n20016, n20018, n20045, n20019, n20020, n20026, n20021, n20024,
    n20023, n20025, n20027, n20037, n20032, n20058, n20057, n20035, n20036,
    n20040, n20041, n20056, n20044, n20042, n20043, n20071, n20069, n20047,
    n20070, n20048, n20054, n20049, n20052, n20051, n20053, n20055, n20064,
    n20061, n20060, n20063, n20104, n20067, n20068, n20093, n20074, n20072,
    n20073, n20075, n20077, n20080, n20079, n20081, n20084, n20083, n20085,
    n20091, n20089, n20087, n20088, n20090, n20092, n20100, n20096, n20101,
    n20098, n20099, n20103, n20111, n20107, n20113, n20109, n20112, n20115,
    n20114, n20116, n20118, n20125, n20123, n20121, n20122, n20124, n20126,
    n20136, n20132, n20133, n20138, n20134, n20135, n20140, n20137, n20139,
    n20143, n20146, n20145, n20151, n20149, n20148, n20150, n20545, n20153,
    n20154, n20157, n20156, n20159, n20158, n20162, n20161, n20173, n20169,
    n20167, n20166, n20168, n20170, n20172, n20171, n20181, n20551, n26228,
    n26274, n20179, n20177, n20176, n20178, n20180, n20183, n20192, n20196,
    n20190, n20188, n20187, n20189, n20191, n20564, n20195, n20194, n20204,
    n20559, n20202, n20200, n20199, n20201, n20203, n20216, n20219, n20214,
    n20212, n20211, n20213, n20215, n20572, n20218, n20217, n20227, n20567,
    n20225, n20223, n20222, n20224, n20226, n20230, n20231, n20232, n20241,
    n20244, n20239, n20237, n20236, n20238, n20240, n20579, n20243, n20242,
    n20252, n20575, n20250, n20248, n20247, n20249, n20251, n20255, n20256,
    n20270, n20262, n20264, n20265, n20582, n20269, n20268, n20272, n20271,
    n20279, n20277, n20275, n20274, n20276, n20278, n20328, n20284, n20285,
    n20286, n20291, n20289, n20288, n20290, n20295, n20592, n20294, n20597,
    n20297, n20296, n20305, n20303, n20301, n20300, n20302, n20304, n20307,
    n20308, n20309, n20314, n20312, n20311, n20313, n20318, n20316, n20600,
    n20317, n20605, n20320, n20319, n20327, n20325, n20323, n20322, n20324,
    n20326, n20329, n20340, n20332, n20341, n20338, n20336, n20335, n20337,
    n20339, n20613, n20608, n20345, n20343, n20344, n20346, n20348, n20347,
    n20351, n20350, n20353, n20358, n20356, n20355, n20357, n20618, n20360,
    n20361, n20365, n20619, n20364, n20368, n20367, n20371, n20370, n20373,
    n20375, n20380, n20378, n20377, n20379, n20626, n20382, n20383, n20390,
    n20386, n20389, n20393, n20392, n20395, n20394, n20397, n20402, n20400,
    n20399, n20401, n20634, n20404, n20403, n20413, n20635, n20411, n20409,
    n20408, n20410, n20412, n20415, n20420, n20418, n20417, n20419, n20642,
    n20422, n20421, n20432, n20643, n20430, n20428, n20426, n20427, n20429,
    n20431, n20434, n20439, n20437, n20436, n20438, n20650, n20441, n20440,
    n20451, n20651, n20449, n20447, n20445, n20446, n20448, n20450, n20453,
    n20458, n20456, n20455, n20457, n20658, n20460, n20459, n20469, n20659,
    n20467, n20465, n20464, n20466, n20468, n20471, n20476, n20474, n20473,
    n20475, n20480, n20664, n20479, n20669, n20483, n20482, n20491, n20489,
    n20487, n20486, n20488, n20490, n20494, n20499, n20497, n20496, n20498,
    n20503, n20502, n20678, n20506, n20505, n20514, n20512, n20510, n20509,
    n20511, n20513, n20516, n20521, n20519, n20518, n20520, n20683, n20523,
    n20522, n20534, n20685, n20532, n20530, n20527, n20529, n20531, n20533,
    n20536, n20690, n20538, n20537, n20541, n20693, n20543, n20542, n20544,
    n20548, n20547, n20696, n20550, n20549, n20554, n20553, n20555, n20699,
    n20558, n20557, n20562, n20561, n20563, n20702, n20566, n20565, n20570,
    n20569, n20571, n20705, n20574, n20573, n20577, n20576, n20578, n20708,
    n20581, n20580, n20584, n20583, n20587, n20586, n20588, n20591, n20590,
    n20595, n20594, n20596, n20713, n20599, n20598, n20603, n20602, n20604,
    n20716, n20607, n20606, n20611, n20610, n20612, n20719, n20615, n20614,
    n20617, n20621, n20620, n20722, n20623, n20622, n20625, n20629, n20628,
    n20725, n20631, n20630, n20633, n20637, n20636, n20728, n20639, n20638,
    n20641, n20645, n20644, n20731, n20647, n20646, n20649, n20653, n20652,
    n20734, n20655, n20654, n20657, n20661, n20660, n20737, n20663, n20662,
    n20667, n20666, n20668, n20740, n20671, n20670, n20676, n20675, n20677,
    n20743, n20680, n20679, n20682, n20687, n20686, n20746, n20689, n20688,
    n20692, n20691, n20695, n20694, n20698, n20697, n20701, n20700, n20704,
    n20703, n20707, n20706, n20710, n20709, n20712, n20711, n20715, n20714,
    n20718, n20717, n20721, n20720, n20724, n20723, n20727, n20726, n20730,
    n20729, n20733, n20732, n20736, n20735, n20739, n20738, n20742, n20741,
    n20745, n20744, n20748, n20747, n20757, n20750, n20751, n20755, n20753,
    n20754, n20756, n20764, n20762, n20761, n20763, n20771, n20769, n20768,
    n20770, n20778, n20776, n20775, n20777, n20784, n20782, n20781, n20783,
    n20791, n20789, n20788, n20790, n20800, n20798, n20797, n20799, n20804,
    n20803, n20817, n20815, n20813, n21498, n20811, n20809, n20808, n20810,
    n20812, n20814, n20816, n20820, n20902, n20822, n20821, n20823, n20833,
    n20825, n24811, n20827, n20826, n20829, n20828, n20831, n20830, n20832,
    n20837, n20838, n20848, n20846, n20840, n20839, n20842, n20841, n20844,
    n20843, n20845, n20847, n20852, n20853, n20862, n20860, n20854, n24915,
    n20856, n20855, n20858, n20857, n20859, n20861, n20864, n20866, n20877,
    n20875, n20869, n20868, n20871, n20870, n20873, n20872, n20874, n20876,
    n20880, n20891, n20889, n20885, n20883, n20882, n20884, n20887, n20886,
    n20888, n20890, n20893, n20895, n21016, n20897, n21015, n20898, n20900,
    n20906, n20904, n20905, n20907, n20916, n20914, n20908, n24854, n20910,
    n20909, n20912, n20911, n20913, n20915, n20919, n20929, n20927, n20921,
    n24879, n20923, n20922, n20925, n20924, n20926, n20928, n20941, n20939,
    n20935, n20933, n20932, n20934, n20937, n20936, n20938, n20940, n20945,
    n20946, n20958, n20947, n20956, n20952, n20950, n20949, n20951, n20954,
    n20953, n20955, n20957, n20962, n20972, n20970, n20966, n20964, n20963,
    n20965, n20968, n20967, n20969, n20971, n20975, n20977, n20982, n20980,
    n20978, n24739, n20979, n20981, n20984, n20983, n20986, n20985, n20989,
    n20999, n20997, n20990, n24895, n20992, n20991, n20995, n20993, n20994,
    n20996, n20998, n21003, n21004, n21014, n21012, n21006, n21005, n21008,
    n21007, n21010, n21009, n21011, n21013, n21018, n21019, n21029, n21022,
    n21020, n24831, n21021, n21024, n21023, n21027, n21026, n21028, n24334,
    n21033, n21034, n21392, n21159, n21369, n21038, n21036, n21041, n21039,
    n21040, n21220, n21046, n21212, n21211, n21044, n21043, n21042, n21210,
    n21045, n21047, n21055, n21049, n21048, n21054, n21051, n21050, n21053,
    n21052, n21057, n21056, n21065, n21060, n21059, n21063, n21062, n21064,
    n21075, n21067, n21066, n21077, n21069, n21068, n21076, n21073, n21079,
    n21078, n21080, n21082, n21081, n21087, n21084, n21083, n21086, n21085,
    n21089, n21088, n21096, n21092, n21091, n21099, n21094, n21093, n21098,
    n21095, n21097, n21101, n21100, n21107, n21103, n21102, n21115, n21105,
    n21104, n21114, n21106, n21108, n21121, n21111, n21110, n21127, n21113,
    n21112, n21126, n21119, n21117, n21116, n21118, n21120, n21140, n21123,
    n21122, n21145, n21125, n21124, n21144, n21131, n21129, n21128, n21130,
    n21138, n21133, n21132, n21142, n21137, n21135, n21134, n21143, n21136,
    n21141, n21139, n21149, n21147, n21146, n21148, n21151, n21150, n21171,
    n21153, n21152, n21170, n21154, n21156, n21155, n21186, n21158, n21157,
    n21185, n21167, n21161, n21341, n21160, n21174, n21165, n21163, n21162,
    n21175, n21164, n21166, n21169, n21179, n21173, n21172, n21177, n21176,
    n21178, n21180, n21182, n21181, n21197, n21184, n21183, n21196, n21190,
    n21188, n21187, n21189, n21191, n21193, n21192, n21205, n21195, n21194,
    n21204, n21201, n21199, n21198, n21200, n21202, n21209, n21207, n21206,
    n21208, n21216, n21214, n21213, n21215, n21217, n21222, n21221, n21230,
    n21224, n21223, n21229, n21226, n21225, n21227, n21231, n21232, n21233,
    n21242, n21236, n21235, n21241, n21238, n21237, n21239, n21243, n21245,
    n21244, n21249, n21247, n21246, n21248, n21251, n21254, n21253, n21260,
    n21258, n21256, n21255, n21257, n21264, n21262, n21261, n21263, n21270,
    n21266, n21265, n21268, n21267, n21269, n21272, n21271, n21281, n21274,
    n21273, n21280, n21275, n21277, n21276, n21285, n21279, n21278, n21284,
    n21283, n21282, n21286, n21288, n21287, n21293, n21290, n21289, n21292,
    n21291, n21295, n21294, n21296, n21299, n21298, n21303, n21302, n21300,
    n21301, n21305, n21304, n21315, n21307, n21306, n21314, n21308, n21311,
    n21310, n21327, n21313, n21312, n21326, n21319, n21317, n21316, n21318,
    n21320, n21322, n21321, n21332, n21325, n21324, n21331, n21329, n21330,
    n21335, n21334, n21349, n21337, n21336, n21348, n21338, n21344, n21342,
    n21343, n21373, n21347, n21346, n21372, n21351, n21350, n21355, n22127,
    n21354, n21358, n21357, n21361, n21360, n25593, n21376, n21362, n21450,
    n21364, n21368, n21385, n21366, n21367, n21382, n21370, n21381, n21375,
    n21374, n21388, n21379, n21378, n21380, n21384, n21383, n21386, n21387,
    n21389, n21390, n21391, n21393, n21399, n21397, n21396, n21398, n24518,
    n21400, n21406, n21404, n21405, n21519, n21442, n21639, n21679, n21827,
    n21869, n21429, n24969, n21428, n21416, n21419, n21418, n21420, n21421,
    n25122, n21422, n21423, n21425, n21424, n21426, n21427, n21844, n21433,
    n21434, n21435, n21743, n21438, n21439, n21443, n21540, n21585, n21448,
    n21452, n21451, n21453, n21458, n21894, n21468, n21895, n21466, n21902,
    n21472, n21464, n21465, n21467, n21901, n21476, n21474, n21471, n21473,
    n21475, n21481, n21479, n21480, n21482, n21485, n21484, n21491, n21489,
    n21488, n21490, n21494, n21493, n21506, n21504, n21502, n21500, n21499,
    n21501, n21503, n21505, n21509, n21510, n21514, n21512, n21511, n21513,
    n21516, n21515, n21531, n21520, n21908, n21529, n21909, n21527, n21525,
    n21523, n21524, n21526, n21528, n21530, n21533, n21537, n21535, n21534,
    n21536, n21927, n21539, n21538, n21554, n21919, n21552, n21543, n21920,
    n21550, n21548, n21546, n21547, n21549, n21551, n21553, n21557, n21567,
    n21570, n21565, n21563, n21562, n21564, n21566, n21938, n21569, n21568,
    n21581, n21930, n21579, n21571, n21931, n21577, n21575, n21573, n21574,
    n21576, n21578, n21580, n21583, n21593, n21596, n21591, n21589, n21588,
    n21590, n21592, n21949, n21595, n21594, n21608, n21941, n21606, n21942,
    n21604, n21602, n21600, n21601, n21603, n21605, n21607, n21610, n21614,
    n21612, n21611, n21613, n21960, n21616, n21615, n21630, n21952, n21628,
    n21953, n21626, n21624, n21622, n21623, n21625, n21627, n21629, n21632,
    n21636, n21634, n21633, n21635, n21971, n21638, n21637, n21651, n21963,
    n21649, n21641, n21964, n21647, n21645, n21643, n21644, n21646, n21648,
    n21650, n21653, n21657, n21655, n21654, n21656, n21981, n21659, n21658,
    n21675, n21974, n21673, n21663, n21665, n21977, n21777, n21671, n21669,
    n21667, n21668, n21670, n21672, n21674, n21677, n21690, n21683, n21680,
    n21682, n21688, n21686, n21685, n21687, n21689, n21992, n21693, n21691,
    n21692, n21704, n21984, n21702, n21985, n21700, n21698, n21696, n21697,
    n21699, n21701, n21703, n21706, n21715, n21719, n21713, n21711, n21710,
    n21712, n21714, n22003, n21718, n21716, n21717, n21731, n21995, n21729,
    n21721, n21996, n21727, n21725, n21724, n21726, n21728, n21730, n21733,
    n21739, n21737, n21736, n21738, n22014, n21742, n21740, n21741, n21754,
    n22006, n21752, n22007, n21750, n21748, n21746, n21747, n21749, n21751,
    n21753, n21756, n21766, n21770, n21764, n21762, n21761, n21763, n21765,
    n22024, n21769, n21767, n21768, n21786, n22017, n21784, n21773, n21776,
    n21775, n22020, n21782, n21780, n21779, n21781, n21783, n21785, n21788,
    n21797, n21801, n21795, n21793, n21792, n21794, n21796, n22035, n21800,
    n21798, n21799, n21814, n22027, n21812, n22028, n21810, n21808, n21806,
    n21807, n21809, n21811, n21813, n21816, n21822, n21820, n21819, n21821,
    n22047, n21825, n21823, n21824, n21840, n22039, n21838, n22040, n21836,
    n21834, n21832, n21833, n21835, n21837, n21839, n21842, n21851, n21858,
    n21849, n21847, n21846, n21848, n21850, n22057, n21852, n21853, n21854,
    n21857, n21855, n21856, n21865, n22050, n21863, n21859, n22051, n21861,
    n21860, n21862, n21864, n21867, n21875, n21879, n21873, n21871, n21870,
    n21872, n21874, n22067, n21878, n21876, n21877, n21893, n22060, n21891,
    n21883, n21881, n21882, n21889, n21884, n21885, n21887, n22061, n21888,
    n21890, n21892, n21898, n21896, n21897, n22070, n21900, n21899, n21905,
    n21903, n21904, n22073, n21907, n21906, n21914, n21912, n21911, n21913,
    n21915, n22079, n21918, n21917, n21925, n21923, n21922, n21924, n21926,
    n22082, n21929, n21928, n21936, n21934, n21933, n21935, n21937, n22085,
    n21940, n21939, n21947, n21945, n21944, n21946, n21948, n22088, n21951,
    n21950, n21958, n21956, n21955, n21957, n21959, n22091, n21962, n21961,
    n21969, n21967, n21966, n21968, n21970, n22094, n21973, n21972, n21979,
    n21976, n21978, n21980, n22097, n21983, n21982, n21990, n21988, n21987,
    n21989, n21991, n22100, n21994, n21993, n22001, n21999, n21998, n22000,
    n22002, n22103, n22005, n22004, n22012, n22010, n22009, n22011, n22013,
    n22106, n22016, n22015, n22022, n22019, n22021, n22023, n22109, n22026,
    n22025, n22033, n22031, n22030, n22032, n22034, n22112, n22037, n22036,
    n22045, n22043, n22042, n22044, n22046, n22115, n22049, n22048, n22055,
    n22053, n22052, n22054, n22056, n22118, n22059, n22058, n22065, n22063,
    n22062, n22064, n22066, n22121, n22069, n22068, n22072, n22071, n22075,
    n22074, n22078, n22077, n22081, n22080, n22084, n22083, n22087, n22086,
    n22090, n22089, n22093, n22092, n22096, n22095, n22099, n22098, n22102,
    n22101, n22105, n22104, n22108, n22107, n22111, n22110, n22114, n22113,
    n22117, n22116, n22120, n22119, n22123, n22122, n22131, n22125, n22126,
    n22129, n22128, n22130, n23123, n22138, n22136, n22134, n22135, n22137,
    n22144, n22142, n22141, n22143, n22149, n24519, n22147, n22146, n22148,
    n23143, n22155, n22153, n22152, n22154, n22162, n22157, n22160, n22159,
    n22161, n23157, n22170, n22168, n22167, n22169, n22173, n22175, n22185,
    n22183, n22181, n22177, n23608, n22179, n22178, n22180, n22182, n22184,
    n22188, n22198, n22196, n22192, n22190, n22189, n22191, n22194, n22193,
    n22195, n22197, n22201, n22369, n22370, n22204, n22205, n22217, n22215,
    n22206, n23534, n22208, n22213, n22211, n23732, n22210, n22212, n22214,
    n22216, n22220, n22222, n22232, n22936, n22230, n22228, n22226, n22224,
    n23731, n22225, n22227, n22229, n22231, n22235, n22236, n22246, n22244,
    n22240, n22238, n22237, n22239, n22242, n22241, n22243, n22245, n22249,
    n22251, n22263, n22261, n22254, n23576, n22256, n22255, n22259, n22258,
    n22260, n22262, n22266, n22276, n22274, n22272, n22270, n22268, n22267,
    n22269, n22271, n22273, n22275, n22278, n22280, n22289, n22287, n22285,
    n22281, n23647, n22283, n22282, n22284, n22286, n22288, n22292, n22294,
    n22305, n22966, n22303, n22681, n22301, n22634, n22299, n22297, n23668,
    n22298, n22300, n22302, n22304, n22308, n22318, n22316, n22314, n22312,
    n22310, n22309, n22311, n22313, n22315, n22317, n22321, n22331, n22329,
    n22327, n22325, n22323, n22322, n22324, n22326, n22328, n22330, n22335,
    n22336, n22347, n22345, n22340, n22338, n23590, n22339, n22343, n22342,
    n22344, n22346, n22350, n22352, n22354, n22353, n22355, n22366, n22364,
    n22362, n22572, n22360, n22358, n22357, n22359, n22361, n22363, n22365,
    n22368, n22373, n22372, n22374, n22375, n22385, n22800, n22383, n22379,
    n22377, n23557, n22378, n22381, n22380, n22382, n22384, n22388, n22398,
    n22396, n22394, n22390, n23687, n22392, n22391, n22393, n22395, n22397,
    n22402, n22403, n22412, n22410, n22408, n22406, n22404, n23635, n22405,
    n22407, n22409, n22411, n22420, n22418, n22415, n22424, n22416, n22417,
    n22419, n22809, n22428, n22426, n22423, n22425, n22427, n22444, n22442,
    n22431, n22430, n22434, n22433, n22438, n22437, n22440, n22439, n22441,
    n22443, n22445, n22449, n22448, n22451, n22456, n22454, n22453, n22455,
    n22460, n22459, n22462, n22461, n22471, n22469, n22818, n22467, n22465,
    n22464, n22466, n22468, n22470, n22828, n22487, n22829, n22473, n22485,
    n22483, n22481, n22475, n22479, n22477, n22476, n22478, n22480, n22482,
    n22484, n22486, n22490, n22489, n22508, n22493, n22846, n22506, n24025,
    n22504, n22502, n22500, n22498, n22497, n22499, n22501, n22503, n22505,
    n22507, n22512, n22856, n22511, n22534, n22520, n22518, n22517, n22519,
    n22525, n22523, n22524, n22868, n22526, n22864, n22530, n22528, n22529,
    n22531, n22533, n22532, n22539, n22861, n22537, n22536, n22538, n22540,
    n22542, n22541, n22563, n22547, n22546, n22872, n22561, n22549, n22873,
    n22559, n22557, n22553, n22552, n22555, n22554, n22556, n22558, n22560,
    n22562, n22567, n22566, n22887, n22584, n22571, n22888, n22582, n22580,
    n22578, n22576, n22574, n22573, n22575, n22577, n22579, n22581, n22583,
    n22587, n22898, n22586, n22903, n22602, n22600, n22598, n22596, n22594,
    n22592, n22591, n22593, n22595, n22597, n22599, n22601, n22606, n22914,
    n22605, n22919, n22623, n22616, n22609, n22608, n22611, n22610, n22614,
    n22613, n22615, n22621, n22619, n22924, n22620, n22622, n22628, n22626,
    n22929, n22627, n22631, n22934, n22647, n22935, n22645, n22643, n22639,
    n22637, n22636, n22638, n22641, n22640, n22642, n22644, n22646, n22651,
    n22945, n22650, n22663, n22654, n22653, n22659, n22657, n22658, n22961,
    n22662, n22661, n22675, n22950, n22673, n22951, n22671, n22669, n22667,
    n22666, n22668, n22670, n22672, n22674, n22964, n22693, n22677, n22679,
    n22965, n22691, n22689, n22685, n22683, n22682, n22684, n22687, n22686,
    n22688, n22690, n22692, n22697, n22975, n22696, n22701, n22700, n22980,
    n22721, n22704, n22981, n22719, n22717, n22712, n22710, n22709, n22711,
    n22715, n22714, n22716, n22718, n22720, n22727, n22724, n22991, n22726,
    n22996, n22744, n22997, n22742, n22740, n22736, n22734, n22733, n22735,
    n22738, n22737, n22739, n22741, n22743, n22748, n23008, n22747, n22751,
    n23013, n22769, n23014, n22767, n22765, n22760, n22758, n22757, n22759,
    n22763, n22762, n22764, n22766, n22768, n22774, n23026, n22773, n23780,
    n22779, n22778, n23746, n23745, n23748, n22781, n23049, n22796, n22785,
    n22787, n22788, n22794, n22792, n22791, n22793, n22795, n23057, n22799,
    n22797, n22798, n22808, n22806, n23050, n22804, n22802, n22801, n22803,
    n22805, n22807, n22814, n22812, n22813, n23063, n22816, n22815, n22823,
    n22821, n22820, n22822, n22825, n23066, n22827, n22826, n22840, n24201,
    n22831, n22838, n22836, n22834, n23953, n22833, n22835, n22837, n22839,
    n22842, n22844, n22843, n22855, n22853, n22851, n22849, n22848, n22850,
    n22852, n22854, n22858, n22857, n23072, n22860, n22859, n22866, n22863,
    n22865, n22867, n23075, n22870, n22869, n24247, n22884, n22882, n22880,
    n22878, n22876, n22875, n22877, n22879, n22881, n22883, n23078, n22886,
    n22885, n22897, n22895, n22893, n22891, n22890, n22892, n22894, n22896,
    n22900, n22899, n23081, n22902, n22901, n22913, n22911, n22909, n22907,
    n22906, n22908, n22910, n22912, n22916, n22915, n23084, n22918, n22917,
    n22928, n22923, n22921, n22920, n22922, n22926, n22925, n22927, n22931,
    n22930, n23087, n22933, n22932, n22944, n22942, n22940, n22938, n22937,
    n22939, n22941, n22943, n22947, n22946, n23090, n22949, n22948, n22959,
    n22957, n22955, n22954, n22956, n22958, n22960, n23093, n22963, n22962,
    n22974, n22972, n22970, n22968, n22967, n22969, n22971, n22973, n22977,
    n22976, n23096, n22979, n22978, n22990, n22988, n22986, n22984, n22983,
    n22985, n22987, n22989, n22993, n22992, n23099, n22995, n22994, n23007,
    n23005, n23003, n23001, n23000, n23002, n23004, n23006, n23010, n23009,
    n23102, n23012, n23011, n23025, n23023, n23021, n23019, n23018, n23020,
    n23022, n23024, n23028, n23027, n23105, n23030, n23029, n23043, n23041,
    n23039, n23037, n23036, n23038, n23040, n23042, n23046, n23045, n23108,
    n23048, n23047, n23055, n23053, n23052, n23054, n23056, n23111, n23059,
    n23058, n23062, n23061, n23065, n23064, n23068, n23067, n23071, n23070,
    n23074, n23073, n23077, n23076, n23080, n23079, n23083, n23082, n23086,
    n23085, n23089, n23088, n23092, n23091, n23095, n23094, n23098, n23097,
    n23101, n23100, n23104, n23103, n23107, n23106, n23110, n23109, n23113,
    n23112, n23122, n23115, n23116, n23120, n23119, n23121, n23129, n23127,
    n23126, n23128, n23131, n23136, n23134, n23133, n23135, n23138, n23142,
    n23140, n23139, n23141, n23148, n23146, n23145, n23147, n23155, n23150,
    n23153, n23152, n23154, n23163, n23158, n23161, n23160, n23162, n23165,
    n23170, n23168, n23169, n23172, n23177, n23175, n23176, n23179, n23182,
    n23186, n23190, n23195, n23193, n23194, n23196, n23200, n23199, n23202,
    n23201, n23209, n23205, n23206, n23208, n23214, n24203, n23212, n23210,
    n23471, n23211, n23213, n23216, n23215, n23927, n23218, n23229, n23223,
    n23224, n23227, n23226, n23228, n23233, n23231, n23230, n23232, n23236,
    n23491, n23249, n23239, n23245, n23240, n23243, n23242, n23244, n23247,
    n23246, n23248, n23251, n23253, n23262, n23256, n23255, n23260, n23258,
    n23257, n23259, n23261, n23263, n23429, n23285, n23270, n23268, n23267,
    n23269, n23291, n23273, n23272, n23290, n23275, n23276, n23283, n23281,
    n23280, n23282, n23284, n23287, n23286, n23289, n23288, n23296, n23292,
    n23294, n23295, n23301, n23297, n23408, n23299, n23298, n23300, n23302,
    n23519, n23306, n23304, n23303, n23305, n23315, n23310, n23313, n23312,
    n23314, n23318, n23328, n23321, n23320, n23326, n23324, n23323, n23325,
    n23327, n23330, n23454, n23349, n23334, n23333, n23347, n23335, n23338,
    n23340, n23341, n23345, n23344, n23346, n23348, n23358, n23352, n23393,
    n23353, n23354, n23355, n23357, n23360, n23359, n23362, n23361, n23370,
    n23365, n23368, n23367, n23369, n23377, n23373, n23375, n23376, n23379,
    n23378, n23387, n23385, n23383, n23384, n23386, n23406, n23388, n23398,
    n24307, n23392, n23395, n23394, n23396, n23397, n23425, n23403, n23402,
    n23404, n23405, n23407, n23423, n23445, n23412, n23411, n23446, n23413,
    n23421, n23418, n23417, n23431, n23430, n23419, n23420, n23422, n23427,
    n23424, n23426, n23428, n23443, n23457, n23441, n23432, n23433, n23434,
    n23463, n23435, n23436, n23438, n23439, n23440, n23442, n23452, n23455,
    n23449, n23447, n23448, n23456, n23450, n23451, n23453, n23469, n23474,
    n23462, n23472, n23459, n23458, n23473, n23460, n23461, n23467, n23484,
    n23482, n23465, n23466, n23468, n23470, n23481, n23476, n23475, n23508,
    n23506, n23477, n23479, n23509, n23478, n23480, n23489, n23485, n23492,
    n23487, n23488, n23490, n23505, n23494, n23495, n23515, n23496, n23497,
    n23498, n23499, n23500, n23503, n23502, n23504, n23514, n23520, n23507,
    n23511, n23510, n23521, n23512, n23513, n23540, n23517, n23531, n23518,
    n23529, n23536, n23524, n23522, n23523, n23535, n23525, n23527, n23526,
    n23528, n23530, n23533, n23551, n23547, n23559, n23538, n23537, n23558,
    n23539, n23546, n23553, n23543, n23542, n23544, n23545, n23549, n23548,
    n23550, n23582, n23554, n23555, n23568, n23556, n23566, n23570, n23561,
    n23560, n23569, n23562, n23564, n23563, n23565, n23567, n23579, n23591,
    n23572, n23571, n23592, n23573, n23578, n23575, n23577, n23581, n23580,
    n23588, n23584, n23598, n23597, n23585, n23586, n23587, n23589, n23603,
    n23613, n23594, n23593, n23612, n23595, n23601, n23622, n23599, n23600,
    n23602, n23605, n23604, n23607, n23610, n23609, n23621, n23611, n23617,
    n23615, n23614, n23616, n23636, n23619, n23618, n23620, n23628, n23631,
    n23630, n23625, n23624, n23626, n23627, n23633, n23644, n23634, n23642,
    n23637, n23648, n23649, n23638, n23640, n23639, n23641, n23643, n23646,
    n23666, n24047, n23670, n23651, n23650, n23669, n23652, n23654, n23653,
    n23664, n23659, n23658, n23679, n23662, n23661, n23663, n23665, n23667,
    n23677, n23692, n23672, n23671, n23691, n23673, n23675, n23674, n23676,
    n23683, n23701, n23680, n23700, n23681, n23682, n23686, n23690, n23689,
    n23699, n24036, n23694, n23693, n23710, n23695, n23713, n23697, n23696,
    n23698, n23705, n23702, n23703, n23704, n23709, n23717, n23712, n23714,
    n23718, n23715, n23716, n23728, n23719, n23727, n23725, n23730, n23734,
    n23733, n23736, n23735, n23761, n23738, n23774, n23741, n23742, n23744,
    n23743, n24246, n23747, n24248, n23757, n23750, n23752, n23755, n23754,
    n24244, n23756, n23758, n23759, n23760, n23764, n23762, n23763, n23766,
    n24235, n23768, n23767, n23787, n23771, n23770, n23784, n23773, n23775,
    n23782, n23778, n23779, n24229, n23781, n23783, n24237, n24009, n23785,
    n23786, n23788, n23791, n23790, n23793, n23792, n23795, n23800, n23810,
    n23798, n23797, n23799, n24225, n24214, n23802, n23809, n23804, n23803,
    n23807, n23806, n23808, n23812, n24221, n23811, n23814, n24217, n23813,
    n23817, n23816, n23822, n23819, n24202, n23821, n23841, n23824, n23835,
    n23827, n23826, n23833, n23830, n24206, n23832, n23834, n24208, n23836,
    n23837, n23839, n23838, n23840, n23844, n23843, n23847, n23846, n23866,
    n24189, n23862, n23850, n23860, n24195, n23858, n23856, n23855, n23857,
    n23859, n24194, n23861, n23864, n23863, n23865, n23869, n23868, n23871,
    n23870, n23896, n24177, n23891, n23877, n23876, n23884, n23879, n23912,
    n23881, n23882, n24183, n23883, n23889, n23887, n23888, n24182, n23890,
    n23894, n23893, n23895, n23899, n23900, n23902, n23901, n24174, n23904,
    n24169, n23909, n24167, n23907, n23908, n23916, n23911, n23913, n24170,
    n23915, n23917, n23918, n23921, n23920, n23923, n23922, n23930, n23928,
    n23929, n24160, n23932, n23935, n23933, n23934, n23938, n23937, n23939,
    n23946, n23943, n24154, n23945, n23948, n23947, n23951, n23952, n23962,
    n23955, n23954, n23960, n23956, n23984, n23957, n24147, n23959, n23961,
    n24149, n23964, n24143, n23965, n23974, n23969, n23968, n23972, n23971,
    n23973, n23975, n23977, n23976, n23979, n23978, n23982, n23981, n24008,
    n23986, n23985, n23997, n24130, n24005, n23987, n23989, n23996, n23992,
    n23994, n23995, n23999, n23998, n24140, n24133, n24134, n24002, n24003,
    n24004, n24006, n24007, n24010, n24018, n24013, n24017, n24016, n24127,
    n24020, n24032, n24024, n24023, n24030, n24028, n24029, n24031, n24035,
    n24116, n24038, n24037, n24040, n24039, n24043, n24042, n24046, n24045,
    n24049, n24048, n24051, n24050, n24055, n24054, n24058, n24057, n24061,
    n24060, n24064, n24063, n24068, n24067, n24071, n24070, n24074, n24073,
    n24077, n24076, n24080, n24079, n24083, n24082, n24087, n24086, n24090,
    n24089, n24093, n24092, n24095, n24094, n24098, n24097, n24100, n24099,
    n24103, n24102, n24105, n24104, n24109, n24108, n24112, n24111, n24115,
    n24118, n24114, n24120, n24119, n24129, n24125, n24124, n24126, n24254,
    n24128, n24142, n24138, n24132, n24136, n24135, n24137, n24139, n24257,
    n24141, n24153, n24146, n24145, n24151, n24148, n24150, n24260, n24152,
    n24164, n24157, n24156, n24162, n24159, n24161, n24263, n24163, n24176,
    n24166, n24168, n24172, n24171, n24173, n24266, n24175, n24188, n24180,
    n24179, n24181, n24186, n24184, n24185, n24269, n24187, n24200, n24192,
    n24191, n24193, n24198, n24196, n24197, n24272, n24199, n24212, n24205,
    n24204, n24210, n24207, n24209, n24275, n24211, n24227, n24215, n24219,
    n24218, n24223, n24222, n24224, n24278, n24226, n24239, n24233, n24232,
    n24234, n24236, n24281, n24238, n24253, n24243, n24245, n24250, n24249,
    n24285, n24252, n24256, n24255, n24259, n24258, n24262, n24261, n24265,
    n24264, n24268, n24267, n24271, n24270, n24274, n24273, n24277, n24276,
    n24280, n24279, n24283, n24282, n24288, n24287, n24291, n24290, n24294,
    n24293, n24297, n24296, n24300, n24299, n24303, n24302, n24306, n24305,
    n24310, n24309, n24313, n24312, n24315, n24314, n24318, n24317, n24322,
    n24321, n24326, n24325, n24329, n24328, n24332, n24331, n24335, n24913,
    n24337, n24657, n24339, n24338, n24348, n24342, n24344, n24343, n24346,
    n24345, n24347, n24352, n24350, n24717, n24351, n24361, n24355, n24359,
    n24357, n24356, n24358, n24360, n24364, n24362, n24575, n24363, n24373,
    n24369, n24367, n24368, n24371, n24370, n24372, n24374, n24682, n24376,
    n24375, n24388, n24380, n24381, n24382, n24384, n24383, n24386, n24385,
    n24387, n24391, n24774, n24393, n24392, n24399, n24397, n24396, n24398,
    n24406, n24403, n24404, n24405, n24409, n24407, n24622, n24408, n24418,
    n24412, n24416, n24414, n24413, n24415, n24417, n25080, n24421, n24419,
    n24596, n24420, n24433, n24428, n24425, n24426, n24427, n24431, n24430,
    n24432, n24437, n24435, n24697, n24436, n24448, n24441, n24442, n24444,
    n24443, n24446, n24445, n24447, n24450, n24451, n24453, n24461, n24457,
    n24456, n24459, n25266, n24458, n24460, n24465, n24463, n24784, n24464,
    n24481, n24468, n24469, n24472, n24479, n24477, n24476, n24478, n24480,
    n24486, n24483, n24485, n24498, n24496, n24494, n24490, n24492, n24493,
    n24495, n24497, n24503, n24501, n24637, n24502, n24515, n24507, n24510,
    n24509, n24513, n24512, n24514, n24896, n24517, n24933, n24523, n24520,
    n24925, n24522, n24524, n24525, n24533, n25283, n24535, n24526, n24545,
    n24527, n24531, n24529, n24528, n24530, n24532, n24559, n24534, n24539,
    n24744, n24536, n24558, n24537, n24538, n24543, n24541, n24540, n24542,
    n24553, n24564, n24544, n24549, n24771, n24546, n24563, n24547, n24548,
    n24551, n24550, n24552, n24555, n24554, n24557, n24556, n24573, n24561,
    n24560, n24579, n24580, n24562, n24571, n24567, n24566, n24585, n24568,
    n24584, n24569, n24570, n24572, n24574, n24578, n24577, n24594, n24582,
    n24581, n24600, n24599, n24583, n24592, n24588, n24587, n24605, n24589,
    n24604, n24590, n24591, n24593, n24595, n24598, n25355, n24597, n24614,
    n24602, n24601, n24626, n24625, n24603, n24612, n24608, n24607, n24616,
    n24609, n24615, n24610, n24611, n24613, n24618, n24617, n24646, n24619,
    n24645, n24620, n24624, n24621, n24623, n24635, n24629, n24628, n24641,
    n24640, n24630, n24633, n24632, n24634, n24636, n24639, n25349, n24638,
    n24655, n24643, n24642, n24667, n24666, n24644, n24653, n24649, n24648,
    n24661, n24650, n24660, n24651, n24652, n24654, n24656, n24659, n25343,
    n24658, n24675, n24663, n24662, n24686, n24664, n24685, n24665, n24673,
    n24670, n24669, n24677, n24676, n24671, n24672, n24674, n24679, n24678,
    n24698, n24699, n24680, n24684, n24681, n24683, n24695, n24689, n24688,
    n24708, n24690, n24709, n24691, n24693, n25340, n24692, n24694, n24712,
    n25331, n24696, n24706, n24704, n24701, n24700, n24727, n24726, n24702,
    n24703, n24705, n24715, n24711, n24710, n24720, n24719, n24713, n24714,
    n24716, n24734, n24718, n24753, n24722, n24721, n24752, n24723, n24732,
    n24724, n24740, n24729, n24728, n24730, n24731, n24733, n24737, n24735,
    n25326, n24736, n24750, n25321, n24738, n24749, n24761, n24743, n24742,
    n24760, n24745, n24747, n24746, n24748, n24758, n24767, n24755, n24754,
    n24766, n24756, n24757, n24794, n24759, n24795, n24763, n24762, n24764,
    n24778, n24769, n24768, n24787, n24785, n24770, n24786, n24772, n24776,
    n24773, n24775, n24777, n24782, n24780, n25316, n24781, n24783, n24806,
    n24792, n24789, n24788, n24791, n24790, n24793, n24818, n24804, n24798,
    n24797, n24801, n24800, n24799, n24802, n24812, n24803, n24805, n24809,
    n24807, n25312, n24808, n24810, n24829, n24813, n24838, n24841, n24839,
    n24814, n24815, n24827, n24816, n25307, n24825, n24822, n24819, n24821,
    n24820, n24823, n24833, n24824, n24826, n24828, n24830, n24849, n24834,
    n24855, n24836, n24835, n24837, n24856, n24847, n24840, n24862, n24844,
    n24843, n24845, n24864, n24846, n24848, n24852, n24850, n24851, n24853,
    n24873, n24874, n24860, n24857, n24859, n24858, n24861, n24882, n24871,
    n24868, n24865, n24867, n24866, n24869, n24887, n24870, n24872, n24877,
    n25303, n24876, n24878, n24881, n25300, n24880, n24893, n24885, n24905,
    n24883, n24904, n24884, n24891, n24900, n24888, n24899, n24889, n24890,
    n24892, n24894, n24898, n25294, n24897, n24912, n24901, n24929, n24902,
    n24910, n24907, n24906, n24920, n24919, n24908, n24909, n24911, n24914,
    n24918, n24917, n24938, n24922, n24921, n24924, n24923, n24926, n24936,
    n24931, n24930, n24932, n24935, n24937, n24940, n24939, n24943, n24942,
    n24963, n25504, n24946, n25510, n24952, n25226, n24945, n24961, n24949,
    n24951, n24954, n24953, n24959, n24957, n24956, n24958, n25514, n24960,
    n24962, n24966, n24965, n24981, n24968, n24975, n25492, n25271, n24973,
    n24972, n24974, n25498, n24977, n25490, n24978, n24979, n24980, n24989,
    n25068, n24985, n24990, n24983, n24984, n25496, n24987, n24986, n24988,
    n24991, n25495, n25483, n24993, n24992, n25007, n24995, n24999, n25478,
    n24998, n25004, n25002, n25001, n25003, n25485, n25005, n25006, n25008,
    n25011, n25010, n25013, n25012, n25015, n25014, n25020, n25060, n25016,
    n25018, n25466, n25019, n25039, n25024, n25023, n25027, n25470, n25026,
    n25032, n25030, n25031, n25472, n25034, n25035, n25037, n25036, n25038,
    n25041, n25044, n25084, n25047, n25046, n25048, n25056, n25453, n25050,
    n25455, n25065, n25053, n25055, n25054, n25058, n25057, n25463, n25062,
    n25061, n25063, n25064, n25066, n25070, n25457, n25069, n25072, n25071,
    n25075, n25074, n25103, n25078, n25082, n25081, n25087, n25446, n25085,
    n25086, n25448, n25089, n25445, n25096, n25094, n25442, n25095, n25097,
    n25098, n25101, n25100, n25102, n25110, n25108, n25107, n25109, n25134,
    n25431, n25117, n25112, n25113, n25115, n25429, n25116, n25132, n25143,
    n25144, n25121, n25123, n25125, n25124, n25130, n25128, n25127, n25129,
    n25438, n25131, n25133, n25171, n25177, n25173, n25138, n25141, n25140,
    n25419, n25147, n25167, n25145, n25146, n25149, n25148, n25154, n25152,
    n25151, n25153, n25426, n25159, n25192, n25157, n25158, n25422, n25164,
    n25162, n25161, n25163, n25165, n25166, n25168, n25170, n25169, n25172,
    n25409, n25180, n25199, n25211, n25176, n25178, n25179, n25182, n25181,
    n25187, n25185, n25184, n25186, n25416, n25191, n25190, n25196, n25193,
    n25412, n25195, n25197, n25198, n25200, n25202, n25201, n25203, n25205,
    n25204, n25232, n25208, n25398, n25207, n25230, n25210, n25212, n25213,
    n25225, n25216, n25215, n25223, n25220, n25404, n25221, n25222, n25224,
    n25403, n25228, n25227, n25229, n25231, n25235, n25234, n25239, n25237,
    n25388, n25236, n25238, n25262, n25242, n25387, n25249, n25259, n25247,
    n25251, n25250, n25258, n25256, n25255, n25257, n25395, n25260, n25261,
    n25265, n25269, n25268, n25288, n25382, n25272, n25276, n25275, n25381,
    n25278, n25280, n25281, n25286, n25285, n25287, n25375, n25369, n25293,
    n25292, n25295, n25299, n25298, n25301, n25304, n25306, n25305, n25308,
    n25310, n25309, n25313, n25315, n25314, n25317, n25319, n25318, n25322,
    n25324, n25323, n25327, n25329, n25328, n25332, n25334, n25333, n25339,
    n25338, n25341, n25345, n25344, n25347, n25346, n25351, n25350, n25353,
    n25352, n25357, n25356, n25359, n25358, n25364, n25363, n25367, n25366,
    n25372, n25371, n25377, n25376, n25386, n25379, n25380, n25384, n25383,
    n25518, n25385, n25397, n25393, n25391, n25390, n25392, n25394, n25521,
    n25396, n25408, n25401, n25400, n25402, n25406, n25405, n25524, n25407,
    n25418, n25414, n25411, n25413, n25415, n25527, n25417, n25428, n25424,
    n25421, n25423, n25425, n25530, n25427, n25440, n25430, n25436, n25434,
    n25433, n25435, n25437, n25533, n25439, n25452, n25443, n25444, n25450,
    n25447, n25449, n25536, n25451, n25465, n25461, n25456, n25459, n25458,
    n25460, n25462, n25539, n25464, n25476, n25469, n25468, n25474, n25471,
    n25473, n25542, n25475, n25487, n25481, n25480, n25482, n25484, n25545,
    n25486, n25502, n25491, n25494, n25493, n25500, n25497, n25499, n25548,
    n25501, n25517, n25508, n25507, n25512, n25511, n25513, n25552, n25516,
    n25520, n25519, n25523, n25522, n25526, n25525, n25529, n25528, n25532,
    n25531, n25535, n25534, n25538, n25537, n25541, n25540, n25544, n25543,
    n25547, n25546, n25550, n25549, n25555, n25554, n25558, n25557, n25561,
    n25560, n25564, n25563, n25567, n25566, n25570, n25569, n25573, n25572,
    n25576, n25575, n25579, n25578, n25582, n25581, n25585, n25584, n25588,
    n25587, n25591, n25590, n25595, n25594, n25596, n25880, n25610, n25599,
    n25708, n25598, n25608, n25601, n25602, n25604, n25606, n25605, n25607,
    n25609, n25613, n25612, n25623, n25614, n25954, n25621, n25617, n25619,
    n25618, n25620, n25622, n25625, n25798, n25637, n25628, n25627, n25635,
    n25631, n25633, n25632, n25634, n25636, n25640, n25639, n25650, n25641,
    n25902, n25648, n25644, n25646, n25645, n25647, n25649, n25653, n25652,
    n25658, n25720, n25656, n25655, n25657, n25665, n25662, n25663, n25664,
    n25668, n25837, n25681, n25670, n25669, n25679, n25674, n25675, n25677,
    n25676, n25678, n25680, n25682, n25686, n25685, n25688, n25687, n25690,
    n25967, n25705, n25694, n25693, n25703, n25696, n25698, n25701, n25700,
    n25702, n25704, n25709, n25719, n25713, n25715, n25717, n25716, n25718,
    n25722, n25721, n25727, n25726, n25740, n25729, n25858, n25738, n25733,
    n25736, n25735, n25737, n25739, n25753, n25743, n25745, n25744, n25749,
    n26010, n25747, n25748, n25760, n25752, n25754, n25756, n25755, n25758,
    n25757, n25759, n25762, n25761, n25770, n25764, n25768, n25766, n25767,
    n25769, n25777, n25772, n26044, n25775, n25774, n25776, n25788, n25781,
    n25786, n25784, n25785, n25787, n25797, n25791, n25795, n25793, n25792,
    n25794, n25796, n25799, n25817, n25801, n25805, n25803, n25804, n25815,
    n25808, n25810, n25813, n25812, n25814, n25816, n25818, n25828, n25826,
    n25824, n25825, n25827, n25836, n25831, n25834, n25833, n25835, n25838,
    n25856, n25840, n25844, n25842, n25843, n25854, n25847, n25849, n25852,
    n25851, n25853, n25855, n25857, n25868, n25861, n25866, n25864, n25865,
    n25867, n25879, n25871, n25872, n25874, n25877, n25876, n25878, n25881,
    n25900, n25883, n25887, n25885, n25886, n25898, n25890, n25892, n25896,
    n25895, n25897, n25899, n25901, n25912, n25905, n25910, n25908, n25909,
    n25911, n25920, n25915, n25918, n25917, n25919, n25922, n25941, n25925,
    n25927, n25926, n25939, n25929, n25937, n25932, n25933, n25935, n25936,
    n25938, n25940, n25944, n25963, n25947, n25961, n25951, n25952, n25959,
    n25953, n25957, n25956, n25958, n25960, n25962, n25965, n25981, n25968,
    n25970, n25969, n25979, n25972, n25977, n25975, n25976, n25978, n25980,
    n25984, n26004, n25987, n25994, n25992, n25989, n25991, n25993, n26002,
    n26000, n25998, n25999, n26001, n26003, n26006, n26025, n26009, n26023,
    n26014, n26021, n26015, n26019, n26018, n26020, n26022, n26024, n26051,
    n26032, n26041, n26034, n26039, n26038, n26040, n26049, n26045, n26047,
    n26048, n26050, n26392, n26056, n26064, n26055, n26058, n26057, n26063,
    n26061, n26060, n26062, n26397, n26065, n26073, n26071, n26069, n26068,
    n26070, n26072, n26077, n26079, n26382, n26080, n26091, n26084, n26082,
    n26083, n26090, n26088, n26087, n26089, n26387, n26092, n26100, n26098,
    n26096, n26095, n26097, n26099, n26103, n26102, n26105, n26104, n26124,
    n26108, n26110, n26374, n26113, n26121, n26115, n26114, n26120, n26118,
    n26117, n26119, n26379, n26122, n26123, n26136, n26128, n26131, n26134,
    n26366, n26132, n26133, n26135, n26139, n26371, n26142, n26144, n26143,
    n26145, n26147, n26146, n26149, n26148, n26154, n26153, n26157, n26156,
    n26173, n26358, n26159, n26170, n26164, n26162, n26163, n26169, n26167,
    n26166, n26168, n26363, n26171, n26172, n26177, n26176, n26180, n26179,
    n26197, n26350, n26186, n26194, n26185, n26188, n26187, n26193, n26191,
    n26190, n26192, n26355, n26195, n26196, n26342, n26202, n26210, n26201,
    n26204, n26203, n26209, n26207, n26206, n26208, n26347, n26211, n26221,
    n26215, n26214, n26219, n26218, n26220, n26223, n26222, n26226, n26225,
    n26244, n26334, n26236, n26241, n26231, n26230, n26240, n26235, n26238,
    n26237, n26239, n26339, n26242, n26243, n26247, n26328, n26246, n26251,
    n26327, n26250, n26266, n26254, n26265, n26257, n26259, n26260, n26263,
    n26261, n26262, n26264, n26331, n26267, n26269, n26268, n26272, n26271,
    n26276, n26320, n26275, n26296, n26321, n26293, n26281, n26285, n26283,
    n26284, n26292, n26290, n26289, n26291, n26324, n26294, n26295, n26299,
    n26298, n26302, n26301, n26309, n26304, n26307, n26317, n26308, n26314,
    n26313, n26319, n26401, n26318, n26326, n26322, n26323, n26404, n26325,
    n26333, n26329, n26330, n26407, n26332, n26341, n26337, n26336, n26338,
    n26410, n26340, n26349, n26345, n26344, n26346, n26413, n26348, n26357,
    n26353, n26352, n26354, n26416, n26356, n26365, n26361, n26360, n26362,
    n26419, n26364, n26373, n26369, n26368, n26370, n26422, n26372, n26381,
    n26377, n26376, n26378, n26425, n26380, n26389, n26385, n26384, n26386,
    n26428, n26388, n26400, n26395, n26394, n26396, n26432, n26399, n26403,
    n26402, n26406, n26405, n26409, n26408, n26412, n26411, n26415, n26414,
    n26418, n26417, n26421, n26420, n26424, n26423, n26427, n26426, n26430,
    n26429, n26435, n26434, n26438, n26437, n26441, n26440, n26444, n26443,
    n26447, n26446, n26450, n26449, n26453, n26452, n26457, n26456, n13665,
    n20481;
  assign n25267 = ~n25233;
  assign n24316 = n15820 | n15819;
  assign n14111 = ~n22847;
  assign n13133 = n14983;
  assign n25489 = ~n17583 | ~n17582;
  assign n25214 = n16698 | n16697;
  assign n21353 = n17502;
  assign n26252 = n16447 | n16446;
  assign n13124 = ~n14877;
  assign n21402 = n17030;
  assign n26152 = n18473 & n17241;
  assign n13116 = ~n26459;
  assign P1_U3086 = ~n13116;
  assign n26459 = ~P1_STATE_REG_SCAN_IN;
  assign n16572 = ~P2_IR_REG_21__SCAN_IN & ~P2_IR_REG_22__SCAN_IN;
  assign n15554 = ~n16809 | ~n13121;
  assign n13134 = n14983;
  assign n19178 = ~n17213;
  assign n14091 = ~P2_IR_REG_0__SCAN_IN;
  assign n14654 = ~n15810;
  assign n15113 = ~n15087 | ~n15086;
  assign n13563 = n13564 & n26280;
  assign n21975 = ~n17682 | ~n17681;
  assign n25264 = ~n25105;
  assign n17487 = ~n14091 | ~n14090;
  assign n23967 = ~n15022 | ~n15021;
  assign n24190 = ~n15155 | ~n15154;
  assign n17312 = n17255 & n13713;
  assign n13866 = n20095 ^ ~n14004;
  assign n20556 = ~n20170 & ~n13563;
  assign n21598 = ~n17721 | ~n24333;
  assign n25104 = ~n25432;
  assign n22889 = ~n17423 | ~n16809;
  assign n23906 = ~n23854;
  assign n22998 = n15465 & n15464;
  assign n24213 = ~n15218 | ~n15217;
  assign n24131 = ~n17352;
  assign n26205 = n16390 | n16389;
  assign n25389 = ~n14430 | ~n14428;
  assign n25284 = ~n25282;
  assign n16928 = ~n13551 | ~n13550;
  assign n13118 = n26030 | P3_REG2_REG_14__SCAN_IN;
  assign n16337 = ~P3_IR_REG_31__SCAN_IN;
  assign n13119 = n14665 & n14396;
  assign n13120 = n17994 ^ n13363;
  assign n14511 = ~n22874;
  assign n15008 = n15007 | n15073;
  assign n13987 = n14435 & n21772;
  assign n18666 = ~n22257;
  assign n14933 = n14925 & n14699;
  assign n14923 = ~n15452 & ~n14921;
  assign n13527 = ~n13529 & ~n13528;
  assign n13123 = ~n18563;
  assign n18563 = ~n18511 | ~n18503;
  assign n24449 = ~n21032 | ~n25378;
  assign n21032 = n17029 & n21407;
  assign n25884 = n19816 ^ ~n25893;
  assign n19816 = ~n13995 | ~n19815;
  assign n19033 = ~n18920;
  assign n25921 = n19985 ^ ~n19984;
  assign n19985 = ~n13945 | ~n19983;
  assign n15111 = n15113 ^ ~n15088;
  assign n13121 = n16232;
  assign n13122 = n16232;
  assign n16232 = ~n17196;
  assign n24516 = n17035 ^ ~n17034;
  assign n22544 = ~n18027 & ~n18026;
  assign n18026 = ~n14511 & ~n22516;
  assign n19334 = ~n26335 & ~n26252;
  assign n26335 = n17222 | n17221;
  assign n16343 = n14836 ^ ~P3_IR_REG_30__SCAN_IN;
  assign n14836 = ~n20752 | ~P3_IR_REG_31__SCAN_IN;
  assign n20065 = n20066 ^ ~n14004;
  assign n20066 = ~n13763 | ~n13760;
  assign n25800 = n13867 ^ ~n25811;
  assign n13867 = ~n19969 | ~n19968;
  assign n22234 = ~n13601 | ~n13600;
  assign n19176 = n19174 & n13231;
  assign n18900 = n18899 & n22457;
  assign n13611 = ~n13609 | ~n13973;
  assign n14630 = n14631 & n17829;
  assign n18805 = ~n14112 | ~n15787;
  assign n21910 = ~n14374 | ~n13135;
  assign n22905 = n15637 & n15636;
  assign n21932 = ~n17734 | ~n17733;
  assign n22618 = ~n15609 | ~n15608;
  assign n15689 = n17346 | n17345;
  assign n22041 = ~n17621 | ~n17620;
  assign n15630 = ~n14163 | ~n14869;
  assign n13582 = ~n15486 | ~n15485;
  assign n23264 = ~n15058 | ~n15057;
  assign n15133 = n15125 ^ ~n15647;
  assign n18649 = ~n15285 | ~n15284;
  assign n21377 = ~n21058;
  assign n23818 = ~n14406 | ~n15185;
  assign n21309 = ~n21058;
  assign n24000 = ~n23254;
  assign n15647 = ~n15859;
  assign n23903 = ~n15099 | ~n15098;
  assign n25420 = ~n13182 | ~n17519;
  assign n13794 = n17948 | n15450;
  assign n24319 = n14949 | n16512;
  assign n15219 = n23124 & n14918;
  assign n15270 = ~n15243 | ~n15271;
  assign n23132 = ~n14914 | ~n23117;
  assign n18501 = n18854 | n23723;
  assign n17049 = ~n13773 | ~n13771;
  assign n23905 = ~n23723;
  assign n17036 = ~n15085;
  assign n13970 = n13969 & n15952;
  assign n13734 = ~n14114 | ~n13910;
  assign n18497 = ~n18142 | ~n18141;
  assign n18141 = n18065 & n13805;
  assign n22076 = ~n17878 | ~n14255;
  assign n22458 = n13626 ^ ~n13625;
  assign n22841 = n14261 ^ ~n18865;
  assign n14255 = n14390 & n13284;
  assign n20589 = ~n13698 | ~n13697;
  assign n13872 = n13952 & n13950;
  assign n13698 = n20582 | n20501;
  assign n20117 = ~n20110 & ~n20109;
  assign n20110 = ~n20082 & ~n20081;
  assign n18080 = ~n14755 | ~n13339;
  assign n14116 = n19082 ^ ~n19098;
  assign n19630 = ~n19185 & ~n19184;
  assign n18904 = ~n18903 | ~n13408;
  assign n13830 = ~n14167 | ~n14600;
  assign n13449 = ~n19008 | ~n19007;
  assign n21676 = ~n17663 | ~n17662;
  assign n22472 = ~n13119 | ~n14400;
  assign n23171 = ~n23174 | ~n17901;
  assign n14848 = ~n19003 | ~n14849;
  assign n23173 = ~n17903 | ~n17902;
  assign n13619 = ~n14037 | ~n14035;
  assign n19003 = ~n14126 | ~n13320;
  assign n21333 = ~n21487;
  assign n22174 = ~n13611 | ~n13610;
  assign n23114 = ~n14292 | ~n14290;
  assign n13668 = n13669 & n14630;
  assign n19095 = ~n15848 | ~n15847;
  assign n14398 = n14667 & n14399;
  assign n22132 = n17980 ^ ~n17979;
  assign n13671 = n13673 & n17826;
  assign n21487 = n17775 & n17774;
  assign n22632 = n14395 & n14392;
  assign n13787 = ~n20918 | ~n20917;
  assign n13503 = ~n13799 & ~n13504;
  assign n22832 = ~n18805;
  assign n14631 = ~n14632 | ~n21556;
  assign n13673 = n14622 | n13674;
  assign n14622 = n14623 & n21617;
  assign n26030 = ~n19996 | ~n19995;
  assign n23137 = ~n17955 | ~n15846;
  assign n20197 = ~n18322 | ~n18321;
  assign n22819 = ~n15812 | ~n15811;
  assign n26005 = n19827 ^ ~n19993;
  assign n19994 = ~n13861 | ~n13860;
  assign n22604 = ~n18050 | ~n18020;
  assign n21921 = ~n17745 | ~n17744;
  assign n13901 = n19289 | n13326;
  assign n22617 = n22633 | n22223;
  assign n22495 = ~n15757 | ~n15756;
  assign n18020 = n22905 | n13716;
  assign n21965 = ~n17694 | ~n17693;
  assign n20976 = ~n13454 | ~n13451;
  assign n21954 = ~n17708 | ~n17707;
  assign n21660 = n21975 ^ ~n21684;
  assign n22728 = ~n22746;
  assign n15637 = n17691 | n15810;
  assign n22862 = ~n15729 | ~n15728;
  assign n24950 = ~n14075 | ~n14074;
  assign n17423 = n15668 ^ ~P2_DATAO_REG_22__SCAN_IN;
  assign n17691 = n13714 ^ ~n15635;
  assign n15693 = ~n15689 | ~n15688;
  assign n17463 = ~n17375 | ~n17374;
  assign n22746 = n18044 & n18011;
  assign n13451 = n13452 & n18954;
  assign n14820 = ~n18189 | ~n14823;
  assign n21986 = ~n14383 | ~n17668;
  assign n21997 = ~n13886 | ~n17660;
  assign n20892 = n18976 | n18975;
  assign n22664 = ~n15558 | ~n15557;
  assign n13714 = ~n13715 | ~n15632;
  assign n17679 = n15629 ^ ~n15661;
  assign n17346 = n15717 ^ ~SI_22_;
  assign n22029 = ~n21037 | ~n21035;
  assign n20349 = ~n13448 | ~n18269;
  assign n14443 = n14444 & n17584;
  assign n23015 = ~n18041;
  assign n15629 = n14278 ^ ~SI_20_;
  assign n22295 = ~n15527 | ~n15526;
  assign n17664 = n15579 ^ ~n15600;
  assign n18041 = ~n15418 | ~n15417;
  assign n14828 = ~n14830 & ~n14829;
  assign n15660 = n15631 & n15630;
  assign n26182 = ~n18404 | ~n19338;
  assign n14446 = n14447 & n17577;
  assign n22018 = ~n17641 | ~n17640;
  assign n23203 = ~n15204 & ~n15203;
  assign n14163 = ~n14106 | ~n14107;
  assign n24982 = n25017 & n17851;
  assign n24473 = ~n17610 | ~n17609;
  assign n23740 = ~n22780 | ~n17399;
  assign n22341 = ~n15383 | ~n15382;
  assign n20209 = ~n26439;
  assign n24308 = ~n15737 | ~n15736;
  assign n24394 = ~n17603 | ~n17602;
  assign n23051 = ~n15323 | ~n15322;
  assign n25506 = ~n17593 | ~n17592;
  assign n23831 = n17363 & n17365;
  assign n13552 = n16543 & n16542;
  assign n15486 = ~n13889 | ~n13196;
  assign n25067 = n13202 & n13142;
  assign n24231 = ~n14653 | ~n15248;
  assign n13142 = n14431 & n25156;
  assign n25479 = ~n13666 | ~n17575;
  assign n13125 = ~n16548;
  assign n14499 = n15372 | n15405;
  assign n25882 = n19980 ^ ~n25893;
  assign n18877 = ~n23278 & ~n24190;
  assign n19980 = ~n13948 | ~n13323;
  assign n13666 = n25330 | n17704;
  assign n25454 = ~n17547 | ~n17546;
  assign n15372 = ~n13586 | ~n13584;
  assign n25240 = n17790 & n17484;
  assign n25330 = n15244 ^ ~n15270;
  assign n25150 = ~n13354 | ~n16733;
  assign n25114 = n25183 | n25420;
  assign n24976 = n16681 | n16680;
  assign n13196 = n13888 & n15448;
  assign n23872 = ~n24178;
  assign n23278 = ~n23875;
  assign n14032 = ~n17359 | ~n17358;
  assign n25689 = ~n26085;
  assign n26212 = ~n26343;
  assign n23753 = n15329 | n15328;
  assign n23825 = n15229 | n15228;
  assign n23853 = n15193 | n15192;
  assign n22790 = n15359 & n15358;
  assign n13583 = n14503 & n15339;
  assign n13888 = n14498 | n15406;
  assign n25021 = n16630 | n16629;
  assign n25049 = n16595 | n16594;
  assign n25126 = n16730 | n16729;
  assign n25432 = ~n17525 | ~n17524;
  assign n25252 = n16617 | n16616;
  assign n25254 = n16773 | n16772;
  assign n25274 = n16784 | n16785;
  assign n15640 = n15610 & P1_REG3_REG_19__SCAN_IN;
  assign n15046 = ~n15860;
  assign n15122 = n17520 | n15450;
  assign n23854 = n15110 | n15109;
  assign n14503 = ~n14103 | ~n13195;
  assign n17357 = n15032 | n15031;
  assign n14991 = n14986 & n14985;
  assign n17382 = ~n13615 | ~n13614;
  assign n23993 = ~n13482 | ~n13480;
  assign n26351 = n18167 | n18166;
  assign n26086 = n16479 | n16478;
  assign n26085 = n16399 | n16398;
  assign n26343 = n17232 | n17231;
  assign n26229 = n16456 | n16457;
  assign n26245 = ~n17212 | ~n17211;
  assign n16941 = n16939 & n16938;
  assign n15021 = n15020 & n15019;
  assign n15860 = ~n14949 | ~n18547;
  assign n13614 = n13616 & n14982;
  assign n13480 = n14917 & n13481;
  assign n25841 = n19975 ^ ~n25850;
  assign n14500 = n14501 & n15408;
  assign n25771 = ~n25751 & ~n25750;
  assign n14810 = n16467 | n16466;
  assign n18385 = ~n18387 & ~n19520;
  assign n15859 = ~n18547 | ~n18501;
  assign n26287 = n16437 | n16438;
  assign n26286 = n16488 | n16487;
  assign n25399 = ~n17497 | ~n17496;
  assign n19975 = ~n13877 | ~n19973;
  assign n14581 = n16314 | P3_ADDR_REG_5__SCAN_IN;
  assign n21356 = n16588 & n22139;
  assign n14109 = n15517 | n14110;
  assign n13915 = ~n14590 | ~n14589;
  assign n16939 = ~n16899 & ~P3_REG3_REG_21__SCAN_IN;
  assign n18547 = ~n18545;
  assign n22139 = ~n16587;
  assign n13129 = ~n14916;
  assign n15559 = ~n13178 & ~n15501;
  assign n16777 = ~n16588 | ~n16587;
  assign n16780 = n22133 & n16587;
  assign n18920 = ~n21395 | ~n17031;
  assign n13525 = ~n16240 | ~P3_ADDR_REG_4__SCAN_IN;
  assign n15036 = n15033 | n15069;
  assign n16460 = n20766 & n16343;
  assign n14175 = ~n21363 & ~n17657;
  assign n14430 = n14426 & n14425;
  assign n14930 = ~n14929 | ~P1_IR_REG_31__SCAN_IN;
  assign n16851 = ~n16501 & ~n13390;
  assign n19868 = ~n19847;
  assign n14100 = n15175 & n15206;
  assign n14935 = n15901 & n15870;
  assign n16484 = n16343 & n16345;
  assign n15033 = n15034 ^ ~SI_2_;
  assign n17502 = ~n24333 | ~n21363;
  assign n17657 = ~n24333;
  assign n15339 = n15313 | SI_11_;
  assign n22133 = n14438 ^ ~n22124;
  assign n25802 = n19809 ^ ~n25811;
  assign n15309 = ~n15276 | ~n15275;
  assign n19847 = n14703 & n14705;
  assign n18861 = ~n14937 | ~n14972;
  assign n24333 = ~n17049 | ~n24516;
  assign n20773 = ~n17182 | ~n13197;
  assign n15371 = n15342 | SI_12_;
  assign n15175 = n15176 ^ ~n18169;
  assign n14580 = ~n16110 | ~n16111;
  assign n15034 = ~n15008 | ~n15074;
  assign n19809 = ~n13992 | ~n19808;
  assign n23156 = ~n13121 & ~P1_STATE_REG_SCAN_IN;
  assign n15387 = n15354 | n22253;
  assign n16110 = ~n16108 | ~n16107;
  assign n18854 = n14146 ^ ~n14973;
  assign n17071 = n17013 & n17016;
  assign n20794 = n16001 ^ ~n15999;
  assign n15206 = n15207 ^ ~n15180;
  assign n15078 = ~n15081 & ~SI_3_;
  assign n15354 = n15353 | n15352;
  assign n13128 = n15037;
  assign n14938 = n14925 & n14701;
  assign n20752 = ~n17177 | ~n14835;
  assign n23723 = n14975 ^ ~P1_IR_REG_19__SCAN_IN;
  assign n17632 = n16878 & n15961;
  assign n16471 = ~n16425 & ~P3_REG3_REG_7__SCAN_IN;
  assign n19840 = n16090 & n19964;
  assign n17597 = ~n16564 & ~n17487;
  assign n15452 = ~n14890 | ~n14889;
  assign n16574 = n16573 & n16572;
  assign n14959 = ~n14958 & ~P3_ADDR_REG_19__SCAN_IN;
  assign n14960 = ~n14957 & ~P2_RD_REG_SCAN_IN;
  assign n14963 = ~n14961 & ~P1_ADDR_REG_19__SCAN_IN;
  assign n13537 = ~n15156 & ~n13538;
  assign n14922 = n14894 & n14893;
  assign n14890 = n15315 & n14886;
  assign n14889 = n14888 & n14887;
  assign n16074 = n23350 & P3_ADDR_REG_0__SCAN_IN;
  assign n15962 = ~P2_IR_REG_18__SCAN_IN & ~P2_IR_REG_16__SCAN_IN;
  assign n15963 = ~P2_IR_REG_17__SCAN_IN & ~P2_IR_REG_19__SCAN_IN;
  assign n15992 = ~P3_IR_REG_23__SCAN_IN & ~P3_IR_REG_22__SCAN_IN;
  assign n14891 = ~P1_IR_REG_16__SCAN_IN & ~P1_IR_REG_17__SCAN_IN;
  assign n14892 = ~P1_IR_REG_18__SCAN_IN & ~P1_IR_REG_15__SCAN_IN;
  assign n15991 = ~P3_IR_REG_16__SCAN_IN & ~P3_IR_REG_11__SCAN_IN;
  assign n14962 = ~P1_RD_REG_SCAN_IN & ~P2_ADDR_REG_19__SCAN_IN;
  assign n19806 = ~P3_IR_REG_0__SCAN_IN & ~P3_IR_REG_1__SCAN_IN;
  assign n15958 = ~P2_IR_REG_14__SCAN_IN & ~P2_IR_REG_13__SCAN_IN;
  assign n15990 = ~P3_IR_REG_19__SCAN_IN & ~P3_IR_REG_20__SCAN_IN;
  assign n15988 = ~P3_IR_REG_17__SCAN_IN & ~P3_IR_REG_14__SCAN_IN;
  assign n14887 = ~P1_IR_REG_12__SCAN_IN & ~P1_IR_REG_10__SCAN_IN;
  assign n14888 = ~P1_IR_REG_7__SCAN_IN & ~P1_IR_REG_11__SCAN_IN;
  assign n14886 = ~P1_IR_REG_14__SCAN_IN & ~P1_IR_REG_13__SCAN_IN;
  assign n14894 = ~P1_IR_REG_5__SCAN_IN & ~P1_IR_REG_3__SCAN_IN;
  assign n14893 = ~P1_IR_REG_4__SCAN_IN & ~P1_IR_REG_6__SCAN_IN;
  assign n15014 = ~P1_IR_REG_2__SCAN_IN;
  assign P2_U3088 = ~P2_STATE_REG_SCAN_IN;
  assign n15668 = n17346 | n13121;
  assign n15011 = n15012 & n15014;
  assign n17359 = n17357 | n23941;
  assign n13126 = ~n16809 | ~n13121;
  assign n13127 = ~n16809 | ~n13121;
  assign n15451 = ~n15379;
  assign n18512 = ~n14916;
  assign n15167 = n15860 | n14976;
  assign n15085 = n14964 & n14965;
  assign n13795 = ~n15036 | ~n15035;
  assign n15865 = n14930 ^ ~P1_IR_REG_26__SCAN_IN;
  assign n13130 = n15421;
  assign n13131 = n15421;
  assign n15421 = n14915 & n14918;
  assign n22817 = n22457 ^ n22450;
  assign n22450 = ~n14125 | ~n18058;
  assign n13132 = ~n15860;
  assign n21460 = n17873 & n13991;
  assign n17873 = ~n13136 & ~n21910;
  assign n18545 = ~n18861 & ~n18860;
  assign n14983 = ~n15024;
  assign n14087 = ~n13589 | ~n13289;
  assign n13589 = ~n13153 | ~n13590;
  assign n14444 = ~n14446 | ~n14445;
  assign n14445 = ~n17576;
  assign n14629 = ~n14630 | ~n21558;
  assign n14073 = ~n21841 | ~n14450;
  assign n14450 = ~n14455 & ~n14451;
  assign n14451 = ~n21431;
  assign n14455 = ~n17623;
  assign n14663 = n18891 & n14661;
  assign n13543 = n13238 & n18900;
  assign n17365 = n23853 | n23818;
  assign n15450 = ~n16809 | ~n17036;
  assign n13545 = n13546 & n15603;
  assign n14329 = ~n17033;
  assign n18627 = ~n18612 | ~n14162;
  assign n14162 = ~n23853 | ~n18829;
  assign n21219 = ~n14596 | ~n14594;
  assign n14594 = ~n14595 & ~n13206;
  assign n14596 = ~n17624 | ~n14598;
  assign n14609 = ~n21240 | ~n21239;
  assign n21240 = n21242 | n21241;
  assign n14565 = n20163 & n20184;
  assign n14837 = ~n14840 & ~n20406;
  assign n19479 = n20220 | n20235;
  assign n13939 = ~n14712 & ~n20442;
  assign n14710 = ~n14712 & ~n20424;
  assign n14823 = ~n26116 | ~n13581;
  assign n13781 = ~n13783;
  assign n14456 = ~n17500 & ~n14457;
  assign n14457 = ~n17485;
  assign n14148 = n14149 & n18813;
  assign n18549 = ~n18544 | ~n24122;
  assign n15719 = n15721 | SI_23_;
  assign n16106 = ~P1_ADDR_REG_2__SCAN_IN;
  assign n13651 = n13652 & n19144;
  assign n13652 = ~n19704;
  assign n20184 = n20197 ^ ~n26439;
  assign n18255 = n19427 | n19674;
  assign n14310 = n14311 & n17794;
  assign n14464 = ~n14088 | ~n14085;
  assign n14085 = n14086 & n14387;
  assign n14088 = ~n14466 | ~n14385;
  assign n14387 = n14388 & n21558;
  assign n13884 = ~n21661 | ~n17821;
  assign n13153 = n14279 & n13373;
  assign n14279 = ~n13158 | ~n14758;
  assign n14758 = ~n17677;
  assign n14640 = n13221 & n17820;
  assign n17814 = ~n21826 | ~n17812;
  assign n14074 = n14077 & n14765;
  assign n14765 = n14766 & n17585;
  assign n14448 = ~n17563;
  assign n24997 = n25479 ^ ~n24971;
  assign n17790 = n25274 | n25389;
  assign n14366 = n14875 & n15961;
  assign n14041 = ~n14785;
  assign n14665 = n14666 & n18057;
  assign n14770 = n14771 & n18036;
  assign n14772 = ~n18034;
  assign n14512 = ~n14513 | ~n22889;
  assign n14513 = ~n14514;
  assign n13623 = n18877 | n14783;
  assign n14783 = ~n17393;
  assign n18876 = ~n23278 | ~n24190;
  assign n14784 = ~n17391 | ~n13213;
  assign n14096 = n14372 & n15716;
  assign n15662 = n15664 | SI_21_;
  assign n15543 = ~n15542;
  assign n13420 = ~n17927 | ~n17928;
  assign n14338 = ~n25615 & ~n14339;
  assign n14339 = ~n19149;
  assign n19253 = ~n19251 & ~n20535;
  assign n17198 = ~n18191;
  assign n19222 = ~n13440 | ~n13439;
  assign n13439 = ~n13303 | ~n19494;
  assign n13440 = ~n13445 | ~n13441;
  assign n14745 = n18440 & n14746;
  assign n14746 = n18438 | n14747;
  assign n20478 = ~n18419 | ~n19397;
  assign n17152 = n17147 | P3_IR_REG_22__SCAN_IN;
  assign n14053 = n14054 & n17075;
  assign n14054 = ~n14056 | ~n14055;
  assign n14055 = ~n16950;
  assign n13434 = ~n14056 | ~n13435;
  assign n13435 = ~n16890;
  assign n13436 = ~n14056;
  assign n13703 = ~n16042;
  assign n17565 = ~P1_DATAO_REG_9__SCAN_IN;
  assign n14489 = ~n16145 | ~n14490;
  assign n14490 = n14491 & n14802;
  assign n14491 = ~n14805 | ~n16144;
  assign n16031 = ~P2_DATAO_REG_5__SCAN_IN;
  assign n14121 = ~n17041 | ~n17046;
  assign n21031 = ~n21402 | ~n17071;
  assign n13984 = ~n13985 & ~n21954;
  assign n13985 = ~n21598 | ~n13986;
  assign n21619 = ~n21965 & ~n21664;
  assign n21323 = ~n13539 | ~n17765;
  assign n13539 = n22150 | n17704;
  assign n14628 = n14629 & n17830;
  assign n21664 = ~n13987 | ~n13988;
  assign n13988 = ~n21975 & ~n21986;
  assign n21744 = ~n13679 | ~n13677;
  assign n13677 = ~n13678 & ~n13304;
  assign n13679 = ~n13675 | ~n21826;
  assign n14072 = ~n14073 | ~n14453;
  assign n14453 = n14454 & n17628;
  assign n13773 = n13777 & n13774;
  assign n13772 = n14084 & n16577;
  assign n17954 = n15841 | SI_28_;
  assign n17014 = ~P2_IR_REG_21__SCAN_IN;
  assign n13881 = ~SI_13_;
  assign n18901 = n18843 ^ ~n24330;
  assign n13721 = ~n23493 | ~n23492;
  assign n13599 = ~n22548 & ~n22862;
  assign n14781 = n22585 & n18021;
  assign n14393 = ~n18048;
  assign n22223 = ~n15583 | ~n15582;
  assign n14395 = ~n13500 | ~n13916;
  assign n13916 = ~n13307 & ~n13917;
  assign n13917 = ~n18892;
  assign n18046 = n22702 | n22999;
  assign n17366 = ~n23829 | ~n17364;
  assign n22457 = ~n18059 | ~n18037;
  assign n23991 = n17404 & n17403;
  assign n14419 = ~n14420 | ~n15904;
  assign n15546 = n15521 | SI_17_;
  assign n16095 = ~n13561 | ~n16074;
  assign n13653 = n13654 & n14187;
  assign n14187 = n14188 & n19596;
  assign n25995 = ~n14270 | ~n14269;
  assign n14269 = ~n25996;
  assign n18351 = n19228;
  assign n19228 = ~n18191 | ~n21363;
  assign n16789 = ~n14808 | ~n16052;
  assign n13705 = ~n17533 | ~P2_DATAO_REG_6__SCAN_IN;
  assign n17058 = ~n17862 & ~n17010;
  assign n13824 = n13825 & n21407;
  assign n13825 = ~n13828 | ~n13830;
  assign n16878 = n15960 & n17597;
  assign n16587 = n16584 & n16583;
  assign n17961 = ~n17955 | ~n17954;
  assign n17955 = ~n14306 | ~n14164;
  assign n14164 = n15843 & n15838;
  assign n15418 = n24052 | n15450;
  assign n13973 = ~n22332;
  assign n13609 = ~n13976 | ~n13974;
  assign n15553 = ~n16809;
  assign n18865 = n18805 ^ ~n14111;
  assign n14297 = n17975 | n14298;
  assign n13889 = ~n15372 | ~n14497;
  assign n15448 = ~n15447 & ~n15446;
  assign n13809 = ~P2_ADDR_REG_7__SCAN_IN;
  assign n13810 = ~n16928;
  assign n23189 = ~n23192 | ~n17939;
  assign n14603 = n13399 | n21458;
  assign n16548 = ~n13484 | ~n13483;
  assign n13483 = ~n13485 | ~n16836;
  assign n13484 = ~n13486 | ~P1_ADDR_REG_6__SCAN_IN;
  assign n13485 = n16546 & n16547;
  assign n17881 = ~n17318 | ~n17317;
  assign n19314 = ~n26287 | ~n14005;
  assign n14556 = ~n19333;
  assign n21071 = n21060 & n21059;
  assign n14012 = n19326 & n14553;
  assign n14027 = ~n13185 | ~n19354;
  assign n13817 = ~n13818 | ~n21141;
  assign n14025 = ~n13139 & ~n13273;
  assign n14599 = ~n21035 | ~n17704;
  assign n14141 = n14142 & n18654;
  assign n21218 = n21046 & n21045;
  assign n19452 = ~n14797 | ~n14796;
  assign n14796 = ~n13227 & ~n13168;
  assign n13469 = n18712 & n13467;
  assign n13905 = ~n26160 & ~n13906;
  assign n14607 = ~n14606 & ~n21249;
  assign n18535 = n22905 | n13123;
  assign n18537 = n22905 | n18779;
  assign n14154 = n14155 & n18755;
  assign n13902 = ~n20362;
  assign n13940 = ~n14723 & ~n13942;
  assign n14360 = n21275 & n21286;
  assign n13834 = ~n13835 | ~n13271;
  assign n13833 = ~n13835;
  assign n21328 = n21326 | n21327;
  assign n21437 = n21435 & n13410;
  assign n13410 = n21743 & n21758;
  assign n14460 = ~n14463 & ~n21556;
  assign n18881 = n18880 & n13693;
  assign n13687 = n22694 & n13688;
  assign n13688 = ~n22723 & ~n13689;
  assign n13689 = ~n22771;
  assign n18279 = n18275 | n20283;
  assign n19460 = n18431 & n20334;
  assign n14853 = n26199 & n13180;
  assign n19315 = n14810 & n26277;
  assign n19312 = ~n14810 & ~n26277;
  assign n15983 = ~P3_IR_REG_9__SCAN_IN & ~P3_IR_REG_5__SCAN_IN;
  assign n14089 = ~n21676 | ~n13234;
  assign n13158 = ~n14760 & ~n21660;
  assign n14760 = ~n17678;
  assign n14183 = ~n14639;
  assign n14316 = n14317 & n17806;
  assign n14318 = ~n17804;
  assign n14768 = ~n17531;
  assign n19248 = ~n19238 & ~n19237;
  assign n13903 = ~n13236 | ~n20184;
  assign n13862 = ~n13864 | ~n25982;
  assign n13759 = n20038 & P3_REG1_REG_15__SCAN_IN;
  assign n20108 = ~n20074 | ~n13394;
  assign n13441 = n14742 & n19494;
  assign n14832 = ~n14227 | ~n14224;
  assign n14224 = ~n14225 & ~n13290;
  assign n13446 = ~n13922 | ~n13924;
  assign n13922 = n13332 & n13923;
  assign n18302 = n20228 & n18303;
  assign n14750 = ~n20330 & ~n14751;
  assign n14751 = ~n18428;
  assign n14842 = n18262 & n18255;
  assign n13576 = ~n14212 | ~n13211;
  assign n13577 = ~n18226 & ~n13283;
  assign n20374 = ~n20372 | ~n20385;
  assign n14216 = n13306 & n14217;
  assign n14218 = ~n18225;
  assign n14841 = ~n19424;
  assign n14202 = n14203 & n18414;
  assign n18202 = n26393 | n25689;
  assign n14821 = ~n13566 | ~n13300;
  assign n13566 = n14822 | n19363;
  assign n14822 = ~n14823;
  assign n18189 = n26130 & n14220;
  assign n14220 = n14221 & n18181;
  assign n19335 = n26252 & n26335;
  assign n19327 = ~n18158 | ~n25707;
  assign n17140 = n15997 & n16013;
  assign n14487 = ~n14878;
  assign n14480 = n14481 & n16323;
  assign n14302 = ~n24401;
  assign n14812 = ~n20973;
  assign n14286 = ~n19018;
  assign n14287 = n20879 & n14288;
  assign n14611 = ~n14614 | ~n13222;
  assign n14267 = ~n21450 | ~n13285;
  assign n13813 = n13815 & n13814;
  assign n14171 = ~n21058 & ~n14172;
  assign n21446 = ~n21443 & ~n14378;
  assign n14642 = n21997 ^ ~n13885;
  assign n17486 = ~P1_DATAO_REG_2__SCAN_IN;
  assign n14755 = ~n13780 | ~n13175;
  assign n14756 = ~n17773;
  assign n14374 = n14375 & n17755;
  assign n14375 = n15786 | n17704;
  assign n14623 = ~n14624 | ~n17824;
  assign n14624 = ~n17823;
  assign n14639 = ~n14642 | ~n17818;
  assign n14180 = ~n14182 & ~n14181;
  assign n14181 = ~n17817;
  assign n17678 = n21986 | n21709;
  assign n21681 = ~n14641 | ~n17820;
  assign n17816 = n22029 | n21818;
  assign n14643 = ~n21789 & ~n14646;
  assign n14646 = ~n17813;
  assign n14764 = ~n21430;
  assign n21868 = ~n14319 | ~n14316;
  assign n14637 = ~n17801;
  assign n17564 = ~n25028 | ~n17562;
  assign n25076 = ~n25083;
  assign n25135 = n25399 | n25252;
  assign n25155 = ~n14433 | ~n14432;
  assign n14432 = ~n25399;
  assign n14433 = ~n25206;
  assign n17508 = ~n17501 | ~n14458;
  assign n13836 = n14139 & n15961;
  assign n18899 = n18895 & n13690;
  assign n13690 = ~n18898 & ~n13691;
  assign n15697 = ~n15640 | ~n13405;
  assign n14043 = ~n18029 & ~n18027;
  assign n18021 = ~n22905 | ~n24298;
  assign n18045 = ~n22729 | ~n22746;
  assign n13636 = ~n18887 | ~n18008;
  assign n14657 = ~n23772 | ~n23776;
  assign n14123 = ~n22457 & ~n14124;
  assign n14124 = ~n18058;
  assign n14400 = ~n13712 | ~n14398;
  assign n14402 = ~n18054;
  assign n13800 = ~n22585 | ~n18052;
  assign n13801 = ~n18049;
  assign n13502 = n13146 & n22625;
  assign n14785 = n13201 & n18014;
  assign n23772 = ~n23777;
  assign n17389 = ~n17388 & ~n14874;
  assign n13629 = ~n24015 | ~n17352;
  assign n15751 = ~n14136 | ~n15748;
  assign n14136 = ~n15724 | ~n14135;
  assign n14135 = ~n13169 & ~SI_24_;
  assign n15805 = n15754 | SI_25_;
  assign n14700 = n14701 & n13319;
  assign n13548 = ~n14493 & ~n15516;
  assign n14493 = ~n15543 | ~n15601;
  assign n14498 = ~n14500 | ~n13219;
  assign n14958 = ~P2_ADDR_REG_19__SCAN_IN;
  assign n14957 = ~P1_ADDR_REG_19__SCAN_IN;
  assign n16094 = ~n16093 | ~P3_ADDR_REG_1__SCAN_IN;
  assign n16093 = ~P1_ADDR_REG_1__SCAN_IN;
  assign n14573 = ~n16106 | ~n14576;
  assign n16314 = ~n14254 | ~n13525;
  assign n13424 = n17942 | n17943;
  assign n17942 = ~n17941 & ~n17940;
  assign n19493 = ~n14256 | ~n26445;
  assign n19494 = ~n20165 | ~n20160;
  assign n14331 = ~n19141 | ~n14534;
  assign n14190 = ~n14191 | ~n14334;
  assign n14334 = ~n14337 & ~n14335;
  assign n14336 = ~n19579 | ~n19446;
  assign n13648 = ~n13651;
  assign n14002 = ~n19807;
  assign n19813 = ~n13993 | ~n19812;
  assign n14234 = n25934 | n25931;
  assign n14241 = ~n19942 | ~n14242;
  assign n14242 = ~n19946;
  assign n14240 = ~n20010;
  assign n18366 = ~n13843 | ~n13842;
  assign n13842 = ~P3_REG3_REG_27__SCAN_IN;
  assign n20152 = P3_REG3_REG_28__SCAN_IN ^ ~n18366;
  assign n13843 = ~n18339 & ~P3_REG3_REG_26__SCAN_IN;
  assign n18339 = ~n13845 | ~n13844;
  assign n13844 = ~P3_REG3_REG_25__SCAN_IN;
  assign n18323 = ~n13845;
  assign n20261 = n20593 | n20267;
  assign n16414 = ~n13851;
  assign n26200 = ~n18161 | ~n18160;
  assign n19257 = ~n20119;
  assign n26282 = ~n20501;
  assign n18455 = n19522 & n20119;
  assign n20129 = ~n26455;
  assign n20185 = ~n18437 | ~n19480;
  assign n18437 = ~n13447 | ~n13930;
  assign n13930 = ~n13932 & ~n13931;
  assign n13447 = ~n13446 | ~n13232;
  assign n20333 = ~n14753 | ~n14750;
  assign n14713 = ~n20424 | ~n19417;
  assign n13921 = ~n18416 | ~n18415;
  assign n14736 = ~n13207 | ~n14734;
  assign n18411 = ~n14868 & ~n18410;
  assign n14868 = ~n26076 & ~n18409;
  assign n19346 = ~n26205 | ~n26351;
  assign n14732 = ~n14731 | ~n19345;
  assign n14731 = ~n26182;
  assign n26258 = ~n19327 | ~n19329;
  assign n18448 = ~n13637 | ~n17135;
  assign n13637 = ~n14528 | ~n14530;
  assign n13642 = ~P3_IR_REG_25__SCAN_IN & ~P3_IR_REG_24__SCAN_IN;
  assign n18306 = ~n18297 | ~n18296;
  assign n18291 = ~n14469 | ~n17457;
  assign n14469 = ~n14071 | ~n13395;
  assign n18443 = ~n17153 | ~n17152;
  assign n17143 = ~P3_IR_REG_21__SCAN_IN;
  assign n17147 = ~n17140 | ~n17143;
  assign n14488 = ~n17270 | ~n17269;
  assign n14808 = ~n16050 | ~n16051;
  assign n14066 = n13144 & n16040;
  assign n14070 = ~n16203;
  assign n16024 = ~P2_DATAO_REG_3__SCAN_IN;
  assign n17039 = n25274 & n24449;
  assign n14860 = ~n18923 & ~n18922;
  assign n17589 = ~P1_DATAO_REG_11__SCAN_IN;
  assign n14863 = ~n24410 | ~n24411;
  assign n21037 = ~n17624 | ~n21352;
  assign n16661 = n16701 | n16604;
  assign n24927 = ~n13897 | ~n24901;
  assign n13991 = ~n21333 & ~n21323;
  assign n21886 = ~n24982 | ~n17852;
  assign n25025 = ~n17799 | ~n17798;
  assign n25083 = n17793 & n25045;
  assign n21395 = ~n21407 | ~n17071;
  assign n21345 = ~n18082 | ~n18081;
  assign n21445 = n21323 ^ ~n19051;
  assign n21409 = ~n14373 | ~n13135;
  assign n14373 = n14374 & n25577;
  assign n13591 = ~n14464 | ~n13592;
  assign n13592 = ~n13594 & ~n14462;
  assign n14632 = ~n17827;
  assign n17745 = n22163 | n17704;
  assign n17708 = n17705 | n17704;
  assign n21772 = ~n21802 & ~n22029;
  assign n21826 = ~n17811 | ~n17810;
  assign n21841 = ~n17604 | ~n21414;
  assign n24947 = n17805 & n17806;
  assign n25017 = n17850 & n25067;
  assign n17863 = ~n25509 & ~n17071;
  assign n15955 = ~P2_IR_REG_6__SCAN_IN & ~P2_IR_REG_8__SCAN_IN;
  assign n16569 = ~P2_IR_REG_25__SCAN_IN & ~P2_IR_REG_24__SCAN_IN;
  assign n14084 = ~n13900 & ~n16575;
  assign n15968 = n15965 | n17032;
  assign n15965 = ~n15979 & ~P2_IR_REG_24__SCAN_IN;
  assign n15970 = ~n15968 | ~n15966;
  assign n15966 = ~P2_IR_REG_25__SCAN_IN;
  assign n15979 = n15974 | P2_IR_REG_23__SCAN_IN;
  assign n14363 = n14364 & n17014;
  assign n14365 = n16878 | n17032;
  assign n13604 = ~n15599;
  assign n23266 = ~n23874;
  assign n15628 = n15623 | n15624;
  assign n14997 = n14994 ^ ~n15859;
  assign n15585 = ~n15559 | ~P1_REG3_REG_17__SCAN_IN;
  assign n15931 = n17442 | n15903;
  assign n13473 = n13474 & n18816;
  assign n14157 = ~n14158 & ~n18841;
  assign n13544 = ~n18060 & ~n19081;
  assign n13733 = ~n23431 | ~n23430;
  assign n19084 = ~n13596 | ~n13595;
  assign n13595 = n13597 & n22535;
  assign n13597 = n14523 & n13598;
  assign n14523 = ~n14524 & ~n19095;
  assign n14524 = ~n22832 | ~n14525;
  assign n22494 = n13599 & n13598;
  assign n14514 = ~n22905 | ~n14515;
  assign n22570 = ~n22617 & ~n14512;
  assign n14779 = ~n18021;
  assign n18018 = n18896 & n22624;
  assign n15609 = n17679 | n15810;
  assign n18896 = n22618 ^ ~n24295;
  assign n14392 = ~n22629 & ~n14394;
  assign n14394 = ~n18047;
  assign n22678 = ~n22705 & ~n22295;
  assign n14777 = ~n18882;
  assign n14520 = ~n13154 | ~n22257;
  assign n17375 = ~n13492 | ~n17373;
  assign n23749 = n23765 & n13914;
  assign n24178 = ~n15122 | ~n15121;
  assign n18843 = ~n17972 | ~n17971;
  assign n15812 = n22150 | n15810;
  assign n13625 = ~n22457;
  assign n13626 = ~n13627 | ~n14770;
  assign n13627 = ~n13628 | ~n14505;
  assign n14510 = ~n14512 & ~n14511;
  assign n22522 = ~n22543 | ~n18028;
  assign n23765 = ~n23820 & ~n24213;
  assign n23851 = ~n18877 & ~n13685;
  assign n13495 = n23926 | n13498;
  assign n13496 = ~n13497 & ~n13270;
  assign n14298 = ~n14299 | ~n17966;
  assign n14299 = ~n17970;
  assign n13462 = n14904 & n14790;
  assign n15806 = ~n13534 | ~n15751;
  assign n13534 = n15750 & n15828;
  assign n15784 = ~n15806 | ~n15805;
  assign n15749 = ~n14095 | ~n14097;
  assign n14097 = ~n13272 & ~n13169;
  assign n14095 = ~n14096 | ~n15630;
  assign n14372 = n15631 & n15659;
  assign n14924 = ~P1_IR_REG_19__SCAN_IN;
  assign n15577 = ~n15575 | ~n15576;
  assign n13879 = n15543 & n15517;
  assign n14496 = ~n15543 | ~n14110;
  assign n14497 = ~n14498;
  assign n15485 = n15438 | SI_15_;
  assign n15315 = ~P1_IR_REG_8__SCAN_IN & ~P1_IR_REG_9__SCAN_IN;
  assign n15069 = ~n15077;
  assign n13508 = n16319 & n16247;
  assign n13523 = ~n14581;
  assign n14582 = ~n16314 | ~P3_ADDR_REG_5__SCAN_IN;
  assign n14586 = n17313 & n13713;
  assign n17918 = ~n13430 | ~n13427;
  assign n13427 = n13428 & n17914;
  assign n19061 = n13424 ^ ~P1_ADDR_REG_17__SCAN_IN;
  assign n14538 = ~n25697 | ~n19153;
  assign n20141 = ~n19493 | ~n19494;
  assign n14184 = ~n14540 | ~n13331;
  assign n14185 = ~n19532;
  assign n25638 = ~n26116;
  assign n25660 = n13639 & n17205;
  assign n20495 = ~n19552;
  assign n19750 = ~n19176 & ~n19175;
  assign n19766 = n19170 | n19674;
  assign n14470 = n14471 & n19522;
  assign n14471 = ~n14473 | ~n14472;
  assign n14715 = ~n19264 & ~n13237;
  assign n19300 = ~n19299 & ~n19298;
  assign n14717 = n19222 | n14718;
  assign n14718 = ~n19268 | ~n14719;
  assign n14719 = ~n19221;
  assign n18326 = ~n16460;
  assign n14003 = ~n19840 | ~n25742;
  assign n13875 = ~n19840 | ~n13966;
  assign n13966 = ~n25746;
  assign n14237 = n25848 | n25846;
  assign n19990 = ~n13859 | ~n19988;
  assign n13859 = ~n13857 | ~n13855;
  assign n13855 = n13856 & n25946;
  assign n19827 = ~n13994 | ~n19826;
  assign n26046 = ~n14238 | ~n13393;
  assign n14238 = ~n25995 | ~n14239;
  assign n14239 = n26011 & n19927;
  assign n20034 = n16894 & n16893;
  assign n20006 = n20007 ^ ~n19999;
  assign n20097 = ~n13866 | ~P3_REG2_REG_17__SCAN_IN;
  assign n13955 = ~n13956 | ~n20103;
  assign n13956 = ~n20101;
  assign n13951 = n13959 | n13957;
  assign n13960 = ~n20097;
  assign n18492 = ~P3_REG3_REG_28__SCAN_IN & ~n18366;
  assign n20174 = ~n14468 | ~n18338;
  assign n14468 = n20779 | n18351;
  assign n18321 = n18176 | n20787;
  assign n18322 = n20785 | n18351;
  assign n26150 = n18173 | n18172;
  assign n20528 = ~n26152;
  assign n26303 = n18455 & n19834;
  assign n18482 = n17101 & n26310;
  assign n17101 = n17134 | P3_D_REG_1__SCAN_IN;
  assign n16338 = ~P3_IR_REG_29__SCAN_IN;
  assign n14044 = ~n19227 | ~n19226;
  assign n17177 = n13575 & n15997;
  assign n13575 = n15996 & n13313;
  assign n14045 = ~n18350 | ~n18349;
  assign n17299 = n17300 ^ ~P1_DATAO_REG_20__SCAN_IN;
  assign n14056 = n14057 & n16952;
  assign n14058 = ~n16057;
  assign n14059 = ~n16058;
  assign n14807 = ~n14808;
  assign n13704 = ~n16043;
  assign n16117 = ~n13705 | ~n16035;
  assign n14792 = ~n14794 & ~n14793;
  assign n21586 = ~n25565;
  assign n14825 = ~n14826 | ~n18950;
  assign n14843 = n14844 & n19032;
  assign n14425 = n24333 | n14424;
  assign n18915 = n17039 | n17040;
  assign n14120 = ~n14121;
  assign n17046 = n24452 & n17045;
  assign n20863 = n19005 | n19004;
  assign n14126 = ~n13459 | ~n14127;
  assign n24389 = ~n21817;
  assign n17525 = n17520 | n17704;
  assign n21845 = ~n24955;
  assign n21560 = ~n25574;
  assign n24471 = n17069 | n17028;
  assign n13829 = ~n13830;
  assign n24521 = ~n24336 | ~n24335;
  assign n21462 = ~n21355 | ~n21354;
  assign n14168 = ~n14175;
  assign n17694 = n17691 | n17704;
  assign n17682 = n17679 | n17704;
  assign n16674 = ~n16686 & ~n16603;
  assign n16590 = P2_REG3_REG_6__SCAN_IN & P2_REG3_REG_7__SCAN_IN;
  assign n18106 = ~n25374 & ~n17007;
  assign n18105 = n17862 | n17861;
  assign n14816 = ~n24454;
  assign n22124 = ~P2_IR_REG_30__SCAN_IN;
  assign n14306 = ~n14307 | ~n15836;
  assign n15836 = n15835 | n15834;
  assign n15843 = n17954 & n15842;
  assign n25194 = n17026 & n13188;
  assign n15273 = ~n15270 & ~n15269;
  assign n13661 = n15239 & n15177;
  assign n15269 = n15210 | SI_8_;
  assign n14406 = n25342 | n15810;
  assign n13610 = ~n22171;
  assign n22187 = n15712 ^ ~n15710;
  assign n13978 = n14691 & n13979;
  assign n14691 = ~n13209 | ~n13145;
  assign n14678 = n14679 & n17996;
  assign n14679 = ~n17995 | ~n14680;
  assign n14689 = ~n14690 | ~n15307;
  assign n22702 = ~n15500 | ~n15499;
  assign n15500 = n25302 | n15810;
  assign n15930 = n14949 & n15928;
  assign n14690 = ~n22371;
  assign n22515 = n15765 & n15764;
  assign n15936 = n15219;
  assign n13616 = ~n13129 | ~P1_REG0_REG_1__SCAN_IN;
  assign n13481 = ~n18512 | ~P1_REG0_REG_0__SCAN_IN;
  assign n13725 = ~n23554;
  assign n23552 = ~n23542 & ~n23543;
  assign n23623 = n14247 & n14246;
  assign n14246 = ~n23598;
  assign n23655 = ~n13729 & ~n23631;
  assign n13729 = ~n23629 & ~n23630;
  assign n23706 = ~n13727 | ~n23702;
  assign n22421 = ~n17982 | ~n17981;
  assign n17982 = n22132 | n15810;
  assign n22422 = ~n19084 & ~n19085;
  assign n22452 = ~n24320;
  assign n22429 = n19084 ^ ~n14526;
  assign n18070 = n15939 ^ ~n13541;
  assign n13541 = ~P1_REG3_REG_28__SCAN_IN;
  assign n15757 = n22163 | n15810;
  assign n14035 = n14036 & n18016;
  assign n22952 = ~n22664;
  assign n14271 = n22725;
  assign n24015 = ~n17382;
  assign n22414 = ~n18843;
  assign n22810 = ~n22421;
  assign n18135 = n13796 ^ ~n18864;
  assign n14653 = ~n14655 | ~n14654;
  assign n24034 = ~n15865 | ~n15869;
  assign n24033 = ~n14949 | ~n16511;
  assign n14300 = ~n17962;
  assign n14293 = n14296 & n14294;
  assign n14294 = ~n17970 | ~n14295;
  assign n14296 = n13387 | n14298;
  assign n14295 = ~n17966;
  assign n17975 = ~n17961 | ~n17960;
  assign n14146 = ~n13295 | ~n14147;
  assign n14587 = ~n15440 | ~n14176;
  assign n14176 = ~n14499 | ~n13293;
  assign n16101 = n13908 ^ ~P1_ADDR_REG_2__SCAN_IN;
  assign n13486 = ~n16836 | ~n16546;
  assign n17315 = ~n17310 | ~n17309;
  assign n23164 = ~n23167 | ~n17888;
  assign n17924 = ~n13711 | ~n23178;
  assign n13516 = ~n13531 | ~n13517;
  assign n13518 = ~n13527;
  assign n13517 = ~n19066;
  assign n20656 = ~n18223 | ~n18222;
  assign n18223 = n18219 | n18351;
  assign n26138 = ~n26189;
  assign n18436 = ~n20801 | ~n18258;
  assign n20665 = ~n18216 | ~n18215;
  assign n18216 = n18212 | n18351;
  assign n20648 = ~n18232 | ~n18231;
  assign n25964 = n19990 ^ ~n19989;
  assign n18253 = n18248 | n18351;
  assign n26297 = ~n26224;
  assign n25093 = ~n25022;
  assign n14602 = ~n14603;
  assign n14327 = n14328 & n16580;
  assign n21456 = ~n17071;
  assign n14112 = ~n23149 | ~n14654;
  assign n23331 = ~n23277;
  assign n14414 = n13684 & n18905;
  assign n13684 = ~n18904 | ~n13408;
  assign n14105 = ~n14414 | ~n14412;
  assign n14412 = ~n18904;
  assign n23493 = ~n14243 | ~n23485;
  assign n14243 = ~n14245 | ~n14244;
  assign n14244 = ~n23482;
  assign n23729 = n16817 & n16815;
  assign n13553 = ~n13552;
  assign n13551 = ~n13552 | ~n13412;
  assign n13412 = ~n13125 | ~n13511;
  assign n23166 = ~n17891 | ~n17890;
  assign n23192 = ~n13513 | ~n13512;
  assign n19313 = ~n19314;
  assign n19333 = ~n19332 & ~n19331;
  assign n21070 = ~n21063 | ~n21062;
  assign n13471 = ~n13472 | ~n13329;
  assign n21090 = ~n25420;
  assign n14368 = n21085 & n21080;
  assign n14410 = ~n18576 & ~n14411;
  assign n14411 = ~n18574;
  assign n14026 = n14027 & n13189;
  assign n14548 = n13223 & n26081;
  assign n18626 = ~n18627;
  assign n14595 = ~n14597 & ~n21035;
  assign n21168 = n13316 & n21169;
  assign n14567 = n19404 & n19410;
  assign n13466 = ~n14140 | ~n13251;
  assign n13464 = n13465 & n18692;
  assign n14798 = ~n14799 & ~n19834;
  assign n14799 = ~n18261;
  assign n19450 = ~n19439 & ~n19438;
  assign n13822 = ~n21230;
  assign n13821 = n21218 & n21229;
  assign n14561 = n19465 & n14791;
  assign n14791 = ~n20292;
  assign n14417 = ~n18730;
  assign n14021 = n14561 & n13190;
  assign n14153 = ~n18754;
  assign n21259 = n21252 & n21251;
  assign n19288 = n19286 & n13904;
  assign n13904 = ~n19287 & ~n13942;
  assign n13411 = n21428 & n21429;
  assign n13478 = ~n13205 | ~n13151;
  assign n13693 = ~n23772 & ~n13694;
  assign n13694 = ~n23740 | ~n13695;
  assign n13695 = ~n14031 & ~n13696;
  assign n14563 = n14564 & n19491;
  assign n14382 = ~n21585;
  assign n13590 = ~n13158 & ~n21411;
  assign n14321 = n14322 & n17805;
  assign n14323 = ~n17803;
  assign n19160 = n19161 | n19644;
  assign n14226 = ~n18317;
  assign n14223 = n18331 & n20205;
  assign n14833 = ~n18332;
  assign n14749 = ~n14884;
  assign n13927 = ~n18424 & ~n13928;
  assign n13926 = ~n14750;
  assign n14214 = ~n18233;
  assign n14215 = ~n14837;
  assign n14212 = ~n14837 | ~n14213;
  assign n14213 = ~n14216;
  assign n14727 = ~n14729 | ~n20461;
  assign n14729 = ~n14730 | ~n19400;
  assign n14730 = ~n19401;
  assign n13569 = ~n13570 & ~n13573;
  assign n13573 = ~n18217;
  assign n13570 = ~n18418;
  assign n13571 = ~n13572 | ~n18217;
  assign n13572 = ~n18417;
  assign n14206 = ~n18202 & ~n14207;
  assign n14207 = ~n18413;
  assign n14813 = ~n24467;
  assign n13832 = ~n13833 | ~n13298;
  assign n14361 = n21291 & n14362;
  assign n14877 = ~n13838 | ~n25194;
  assign n13838 = ~n21395 & ~n21402;
  assign n14614 = ~n14615 | ~n21320;
  assign n14358 = ~n13208 | ~n21303;
  assign n21365 = n21034 & n21392;
  assign n14172 = ~n14175 & ~n14174;
  assign n21441 = ~n21440 & ~n21660;
  assign n21440 = n21639 | n21439;
  assign n14378 = ~n21444 | ~n14379;
  assign n14379 = ~n21540 & ~n14380;
  assign n14380 = ~n14382 | ~n14381;
  assign n14381 = ~n21617;
  assign n14461 = ~n17754 | ~n14462;
  assign n13549 = ~n14757 & ~n21445;
  assign n14757 = ~n21409;
  assign n14388 = ~n13785 | ~n17731;
  assign n14466 = ~n14089;
  assign n14385 = ~n13786 & ~n14386;
  assign n14386 = ~n17717;
  assign n14644 = ~n17816;
  assign n14766 = ~n24947;
  assign n14077 = ~n14443 | ~n14078;
  assign n14078 = ~n14446;
  assign n14459 = ~n25245 | ~n25244;
  assign n13778 = ~P2_IR_REG_28__SCAN_IN | ~P2_IR_REG_31__SCAN_IN;
  assign n18893 = ~n18890 & ~n13686;
  assign n13686 = ~n22629 | ~n13687;
  assign n13691 = ~n22544 | ~n13692;
  assign n13692 = ~n18897 & ~n14658;
  assign n14667 = n22491 & n18056;
  assign n14659 = ~n18013;
  assign n14660 = n18046 & n18044;
  assign n17400 = n23740 & n23739;
  assign n14572 = n16094 & n16106;
  assign n19177 = ~n19176;
  assign n14534 = ~n14535;
  assign n14189 = ~n14882;
  assign n14335 = ~n19766;
  assign n14800 = n19507 & n19512;
  assign n13947 = ~n19976;
  assign n13770 = ~P3_REG1_REG_7__SCAN_IN;
  assign n13845 = ~n17091 & ~P3_REG3_REG_24__SCAN_IN;
  assign n13840 = ~n16528 | ~n13841;
  assign n13841 = ~P3_REG3_REG_16__SCAN_IN;
  assign n13851 = ~n13177 & ~n13846;
  assign n13846 = ~n13847 | ~n16363;
  assign n13847 = ~n13848;
  assign n19364 = n18443 | n19306;
  assign n13445 = ~n20185;
  assign n13932 = ~n13933 & ~n19270;
  assign n13931 = ~n19479;
  assign n13933 = ~n18435 & ~n19271;
  assign n20208 = n19479 & n19480;
  assign n18283 = n18282 | n18281;
  assign n20282 = n20330 & n14881;
  assign n13707 = ~n13936 | ~n13935;
  assign n13936 = n13937 & n14708;
  assign n14723 = ~n14725 & ~n14724;
  assign n14724 = ~n19405;
  assign n14725 = ~n14727 & ~n19400;
  assign n14722 = ~n20478 | ~n14726;
  assign n14726 = ~n14727;
  assign n14734 = ~n14737 | ~n20524;
  assign n14819 = ~n14821 & ~n26053;
  assign n14854 = ~n14855 | ~n13180;
  assign n19338 = ~n25624 | ~n26212;
  assign n14200 = ~n26256;
  assign n14705 = ~n14706 | ~n13347;
  assign n14703 = ~n14704 & ~n13315;
  assign n18297 = ~n18291 | ~n18290;
  assign n16954 = n16011 | n16010;
  assign n15987 = ~n15985 & ~n15984;
  assign n14802 = ~n16036 & ~n14803;
  assign n14803 = ~n13705;
  assign n13452 = n14825 | n13453;
  assign n14313 = ~n25432 & ~n14314;
  assign n21444 = ~n18113;
  assign n13674 = ~n17825;
  assign n17734 = n17732 | n17704;
  assign n14619 = ~n14625 & ~n14620;
  assign n14620 = ~n17822;
  assign n14625 = ~n17824;
  assign n14465 = ~n14087;
  assign n13675 = ~n13203 & ~n13676;
  assign n13676 = ~n17812;
  assign n13678 = ~n14643 & ~n13203;
  assign n14454 = ~n14763 | ~n17623;
  assign n13682 = n17807 | n13683;
  assign n14440 = ~n14441 | ~n17539;
  assign n14441 = n14768 | n25083;
  assign n25045 = ~n13779 | ~n13983;
  assign n25120 = ~n14079 | ~n25420;
  assign n14617 = ~n25219 | ~n17791;
  assign n25209 = ~n14459 | ~n17485;
  assign n14081 = n14083 & n14080;
  assign n14083 = ~n16576;
  assign n14080 = ~n17596 & ~P2_IR_REG_27__SCAN_IN;
  assign n13774 = ~n13776 & ~n13775;
  assign n13775 = ~P2_IR_REG_28__SCAN_IN & ~P2_IR_REG_31__SCAN_IN;
  assign n13776 = ~n14084 & ~n13778;
  assign n13777 = n14081 | n13778;
  assign n15961 = ~P2_IR_REG_15__SCAN_IN;
  assign n14139 = ~n13160 & ~P2_IR_REG_16__SCAN_IN;
  assign n15959 = ~P2_IR_REG_3__SCAN_IN & ~P2_IR_REG_2__SCAN_IN;
  assign n14282 = ~P2_IR_REG_4__SCAN_IN & ~P2_IR_REG_5__SCAN_IN;
  assign n16037 = ~P2_DATAO_REG_7__SCAN_IN;
  assign n15123 = n15860 | n23872;
  assign n14150 = ~n18813;
  assign n14407 = ~n18795 | ~n13324;
  assign n14506 = ~n14769 | ~n14507;
  assign n14507 = ~n18032;
  assign n15851 = n15815 & P1_REG3_REG_26__SCAN_IN;
  assign n13492 = ~n14656 | ~n22775;
  assign n14505 = ~n14506;
  assign n23777 = ~n17368 | ~n22777;
  assign n13621 = n14033 & n13213;
  assign n13498 = ~n17359;
  assign n14030 = n17358 & n17357;
  assign n23926 = ~n13899 | ~n17356;
  assign n15750 = ~n15749 | ~SI_24_;
  assign n14098 = ~n15667;
  assign n15716 = n15715 & n15719;
  assign n14699 = n14700 & n15907;
  assign n13432 = ~n17896;
  assign n13429 = ~n17904;
  assign n19138 = n26367 ^ ~n17213;
  assign n14535 = n19135 & n19133;
  assign n19135 = n25731 & n25603;
  assign n13641 = n17213 ^ ~n25651;
  assign n14188 = ~n19719 | ~n14189;
  assign n13657 = ~n13658 | ~n19719;
  assign n13658 = ~n14190 | ~n14336;
  assign n13654 = n13657 | n14336;
  assign n13643 = n17235 & n17226;
  assign n13907 = ~n19295 & ~n14834;
  assign n13877 = ~n13962 | ~n13198;
  assign n14235 = ~n25870 & ~n14236;
  assign n13858 = ~n25921;
  assign n19822 = ~n13757 | ~n19821;
  assign n25974 = ~n14231 | ~n14232;
  assign n14232 = n14233 & n19913;
  assign n14233 = ~n13191 | ~n25931;
  assign n13860 = ~n25964 | ~n13863;
  assign n13861 = n13862 & n19992;
  assign n13863 = n25982 & P3_REG2_REG_11__SCAN_IN;
  assign n16063 = n16872 | P3_IR_REG_15__SCAN_IN;
  assign n13760 = n13761 & n20040;
  assign n13763 = ~n20006 | ~n13759;
  assign n20082 = ~n20077 | ~n20108;
  assign n13753 = ~P3_REG1_REG_17__SCAN_IN;
  assign n17091 = ~n16941 | ~n16909;
  assign n16899 = n16852 | P3_REG3_REG_20__SCAN_IN;
  assign n16798 = ~n16501 & ~n13840;
  assign n16529 = ~n16501 & ~P3_REG3_REG_16__SCAN_IN;
  assign n16501 = n16491 | P3_REG3_REG_15__SCAN_IN;
  assign n16491 = ~n13851 | ~n13850;
  assign n13850 = ~P3_REG3_REG_14__SCAN_IN;
  assign n16363 = ~P3_REG3_REG_13__SCAN_IN;
  assign n14198 = ~n18209 | ~n13121;
  assign n16373 = ~P3_REG3_REG_12__SCAN_IN;
  assign n16376 = ~n13177 & ~n13848;
  assign n16425 = ~n13852 | ~n16452;
  assign n13852 = n25667 & n13853;
  assign n26256 = ~n18159 | ~n26277;
  assign n26279 = ~n19274;
  assign n19503 = ~n18365 | ~n18364;
  assign n18365 = n20765 | n19228;
  assign n20144 = n14832 & n14831;
  assign n14831 = n20141 & n13138;
  assign n19295 = ~n19499;
  assign n20142 = n14832 & n13138;
  assign n14742 = n14743 & n18441;
  assign n13562 = ~n18305 | ~n14861;
  assign n14861 = ~n13152 & ~n13242;
  assign n20205 = ~n20208;
  assign n20233 = ~n19271 & ~n19270;
  assign n20293 = ~n13708 | ~n20259;
  assign n20331 = ~n14753 | ~n18428;
  assign n20352 = ~n20374 | ~n18255;
  assign n20385 = n18255 & n18254;
  assign n20387 = ~n13707 | ~n13706;
  assign n13706 = n18424 & n18423;
  assign n18425 = n13707 & n18423;
  assign n14838 = ~n14211 | ~n14216;
  assign n13574 = ~n20492 | ~n18418;
  assign n14740 = ~n14733 & ~n19388;
  assign n14733 = ~n18411 & ~n14741;
  assign n26054 = n14820 & n14818;
  assign n14818 = ~n14821;
  assign n26076 = n13943 & n18408;
  assign n26126 = ~n18385;
  assign n26233 = ~n18157 | ~n18402;
  assign n26273 = ~n19304 | ~n26316;
  assign n14549 = n14550 & P3_IR_REG_29__SCAN_IN;
  assign n14550 = ~P3_IR_REG_31__SCAN_IN | ~P3_IR_REG_28__SCAN_IN;
  assign n14330 = ~n16955 & ~n16954;
  assign n14483 = ~n16054;
  assign n14476 = n14477 & n16048;
  assign n14478 = ~n16047;
  assign n16039 = ~P2_DATAO_REG_8__SCAN_IN;
  assign n16034 = ~P2_DATAO_REG_6__SCAN_IN;
  assign n16027 = ~P2_DATAO_REG_4__SCAN_IN;
  assign n14793 = ~n16130;
  assign n14794 = ~n16026;
  assign n16021 = ~P2_DATAO_REG_2__SCAN_IN;
  assign n18939 = n25454 ^ ~n18920;
  assign n18937 = ~n13458 | ~n13457;
  assign n13458 = ~n18935;
  assign n14846 = ~n20805 & ~n14847;
  assign n14847 = ~n19029;
  assign n14132 = ~n20851;
  assign n14127 = ~n14129 & ~n14128;
  assign n14128 = ~n18994;
  assign n14129 = ~n20850;
  assign n14301 = ~n13163 | ~n14302;
  assign n13459 = ~n13787 | ~n13328;
  assign n14849 = ~n14851 & ~n14850;
  assign n14851 = ~n13388;
  assign n14850 = ~n20943;
  assign n24489 = ~n14121 | ~n18915;
  assign n24488 = n18919 & n14119;
  assign n18936 = n25090 ^ ~n19033;
  assign n17533 = ~P1_DATAO_REG_6__SCAN_IN;
  assign n14283 = ~n14118 | ~n14287;
  assign n14284 = n14285 & n19022;
  assign n14165 = ~n14613 | ~n14166;
  assign n14166 = ~n14267 & ~n13287;
  assign n14167 = ~n13156 | ~n13267;
  assign n13828 = n13149 | n21389;
  assign n21455 = ~n21452 & ~n21451;
  assign n21449 = ~n21448 & ~n21447;
  assign n24741 = ~n24729 & ~n24728;
  assign n15957 = ~P2_IR_REG_12__SCAN_IN;
  assign n17758 = n17746 & P2_REG3_REG_24__SCAN_IN;
  assign n21597 = ~n21619 | ~n21620;
  assign n17737 = n17722 & P2_REG3_REG_22__SCAN_IN;
  assign n17722 = n17711 & P2_REG3_REG_21__SCAN_IN;
  assign n17711 = n17695 & P2_REG3_REG_20__SCAN_IN;
  assign n17685 = n17671 & P2_REG3_REG_18__SCAN_IN;
  assign n16751 = ~n16661 & ~n16605;
  assign n17578 = ~P1_DATAO_REG_10__SCAN_IN;
  assign n25245 = ~n25240;
  assign n21609 = ~n17703 | ~n21412;
  assign n21631 = ~n14467 | ~n13153;
  assign n21661 = ~n14179 | ~n14177;
  assign n14177 = n14178 & n21678;
  assign n21694 = n21683 & n21682;
  assign n21757 = ~n14645 | ~n17816;
  assign n21790 = ~n17814 | ~n17813;
  assign n21843 = ~n13681 | ~n17808;
  assign n13681 = ~n21868 | ~n17807;
  assign n14634 = n14635 & n17802;
  assign n24948 = ~n14767 | ~n17585;
  assign n14449 = ~n17564;
  assign n25077 = ~n17532 | ~n17531;
  assign n14431 = ~n25155 & ~n25420;
  assign n25219 = ~n25218 | ~n25217;
  assign n25217 = ~n25174;
  assign n14817 = ~n25254 | ~n24454;
  assign n25241 = ~n14817 | ~n25240;
  assign n15830 = n15831 | n15827;
  assign n14138 = n14139 & n17017;
  assign n17613 = n17605 | P2_IR_REG_12__SCAN_IN;
  assign n15267 = ~n15270 & ~n15266;
  assign n17569 = n17556 | P2_IR_REG_8__SCAN_IN;
  assign n13975 = ~n22248;
  assign n15730 = ~n15697 & ~n15696;
  assign n14692 = ~n22290;
  assign n13979 = ~n13305 | ~n22279;
  assign n14680 = ~n15776;
  assign n14677 = ~n22265;
  assign n14673 = n13314 & n14674;
  assign n15646 = n22905 | n15860;
  assign n15654 = n15650 & n15649;
  assign n15650 = n22905 | n15823;
  assign n15353 = ~n15288 | ~P1_REG3_REG_10__SCAN_IN;
  assign n14697 = ~n13155 | ~n14698;
  assign n15815 = n15788 & P1_REG3_REG_25__SCAN_IN;
  assign n15766 = ~n15167;
  assign n15481 = ~n22174 | ~n14865;
  assign n15758 = n15730 & P1_REG3_REG_23__SCAN_IN;
  assign n15610 = ~n15585 & ~n15584;
  assign n14042 = n14770 & n14043;
  assign n15939 = n15851 & P1_REG3_REG_27__SCAN_IN;
  assign n14038 = ~n18015;
  assign n13912 = ~n22730 & ~n18702;
  assign n22705 = ~n13912 | ~n13617;
  assign n22729 = ~n13499 | ~n13797;
  assign n13499 = ~n13798 | ~n14650;
  assign n13798 = n14648 & n18043;
  assign n22753 = n23749 & n14518;
  assign n14518 = ~n14520 & ~n22341;
  assign n14650 = ~n17463 | ~n17464;
  assign n14350 = ~n17402;
  assign n22777 = ~n13914 | ~n23241;
  assign n15223 = ~n13535 | ~n13536;
  assign n13535 = n13537 & P1_REG3_REG_7__SCAN_IN;
  assign n13536 = ~n15157;
  assign n13804 = ~n17361;
  assign n14516 = n24155 & n24165;
  assign n15020 = n15554 | n16021;
  assign n13796 = ~n13506 | ~n13299;
  assign n13506 = ~n13288 | ~n13119;
  assign n14122 = ~n14123 | ~n18865;
  assign n13712 = ~n13503 | ~n13501;
  assign n22780 = ~n14345 | ~n14344;
  assign n14345 = ~n18649;
  assign n23751 = ~n23749 | ~n24242;
  assign n23823 = n14034 & n18876;
  assign n14782 = ~n13623;
  assign n23849 = ~n14784 | ~n17393;
  assign n23886 = n17391 & n17390;
  assign n23924 = ~n23949 | ~n17387;
  assign n15777 = ~n15751 | ~n15750;
  assign n15828 = n15805 & n15755;
  assign n15905 = n14925 & n14700;
  assign n15907 = ~P1_IR_REG_23__SCAN_IN;
  assign n15446 = n15445 & SI_14_;
  assign n14502 = ~n15371;
  assign n15012 = ~P1_IR_REG_0__SCAN_IN & ~P1_IR_REG_1__SCAN_IN;
  assign n14574 = n16094 & n14576;
  assign n13811 = ~n13894 | ~P3_ADDR_REG_2__SCAN_IN;
  assign n13416 = ~n13555 | ~n13557;
  assign n13557 = ~P1_ADDR_REG_6__SCAN_IN | ~n16545;
  assign n13555 = ~n14582 | ~n13558;
  assign n13558 = ~P3_ADDR_REG_6__SCAN_IN | ~n16547;
  assign n13415 = ~n14581 | ~n13556;
  assign n13556 = n13559 & n16315;
  assign n13559 = ~P1_ADDR_REG_6__SCAN_IN | ~n16545;
  assign n13425 = ~n16923 | ~P3_ADDR_REG_8__SCAN_IN;
  assign n17940 = n13421 & n17936;
  assign n13421 = ~n13420 | ~n13418;
  assign n13418 = n13419 & n17933;
  assign n19065 = n19063 | n19062;
  assign n19064 = ~n13424;
  assign n25603 = n19138 ^ ~n19134;
  assign n14539 = ~n13302 | ~n19194;
  assign n14540 = ~n19630 | ~n14541;
  assign n14541 = ~n19195 & ~n19190;
  assign n19547 = ~n19157 | ~n14196;
  assign n14196 = ~n19126 | ~n19735;
  assign n25616 = ~n19706 | ~n19149;
  assign n25651 = ~n26277;
  assign n19597 = n19173 | n19752;
  assign n19413 = ~n18242 | ~n18241;
  assign n20454 = ~n19646;
  assign n19666 = ~n19652 & ~n19121;
  assign n16452 = ~P3_REG3_REG_4__SCAN_IN & ~P3_REG3_REG_3__SCAN_IN;
  assign n16473 = n16471 & n16470;
  assign n19708 = ~P3_REG3_REG_9__SCAN_IN;
  assign n26125 = ~n26086;
  assign n19703 = ~n19145 | ~n19144;
  assign n19304 = ~n26287;
  assign n19721 = ~n13656 | ~n14336;
  assign n19735 = ~n19156 | ~n20517;
  assign n13646 = n13647 & n19152;
  assign n25730 = n25673 & n19133;
  assign n20165 = n18356 & n13839;
  assign n13839 = ~n18359 & ~n13385;
  assign n20310 = n16947 & n16946;
  assign n20334 = n16906 & n16905;
  assign n20398 = n16805 & n16804;
  assign n25773 = ~n19840;
  assign n25780 = n19967 ^ ~P3_REG1_REG_2__SCAN_IN;
  assign n13745 = ~n14000 | ~n14003;
  assign n14000 = ~n14002 & ~n14001;
  assign n14001 = ~P3_REG1_REG_1__SCAN_IN;
  assign n25783 = ~n13876 | ~n19966;
  assign n13876 = ~n13875 | ~n13873;
  assign n13873 = ~n19965 & ~n13874;
  assign n13739 = ~n19811 | ~n19810;
  assign n25839 = n19813 ^ ~n25850;
  assign n25928 = n19819 ^ ~n19984;
  assign n25950 = ~n14234 | ~n13191;
  assign n25949 = n14234 & n25930;
  assign n25971 = n19822 ^ ~n19989;
  assign n26012 = n25995 & n19927;
  assign n19947 = ~n20010 | ~n19942;
  assign n19269 = ~n14060 | ~n13404;
  assign n14061 = ~n19245 | ~n13121;
  assign n18355 = ~n13843;
  assign n20220 = ~n18310 | ~n18309;
  assign n18310 = n20793 | n18351;
  assign n18431 = ~n18273 | ~n18272;
  assign n18273 = n18270 | n19228;
  assign n20526 = n20481 & n20388;
  assign n26174 = ~n26351;
  assign n20540 = n20130 | n20129;
  assign n19501 = ~n19503;
  assign n18495 = n19222 ^ ~n19295;
  assign n20585 = ~n18288 | ~n18287;
  assign n18288 = n18285 | n18351;
  assign n13697 = n20270 & n13391;
  assign n20462 = ~n14728 | ~n19400;
  assign n26158 = ~n14732 | ~n19346;
  assign n26391 = n26278 | n19305;
  assign n17178 = n17177 | n16337;
  assign n18348 = ~n18337 | ~n18336;
  assign n14063 = n14064 & n18334;
  assign n16286 = n17172 ^ ~P3_IR_REG_26__SCAN_IN;
  assign n16014 = ~P3_IR_REG_23__SCAN_IN;
  assign n19308 = n17146 & n17147;
  assign n17300 = ~n14488 | ~n17272;
  assign n17302 = n17299 | P2_DATAO_REG_20__SCAN_IN;
  assign n17270 = ~n13437 | ~n17078;
  assign n13437 = ~n13157 | ~n13344;
  assign n16872 = n16790 | P3_IR_REG_14__SCAN_IN;
  assign n16254 = ~n16204;
  assign n16043 = ~n13438 | ~n14068;
  assign n14068 = n16041 & n14069;
  assign n13438 = ~n14489 | ~n14066;
  assign n16203 = P1_DATAO_REG_8__SCAN_IN ^ ~P2_DATAO_REG_8__SCAN_IN;
  assign n16138 = P1_DATAO_REG_7__SCAN_IN ^ ~P2_DATAO_REG_7__SCAN_IN;
  assign n14805 = ~n13710;
  assign n16204 = n16124 | P3_IR_REG_6__SCAN_IN;
  assign n18169 = ~SI_6_;
  assign n16146 = ~P3_IR_REG_4__SCAN_IN;
  assign n16154 = n16026 & n16025;
  assign n16082 = P1_DATAO_REG_1__SCAN_IN ^ ~P2_DATAO_REG_1__SCAN_IN;
  assign n16175 = n16076 & P2_DATAO_REG_0__SCAN_IN;
  assign n24341 = n18939 ^ ~n18940;
  assign n17621 = n24052 | n17704;
  assign n14383 = ~n17664 | ~n21352;
  assign n21684 = ~n25559;
  assign n17603 = n24065 | n17704;
  assign n17641 = n25302 | n17704;
  assign n14857 = ~n14860 & ~n14858;
  assign n14858 = ~n24422;
  assign n17651 = n25296 | n17704;
  assign n25079 = n21031 | n17049;
  assign n24491 = ~n24488 | ~n24489;
  assign n13886 = n25290 | n17704;
  assign n21478 = n18126 & n17779;
  assign n16615 = ~n21356 | ~P2_REG2_REG_2__SCAN_IN;
  assign n14324 = n22139 & P2_REG2_REG_1__SCAN_IN;
  assign n24796 = ~n24763 & ~n24762;
  assign n21521 = ~n21910;
  assign n21542 = ~n21619 | ~n13984;
  assign n16676 = n16674 & P2_REG3_REG_11__SCAN_IN;
  assign n16686 = n16714 | n16602;
  assign n16725 = ~n16742 & ~n16589;
  assign n17497 = n25361 | n17704;
  assign n17494 = n24333 | n13793;
  assign n25273 = ~n25092;
  assign n25233 = n25373 & n17863;
  assign n25277 = ~n21395 & ~n17029;
  assign n18150 = n18122 ^ ~n21447;
  assign n18121 = n18120 | n18119;
  assign n21477 = n21460 | n17855;
  assign n14390 = ~n14093 | ~n25246;
  assign n14093 = n14094 ^ ~n21445;
  assign n14094 = ~n13591 | ~n13322;
  assign n21541 = ~n14627 | ~n14630;
  assign n14627 = ~n14633 | ~n21556;
  assign n14633 = ~n17828;
  assign n21618 = ~n14621 | ~n17824;
  assign n14621 = ~n21640 | ~n17823;
  assign n21662 = ~n13171 | ~n14435;
  assign n18146 = ~n17865 | ~n17864;
  assign n17059 = n17011 & n17447;
  assign n14328 = n16577 & n17034;
  assign n16580 = ~P2_IR_REG_29__SCAN_IN;
  assign n17033 = ~n14084 | ~n14082;
  assign n22156 = n15967 ^ ~P2_IR_REG_26__SCAN_IN;
  assign n17008 = n15972 ^ ~P2_IR_REG_24__SCAN_IN;
  assign n17015 = ~n17021 | ~P2_IR_REG_31__SCAN_IN;
  assign n15661 = ~n15607 | ~n15606;
  assign n21407 = ~n17022 | ~n17021;
  assign n17022 = ~n17020 | ~n17019;
  assign n13584 = ~n13585 & ~n15369;
  assign n13585 = ~n13179 & ~n13588;
  assign n17521 = ~P1_DATAO_REG_5__SCAN_IN;
  assign n17503 = ~P1_DATAO_REG_3__SCAN_IN;
  assign n22874 = n15695 & n15694;
  assign n23235 = ~P1_REG3_REG_8__SCAN_IN;
  assign n13601 = n13602 & n15628;
  assign n13600 = ~n22219 | ~n13218;
  assign n13602 = ~n13218 | ~n13604;
  assign n15527 = n25296 | n15810;
  assign n15386 = ~P1_REG3_REG_13__SCAN_IN;
  assign n14684 = ~n14688 & ~n14685;
  assign n14685 = ~n22247;
  assign n15323 = n25320 | n15810;
  assign n14265 = ~n15023 | ~n14260;
  assign n14260 = ~n23967 | ~n15046;
  assign n15023 = n24000 | n15823;
  assign n22293 = n13980 & n13143;
  assign n13980 = ~n13982 | ~n13981;
  assign n13982 = ~n22278;
  assign n23332 = ~n23279;
  assign n17377 = ~n18856;
  assign n18856 = n18854 | n18861;
  assign n14156 = n18842 & n14161;
  assign n14159 = ~n18842 | ~n14157;
  assign n13542 = n13544 & n18901;
  assign n18863 = n15943 & n15942;
  assign n22516 = n15704 & n15703;
  assign n22551 = n15675 & n15674;
  assign n16511 = n16808 & P1_STATE_REG_SCAN_IN;
  assign n13731 = ~n23436 & ~n13732;
  assign n23437 = ~n13733 | ~n23433;
  assign n23483 = ~n23464 | ~n23463;
  assign n14245 = ~n23483;
  assign n23516 = ~n13721 | ~n13719;
  assign n23660 = ~n23658 & ~n14252;
  assign n14252 = ~n23657 & ~P1_REG1_REG_15__SCAN_IN;
  assign n23721 = n14251 ^ ~n14250;
  assign n14250 = ~P1_REG1_REG_19__SCAN_IN;
  assign n14251 = ~n23708 | ~n23709;
  assign n14522 = ~n14524;
  assign n22492 = ~n13599;
  assign n22845 = n13918 ^ ~n22509;
  assign n13918 = ~n14668 | ~n18056;
  assign n14668 = n22513 | n22514;
  assign n22569 = ~n22617 & ~n14514;
  assign n22565 = ~n14780 & ~n14779;
  assign n14786 = n14787 & n18019;
  assign n22625 = ~n18896;
  assign n13630 = n13631 & n18010;
  assign n14519 = ~n14520;
  assign n14651 = ~n17463;
  assign n22568 = n24021 | n23991;
  assign n17466 = ~n23749 | ~n13154;
  assign n15252 = ~n15223 & ~n23235;
  assign n15288 = n15252 & P1_REG3_REG_9__SCAN_IN;
  assign n23820 = ~n13606 | ~n13605;
  assign n13605 = ~n13608 & ~n23818;
  assign n13606 = ~n13607;
  assign n15189 = ~n15157 & ~n15156;
  assign n13618 = ~n23967 & ~n24122;
  assign n24027 = ~n24122;
  assign n22824 = ~n22460 & ~n22459;
  assign n24241 = ~n24230;
  assign n24123 = n18854 & n18861;
  assign n15933 = ~n14955 | ~n14909;
  assign n14955 = ~n14954 | ~n14953;
  assign n22150 = n13540 ^ ~n13381;
  assign n15781 = ~n15784;
  assign n22163 = n15777 ^ ~n15828;
  assign n15870 = n14934 ^ ~P1_IR_REG_24__SCAN_IN;
  assign n14934 = ~n15911 | ~P1_IR_REG_31__SCAN_IN;
  assign n14420 = n14421 & n14936;
  assign n14936 = ~P1_IR_REG_21__SCAN_IN;
  assign n15664 = ~n15634 | ~n15633;
  assign n13715 = ~n15629 | ~n15661;
  assign n15604 = ~n15578 | ~n15603;
  assign n14107 = n14108 & n15545;
  assign n14106 = ~n13582 | ~n13297;
  assign n13887 = ~n15602 | ~n18249;
  assign n15602 = ~n14492 | ~n14494;
  assign n15344 = n15318 | n15317;
  assign n13460 = ~n14104 | ~n15177;
  assign n13659 = n14391 ^ ~n15117;
  assign n14276 = n15083 & n15082;
  assign n16823 = n14984 ^ ~n14248;
  assign n14248 = ~P1_IR_REG_31__SCAN_IN | ~P1_IR_REG_0__SCAN_IN;
  assign n23350 = ~P1_ADDR_REG_0__SCAN_IN;
  assign n16239 = n14580 | n14579;
  assign n16540 = ~n13507 | ~n13807;
  assign n13807 = ~n16321 | ~P2_ADDR_REG_4__SCAN_IN;
  assign n13507 = ~n13508 | ~n13509;
  assign n16546 = ~n13533 | ~n13560;
  assign n13533 = n14582 & n16545;
  assign n13560 = ~n14581 | ~n16315;
  assign n16836 = ~n13522 | ~n13520;
  assign n13520 = n13521 & P3_ADDR_REG_6__SCAN_IN;
  assign n13522 = ~n13523 | ~n14582;
  assign n17316 = n14586 ^ ~n13400;
  assign n17915 = ~n13426 | ~n13401;
  assign n13530 = ~n14577 & ~n17946;
  assign n19581 = ~n19763 | ~n19766;
  assign n20601 = ~n18431;
  assign n25666 = ~n17238 | ~n17183;
  assign n20632 = ~n18247 | ~n18246;
  assign n18247 = n18243 | n18351;
  assign n20593 = ~n18266 | ~n18258;
  assign n26359 = ~n26150;
  assign n20560 = ~n20197;
  assign n19781 = n14340 ^ ~n13282;
  assign n14342 = ~n19629;
  assign n25725 = n17242 & n20528;
  assign n14018 = n14016 & n13356;
  assign n14714 = n14716 & n14715;
  assign n14720 = ~n14721 & ~n19835;
  assign n14721 = ~n19531;
  assign n26455 = n19236 | n19235;
  assign n26451 = n18384 | n18383;
  assign n26448 = n18372 | n18371;
  assign n26445 = ~n20165;
  assign n26439 = ~n18330 | ~n18329;
  assign n26436 = ~n18316 | ~n18315;
  assign n20267 = ~n20310;
  assign n19674 = ~n20398;
  assign n19406 = n16419 | n16418;
  assign n19552 = n16368 | n16367;
  assign n26059 = n16349 | n16348;
  assign n26116 = n16409 | n16408;
  assign n26189 = n16358 | n16357;
  assign n16483 = ~n16460 | ~P3_REG2_REG_2__SCAN_IN;
  assign n26454 = ~P3_U3897;
  assign n25765 = ~n14003 | ~n19807;
  assign n25763 = n13875 & n19966;
  assign n25873 = ~n14237 | ~n25845;
  assign n13865 = ~n25964 | ~P3_REG2_REG_11__SCAN_IN;
  assign n13740 = ~n19829 | ~n19828;
  assign n26043 = n14238 & n19932;
  assign n13764 = ~n20006 | ~P3_REG1_REG_15__SCAN_IN;
  assign n13950 = ~n13951 | ~n13954;
  assign n13954 = n13955 & n20111;
  assign n13870 = ~n13960 | ~n20101;
  assign n20535 = ~n19269;
  assign n19230 = n20758 | n18351;
  assign n18354 = n20772 | n18351;
  assign n13448 = n18267 | n19228;
  assign n20369 = ~n14795 | ~n18261;
  assign n14795 = n18256 | n18351;
  assign n26393 = ~n18200 | ~n18199;
  assign n26224 = ~n18491 | ~n18490;
  assign n26431 = ~n18487 | ~n18462;
  assign n26390 = ~n18474 | ~n18473;
  assign n14835 = n17179 & n16338;
  assign n20759 = ~n16343;
  assign n20779 = n18348 ^ ~n18347;
  assign n18335 = ~n14062 | ~n18320;
  assign n14062 = n18319 | n18318;
  assign n20801 = ~n18301 | ~n18300;
  assign n18301 = n18299 | n13121;
  assign n19306 = ~n19308;
  assign n17138 = ~P3_IR_REG_20__SCAN_IN;
  assign n17076 = ~n14052 | ~n14056;
  assign n14052 = ~n14059 | ~n16950;
  assign n16053 = ~n16789;
  assign n18219 = n16789 ^ ~n16788;
  assign n16519 = ~n14807 | ~n16052;
  assign n14479 = ~n16275 | ~n16046;
  assign n18203 = n16275 ^ ~n16276;
  assign n16118 = ~n16033 | ~n16032;
  assign n20806 = n14134 ^ ~n14133;
  assign n14133 = ~n20805;
  assign n14134 = ~n21000 | ~n19029;
  assign n21830 = ~n22041;
  assign n13455 = ~n13137 | ~n13790;
  assign n24455 = n17058 & n17051;
  assign n14428 = ~n14429 | ~P1_DATAO_REG_1__SCAN_IN;
  assign n18916 = ~n14120 | ~n18915;
  assign n20865 = ~n19003 | ~n20943;
  assign n20878 = ~n13461 | ~n19018;
  assign n24452 = ~n25254 | ~n14815;
  assign n14815 = ~n18125 & ~n14816;
  assign n24470 = ~n14814 | ~n24402;
  assign n24499 = ~n24455;
  assign n25580 = n17772 | n17771;
  assign n25574 = n17753 | n17752;
  assign n25571 = n17742 | n17741;
  assign n25568 = n17729 | n17728;
  assign n25565 = n17716 | n17715;
  assign n25562 = n17702 | n17701;
  assign n25556 = n17676 | n17675;
  assign n21436 = n16650 | n16649;
  assign n21735 = n16757 | n16756;
  assign n21818 = n16669 | n16668;
  assign n21413 = n16638 | n16637;
  assign n21817 = n16707 | n16706;
  assign n24955 = n16658 | n16657;
  assign n25000 = n16690 | n16689;
  assign n25022 = n16720 | n16719;
  assign n24934 = n24932 ^ ~n13898;
  assign n13898 = n25194 ^ ~n21691;
  assign n21461 = n17873 & n13989;
  assign n13989 = n13161 & n13990;
  assign n21470 = ~n17873 | ~n13161;
  assign n25105 = ~n25284 | ~n25189;
  assign n25551 = n18146 | n18109;
  assign n25515 = ~n25488;
  assign n25373 = n17059 & P2_STATE_REG_SCAN_IN;
  assign n14438 = ~n16583 | ~P2_IR_REG_31__SCAN_IN;
  assign n23130 = ~n17976 | ~n17975;
  assign n17974 = ~n17961;
  assign n15845 = ~n14306 | ~n15838;
  assign n22165 = ~n17006;
  assign n17324 = ~n17008;
  assign n25297 = ~P1_DATAO_REG_17__SCAN_IN;
  assign n25325 = n14351 ^ ~n15277;
  assign n15244 = ~n13664 | ~n13662;
  assign n13662 = n13660 & n15269;
  assign n22172 = ~n13611;
  assign n22186 = n14675 & n15685;
  assign n14683 = ~n14688;
  assign n23311 = ~P1_STATE_REG_SCAN_IN | ~n15929;
  assign n15558 = n25290 | n15810;
  assign n23277 = n15924 & n23936;
  assign n24320 = n15855 | n15854;
  assign n24311 = ~n22515;
  assign n24304 = ~n22516;
  assign n24301 = ~n22551;
  assign n22999 = n15508 | n15507;
  assign n23034 = ~n22790;
  assign n23874 = n15068 | n15067;
  assign n13615 = ~n13200 & ~n13613;
  assign n13482 = n14919 & n14920;
  assign n13718 = ~n13720 | ~n23515;
  assign n13717 = ~n23493 | ~n13212;
  assign n23583 = ~n13726 | ~n23554;
  assign n13726 = ~n23552 | ~n23553;
  assign n13724 = ~n23582 & ~n13725;
  assign n23629 = ~n13730 | ~n23624;
  assign n13730 = ~n23623 | ~n23622;
  assign n23657 = n23655 ^ ~n23656;
  assign n23707 = n23706 ^ ~n24036;
  assign n22413 = n17983 ^ ~n22414;
  assign n22446 = n14116 & n13493;
  assign n14261 = ~n14773 | ~n18034;
  assign n14405 = ~n22588;
  assign n22695 = ~n14271 | ~n18014;
  assign n23936 = n24033 | n17436;
  assign n24284 = n17443 | n17442;
  assign n13910 = n14113 & n13240;
  assign n24240 = n17443 | n17439;
  assign n14292 = n14297 & n14293;
  assign n14291 = n13387 & n17970;
  assign n23351 = n15933;
  assign n15442 = n14587 | n15445;
  assign n24053 = ~P2_DATAO_REG_14__SCAN_IN;
  assign n24066 = ~P2_DATAO_REG_12__SCAN_IN;
  assign n24072 = ~P2_DATAO_REG_11__SCAN_IN;
  assign n24078 = ~P2_DATAO_REG_10__SCAN_IN;
  assign n24084 = ~P2_DATAO_REG_9__SCAN_IN;
  assign n16115 = ~n13578 | ~n13580;
  assign n16243 = n16245 ^ ~n16244;
  assign n13909 = n16930 & n16931;
  assign n13808 = ~n16932;
  assign n13728 = ~n14272 | ~n14273;
  assign n14571 = n17881 & n17889;
  assign n17899 = ~n17902;
  assign n14584 = n23184 & n17931;
  assign n13532 = ~n13890;
  assign n19219 = n14186 & n13310;
  assign n14601 = ~n14603 | ~n14604;
  assign n14885 = n19106 | n15914;
  assign n13911 = n14105 & n18914;
  assign n14253 = n23730 & n23731;
  assign n16834 = ~n13553 | ~n13125;
  assign n14598 = n13124 & n14599;
  assign n15391 = ~n15186;
  assign n13135 = n15785 | n17704;
  assign n18829 = ~n18779;
  assign n18159 = ~n14809;
  assign n13136 = ~n13358 | ~n21619;
  assign n21058 = ~n21159;
  assign n13137 = n13788 & n13317;
  assign n21556 = ~n21558;
  assign n13138 = n20174 | n26442;
  assign n14597 = ~n14598;
  assign n13139 = ~n19394 & ~n19393;
  assign n16003 = ~P3_IR_REG_24__SCAN_IN;
  assign n13140 = n13789 & n18942;
  assign n13141 = ~n22349 & ~n15684;
  assign n19446 = ~n20376;
  assign n13906 = ~n26106;
  assign n19427 = ~n18253 | ~n18252;
  assign n13143 = n15515 | n15514;
  assign n17196 = n15037;
  assign n13144 = n13709 & n16038;
  assign n13145 = n15572 | n15571;
  assign n13146 = ~n18051 & ~n18053;
  assign n13147 = ~n15171 | ~n15172;
  assign n13148 = n15274 & n13261;
  assign n13149 = n21384 | n21383;
  assign n13150 = n14349 & n13374;
  assign n13151 = n18761 & n14154;
  assign n13152 = ~n18304 & ~n20229;
  assign n13154 = n24242 & n14521;
  assign n13155 = n23237 | n15204;
  assign n13156 = n21375 | n21374;
  assign n13157 = n16889 | n13436;
  assign n13159 = n18488 | n26270;
  assign n13160 = P2_IR_REG_17__SCAN_IN | P2_IR_REG_18__SCAN_IN;
  assign n24298 = n15644 | n15643;
  assign n13716 = ~n24298;
  assign n14752 = n20349 ^ ~n19602;
  assign n13161 = n13991 & n21459;
  assign n13162 = n19459 | n19834;
  assign n13163 = n13325 & n14811;
  assign n13164 = ~n18808 & ~n14148;
  assign n13779 = ~n25126;
  assign n13165 = n14353 & n14605;
  assign n13166 = n13335 & n14022;
  assign n13167 = n13301 & n19719;
  assign n13168 = n14798 & n18351;
  assign n15518 = n15489 | SI_16_;
  assign n23801 = n15258 | n15257;
  assign n13169 = ~n15723 | ~n15722;
  assign n13170 = n19514 & n14472;
  assign n13171 = n21772 & n14434;
  assign n13172 = n13702 & n16045;
  assign n13981 = ~n22279;
  assign n22589 = n15617 & n15616;
  assign n24295 = ~n22589;
  assign n17029 = ~n25194;
  assign n13173 = n14741 | n19391;
  assign n13174 = n13783 | n17731;
  assign n13175 = n13174 & n13345;
  assign n13176 = n14436 & n21771;
  assign n17897 = ~n17894 | ~n17893;
  assign n14662 = ~n18046 | ~n18013;
  assign n15530 = n14915 & n23132;
  assign n18050 = ~n15637 | ~n13294;
  assign n13177 = n16403 | P3_REG3_REG_10__SCAN_IN;
  assign n18125 = ~n24449;
  assign n13178 = n15467 | n15466;
  assign n13179 = n15338 & n15310;
  assign n13180 = n26205 | n26174;
  assign n14709 = ~n20406;
  assign n13181 = n16544 & n16317;
  assign n24052 = n14587 ^ ~n15443;
  assign n18176 = ~n18191 | ~n13121;
  assign n13182 = n17518 & n17517;
  assign n13183 = n21954 | n21586;
  assign n23254 = ~n15006 | ~n15005;
  assign n13184 = n13519 & n19066;
  assign n14289 = ~n20930;
  assign n18340 = n20759 & n20766;
  assign n19273 = n19321 & n19322;
  assign n17704 = ~n24333 | ~n13121;
  assign n26442 = ~n18346 | ~n18345;
  assign n13185 = n26106 & n19359;
  assign n21359 = n16781;
  assign n25697 = ~n13649 | ~n13646;
  assign n13186 = n14241 & n20010;
  assign n18860 = ~n18853;
  assign n19545 = n14538 & n19155;
  assign n13187 = n19460 | n19520;
  assign n13188 = ~n17632 | ~n14138;
  assign n13189 = n19369 & n19368;
  assign n13190 = n18431 ^ n20334;
  assign n20461 = n20656 ^ ~n20472;
  assign n14570 = ~n20461;
  assign n13191 = n25948 & n25930;
  assign n13192 = n14201 & n14199;
  assign n13193 = n20588 | n20589;
  assign n13194 = n16781 & P2_REG0_REG_5__SCAN_IN;
  assign n13195 = n14101 & n15267;
  assign n13197 = ~n17177 | ~n17179;
  assign n13198 = n13961 & n25822;
  assign n13199 = n17940 ^ n17938;
  assign n13200 = n13131 & P1_REG3_REG_1__SCAN_IN;
  assign n20163 = n20174 ^ ~n26442;
  assign n14834 = ~n20163;
  assign n13201 = ~n22295 | ~n22706;
  assign n13202 = n25104 & n13983;
  assign n14577 = n19061 ^ ~n19062;
  assign n17944 = ~n14577;
  assign n13203 = n21758 | n14644;
  assign n20539 = ~n19230 | ~n19229;
  assign n13596 = ~n22548;
  assign n18887 = n22750 & n17465;
  assign n13204 = n13145 & n22291;
  assign n13205 = n18744 & n18743;
  assign n13206 = n21369 & n21818;
  assign n13207 = n18411 | n13173;
  assign n18544 = ~n23993;
  assign n14463 = ~n17754;
  assign n13208 = n21302 | n21301;
  assign n13209 = n22387 | n14692;
  assign n13210 = n17174 | P3_IR_REG_26__SCAN_IN;
  assign n13211 = n20632 | n20416;
  assign n21582 = ~n14754 | ~n17717;
  assign n22264 = ~n15747 | ~n15746;
  assign n20405 = ~n14707 | ~n14711;
  assign n13212 = n23492 & n23515;
  assign n14462 = ~n17743;
  assign n14384 = ~n21411;
  assign n13213 = n17390 & n17392;
  assign n13214 = ~n15640 | ~P1_REG3_REG_20__SCAN_IN;
  assign n13215 = n22655 & n14040;
  assign n13216 = n25029 & n24997;
  assign n13217 = n14404 & n18050;
  assign n13218 = n22319 & n13603;
  assign n21544 = ~n21921;
  assign n13219 = n15445 | SI_14_;
  assign n13220 = n19563 | n19692;
  assign n13221 = n21986 | n25556;
  assign n13222 = n21332 | n21331;
  assign n13223 = n19371 | n19370;
  assign n22491 = n22495 ^ ~n22515;
  assign n13224 = n19841 & n19844;
  assign n14525 = ~n22819;
  assign n13225 = n19454 | n19453;
  assign n13226 = n18150 | n22038;
  assign n13227 = n20376 & n19834;
  assign n13228 = n21283 | n21282;
  assign n13229 = n19458 | n19457;
  assign n16583 = ~n14329 | ~n14327;
  assign n22535 = ~n22862;
  assign n26383 = ~n18195 | ~n18194;
  assign n13581 = ~n26383;
  assign n13230 = n14486 & n16870;
  assign n23769 = n15293 | n15292;
  assign n14344 = ~n23769;
  assign n13231 = n20593 ^ n17213;
  assign n13232 = n18434 & n19472;
  assign n13233 = n19246 & n19516;
  assign n13234 = n13153 & n14384;
  assign n13235 = n16052 & n13230;
  assign n13236 = n20233 & n20208;
  assign n13237 = n13233 & n19221;
  assign n13238 = n24327 ^ ~n22421;
  assign n20881 = ~n25577;
  assign n25577 = n17763 | n17762;
  assign n13239 = n18153 & n18152;
  assign n13240 = n19091 & n19090;
  assign n13786 = ~n17731;
  assign n14158 = ~n14161;
  assign n13241 = n15336 | n15335;
  assign n13242 = n20245 & n20266;
  assign n13243 = n18258 & n14198;
  assign n13244 = n13765 & n25903;
  assign n13245 = n22771 | n18042;
  assign n13246 = n13754 & n25942;
  assign n13247 = n14331 & n25643;
  assign n14266 = n24178;
  assign n25692 = ~n20517;
  assign n20517 = ~n16380 & ~n16379;
  assign n13248 = n14443 & n17562;
  assign n13249 = n15860 | n24027;
  assign n13250 = n19160 & n19153;
  assign n13251 = n18687 & n18665;
  assign n13252 = n19343 | n19342;
  assign n13253 = n19337 | n19336;
  assign n13254 = ~n18620 | ~n18619;
  assign n13255 = n13819 & n21227;
  assign n13256 = n14641 & n14640;
  assign n13257 = n18064 | n18063;
  assign n13258 = n21180 & n21191;
  assign n13259 = n16238 & n14578;
  assign n14515 = ~n22618;
  assign n13260 = n19177 & n13220;
  assign n13261 = n15309 | SI_10_;
  assign n13262 = ~n14152 | ~n18760;
  assign n13263 = ~n14938 & ~n15904;
  assign n13264 = n14582 & n16315;
  assign n13265 = n19064 | P1_ADDR_REG_17__SCAN_IN;
  assign n13266 = n23553 & n13723;
  assign n14615 = ~n21330;
  assign n13267 = n21388 | n21380;
  assign n13268 = n19278 & n19277;
  assign n19092 = ~n19095;
  assign n13269 = n19293 | n13903;
  assign n13270 = ~n18871 | ~n18866;
  assign n13271 = n21266 & n21265;
  assign n13272 = n15716 & n14098;
  assign n13273 = n19399 & n19398;
  assign n13274 = n25114 & n14315;
  assign n13275 = n19839 & n19840;
  assign n13276 = n15009 & n17207;
  assign n13277 = n17529 & n17539;
  assign n13278 = ~n16110 | ~n16238;
  assign n13279 = ~n18676 | ~n18675;
  assign n14711 = ~n14712;
  assign n14712 = ~n14713 | ~n18422;
  assign n20160 = ~n18354 | ~n18353;
  assign n14256 = ~n20160;
  assign n13280 = n13466 & n13464;
  assign n13281 = n21408 | n21393;
  assign n26316 = n17203 | n17202;
  assign n14005 = ~n26316;
  assign n13282 = n19194 & n19193;
  assign n13283 = n14215 | n14214;
  assign n20524 = ~n19391;
  assign n19391 = n18414 & n18413;
  assign n13284 = n17871 & n17870;
  assign n13285 = n21351 & n21350;
  assign n16144 = n17521 ^ ~P2_DATAO_REG_5__SCAN_IN;
  assign n13986 = ~n21932;
  assign n13683 = ~n17808;
  assign n13286 = ~n19838 | ~n19839;
  assign n13287 = n14612 & n14611;
  assign n13914 = ~n24231;
  assign n19085 = ~n17978 | ~n17977;
  assign n14526 = ~n19085;
  assign n13288 = n14400 & n14123;
  assign n13289 = n13183 & n21412;
  assign n13290 = n20163 | n14833;
  assign n13291 = n17367 & n17365;
  assign n13292 = n17764 & n17773;
  assign n13293 = n14500 & SI_14_;
  assign n13294 = n13716 & n15636;
  assign n13295 = n14419 & P1_IR_REG_31__SCAN_IN;
  assign n13296 = n19215 & n19199;
  assign n14257 = ~n21445;
  assign n18059 = n22819 | n24316;
  assign n17174 = ~P3_IR_REG_27__SCAN_IN;
  assign n13423 = ~n17927;
  assign n17927 = ~n17918 | ~n17917;
  assign n13297 = n14109 & n15543;
  assign n13298 = ~n14360 | ~n13271;
  assign n13299 = n14122 & n18059;
  assign n17179 = ~P3_IR_REG_28__SCAN_IN;
  assign n24059 = ~P2_DATAO_REG_13__SCAN_IN;
  assign n13300 = n13581 | n26116;
  assign n13301 = n19721 | n14189;
  assign n13302 = ~n13282 | ~n14542;
  assign n13303 = ~n13443 | ~n19493;
  assign n13304 = n22018 & n21735;
  assign n13719 = ~n13720;
  assign n13720 = ~n23497 | ~n23494;
  assign n22513 = ~n14401 | ~n18055;
  assign n14762 = ~n14763;
  assign n14763 = n17622 | n14764;
  assign n22488 = ~n18865;
  assign n13305 = n13204 & n13143;
  assign n26199 = ~n19340 | ~n19338;
  assign n13306 = n19424 & n18234;
  assign n13307 = ~n22664 & ~n24289;
  assign n21469 = ~n14170 | ~n14173;
  assign n13990 = ~n21469;
  assign n13308 = n13742 & n25859;
  assign n13309 = n17833 & n21445;
  assign n13310 = n19214 & n19213;
  assign n13311 = ~n24190 & ~n23875;
  assign n13312 = n14007 & n14006;
  assign n13313 = n16336 & n16335;
  assign n13314 = n22187 & n15685;
  assign n13315 = n17176 & n17175;
  assign n13316 = n13817 & n21154;
  assign n13317 = n24379 & n18950;
  assign n13318 = n14565 & n20208;
  assign n20330 = ~n14752;
  assign n13319 = ~P1_IR_REG_22__SCAN_IN & ~P1_IR_REG_21__SCAN_IN;
  assign n13320 = n20944 & n14131;
  assign n13321 = n22617 | n22618;
  assign n16345 = n16340 & n20752;
  assign n13322 = n13593 & n21409;
  assign n13323 = n13946 & n19978;
  assign n13324 = n18794 & n18800;
  assign n13325 = n14813 & n24402;
  assign n13326 = n14709 | n13902;
  assign n13327 = n13571 & n18218;
  assign n13328 = n18991 & n18990;
  assign n13329 = n18563 & n18548;
  assign n13330 = n23818 | n23234;
  assign n13331 = n14539 & n14185;
  assign n13332 = n18430 & n14748;
  assign n14956 = ~P1_IR_REG_27__SCAN_IN;
  assign n15603 = n15577 | SI_19_;
  assign n13333 = n13416 & n16837;
  assign n13334 = n20863 & n19006;
  assign n13335 = n14562 & n19470;
  assign n13336 = n18005 & n18004;
  assign n13337 = n17826 & n13674;
  assign n13338 = ~n18399 | ~n19325;
  assign n13339 = n13549 | n14756;
  assign n14839 = ~n14840;
  assign n14840 = ~n19287 & ~n14841;
  assign n13340 = n18009 & n13632;
  assign n13341 = n19028 & n14284;
  assign n13342 = n18838 & n18837;
  assign n13343 = n14417 & n18723;
  assign n17399 = ~n18649 | ~n23769;
  assign n13344 = n14053 & n13434;
  assign n13345 = n13292 & n14461;
  assign n13346 = n19482 & n19481;
  assign n13347 = P3_IR_REG_31__SCAN_IN & n17174;
  assign n13348 = n18701 & n18700;
  assign n13349 = n19486 & n19485;
  assign n13350 = n14040 & n14038;
  assign n13351 = n18115 & n17833;
  assign n13352 = ~n19159 | ~n19155;
  assign n14033 = n18876 & n17394;
  assign n13353 = n14504 & n22457;
  assign n13354 = ~n16736 & ~n13194;
  assign n13355 = n13806 & n17945;
  assign n13356 = n14470 & n19832;
  assign n13357 = n19688 & n19182;
  assign n13358 = n13984 & n21544;
  assign n13359 = n14876 & n19346;
  assign n13360 = n15240 & n14309;
  assign n13361 = ~n14681 & ~n14677;
  assign n13362 = ~n14281 | ~n18575;
  assign n13363 = ~n17996 | ~n17995;
  assign n14193 = ~n14194;
  assign n14194 = ~n19168 | ~n19765;
  assign n13364 = n24516 & P2_IR_REG_0__SCAN_IN;
  assign n13365 = n14482 & n16055;
  assign n14790 = ~P1_IR_REG_28__SCAN_IN & ~P1_IR_REG_27__SCAN_IN;
  assign n13366 = ~n19464 & ~n19463;
  assign n13367 = n14304 & P2_IR_REG_20__SCAN_IN;
  assign n13368 = n13700 & n14480;
  assign n13369 = n17809 & n13682;
  assign n13370 = n14150 & n18809;
  assign n13371 = n14301 & n24466;
  assign n13372 = n14159 & n18852;
  assign n13373 = ~n21975 | ~n21684;
  assign n13374 = ~n22257 | ~n23034;
  assign n13375 = n13210 | P3_IR_REG_25__SCAN_IN;
  assign n13376 = n13187 & n13162;
  assign n13377 = n14316 & n17808;
  assign n20257 = n13446 & n18434;
  assign n13934 = ~n20257;
  assign n13378 = n17945 & n17946;
  assign n13379 = n14476 & P2_DATAO_REG_13__SCAN_IN;
  assign n13380 = n14241 | n14240;
  assign n14701 = ~n14702;
  assign n14702 = ~n14924 | ~n14941;
  assign n14494 = ~n14495;
  assign n14495 = ~n14496 | ~n15546;
  assign n15904 = ~P1_IR_REG_31__SCAN_IN;
  assign n14090 = ~P2_IR_REG_1__SCAN_IN;
  assign n13885 = ~n21734;
  assign n13381 = n15837 ^ SI_27_;
  assign n13538 = ~P1_REG3_REG_6__SCAN_IN;
  assign n13598 = ~n22495;
  assign n13493 = ~n22752;
  assign n22008 = ~n17651 | ~n17650;
  assign n18779 = n18522 & n18508;
  assign n14434 = ~n21986;
  assign n25673 = ~n25672 | ~n25671;
  assign n22775 = ~n17366 | ~n13291;
  assign n15901 = n14932 ^ ~P1_IR_REG_25__SCAN_IN;
  assign n17631 = ~n17632 | ~n17634;
  assign n20492 = ~n14204 | ~n14202;
  assign n25028 = ~n17550 | ~n17549;
  assign n20452 = ~n13568 | ~n13327;
  assign n22745 = ~n13633 | ~n13630;
  assign n23794 = ~n13624 | ~n13622;
  assign n24967 = ~n14442 | ~n14446;
  assign n24365 = n24491 & n18919;
  assign n25118 = ~n17508 & ~n25136;
  assign n13382 = ~n18189 & ~n18188;
  assign n13383 = n23749 & n14519;
  assign n13384 = n20481 | P3_REG2_REG_29__SCAN_IN;
  assign n13385 = n16422 & P3_REG2_REG_28__SCAN_IN;
  assign n16076 = ~P1_DATAO_REG_0__SCAN_IN;
  assign n20376 = n16848 & n16847;
  assign n13386 = n21772 & n13176;
  assign n15443 = n15410 & n15409;
  assign n15445 = ~n15443;
  assign n13387 = ~n17979 & ~n14300;
  assign n13388 = ~n19005 | ~n19004;
  assign n13723 = ~n23584;
  assign n13389 = ~n14195 | ~n19168;
  assign n13390 = n13840 | P3_REG3_REG_18__SCAN_IN;
  assign n13511 = ~P2_ADDR_REG_6__SCAN_IN;
  assign n17037 = ~P1_DATAO_REG_1__SCAN_IN;
  assign n13391 = n20269 & n20268;
  assign n13392 = n14687 & n14690;
  assign n13393 = n19932 & n26042;
  assign n26053 = ~n18202 | ~n18201;
  assign n13394 = n20073 & n20075;
  assign n13874 = ~P3_REG2_REG_1__SCAN_IN;
  assign n13395 = n17455 & n17282;
  assign n13396 = n17366 & n17365;
  assign n13397 = n14867 & n17272;
  assign n13398 = n13724 | n23584;
  assign n15605 = ~n15573;
  assign n15573 = n15548 & n15547;
  assign n14688 = ~n14689 | ~n13241;
  assign n14809 = n14810;
  assign n25270 = ~n25246;
  assign n25246 = ~n21394 | ~n17788;
  assign n13399 = n21406 | n21405;
  assign n13400 = P3_ADDR_REG_10__SCAN_IN ^ P1_ADDR_REG_10__SCAN_IN;
  assign n14236 = ~n25845;
  assign n14137 = ~SI_24_;
  assign n13401 = n13431 & n17907;
  assign n14079 = ~n25183;
  assign n14521 = ~n23051;
  assign n13402 = n20111 & n20101;
  assign n23940 = ~n14517;
  assign n23949 = ~n23958 | ~n23950;
  assign n13403 = ~n13721 | ~n23494;
  assign n13404 = n18258 & n14061;
  assign n14604 = ~n14605 | ~n21456;
  assign n14173 = ~n14174;
  assign n14174 = ~n21364 & ~n17657;
  assign n26129 = n18373 & n19252;
  assign n13405 = P1_REG3_REG_20__SCAN_IN & P1_REG3_REG_21__SCAN_IN;
  assign n14605 = ~n21458;
  assign n13406 = n18915 & n17041;
  assign n13407 = n13607 | n13608;
  assign n19835 = n16015 ^ ~n16014;
  assign n13408 = n18861 & n18860;
  assign n13409 = n13509 & n16247;
  assign n13793 = ~n24586;
  assign n24565 = n16168 & n17487;
  assign n14424 = ~n24565;
  assign n14568 = n14569 & n20442;
  assign n14004 = ~n20094;
  assign n25503 = n25378 & n21407;
  assign n25378 = n21456 & n21030;
  assign n21916 = ~n21514 & ~n21513;
  assign n13992 = ~n25779 | ~n25780;
  assign n13995 = ~n13744 | ~n13308;
  assign n13413 = ~n25839;
  assign n14108 = ~n13297 | ~n14110;
  assign n21532 = ~n14464 | ~n17743;
  assign n17310 = ~n13728 | ~P2_ADDR_REG_9__SCAN_IN;
  assign n13711 = ~n17912 | ~n17911;
  assign n13567 = n16540 ^ ~n13181;
  assign n13554 = ~n13893 | ~n13425;
  assign n21432 = ~n21427 | ~n13411;
  assign n14376 = ~n14377 & ~n14602;
  assign n20007 = ~n13996 | ~n19830;
  assign n19819 = ~n13768 | ~n19818;
  assign n13744 = ~n13413 | ~n19814;
  assign P3_U3201 = ~n13414 | ~n20128;
  assign n13414 = ~n20127 & ~n20126;
  assign n13999 = ~n13747 | ~n20107;
  assign n25779 = ~n13745 | ~n19807;
  assign n13586 = ~n13583 | ~n13148;
  assign n14357 = n14610 & n14358;
  assign n17259 = n17312 ^ ~n17311;
  assign n16838 = ~n13415 | ~n13416;
  assign n16839 = ~n13333 | ~n13415;
  assign n17934 = ~n13417 | ~n17928;
  assign n13417 = ~n13423 | ~n13422;
  assign n13419 = ~n17926 | ~n17928;
  assign n13422 = ~n17926;
  assign n16926 = ~n13425 | ~n16924;
  assign n13893 = ~n13735 | ~n13425;
  assign n13426 = ~n13433 | ~n17904;
  assign n13428 = ~n13401 | ~n13429;
  assign n13430 = ~n17897 | ~n13401;
  assign n17905 = ~n17897 | ~n17896;
  assign n13431 = ~n13432 | ~n17904;
  assign n13433 = ~n17897;
  assign n16049 = ~n14475 | ~n14476;
  assign n16052 = ~n14475 | ~n13379;
  assign n14484 = ~n14808 | ~n13235;
  assign n16058 = ~n16889 | ~n16890;
  assign n13701 = ~n16043 | ~n13172;
  assign n13919 = ~n13442 | ~n14742;
  assign n13442 = ~n20185 | ~n14745;
  assign n13443 = ~n14742 | ~n13444;
  assign n13444 = ~n14745;
  assign n19013 = n13449 & n19012;
  assign n19009 = ~n19010 | ~n13449;
  assign n20960 = ~n20959 | ~n13449;
  assign n13454 = ~n13137 | ~n13450;
  assign n13450 = n13790 & n24353;
  assign n24354 = ~n13455 | ~n14825;
  assign n13453 = ~n24353;
  assign n13789 = ~n24341 | ~n13456;
  assign n13456 = ~n18937;
  assign n13457 = ~n18936;
  assign n20849 = ~n13459 | ~n18994;
  assign n15268 = ~n13460 | ~n15206;
  assign n25342 = n13460 ^ ~n15206;
  assign n13461 = ~n14118 | ~n20930;
  assign n13463 = ~n14905 | ~n14904;
  assign n14909 = ~n13462 | ~n14905;
  assign n14950 = n13463 | P1_IR_REG_27__SCAN_IN;
  assign n14527 = ~n13463 | ~P1_IR_REG_31__SCAN_IN;
  assign n13465 = ~n13279 | ~n18687;
  assign n13467 = ~n18707 | ~n13348;
  assign n13470 = ~n13280 | ~n13468;
  assign n13468 = n18707 & n18697;
  assign n18718 = ~n13470 | ~n13469;
  assign n18551 = ~n18550 | ~n13471;
  assign n13472 = ~n18546 | ~n24027;
  assign n18822 = ~n13475 | ~n13473;
  assign n13474 = ~n13164 | ~n13370;
  assign n13475 = ~n18810 | ~n13164;
  assign n18772 = ~n13478 | ~n13476;
  assign n13476 = n18766 & n13477;
  assign n13477 = ~n18761 | ~n13262;
  assign n13513 = ~n13479;
  assign n23191 = ~n13479 | ~n13199;
  assign n13479 = ~n14277 | ~n13510;
  assign n18599 = ~n13487 | ~n18587;
  assign n13487 = ~n13490 | ~n13488;
  assign n13488 = n13489 & n18572;
  assign n13489 = ~n14410 | ~n18573;
  assign n13490 = ~n13491 | ~n18567;
  assign n13491 = ~n18561 | ~n18560;
  assign n23878 = ~n13494 | ~n17359;
  assign n13494 = ~n23926 | ~n14031;
  assign n17362 = ~n13496 | ~n13495;
  assign n13497 = ~n14031 & ~n13498;
  assign n22652 = ~n13500 | ~n18892;
  assign n13500 = ~n14664 | ~n14663;
  assign n13501 = ~n22607 | ~n13502;
  assign n13504 = ~n13505 | ~n13800;
  assign n13802 = ~n22607 | ~n22625;
  assign n13505 = ~n13146 | ~n13801;
  assign n19078 = ~n13796;
  assign n13509 = ~n16243 | ~n16242;
  assign n23188 = ~n13510 | ~n23187;
  assign n13510 = ~n14583 | ~n17932;
  assign n13512 = ~n13199;
  assign n16320 = n13514 ^ ~n16313;
  assign n13514 = ~n13525 | ~n16241;
  assign n13561 = P3_ADDR_REG_1__SCAN_IN ^ ~P1_ADDR_REG_1__SCAN_IN;
  assign n13896 = ~n13515 | ~n14573;
  assign n13515 = ~n16095 | ~n14572;
  assign n13519 = ~n13527 | ~n13531;
  assign n23198 = ~n13518 & ~n13516;
  assign n13521 = ~n14582 | ~P1_ADDR_REG_5__SCAN_IN;
  assign n17257 = ~n13524 | ~P2_ADDR_REG_8__SCAN_IN;
  assign n16937 = ~n17256 | ~n13524;
  assign n13524 = ~n16929 | ~n13909;
  assign n13550 = ~n16548 | ~P2_ADDR_REG_6__SCAN_IN;
  assign n13529 = ~n23189 & ~n13530;
  assign n13806 = ~n13526 | ~n14577;
  assign n13526 = ~n23189 | ~n23191;
  assign n13528 = ~n23191 & ~n17944;
  assign n13531 = ~n13890 | ~n17946;
  assign n17945 = ~n13532 | ~n23189;
  assign n15222 = ~n13536 | ~n13537;
  assign n13540 = ~n15807 | ~n15827;
  assign n15600 = ~n15604;
  assign n18902 = ~n13543 | ~n13542;
  assign n15631 = n13547 & n13545;
  assign n13546 = ~n14495 | ~n15601;
  assign n13547 = ~n13582 | ~n13548;
  assign n16835 = ~n13552 | ~n16548;
  assign n16316 = ~n14581 | ~n14582;
  assign n13713 = ~n13554 | ~P3_ADDR_REG_9__SCAN_IN;
  assign n17254 = ~n13554;
  assign n16073 = ~n13561;
  assign n14228 = ~n13562 | ~n20205;
  assign n14227 = ~n13562 | ~n14223;
  assign n20206 = n13562 ^ ~n20205;
  assign n13564 = n13565 ^ ~n20163;
  assign n13565 = ~n18333 | ~n18332;
  assign n16539 = ~n13567;
  assign n16543 = ~n13567 | ~n13913;
  assign n13568 = ~n20492 | ~n13569;
  assign n20470 = ~n13574 | ~n18417;
  assign n15998 = n15997 & n15996;
  assign n16002 = n15998 | n16337;
  assign n14219 = ~n18226;
  assign n20372 = ~n13577 & ~n13576;
  assign n16114 = ~n13579 | ~n16101;
  assign n13579 = ~n16100 | ~n16099;
  assign n13578 = ~n13579;
  assign n13580 = ~n16101;
  assign n13878 = ~n13582 | ~n15517;
  assign n14492 = ~n13582 | ~n13879;
  assign n25302 = n13582 ^ ~n15516;
  assign n14117 = ~n13148 | ~n14503;
  assign n15370 = ~n13587 | ~n15339;
  assign n13587 = ~n14117 | ~n13179;
  assign n13588 = ~n15339;
  assign n21507 = ~n21532 | ~n17754;
  assign n13593 = ~n17764 | ~n14463;
  assign n13594 = ~n17764;
  assign n13603 = n22218 | n13604;
  assign n22320 = ~n22221 | ~n15599;
  assign n22221 = ~n22219 | ~n22218;
  assign n13607 = ~n23940 | ~n23845;
  assign n23848 = ~n14517 & ~n13608;
  assign n23873 = ~n23940 | ~n14516;
  assign n13608 = ~n14516 | ~n23872;
  assign n15308 = ~n13612 & ~n15300;
  assign n22200 = ~n13612 & ~n22199;
  assign n23307 = n13612 ^ ~n22199;
  assign n13612 = ~n14695 | ~n14697;
  assign n13613 = n15219 & P1_REG1_REG_1__SCAN_IN;
  assign n22703 = ~n13912;
  assign n22633 = ~n22678 | ~n22952;
  assign n13617 = ~n22702;
  assign n14517 = ~n24131 | ~n13618;
  assign n14788 = ~n13619 | ~n18018;
  assign n22649 = n13619 | n14789;
  assign n22648 = ~n13619 | ~n14789;
  assign n13622 = n13620 & n13330;
  assign n13620 = ~n14033 | ~n13623;
  assign n13624 = ~n17391 | ~n13621;
  assign n13628 = ~n18033;
  assign n17384 = ~n18549 | ~n13629;
  assign n13633 = ~n13634 | ~n18007;
  assign n13631 = ~n13636 | ~n13340;
  assign n13632 = ~n18008;
  assign n13634 = n13636 & n18009;
  assign n22770 = ~n13635 | ~n18008;
  assign n13635 = ~n18007 | ~n18006;
  assign n14530 = ~n20794 | ~n13638;
  assign n13638 = n16287 ^ ~P3_B_REG_SCAN_IN;
  assign n17205 = ~n18159 | ~n13641;
  assign n13639 = ~n14809 | ~n13640;
  assign n13640 = ~n13641;
  assign n17213 = ~n17192 | ~n17191;
  assign n16000 = ~n15998 | ~n16003;
  assign n14706 = ~n15998 | ~n13642;
  assign n14704 = ~n16000 & ~n13375;
  assign n13645 = ~n17227 | ~n17226;
  assign n19130 = ~n17227 | ~n13643;
  assign n17236 = ~n13645 | ~n13644;
  assign n13644 = ~n17235;
  assign n13650 = ~n19145;
  assign n19706 = ~n19145 | ~n13651;
  assign n13647 = ~n13648 | ~n14338;
  assign n13649 = ~n13650 | ~n14338;
  assign n19594 = ~n13655 | ~n13653;
  assign n13655 = n14192 | n13657;
  assign n13656 = n14192 | n14190;
  assign n14588 = ~n13659 | ~n14592;
  assign n14591 = n13659 & n15111;
  assign n17520 = n15138 ^ ~n13659;
  assign n13660 = ~n15239 | ~n13663;
  assign n13664 = ~n13661 | ~n14104;
  assign n13663 = ~n15206;
  assign n14439 = ~n18477 | ~n25553;
  assign n18477 = ~n13665 | ~n13226;
  assign n13670 = ~n13671 | ~n14618;
  assign n17828 = ~n13667 | ~n13671;
  assign n13667 = n14618 | n13674;
  assign n14626 = ~n13670 | ~n13668;
  assign n13669 = ~n13673 | ~n13337;
  assign n21584 = ~n13672 | ~n17825;
  assign n13672 = ~n14618 | ~n14622;
  assign n14645 = ~n17814 | ~n14643;
  assign n13680 = ~n14319 | ~n13377;
  assign n17811 = ~n13680 | ~n13369;
  assign n13685 = ~n18876;
  assign n23845 = ~n24190;
  assign n13696 = ~n23958;
  assign n16275 = ~n13699 | ~n13172;
  assign n13699 = ~n13704 | ~n16044;
  assign n14475 = ~n13701 | ~n13368;
  assign n13700 = ~n13172 | ~n16250;
  assign n16249 = ~n16043 | ~n16042;
  assign n13702 = ~n16044 | ~n13703;
  assign n16050 = ~n16049 | ~n24059;
  assign n16137 = ~n14804 | ~n13705;
  assign n20384 = ~n18425;
  assign n13708 = ~n20333 | ~n20258;
  assign n13710 = ~n14806 | ~n16032;
  assign n13709 = ~n13710 | ~n14802;
  assign n23181 = ~n13711 | ~n23180;
  assign n23183 = ~n23179 | ~n13711;
  assign n14401 = ~n13712 | ~n18054;
  assign n22871 = n13712 ^ ~n22544;
  assign n22904 = n13321 ^ ~n22905;
  assign n23541 = ~n13717 | ~n13718;
  assign n13722 = ~n23552 | ~n13266;
  assign n23596 = ~n13722 | ~n13398;
  assign n23708 = ~n23707 | ~P1_REG1_REG_18__SCAN_IN;
  assign n13727 = ~n23700 | ~n23701;
  assign n17260 = ~n13728 | ~n17309;
  assign n13732 = ~n23433;
  assign n23464 = ~n13731 | ~n13733;
  assign n14508 = ~n13734 | ~n24251;
  assign n19100 = ~n13734 | ~n24286;
  assign n13735 = n16924 & n16925;
  assign P1_U3262 = ~n13736 | ~n14253;
  assign n13736 = ~n23728 | ~n13737;
  assign n13737 = ~n23726 | ~n13738;
  assign n13738 = n23727 & n23725;
  assign n13993 = ~n13739 | ~n25820;
  assign n25821 = n13739 ^ ~n25820;
  assign n13996 = ~n13740 | ~n26026;
  assign n26028 = n13740 ^ ~n26026;
  assign n25860 = ~n13741 | ~n19814;
  assign n13741 = ~n25839 | ~P3_REG1_REG_5__SCAN_IN;
  assign n13742 = ~n19814 | ~n13743;
  assign n13743 = ~P3_REG1_REG_5__SCAN_IN;
  assign n19967 = n13746 ^ ~n16158;
  assign n13746 = ~n19806 & ~n16337;
  assign n13751 = ~n20065;
  assign n13747 = ~n13749 | ~n13748;
  assign n13748 = ~n13751 | ~n20067;
  assign n13749 = n13750 & n20104;
  assign n13750 = ~n20067 | ~n13753;
  assign n20105 = ~n13752 | ~n20067;
  assign n13752 = ~n20065 | ~P3_REG1_REG_17__SCAN_IN;
  assign n13757 = ~n13755 | ~n13246;
  assign n13754 = ~n19820 | ~n19901;
  assign n13755 = ~n13756 | ~n19820;
  assign n13756 = ~n25928;
  assign n25943 = ~n13758 | ~n19820;
  assign n13758 = ~n25928 | ~P3_REG1_REG_9__SCAN_IN;
  assign n13762 = ~n20008;
  assign n20039 = ~n13764 | ~n20008;
  assign n13761 = ~n13762 | ~n20038;
  assign n13768 = ~n13766 | ~n13244;
  assign n13765 = ~n19817 | ~n13770;
  assign n13766 = ~n13767 | ~n19817;
  assign n13767 = ~n25884;
  assign n25904 = ~n13769 | ~n19817;
  assign n13769 = ~n25884 | ~P3_REG1_REG_7__SCAN_IN;
  assign n17611 = ~n21841 | ~n21431;
  assign n13771 = ~n14081 | ~n13772;
  assign n14759 = ~n21676;
  assign n14075 = ~n25028 | ~n13248;
  assign n13780 = ~n21582 | ~n13781;
  assign n21555 = ~n13782 | ~n17731;
  assign n13782 = ~n21582 | ~n17730;
  assign n13783 = ~n14460 | ~n13784;
  assign n13784 = ~n17731 | ~n13785;
  assign n13785 = ~n17730;
  assign n20988 = ~n13787 | ~n18990;
  assign n20920 = ~n20919 | ~n13787;
  assign n13788 = ~n13140 | ~n13792;
  assign n13790 = ~n18938 | ~n13140;
  assign n24377 = ~n13791 | ~n13140;
  assign n13791 = n18938 | n13792;
  assign n24340 = ~n18938 | ~n18937;
  assign n13792 = ~n24341;
  assign n21000 = ~n14283 | ~n13341;
  assign n21001 = ~n14283 | ~n14284;
  assign n23941 = ~n13794 | ~n15045;
  assign n17948 = n13795 ^ ~n15041;
  assign n22749 = ~n14650 | ~n14648;
  assign n13797 = ~n13245 | ~n18043;
  assign n13799 = n14403 & n18052;
  assign n22588 = ~n13802 | ~n18049;
  assign n23852 = ~n17362 | ~n17361;
  assign n23829 = ~n17362 | ~n13803;
  assign n13803 = ~n13311 & ~n13804;
  assign n18144 = ~n18497 | ~n24286;
  assign n13805 = ~n18066 & ~n13257;
  assign n19060 = ~n13378 | ~n13806;
  assign n16929 = ~n16933 | ~n13808;
  assign n16933 = ~n13810 | ~n13809;
  assign n13908 = ~n13811 | ~n14575;
  assign n16109 = ~n13895 | ~n13811;
  assign n14613 = ~n13813 | ~n13812;
  assign n13812 = ~n13816 | ~n13208;
  assign n13814 = n14357 & n21308;
  assign n13815 = ~n13816 | ~n21303;
  assign n13816 = ~n21297 | ~n21296;
  assign n13818 = ~n21149 | ~n21148;
  assign n21234 = ~n13820 | ~n13255;
  assign n13819 = ~n13822 | ~n21229;
  assign n13820 = ~n21217 | ~n13821;
  assign n21228 = ~n21217 | ~n21218;
  assign n21408 = ~n13823 | ~n13828;
  assign n13823 = ~n14165 | ~n13829;
  assign n21454 = ~n13826 | ~n13824;
  assign n13826 = ~n13827 | ~n13828;
  assign n13827 = ~n14165;
  assign n13831 = ~n21270 | ~n13834;
  assign n14359 = ~n13831 | ~n13832;
  assign n13835 = n14360 & n21269;
  assign n17023 = ~n16878 | ~n13836;
  assign n13837 = ~n17023 | ~P2_IR_REG_31__SCAN_IN;
  assign n17025 = ~n13837 | ~P2_IR_REG_19__SCAN_IN;
  assign n16852 = ~n16851 | ~n19583;
  assign n16374 = ~n13177 & ~P3_REG3_REG_11__SCAN_IN;
  assign n13848 = ~n16373 | ~n13849;
  assign n13849 = ~P3_REG3_REG_11__SCAN_IN;
  assign n16386 = ~n16452 | ~n25667;
  assign n13853 = ~P3_REG3_REG_6__SCAN_IN;
  assign n25945 = ~n13854 | ~n19986;
  assign n13854 = ~n25921 | ~P3_REG2_REG_9__SCAN_IN;
  assign n13856 = ~n19986 | ~n26093;
  assign n13857 = ~n13858 | ~n19986;
  assign n25983 = ~n13865 | ~n19991;
  assign n13864 = ~n19991;
  assign n20062 = n13866 ^ ~P3_REG2_REG_17__SCAN_IN;
  assign n19971 = ~n13867 | ~n19970;
  assign n16089 = ~P3_IR_REG_31__SCAN_IN | ~n16086;
  assign n16339 = ~P3_IR_REG_31__SCAN_IN | ~n16338;
  assign n17180 = ~P3_IR_REG_31__SCAN_IN | ~n17179;
  assign n16958 = ~P3_IR_REG_31__SCAN_IN | ~n16960;
  assign n16160 = ~n16159 | ~P3_IR_REG_31__SCAN_IN;
  assign n16139 = ~n16204 | ~P3_IR_REG_31__SCAN_IN;
  assign n20128 = ~n13868 | ~n26031;
  assign n13868 = ~n13869 | ~n13872;
  assign n13869 = ~n13871 | ~n13870;
  assign n13871 = ~n13958 & ~n20111;
  assign n19977 = ~n25841 | ~P3_REG2_REG_5__SCAN_IN;
  assign n15544 = ~n13878 | ~n15518;
  assign n13880 = ~n14325 | ~n17833;
  assign n17834 = ~n14325 | ~n13309;
  assign n17872 = n13880 ^ ~n21445;
  assign n15408 = ~n13882 | ~n13881;
  assign n13882 = ~n13883;
  assign n15375 = ~n13883 | ~SI_13_;
  assign n13883 = ~n15374 | ~n15373;
  assign n14618 = ~n13884 | ~n14619;
  assign n21640 = ~n13884 | ~n17822;
  assign n21707 = ~n14642;
  assign n15574 = ~n13887 | ~n14163;
  assign n15579 = ~n13887 | ~n14389;
  assign n13890 = ~n23191 | ~n17944;
  assign n16923 = ~n13892 | ~n16921;
  assign n16924 = ~n13892 | ~n13891;
  assign n13891 = n16921 & n16922;
  assign n13892 = ~n16920 | ~n16919;
  assign n16930 = n16927 & n13893;
  assign n13894 = ~n16095 | ~n16094;
  assign n13895 = ~n13896 | ~n14575;
  assign n14575 = ~n14574 | ~n16095;
  assign n17894 = ~n17886 | ~n17885;
  assign n23178 = ~n23180 | ~n17909;
  assign n17925 = ~n23185 | ~n17922;
  assign n17903 = ~n23164 | ~n23166;
  assign n23167 = ~n14571 | ~n17882;
  assign n19077 = ~n23197 & ~n13184;
  assign n23204 = ~n13968 | ~n23337;
  assign n19106 = ~n19101 | ~n19102;
  assign n14016 = ~n14268 | ~n13170;
  assign n14268 = ~n14545 | ~n14543;
  assign n14051 = ~n14018 | ~n14017;
  assign n26255 = ~n19273 & ~n26279;
  assign n18393 = ~n20144 & ~n18376;
  assign n14013 = n14563 & n14014;
  assign n13920 = ~n18446 | ~n18447;
  assign n13897 = ~n24899 | ~n24900;
  assign n13899 = n17354 | n17353;
  assign n15724 = ~n15717 | ~n15716;
  assign n13900 = ~n16567 | ~n16566;
  assign n21483 = ~n17848 & ~n17847;
  assign n14319 = ~n24970 | ~n14321;
  assign n14047 = ~n14048 | ~n19303;
  assign n19279 = ~n13268 | ~n13905;
  assign n19297 = n19294 & n13907;
  assign n14332 = ~n14333 | ~n19141;
  assign n14192 = ~n19166 & ~n14194;
  assign n14254 = ~n16241 | ~n16313;
  assign n16245 = ~n16116 | ~n16115;
  assign n16564 = ~n14282 | ~n15959;
  assign n14092 = ~n13277 | ~n17530;
  assign n21866 = ~n24950 | ~n17594;
  assign P1_U3242 = ~n13911 | ~n14413;
  assign n25467 = ~n17561 | ~n17560;
  assign n14118 = ~n19014 | ~n20835;
  assign n17991 = ~n22413 | ~n24216;
  assign n19049 = ~n19041 & ~n19040;
  assign n14830 = ~n24438;
  assign n14826 = ~n14828;
  assign n15717 = ~n14099 | ~n15667;
  assign n14125 = ~n22472 | ~n22488;
  assign n13913 = ~P2_ADDR_REG_5__SCAN_IN;
  assign n14579 = ~n16238;
  assign n14104 = ~n13915 | ~n15175;
  assign n14103 = ~n14100 | ~n13915;
  assign n25348 = n13915 ^ ~n15175;
  assign n20546 = n13919 ^ ~n20155;
  assign n18464 = ~n13920 | ~n26433;
  assign n18476 = ~n13920 | ~n26398;
  assign n18419 = ~n13921 | ~n20493;
  assign n20672 = n13921 ^ ~n20500;
  assign n13924 = ~n18425 | ~n13925;
  assign n13923 = ~n13925 | ~n13928;
  assign n13925 = ~n13927 & ~n13926;
  assign n13928 = ~n18426;
  assign n20363 = ~n20387 | ~n18426;
  assign n20207 = ~n13929 | ~n19472;
  assign n13929 = ~n13934 | ~n13933;
  assign n20234 = ~n20257 & ~n18435;
  assign n13935 = ~n13941 | ~n14722;
  assign n13937 = ~n13938 | ~n13939;
  assign n13938 = ~n13940;
  assign n13941 = ~n13940 & ~n14712;
  assign n13942 = ~n20442;
  assign n18421 = ~n20443 | ~n20442;
  assign n20443 = ~n14722 | ~n14723;
  assign n26109 = ~n26111;
  assign n13943 = ~n13944 | ~n26111;
  assign n13944 = ~n26107;
  assign n13945 = ~n25907 | ~n25906;
  assign n25863 = ~n19977 | ~n19976;
  assign n13946 = ~n13947 | ~n25862;
  assign n13948 = ~n13949 | ~n25862;
  assign n13949 = ~n19977;
  assign n13952 = ~n13960 | ~n13402;
  assign n13958 = ~n13953 | ~n20103;
  assign n13953 = ~n13959 | ~n20101;
  assign n13957 = ~n20103;
  assign n20102 = ~n20097 | ~n20096;
  assign n13959 = ~n20096;
  assign n13961 = ~n19971 | ~n13965;
  assign n13962 = ~n13963 | ~n19971;
  assign n13963 = ~n25800;
  assign n25823 = ~n13964 | ~n19971;
  assign n13964 = ~n25800 | ~P3_REG2_REG_3__SCAN_IN;
  assign n13965 = ~P3_REG2_REG_3__SCAN_IN;
  assign n20033 = ~n20029 | ~P3_REG2_REG_15__SCAN_IN;
  assign n20029 = n20031 ^ ~n19999;
  assign n20031 = ~n13967 | ~n19998;
  assign n13967 = ~n13118 | ~n26036;
  assign n14895 = ~n14921;
  assign n14921 = ~n14892 | ~n14891;
  assign n23342 = ~n13968 & ~n23335;
  assign n13968 = ~n15170 | ~n13147;
  assign n13969 = ~n19106 | ~n15918;
  assign P1_U3220 = ~n14885 | ~n13970;
  assign n22306 = ~n13971 | ~n15713;
  assign n13971 = ~n13972 | ~n14673;
  assign n13972 = ~n22234 | ~n13141;
  assign n13976 = ~n14686 | ~n14684;
  assign n22334 = ~n13976 | ~n22248;
  assign n13974 = ~n22333 & ~n13975;
  assign n22219 = ~n13978 | ~n13977;
  assign n13977 = ~n22277 | ~n13305;
  assign n25361 = n15033 ^ ~n15069;
  assign n25088 = ~n13142 | ~n25104;
  assign n13983 = ~n25090;
  assign n17853 = ~n17873 | ~n21497;
  assign n19811 = ~n25802 | ~P3_REG1_REG_3__SCAN_IN;
  assign n19824 = ~n25971 | ~P3_REG1_REG_11__SCAN_IN;
  assign n19829 = ~n26005 | ~P3_REG1_REG_13__SCAN_IN;
  assign n13994 = ~n25986 | ~n25985;
  assign n20127 = n13997 & n26027;
  assign n13997 = n13999 ^ ~n13998;
  assign n13998 = ~n20113;
  assign n14006 = ~n19433 & ~n14709;
  assign n14007 = ~n14008 | ~n19426;
  assign n14008 = ~n19423 | ~n19422;
  assign n19344 = ~n14012 & ~n14009;
  assign n14009 = ~n14010 | ~n13252;
  assign n14010 = ~n14011 | ~n14555;
  assign n14011 = ~n14554 | ~n13253;
  assign n19492 = ~n14015 | ~n14013;
  assign n14014 = ~n14565 | ~n13346;
  assign n14015 = ~n19478 | ~n13318;
  assign n14019 = ~n14268 | ~n19514;
  assign n14017 = ~n14019 | ~n14474;
  assign n19471 = ~n14020 | ~n13166;
  assign n14020 = ~n14557 | ~n14021;
  assign n14022 = ~n14561 | ~n13376;
  assign n14566 = ~n14023 | ~n14567;
  assign n14023 = ~n14024 | ~n20477;
  assign n14024 = ~n19395 | ~n14025;
  assign n14028 = ~n19355 | ~n13185;
  assign n14029 = ~n14028 | ~n14026;
  assign n14547 = ~n14029 | ~n14548;
  assign n18007 = ~n14774 | ~n13150;
  assign n23897 = ~n14030 | ~n17359;
  assign n14031 = ~n14032;
  assign n24158 = n23926 ^ ~n14032;
  assign n23925 = n23924 ^ ~n14032;
  assign n14034 = ~n14784 | ~n14782;
  assign n14036 = ~n22655 | ~n13350;
  assign n14037 = ~n22725 | ~n13215;
  assign n22656 = ~n14039 | ~n18015;
  assign n14039 = ~n22725 | ~n14785;
  assign n14040 = ~n14041 | ~n18015;
  assign n22543 = ~n22545 | ~n22544;
  assign n18033 = n22543 & n14043;
  assign n14348 = ~n22543 | ~n14042;
  assign n19242 = ~n14044 | ~n19240;
  assign n20758 = n14044 ^ ~n19240;
  assign n18363 = ~n14045 | ~n18360;
  assign n20772 = n14045 ^ ~n18360;
  assign P3_U3296 = ~n14049 | ~n14046;
  assign n14046 = ~n14047 | ~n14720;
  assign n14048 = ~n14714 | ~n14717;
  assign n14049 = ~n14050 | ~n19531;
  assign n14050 = ~n14051 | ~n19528;
  assign n16951 = ~n16058 | ~n16057;
  assign n14057 = ~n14058 | ~n16950;
  assign n20749 = n19244 ^ ~n19243;
  assign n14060 = ~n20749 | ~n19245;
  assign n18337 = ~n14065 | ~n14063;
  assign n14064 = ~n18318 | ~n18320;
  assign n14065 = ~n18319 | ~n18320;
  assign n16202 = ~n14489 | ~n13144;
  assign n16223 = ~n14067 | ~n16040;
  assign n14067 = ~n16202 | ~n16203;
  assign n14069 = ~n14070 | ~n16040;
  assign n17456 = ~n14071 | ~n17282;
  assign n14071 = ~n17280 | ~n17279;
  assign n21755 = ~n14072 | ~n17629;
  assign n14767 = ~n14076 | ~n14443;
  assign n14076 = ~n17564 | ~n14446;
  assign n14082 = ~n16576 & ~n17596;
  assign n14754 = ~n14089 | ~n14465;
  assign n14086 = ~n14087 | ~n14385;
  assign n14437 = ~n17487;
  assign n17550 = ~n25051 | ~n17548;
  assign n25051 = ~n14440 | ~n14092;
  assign n14099 = ~n15630 | ~n14372;
  assign n14101 = ~n15206 | ~n14102;
  assign n14102 = ~n15177;
  assign n14110 = ~n15518;
  assign n14113 = ~n22447 | ~n24011;
  assign n22447 = n14115 ^ ~n19098;
  assign n14114 = ~n14116 | ~n24247;
  assign n14115 = ~n19097 | ~n19096;
  assign n15337 = ~n14117 | ~n15310;
  assign n20931 = n14118 ^ ~n14289;
  assign n14119 = ~n18918 | ~n18917;
  assign n20942 = ~n14130 | ~n20850;
  assign n14130 = ~n20849 | ~n20851;
  assign n14131 = ~n20850 | ~n14132;
  assign n14140 = ~n14143 | ~n14141;
  assign n14142 = ~n14422 | ~n18642;
  assign n14143 = ~n14145 | ~n14144;
  assign n14144 = n14423 & n18642;
  assign n14145 = ~n18611 | ~n18610;
  assign n14147 = ~n14925 | ~n14420;
  assign n14149 = ~n18809;
  assign n18731 = ~n18724 | ~n18723;
  assign n14151 = ~n18724 | ~n13343;
  assign n14416 = ~n14151 | ~n18729;
  assign n14152 = ~n14154 | ~n14153;
  assign n14155 = ~n18749 | ~n18754;
  assign n14160 = ~n18834 | ~n14156;
  assign n18859 = ~n14160 | ~n13372;
  assign n14161 = ~n18841 | ~n13342;
  assign n14389 = ~n14163 | ~n15573;
  assign n21371 = ~n14169 | ~n14171;
  assign n14169 = ~n22132 | ~n14173;
  assign n14170 = n22132 | n14168;
  assign n15444 = ~n14499 | ~n14500;
  assign n17624 = ~n15449 | ~n15486;
  assign n14178 = ~n14639 | ~n14640;
  assign n14179 = ~n14180 | ~n21744;
  assign n14182 = ~n14640;
  assign n17819 = ~n21744 | ~n17817;
  assign n14641 = ~n17819 | ~n14183;
  assign n14186 = ~n14184 | ~n13296;
  assign n19533 = ~n14540 | ~n14539;
  assign n19217 = ~n14184;
  assign n14191 = n19165 | n14194;
  assign n19763 = ~n14195 | ~n14193;
  assign n14195 = ~n19166 | ~n19165;
  assign n18208 = n16322 ^ ~n16323;
  assign n14197 = ~n18208 | ~n18209;
  assign n18211 = ~n14197 | ~n13243;
  assign n14201 = ~n26255 | ~n26258;
  assign n18399 = ~n26258;
  assign n14199 = ~n26258 | ~n14200;
  assign n14203 = ~n14209 | ~n14206;
  assign n14204 = ~n14205 | ~n14820;
  assign n14205 = n14209 & n18413;
  assign n20515 = ~n14208 | ~n18202;
  assign n14208 = ~n14819 | ~n14820;
  assign n14209 = n14819 | n14210;
  assign n14210 = ~n18202;
  assign n14211 = ~n14219 | ~n18233;
  assign n14217 = ~n14218 | ~n18233;
  assign n18235 = ~n20433 | ~n18233;
  assign n20433 = ~n18226 | ~n18225;
  assign n14222 = ~n26130 | ~n18181;
  assign n14221 = ~n19371;
  assign n26112 = n14222 ^ ~n26111;
  assign n14225 = n18331 & n14226;
  assign n18333 = ~n20182 | ~n18331;
  assign n20182 = ~n14228 | ~n18317;
  assign P3_U3204 = ~n14230 | ~n14229;
  assign n14229 = ~n13159 | ~n13384;
  assign n14230 = n18496 & n18494;
  assign n19844 = ~n13275 | ~n19838;
  assign n19845 = ~n13224 | ~n25771;
  assign n20076 = ~n20074 | ~n20073;
  assign n14231 = ~n25934 | ~n13191;
  assign n19883 = ~n14237 | ~n14235;
  assign n14247 = n23596 | n23597;
  assign n23726 = ~n14249 | ~n23722;
  assign n14249 = ~n23721;
  assign n25848 = ~n19867 | ~n19866;
  assign n25934 = ~n19900 | ~n19899;
  assign n20095 = ~n20061 | ~n20060;
  assign n19940 = ~n19941;
  assign n19941 = ~n26046 | ~n19939;
  assign n14855 = ~n26181 | ~n18162;
  assign n20281 = ~n20374 | ~n14842;
  assign n26130 = ~n26127 | ~n13906;
  assign n14259 = ~n23250;
  assign n14672 = ~n14981 | ~n14980;
  assign n18174 = ~n26161 | ~n26160;
  assign n26161 = ~n14852 | ~n14854;
  assign n15001 = ~n14259 | ~n14258;
  assign n14258 = ~n23252;
  assign n23252 = ~n14669 | ~n14670;
  assign n23124 = ~n14915;
  assign n19321 = ~n19312;
  assign n16467 = ~n16462 | ~n16461;
  assign n14696 = ~n14694 & ~n15237;
  assign n14666 = ~n14667 | ~n22514;
  assign n15056 = n15049 ^ ~n15647;
  assign n15070 = ~n14880 | ~n14987;
  assign n18022 = ~n22603 | ~n22604;
  assign n22725 = ~n14262 | ~n14662;
  assign n14262 = ~n22722;
  assign n14263 = ~n23924;
  assign n23898 = ~n14263 | ~n13362;
  assign n23069 = ~n14264 | ~n22842;
  assign n14264 = ~n22841 | ~n24011;
  assign n17391 = ~n23898 | ~n17389;
  assign n22722 = ~n14346 | ~n18012;
  assign n14281 = n23941;
  assign n23336 = ~n15137 | ~n15136;
  assign n15054 = n14265 ^ ~n15647;
  assign n23274 = n15133 ^ ~n15131;
  assign n17886 = ~n14586 | ~n17883;
  assign n14353 = ~n21408 | ~n14871;
  assign n14560 = n13312 | n19451;
  assign n14554 = ~n14556 | ~n13338;
  assign n22607 = ~n22632 & ~n14393;
  assign n14270 = ~n25997;
  assign n25997 = ~n19920 | ~n19919;
  assign n18039 = n19094 ^ ~n18060;
  assign n19094 = ~n14347 | ~n18038;
  assign n22545 = ~n22564 | ~n18025;
  assign n14272 = ~n17258;
  assign n14273 = ~n17259;
  assign n14501 = ~n15406 | ~n14502;
  assign n23250 = n14998 ^ ~n14997;
  assign P1_U3240 = ~n14274 | ~n13336;
  assign n14274 = ~n13120 | ~n23339;
  assign n14391 = ~n15115 | ~n15116;
  assign n15039 = ~n15085 | ~P1_DATAO_REG_3__SCAN_IN;
  assign n18810 = ~n14408 | ~n14407;
  assign n20472 = ~n19406;
  assign n14592 = ~n15114;
  assign n17352 = ~n14991 | ~n14990;
  assign n14806 = ~n16117;
  assign SUB_1596_U62 = ~n14275 | ~n23200;
  assign n14275 = ~n23199 | ~P2_ADDR_REG_18__SCAN_IN;
  assign n14993 = ~n17382 | ~n14983;
  assign n15652 = ~n22234;
  assign n15112 = ~n14276 | ~n15084;
  assign n15037 = ~n15085;
  assign n24970 = ~n14636 | ~n14634;
  assign n14277 = ~n23187 | ~n17930;
  assign n14278 = ~n15630 | ~n15631;
  assign n15302 = ~n14280;
  assign n15304 = ~n14280 | ~n22202;
  assign n14280 = n23308 | n22199;
  assign n23187 = ~n17925 | ~n14584;
  assign n16108 = ~n16109;
  assign n23180 = ~n23171 | ~n14585;
  assign n14408 = ~n14409 | ~n18800;
  assign n14285 = ~n14287 | ~n14286;
  assign n14288 = ~n14289 | ~n19018;
  assign n17980 = ~n17975 | ~n17962;
  assign n14290 = ~n17975 | ~n14291;
  assign n20818 = ~n14303 | ~n13371;
  assign n14303 = ~n18959 | ~n13163;
  assign n17020 = ~n14305 | ~n13367;
  assign n14304 = ~P2_IR_REG_19__SCAN_IN | ~P2_IR_REG_31__SCAN_IN;
  assign n14305 = ~n17023 | ~P2_IR_REG_31__SCAN_IN;
  assign n14307 = ~n14308 | ~n15829;
  assign n14308 = ~n15777;
  assign n19008 = ~n14848 | ~n20863;
  assign n15271 = ~n15241 | ~n13360;
  assign n15242 = ~n15241 | ~n15240;
  assign n14309 = ~SI_9_;
  assign n14312 = ~n17795 | ~n14310;
  assign n14311 = ~n13274 | ~n25040;
  assign n17799 = ~n14312 | ~n17797;
  assign n14314 = ~n16733;
  assign n14315 = ~n13354 | ~n14313;
  assign n14317 = ~n14321 | ~n14318;
  assign n24944 = ~n14320 | ~n17804;
  assign n14320 = ~n24970 | ~n17803;
  assign n14322 = ~n14323 | ~n17804;
  assign n16778 = ~n14324 | ~n16588;
  assign n16771 = ~n21356 | ~P2_REG2_REG_0__SCAN_IN;
  assign n14325 = ~n21518 | ~n17832;
  assign n14326 = ~n14325 | ~n13351;
  assign n18122 = ~n14326 | ~n18121;
  assign n16578 = ~n14329 | ~n14328;
  assign n19174 = ~n19594 | ~n19597;
  assign n16956 = ~n14330;
  assign n17084 = ~n14330 | ~n16960;
  assign n19145 = ~n14332 | ~n13247;
  assign n14333 = ~n25673;
  assign n14337 = ~n19579 & ~n19446;
  assign n14340 = ~n14341 | ~n19189;
  assign n14341 = ~n14343 | ~n14342;
  assign n14343 = ~n19630;
  assign n14346 = ~n22745 | ~n22728;
  assign n14347 = ~n14348 | ~n13353;
  assign n14349 = ~n14350 | ~n14776;
  assign n14351 = ~n14503 | ~n15274;
  assign P2_U3328 = ~n14354 | ~n14352;
  assign n14352 = ~n13281 | ~n13165;
  assign n14354 = ~n14355 | ~n14601;
  assign n14355 = ~n14356 | ~n14376;
  assign n14356 = ~n21454 | ~n21453;
  assign n21072 = ~n21071 & ~n21070;
  assign n21297 = ~n14359 | ~n14361;
  assign n14362 = ~n13228 | ~n21286;
  assign n17013 = ~n14365 | ~n14363;
  assign n14364 = n14366 | n17032;
  assign n17021 = ~n16878 | ~n14366;
  assign n21109 = ~n14367 | ~n21097;
  assign n14367 = ~n14369 | ~n14368;
  assign n14369 = ~n21074 | ~n21075;
  assign n21203 = ~n14370 | ~n13258;
  assign n14370 = ~n21168 | ~n14371;
  assign n14371 = ~n21140 | ~n21139;
  assign n23149 = ~n15785 | ~n15786;
  assign n14377 = n21455 & n17029;
  assign n21492 = n14390 & n13284;
  assign n15139 = ~n14391 | ~SI_5_;
  assign n22630 = ~n14395 | ~n18047;
  assign n14396 = ~n14667 | ~n14397;
  assign n14397 = ~n18055;
  assign n14399 = ~n18055 | ~n14402;
  assign n14403 = ~n14658 & ~n18051;
  assign n14404 = ~n14405 | ~n14658;
  assign n14409 = ~n18787 | ~n18786;
  assign n18583 = ~n18573 | ~n18574;
  assign n14413 = ~n18862 | ~n14414;
  assign n18744 = ~n14415 | ~n18738;
  assign n14415 = ~n14416 | ~n18732;
  assign n14421 = ~n14702 | ~P1_IR_REG_31__SCAN_IN;
  assign n14972 = ~n14418 | ~n14420;
  assign n14418 = n14925 | n15904;
  assign n14423 = ~n18631 | ~n13254;
  assign n14422 = ~n18631;
  assign n14429 = ~n17502;
  assign n14426 = ~n14427 | ~n24333;
  assign n14427 = ~n17038 & ~n13128;
  assign n25206 = ~n21061 | ~n14816;
  assign n21720 = ~n14435 | ~n21772;
  assign n14435 = n21722 & n13176;
  assign n21774 = ~n21772 | ~n21771;
  assign n14436 = ~n22008;
  assign n16575 = ~n16574 | ~n14437;
  assign P2_U3528 = ~n14439 | ~n18478;
  assign n17532 = ~n17530 | ~n17529;
  assign n14442 = ~n14449 | ~n17576;
  assign n24994 = ~n17564 | ~n17563;
  assign n14447 = ~n14448 | ~n17576;
  assign n21787 = ~n14452 | ~n17623;
  assign n14452 = ~n17611 | ~n14762;
  assign n14458 = ~n14459 | ~n14456;
  assign n17703 = ~n14467 | ~n13234;
  assign n14467 = ~n14759 | ~n13158;
  assign n14472 = ~n19521;
  assign n14473 = ~n19519;
  assign n14474 = n19519 & n19521;
  assign n14477 = ~n14480 | ~n14478;
  assign n16322 = ~n14479 | ~n16047;
  assign n14481 = ~n16276 | ~n16047;
  assign n16889 = ~n14484 | ~n13365;
  assign n14482 = ~n13230 | ~n14483;
  assign n16871 = ~n14485 | ~n16054;
  assign n14485 = ~n16053 | ~n14878;
  assign n14486 = ~n14487 | ~n16054;
  assign n17280 = ~n14488 | ~n13397;
  assign n14804 = ~n16033 | ~n14805;
  assign n16033 = ~n16145 | ~n16030;
  assign n16029 = ~n16157 | ~n14792;
  assign n16131 = ~n16157 | ~n16026;
  assign n16157 = ~n16155 | ~n16154;
  assign n15407 = ~n15372 | ~n15371;
  assign n14504 = ~n14506 | ~n14770;
  assign n22510 = ~n18033 & ~n18032;
  assign P1_U3525 = ~n14508 | ~n19220;
  assign n14509 = ~n22617;
  assign n22548 = ~n14510 | ~n14509;
  assign n23942 = ~n23940 | ~n24155;
  assign n23963 = ~n24131 | ~n24027;
  assign n22830 = ~n22494 | ~n22832;
  assign n18069 = n22494 & n14522;
  assign n16818 = n14527 ^ ~n14956;
  assign n14528 = n16286 & n14529;
  assign n17134 = ~n14530 | ~n16286;
  assign n14529 = ~P3_D_REG_0__SCAN_IN;
  assign n14531 = ~n14532 | ~n13260;
  assign n14532 = ~n19750 | ~n20310;
  assign n19185 = n14531 & n13357;
  assign n19565 = ~n14532 | ~n19177;
  assign n25642 = ~n14533 | ~n19141;
  assign n14533 = ~n25673 | ~n14535;
  assign n14537 = ~n25697 | ~n13250;
  assign n19166 = ~n14537 | ~n14536;
  assign n14536 = ~n13352 | ~n19160;
  assign n14542 = ~n19189 | ~n19629;
  assign n14543 = ~n14544 | ~n19834;
  assign n14544 = ~n19510 | ~n19511;
  assign n14545 = ~n14546 | ~n19520;
  assign n14546 = ~n19513 | ~n19512;
  assign n19384 = ~n14547 | ~n19376;
  assign n14552 = ~n14551 | ~n14549;
  assign n14551 = n17177 | n16337;
  assign n16340 = ~n14552 | ~n16339;
  assign n14555 = ~n26199;
  assign n14553 = ~n26199 & ~n19333;
  assign n14557 = ~n14558 | ~n13229;
  assign n14558 = ~n14559 | ~n14752;
  assign n14559 = ~n14560 | ~n13225;
  assign n14562 = ~n13366 | ~n19465;
  assign n14564 = ~n13349 | ~n20163;
  assign n19423 = ~n14566 | ~n14568;
  assign n14569 = ~n19410 | ~n14570;
  assign n17891 = ~n17882 | ~n17881;
  assign n14576 = ~P3_ADDR_REG_2__SCAN_IN;
  assign n16240 = ~n16238 | ~n14580;
  assign n16241 = ~n13259 | ~n14580;
  assign n14578 = ~P3_ADDR_REG_4__SCAN_IN;
  assign n16544 = ~n13264 | ~n14581;
  assign n14583 = ~n17925 | ~n23184;
  assign n17912 = ~n23171 | ~n23173;
  assign n14585 = n23173 & n17910;
  assign n23174 = ~n17900 | ~n17899;
  assign n23185 = ~n17921 | ~n17920;
  assign n25661 = ~n25660 | ~n25659;
  assign n14589 = n14588 & n15139;
  assign n14590 = ~n14591 | ~n15112;
  assign n14593 = ~n15112 | ~n15111;
  assign n15138 = ~n14593 | ~n15114;
  assign n14600 = ~n21389;
  assign n14606 = ~n21243;
  assign n21250 = ~n14609 | ~n21243;
  assign n14608 = ~n14607 | ~n14609;
  assign n21252 = ~n14608 | ~n21248;
  assign n14610 = ~n21338 & ~n21330;
  assign n14612 = ~n21338;
  assign n17795 = ~n14616 | ~n13274;
  assign n14616 = ~n14617;
  assign n25042 = ~n14617 | ~n25041;
  assign n25139 = ~n25113 | ~n14617;
  assign n21518 = ~n14626 | ~n14628;
  assign n21559 = ~n17828 | ~n17827;
  assign n14635 = ~n14637 | ~n24997;
  assign n14636 = ~n13216 | ~n25025;
  assign n14638 = ~n25025 | ~n25029;
  assign n24996 = ~n14638 | ~n17801;
  assign n21708 = ~n17819 | ~n17818;
  assign n18040 = ~n14647 | ~n17464;
  assign n14647 = ~n14651 | ~n17480;
  assign n14648 = n14649 & n18887;
  assign n14649 = ~n18885 | ~n17464;
  assign n14652 = ~n13276 | ~n15010;
  assign n15077 = ~n15010 | ~n15009;
  assign n15072 = ~n15071 | ~n14652;
  assign n14655 = ~n25330;
  assign n14656 = ~n17369 & ~n14657;
  assign n22776 = ~n14657;
  assign n14658 = ~n22604;
  assign n14664 = ~n18045 | ~n14660;
  assign n14661 = ~n14659 | ~n18046;
  assign n22699 = ~n18045 | ~n18044;
  assign n22723 = ~n14662;
  assign n22676 = ~n22698 | ~n18046;
  assign n22698 = ~n22699 | ~n22723;
  assign n16968 = ~n14672;
  assign n14669 = ~n14672 | ~n16969;
  assign n14670 = ~n14671 | ~n15647;
  assign n14671 = ~n16969;
  assign n16969 = ~n14971 | ~n13249;
  assign n14674 = ~n13141 | ~n22233;
  assign n14675 = ~n22348 | ~n13141;
  assign n22348 = ~n15652 | ~n15651;
  assign n19101 = ~n14676 | ~n14678;
  assign n14676 = ~n22264 | ~n13361;
  assign n14682 = ~n22264 | ~n22265;
  assign n17994 = ~n14682 | ~n15776;
  assign n14681 = ~n17995;
  assign n22250 = n14686 & n14683;
  assign n14686 = ~n15308 | ~n14690;
  assign n14687 = n15308 | n15307;
  assign n14693 = ~n22293 | ~n22291;
  assign n22386 = ~n14693 | ~n22290;
  assign n14698 = ~n15237;
  assign n14694 = ~n23203;
  assign n23207 = ~n23204 | ~n23203;
  assign n14695 = ~n23204 | ~n14696;
  assign n23238 = ~n23207 | ~n15205;
  assign n14939 = ~n14925 | ~n14924;
  assign n17172 = ~n14706 | ~P3_IR_REG_31__SCAN_IN;
  assign n14707 = n18421 | n19287;
  assign n14708 = ~n14710 & ~n14709;
  assign n20423 = ~n18421 | ~n18420;
  assign n14716 = ~n19222 | ~n13233;
  assign n14728 = ~n20478 | ~n19401;
  assign n18406 = ~n14732 | ~n13359;
  assign n14739 = ~n18412 | ~n14740;
  assign n20525 = ~n14735 | ~n14740;
  assign n14735 = n18412 | n14741;
  assign n18416 = ~n14739 | ~n14736;
  assign n14737 = ~n14741 | ~n14738;
  assign n14738 = ~n19388;
  assign n26052 = ~n18412 | ~n18411;
  assign n14741 = ~n26053;
  assign n14743 = ~n14745 | ~n14747;
  assign n20164 = ~n14744 | ~n18439;
  assign n14744 = ~n20185 | ~n18438;
  assign n14747 = ~n18439;
  assign n14748 = ~n14750 | ~n14749;
  assign n14753 = ~n18427 | ~n14884;
  assign n14761 = ~n21676 | ~n17677;
  assign n21652 = ~n14761 | ~n17678;
  assign n21815 = ~n17611 | ~n21430;
  assign n17044 = ~n17049 | ~n13364;
  assign n14905 = ~n15452 & ~n14896;
  assign n14773 = ~n22510 | ~n22509;
  assign n14769 = n18035 & n22509;
  assign n14771 = ~n18035 | ~n14772;
  assign n14778 = ~n22782 | ~n17402;
  assign n14774 = ~n14775 | ~n14776;
  assign n14775 = ~n22782;
  assign n17481 = ~n14778 | ~n18882;
  assign n14776 = ~n17480 & ~n14777;
  assign n14780 = ~n18022;
  assign n22564 = ~n18022 | ~n14781;
  assign n14787 = ~n18018 | ~n14789;
  assign n22603 = ~n14788 | ~n14786;
  assign n14789 = ~n22629;
  assign n14907 = ~n14909;
  assign n14797 = ~n18256 | ~n14798;
  assign n19510 = ~n19508 | ~n14800;
  assign n19513 = ~n19508 | ~n14801;
  assign n14801 = n19511 & n19507;
  assign n16520 = ~n16052 | ~n16050;
  assign n18161 = ~n13192 | ~n14872;
  assign n26234 = ~n13192 | ~n26232;
  assign n16469 = ~n14809 | ~P3_U3897;
  assign n26306 = ~n18385 | ~n14809;
  assign n25683 = ~n25728 | ~n14809;
  assign n25710 = ~n25706 | ~n14809;
  assign n26253 = ~n26288 | ~n14809;
  assign n14811 = ~n14812 | ~n24401;
  assign n14814 = ~n24400 | ~n24401;
  assign n24400 = ~n18959 | ~n20973;
  assign n25279 = ~n21416 | ~n14817;
  assign n25243 = ~n25240 & ~n14817;
  assign n24440 = ~n14824 | ~n14828;
  assign n14824 = ~n24377 | ~n24379;
  assign n24439 = ~n14827 | ~n24379;
  assign n14827 = n24377 | n24378;
  assign n14829 = n24378 & n24379;
  assign n20396 = ~n14838 | ~n14839;
  assign n20414 = ~n18235 | ~n18234;
  assign n14845 = ~n21001 | ~n14846;
  assign n19042 = ~n14845 | ~n14843;
  assign n14844 = ~n14846 | ~n21002;
  assign n20959 = ~n14848 | ~n13334;
  assign n14856 = ~n26200 | ~n26199;
  assign n14852 = ~n26200 | ~n14853;
  assign n26184 = ~n14856 | ~n18162;
  assign n18927 = ~n18924 | ~n14857;
  assign n24424 = ~n14859 & ~n14860;
  assign n14859 = ~n18924;
  assign n18938 = ~n14863 | ~n14862;
  assign n24504 = ~n14863 | ~n18933;
  assign n14862 = n18934 & n18933;
  assign n14949 = ~n15865 | ~n14935;
  assign n14981 = n15167 | n18544;
  assign n15454 = n14922 & n15011;
  assign n20245 = ~n18436;
  assign n23983 = ~n23993 | ~n24122;
  assign n15866 = n15901 | n15870;
  assign n25174 = ~n25135 | ~n17499;
  assign n16588 = ~n22133;
  assign n14864 = n16570 & n16569;
  assign n24021 = n22436 & n23936;
  assign n14865 = n15435 | n15434;
  assign n24012 = n23914 & n23905;
  assign n14866 = n15219 & P1_REG1_REG_2__SCAN_IN;
  assign n14867 = n17680 | P2_DATAO_REG_20__SCAN_IN;
  assign n14869 = ~n15605 & ~n15604;
  assign n14870 = ~n15000 | ~n14999;
  assign n14871 = n21399 | n21398;
  assign n18424 = ~n20385;
  assign n14872 = n26233 & n26232;
  assign n14873 = n23293 & n15130;
  assign n14874 = n23874 & n24165;
  assign n16051 = ~P1_DATAO_REG_13__SCAN_IN;
  assign n26315 = n18443 & n19306;
  assign n23016 = ~n22176;
  assign n14875 = ~n16565 & ~P2_IR_REG_20__SCAN_IN;
  assign n17017 = ~P2_IR_REG_19__SCAN_IN;
  assign n14876 = ~n26189 | ~n26359;
  assign n14878 = n24053 | P1_DATAO_REG_14__SCAN_IN;
  assign n14879 = n26316 & n26315;
  assign n14880 = ~n15085 | ~P1_DATAO_REG_1__SCAN_IN;
  assign n14881 = ~n20601 | ~n20334;
  assign n14882 = ~n19171 | ~n19602;
  assign n14883 = ~n20306 | ~n18274;
  assign n14884 = n20369 | n20376;
  assign n21074 = ~n21073 & ~n21072;
  assign n19441 = ~n19440 & ~n20624;
  assign n19431 = ~n19429 | ~n19428;
  assign n19449 = ~n19448 & ~n19447;
  assign n19465 = ~n20263;
  assign n15048 = n18575 | n15823;
  assign n15129 = n15128 & n23274;
  assign n18410 = ~n19372;
  assign n17040 = n18920 ^ ~n25389;
  assign n15953 = ~P2_IR_REG_7__SCAN_IN & ~P2_IR_REG_10__SCAN_IN;
  assign n15049 = ~n15048 | ~n15047;
  assign n23737 = ~n17398 | ~n17397;
  assign n26227 = ~n18400 | ~n19327;
  assign n17787 = n21487 | n25583;
  assign n17634 = ~P2_IR_REG_16__SCAN_IN;
  assign n15352 = ~P1_REG3_REG_11__SCAN_IN;
  assign n14952 = ~P1_IR_REG_28__SCAN_IN;
  assign n15659 = n15658 & n15662;
  assign n15999 = ~P3_IR_REG_25__SCAN_IN;
  assign n26198 = ~n18403 | ~n18402;
  assign n26288 = ~n26137;
  assign n16326 = ~P3_IR_REG_12__SCAN_IN;
  assign n15986 = ~P3_IR_REG_3__SCAN_IN & ~P3_IR_REG_2__SCAN_IN;
  assign n17746 = n17737 & P2_REG3_REG_23__SCAN_IN;
  assign n17695 = n17685 & P2_REG3_REG_19__SCAN_IN;
  assign n17768 = n17758 & P2_REG3_REG_25__SCAN_IN;
  assign n16603 = ~P2_REG3_REG_10__SCAN_IN;
  assign n25253 = ~n25079;
  assign n23222 = n15056 ^ ~n15057;
  assign n15788 = n15758 & P1_REG3_REG_24__SCAN_IN;
  assign n15102 = ~n23874 | ~n13134;
  assign n18062 = ~n24316;
  assign n22761 = ~n22707;
  assign n15156 = ~P1_REG3_REG_5__SCAN_IN;
  assign n23958 = ~n17386 | ~n17385;
  assign n14926 = ~P1_IR_REG_24__SCAN_IN;
  assign n15667 = n15666 & n15665;
  assign n15517 = ~n15516;
  assign n20354 = ~n19602;
  assign n20235 = ~n26436;
  assign n16470 = ~P3_REG3_REG_8__SCAN_IN;
  assign n26280 = ~n26129;
  assign n26137 = ~n18387 | ~n19834;
  assign n16960 = ~P3_IR_REG_18__SCAN_IN;
  assign n19051 = ~n25580;
  assign n19029 = n19023 | n19024;
  assign n17671 = n16751 & n16606;
  assign n15960 = ~n17596 & ~n16568;
  assign n21352 = ~n17704;
  assign n21412 = n21965 | n20948;
  assign n25248 = n17836 & n17029;
  assign n16589 = ~P2_REG3_REG_5__SCAN_IN;
  assign n25509 = n17070 | n21402;
  assign n22253 = ~P1_REG3_REG_12__SCAN_IN;
  assign n15810 = n15450;
  assign n23796 = ~n17395;
  assign n23988 = ~n22789;
  assign n17962 = n17958 | SI_29_;
  assign n20416 = ~n19771;
  assign n25706 = ~n25724;
  assign n20186 = ~n26442;
  assign n26013 = P3_U3897 & n20773;
  assign n20501 = n18445 & n18452;
  assign n20627 = n20387 & n20386;
  assign n26140 = n26136 | n26135;
  assign n18307 = ~n18306 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n16181 = n16023 & n16022;
  assign n24500 = ~n24484;
  assign n24475 = ~n24511;
  assign n16779 = n16777 | n16776;
  assign n17864 = ~n18105 & ~n17863;
  assign n15967 = ~n15970 | ~P2_IR_REG_31__SCAN_IN;
  assign n17345 = n15687 & n15686;
  assign n23322 = n23217 & n23391;
  assign n24230 = n24123 & n15912;
  assign n18060 = ~n18864;
  assign n15871 = n24034 | P1_D_REG_0__SCAN_IN;
  assign n24011 = ~n23991;
  assign n24228 = n18854 & n15923;
  assign n15867 = n15870 | P1_B_REG_SCAN_IN;
  assign n14932 = ~n14931 | ~P1_IR_REG_31__SCAN_IN;
  assign n23656 = n15461 & n15460;
  assign n15338 = n15339 & n15314;
  assign n15212 = ~P1_IR_REG_7__SCAN_IN;
  assign n16008 = n16007 & n20802;
  assign n20552 = ~n20174;
  assign n25611 = ~n26059;
  assign n16403 = ~n16473 | ~n19708;
  assign n25667 = ~P3_REG3_REG_5__SCAN_IN;
  assign n18487 = n18451 & n18450;
  assign n18473 = n17461 & n19831;
  assign n19224 = ~n18363 | ~n18362;
  assign n24511 = n17066 & n17065;
  assign n21025 = n17072 & n25267;
  assign n16617 = ~n16612 | ~n16611;
  assign n24916 = n24896 | P2_U3088;
  assign n21828 = n25099 & n18124;
  assign n25099 = ~n25284 | ~n25277;
  assign n18145 = ~n25370 & ~n17009;
  assign n17006 = n15971 & n15970;
  assign n23329 = ~n23322;
  assign n18907 = n15930 & P1_STATE_REG_SCAN_IN;
  assign n22847 = n15794 & n15793;
  assign n23724 = n23356 | n23391;
  assign n23684 = ~n23729;
  assign n23892 = n24021 | n23970;
  assign n23944 = n24021 | n24001;
  assign n17442 = ~n15871 | ~n24113;
  assign n17443 = n17438 | n17437;
  assign n16313 = ~P1_ADDR_REG_4__SCAN_IN;
  assign n25734 = ~n17169 | ~n17168;
  assign n19752 = ~n20334;
  assign n26027 = ~n25741;
  assign n26031 = n20002 & n20001;
  assign n26270 = n18489 & n20528;
  assign n26433 = ~n26431;
  assign n26398 = ~n26390;
  assign n17285 = ~n20792;
  assign n24336 = n17011 | n21339;
  assign n24508 = ~n21025;
  assign n24506 = ~n24471;
  assign n25583 = ~n17786 | ~n17785;
  assign n25559 = n17690 | n17689;
  assign n24875 = ~n24896;
  assign n25263 = n21803;
  assign n25282 = n18110 & n25267;
  assign n25553 = ~n25551;
  assign n25289 = ~n16976 | ~n22156;
  assign n24707 = n17557 & n17569;
  assign n22164 = n13121 & P2_U3088;
  assign n23343 = ~n23311;
  assign n23309 = ~n23339;
  assign n23688 = ~n23724;
  assign n23722 = ~n23501;
  assign n22772 = ~n22568;
  assign n24026 = ~n23944;
  assign n24019 = ~n24021;
  assign n24286 = ~n24284;
  assign n24251 = ~n24240;
  assign n24113 = n15865 | n15870;
  assign n24106 = ~n23156;
  assign n17461 = n19835 & P3_STATE_REG_SCAN_IN;
  assign n25592 = n24336 | P2_U3088;
  assign n25368 = ~n25373 | ~n25289;
  assign P3_U3897 = n16016 & n17461;
  assign P2_U3947 = ~n25592;
  assign n14896 = ~n14895 | ~n14922;
  assign n14898 = ~P1_IR_REG_26__SCAN_IN & ~P1_IR_REG_25__SCAN_IN;
  assign n14897 = ~P1_IR_REG_23__SCAN_IN & ~P1_IR_REG_22__SCAN_IN;
  assign n14902 = ~n14898 | ~n14897;
  assign n14900 = ~P1_IR_REG_20__SCAN_IN & ~P1_IR_REG_21__SCAN_IN;
  assign n14899 = ~P1_IR_REG_24__SCAN_IN & ~P1_IR_REG_19__SCAN_IN;
  assign n14901 = ~n14900 | ~n14899;
  assign n14903 = ~n14902 & ~n14901;
  assign n14904 = n15011 & n14903;
  assign n14906 = ~P1_IR_REG_29__SCAN_IN;
  assign n14913 = ~n14907 | ~n14906;
  assign n14908 = ~n14913 | ~P1_IR_REG_31__SCAN_IN;
  assign n14915 = n14908 ^ ~P1_IR_REG_30__SCAN_IN;
  assign n14910 = ~n14909 | ~P1_IR_REG_31__SCAN_IN;
  assign n14912 = ~n14910 | ~P1_IR_REG_29__SCAN_IN;
  assign n14911 = ~n14906 | ~P1_IR_REG_31__SCAN_IN;
  assign n14914 = ~n14912 | ~n14911;
  assign n23117 = n14913;
  assign n14918 = ~n23132;
  assign n14917 = ~n13131 | ~P1_REG3_REG_0__SCAN_IN;
  assign n14916 = ~n23124 | ~n23132;
  assign n14920 = ~n15530 | ~P1_REG2_REG_0__SCAN_IN;
  assign n14919 = ~n15219 | ~P1_REG1_REG_0__SCAN_IN;
  assign n14974 = ~n14923 | ~n15454;
  assign n14925 = ~n14974;
  assign n14931 = ~n14933 | ~n14926;
  assign n14928 = ~n14931;
  assign n14927 = ~P1_IR_REG_25__SCAN_IN;
  assign n14929 = ~n14928 | ~n14927;
  assign n15911 = ~n14933;
  assign n14937 = ~n13263 | ~P1_IR_REG_21__SCAN_IN;
  assign n14945 = ~n14938;
  assign n14940 = ~n14939 | ~P1_IR_REG_31__SCAN_IN;
  assign n14943 = ~n14940 | ~P1_IR_REG_20__SCAN_IN;
  assign n14941 = ~P1_IR_REG_20__SCAN_IN;
  assign n14942 = ~n14941 | ~P1_IR_REG_31__SCAN_IN;
  assign n14944 = ~n14943 | ~n14942;
  assign n18853 = ~n14944 | ~n14945;
  assign n15024 = ~n14949 | ~n18545;
  assign n14948 = ~n23993 | ~n14983;
  assign n14946 = ~P1_REG1_REG_0__SCAN_IN;
  assign n14947 = n14949 | n14946;
  assign n14971 = n14948 & n14947;
  assign n14951 = ~n14950 | ~P1_IR_REG_31__SCAN_IN;
  assign n14954 = ~n14951 | ~P1_IR_REG_28__SCAN_IN;
  assign n14953 = ~n14952 | ~P1_IR_REG_31__SCAN_IN;
  assign n16809 = ~n15933 | ~n16818;
  assign n14977 = ~P1_IR_REG_0__SCAN_IN;
  assign n14970 = n16809 | n14977;
  assign n14965 = ~n14960 | ~n14959;
  assign n14961 = ~P3_ADDR_REG_19__SCAN_IN;
  assign n14964 = ~n14963 | ~n14962;
  assign n14966 = ~n21363 | ~SI_0_;
  assign n16176 = ~P2_DATAO_REG_0__SCAN_IN;
  assign n14968 = ~n14966 | ~n16176;
  assign n14967 = P2_DATAO_REG_0__SCAN_IN & SI_0_;
  assign n14989 = ~n15037 | ~n14967;
  assign n16103 = n14968 & n14989;
  assign n14969 = ~n16809 | ~n16103;
  assign n24122 = ~n14970 | ~n14969;
  assign n14973 = ~P1_IR_REG_22__SCAN_IN;
  assign n14975 = ~n14974 | ~P1_IR_REG_31__SCAN_IN;
  assign n15912 = ~n23905 | ~n18853;
  assign n15925 = ~n15912;
  assign n24001 = ~n24123 | ~n15925;
  assign n14976 = ~n24001;
  assign n14979 = n15024 | n24027;
  assign n14978 = n14949 | n14977;
  assign n14980 = n14979 & n14978;
  assign n14982 = ~n15530 | ~P1_REG2_REG_1__SCAN_IN;
  assign n14986 = ~n15379 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n14984 = ~P1_IR_REG_1__SCAN_IN;
  assign n14985 = n16809 | n16823;
  assign n14987 = ~n17036 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n15007 = n15070 ^ ~SI_1_;
  assign n14988 = SI_0_ & P1_DATAO_REG_0__SCAN_IN;
  assign n16078 = ~n15085 | ~n14988;
  assign n15073 = n16078 & n14989;
  assign n17038 = n15007 ^ ~n15073;
  assign n14990 = n15450 | n17038;
  assign n14992 = ~n17352 | ~n13132;
  assign n14994 = ~n14993 | ~n14992;
  assign n14996 = n15167 | n24015;
  assign n14995 = n15823 | n24131;
  assign n14998 = ~n14996 | ~n14995;
  assign n15000 = ~n14997;
  assign n14999 = ~n14998;
  assign n23316 = ~n15001 | ~n14870;
  assign n15003 = ~n15530 | ~P1_REG2_REG_2__SCAN_IN;
  assign n15002 = ~n15421 | ~P1_REG3_REG_2__SCAN_IN;
  assign n15004 = ~n15003 | ~n15002;
  assign n15006 = ~n15004 & ~n14866;
  assign n15005 = ~n18512 | ~P1_REG0_REG_2__SCAN_IN;
  assign n15074 = ~n15070 | ~SI_1_;
  assign n15010 = ~n15085 | ~P1_DATAO_REG_2__SCAN_IN;
  assign n15009 = ~n15037 | ~P2_DATAO_REG_2__SCAN_IN;
  assign n15022 = n25361 | n15450;
  assign n15018 = ~n15011;
  assign n15013 = n15012 | n15904;
  assign n15016 = ~n15013 | ~P1_IR_REG_2__SCAN_IN;
  assign n15015 = ~n15014 | ~P1_IR_REG_31__SCAN_IN;
  assign n15017 = ~n15016 | ~n15015;
  assign n24107 = ~n15018 | ~n15017;
  assign n15019 = n16809 | n24107;
  assign n24144 = ~n23967;
  assign n15026 = n15167 | n24000;
  assign n15823 = n15024;
  assign n15025 = n15823 | n24144;
  assign n15052 = ~n15026 | ~n15025;
  assign n23317 = n15054 ^ ~n15052;
  assign n23221 = ~n23316 | ~n23317;
  assign n15028 = ~n15219 | ~P1_REG1_REG_3__SCAN_IN;
  assign n15027 = ~n13129 | ~P1_REG0_REG_3__SCAN_IN;
  assign n15032 = ~n15028 | ~n15027;
  assign n15030 = ~n15530 | ~P1_REG2_REG_3__SCAN_IN;
  assign n15062 = ~P1_REG3_REG_3__SCAN_IN;
  assign n15029 = ~n15421 | ~n15062;
  assign n15031 = ~n15030 | ~n15029;
  assign n18575 = ~n17357;
  assign n15035 = ~n15034 | ~SI_2_;
  assign n15038 = ~n15037 | ~P2_DATAO_REG_3__SCAN_IN;
  assign n15081 = ~n15039 | ~n15038;
  assign n15040 = ~SI_3_;
  assign n15041 = n15081 ^ ~n15040;
  assign n15044 = n15554 | n16024;
  assign n15042 = n15011 | n15904;
  assign n15089 = ~P1_IR_REG_3__SCAN_IN;
  assign n17949 = n15042 ^ ~n15089;
  assign n15043 = n16809 | n17949;
  assign n15045 = n15044 & n15043;
  assign n15047 = ~n15046 | ~n23941;
  assign n15051 = n15167 | n18575;
  assign n15050 = ~n13133 | ~n14281;
  assign n15057 = ~n15051 | ~n15050;
  assign n15053 = ~n15052;
  assign n23220 = ~n15054 | ~n15053;
  assign n15055 = n23222 & n23220;
  assign n23225 = ~n23221 | ~n15055;
  assign n15058 = ~n15056;
  assign n15060 = ~n15936 | ~P1_REG1_REG_4__SCAN_IN;
  assign n15059 = ~n13129 | ~P1_REG0_REG_4__SCAN_IN;
  assign n15068 = ~n15060 | ~n15059;
  assign n15066 = ~n15530 | ~P1_REG2_REG_4__SCAN_IN;
  assign n15061 = ~P1_REG3_REG_4__SCAN_IN;
  assign n15063 = ~n15062 | ~n15061;
  assign n15157 = ~P1_REG3_REG_4__SCAN_IN | ~P1_REG3_REG_3__SCAN_IN;
  assign n23919 = ~n15063 | ~n15157;
  assign n15064 = ~n23919;
  assign n15065 = ~n13130 | ~n15064;
  assign n15067 = ~n15066 | ~n15065;
  assign n15100 = n15167 | n23266;
  assign n17207 = ~SI_2_;
  assign n15071 = n15070 | SI_1_;
  assign n15076 = ~n15072 & ~n15078;
  assign n15075 = ~n15074 | ~n15073;
  assign n15084 = ~n15076 | ~n15075;
  assign n15080 = n15077 & SI_2_;
  assign n15079 = ~n15078;
  assign n15083 = ~n15080 | ~n15079;
  assign n15082 = ~n15081 | ~SI_3_;
  assign n15087 = ~n15085 | ~P1_DATAO_REG_4__SCAN_IN;
  assign n15086 = ~n13128 | ~P2_DATAO_REG_4__SCAN_IN;
  assign n15088 = ~SI_4_;
  assign n25354 = n15111 ^ ~n15112;
  assign n15099 = n25354 | n15450;
  assign n15097 = n13126 | n16027;
  assign n15094 = ~n15011 | ~n15089;
  assign n15090 = ~n15094 | ~P1_IR_REG_31__SCAN_IN;
  assign n15093 = ~n15090 | ~P1_IR_REG_4__SCAN_IN;
  assign n15091 = ~P1_IR_REG_4__SCAN_IN;
  assign n15092 = ~n15091 | ~P1_IR_REG_31__SCAN_IN;
  assign n15095 = ~n15093 | ~n15092;
  assign n15142 = n15094 | P1_IR_REG_4__SCAN_IN;
  assign n24101 = ~n15095 | ~n15142;
  assign n15096 = n16809 | n24101;
  assign n15098 = n15097 & n15096;
  assign n24165 = ~n23903;
  assign n23265 = n15823 | n24165;
  assign n15130 = n15100 & n23265;
  assign n23271 = ~n23264 | ~n15130;
  assign n15101 = n15860 | n24165;
  assign n15103 = ~n15102 | ~n15101;
  assign n23293 = n15103 ^ ~n15647;
  assign n15104 = ~n23264 | ~n23293;
  assign n15128 = ~n23271 | ~n15104;
  assign n15106 = ~n15530 | ~P1_REG2_REG_5__SCAN_IN;
  assign n15105 = ~n13129 | ~P1_REG0_REG_5__SCAN_IN;
  assign n15110 = ~n15106 | ~n15105;
  assign n23867 = n15157 ^ ~P1_REG3_REG_5__SCAN_IN;
  assign n15108 = ~n13130 | ~n23867;
  assign n15107 = ~n15219 | ~P1_REG1_REG_5__SCAN_IN;
  assign n15109 = ~n15108 | ~n15107;
  assign n15124 = n23906 | n15823;
  assign n15114 = ~n15113 | ~SI_4_;
  assign n15116 = ~n15085 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n15115 = ~n17196 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n15117 = ~SI_5_;
  assign n15120 = n13127 | n16031;
  assign n15118 = ~n15142 | ~P1_IR_REG_31__SCAN_IN;
  assign n15143 = ~P1_IR_REG_5__SCAN_IN;
  assign n23444 = n15118 ^ ~n15143;
  assign n15119 = n16809 | n23444;
  assign n15121 = n15120 & n15119;
  assign n15125 = ~n15124 | ~n15123;
  assign n15127 = n15167 | n23906;
  assign n15126 = n15823 | n23872;
  assign n15131 = ~n15127 | ~n15126;
  assign n15137 = ~n23225 | ~n15129;
  assign n15135 = ~n14873 | ~n23274;
  assign n15132 = ~n15131;
  assign n15134 = ~n15133 | ~n15132;
  assign n15136 = n15135 & n15134;
  assign n15170 = ~n23336;
  assign n15141 = ~n16232 | ~P1_DATAO_REG_6__SCAN_IN;
  assign n15140 = ~n13128 | ~P2_DATAO_REG_6__SCAN_IN;
  assign n15176 = ~n15141 | ~n15140;
  assign n15155 = n25348 | n15810;
  assign n15153 = n15451 | n16034;
  assign n15144 = ~n15142;
  assign n15145 = ~n15144 | ~n15143;
  assign n15146 = ~n15145 | ~P1_IR_REG_31__SCAN_IN;
  assign n15149 = ~n15146 | ~P1_IR_REG_6__SCAN_IN;
  assign n15147 = ~P1_IR_REG_6__SCAN_IN;
  assign n15148 = ~n15147 | ~P1_IR_REG_31__SCAN_IN;
  assign n15151 = ~n15149 | ~n15148;
  assign n15150 = ~n15454;
  assign n24096 = ~n15151 | ~n15150;
  assign n15152 = n16809 | n24096;
  assign n15154 = n15153 & n15152;
  assign n15165 = n23845 | n15860;
  assign n15186 = ~n15530;
  assign n15159 = ~n15251 | ~P1_REG2_REG_6__SCAN_IN;
  assign n23842 = n15189 ^ ~n13538;
  assign n15158 = ~n13131 | ~n23842;
  assign n15163 = ~n15159 | ~n15158;
  assign n15669 = n15219;
  assign n15161 = ~n15669 | ~P1_REG1_REG_6__SCAN_IN;
  assign n15160 = ~n13129 | ~P1_REG0_REG_6__SCAN_IN;
  assign n15162 = ~n15161 | ~n15160;
  assign n23875 = n15163 | n15162;
  assign n15164 = n23278 | n15823;
  assign n15166 = ~n15165 | ~n15164;
  assign n15171 = n15166 ^ ~n15647;
  assign n15169 = n15167 | n23278;
  assign n15168 = n23845 | n15823;
  assign n15172 = n15169 & n15168;
  assign n15174 = ~n15171;
  assign n15173 = ~n15172;
  assign n23337 = ~n15174 | ~n15173;
  assign n15177 = ~n15176 | ~SI_6_;
  assign n15179 = ~n15085 | ~P1_DATAO_REG_7__SCAN_IN;
  assign n15178 = ~n17036 | ~P2_DATAO_REG_7__SCAN_IN;
  assign n15207 = ~n15179 | ~n15178;
  assign n15180 = ~SI_7_;
  assign n15184 = n15451 | n16037;
  assign n15182 = n15454 | n15904;
  assign n23486 = n15182 ^ ~n15212;
  assign n15183 = n16809 | n23486;
  assign n15185 = n15184 & n15183;
  assign n15195 = ~n23818 | ~n15046;
  assign n15251 = ~n15186;
  assign n15188 = ~n15251 | ~P1_REG2_REG_7__SCAN_IN;
  assign n15187 = ~n18512 | ~P1_REG0_REG_7__SCAN_IN;
  assign n15193 = ~n15188 | ~n15187;
  assign n23815 = n15222 ^ ~P1_REG3_REG_7__SCAN_IN;
  assign n15191 = ~n13130 | ~n23815;
  assign n15190 = ~n15936 | ~P1_REG1_REG_7__SCAN_IN;
  assign n15192 = ~n15191 | ~n15190;
  assign n23234 = ~n23853;
  assign n15194 = n23234 | n15823;
  assign n15196 = ~n15195 | ~n15194;
  assign n15199 = n15196 ^ ~n15647;
  assign n15198 = n15167 | n23234;
  assign n15197 = ~n23818 | ~n13134;
  assign n15200 = n15198 & n15197;
  assign n15204 = ~n15199 & ~n15200;
  assign n15202 = ~n15199;
  assign n15201 = ~n15200;
  assign n15203 = ~n15202 & ~n15201;
  assign n15205 = ~n15204;
  assign n15264 = ~n15207 | ~SI_7_;
  assign n15211 = ~n15268 | ~n15264;
  assign n15209 = ~n15085 | ~P1_DATAO_REG_8__SCAN_IN;
  assign n15208 = ~n17036 | ~P2_DATAO_REG_8__SCAN_IN;
  assign n15210 = ~n15209 | ~n15208;
  assign n15265 = ~n15210 | ~SI_8_;
  assign n15238 = n15269 & n15265;
  assign n25335 = n15211 ^ ~n15238;
  assign n15218 = n25335 | n15810;
  assign n15216 = n15451 | n16039;
  assign n15318 = ~n15454 | ~n15212;
  assign n15214 = ~n15318 | ~P1_IR_REG_31__SCAN_IN;
  assign n15213 = ~P1_IR_REG_8__SCAN_IN;
  assign n24091 = n15214 ^ ~n15213;
  assign n15215 = n16809 | n24091;
  assign n15217 = n15216 & n15215;
  assign n15231 = ~n24213 | ~n15046;
  assign n15221 = ~n15936 | ~P1_REG1_REG_8__SCAN_IN;
  assign n15220 = ~n18512 | ~P1_REG0_REG_8__SCAN_IN;
  assign n15229 = ~n15221 | ~n15220;
  assign n15227 = ~n15391 | ~P1_REG2_REG_8__SCAN_IN;
  assign n15224 = n15223 & n23235;
  assign n23805 = n15224 | n15252;
  assign n15225 = ~n23805;
  assign n15226 = ~n13130 | ~n15225;
  assign n15228 = ~n15227 | ~n15226;
  assign n17396 = ~n23825;
  assign n15230 = n17396 | n15823;
  assign n15232 = ~n15231 | ~n15230;
  assign n15236 = n15232 ^ ~n15859;
  assign n15234 = ~n24213 | ~n13133;
  assign n15233 = ~n15766 | ~n23825;
  assign n15235 = ~n15234 | ~n15233;
  assign n23237 = n15236 ^ ~n15235;
  assign n15237 = ~n15236 & ~n15235;
  assign n15239 = n15238 & n15264;
  assign n15241 = ~n13122 | ~P1_DATAO_REG_9__SCAN_IN;
  assign n15240 = ~n13128 | ~P2_DATAO_REG_9__SCAN_IN;
  assign n15243 = ~n15242 | ~SI_9_;
  assign n15247 = n15451 | n24084;
  assign n15245 = n15318 | P1_IR_REG_8__SCAN_IN;
  assign n15279 = ~n15245 | ~P1_IR_REG_31__SCAN_IN;
  assign n24088 = n15279 ^ ~P1_IR_REG_9__SCAN_IN;
  assign n15246 = ~n15553 | ~n24088;
  assign n15248 = n15247 & n15246;
  assign n15260 = ~n24231 | ~n15046;
  assign n15250 = ~n15669 | ~P1_REG1_REG_9__SCAN_IN;
  assign n15249 = ~n13129 | ~P1_REG0_REG_9__SCAN_IN;
  assign n15258 = ~n15250 | ~n15249;
  assign n15256 = ~n15251 | ~P1_REG2_REG_9__SCAN_IN;
  assign n15253 = ~n15252 & ~P1_REG3_REG_9__SCAN_IN;
  assign n23789 = n15288 | n15253;
  assign n15254 = ~n23789;
  assign n15255 = ~n13131 | ~n15254;
  assign n15257 = ~n15256 | ~n15255;
  assign n23241 = ~n23801;
  assign n15259 = n23241 | n15823;
  assign n15261 = ~n15260 | ~n15259;
  assign n23308 = n15261 ^ ~n15859;
  assign n15263 = ~n24231 | ~n13134;
  assign n15262 = n15167 | n23241;
  assign n22199 = ~n15263 | ~n15262;
  assign n15299 = ~n23308 | ~n22199;
  assign n15266 = ~n15265 | ~n15264;
  assign n15272 = ~n15271;
  assign n15274 = ~n15273 & ~n15272;
  assign n15276 = ~n13121 | ~P1_DATAO_REG_10__SCAN_IN;
  assign n15275 = ~n21363 | ~P2_DATAO_REG_10__SCAN_IN;
  assign n15277 = n15309 ^ ~SI_10_;
  assign n15285 = n25325 | n15810;
  assign n15283 = n15451 | n24078;
  assign n15278 = ~P1_IR_REG_9__SCAN_IN;
  assign n15280 = ~n15279 | ~n15278;
  assign n15281 = ~n15280 | ~P1_IR_REG_31__SCAN_IN;
  assign n24081 = n15281 ^ ~P1_IR_REG_10__SCAN_IN;
  assign n15282 = ~n24081 | ~n15553;
  assign n15284 = n15283 & n15282;
  assign n15295 = ~n18649 | ~n15046;
  assign n15287 = ~n15669 | ~P1_REG1_REG_10__SCAN_IN;
  assign n15286 = ~n18512 | ~P1_REG0_REG_10__SCAN_IN;
  assign n15293 = ~n15287 | ~n15286;
  assign n15289 = n15288 | P1_REG3_REG_10__SCAN_IN;
  assign n22209 = n15353 & n15289;
  assign n15291 = ~n13131 | ~n22209;
  assign n15290 = ~n15391 | ~P1_REG2_REG_10__SCAN_IN;
  assign n15292 = ~n15291 | ~n15290;
  assign n15294 = n14344 | n15823;
  assign n15296 = ~n15295 | ~n15294;
  assign n22203 = n15296 ^ ~n15859;
  assign n15298 = ~n18649 | ~n13134;
  assign n15297 = n15167 | n14344;
  assign n22202 = ~n15298 | ~n15297;
  assign n22367 = ~n22203 | ~n22202;
  assign n15300 = ~n15299 | ~n22367;
  assign n15301 = ~n22202;
  assign n15306 = ~n15302 | ~n15301;
  assign n15303 = ~n22203;
  assign n15305 = ~n15304 | ~n15303;
  assign n15307 = ~n15306 | ~n15305;
  assign n15310 = ~n15309 | ~SI_10_;
  assign n15312 = ~n13122 | ~P1_DATAO_REG_11__SCAN_IN;
  assign n15311 = ~n17196 | ~P2_DATAO_REG_11__SCAN_IN;
  assign n15313 = ~n15312 | ~n15311;
  assign n15314 = ~n15313 | ~SI_11_;
  assign n25320 = n15337 ^ ~n15338;
  assign n15321 = n15451 | n24072;
  assign n15316 = ~P1_IR_REG_10__SCAN_IN;
  assign n15317 = ~n15315 | ~n15316;
  assign n15319 = ~n15344 | ~P1_IR_REG_31__SCAN_IN;
  assign n24075 = n15319 ^ ~P1_IR_REG_11__SCAN_IN;
  assign n15320 = ~n15553 | ~n24075;
  assign n15322 = n15321 & n15320;
  assign n15331 = ~n23051 | ~n15046;
  assign n15325 = ~n15669 | ~P1_REG1_REG_11__SCAN_IN;
  assign n15324 = ~n18512 | ~P1_REG0_REG_11__SCAN_IN;
  assign n15329 = ~n15325 | ~n15324;
  assign n22376 = n15353 ^ ~P1_REG3_REG_11__SCAN_IN;
  assign n15327 = ~n13130 | ~n22376;
  assign n15326 = ~n15391 | ~P1_REG2_REG_11__SCAN_IN;
  assign n15328 = ~n15327 | ~n15326;
  assign n22207 = ~n23753;
  assign n15330 = n22207 | n15823;
  assign n15332 = ~n15331 | ~n15330;
  assign n15336 = n15332 ^ ~n15859;
  assign n15334 = ~n23051 | ~n13133;
  assign n15333 = ~n15766 | ~n23753;
  assign n15335 = ~n15334 | ~n15333;
  assign n22371 = n15336 ^ ~n15335;
  assign n15341 = ~n13122 | ~P1_DATAO_REG_12__SCAN_IN;
  assign n15340 = ~n13128 | ~P2_DATAO_REG_12__SCAN_IN;
  assign n15342 = ~n15341 | ~n15340;
  assign n15343 = ~n15342 | ~SI_12_;
  assign n15369 = ~n15371 | ~n15343;
  assign n24065 = n15370 ^ ~n15369;
  assign n15349 = n24065 | n15810;
  assign n15377 = ~n15344 & ~P1_IR_REG_11__SCAN_IN;
  assign n15345 = n15377 | n15904;
  assign n24069 = n15345 ^ ~P1_IR_REG_12__SCAN_IN;
  assign n15347 = ~n24069 | ~n15553;
  assign n15346 = n15451 | n24066;
  assign n15348 = n15347 & n15346;
  assign n22257 = n15349 & n15348;
  assign n15361 = ~n22257 & ~n15860;
  assign n15351 = ~n15669 | ~P1_REG1_REG_12__SCAN_IN;
  assign n15350 = ~n13129 | ~P1_REG0_REG_12__SCAN_IN;
  assign n15359 = n15351 & n15350;
  assign n15355 = ~n15354 | ~n22253;
  assign n17414 = ~n15387 | ~n15355;
  assign n22252 = ~n17414;
  assign n15357 = ~n13130 | ~n22252;
  assign n15356 = ~n15391 | ~P1_REG2_REG_12__SCAN_IN;
  assign n15358 = n15357 & n15356;
  assign n15360 = ~n15823 & ~n22790;
  assign n15362 = n15361 | n15360;
  assign n15365 = n15362 ^ ~n15647;
  assign n15364 = ~n18666 | ~n13134;
  assign n15363 = n15167 | n22790;
  assign n15366 = n15364 & n15363;
  assign n22247 = ~n15365 | ~n15366;
  assign n15368 = ~n15365;
  assign n15367 = ~n15366;
  assign n22248 = ~n15368 | ~n15367;
  assign n15374 = ~n13122 | ~P1_DATAO_REG_13__SCAN_IN;
  assign n15373 = ~n13128 | ~P2_DATAO_REG_13__SCAN_IN;
  assign n15405 = ~n15408 | ~n15375;
  assign n25311 = n15405 ^ ~n15407;
  assign n15383 = n25311 | n15810;
  assign n15376 = ~P1_IR_REG_12__SCAN_IN;
  assign n15378 = ~n15377 | ~n15376;
  assign n15412 = ~n15378 | ~P1_IR_REG_31__SCAN_IN;
  assign n24062 = n15412 ^ ~P1_IR_REG_13__SCAN_IN;
  assign n15381 = ~n24062 | ~n15553;
  assign n15379 = ~n15554;
  assign n15380 = n15451 | n24059;
  assign n15382 = n15381 & n15380;
  assign n15397 = ~n22341 | ~n15046;
  assign n15385 = ~n15669 | ~P1_REG1_REG_13__SCAN_IN;
  assign n15384 = ~n13129 | ~P1_REG0_REG_13__SCAN_IN;
  assign n15395 = n15385 & n15384;
  assign n15390 = ~n13131;
  assign n15419 = ~n15387 & ~n15386;
  assign n15389 = ~n15419;
  assign n15388 = ~n15387 | ~n15386;
  assign n22337 = ~n15389 | ~n15388;
  assign n15393 = n15390 | n22337;
  assign n15392 = ~n15391 | ~P1_REG2_REG_13__SCAN_IN;
  assign n15394 = n15393 & n15392;
  assign n23017 = ~n15395 | ~n15394;
  assign n22754 = ~n23017;
  assign n15396 = n22754 | n15823;
  assign n15398 = ~n15397 | ~n15396;
  assign n15401 = n15398 ^ ~n15647;
  assign n15400 = ~n22341 | ~n13133;
  assign n15399 = n15167 | n22754;
  assign n15402 = n15400 & n15399;
  assign n22333 = ~n15401 & ~n15402;
  assign n15404 = ~n15401;
  assign n15403 = ~n15402;
  assign n22332 = ~n15404 & ~n15403;
  assign n15406 = ~n15405;
  assign n16792 = ~SI_14_;
  assign n15440 = ~n15444 | ~n16792;
  assign n15410 = ~n13121 | ~P1_DATAO_REG_14__SCAN_IN;
  assign n21363 = n13128;
  assign n15409 = ~n21363 | ~P2_DATAO_REG_14__SCAN_IN;
  assign n15411 = ~P1_IR_REG_13__SCAN_IN;
  assign n15413 = ~n15412 | ~n15411;
  assign n15414 = ~n15413 | ~P1_IR_REG_31__SCAN_IN;
  assign n24056 = n15414 ^ ~P1_IR_REG_14__SCAN_IN;
  assign n15416 = ~n24056 | ~n15553;
  assign n15415 = n15451 | n24053;
  assign n15417 = n15416 & n15415;
  assign n15429 = ~n23015 & ~n15823;
  assign n15420 = n15419 | P1_REG3_REG_14__SCAN_IN;
  assign n15467 = ~n15419 | ~P1_REG3_REG_14__SCAN_IN;
  assign n22756 = n15420 & n15467;
  assign n15423 = ~n22756 | ~n13131;
  assign n15422 = ~n15391 | ~P1_REG2_REG_14__SCAN_IN;
  assign n15427 = n15423 & n15422;
  assign n15425 = ~n15669 | ~P1_REG1_REG_14__SCAN_IN;
  assign n15424 = ~n18512 | ~P1_REG0_REG_14__SCAN_IN;
  assign n15426 = n15425 & n15424;
  assign n23035 = ~n15427 | ~n15426;
  assign n22731 = ~n23035;
  assign n15428 = ~n15167 & ~n22731;
  assign n15433 = ~n15429 & ~n15428;
  assign n15431 = ~n18041 | ~n15046;
  assign n15430 = ~n13133 | ~n23035;
  assign n15432 = ~n15431 | ~n15430;
  assign n15435 = n15432 ^ ~n15859;
  assign n22171 = n15433 ^ n15435;
  assign n15434 = ~n15433;
  assign n15437 = ~n13122 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n15436 = ~n21363 | ~P2_DATAO_REG_15__SCAN_IN;
  assign n15438 = ~n15437 | ~n15436;
  assign n15439 = ~n15438 | ~SI_15_;
  assign n15447 = ~n15485 | ~n15439;
  assign n15441 = n15440 & n15447;
  assign n15449 = ~n15442 | ~n15441;
  assign n15465 = ~n17624 | ~n14654;
  assign n16884 = ~P2_DATAO_REG_15__SCAN_IN;
  assign n15463 = n15451 | n16884;
  assign n15453 = ~n15452;
  assign n15455 = ~n15454 | ~n15453;
  assign n15495 = ~n15455 & ~P1_IR_REG_15__SCAN_IN;
  assign n15461 = ~n15495;
  assign n15456 = ~n15455 | ~P1_IR_REG_31__SCAN_IN;
  assign n15459 = ~n15456 | ~P1_IR_REG_15__SCAN_IN;
  assign n15457 = ~P1_IR_REG_15__SCAN_IN;
  assign n15458 = ~n15457 | ~P1_IR_REG_31__SCAN_IN;
  assign n15460 = ~n15459 | ~n15458;
  assign n23632 = ~n23656;
  assign n15462 = n16809 | n23632;
  assign n15464 = n15463 & n15462;
  assign n15476 = ~n22998 & ~n15860;
  assign n15466 = ~P1_REG3_REG_15__SCAN_IN;
  assign n15468 = ~n15467 | ~n15466;
  assign n22732 = n13178 & n15468;
  assign n15470 = ~n22732 | ~n13130;
  assign n15469 = ~n15391 | ~P1_REG2_REG_15__SCAN_IN;
  assign n15474 = ~n15470 | ~n15469;
  assign n15472 = ~n15669 | ~P1_REG1_REG_15__SCAN_IN;
  assign n15471 = ~n13129 | ~P1_REG0_REG_15__SCAN_IN;
  assign n15473 = ~n15472 | ~n15471;
  assign n22176 = ~n15474 & ~n15473;
  assign n15475 = ~n22176 & ~n15823;
  assign n15477 = ~n15476 & ~n15475;
  assign n15482 = n15859 ^ n15477;
  assign n15478 = ~n15482;
  assign n22399 = ~n15481 | ~n15478;
  assign n18702 = ~n22998;
  assign n15480 = ~n18702 | ~n13133;
  assign n15479 = ~n15766 | ~n23016;
  assign n22401 = ~n15480 | ~n15479;
  assign n15484 = ~n22399 | ~n22401;
  assign n15483 = ~n15481;
  assign n22400 = ~n15483 | ~n15482;
  assign n22277 = ~n15484 | ~n22400;
  assign n15488 = ~n13121 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n15487 = ~n21363 | ~P2_DATAO_REG_16__SCAN_IN;
  assign n15489 = ~n15488 | ~n15487;
  assign n15490 = ~n15489 | ~SI_16_;
  assign n15516 = ~n15518 | ~n15490;
  assign n16056 = ~P2_DATAO_REG_16__SCAN_IN;
  assign n15498 = n15451 | n16056;
  assign n15491 = n15495 | n15904;
  assign n15493 = ~n15491 | ~P1_IR_REG_16__SCAN_IN;
  assign n15494 = ~P1_IR_REG_16__SCAN_IN;
  assign n15492 = ~n15494 | ~P1_IR_REG_31__SCAN_IN;
  assign n15496 = ~n15493 | ~n15492;
  assign n15523 = ~n15495 | ~n15494;
  assign n23678 = n15496 & n15523;
  assign n15497 = ~n15553 | ~n23678;
  assign n15499 = n15498 & n15497;
  assign n15510 = ~n22702 | ~n15046;
  assign n15501 = ~P1_REG3_REG_16__SCAN_IN;
  assign n15502 = n13178 & n15501;
  assign n22708 = ~n15559 & ~n15502;
  assign n15504 = ~n22708 | ~n13131;
  assign n15503 = ~n15391 | ~P1_REG2_REG_16__SCAN_IN;
  assign n15508 = ~n15504 | ~n15503;
  assign n15506 = ~n15669 | ~P1_REG1_REG_16__SCAN_IN;
  assign n15505 = ~n13129 | ~P1_REG0_REG_16__SCAN_IN;
  assign n15507 = ~n15506 | ~n15505;
  assign n15509 = ~n22999 | ~n13134;
  assign n15511 = ~n15510 | ~n15509;
  assign n15515 = n15511 ^ ~n15859;
  assign n15513 = ~n22702 | ~n13133;
  assign n15512 = ~n22999 | ~n15766;
  assign n15514 = ~n15513 | ~n15512;
  assign n22279 = n15515 ^ ~n15514;
  assign n15520 = ~n13121 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n15519 = ~n21363 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n15521 = ~n15520 | ~n15519;
  assign n15522 = ~n15521 | ~SI_17_;
  assign n15542 = ~n15546 | ~n15522;
  assign n25296 = n15544 ^ ~n15542;
  assign n15550 = ~n15523 | ~P1_IR_REG_31__SCAN_IN;
  assign n24044 = n15550 ^ ~P1_IR_REG_17__SCAN_IN;
  assign n15525 = ~n24044 | ~n15553;
  assign n24041 = ~P2_DATAO_REG_17__SCAN_IN;
  assign n15524 = n15451 | n24041;
  assign n15526 = n15525 & n15524;
  assign n15536 = ~n22295 | ~n15046;
  assign n22296 = n15559 ^ ~P1_REG3_REG_17__SCAN_IN;
  assign n15534 = n22296 | n15390;
  assign n15529 = ~n15669 | ~P1_REG1_REG_17__SCAN_IN;
  assign n15528 = ~n13129 | ~P1_REG0_REG_17__SCAN_IN;
  assign n15532 = ~n15529 | ~n15528;
  assign n15531 = n15391 & P1_REG2_REG_17__SCAN_IN;
  assign n15533 = ~n15532 & ~n15531;
  assign n22982 = ~n15534 | ~n15533;
  assign n15535 = ~n22982 | ~n13133;
  assign n15537 = ~n15536 | ~n15535;
  assign n15541 = n15537 ^ ~n15647;
  assign n15539 = ~n22295 | ~n13134;
  assign n15538 = ~n22982 | ~n15766;
  assign n15540 = n15539 & n15538;
  assign n22291 = ~n15541 | ~n15540;
  assign n22290 = n15541 | n15540;
  assign n15545 = SI_18_ & n15546;
  assign n18249 = ~SI_18_;
  assign n15548 = ~n13121 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n15547 = ~n21363 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n25290 = n15574 ^ ~n15573;
  assign n15549 = ~P1_IR_REG_31__SCAN_IN | ~P1_IR_REG_17__SCAN_IN;
  assign n15552 = ~n15550 | ~n15549;
  assign n15551 = ~P1_IR_REG_18__SCAN_IN;
  assign n23711 = n15552 ^ ~n15551;
  assign n15556 = ~n23711 | ~n15553;
  assign n17077 = ~P2_DATAO_REG_18__SCAN_IN;
  assign n15555 = n15451 | n17077;
  assign n15557 = n15556 & n15555;
  assign n15567 = ~n22664 | ~n15046;
  assign n22389 = P1_REG3_REG_18__SCAN_IN ^ n15585;
  assign n22665 = ~n22389;
  assign n15565 = ~n22665 | ~n13130;
  assign n15561 = ~n15936 | ~P1_REG1_REG_18__SCAN_IN;
  assign n15560 = ~n18512 | ~P1_REG0_REG_18__SCAN_IN;
  assign n15563 = ~n15561 | ~n15560;
  assign n22660 = ~P1_REG2_REG_18__SCAN_IN;
  assign n15562 = ~n15186 & ~n22660;
  assign n15564 = ~n15563 & ~n15562;
  assign n24289 = ~n15565 | ~n15564;
  assign n15566 = ~n24289 | ~n13134;
  assign n15568 = ~n15567 | ~n15566;
  assign n15572 = n15568 ^ ~n15859;
  assign n15570 = ~n22664 | ~n13133;
  assign n15569 = ~n24289 | ~n15766;
  assign n15571 = ~n15570 | ~n15569;
  assign n22387 = n15572 ^ ~n15571;
  assign n15576 = ~n13122 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n15575 = ~n21363 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n15578 = ~n15577 | ~SI_19_;
  assign n15583 = ~n17664 | ~n14654;
  assign n17271 = ~P2_DATAO_REG_19__SCAN_IN;
  assign n15581 = n15451 | n17271;
  assign n15580 = n16809 | n23905;
  assign n15582 = n15581 & n15580;
  assign n15593 = ~n22223 | ~n13133;
  assign n15584 = ~P1_REG3_REG_18__SCAN_IN;
  assign n22635 = P1_REG3_REG_19__SCAN_IN ^ n15610;
  assign n15591 = ~n22635 | ~n13131;
  assign n15587 = ~n15391 | ~P1_REG2_REG_19__SCAN_IN;
  assign n15586 = ~n15669 | ~P1_REG1_REG_19__SCAN_IN;
  assign n15589 = ~n15587 | ~n15586;
  assign n15588 = n18512 & P1_REG0_REG_19__SCAN_IN;
  assign n15590 = ~n15589 & ~n15588;
  assign n24292 = ~n15591 | ~n15590;
  assign n15592 = ~n24292 | ~n15766;
  assign n15597 = ~n15593 | ~n15592;
  assign n15595 = ~n22223 | ~n15046;
  assign n15594 = ~n24292 | ~n13134;
  assign n15596 = ~n15595 | ~n15594;
  assign n15598 = n15596 ^ ~n15859;
  assign n22218 = n15597 ^ n15598;
  assign n15599 = ~n15598 | ~n15597;
  assign n15601 = ~n15604 & ~SI_18_;
  assign n15607 = ~n13122 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n15606 = ~n21363 | ~P2_DATAO_REG_20__SCAN_IN;
  assign n17294 = ~P2_DATAO_REG_20__SCAN_IN;
  assign n15608 = n15451 | n17294;
  assign n15619 = ~n22618 | ~n15046;
  assign n15611 = ~P1_REG3_REG_20__SCAN_IN;
  assign n22612 = n15640 ^ ~n15611;
  assign n15617 = ~n22612 | ~n13131;
  assign n15613 = ~n15669 | ~P1_REG1_REG_20__SCAN_IN;
  assign n15612 = ~n18512 | ~P1_REG0_REG_20__SCAN_IN;
  assign n15615 = ~n15613 | ~n15612;
  assign n15614 = n15251 & P1_REG2_REG_20__SCAN_IN;
  assign n15616 = ~n15615 & ~n15614;
  assign n15618 = ~n24295 | ~n13133;
  assign n15620 = ~n15619 | ~n15618;
  assign n15623 = n15620 ^ ~n15647;
  assign n15622 = ~n22618 | ~n13134;
  assign n15621 = n22589 | n15167;
  assign n15624 = n15622 & n15621;
  assign n15626 = ~n15623;
  assign n15625 = ~n15624;
  assign n15627 = n15626 | n15625;
  assign n22319 = n15628 & n15627;
  assign n15632 = ~n15660 | ~SI_20_;
  assign n15634 = ~n13121 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n15633 = ~n21363 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n18271 = ~SI_21_;
  assign n15635 = n15664 ^ ~n18271;
  assign n17281 = ~P2_DATAO_REG_21__SCAN_IN;
  assign n15636 = n15451 | n17281;
  assign n15639 = ~n15669 | ~P1_REG1_REG_21__SCAN_IN;
  assign n15638 = ~n18512 | ~P1_REG0_REG_21__SCAN_IN;
  assign n15644 = ~n15639 | ~n15638;
  assign n22590 = P1_REG3_REG_21__SCAN_IN ^ ~n13214;
  assign n15642 = ~n13130 | ~n22590;
  assign n15641 = ~n15391 | ~P1_REG2_REG_21__SCAN_IN;
  assign n15643 = ~n15642 | ~n15641;
  assign n15645 = n13716 | n15823;
  assign n15648 = ~n15646 | ~n15645;
  assign n15653 = n15648 ^ ~n15647;
  assign n15649 = n15167 | n13716;
  assign n22233 = ~n15653 & ~n15654;
  assign n15651 = ~n22233;
  assign n15656 = ~n15653;
  assign n15655 = ~n15654;
  assign n22349 = ~n15656 & ~n15655;
  assign n15657 = ~n15661;
  assign n18268 = ~SI_20_;
  assign n15658 = ~n15657 | ~n18268;
  assign n15663 = n15661 & SI_20_;
  assign n15666 = ~n15663 | ~n15662;
  assign n15665 = ~n15664 | ~SI_21_;
  assign n15677 = n22889 | n15860;
  assign n22356 = P1_REG3_REG_22__SCAN_IN ^ ~n15697;
  assign n15675 = ~n22356 | ~n13131;
  assign n15671 = ~n15251 | ~P1_REG2_REG_22__SCAN_IN;
  assign n15670 = ~n15669 | ~P1_REG1_REG_22__SCAN_IN;
  assign n15673 = ~n15671 | ~n15670;
  assign n15672 = n18512 & P1_REG0_REG_22__SCAN_IN;
  assign n15674 = ~n15673 & ~n15672;
  assign n15676 = ~n24301 | ~n13134;
  assign n15678 = ~n15677 | ~n15676;
  assign n15683 = n15678 ^ ~n15859;
  assign n15681 = ~n15683;
  assign n15680 = ~n22889 & ~n15823;
  assign n15679 = ~n22551 & ~n15167;
  assign n15682 = ~n15680 & ~n15679;
  assign n15684 = n15681 & n15682;
  assign n22351 = n15683 ^ ~n15682;
  assign n15685 = n15684 | n22351;
  assign n15687 = ~n13121 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n15686 = ~n21363 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n15688 = ~n15717 | ~SI_22_;
  assign n15691 = ~n13121 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n15690 = ~n21363 | ~P2_DATAO_REG_23__SCAN_IN;
  assign n15721 = ~n15691 | ~n15690;
  assign n15692 = n15721 ^ ~SI_23_;
  assign n17718 = n15693 ^ ~n15692;
  assign n15695 = ~n17718 | ~n14654;
  assign n17451 = ~P2_DATAO_REG_23__SCAN_IN;
  assign n15694 = n15451 | n17451;
  assign n15706 = ~n22874 & ~n15860;
  assign n15696 = ~P1_REG3_REG_22__SCAN_IN;
  assign n22550 = P1_REG3_REG_23__SCAN_IN ^ ~n15730;
  assign n15698 = ~n22550;
  assign n15704 = ~n15698 | ~n13130;
  assign n15700 = ~n15936 | ~P1_REG1_REG_23__SCAN_IN;
  assign n15699 = ~n13129 | ~P1_REG0_REG_23__SCAN_IN;
  assign n15702 = ~n15700 | ~n15699;
  assign n15701 = n15251 & P1_REG2_REG_23__SCAN_IN;
  assign n15703 = ~n15702 & ~n15701;
  assign n15705 = ~n22516 & ~n15823;
  assign n15707 = ~n15706 & ~n15705;
  assign n15712 = n15707 ^ ~n15859;
  assign n15709 = n22874 | n15823;
  assign n15708 = ~n24304 | ~n15766;
  assign n15710 = ~n15709 | ~n15708;
  assign n15711 = ~n15710;
  assign n15713 = ~n15712 | ~n15711;
  assign n15714 = ~SI_22_;
  assign n15715 = ~n17345 | ~n15714;
  assign n15718 = ~n17345;
  assign n15720 = n15718 & SI_22_;
  assign n15723 = ~n15720 | ~n15719;
  assign n15722 = ~n15721 | ~SI_23_;
  assign n15726 = ~n13121 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n15725 = ~n21363 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n15748 = ~n15726 | ~n15725;
  assign n15727 = n15748 ^ ~n14137;
  assign n17732 = n15749 ^ ~n15727;
  assign n15729 = n17732 | n15810;
  assign n17331 = ~P2_DATAO_REG_24__SCAN_IN;
  assign n15728 = n15451 | n17331;
  assign n15739 = ~n22862 | ~n15046;
  assign n15731 = ~P1_REG3_REG_24__SCAN_IN;
  assign n22527 = n15758 ^ ~n15731;
  assign n15737 = ~n22527 | ~n13131;
  assign n15733 = ~n15936 | ~P1_REG1_REG_24__SCAN_IN;
  assign n15732 = ~n13129 | ~P1_REG0_REG_24__SCAN_IN;
  assign n15735 = ~n15733 | ~n15732;
  assign n15734 = n15391 & P1_REG2_REG_24__SCAN_IN;
  assign n15736 = ~n15735 & ~n15734;
  assign n15738 = ~n24308 | ~n13133;
  assign n15740 = ~n15739 | ~n15738;
  assign n15743 = n15740 ^ ~n15859;
  assign n15742 = ~n22535 & ~n15823;
  assign n18031 = ~n24308;
  assign n15741 = ~n18031 & ~n15167;
  assign n15744 = ~n15742 & ~n15741;
  assign n22307 = n15743 ^ ~n15744;
  assign n15747 = ~n22306 | ~n22307;
  assign n15745 = ~n15743;
  assign n15746 = ~n15745 | ~n15744;
  assign n15753 = ~n13121 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n15752 = ~n21363 | ~P2_DATAO_REG_25__SCAN_IN;
  assign n15754 = ~n15753 | ~n15752;
  assign n15755 = ~n15754 | ~SI_25_;
  assign n23159 = ~P2_DATAO_REG_25__SCAN_IN;
  assign n15756 = n15451 | n23159;
  assign n15768 = ~n22495 | ~n13134;
  assign n22496 = P1_REG3_REG_25__SCAN_IN ^ ~n15788;
  assign n15759 = ~n22496;
  assign n15765 = ~n15759 | ~n13130;
  assign n15761 = ~n15936 | ~P1_REG1_REG_25__SCAN_IN;
  assign n15760 = ~n18512 | ~P1_REG0_REG_25__SCAN_IN;
  assign n15763 = ~n15761 | ~n15760;
  assign n15762 = n15391 & P1_REG2_REG_25__SCAN_IN;
  assign n15764 = ~n15763 & ~n15762;
  assign n15767 = ~n24311 | ~n15766;
  assign n15773 = ~n15768 | ~n15767;
  assign n15770 = ~n22495 | ~n15046;
  assign n15769 = ~n24311 | ~n13134;
  assign n15771 = ~n15770 | ~n15769;
  assign n15772 = n15771 ^ ~n15859;
  assign n22265 = n15773 ^ n15772;
  assign n15775 = ~n15772;
  assign n15774 = ~n15773;
  assign n15776 = ~n15775 | ~n15774;
  assign n15779 = ~n13122 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n15778 = ~n21363 | ~P2_DATAO_REG_26__SCAN_IN;
  assign n15780 = ~n15779 | ~n15778;
  assign n15804 = n15780 | SI_26_;
  assign n15827 = ~n15780 | ~SI_26_;
  assign n15782 = ~n15804 | ~n15827;
  assign n15786 = ~n15781 | ~n15782;
  assign n15783 = ~n15782;
  assign n15785 = ~n15784 | ~n15783;
  assign n23151 = ~P2_DATAO_REG_26__SCAN_IN;
  assign n15787 = n15451 | n23151;
  assign n15796 = ~n18805 | ~n13132;
  assign n17997 = ~P1_REG3_REG_26__SCAN_IN;
  assign n22474 = n15815 ^ ~n17997;
  assign n15794 = ~n22474 | ~n13130;
  assign n15790 = ~n15936 | ~P1_REG1_REG_26__SCAN_IN;
  assign n15789 = ~n18512 | ~P1_REG0_REG_26__SCAN_IN;
  assign n15792 = ~n15790 | ~n15789;
  assign n15791 = n15251 & P1_REG2_REG_26__SCAN_IN;
  assign n15793 = ~n15792 & ~n15791;
  assign n15795 = ~n14111 | ~n13133;
  assign n15797 = ~n15796 | ~n15795;
  assign n15800 = n15797 ^ ~n15859;
  assign n15799 = ~n18805 | ~n13134;
  assign n15798 = n22847 | n15167;
  assign n15801 = ~n15799 | ~n15798;
  assign n17995 = ~n15800 | ~n15801;
  assign n15803 = ~n15800;
  assign n15802 = ~n15801;
  assign n17996 = ~n15803 | ~n15802;
  assign n15833 = n15805 & n15804;
  assign n15807 = ~n15806 | ~n15833;
  assign n15809 = ~n13121 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n15808 = ~n21363 | ~P2_DATAO_REG_27__SCAN_IN;
  assign n15837 = ~n15809 | ~n15808;
  assign n23144 = ~P2_DATAO_REG_27__SCAN_IN;
  assign n15811 = n15451 | n23144;
  assign n15822 = ~n22819 | ~n13133;
  assign n15814 = ~n15669 | ~P1_REG1_REG_27__SCAN_IN;
  assign n15813 = ~n13129 | ~P1_REG0_REG_27__SCAN_IN;
  assign n15820 = ~n15814 | ~n15813;
  assign n15816 = ~n15851;
  assign n19108 = P1_REG3_REG_27__SCAN_IN ^ ~n15816;
  assign n15818 = ~n13131 | ~n19108;
  assign n15817 = ~n15251 | ~P1_REG2_REG_27__SCAN_IN;
  assign n15819 = ~n15818 | ~n15817;
  assign n15821 = n15167 | n18062;
  assign n15915 = ~n15822 | ~n15821;
  assign n15825 = ~n22819 | ~n13132;
  assign n15824 = n18062 | n15823;
  assign n15826 = ~n15825 | ~n15824;
  assign n15916 = n15826 ^ ~n15859;
  assign n19102 = n15915 ^ n15916;
  assign n15831 = ~n15837 & ~SI_27_;
  assign n15829 = n15828 & n15830;
  assign n15835 = ~n15830;
  assign n15832 = ~n15831;
  assign n15834 = n15833 & n15832;
  assign n15838 = ~n15837 | ~SI_27_;
  assign n15840 = ~n13121 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n15839 = ~n21363 | ~P2_DATAO_REG_28__SCAN_IN;
  assign n15841 = ~n15840 | ~n15839;
  assign n15842 = ~n15841 | ~SI_28_;
  assign n15844 = ~n15843;
  assign n15846 = ~n15845 | ~n15844;
  assign n15848 = ~n23137 | ~n14654;
  assign n18361 = ~P2_DATAO_REG_28__SCAN_IN;
  assign n15847 = n15451 | n18361;
  assign n15857 = ~n19092 & ~n15823;
  assign n15850 = ~n15936 | ~P1_REG1_REG_28__SCAN_IN;
  assign n15849 = ~n18512 | ~P1_REG0_REG_28__SCAN_IN;
  assign n15855 = ~n15850 | ~n15849;
  assign n15853 = ~n13130 | ~n18070;
  assign n15852 = ~n15391 | ~P1_REG2_REG_28__SCAN_IN;
  assign n15854 = ~n15853 | ~n15852;
  assign n15856 = ~n15167 & ~n22452;
  assign n15858 = ~n15857 & ~n15856;
  assign n15864 = n15859 ^ n15858;
  assign n15862 = ~n19092 & ~n15860;
  assign n15861 = ~n22452 & ~n15823;
  assign n15863 = ~n15862 & ~n15861;
  assign n15921 = n15864 ^ ~n15863;
  assign n15868 = ~n15866 | ~P1_B_REG_SCAN_IN;
  assign n15869 = ~n15868 | ~n15867;
  assign n15877 = ~P1_D_REG_6__SCAN_IN & ~P1_D_REG_7__SCAN_IN;
  assign n15875 = P1_D_REG_8__SCAN_IN | P1_D_REG_9__SCAN_IN;
  assign n15873 = ~P1_D_REG_10__SCAN_IN & ~P1_D_REG_11__SCAN_IN;
  assign n15872 = ~P1_D_REG_12__SCAN_IN & ~P1_D_REG_13__SCAN_IN;
  assign n15874 = ~n15873 | ~n15872;
  assign n15876 = ~n15875 & ~n15874;
  assign n15893 = ~n15877 | ~n15876;
  assign n15879 = ~P1_D_REG_18__SCAN_IN & ~P1_D_REG_19__SCAN_IN;
  assign n15878 = ~P1_D_REG_20__SCAN_IN & ~P1_D_REG_21__SCAN_IN;
  assign n15883 = ~n15879 | ~n15878;
  assign n15881 = ~P1_D_REG_16__SCAN_IN & ~P1_D_REG_14__SCAN_IN;
  assign n15880 = ~P1_D_REG_15__SCAN_IN & ~P1_D_REG_17__SCAN_IN;
  assign n15882 = ~n15881 | ~n15880;
  assign n15891 = ~n15883 & ~n15882;
  assign n15885 = ~P1_D_REG_26__SCAN_IN & ~P1_D_REG_27__SCAN_IN;
  assign n15884 = ~P1_D_REG_28__SCAN_IN & ~P1_D_REG_31__SCAN_IN;
  assign n15889 = ~n15885 | ~n15884;
  assign n15887 = ~P1_D_REG_22__SCAN_IN & ~P1_D_REG_23__SCAN_IN;
  assign n15886 = ~P1_D_REG_24__SCAN_IN & ~P1_D_REG_25__SCAN_IN;
  assign n15888 = ~n15887 | ~n15886;
  assign n15890 = ~n15889 & ~n15888;
  assign n15892 = ~n15891 | ~n15890;
  assign n15898 = ~n15893 & ~n15892;
  assign n15895 = ~P1_D_REG_2__SCAN_IN & ~P1_D_REG_3__SCAN_IN;
  assign n15894 = ~P1_D_REG_4__SCAN_IN & ~P1_D_REG_5__SCAN_IN;
  assign n15896 = ~n15895 | ~n15894;
  assign n15897 = ~P1_D_REG_30__SCAN_IN & ~n15896;
  assign n15899 = ~n15898 | ~n15897;
  assign n15900 = ~P1_D_REG_29__SCAN_IN & ~n15899;
  assign n17438 = ~n24034 & ~n15900;
  assign n24117 = n15865 | n15901;
  assign n15902 = P1_D_REG_1__SCAN_IN | n24034;
  assign n17434 = ~n24117 | ~n15902;
  assign n17408 = ~n17438 & ~n17434;
  assign n15903 = ~n17408;
  assign n15906 = n15905 | n15904;
  assign n15909 = ~n15906 | ~P1_IR_REG_23__SCAN_IN;
  assign n15908 = ~n15907 | ~P1_IR_REG_31__SCAN_IN;
  assign n15910 = ~n15909 | ~n15908;
  assign n16808 = ~n15911 | ~n15910;
  assign n15922 = ~n15931 & ~n24033;
  assign n15913 = ~n24230 & ~n17377;
  assign n23339 = n15922 & n15913;
  assign n15914 = ~n15921 | ~n23339;
  assign n15919 = n15916 | n15915;
  assign n15917 = ~n15919 | ~n23339;
  assign n15918 = ~n15921 & ~n15917;
  assign n15920 = ~n15919 & ~n23309;
  assign n15951 = ~n15921 | ~n15920;
  assign n23931 = ~n24123 | ~n18860;
  assign n23966 = ~n23931;
  assign n15924 = ~n15922 | ~n23966;
  assign n15923 = n18853 & n23723;
  assign n17436 = ~n24228 | ~n18861;
  assign n15949 = ~n19092 & ~n23277;
  assign n15927 = ~n18856 & ~n15925;
  assign n15926 = ~n16808;
  assign n15928 = ~n15927 & ~n15926;
  assign n16972 = ~n15931 | ~n17436;
  assign n15929 = ~n15930 | ~n16972;
  assign n15947 = ~n23343 | ~n18070;
  assign n15932 = ~n18907 | ~n17377;
  assign n23217 = ~n15932 & ~n15931;
  assign n23391 = ~n23351;
  assign n15935 = ~n23322 | ~n24316;
  assign n15934 = ~P1_U3086 | ~P1_REG3_REG_28__SCAN_IN;
  assign n15945 = ~n15935 | ~n15934;
  assign n23279 = ~n23217 | ~n23351;
  assign n15938 = ~n15936 | ~P1_REG1_REG_29__SCAN_IN;
  assign n15937 = ~n18512 | ~P1_REG0_REG_29__SCAN_IN;
  assign n15943 = n15938 & n15937;
  assign n15941 = ~n15391 | ~P1_REG2_REG_29__SCAN_IN;
  assign n22432 = ~n15939 | ~P1_REG3_REG_28__SCAN_IN;
  assign n15940 = n15390 | n22432;
  assign n15942 = n15941 & n15940;
  assign n15944 = ~n23279 & ~n18863;
  assign n15946 = ~n15945 & ~n15944;
  assign n15948 = ~n15947 | ~n15946;
  assign n15950 = ~n15949 & ~n15948;
  assign n15952 = n15951 & n15950;
  assign n15954 = ~P2_IR_REG_9__SCAN_IN & ~P2_IR_REG_11__SCAN_IN;
  assign n15956 = n15954 & n15953;
  assign n17596 = ~n15956 | ~n15955;
  assign n16568 = ~n15958 | ~n15957;
  assign n16565 = ~n15963 | ~n15962;
  assign n15964 = ~n17021;
  assign n15974 = ~n15964 | ~n16572;
  assign n15969 = ~n15968;
  assign n15971 = ~n15969 | ~P2_IR_REG_25__SCAN_IN;
  assign n15972 = ~n15979 | ~P2_IR_REG_31__SCAN_IN;
  assign n15973 = ~n22165 & ~n17324;
  assign n17011 = ~n22156 | ~n15973;
  assign n15975 = ~n15974 | ~P2_IR_REG_31__SCAN_IN;
  assign n15978 = ~n15975 | ~P2_IR_REG_23__SCAN_IN;
  assign n15976 = ~P2_IR_REG_23__SCAN_IN;
  assign n15977 = ~n15976 | ~P2_IR_REG_31__SCAN_IN;
  assign n15980 = ~n15978 | ~n15977;
  assign n17447 = ~n15980 | ~n15979;
  assign n21339 = ~n17447;
  assign n15982 = ~P3_IR_REG_8__SCAN_IN & ~P3_IR_REG_6__SCAN_IN;
  assign n15981 = ~P3_IR_REG_7__SCAN_IN & ~P3_IR_REG_10__SCAN_IN;
  assign n15985 = ~n15982 | ~n15981;
  assign n15984 = ~n15983 | ~n16146;
  assign n16132 = n19806 & n15986;
  assign n16009 = ~n15987 | ~n16132;
  assign n15997 = ~n16009;
  assign n15989 = ~P3_IR_REG_15__SCAN_IN & ~P3_IR_REG_13__SCAN_IN;
  assign n16010 = ~n15989 | ~n15988;
  assign n16012 = ~n15990 | ~n16960;
  assign n15995 = ~n16010 & ~n16012;
  assign n16011 = ~n15991 | ~n16326;
  assign n15993 = ~n15992 | ~n17143;
  assign n15994 = ~n16011 & ~n15993;
  assign n15996 = n15995 & n15994;
  assign n16001 = ~n16000 | ~P3_IR_REG_31__SCAN_IN;
  assign n16007 = ~n20794;
  assign n16005 = ~n16002 | ~P3_IR_REG_24__SCAN_IN;
  assign n16004 = ~n16003 | ~P3_IR_REG_31__SCAN_IN;
  assign n16006 = ~n16005 | ~n16004;
  assign n16287 = ~n16006 | ~n16000;
  assign n20802 = ~n16287;
  assign n19831 = ~n16286 | ~n16008;
  assign n16016 = ~n19831;
  assign n16955 = n16009;
  assign n16013 = ~n16954 & ~n16012;
  assign n16015 = ~n17152 | ~P3_IR_REG_31__SCAN_IN;
  assign P3_U3151 = ~P3_STATE_REG_SCAN_IN;
  assign n16017 = P1_WR_REG_SCAN_IN ^ ~P2_WR_REG_SCAN_IN;
  assign U28 = P3_WR_REG_SCAN_IN | n16017;
  assign n16018 = P2_RD_REG_SCAN_IN ^ ~P1_RD_REG_SCAN_IN;
  assign U29 = P3_RD_REG_SCAN_IN | n16018;
  assign n16020 = ~n16082 | ~n16175;
  assign n16019 = ~n17037 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n16182 = ~n16020 | ~n16019;
  assign n16023 = ~n17486 | ~P2_DATAO_REG_2__SCAN_IN;
  assign n16022 = ~n16021 | ~P1_DATAO_REG_2__SCAN_IN;
  assign n16184 = ~n16182 | ~n16181;
  assign n16155 = ~n16184 | ~n16023;
  assign n16026 = ~n17503 | ~P2_DATAO_REG_3__SCAN_IN;
  assign n16025 = ~n16024 | ~P1_DATAO_REG_3__SCAN_IN;
  assign n16130 = P1_DATAO_REG_4__SCAN_IN ^ ~P2_DATAO_REG_4__SCAN_IN;
  assign n16028 = ~n16027 | ~P1_DATAO_REG_4__SCAN_IN;
  assign n16145 = ~n16029 | ~n16028;
  assign n16030 = ~n16144;
  assign n16032 = ~n16031 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n16035 = ~n16034 | ~P1_DATAO_REG_6__SCAN_IN;
  assign n16036 = ~n16138;
  assign n16038 = ~n16037 | ~P1_DATAO_REG_7__SCAN_IN;
  assign n16040 = ~n16039 | ~P1_DATAO_REG_8__SCAN_IN;
  assign n16224 = n17565 ^ ~P2_DATAO_REG_9__SCAN_IN;
  assign n16041 = ~n16224;
  assign n16042 = ~n24084 | ~P1_DATAO_REG_9__SCAN_IN;
  assign n16250 = n17578 ^ ~P2_DATAO_REG_10__SCAN_IN;
  assign n16044 = ~n16250;
  assign n16045 = ~n24078 | ~P1_DATAO_REG_10__SCAN_IN;
  assign n16276 = n17589 ^ ~P2_DATAO_REG_11__SCAN_IN;
  assign n16046 = ~n16276;
  assign n16047 = ~n24072 | ~P1_DATAO_REG_11__SCAN_IN;
  assign n16323 = P1_DATAO_REG_12__SCAN_IN ^ ~P2_DATAO_REG_12__SCAN_IN;
  assign n16048 = ~n24066 | ~P1_DATAO_REG_12__SCAN_IN;
  assign n16054 = ~n24053 | ~P1_DATAO_REG_14__SCAN_IN;
  assign n16870 = P1_DATAO_REG_15__SCAN_IN ^ ~P2_DATAO_REG_15__SCAN_IN;
  assign n16055 = ~n16884 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n16890 = P1_DATAO_REG_16__SCAN_IN ^ ~P2_DATAO_REG_16__SCAN_IN;
  assign n16057 = ~n16056 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n16059 = n25297 ^ ~P2_DATAO_REG_17__SCAN_IN;
  assign n18243 = n16951 ^ ~n16059;
  assign n20792 = ~n21363 | ~P3_U3151;
  assign n16070 = n18243 & n17285;
  assign n16324 = n16955 | P3_IR_REG_11__SCAN_IN;
  assign n16060 = ~n16324;
  assign n16522 = ~n16060 | ~n16326;
  assign n16062 = ~n16522;
  assign n16061 = ~P3_IR_REG_13__SCAN_IN;
  assign n16790 = ~n16062 | ~n16061;
  assign n16891 = ~n16063 | ~P3_IR_REG_31__SCAN_IN;
  assign n16064 = ~P3_IR_REG_16__SCAN_IN;
  assign n16893 = ~n16891 | ~n16064;
  assign n16066 = ~n16893 | ~P3_IR_REG_31__SCAN_IN;
  assign n16065 = ~P3_IR_REG_17__SCAN_IN;
  assign n20094 = n16066 ^ ~n16065;
  assign n16068 = n20094 | P3_U3151;
  assign n20796 = ~n13121 | ~P3_U3151;
  assign n20774 = ~n20796;
  assign n16067 = ~n20774 | ~SI_17_;
  assign n16069 = ~n16068 | ~n16067;
  assign P3_U3278 = n16070 | n16069;
  assign n16071 = n23350 ^ ~P3_ADDR_REG_0__SCAN_IN;
  assign SUB_1596_U53 = P2_ADDR_REG_0__SCAN_IN ^ n16071;
  assign n16096 = ~n16071 | ~P2_ADDR_REG_0__SCAN_IN;
  assign n16072 = ~n16074;
  assign n16075 = ~n16073 | ~n16072;
  assign n16098 = ~n16075 | ~n16095;
  assign n16097 = n16098 ^ ~P2_ADDR_REG_1__SCAN_IN;
  assign SUB_1596_U5 = n16097 ^ n16096;
  assign n16077 = ~n13121 | ~SI_0_;
  assign n16079 = ~n16077 | ~n16076;
  assign n17042 = n16079 & n16078;
  assign n16081 = ~n17042 | ~P2_U3088;
  assign n16080 = ~P2_IR_REG_0__SCAN_IN | ~P2_STATE_REG_SCAN_IN;
  assign P2_U3327 = ~n16081 | ~n16080;
  assign n16083 = n16082 ^ ~n16175;
  assign n16085 = ~n16083 | ~n21363;
  assign n16084 = ~n13121 | ~SI_1_;
  assign n17193 = n16085 & n16084;
  assign n16092 = n17193 | P3_STATE_REG_SCAN_IN;
  assign n19964 = ~n19806;
  assign n16086 = ~P3_IR_REG_1__SCAN_IN;
  assign n16087 = ~P3_IR_REG_31__SCAN_IN | ~P3_IR_REG_0__SCAN_IN;
  assign n16088 = ~n16087 | ~P3_IR_REG_1__SCAN_IN;
  assign n16090 = ~n16089 | ~n16088;
  assign n16091 = ~n19840 | ~P3_STATE_REG_SCAN_IN;
  assign P3_U3294 = ~n16092 | ~n16091;
  assign n16100 = n16097 | n16096;
  assign n16099 = ~n16098 | ~P2_ADDR_REG_1__SCAN_IN;
  assign n16102 = ~n16115 | ~n16114;
  assign SUB_1596_U61 = n16102 ^ ~P2_ADDR_REG_2__SCAN_IN;
  assign n16105 = ~n16103 | ~P1_U3086;
  assign n16104 = ~P1_IR_REG_0__SCAN_IN | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3355 = ~n16105 | ~n16104;
  assign n16107 = ~P3_ADDR_REG_3__SCAN_IN;
  assign n16238 = ~n16109 | ~P3_ADDR_REG_3__SCAN_IN;
  assign n16111 = ~P1_ADDR_REG_3__SCAN_IN;
  assign n16112 = ~n13278 | ~P1_ADDR_REG_3__SCAN_IN;
  assign n16244 = ~n16239 | ~n16112;
  assign n16113 = ~P2_ADDR_REG_2__SCAN_IN;
  assign n16116 = ~n16114 | ~n16113;
  assign n16242 = ~P2_ADDR_REG_3__SCAN_IN;
  assign SUB_1596_U60 = n16243 ^ ~n16242;
  assign n18168 = n16118 ^ ~n16117;
  assign n16129 = ~n18168 | ~n17285;
  assign n16119 = ~P3_IR_REG_4__SCAN_IN & ~P3_IR_REG_5__SCAN_IN;
  assign n16124 = ~n16132 | ~n16119;
  assign n16120 = ~n16124 | ~P3_IR_REG_31__SCAN_IN;
  assign n16123 = ~n16120 | ~P3_IR_REG_6__SCAN_IN;
  assign n16121 = ~P3_IR_REG_6__SCAN_IN;
  assign n16122 = ~n16121 | ~P3_IR_REG_31__SCAN_IN;
  assign n16125 = ~n16123 | ~n16122;
  assign n25875 = ~n16125 | ~n16204;
  assign n16127 = ~n25875 & ~P3_U3151;
  assign n16126 = ~n20796 & ~n18169;
  assign n16128 = ~n16127 & ~n16126;
  assign P3_U3289 = ~n16129 | ~n16128;
  assign n17230 = n16131 ^ ~n16130;
  assign n16136 = ~n17230 | ~n17285;
  assign n16147 = n16132 | n16337;
  assign n19972 = n16147 ^ ~P3_IR_REG_4__SCAN_IN;
  assign n16134 = ~n19972 | ~P3_STATE_REG_SCAN_IN;
  assign n16133 = ~n20774 | ~SI_4_;
  assign n16135 = n16134 & n16133;
  assign P3_U3291 = ~n16136 | ~n16135;
  assign n18175 = n16137 ^ ~n16138;
  assign n16143 = ~n18175 | ~n17285;
  assign n25893 = n16139 ^ ~P3_IR_REG_7__SCAN_IN;
  assign n16141 = ~n25893 | ~P3_STATE_REG_SCAN_IN;
  assign n16140 = ~n20774 | ~SI_7_;
  assign n16142 = n16141 & n16140;
  assign P3_U3288 = ~n16143 | ~n16142;
  assign n18165 = n16145 ^ ~n16144;
  assign n16153 = ~n18165 | ~n17285;
  assign n16148 = ~n16147 | ~n16146;
  assign n16149 = ~n16148 | ~P3_IR_REG_31__SCAN_IN;
  assign n25850 = n16149 ^ ~P3_IR_REG_5__SCAN_IN;
  assign n16151 = ~n25850 | ~P3_STATE_REG_SCAN_IN;
  assign n16150 = ~n20774 | ~SI_5_;
  assign n16152 = n16151 & n16150;
  assign P3_U3290 = ~n16153 | ~n16152;
  assign n16156 = n16155 | n16154;
  assign n17218 = ~n16157 | ~n16156;
  assign n16164 = ~n17218 | ~n17285;
  assign n16158 = ~P3_IR_REG_2__SCAN_IN;
  assign n16159 = ~n19806 | ~n16158;
  assign n25811 = n16160 ^ ~P3_IR_REG_3__SCAN_IN;
  assign n16162 = ~n25811 | ~P3_STATE_REG_SCAN_IN;
  assign n16161 = ~n20774 | ~SI_3_;
  assign n16163 = n16162 & n16161;
  assign P3_U3292 = ~n16164 | ~n16163;
  assign n25360 = ~n22164;
  assign n16172 = ~n17038 & ~n25360;
  assign n25337 = ~n21363 | ~P2_U3088;
  assign n16170 = n25337 | n17037;
  assign n16167 = ~n14090 | ~P2_IR_REG_31__SCAN_IN;
  assign n16165 = ~P2_IR_REG_31__SCAN_IN | ~P2_IR_REG_0__SCAN_IN;
  assign n16166 = ~n16165 | ~P2_IR_REG_1__SCAN_IN;
  assign n16168 = ~n16167 | ~n16166;
  assign n16169 = ~n24565 | ~P2_STATE_REG_SCAN_IN;
  assign n16171 = ~n16170 | ~n16169;
  assign P2_U3326 = n16172 | n16171;
  assign n16174 = ~n20774 | ~SI_0_;
  assign n16173 = ~P3_STATE_REG_SCAN_IN | ~P3_IR_REG_0__SCAN_IN;
  assign n16180 = ~n16174 | ~n16173;
  assign n16178 = ~n16175;
  assign n16177 = ~n16176 | ~P1_DATAO_REG_0__SCAN_IN;
  assign n17197 = n16178 & n16177;
  assign n16179 = ~n20792 & ~n17197;
  assign P3_U3295 = n16180 | n16179;
  assign n16183 = n16182 | n16181;
  assign n17206 = n16184 & n16183;
  assign n16188 = ~n17206 & ~n20792;
  assign n16186 = ~n19967 | ~P3_STATE_REG_SCAN_IN;
  assign n16185 = ~n20774 | ~SI_2_;
  assign n16187 = ~n16186 | ~n16185;
  assign P3_U3293 = n16188 | n16187;
  assign n16189 = ~n17520;
  assign n16201 = ~n16189 | ~n22164;
  assign n17492 = n17487 | P2_IR_REG_2__SCAN_IN;
  assign n16190 = ~n17492;
  assign n16215 = ~P2_IR_REG_3__SCAN_IN;
  assign n17510 = ~n16190 | ~n16215;
  assign n16191 = ~n17510;
  assign n17512 = ~P2_IR_REG_4__SCAN_IN;
  assign n17515 = ~n16191 | ~n17512;
  assign n16192 = ~n17515 | ~P2_IR_REG_31__SCAN_IN;
  assign n16195 = ~n16192 | ~P2_IR_REG_5__SCAN_IN;
  assign n16193 = ~P2_IR_REG_5__SCAN_IN;
  assign n16194 = ~n16193 | ~P2_IR_REG_31__SCAN_IN;
  assign n16197 = ~n16195 | ~n16194;
  assign n16196 = ~n17597;
  assign n24647 = n16197 & n16196;
  assign n24631 = ~n24647;
  assign n16199 = ~n24631 & ~P2_U3088;
  assign n16198 = ~n25337 & ~n17521;
  assign n16200 = ~n16199 & ~n16198;
  assign P2_U3322 = ~n16201 | ~n16200;
  assign n18182 = n16202 ^ ~n16203;
  assign n16212 = n18182 | n20792;
  assign n16251 = ~P3_IR_REG_7__SCAN_IN;
  assign n16205 = ~n16254 | ~n16251;
  assign n16207 = ~n16205 | ~P3_IR_REG_31__SCAN_IN;
  assign n16206 = ~P3_IR_REG_8__SCAN_IN;
  assign n16208 = n16207 | n16206;
  assign n16225 = ~n16207 | ~n16206;
  assign n25916 = ~n16208 | ~n16225;
  assign n16210 = ~n25916 & ~P3_U3151;
  assign n18183 = ~SI_8_;
  assign n16209 = ~n20796 & ~n18183;
  assign n16211 = ~n16210 & ~n16209;
  assign P3_U3287 = ~n16212 | ~n16211;
  assign n16213 = ~n17948;
  assign n16222 = ~n16213 | ~n22164;
  assign n16214 = ~n17492 | ~P2_IR_REG_31__SCAN_IN;
  assign n16217 = ~n16214 | ~P2_IR_REG_3__SCAN_IN;
  assign n16216 = ~n16215 | ~P2_IR_REG_31__SCAN_IN;
  assign n16218 = ~n16217 | ~n16216;
  assign n24606 = n16218 & n17510;
  assign n24576 = ~n24606;
  assign n16220 = ~n24576 & ~P2_U3088;
  assign n16219 = ~n25337 & ~n17503;
  assign n16221 = ~n16220 & ~n16219;
  assign P2_U3324 = ~n16222 | ~n16221;
  assign n18190 = n16223 ^ ~n16224;
  assign n16230 = ~n18190 | ~n17285;
  assign n16226 = ~n16225 | ~P3_IR_REG_31__SCAN_IN;
  assign n19984 = n16226 ^ ~P3_IR_REG_9__SCAN_IN;
  assign n16228 = ~n19984 | ~P3_STATE_REG_SCAN_IN;
  assign n16227 = ~n20774 | ~SI_9_;
  assign n16229 = n16228 & n16227;
  assign P3_U3286 = ~n16230 | ~n16229;
  assign n16231 = ~n17038;
  assign n16237 = ~n16231 | ~n23156;
  assign n24085 = ~n13122 | ~P1_U3086;
  assign n16233 = ~P2_DATAO_REG_1__SCAN_IN;
  assign n16235 = ~n24085 & ~n16233;
  assign n16234 = ~n16823 & ~P1_U3086;
  assign n16236 = ~n16235 & ~n16234;
  assign P1_U3354 = ~n16237 | ~n16236;
  assign n16318 = ~P2_ADDR_REG_4__SCAN_IN;
  assign n16248 = n16320 ^ ~n16318;
  assign n16246 = ~n16244;
  assign n16247 = ~n16246 | ~n16245;
  assign SUB_1596_U59 = n13409 ^ ~n16248;
  assign n18196 = n16249 ^ ~n16250;
  assign n16260 = ~n18196 | ~n17285;
  assign n16252 = ~P3_IR_REG_9__SCAN_IN & ~P3_IR_REG_8__SCAN_IN;
  assign n16253 = n16252 & n16251;
  assign n16255 = ~n16254 | ~n16253;
  assign n16256 = ~n16255 | ~P3_IR_REG_31__SCAN_IN;
  assign n19987 = n16256 ^ ~P3_IR_REG_10__SCAN_IN;
  assign n16258 = ~n19987 | ~P3_STATE_REG_SCAN_IN;
  assign n16257 = ~n20774 | ~SI_10_;
  assign n16259 = n16258 & n16257;
  assign P3_U3285 = ~n16260 | ~n16259;
  assign n16264 = ~n17520 & ~n24106;
  assign n16262 = n23444 | P1_U3086;
  assign n24110 = ~n24085;
  assign n16261 = ~n24110 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n16263 = ~n16262 | ~n16261;
  assign P1_U3350 = n16264 | n16263;
  assign n26311 = ~n17461;
  assign n17133 = ~n17134;
  assign n16290 = ~n26311 & ~n17133;
  assign n16265 = ~P3_D_REG_7__SCAN_IN;
  assign P3_U3258 = ~n26312 & ~n16265;
  assign n17106 = ~P3_D_REG_8__SCAN_IN;
  assign P3_U3257 = ~n26312 & ~n17106;
  assign n16266 = ~P3_D_REG_2__SCAN_IN;
  assign P3_U3263 = ~n16290 & ~n16266;
  assign n16267 = ~P3_D_REG_4__SCAN_IN;
  assign P3_U3261 = ~n16290 & ~n16267;
  assign n16268 = ~P3_D_REG_5__SCAN_IN;
  assign P3_U3260 = ~n16290 & ~n16268;
  assign n16269 = ~P3_D_REG_3__SCAN_IN;
  assign P3_U3262 = ~n16290 & ~n16269;
  assign n16270 = ~P3_D_REG_6__SCAN_IN;
  assign P3_U3259 = ~n16290 & ~n16270;
  assign n16274 = ~n25342 & ~n24106;
  assign n16272 = n23486 | P1_U3086;
  assign n16271 = ~n24110 | ~P2_DATAO_REG_7__SCAN_IN;
  assign n16273 = ~n16272 | ~n16271;
  assign P1_U3348 = n16274 | n16273;
  assign n16285 = ~n18203 | ~n17285;
  assign n16277 = ~n16955 | ~P3_IR_REG_31__SCAN_IN;
  assign n16280 = ~n16277 | ~P3_IR_REG_11__SCAN_IN;
  assign n16278 = ~P3_IR_REG_11__SCAN_IN;
  assign n16279 = ~n16278 | ~P3_IR_REG_31__SCAN_IN;
  assign n16281 = ~n16280 | ~n16279;
  assign n19989 = n16281 & n16324;
  assign n16283 = ~n19989 | ~P3_STATE_REG_SCAN_IN;
  assign n16282 = ~n20774 | ~SI_11_;
  assign n16284 = n16283 & n16282;
  assign P3_U3284 = ~n16285 | ~n16284;
  assign n16289 = ~n26312 & ~P3_D_REG_0__SCAN_IN;
  assign n20786 = ~n16286;
  assign n17135 = ~n20786 | ~n16287;
  assign n16288 = ~n26311 & ~n17135;
  assign P3_U3376 = ~n16289 & ~n16288;
  assign n26312 = n16290;
  assign n16291 = ~P3_D_REG_23__SCAN_IN;
  assign P3_U3242 = ~n26312 & ~n16291;
  assign n16292 = ~P3_D_REG_28__SCAN_IN;
  assign P3_U3237 = ~n26312 & ~n16292;
  assign n16293 = ~P3_D_REG_13__SCAN_IN;
  assign P3_U3252 = ~n26312 & ~n16293;
  assign n16294 = ~P3_D_REG_30__SCAN_IN;
  assign P3_U3235 = ~n26312 & ~n16294;
  assign n16295 = ~P3_D_REG_15__SCAN_IN;
  assign P3_U3250 = ~n26312 & ~n16295;
  assign n16296 = ~P3_D_REG_16__SCAN_IN;
  assign P3_U3249 = ~n26312 & ~n16296;
  assign n17105 = ~P3_D_REG_9__SCAN_IN;
  assign P3_U3256 = ~n26312 & ~n17105;
  assign n16297 = ~P3_D_REG_26__SCAN_IN;
  assign P3_U3239 = ~n26312 & ~n16297;
  assign n16298 = ~P3_D_REG_11__SCAN_IN;
  assign P3_U3254 = ~n26312 & ~n16298;
  assign n16299 = ~P3_D_REG_12__SCAN_IN;
  assign P3_U3253 = ~n26312 & ~n16299;
  assign n16300 = ~P3_D_REG_21__SCAN_IN;
  assign P3_U3244 = ~n26312 & ~n16300;
  assign n16301 = ~P3_D_REG_14__SCAN_IN;
  assign P3_U3251 = ~n26312 & ~n16301;
  assign n16302 = ~P3_D_REG_31__SCAN_IN;
  assign P3_U3234 = ~n26312 & ~n16302;
  assign n16303 = ~P3_D_REG_10__SCAN_IN;
  assign P3_U3255 = ~n26312 & ~n16303;
  assign n16304 = ~P3_D_REG_29__SCAN_IN;
  assign P3_U3236 = ~n26312 & ~n16304;
  assign n16305 = ~P3_D_REG_24__SCAN_IN;
  assign P3_U3241 = ~n26312 & ~n16305;
  assign n16306 = ~P3_D_REG_27__SCAN_IN;
  assign P3_U3238 = ~n26312 & ~n16306;
  assign n16307 = ~P3_D_REG_18__SCAN_IN;
  assign P3_U3247 = ~n26312 & ~n16307;
  assign n16308 = ~P3_D_REG_19__SCAN_IN;
  assign P3_U3246 = ~n26312 & ~n16308;
  assign n16309 = ~P3_D_REG_20__SCAN_IN;
  assign P3_U3245 = ~n26312 & ~n16309;
  assign n16310 = ~P3_D_REG_25__SCAN_IN;
  assign P3_U3240 = ~n26312 & ~n16310;
  assign n16311 = ~P3_D_REG_22__SCAN_IN;
  assign P3_U3243 = ~n26312 & ~n16311;
  assign n16312 = ~P3_D_REG_17__SCAN_IN;
  assign P3_U3248 = ~n26312 & ~n16312;
  assign n16315 = ~P1_ADDR_REG_5__SCAN_IN;
  assign n16317 = ~n16316 | ~P1_ADDR_REG_5__SCAN_IN;
  assign n16319 = ~n16320 | ~n16318;
  assign n16321 = ~n16320;
  assign SUB_1596_U58 = n16539 ^ ~P2_ADDR_REG_5__SCAN_IN;
  assign n16334 = ~n18208 & ~n20792;
  assign n16325 = ~n16324 | ~P3_IR_REG_31__SCAN_IN;
  assign n16328 = ~n16325 | ~P3_IR_REG_12__SCAN_IN;
  assign n16327 = ~n16326 | ~P3_IR_REG_31__SCAN_IN;
  assign n16329 = ~n16328 | ~n16327;
  assign n25988 = ~n16329 | ~n16522;
  assign n16330 = ~n25988;
  assign n16332 = ~n16330 | ~P3_STATE_REG_SCAN_IN;
  assign n16331 = ~n20774 | ~SI_12_;
  assign n16333 = ~n16332 | ~n16331;
  assign P3_U3283 = n16334 | n16333;
  assign n16336 = ~P3_IR_REG_26__SCAN_IN & ~P3_IR_REG_27__SCAN_IN;
  assign n16335 = ~P3_IR_REG_25__SCAN_IN & ~P3_IR_REG_24__SCAN_IN;
  assign n16422 = n16460;
  assign n16342 = ~n16422 | ~P3_REG2_REG_11__SCAN_IN;
  assign n20766 = ~n16345;
  assign n16341 = ~n18380 | ~P3_REG0_REG_11__SCAN_IN;
  assign n16349 = ~n16342 | ~n16341;
  assign n16344 = n13177 & P3_REG3_REG_11__SCAN_IN;
  assign n25699 = n16344 | n16374;
  assign n16347 = ~n16484 | ~n25699;
  assign n16463 = n20759 & n16345;
  assign n18368 = n16463;
  assign n16346 = ~n18368 | ~P3_REG1_REG_11__SCAN_IN;
  assign n16348 = ~n16347 | ~n16346;
  assign n16351 = ~n26059 | ~P3_U3897;
  assign n16350 = ~n26454 | ~P3_DATAO_REG_11__SCAN_IN;
  assign P3_U3502 = ~n16351 | ~n16350;
  assign n16353 = ~n16422 | ~P3_REG2_REG_6__SCAN_IN;
  assign n16352 = ~n18368 | ~P3_REG1_REG_6__SCAN_IN;
  assign n16358 = ~n16353 | ~n16352;
  assign n16354 = ~n16386 | ~P3_REG3_REG_6__SCAN_IN;
  assign n26151 = ~n16425 | ~n16354;
  assign n16356 = ~n16484 | ~n26151;
  assign n16355 = ~n18380 | ~P3_REG0_REG_6__SCAN_IN;
  assign n16357 = ~n16356 | ~n16355;
  assign n16360 = ~n26189 | ~P3_U3897;
  assign n16359 = ~n26454 | ~P3_DATAO_REG_6__SCAN_IN;
  assign P3_U3497 = ~n16360 | ~n16359;
  assign n16362 = ~n16422 | ~P3_REG2_REG_13__SCAN_IN;
  assign n16361 = ~n18380 | ~P3_REG0_REG_13__SCAN_IN;
  assign n16368 = ~n16362 | ~n16361;
  assign n16364 = n16376 | n16363;
  assign n20485 = ~n16414 | ~n16364;
  assign n16366 = ~n16484 | ~n20485;
  assign n16365 = ~n18368 | ~P3_REG1_REG_13__SCAN_IN;
  assign n16367 = ~n16366 | ~n16365;
  assign n16370 = ~n19552 | ~P3_U3897;
  assign n16369 = ~n26454 | ~P3_DATAO_REG_13__SCAN_IN;
  assign P3_U3504 = ~n16370 | ~n16369;
  assign n16372 = ~n16422 | ~P3_REG2_REG_12__SCAN_IN;
  assign n16371 = ~n16463 | ~P3_REG1_REG_12__SCAN_IN;
  assign n16380 = ~n16372 | ~n16371;
  assign n16375 = ~n16374 & ~n16373;
  assign n20508 = n16376 | n16375;
  assign n16378 = ~n16484 | ~n20508;
  assign n16377 = ~n18380 | ~P3_REG0_REG_12__SCAN_IN;
  assign n16379 = ~n16378 | ~n16377;
  assign n16382 = ~n25692 | ~P3_U3897;
  assign n16381 = ~n26454 | ~P3_DATAO_REG_12__SCAN_IN;
  assign P3_U3503 = ~n16382 | ~n16381;
  assign n16384 = ~n16422 | ~P3_REG2_REG_5__SCAN_IN;
  assign n16383 = ~n16463 | ~P3_REG1_REG_5__SCAN_IN;
  assign n16390 = ~n16384 | ~n16383;
  assign n16385 = n16452 | n25667;
  assign n26175 = ~n16386 | ~n16385;
  assign n16388 = ~n16484 | ~n26175;
  assign n16387 = ~n18380 | ~P3_REG0_REG_5__SCAN_IN;
  assign n16389 = ~n16388 | ~n16387;
  assign n16392 = ~n26205 | ~P3_U3897;
  assign n16391 = ~n26454 | ~P3_DATAO_REG_5__SCAN_IN;
  assign P3_U3496 = ~n16392 | ~n16391;
  assign n16394 = ~n16422 | ~P3_REG2_REG_10__SCAN_IN;
  assign n16393 = ~n18380 | ~P3_REG0_REG_10__SCAN_IN;
  assign n16399 = ~n16394 | ~n16393;
  assign n16395 = ~n16403 | ~P3_REG3_REG_10__SCAN_IN;
  assign n26067 = ~n13177 | ~n16395;
  assign n16397 = ~n16484 | ~n26067;
  assign n16396 = ~n18368 | ~P3_REG1_REG_10__SCAN_IN;
  assign n16398 = ~n16397 | ~n16396;
  assign n16401 = ~n26085 | ~P3_U3897;
  assign n16400 = ~n26454 | ~P3_DATAO_REG_10__SCAN_IN;
  assign P3_U3501 = ~n16401 | ~n16400;
  assign n16405 = ~n16422 | ~P3_REG2_REG_9__SCAN_IN;
  assign n16402 = n16473 | n19708;
  assign n26094 = ~n16403 | ~n16402;
  assign n16404 = ~n16484 | ~n26094;
  assign n16409 = ~n16405 | ~n16404;
  assign n16407 = ~n16463 | ~P3_REG1_REG_9__SCAN_IN;
  assign n16406 = ~n18380 | ~P3_REG0_REG_9__SCAN_IN;
  assign n16408 = ~n16407 | ~n16406;
  assign n16411 = ~n26116 | ~P3_U3897;
  assign n16410 = ~n26454 | ~P3_DATAO_REG_9__SCAN_IN;
  assign P3_U3500 = ~n16411 | ~n16410;
  assign n16413 = ~n16422 | ~P3_REG2_REG_14__SCAN_IN;
  assign n16412 = ~n18368 | ~P3_REG1_REG_14__SCAN_IN;
  assign n16419 = ~n16413 | ~n16412;
  assign n16415 = ~n16414 | ~P3_REG3_REG_14__SCAN_IN;
  assign n20463 = ~n16491 | ~n16415;
  assign n16417 = ~n20463 | ~n16484;
  assign n16416 = ~n18380 | ~P3_REG0_REG_14__SCAN_IN;
  assign n16418 = ~n16417 | ~n16416;
  assign n16421 = ~n19406 | ~P3_U3897;
  assign n16420 = ~n26454 | ~P3_DATAO_REG_14__SCAN_IN;
  assign P3_U3505 = ~n16421 | ~n16420;
  assign n16424 = ~n16422 | ~P3_REG2_REG_7__SCAN_IN;
  assign n18380 = n18340;
  assign n16423 = ~n18380 | ~P3_REG0_REG_7__SCAN_IN;
  assign n16430 = ~n16424 | ~n16423;
  assign n16426 = n16425 & P3_REG3_REG_7__SCAN_IN;
  assign n26141 = n16426 | n16471;
  assign n16428 = ~n16484 | ~n26141;
  assign n16427 = ~n16463 | ~P3_REG1_REG_7__SCAN_IN;
  assign n16429 = ~n16428 | ~n16427;
  assign n19134 = ~n16430 & ~n16429;
  assign n26165 = ~n19134;
  assign n16432 = ~n26165 | ~P3_U3897;
  assign n16431 = ~n26454 | ~P3_DATAO_REG_7__SCAN_IN;
  assign P3_U3498 = ~n16432 | ~n16431;
  assign n16434 = ~n16460 | ~P3_REG2_REG_0__SCAN_IN;
  assign n16433 = ~n16484 | ~P3_REG3_REG_0__SCAN_IN;
  assign n16438 = ~n16434 | ~n16433;
  assign n16436 = ~n16463 | ~P3_REG1_REG_0__SCAN_IN;
  assign n16435 = ~n18340 | ~P3_REG0_REG_0__SCAN_IN;
  assign n16437 = ~n16436 | ~n16435;
  assign n16440 = ~n26287 | ~P3_U3897;
  assign n16439 = ~n26454 | ~P3_DATAO_REG_0__SCAN_IN;
  assign P3_U3491 = ~n16440 | ~n16439;
  assign n16442 = ~n16463 | ~P3_REG1_REG_3__SCAN_IN;
  assign n16441 = ~n18340 | ~P3_REG0_REG_3__SCAN_IN;
  assign n16447 = ~n16442 | ~n16441;
  assign n16445 = ~n16460 | ~P3_REG2_REG_3__SCAN_IN;
  assign n16443 = ~P3_REG3_REG_3__SCAN_IN;
  assign n16444 = ~n16484 | ~n16443;
  assign n16446 = ~n16445 | ~n16444;
  assign n16449 = ~n26252 | ~P3_U3897;
  assign n16448 = ~n26454 | ~P3_DATAO_REG_3__SCAN_IN;
  assign P3_U3494 = ~n16449 | ~n16448;
  assign n16451 = ~n16422 | ~P3_REG2_REG_4__SCAN_IN;
  assign n16450 = ~n18380 | ~P3_REG0_REG_4__SCAN_IN;
  assign n16457 = ~n16451 | ~n16450;
  assign n16453 = P3_REG3_REG_4__SCAN_IN & P3_REG3_REG_3__SCAN_IN;
  assign n26213 = n16453 | n16452;
  assign n16455 = ~n16484 | ~n26213;
  assign n16454 = ~n16463 | ~P3_REG1_REG_4__SCAN_IN;
  assign n16456 = ~n16455 | ~n16454;
  assign n16459 = ~n26229 | ~P3_U3897;
  assign n16458 = ~n26454 | ~P3_DATAO_REG_4__SCAN_IN;
  assign P3_U3495 = ~n16459 | ~n16458;
  assign n16462 = ~n16460 | ~P3_REG2_REG_1__SCAN_IN;
  assign n16461 = ~n16484 | ~P3_REG3_REG_1__SCAN_IN;
  assign n16465 = ~n18340 | ~P3_REG0_REG_1__SCAN_IN;
  assign n16464 = ~n16463 | ~P3_REG1_REG_1__SCAN_IN;
  assign n16466 = ~n16465 | ~n16464;
  assign n16468 = ~n26454 | ~P3_DATAO_REG_1__SCAN_IN;
  assign P3_U3492 = ~n16469 | ~n16468;
  assign n16475 = ~n16422 | ~P3_REG2_REG_8__SCAN_IN;
  assign n16472 = ~n16471 & ~n16470;
  assign n26101 = n16473 | n16472;
  assign n16474 = ~n16484 | ~n26101;
  assign n16479 = ~n16475 | ~n16474;
  assign n16477 = ~n18368 | ~P3_REG1_REG_8__SCAN_IN;
  assign n16476 = ~n18380 | ~P3_REG0_REG_8__SCAN_IN;
  assign n16478 = ~n16477 | ~n16476;
  assign n16481 = ~n26086 | ~P3_U3897;
  assign n16480 = ~n26454 | ~P3_DATAO_REG_8__SCAN_IN;
  assign P3_U3499 = ~n16481 | ~n16480;
  assign n16482 = ~n16463 | ~P3_REG1_REG_2__SCAN_IN;
  assign n16488 = ~n16483 | ~n16482;
  assign n16486 = ~n16484 | ~P3_REG3_REG_2__SCAN_IN;
  assign n16485 = ~n18340 | ~P3_REG0_REG_2__SCAN_IN;
  assign n16487 = ~n16486 | ~n16485;
  assign n16490 = ~n26286 | ~P3_U3897;
  assign n16489 = ~n26454 | ~P3_DATAO_REG_2__SCAN_IN;
  assign P3_U3493 = ~n16490 | ~n16489;
  assign n16492 = ~n16491 | ~P3_REG3_REG_15__SCAN_IN;
  assign n20444 = ~n16501 | ~n16492;
  assign n16494 = ~n20444 | ~n16484;
  assign n16493 = ~n16422 | ~P3_REG2_REG_15__SCAN_IN;
  assign n16498 = n16494 & n16493;
  assign n16496 = ~n18368 | ~P3_REG1_REG_15__SCAN_IN;
  assign n16495 = ~n18380 | ~P3_REG0_REG_15__SCAN_IN;
  assign n16497 = n16496 & n16495;
  assign n19646 = ~n16498 | ~n16497;
  assign n16500 = ~n19646 | ~P3_U3897;
  assign n16499 = ~n26454 | ~P3_DATAO_REG_15__SCAN_IN;
  assign P3_U3506 = ~n16500 | ~n16499;
  assign n16502 = n16501 & P3_REG3_REG_16__SCAN_IN;
  assign n20425 = n16502 | n16529;
  assign n16508 = ~n20425 | ~n16484;
  assign n16504 = ~n16422 | ~P3_REG2_REG_16__SCAN_IN;
  assign n16503 = ~n16463 | ~P3_REG1_REG_16__SCAN_IN;
  assign n16506 = ~n16504 | ~n16503;
  assign n16505 = n18380 & P3_REG0_REG_16__SCAN_IN;
  assign n16507 = ~n16506 & ~n16505;
  assign n19795 = ~n16508 | ~n16507;
  assign n16510 = ~n19795 | ~P3_U3897;
  assign n16509 = ~n26454 | ~P3_DATAO_REG_16__SCAN_IN;
  assign P3_U3507 = ~n16510 | ~n16509;
  assign n16512 = ~n16511;
  assign n16514 = ~P1_U4016 | ~n17382;
  assign n16513 = ~n24319 | ~P1_DATAO_REG_1__SCAN_IN;
  assign P1_U3561 = ~n16514 | ~n16513;
  assign n16516 = ~P1_U4016 | ~n23034;
  assign n16515 = ~n24319 | ~P1_DATAO_REG_12__SCAN_IN;
  assign P1_U3572 = ~n16516 | ~n16515;
  assign n16518 = ~P1_U4016 | ~n23854;
  assign n16517 = ~n24319 | ~P1_DATAO_REG_5__SCAN_IN;
  assign P1_U3565 = ~n16518 | ~n16517;
  assign n16521 = ~n16520 | ~P1_DATAO_REG_13__SCAN_IN;
  assign n18212 = ~n16519 | ~n16521;
  assign n16527 = ~n18212 | ~n17285;
  assign n16523 = ~n16522 | ~P3_IR_REG_31__SCAN_IN;
  assign n19993 = n16523 ^ ~P3_IR_REG_13__SCAN_IN;
  assign n16525 = ~n19993 | ~P3_STATE_REG_SCAN_IN;
  assign n16524 = ~n20774 | ~SI_13_;
  assign n16526 = n16525 & n16524;
  assign P3_U3282 = ~n16527 | ~n16526;
  assign n16528 = ~P3_REG3_REG_17__SCAN_IN;
  assign n16530 = ~n16529 & ~n16528;
  assign n20407 = n16798 | n16530;
  assign n16536 = ~n20407 | ~n16484;
  assign n16532 = ~n16422 | ~P3_REG2_REG_17__SCAN_IN;
  assign n16531 = ~n18368 | ~P3_REG1_REG_17__SCAN_IN;
  assign n16534 = ~n16532 | ~n16531;
  assign n16533 = n18380 & P3_REG0_REG_17__SCAN_IN;
  assign n16535 = ~n16534 & ~n16533;
  assign n19771 = ~n16536 | ~n16535;
  assign n16538 = ~n19771 | ~P3_U3897;
  assign n16537 = ~n26454 | ~P3_DATAO_REG_17__SCAN_IN;
  assign P3_U3508 = ~n16538 | ~n16537;
  assign n16541 = ~n16540;
  assign n16542 = ~n13181 | ~n16541;
  assign n16545 = ~P3_ADDR_REG_6__SCAN_IN;
  assign n16547 = ~P1_ADDR_REG_6__SCAN_IN;
  assign n16549 = ~n16835 | ~n16834;
  assign SUB_1596_U57 = n16549 ^ ~P2_ADDR_REG_6__SCAN_IN;
  assign n16551 = ~P1_U4016 | ~n23017;
  assign n16550 = ~n24319 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P1_U3573 = ~n16551 | ~n16550;
  assign n16553 = ~P1_U4016 | ~n23035;
  assign n16552 = ~n24319 | ~P1_DATAO_REG_14__SCAN_IN;
  assign P1_U3574 = ~n16553 | ~n16552;
  assign n16555 = ~P1_U4016 | ~n23753;
  assign n16554 = ~n24319 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P1_U3571 = ~n16555 | ~n16554;
  assign P1_U4016 = ~n24319;
  assign n16557 = ~P1_U4016 | ~n23825;
  assign n16556 = ~n24319 | ~P1_DATAO_REG_8__SCAN_IN;
  assign P1_U3568 = ~n16557 | ~n16556;
  assign n16559 = ~P1_U4016 | ~n23769;
  assign n16558 = ~n24319 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P1_U3570 = ~n16559 | ~n16558;
  assign n16561 = ~P1_U4016 | ~n17357;
  assign n16560 = ~n24319 | ~P1_DATAO_REG_3__SCAN_IN;
  assign P1_U3563 = ~n16561 | ~n16560;
  assign n16563 = ~n22982 | ~P1_U4016;
  assign n16562 = ~n24319 | ~P1_DATAO_REG_17__SCAN_IN;
  assign P1_U3577 = ~n16563 | ~n16562;
  assign n16567 = ~n16564;
  assign n16566 = ~n16565;
  assign n16571 = ~n16568;
  assign n16570 = ~P2_IR_REG_23__SCAN_IN & ~P2_IR_REG_26__SCAN_IN;
  assign n16576 = ~n16571 | ~n14864;
  assign n16573 = ~P2_IR_REG_15__SCAN_IN & ~P2_IR_REG_20__SCAN_IN;
  assign n16577 = ~P2_IR_REG_28__SCAN_IN;
  assign n16579 = ~n16578 | ~P2_IR_REG_31__SCAN_IN;
  assign n16582 = ~n16579 | ~P2_IR_REG_29__SCAN_IN;
  assign n16581 = ~n16580 | ~P2_IR_REG_31__SCAN_IN;
  assign n16584 = ~n16582 | ~n16581;
  assign n16586 = ~n16780 | ~P2_REG1_REG_8__SCAN_IN;
  assign n16781 = n22133 & n22139;
  assign n16585 = ~n16781 | ~P2_REG0_REG_8__SCAN_IN;
  assign n16595 = ~n16586 | ~n16585;
  assign n16593 = ~n21356 | ~P2_REG2_REG_8__SCAN_IN;
  assign n16742 = ~P2_REG3_REG_4__SCAN_IN | ~P2_REG3_REG_3__SCAN_IN;
  assign n16714 = ~n16725 | ~n16590;
  assign n16622 = ~P2_REG3_REG_8__SCAN_IN;
  assign n25033 = n16714 ^ ~n16622;
  assign n16591 = ~n25033;
  assign n16592 = ~n17780 | ~n16591;
  assign n16594 = ~n16593 | ~n16592;
  assign n16597 = ~P2_U3947 | ~n25049;
  assign n16596 = ~n25592 | ~P2_DATAO_REG_8__SCAN_IN;
  assign P2_U3539 = ~n16597 | ~n16596;
  assign n16599 = ~n21359 | ~P2_REG0_REG_18__SCAN_IN;
  assign n16598 = ~n21356 | ~P2_REG2_REG_18__SCAN_IN;
  assign n16601 = ~n16599 | ~n16598;
  assign n16600 = n16780 & P2_REG1_REG_18__SCAN_IN;
  assign n16608 = ~n16601 & ~n16600;
  assign n16602 = ~P2_REG3_REG_8__SCAN_IN | ~P2_REG3_REG_9__SCAN_IN;
  assign n16701 = ~n16676 | ~P2_REG3_REG_12__SCAN_IN;
  assign n16604 = ~P2_REG3_REG_13__SCAN_IN;
  assign n16605 = ~P2_REG3_REG_14__SCAN_IN | ~P2_REG3_REG_15__SCAN_IN;
  assign n16606 = P2_REG3_REG_17__SCAN_IN & P2_REG3_REG_16__SCAN_IN;
  assign n21723 = n17671 ^ ~P2_REG3_REG_18__SCAN_IN;
  assign n16607 = n21723 | n16777;
  assign n21734 = ~n16608 | ~n16607;
  assign n16610 = ~P2_U3947 | ~n21734;
  assign n16609 = ~n25592 | ~P2_DATAO_REG_18__SCAN_IN;
  assign P2_U3549 = ~n16610 | ~n16609;
  assign n16612 = ~n16780 | ~P2_REG1_REG_2__SCAN_IN;
  assign n16611 = ~n16781 | ~P2_REG0_REG_2__SCAN_IN;
  assign n16613 = ~P2_REG3_REG_2__SCAN_IN;
  assign n16614 = n16777 | n16613;
  assign n16616 = ~n16615 | ~n16614;
  assign n16619 = ~P2_U3947 | ~n25252;
  assign n16618 = ~n25592 | ~P2_DATAO_REG_2__SCAN_IN;
  assign P2_U3533 = ~n16619 | ~n16618;
  assign n16621 = ~n16780 | ~P2_REG1_REG_9__SCAN_IN;
  assign n16620 = ~n16781 | ~P2_REG0_REG_9__SCAN_IN;
  assign n16630 = ~n16621 | ~n16620;
  assign n16628 = ~n21356 | ~P2_REG2_REG_9__SCAN_IN;
  assign n17780 = ~n16777;
  assign n16624 = n16714 | n16622;
  assign n16623 = ~P2_REG3_REG_9__SCAN_IN;
  assign n16625 = ~n16624 | ~n16623;
  assign n25009 = ~n16625 | ~n16686;
  assign n16626 = ~n25009;
  assign n16627 = ~n17780 | ~n16626;
  assign n16629 = ~n16628 | ~n16627;
  assign n16632 = ~P2_U3947 | ~n25021;
  assign n16631 = ~n25592 | ~P2_DATAO_REG_9__SCAN_IN;
  assign P2_U3540 = ~n16632 | ~n16631;
  assign n16634 = ~n16780 | ~P2_REG1_REG_14__SCAN_IN;
  assign n16633 = ~n16781 | ~P2_REG0_REG_14__SCAN_IN;
  assign n16638 = ~n16634 | ~n16633;
  assign n21831 = n16661 ^ ~P2_REG3_REG_14__SCAN_IN;
  assign n16636 = ~n17780 | ~n21831;
  assign n16635 = ~n21356 | ~P2_REG2_REG_14__SCAN_IN;
  assign n16637 = ~n16636 | ~n16635;
  assign n16640 = ~P2_U3947 | ~n21413;
  assign n16639 = ~n25592 | ~P2_DATAO_REG_14__SCAN_IN;
  assign P2_U3545 = ~n16640 | ~n16639;
  assign n16644 = ~n17671;
  assign n16642 = ~n16751 | ~P2_REG3_REG_16__SCAN_IN;
  assign n16641 = ~P2_REG3_REG_17__SCAN_IN;
  assign n16643 = ~n16642 | ~n16641;
  assign n21745 = n16644 & n16643;
  assign n16646 = ~n21745 | ~n17780;
  assign n16645 = ~n21356 | ~P2_REG2_REG_17__SCAN_IN;
  assign n16650 = ~n16646 | ~n16645;
  assign n16648 = ~n16780 | ~P2_REG1_REG_17__SCAN_IN;
  assign n16647 = ~n21359 | ~P2_REG0_REG_17__SCAN_IN;
  assign n16649 = ~n16648 | ~n16647;
  assign n16652 = ~P2_U3947 | ~n21436;
  assign n16651 = ~n25592 | ~P2_DATAO_REG_17__SCAN_IN;
  assign P2_U3548 = ~n16652 | ~n16651;
  assign n16654 = ~n21356 | ~P2_REG2_REG_12__SCAN_IN;
  assign n16653 = ~n21359 | ~P2_REG0_REG_12__SCAN_IN;
  assign n16658 = ~n16654 | ~n16653;
  assign n24390 = ~P2_REG3_REG_12__SCAN_IN;
  assign n24395 = n16676 ^ ~n24390;
  assign n16656 = ~n17780 | ~n24395;
  assign n16655 = ~n16780 | ~P2_REG1_REG_12__SCAN_IN;
  assign n16657 = ~n16656 | ~n16655;
  assign n16660 = ~P2_U3947 | ~n24955;
  assign n16659 = ~n25592 | ~P2_DATAO_REG_12__SCAN_IN;
  assign P2_U3543 = ~n16660 | ~n16659;
  assign n20824 = ~P2_REG3_REG_14__SCAN_IN;
  assign n16663 = ~n16661 & ~n20824;
  assign n16662 = ~P2_REG3_REG_15__SCAN_IN;
  assign n21805 = n16663 ^ ~n16662;
  assign n16665 = ~n17780 | ~n21805;
  assign n16664 = ~n21356 | ~P2_REG2_REG_15__SCAN_IN;
  assign n16669 = ~n16665 | ~n16664;
  assign n16667 = ~n16780 | ~P2_REG1_REG_15__SCAN_IN;
  assign n16666 = ~n16781 | ~P2_REG0_REG_15__SCAN_IN;
  assign n16668 = ~n16667 | ~n16666;
  assign n16671 = ~P2_U3947 | ~n21818;
  assign n16670 = ~n25592 | ~P2_DATAO_REG_15__SCAN_IN;
  assign P2_U3546 = ~n16671 | ~n16670;
  assign n16673 = ~n16780 | ~P2_REG1_REG_11__SCAN_IN;
  assign n16672 = ~n21359 | ~P2_REG0_REG_11__SCAN_IN;
  assign n16681 = ~n16673 | ~n16672;
  assign n16679 = ~n21356 | ~P2_REG2_REG_11__SCAN_IN;
  assign n16675 = ~n16674 & ~P2_REG3_REG_11__SCAN_IN;
  assign n24941 = n16676 | n16675;
  assign n16677 = ~n24941;
  assign n16678 = ~n17780 | ~n16677;
  assign n16680 = ~n16679 | ~n16678;
  assign n16683 = ~P2_U3947 | ~n24976;
  assign n16682 = ~n25592 | ~P2_DATAO_REG_11__SCAN_IN;
  assign P2_U3542 = ~n16683 | ~n16682;
  assign n16685 = ~n16780 | ~P2_REG1_REG_10__SCAN_IN;
  assign n16684 = ~n16781 | ~P2_REG0_REG_10__SCAN_IN;
  assign n16690 = ~n16685 | ~n16684;
  assign n16688 = ~n21356 | ~P2_REG2_REG_10__SCAN_IN;
  assign n24964 = n16686 ^ ~P2_REG3_REG_10__SCAN_IN;
  assign n16687 = ~n17780 | ~n24964;
  assign n16689 = ~n16688 | ~n16687;
  assign n16692 = ~P2_U3947 | ~n25000;
  assign n16691 = ~n25592 | ~P2_DATAO_REG_10__SCAN_IN;
  assign P2_U3541 = ~n16692 | ~n16691;
  assign n16694 = ~n16780 | ~P2_REG1_REG_3__SCAN_IN;
  assign n16693 = ~n16781 | ~P2_REG0_REG_3__SCAN_IN;
  assign n16698 = ~n16694 | ~n16693;
  assign n16696 = ~n21356 | ~P2_REG2_REG_3__SCAN_IN;
  assign n25188 = ~P2_REG3_REG_3__SCAN_IN;
  assign n16695 = ~n17780 | ~n25188;
  assign n16697 = ~n16696 | ~n16695;
  assign n16700 = ~P2_U3947 | ~n25214;
  assign n16699 = ~n25592 | ~P2_DATAO_REG_3__SCAN_IN;
  assign P2_U3534 = ~n16700 | ~n16699;
  assign n24474 = n16701 ^ ~P2_REG3_REG_13__SCAN_IN;
  assign n16703 = ~n17780 | ~n24474;
  assign n16702 = ~n16780 | ~P2_REG1_REG_13__SCAN_IN;
  assign n16707 = ~n16703 | ~n16702;
  assign n16705 = ~n21356 | ~P2_REG2_REG_13__SCAN_IN;
  assign n16704 = ~n16781 | ~P2_REG0_REG_13__SCAN_IN;
  assign n16706 = ~n16705 | ~n16704;
  assign n16709 = ~P2_U3947 | ~n21817;
  assign n16708 = ~n25592 | ~P2_DATAO_REG_13__SCAN_IN;
  assign P2_U3544 = ~n16709 | ~n16708;
  assign n16711 = ~n16780 | ~P2_REG1_REG_7__SCAN_IN;
  assign n16710 = ~n16781 | ~P2_REG0_REG_7__SCAN_IN;
  assign n16720 = ~n16711 | ~n16710;
  assign n16718 = ~n21356 | ~P2_REG2_REG_7__SCAN_IN;
  assign n16713 = ~n16725 | ~P2_REG3_REG_6__SCAN_IN;
  assign n16712 = ~P2_REG3_REG_7__SCAN_IN;
  assign n16715 = ~n16713 | ~n16712;
  assign n25059 = ~n16715 | ~n16714;
  assign n16716 = ~n25059;
  assign n16717 = ~n17780 | ~n16716;
  assign n16719 = ~n16718 | ~n16717;
  assign n16722 = ~P2_U3947 | ~n25022;
  assign n16721 = ~n25592 | ~P2_DATAO_REG_7__SCAN_IN;
  assign P2_U3538 = ~n16722 | ~n16721;
  assign n16724 = ~n16780 | ~P2_REG1_REG_6__SCAN_IN;
  assign n16723 = ~n16781 | ~P2_REG0_REG_6__SCAN_IN;
  assign n16730 = ~n16724 | ~n16723;
  assign n16728 = ~n21356 | ~P2_REG2_REG_6__SCAN_IN;
  assign n25073 = n16725 ^ ~P2_REG3_REG_6__SCAN_IN;
  assign n16726 = ~n25073;
  assign n16727 = ~n17780 | ~n16726;
  assign n16729 = ~n16728 | ~n16727;
  assign n16732 = ~P2_U3947 | ~n25126;
  assign n16731 = ~n25592 | ~P2_DATAO_REG_6__SCAN_IN;
  assign P2_U3537 = ~n16732 | ~n16731;
  assign n16733 = ~n21356 | ~P2_REG2_REG_5__SCAN_IN;
  assign n25106 = n16742 ^ ~P2_REG3_REG_5__SCAN_IN;
  assign n16735 = ~n17780 | ~n25106;
  assign n16734 = ~n16780 | ~P2_REG1_REG_5__SCAN_IN;
  assign n16736 = ~n16735 | ~n16734;
  assign n16738 = ~P2_U3947 | ~n25150;
  assign n16737 = ~n25592 | ~P2_DATAO_REG_5__SCAN_IN;
  assign P2_U3536 = ~n16738 | ~n16737;
  assign n16740 = ~n16780 | ~P2_REG1_REG_4__SCAN_IN;
  assign n16739 = ~n16781 | ~P2_REG0_REG_4__SCAN_IN;
  assign n16747 = ~n16740 | ~n16739;
  assign n16745 = ~n21356 | ~P2_REG2_REG_4__SCAN_IN;
  assign n16741 = ~P2_REG3_REG_4__SCAN_IN;
  assign n16743 = ~n25188 | ~n16741;
  assign n24429 = ~n16743 | ~n16742;
  assign n25160 = ~n24429;
  assign n16744 = ~n17780 | ~n25160;
  assign n16746 = ~n16745 | ~n16744;
  assign n25183 = n16747 | n16746;
  assign n16749 = ~P2_U3947 | ~n25183;
  assign n16748 = ~n25592 | ~P2_DATAO_REG_4__SCAN_IN;
  assign P2_U3535 = ~n16749 | ~n16748;
  assign n16750 = ~P2_REG3_REG_16__SCAN_IN;
  assign n21778 = n16751 ^ ~n16750;
  assign n16753 = ~n21778 | ~n17780;
  assign n16752 = ~n21356 | ~P2_REG2_REG_16__SCAN_IN;
  assign n16757 = ~n16753 | ~n16752;
  assign n16755 = ~n16780 | ~P2_REG1_REG_16__SCAN_IN;
  assign n16754 = ~n16781 | ~P2_REG0_REG_16__SCAN_IN;
  assign n16756 = ~n16755 | ~n16754;
  assign n16759 = ~P2_U3947 | ~n21735;
  assign n16758 = ~n25592 | ~P2_DATAO_REG_16__SCAN_IN;
  assign P2_U3547 = ~n16759 | ~n16758;
  assign n16761 = ~P1_U4016 | ~n23853;
  assign n16760 = ~n24319 | ~P1_DATAO_REG_7__SCAN_IN;
  assign P1_U3567 = ~n16761 | ~n16760;
  assign n16763 = ~P1_U4016 | ~n23875;
  assign n16762 = ~n24319 | ~P1_DATAO_REG_6__SCAN_IN;
  assign P1_U3566 = ~n16763 | ~n16762;
  assign n16765 = ~P1_U4016 | ~n23801;
  assign n16764 = ~n24319 | ~P1_DATAO_REG_9__SCAN_IN;
  assign P1_U3569 = ~n16765 | ~n16764;
  assign n16767 = ~P1_U4016 | ~n23874;
  assign n16766 = ~n24319 | ~P1_DATAO_REG_4__SCAN_IN;
  assign P1_U3564 = ~n16767 | ~n16766;
  assign n16769 = ~n17780 | ~P2_REG3_REG_0__SCAN_IN;
  assign n16768 = ~n16780 | ~P2_REG1_REG_0__SCAN_IN;
  assign n16773 = ~n16769 | ~n16768;
  assign n16770 = ~n16781 | ~P2_REG0_REG_0__SCAN_IN;
  assign n16772 = ~n16771 | ~n16770;
  assign n16775 = ~P2_U3947 | ~n25254;
  assign n16774 = ~n25592 | ~P2_DATAO_REG_0__SCAN_IN;
  assign P2_U3531 = ~n16775 | ~n16774;
  assign n16776 = ~P2_REG3_REG_1__SCAN_IN;
  assign n16785 = ~n16779 | ~n16778;
  assign n16783 = ~n16780 | ~P2_REG1_REG_1__SCAN_IN;
  assign n16782 = ~n16781 | ~P2_REG0_REG_1__SCAN_IN;
  assign n16784 = ~n16783 | ~n16782;
  assign n16787 = ~P2_U3947 | ~n25274;
  assign n16786 = ~n25592 | ~P2_DATAO_REG_1__SCAN_IN;
  assign P2_U3532 = ~n16787 | ~n16786;
  assign n16788 = P1_DATAO_REG_14__SCAN_IN ^ ~P2_DATAO_REG_14__SCAN_IN;
  assign n16796 = ~n18219 | ~n17285;
  assign n16791 = ~n16790 | ~P3_IR_REG_31__SCAN_IN;
  assign n19997 = n16791 ^ ~P3_IR_REG_14__SCAN_IN;
  assign n26036 = ~n19997;
  assign n16794 = ~n26036 & ~P3_U3151;
  assign n16793 = ~n20796 & ~n16792;
  assign n16795 = ~n16794 & ~n16793;
  assign P3_U3281 = ~n16796 | ~n16795;
  assign n16797 = ~P3_REG3_REG_18__SCAN_IN;
  assign n16799 = ~n16798 & ~n16797;
  assign n20381 = n16851 | n16799;
  assign n16805 = ~n20381 | ~n16484;
  assign n16801 = ~n16463 | ~P3_REG1_REG_18__SCAN_IN;
  assign n16800 = ~n18380 | ~P3_REG0_REG_18__SCAN_IN;
  assign n16803 = ~n16801 | ~n16800;
  assign n20391 = ~P3_REG2_REG_18__SCAN_IN;
  assign n16802 = ~n18326 & ~n20391;
  assign n16804 = ~n16803 & ~n16802;
  assign n16807 = ~n19674 | ~P3_U3897;
  assign n16806 = ~n26454 | ~P3_DATAO_REG_18__SCAN_IN;
  assign P3_U3509 = ~n16807 | ~n16806;
  assign n23219 = ~P1_REG3_REG_3__SCAN_IN | ~P1_U3086;
  assign n18905 = ~n16808 & ~P1_U3086;
  assign n18908 = ~n18905;
  assign n16817 = ~n24033 | ~n18908;
  assign n16810 = ~n17377 | ~n16808;
  assign n16815 = ~n16810 | ~n16809;
  assign n16811 = ~P1_ADDR_REG_3__SCAN_IN | ~n23729;
  assign n16831 = ~n23219 | ~n16811;
  assign n23409 = n17949 ^ ~P1_REG2_REG_3__SCAN_IN;
  assign n23364 = n16823 ^ ~P1_REG2_REG_1__SCAN_IN;
  assign n23363 = ~P1_IR_REG_0__SCAN_IN | ~P1_REG2_REG_0__SCAN_IN;
  assign n23390 = ~n23363;
  assign n16813 = ~n23364 | ~n23390;
  assign n23366 = ~n16823;
  assign n16812 = ~n23366 | ~P1_REG2_REG_1__SCAN_IN;
  assign n23401 = ~n16813 | ~n16812;
  assign n23400 = n24107 ^ ~P1_REG2_REG_2__SCAN_IN;
  assign n23399 = ~n23401 | ~n23400;
  assign n23380 = ~n24107;
  assign n16814 = ~n23380 | ~P1_REG2_REG_2__SCAN_IN;
  assign n23410 = ~n23399 | ~n16814;
  assign n16820 = n23409 ^ n23410;
  assign n16816 = ~n16815;
  assign n23356 = ~n16817 | ~n16816;
  assign n16819 = n23351 | n16818;
  assign n23720 = ~n23356 & ~n16819;
  assign n16829 = ~n16820 | ~n23720;
  assign n16821 = ~n16818;
  assign n23501 = n23356 | n16821;
  assign n16822 = ~P1_REG1_REG_1__SCAN_IN;
  assign n23372 = n16823 ^ ~n16822;
  assign n23371 = ~P1_IR_REG_0__SCAN_IN | ~P1_REG1_REG_0__SCAN_IN;
  assign n23374 = n23372 | n23371;
  assign n16824 = n16823 | n16822;
  assign n23382 = ~n23374 | ~n16824;
  assign n23381 = n24107 ^ ~P1_REG1_REG_2__SCAN_IN;
  assign n16826 = ~n23382 | ~n23381;
  assign n16825 = ~n23380 | ~P1_REG1_REG_2__SCAN_IN;
  assign n23414 = ~n16826 | ~n16825;
  assign n23415 = n17949 ^ ~P1_REG1_REG_3__SCAN_IN;
  assign n16827 = n23414 ^ n23415;
  assign n16828 = ~n23722 | ~n16827;
  assign n16830 = ~n16829 | ~n16828;
  assign n16833 = ~n16831 & ~n16830;
  assign n23416 = ~n17949;
  assign n16832 = ~n23688 | ~n23416;
  assign P1_U3246 = ~n16833 | ~n16832;
  assign n16841 = n16928 ^ P2_ADDR_REG_7__SCAN_IN;
  assign n16837 = ~P3_ADDR_REG_7__SCAN_IN;
  assign n16921 = ~n16838 | ~P3_ADDR_REG_7__SCAN_IN;
  assign n16920 = n16839 & n16921;
  assign n16840 = ~n16920;
  assign n16919 = ~P1_ADDR_REG_7__SCAN_IN;
  assign n16932 = n16840 ^ ~n16919;
  assign SUB_1596_U56 = n16841 ^ ~n16932;
  assign P1_U3085 = ~n23729 & ~n24307;
  assign n19587 = n16851 ^ ~P3_REG3_REG_19__SCAN_IN;
  assign n16842 = ~n16484;
  assign n16848 = n19587 | n16842;
  assign n16844 = ~n18368 | ~P3_REG1_REG_19__SCAN_IN;
  assign n16843 = ~n18380 | ~P3_REG0_REG_19__SCAN_IN;
  assign n16846 = ~n16844 | ~n16843;
  assign n20366 = ~P3_REG2_REG_19__SCAN_IN;
  assign n16845 = ~n18326 & ~n20366;
  assign n16847 = ~n16846 & ~n16845;
  assign n16850 = ~n19446 | ~P3_U3897;
  assign n16849 = ~n26454 | ~P3_DATAO_REG_19__SCAN_IN;
  assign P3_U3510 = ~n16850 | ~n16849;
  assign n19583 = ~P3_REG3_REG_19__SCAN_IN;
  assign n16853 = ~n16852 | ~P3_REG3_REG_20__SCAN_IN;
  assign n20342 = ~n16899 | ~n16853;
  assign n16859 = ~n20342 | ~n16484;
  assign n16855 = ~n16422 | ~P3_REG2_REG_20__SCAN_IN;
  assign n16854 = ~n18368 | ~P3_REG1_REG_20__SCAN_IN;
  assign n16857 = ~n16855 | ~n16854;
  assign n16856 = n18380 & P3_REG0_REG_20__SCAN_IN;
  assign n16858 = ~n16857 & ~n16856;
  assign n19602 = ~n16859 | ~n16858;
  assign n16861 = ~n19602 | ~P3_U3897;
  assign n16860 = ~n26454 | ~P3_DATAO_REG_20__SCAN_IN;
  assign P3_U3511 = ~n16861 | ~n16860;
  assign n16863 = ~n23016 | ~P1_U4016;
  assign n16862 = ~n24319 | ~P1_DATAO_REG_15__SCAN_IN;
  assign P1_U3575 = ~n16863 | ~n16862;
  assign n16865 = ~n22999 | ~n24307;
  assign n16864 = ~n24319 | ~P1_DATAO_REG_16__SCAN_IN;
  assign P1_U3576 = ~n16865 | ~n16864;
  assign n16867 = ~n24307 | ~n23254;
  assign n16866 = ~n24319 | ~P1_DATAO_REG_2__SCAN_IN;
  assign P1_U3562 = ~n16867 | ~n16866;
  assign n16869 = ~n24307 | ~n23993;
  assign n16868 = ~n24319 | ~P1_DATAO_REG_0__SCAN_IN;
  assign P1_U3560 = ~n16869 | ~n16868;
  assign n18228 = n16871 ^ ~n16870;
  assign n16877 = ~n18228 & ~n20792;
  assign n16873 = ~n16872 | ~P3_IR_REG_31__SCAN_IN;
  assign n19999 = n16873 ^ ~P3_IR_REG_15__SCAN_IN;
  assign n16875 = ~n19999 | ~P3_STATE_REG_SCAN_IN;
  assign n16874 = ~n20774 | ~SI_15_;
  assign n16876 = ~n16875 | ~n16874;
  assign P3_U3280 = n16877 | n16876;
  assign n16883 = ~n17624 | ~n22164;
  assign n16879 = n16878 | n17032;
  assign n24863 = n16879 ^ ~P2_IR_REG_15__SCAN_IN;
  assign n24842 = ~n24863;
  assign n16881 = ~n24842 & ~P2_U3088;
  assign n17625 = ~P1_DATAO_REG_15__SCAN_IN;
  assign n16880 = ~n25337 & ~n17625;
  assign n16882 = ~n16881 & ~n16880;
  assign P2_U3312 = ~n16883 | ~n16882;
  assign n16888 = ~n17624 | ~n23156;
  assign n16886 = ~n24085 & ~n16884;
  assign n16885 = ~n23632 & ~P1_U3086;
  assign n16887 = ~n16886 & ~n16885;
  assign P1_U3340 = ~n16888 | ~n16887;
  assign n18236 = n16889 ^ ~n16890;
  assign n16898 = n18236 | n20792;
  assign n16892 = ~n16891;
  assign n16894 = ~n16892 | ~P3_IR_REG_16__SCAN_IN;
  assign n20059 = ~n20034;
  assign n16896 = ~n20059 & ~P3_U3151;
  assign n18238 = ~SI_16_;
  assign n16895 = ~n20796 & ~n18238;
  assign n16897 = ~n16896 & ~n16895;
  assign P3_U3279 = ~n16898 | ~n16897;
  assign n16900 = n16899 & P3_REG3_REG_21__SCAN_IN;
  assign n20321 = n16900 | n16939;
  assign n16906 = ~n20321 | ~n16484;
  assign n16902 = ~n16460 | ~P3_REG2_REG_21__SCAN_IN;
  assign n16901 = ~n18380 | ~P3_REG0_REG_21__SCAN_IN;
  assign n16904 = ~n16902 | ~n16901;
  assign n16903 = n18368 & P3_REG1_REG_21__SCAN_IN;
  assign n16905 = ~n16904 & ~n16903;
  assign n16908 = ~n19752 | ~P3_U3897;
  assign n16907 = ~n26454 | ~P3_DATAO_REG_21__SCAN_IN;
  assign P3_U3512 = ~n16908 | ~n16907;
  assign n16938 = ~P3_REG3_REG_22__SCAN_IN;
  assign n16909 = ~P3_REG3_REG_23__SCAN_IN;
  assign n16910 = n16941 | n16909;
  assign n20273 = ~n17091 | ~n16910;
  assign n16916 = ~n20273 | ~n16484;
  assign n16912 = ~n16460 | ~P3_REG2_REG_23__SCAN_IN;
  assign n16911 = ~n16463 | ~P3_REG1_REG_23__SCAN_IN;
  assign n16914 = ~n16912 | ~n16911;
  assign n16913 = n18380 & P3_REG0_REG_23__SCAN_IN;
  assign n16915 = ~n16914 & ~n16913;
  assign n19692 = ~n16916 | ~n16915;
  assign n16918 = ~n19692 | ~P3_U3897;
  assign n16917 = ~n26454 | ~P3_DATAO_REG_23__SCAN_IN;
  assign P3_U3514 = ~n16918 | ~n16917;
  assign n16922 = ~P3_ADDR_REG_8__SCAN_IN;
  assign n16925 = ~P1_ADDR_REG_8__SCAN_IN;
  assign n16927 = ~n16926 | ~P1_ADDR_REG_8__SCAN_IN;
  assign n16931 = ~n16928 | ~P2_ADDR_REG_7__SCAN_IN;
  assign n16936 = ~n16930;
  assign n16934 = ~n16932 | ~n16931;
  assign n16935 = n16934 & n16933;
  assign n17256 = ~n16936 | ~n16935;
  assign SUB_1596_U55 = n16937 ^ ~P2_ADDR_REG_8__SCAN_IN;
  assign n16940 = ~n16939 & ~n16938;
  assign n20299 = n16941 | n16940;
  assign n16947 = ~n20299 | ~n16484;
  assign n16943 = ~n16422 | ~P3_REG2_REG_22__SCAN_IN;
  assign n16942 = ~n18380 | ~P3_REG0_REG_22__SCAN_IN;
  assign n16945 = ~n16943 | ~n16942;
  assign n16944 = n18368 & P3_REG1_REG_22__SCAN_IN;
  assign n16946 = ~n16945 & ~n16944;
  assign n16949 = ~n20267 | ~P3_U3897;
  assign n16948 = ~n26454 | ~P3_DATAO_REG_22__SCAN_IN;
  assign P3_U3513 = ~n16949 | ~n16948;
  assign n16950 = ~n25297 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n16952 = ~n24041 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n16953 = P1_DATAO_REG_18__SCAN_IN ^ ~P2_DATAO_REG_18__SCAN_IN;
  assign n18248 = n17076 ^ ~n16953;
  assign n16965 = n18248 | n20792;
  assign n16957 = ~n16956 | ~P3_IR_REG_31__SCAN_IN;
  assign n16959 = ~n16957 | ~P3_IR_REG_18__SCAN_IN;
  assign n16961 = ~n16959 | ~n16958;
  assign n20106 = ~n16961 | ~n17084;
  assign n16963 = ~n20106 & ~P3_U3151;
  assign n16962 = ~n20796 & ~n18249;
  assign n16964 = ~n16963 & ~n16962;
  assign P3_U3277 = ~n16965 | ~n16964;
  assign n16967 = ~n23331 | ~n24122;
  assign n16966 = ~n23332 | ~n17382;
  assign n16971 = ~n16967 | ~n16966;
  assign n23389 = n16969 ^ ~n16968;
  assign n16970 = n23389 & n23339;
  assign n16974 = ~n16971 & ~n16970;
  assign n23319 = ~n18907 | ~n16972;
  assign n16973 = ~P1_REG3_REG_0__SCAN_IN | ~n23319;
  assign P1_U3232 = ~n16974 | ~n16973;
  assign n16975 = n17324 ^ ~P2_B_REG_SCAN_IN;
  assign n16976 = ~n16975 | ~n22165;
  assign n16982 = ~P2_D_REG_6__SCAN_IN & ~P2_D_REG_7__SCAN_IN;
  assign n16980 = P2_D_REG_8__SCAN_IN | P2_D_REG_9__SCAN_IN;
  assign n16978 = ~P2_D_REG_10__SCAN_IN & ~P2_D_REG_11__SCAN_IN;
  assign n16977 = ~P2_D_REG_12__SCAN_IN & ~P2_D_REG_13__SCAN_IN;
  assign n16979 = ~n16978 | ~n16977;
  assign n16981 = ~n16980 & ~n16979;
  assign n16998 = ~n16982 | ~n16981;
  assign n16984 = ~P2_D_REG_18__SCAN_IN & ~P2_D_REG_19__SCAN_IN;
  assign n16983 = ~P2_D_REG_20__SCAN_IN & ~P2_D_REG_21__SCAN_IN;
  assign n16988 = ~n16984 | ~n16983;
  assign n16986 = ~P2_D_REG_16__SCAN_IN & ~P2_D_REG_14__SCAN_IN;
  assign n16985 = ~P2_D_REG_15__SCAN_IN & ~P2_D_REG_17__SCAN_IN;
  assign n16987 = ~n16986 | ~n16985;
  assign n16996 = ~n16988 & ~n16987;
  assign n16990 = ~P2_D_REG_26__SCAN_IN & ~P2_D_REG_27__SCAN_IN;
  assign n16989 = ~P2_D_REG_28__SCAN_IN & ~P2_D_REG_31__SCAN_IN;
  assign n16994 = ~n16990 | ~n16989;
  assign n16992 = ~P2_D_REG_22__SCAN_IN & ~P2_D_REG_23__SCAN_IN;
  assign n16991 = ~P2_D_REG_24__SCAN_IN & ~P2_D_REG_25__SCAN_IN;
  assign n16993 = ~n16992 | ~n16991;
  assign n16995 = ~n16994 & ~n16993;
  assign n16997 = ~n16996 | ~n16995;
  assign n17003 = ~n16998 & ~n16997;
  assign n17000 = ~P2_D_REG_2__SCAN_IN & ~P2_D_REG_3__SCAN_IN;
  assign n16999 = ~P2_D_REG_4__SCAN_IN & ~P2_D_REG_5__SCAN_IN;
  assign n17001 = ~n17000 | ~n16999;
  assign n17002 = ~P2_D_REG_30__SCAN_IN & ~n17001;
  assign n17004 = ~n17003 | ~n17002;
  assign n17005 = ~P2_D_REG_29__SCAN_IN & ~n17004;
  assign n17862 = ~n25289 & ~n17005;
  assign n25374 = ~n22156 & ~n17006;
  assign n17007 = ~P2_D_REG_1__SCAN_IN & ~n25289;
  assign n25370 = ~n22156 & ~n17008;
  assign n17009 = ~P2_D_REG_0__SCAN_IN & ~n25289;
  assign n17010 = ~n18106 | ~n18145;
  assign n17069 = ~n17058 | ~n25373;
  assign n17012 = ~n17013 | ~P2_IR_REG_31__SCAN_IN;
  assign n17030 = n17012 ^ ~P2_IR_REG_22__SCAN_IN;
  assign n21030 = ~n17030;
  assign n17016 = n17015 | n17014;
  assign n17018 = ~P2_IR_REG_20__SCAN_IN;
  assign n17019 = ~n17018 | ~P2_IR_REG_31__SCAN_IN;
  assign n17024 = ~n17017 | ~P2_IR_REG_31__SCAN_IN;
  assign n17026 = ~n17025 | ~n17024;
  assign n17027 = ~n21032;
  assign n25441 = ~n25378 | ~n17027;
  assign n17028 = ~n25441 | ~n21031;
  assign n17031 = ~n17030 | ~n17029;
  assign n17032 = ~P2_IR_REG_31__SCAN_IN;
  assign n17035 = ~n17033 | ~P2_IR_REG_31__SCAN_IN;
  assign n17034 = ~P2_IR_REG_27__SCAN_IN;
  assign n17041 = ~n17040 | ~n17039;
  assign n17043 = ~n24333 | ~n17042;
  assign n24454 = ~n17044 | ~n17043;
  assign n17045 = ~n19033 | ~n14816;
  assign n17047 = n13406 | n17046;
  assign n17048 = ~n17047 | ~n18916;
  assign n17057 = ~n24506 | ~n17048;
  assign n21401 = ~n25373 | ~n21032;
  assign n17050 = ~n21031;
  assign n25092 = ~n17050 | ~n17049;
  assign n17051 = ~n21401 & ~n25092;
  assign n17498 = ~n25252;
  assign n17055 = ~n24499 & ~n17498;
  assign n17052 = ~n21401 & ~n25079;
  assign n24484 = ~n17058 | ~n17052;
  assign n17053 = ~n25254;
  assign n17054 = ~n24484 & ~n17053;
  assign n17056 = ~n17055 & ~n17054;
  assign n17068 = ~n17057 | ~n17056;
  assign n17063 = ~n17058;
  assign n17061 = ~n17063 | ~n25441;
  assign n17860 = n21031 | n21032;
  assign n17060 = n17059 & n17860;
  assign n17062 = ~n17061 | ~n17060;
  assign n17066 = ~n17062 | ~P2_STATE_REG_SCAN_IN;
  assign n17290 = n21407 | P2_U3088;
  assign n17064 = ~n17290;
  assign n17065 = ~n17064 | ~n17063;
  assign n24487 = ~n24475 & ~P2_U3088;
  assign n17067 = ~n24487 & ~n16776;
  assign n17074 = ~n17068 & ~n17067;
  assign n21417 = ~n21407;
  assign n25091 = ~n25378 | ~n21417;
  assign n17072 = n17069 | n25091;
  assign n17070 = ~n21407 | ~n25194;
  assign n17073 = ~n24508 | ~n25389;
  assign P2_U3194 = ~n17074 | ~n17073;
  assign n25291 = ~P1_DATAO_REG_18__SCAN_IN;
  assign n17075 = ~n25291 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n17078 = ~n17077 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n17079 = P1_DATAO_REG_19__SCAN_IN ^ ~P2_DATAO_REG_19__SCAN_IN;
  assign n18256 = n17270 ^ ~n17079;
  assign n17090 = n18256 | n20792;
  assign n17080 = ~n17084 | ~P3_IR_REG_31__SCAN_IN;
  assign n17083 = ~n17080 | ~P3_IR_REG_19__SCAN_IN;
  assign n17081 = ~P3_IR_REG_19__SCAN_IN;
  assign n17082 = ~n17081 | ~P3_IR_REG_31__SCAN_IN;
  assign n17086 = ~n17083 | ~n17082;
  assign n17085 = ~n17084;
  assign n17137 = ~n17085 | ~n17081;
  assign n20119 = ~n17086 | ~n17137;
  assign n17088 = ~n20119 & ~P3_U3151;
  assign n18257 = ~SI_19_;
  assign n17087 = ~n20796 & ~n18257;
  assign n17089 = ~n17088 & ~n17087;
  assign P3_U3276 = ~n17090 | ~n17089;
  assign n17092 = ~n17091 | ~P3_REG3_REG_24__SCAN_IN;
  assign n20246 = ~n18323 | ~n17092;
  assign n17098 = ~n20246 | ~n16484;
  assign n17094 = ~n16422 | ~P3_REG2_REG_24__SCAN_IN;
  assign n17093 = ~n18368 | ~P3_REG1_REG_24__SCAN_IN;
  assign n17096 = ~n17094 | ~n17093;
  assign n17095 = n18380 & P3_REG0_REG_24__SCAN_IN;
  assign n17097 = ~n17096 & ~n17095;
  assign n20266 = ~n17098 | ~n17097;
  assign n17100 = ~n20266 | ~P3_U3897;
  assign n17099 = ~n26454 | ~P3_DATAO_REG_24__SCAN_IN;
  assign P3_U3515 = ~n17100 | ~n17099;
  assign n26310 = ~n20786 | ~n20794;
  assign n17103 = ~P3_D_REG_2__SCAN_IN & ~P3_D_REG_3__SCAN_IN;
  assign n17102 = ~P3_D_REG_4__SCAN_IN & ~P3_D_REG_5__SCAN_IN;
  assign n17104 = ~n17103 | ~n17102;
  assign n17130 = ~P3_D_REG_30__SCAN_IN & ~n17104;
  assign n17112 = ~P3_D_REG_6__SCAN_IN & ~P3_D_REG_7__SCAN_IN;
  assign n17110 = ~n17106 | ~n17105;
  assign n17108 = ~P3_D_REG_10__SCAN_IN & ~P3_D_REG_11__SCAN_IN;
  assign n17107 = ~P3_D_REG_12__SCAN_IN & ~P3_D_REG_13__SCAN_IN;
  assign n17109 = ~n17108 | ~n17107;
  assign n17111 = ~n17110 & ~n17109;
  assign n17128 = ~n17112 | ~n17111;
  assign n17114 = ~P3_D_REG_18__SCAN_IN & ~P3_D_REG_19__SCAN_IN;
  assign n17113 = ~P3_D_REG_20__SCAN_IN & ~P3_D_REG_21__SCAN_IN;
  assign n17118 = ~n17114 | ~n17113;
  assign n17116 = ~P3_D_REG_16__SCAN_IN & ~P3_D_REG_14__SCAN_IN;
  assign n17115 = ~P3_D_REG_15__SCAN_IN & ~P3_D_REG_17__SCAN_IN;
  assign n17117 = ~n17116 | ~n17115;
  assign n17126 = ~n17118 & ~n17117;
  assign n17120 = ~P3_D_REG_26__SCAN_IN & ~P3_D_REG_27__SCAN_IN;
  assign n17119 = ~P3_D_REG_28__SCAN_IN & ~P3_D_REG_31__SCAN_IN;
  assign n17124 = ~n17120 | ~n17119;
  assign n17122 = ~P3_D_REG_22__SCAN_IN & ~P3_D_REG_23__SCAN_IN;
  assign n17121 = ~P3_D_REG_24__SCAN_IN & ~P3_D_REG_25__SCAN_IN;
  assign n17123 = ~n17122 | ~n17121;
  assign n17125 = ~n17124 & ~n17123;
  assign n17127 = ~n17126 | ~n17125;
  assign n17129 = ~n17128 & ~n17127;
  assign n17131 = ~n17130 | ~n17129;
  assign n17132 = P3_D_REG_29__SCAN_IN | n17131;
  assign n17155 = n17133 & n17132;
  assign n18449 = ~n17155;
  assign n17136 = ~n18449 | ~n18448;
  assign n17171 = n18482 | n17136;
  assign n18467 = ~n17171;
  assign n17139 = ~n17137 | ~P3_IR_REG_31__SCAN_IN;
  assign n19522 = n17139 ^ ~n17138;
  assign n17190 = ~n19522;
  assign n17141 = ~n17140;
  assign n17142 = ~n17141 | ~P3_IR_REG_31__SCAN_IN;
  assign n17145 = ~n17142 | ~P3_IR_REG_21__SCAN_IN;
  assign n17144 = ~n17143 | ~P3_IR_REG_31__SCAN_IN;
  assign n17146 = ~n17145 | ~n17144;
  assign n19301 = n17190 & n19306;
  assign n17148 = ~n17147 | ~P3_IR_REG_31__SCAN_IN;
  assign n17151 = ~n17148 | ~P3_IR_REG_22__SCAN_IN;
  assign n17149 = ~P3_IR_REG_22__SCAN_IN;
  assign n17150 = ~n17149 | ~P3_IR_REG_31__SCAN_IN;
  assign n17153 = ~n17151 | ~n17150;
  assign n18454 = ~n18443 & ~n20119;
  assign n18468 = n19301 & n18454;
  assign n17154 = ~n18468;
  assign n17164 = ~n18467 & ~n17154;
  assign n17156 = ~n18448 & ~n17155;
  assign n18470 = n17156 & n18482;
  assign n17157 = ~n18443 & ~n19308;
  assign n17159 = ~n19522 | ~n17157;
  assign n17158 = ~n20119 | ~n19306;
  assign n17161 = n17159 & n17158;
  assign n17160 = n17190 | n19308;
  assign n18457 = ~n17160 | ~n18443;
  assign n18465 = n17161 & n18457;
  assign n17162 = n18470 | n18465;
  assign n17163 = ~n19831 | ~n17162;
  assign n17166 = ~n17164 & ~n17163;
  assign n18453 = n19520 | n18455;
  assign n17165 = n18453 & n19835;
  assign n17167 = ~n17166 | ~n17165;
  assign n17169 = ~P3_STATE_REG_SCAN_IN | ~n17167;
  assign n19834 = ~n19364;
  assign n19524 = n18473 & n26303;
  assign n17168 = ~n17171 | ~n19524;
  assign n17252 = ~n25734 | ~n26213;
  assign n17170 = ~n19524;
  assign n17238 = ~n17171 & ~n17170;
  assign n17173 = ~n17174 | ~P3_IR_REG_26__SCAN_IN;
  assign n17176 = ~n17173 | ~P3_IR_REG_31__SCAN_IN;
  assign n17175 = ~n17174 | ~n16337;
  assign n17181 = ~n17178 | ~P3_IR_REG_28__SCAN_IN;
  assign n17182 = ~n17181 | ~n17180;
  assign n20000 = n20078 | n20773;
  assign n18191 = ~n19847 | ~n20773;
  assign n18258 = ~n17198;
  assign n18387 = n20000 & n18258;
  assign n17183 = ~n18387;
  assign n25728 = ~n25666;
  assign n17250 = ~n25728 | ~n26205;
  assign n25819 = ~P3_REG3_REG_4__SCAN_IN | ~P3_U3151;
  assign n17248 = ~n25819;
  assign n17186 = ~n18467 | ~n18468;
  assign n17184 = ~n18465 & ~n26315;
  assign n17185 = ~n18470 | ~n17184;
  assign n17187 = ~n17186 | ~n17185;
  assign n25732 = n17187 & n18473;
  assign n17188 = ~n18448;
  assign n17192 = ~n17188 | ~n19301;
  assign n17189 = ~n20119 & ~n19308;
  assign n17191 = n17190 | n17189;
  assign n17195 = n18191 | n19840;
  assign n17194 = ~n18191 | ~n17193;
  assign n26277 = ~n17195 | ~n17194;
  assign n17200 = n19228 | n17197;
  assign n17199 = ~n17198 | ~P3_IR_REG_0__SCAN_IN;
  assign n17203 = ~n17200 | ~n17199;
  assign n17201 = ~SI_0_;
  assign n17202 = ~n18176 & ~n17201;
  assign n17204 = ~n19178 | ~n14005;
  assign n25659 = ~n26273 | ~n17204;
  assign n25712 = ~n25661 | ~n17205;
  assign n17212 = n18191 | n19967;
  assign n17209 = ~n17206 | ~n17036;
  assign n17208 = ~n13122 | ~n17207;
  assign n17210 = ~n17209 | ~n17208;
  assign n17211 = ~n18258 | ~n17210;
  assign n17214 = n17213 ^ ~n26245;
  assign n17217 = n17214 | n26286;
  assign n17215 = ~n17214;
  assign n18158 = ~n26286;
  assign n17216 = n17215 | n18158;
  assign n25711 = n17217 & n17216;
  assign n25714 = ~n25712 | ~n25711;
  assign n25629 = ~n25714 | ~n17217;
  assign n17224 = ~n25629;
  assign n17220 = n19228 | n17218;
  assign n17219 = n18258 | n25811;
  assign n17222 = ~n17220 | ~n17219;
  assign n17221 = ~n18176 & ~SI_3_;
  assign n17225 = n17213 ^ ~n26335;
  assign n25630 = n17225 ^ ~n26252;
  assign n17223 = ~n25630;
  assign n17227 = ~n17224 | ~n17223;
  assign n17226 = ~n17225 | ~n26252;
  assign n17229 = n18176 | SI_4_;
  assign n17228 = n18258 | n19972;
  assign n17232 = ~n17229 | ~n17228;
  assign n17231 = ~n19228 & ~n17230;
  assign n17233 = n17213 ^ ~n26343;
  assign n19129 = n17233 | n26229;
  assign n17234 = ~n17233 | ~n26229;
  assign n17235 = n19129 & n17234;
  assign n17237 = ~n19130 | ~n17236;
  assign n17246 = ~n25732 | ~n17237;
  assign n17239 = ~n26252;
  assign n25724 = ~n17238 | ~n18387;
  assign n17244 = ~n17239 & ~n25724;
  assign n17240 = n18473 & n26315;
  assign n17242 = ~n18470 | ~n17240;
  assign n26278 = ~n19522 | ~n19257;
  assign n20673 = ~n26315;
  assign n17241 = ~n26278 & ~n20673;
  assign n17243 = ~n25725 & ~n26343;
  assign n17245 = ~n17244 & ~n17243;
  assign n17247 = ~n17246 | ~n17245;
  assign n17249 = ~n17248 & ~n17247;
  assign n17251 = n17250 & n17249;
  assign P3_U3170 = ~n17252 | ~n17251;
  assign n17253 = ~P3_ADDR_REG_9__SCAN_IN;
  assign n17255 = ~n17254 | ~n17253;
  assign n17258 = ~n17257 | ~n17256;
  assign n17309 = ~n17259 | ~n17258;
  assign SUB_1596_U54 = n17260 ^ ~P2_ADDR_REG_9__SCAN_IN;
  assign n17264 = ~n17664 | ~n23156;
  assign n17262 = ~n23905 & ~P1_U3086;
  assign n17261 = ~n24085 & ~n17271;
  assign n17263 = ~n17262 & ~n17261;
  assign P1_U3336 = ~n17264 | ~n17263;
  assign n17268 = ~n17664 | ~n22164;
  assign n17266 = ~n17029 & ~P2_U3088;
  assign n17665 = ~P1_DATAO_REG_19__SCAN_IN;
  assign n17265 = ~n25337 & ~n17665;
  assign n17267 = ~n17266 & ~n17265;
  assign P2_U3308 = ~n17268 | ~n17267;
  assign n17269 = ~n17665 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n17272 = ~n17271 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n18267 = n17299 ^ ~P2_DATAO_REG_20__SCAN_IN;
  assign n17276 = n18267 | n20792;
  assign n17274 = ~n19522 & ~P3_U3151;
  assign n17273 = ~n20796 & ~n18268;
  assign n17275 = ~n17274 & ~n17273;
  assign P3_U3275 = ~n17276 | ~n17275;
  assign n17680 = ~P1_DATAO_REG_20__SCAN_IN;
  assign n17278 = ~n17680 | ~P2_DATAO_REG_20__SCAN_IN;
  assign n17692 = ~P1_DATAO_REG_21__SCAN_IN;
  assign n17277 = ~n17692 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n17279 = n17278 & n17277;
  assign n17282 = ~n17281 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n17706 = ~P1_DATAO_REG_22__SCAN_IN;
  assign n17457 = ~n17706 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n17283 = ~P2_DATAO_REG_22__SCAN_IN;
  assign n17284 = ~n17283 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n17455 = n17457 & n17284;
  assign n18263 = n17456 ^ ~n17455;
  assign n17288 = ~n18263 | ~n17285;
  assign n19305 = ~n18443;
  assign n19526 = ~n19305 & ~P3_U3151;
  assign n17286 = ~n20796 & ~SI_22_;
  assign n17287 = ~n19526 & ~n17286;
  assign P3_U3273 = n17288 & n17287;
  assign n17292 = ~n17679 & ~n25360;
  assign n25365 = ~n25337;
  assign n17289 = ~n25365 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n17291 = ~n17290 | ~n17289;
  assign P2_U3307 = n17292 | n17291;
  assign n17293 = ~n17679;
  assign n17298 = ~n17293 | ~n23156;
  assign n17296 = ~n18853 & ~P1_U3086;
  assign n17295 = ~n24085 & ~n17294;
  assign n17297 = ~n17296 & ~n17295;
  assign P1_U3335 = ~n17298 | ~n17297;
  assign n17301 = ~n17300 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n17304 = ~n17302 | ~n17301;
  assign n17303 = P1_DATAO_REG_21__SCAN_IN ^ ~P2_DATAO_REG_21__SCAN_IN;
  assign n18270 = n17304 ^ ~n17303;
  assign n17308 = n18270 | n20792;
  assign n17306 = ~n19306 & ~P3_U3151;
  assign n17305 = ~n20796 & ~n18271;
  assign n17307 = ~n17306 & ~n17305;
  assign P3_U3274 = ~n17308 | ~n17307;
  assign n17311 = ~P1_ADDR_REG_9__SCAN_IN;
  assign n17313 = ~n17312 | ~n17311;
  assign n17320 = ~n17315 | ~n17316;
  assign n17314 = ~P2_ADDR_REG_10__SCAN_IN;
  assign n17882 = ~n17320 | ~n17314;
  assign n17319 = ~n17882;
  assign n17318 = ~n17315;
  assign n17317 = ~n17316;
  assign n17323 = ~n17319 | ~n17881;
  assign n17321 = ~n17881 | ~n17320;
  assign n17322 = ~n17321 | ~P2_ADDR_REG_10__SCAN_IN;
  assign SUB_1596_U70 = ~n17323 | ~n17322;
  assign n17329 = ~n17732;
  assign n17328 = ~n17329 | ~n22164;
  assign n17326 = ~n17324 & ~P2_U3088;
  assign n18293 = ~P1_DATAO_REG_24__SCAN_IN;
  assign n17325 = ~n25337 & ~n18293;
  assign n17327 = ~n17326 & ~n17325;
  assign P2_U3303 = ~n17328 | ~n17327;
  assign n17335 = ~n17329 | ~n23156;
  assign n17330 = ~n15870;
  assign n17333 = ~n17330 & ~P1_U3086;
  assign n17332 = ~n24085 & ~n17331;
  assign n17334 = ~n17333 & ~n17332;
  assign P1_U3331 = ~n17335 | ~n17334;
  assign n17339 = ~n17691 & ~n24106;
  assign n17337 = n18861 | P1_U3086;
  assign n17336 = ~n24110 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n17338 = ~n17337 | ~n17336;
  assign P1_U3334 = n17339 | n17338;
  assign n17340 = ~n17691;
  assign n17344 = ~n17340 | ~n22164;
  assign n17342 = ~n21456 & ~P2_U3088;
  assign n17341 = ~n25337 & ~n17692;
  assign n17343 = ~n17342 & ~n17341;
  assign P2_U3306 = ~n17344 | ~n17343;
  assign n17705 = n17346 ^ ~n17345;
  assign n17347 = ~n17705;
  assign n17351 = ~n17347 | ~n22164;
  assign n17349 = ~n21030 & ~P2_U3088;
  assign n17348 = ~n25337 & ~n17706;
  assign n17350 = ~n17349 & ~n17348;
  assign P2_U3305 = ~n17351 | ~n17350;
  assign n18868 = ~n17382 | ~n17352;
  assign n17354 = ~n23983 | ~n18868;
  assign n17353 = n23254 & n23967;
  assign n17386 = ~n24000 | ~n24144;
  assign n18869 = ~n17382 & ~n17352;
  assign n17385 = ~n23254 | ~n23967;
  assign n17355 = ~n18869 | ~n17385;
  assign n17356 = n17386 & n17355;
  assign n17358 = ~n23941 | ~n17357;
  assign n18871 = ~n23854 | ~n14266;
  assign n18866 = ~n23874 | ~n23903;
  assign n23880 = ~n23874 & ~n23903;
  assign n17360 = ~n23880 | ~n18871;
  assign n18872 = ~n23906 | ~n23872;
  assign n17361 = n17360 & n18872;
  assign n23828 = ~n24190 | ~n23875;
  assign n17363 = ~n23818 | ~n23853;
  assign n17364 = n23828 & n23831;
  assign n17367 = n24213 | n23825;
  assign n17368 = ~n24231 | ~n23801;
  assign n17395 = n24213 ^ ~n17396;
  assign n23776 = n17395 | n17396;
  assign n17369 = ~n17399;
  assign n17372 = ~n22777 & ~n17369;
  assign n17370 = n23051 | n23753;
  assign n17371 = ~n17370 | ~n22780;
  assign n17373 = ~n17372 & ~n17371;
  assign n17374 = ~n23051 | ~n23753;
  assign n17464 = ~n22257 | ~n22790;
  assign n17376 = ~n18666 | ~n23034;
  assign n18885 = ~n17464 | ~n17376;
  assign n17413 = n17463 ^ ~n18885;
  assign n23914 = n18545 ^ ~n18501;
  assign n17381 = ~n17413 | ~n24012;
  assign n24014 = ~n17377 | ~n23351;
  assign n17379 = ~n22754 & ~n24014;
  assign n22789 = ~n17377 | ~n23391;
  assign n17378 = ~n22207 & ~n22789;
  assign n17380 = ~n17379 & ~n17378;
  assign n17407 = ~n17381 | ~n17380;
  assign n17383 = ~n17382 | ~n24131;
  assign n23950 = n17384 & n17383;
  assign n17387 = ~n24000 | ~n23967;
  assign n17388 = ~n23897;
  assign n17390 = ~n23266 | ~n23903;
  assign n17392 = ~n23906 | ~n14266;
  assign n17393 = ~n23854 | ~n23872;
  assign n17394 = ~n23818 | ~n23234;
  assign n17398 = ~n23794 | ~n23796;
  assign n17397 = n24213 | n17396;
  assign n23739 = ~n24231 | ~n23241;
  assign n22782 = ~n23737 | ~n17400;
  assign n22784 = ~n17400 | ~n23772;
  assign n18883 = n23051 | n22207;
  assign n22783 = n18649 | n14344;
  assign n17401 = n18883 & n22783;
  assign n17402 = n22784 & n17401;
  assign n18882 = ~n23051 | ~n22207;
  assign n17480 = ~n18885;
  assign n17405 = n17481 ^ ~n17480;
  assign n17404 = n18854 | n23905;
  assign n17403 = n18861 | n18853;
  assign n17406 = ~n17405 & ~n23991;
  assign n17433 = ~n17407 & ~n17406;
  assign n17409 = n18907 & n17408;
  assign n22436 = ~n17442 | ~n17409;
  assign n17412 = ~n17433 | ~n24019;
  assign n17410 = ~P1_REG2_REG_12__SCAN_IN;
  assign n17411 = ~n24021 | ~n17410;
  assign n17422 = ~n17412 | ~n17411;
  assign n17426 = ~n17413;
  assign n23970 = ~n18545 | ~n23723;
  assign n17420 = ~n17426 & ~n23892;
  assign n24155 = ~n23941;
  assign n24242 = ~n18649;
  assign n17427 = n17466 ^ ~n22257;
  assign n17418 = ~n17427 | ~n24026;
  assign n23980 = n24021 | n23931;
  assign n17416 = ~n22257 & ~n23980;
  assign n17415 = ~n23936 & ~n17414;
  assign n17417 = ~n17416 & ~n17415;
  assign n17419 = ~n17418 | ~n17417;
  assign n17421 = ~n17420 & ~n17419;
  assign P1_U3281 = ~n17422 | ~n17421;
  assign n17425 = ~n17423 | ~P1_U3086;
  assign n18909 = ~n18854;
  assign n17424 = ~n18909 | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3333 = ~n17425 | ~n17424;
  assign n24220 = ~n24228;
  assign n17431 = ~n17426 & ~n24220;
  assign n24216 = n24123 & n18853;
  assign n17429 = ~n17427 | ~n24216;
  assign n17428 = ~n18666 | ~n24230;
  assign n17430 = ~n17429 | ~n17428;
  assign n17432 = ~n17431 & ~n17430;
  assign n17444 = ~n17433 | ~n17432;
  assign n17435 = n18907 & n17434;
  assign n17437 = ~n17436 | ~n17435;
  assign n17439 = ~n17442;
  assign n17441 = ~n17444 | ~n24251;
  assign n17440 = ~n24240 | ~P1_REG0_REG_12__SCAN_IN;
  assign P1_U3495 = ~n17441 | ~n17440;
  assign n17446 = ~n17444 | ~n24286;
  assign n17445 = ~n24284 | ~P1_REG1_REG_12__SCAN_IN;
  assign P1_U3540 = ~n17446 | ~n17445;
  assign n17450 = ~n17718 | ~n22164;
  assign n21403 = n17447 | P2_U3088;
  assign n21457 = ~n21403;
  assign n18292 = ~P1_DATAO_REG_23__SCAN_IN;
  assign n17448 = ~n25337 & ~n18292;
  assign n17449 = ~n21457 & ~n17448;
  assign P2_U3304 = ~n17450 | ~n17449;
  assign n17454 = ~n17718 | ~n23156;
  assign n17452 = ~n24085 & ~n17451;
  assign n17453 = ~n18905 & ~n17452;
  assign P1_U3332 = ~n17454 | ~n17453;
  assign n18289 = n18292 ^ ~P2_DATAO_REG_23__SCAN_IN;
  assign n18285 = n18291 ^ ~n18289;
  assign n17459 = n18285 & n21363;
  assign n17458 = ~n21363 & ~SI_23_;
  assign n17460 = ~n17459 & ~n17458;
  assign n17462 = ~n17460 & ~P3_STATE_REG_SCAN_IN;
  assign P3_U3272 = ~n17462 & ~n17461;
  assign n22750 = n22341 | n23017;
  assign n17465 = ~n22341 | ~n23017;
  assign n18006 = ~n18887;
  assign n23031 = n18040 ^ ~n18006;
  assign n22752 = ~n24019 | ~n23914;
  assign n17479 = ~n23031 & ~n22752;
  assign n23032 = n13383 ^ ~n22341;
  assign n17477 = ~n23032 | ~n24026;
  assign n23033 = ~n22341;
  assign n17475 = ~n23033 & ~n23980;
  assign n22707 = n24021 | n24014;
  assign n17471 = ~n22707 & ~n22731;
  assign n17469 = ~n24021 | ~P1_REG2_REG_13__SCAN_IN;
  assign n24022 = ~n23936;
  assign n17467 = ~n22337;
  assign n17468 = ~n24022 | ~n17467;
  assign n17470 = ~n17469 | ~n17468;
  assign n17473 = ~n17471 & ~n17470;
  assign n22755 = n24021 | n22789;
  assign n22713 = ~n22755;
  assign n17472 = ~n22713 | ~n23034;
  assign n17474 = ~n17473 | ~n17472;
  assign n17476 = ~n17475 & ~n17474;
  assign n17478 = ~n17477 | ~n17476;
  assign n17483 = ~n17479 & ~n17478;
  assign n23044 = n18007 ^ ~n18887;
  assign n17482 = ~n23044 | ~n22772;
  assign P1_U3280 = ~n17483 | ~n17482;
  assign n17484 = ~n25274 | ~n25389;
  assign n25244 = ~n25254 & ~n14816;
  assign n21061 = ~n25389;
  assign n17485 = n25274 | n21061;
  assign n17495 = n17502 | n17486;
  assign n17488 = ~n17487 | ~P2_IR_REG_31__SCAN_IN;
  assign n17491 = ~n17488 | ~P2_IR_REG_2__SCAN_IN;
  assign n17489 = ~P2_IR_REG_2__SCAN_IN;
  assign n17490 = ~n17489 | ~P2_IR_REG_31__SCAN_IN;
  assign n17493 = ~n17491 | ~n17490;
  assign n24586 = n17493 & n17492;
  assign n17496 = n17495 & n17494;
  assign n17500 = n17498 & n25399;
  assign n17499 = ~n25399 | ~n25252;
  assign n25175 = ~n17500;
  assign n17501 = ~n25217 | ~n25175;
  assign n17507 = n17948 | n17704;
  assign n17505 = n17502 | n17503;
  assign n17504 = ~n17657 | ~n24606;
  assign n17506 = n17505 & n17504;
  assign n25410 = ~n17507 | ~n17506;
  assign n25137 = n25410 | n25214;
  assign n25111 = ~n25410 | ~n25214;
  assign n25136 = n25137 & n25111;
  assign n17509 = ~P1_DATAO_REG_4__SCAN_IN;
  assign n17518 = n17502 | n17509;
  assign n17511 = ~n17510 | ~P2_IR_REG_31__SCAN_IN;
  assign n17514 = ~n17511 | ~P2_IR_REG_4__SCAN_IN;
  assign n17513 = ~n17512 | ~P2_IR_REG_31__SCAN_IN;
  assign n17516 = ~n17514 | ~n17513;
  assign n24627 = n17516 & n17515;
  assign n17517 = ~n17657 | ~n24627;
  assign n17519 = n25354 | n17704;
  assign n17792 = ~n25183 | ~n25420;
  assign n25142 = ~n25114 | ~n17792;
  assign n17530 = ~n25118 | ~n25142;
  assign n24482 = ~n25214;
  assign n25119 = n25410 & n24482;
  assign n17528 = ~n25119 | ~n25142;
  assign n17523 = n17502 | n17521;
  assign n17522 = ~n17657 | ~n24647;
  assign n17524 = n17523 & n17522;
  assign n17526 = n25104 | n25150;
  assign n17527 = n17526 & n25120;
  assign n17529 = n17528 & n17527;
  assign n17531 = ~n25104 | ~n25150;
  assign n17538 = n25348 | n17704;
  assign n17536 = n17502 | n17533;
  assign n17534 = n17597 | n17032;
  assign n24668 = n17534 ^ ~P2_IR_REG_6__SCAN_IN;
  assign n17535 = ~n17657 | ~n24668;
  assign n17537 = n17536 & n17535;
  assign n25090 = ~n17538 | ~n17537;
  assign n17793 = ~n25090 | ~n25126;
  assign n17539 = ~n25090 | ~n13779;
  assign n17547 = n25342 | n17704;
  assign n17540 = ~P1_DATAO_REG_7__SCAN_IN;
  assign n17545 = n17502 | n17540;
  assign n17541 = ~P2_IR_REG_6__SCAN_IN;
  assign n17542 = ~n17597 | ~n17541;
  assign n17543 = ~n17542 | ~P2_IR_REG_31__SCAN_IN;
  assign n24687 = n17543 ^ ~P2_IR_REG_7__SCAN_IN;
  assign n17544 = ~n17657 | ~n24687;
  assign n17546 = n17545 & n17544;
  assign n17548 = ~n25454 | ~n25093;
  assign n17549 = n25454 | n25093;
  assign n17561 = n25335 | n17704;
  assign n25336 = ~P1_DATAO_REG_8__SCAN_IN;
  assign n17559 = n21353 | n25336;
  assign n17551 = ~P2_IR_REG_6__SCAN_IN & ~P2_IR_REG_7__SCAN_IN;
  assign n17556 = ~n17597 | ~n17551;
  assign n17552 = ~n17556 | ~P2_IR_REG_31__SCAN_IN;
  assign n17555 = ~n17552 | ~P2_IR_REG_8__SCAN_IN;
  assign n17553 = ~P2_IR_REG_8__SCAN_IN;
  assign n17554 = ~n17553 | ~P2_IR_REG_31__SCAN_IN;
  assign n17557 = ~n17555 | ~n17554;
  assign n17558 = ~n17657 | ~n24707;
  assign n17560 = n17559 & n17558;
  assign n17800 = ~n25049;
  assign n17562 = ~n25467 | ~n17800;
  assign n17563 = n25467 | n17800;
  assign n17574 = n21353 | n17565;
  assign n17566 = ~n17569 | ~P2_IR_REG_31__SCAN_IN;
  assign n17568 = ~n17566 | ~P2_IR_REG_9__SCAN_IN;
  assign n17570 = ~P2_IR_REG_9__SCAN_IN;
  assign n17567 = ~n17570 | ~P2_IR_REG_31__SCAN_IN;
  assign n17572 = ~n17568 | ~n17567;
  assign n17571 = ~n17569;
  assign n17586 = ~n17571 | ~n17570;
  assign n24725 = n17572 & n17586;
  assign n17573 = ~n17657 | ~n24725;
  assign n17575 = n17574 & n17573;
  assign n24971 = ~n25021;
  assign n17576 = ~n25479 | ~n24971;
  assign n17577 = n25479 | n24971;
  assign n17583 = n25325 | n17704;
  assign n17581 = n17502 | n17578;
  assign n17579 = ~n17586 | ~P2_IR_REG_31__SCAN_IN;
  assign n24751 = n17579 ^ ~P2_IR_REG_10__SCAN_IN;
  assign n17580 = ~n17657 | ~n24751;
  assign n17582 = n17581 & n17580;
  assign n24434 = ~n25000;
  assign n17584 = ~n25489 | ~n24434;
  assign n17585 = n25489 | n24434;
  assign n17593 = n25320 | n17704;
  assign n17587 = n17586 | P2_IR_REG_10__SCAN_IN;
  assign n17588 = ~n17587 | ~P2_IR_REG_31__SCAN_IN;
  assign n24765 = n17588 ^ ~P2_IR_REG_11__SCAN_IN;
  assign n17591 = ~n24765 | ~n17657;
  assign n17590 = n21353 | n17589;
  assign n17592 = n17591 & n17590;
  assign n17805 = n25506 | n24976;
  assign n17806 = ~n25506 | ~n24976;
  assign n24349 = ~n24976;
  assign n17594 = ~n25506 | ~n24349;
  assign n17595 = ~P1_DATAO_REG_12__SCAN_IN;
  assign n17601 = n21353 | n17595;
  assign n17598 = ~n17596;
  assign n17605 = ~n17598 | ~n17597;
  assign n17599 = ~n17605 | ~P2_IR_REG_31__SCAN_IN;
  assign n24779 = n17599 ^ ~P2_IR_REG_12__SCAN_IN;
  assign n17600 = ~n17657 | ~n24779;
  assign n17602 = n17601 & n17600;
  assign n21415 = n24394 | n21845;
  assign n17604 = ~n21866 | ~n21415;
  assign n21414 = ~n24394 | ~n21845;
  assign n17610 = n25311 | n17704;
  assign n17608 = n17502 | n16051;
  assign n17606 = ~n17613 | ~P2_IR_REG_31__SCAN_IN;
  assign n24817 = n17606 ^ ~P2_IR_REG_13__SCAN_IN;
  assign n17607 = ~n17657 | ~n24817;
  assign n17609 = n17608 & n17607;
  assign n21431 = n24473 | n24389;
  assign n21430 = ~n24473 | ~n24389;
  assign n17612 = ~P1_DATAO_REG_14__SCAN_IN;
  assign n17619 = n21353 | n17612;
  assign n17615 = ~n17613;
  assign n17614 = ~P2_IR_REG_13__SCAN_IN;
  assign n17616 = ~n17615 | ~n17614;
  assign n17617 = ~n17616 | ~P2_IR_REG_31__SCAN_IN;
  assign n24832 = n17617 ^ ~P2_IR_REG_14__SCAN_IN;
  assign n17618 = ~n24832 | ~n17657;
  assign n17620 = n17619 & n17618;
  assign n24462 = ~n21413;
  assign n17622 = n22041 & n24462;
  assign n17623 = ~n21830 | ~n21413;
  assign n17627 = n21353 | n17625;
  assign n17626 = ~n17657 | ~n24863;
  assign n21035 = n17627 & n17626;
  assign n21760 = ~n21818;
  assign n17628 = ~n22029 | ~n21760;
  assign n21804 = ~n22029;
  assign n17629 = ~n21804 | ~n21818;
  assign n17630 = ~P1_DATAO_REG_16__SCAN_IN;
  assign n17639 = n21353 | n17630;
  assign n17633 = n17632 | n17032;
  assign n17636 = ~n17633 | ~P2_IR_REG_16__SCAN_IN;
  assign n17635 = ~n17634 | ~P2_IR_REG_31__SCAN_IN;
  assign n17637 = ~n17636 | ~n17635;
  assign n24886 = n17631 & n17637;
  assign n17638 = ~n17657 | ~n24886;
  assign n17640 = n17639 & n17638;
  assign n21791 = ~n21735;
  assign n17642 = ~n22018 | ~n21791;
  assign n17644 = ~n21755 | ~n17642;
  assign n17643 = n22018 | n21791;
  assign n21732 = ~n17644 | ~n17643;
  assign n17649 = n21353 | n25297;
  assign n17646 = ~n17631 | ~P2_IR_REG_31__SCAN_IN;
  assign n17645 = ~P2_IR_REG_17__SCAN_IN;
  assign n17655 = ~n17646 | ~n17645;
  assign n17647 = n17646 | n17645;
  assign n24903 = n17655 & n17647;
  assign n17648 = ~n17657 | ~n24903;
  assign n17650 = n17649 & n17648;
  assign n21759 = ~n21436;
  assign n17652 = ~n22008 | ~n21759;
  assign n17654 = ~n21732 | ~n17652;
  assign n17653 = n22008 | n21759;
  assign n21705 = ~n17654 | ~n17653;
  assign n17656 = ~n17655 | ~P2_IR_REG_31__SCAN_IN;
  assign n24928 = n17656 ^ ~P2_IR_REG_18__SCAN_IN;
  assign n17659 = ~n24928 | ~n17657;
  assign n17658 = n21353 | n25291;
  assign n17660 = n17659 & n17658;
  assign n17661 = ~n21997 | ~n13885;
  assign n17663 = ~n21705 | ~n17661;
  assign n17662 = n21997 | n13885;
  assign n17667 = n21353 | n17665;
  assign n17666 = n17029 | n24333;
  assign n17668 = n17667 & n17666;
  assign n17670 = ~n21356 | ~P2_REG2_REG_19__SCAN_IN;
  assign n17669 = ~n21359 | ~P2_REG0_REG_19__SCAN_IN;
  assign n17676 = ~n17670 | ~n17669;
  assign n17672 = ~n17685;
  assign n21695 = P2_REG3_REG_19__SCAN_IN ^ ~n17672;
  assign n17674 = ~n17780 | ~n21695;
  assign n17673 = ~n16780 | ~P2_REG1_REG_19__SCAN_IN;
  assign n17675 = ~n17674 | ~n17673;
  assign n21709 = ~n25556;
  assign n17677 = ~n21986 | ~n21709;
  assign n17681 = n21353 | n17680;
  assign n17684 = ~n16780 | ~P2_REG1_REG_20__SCAN_IN;
  assign n17683 = ~n21359 | ~P2_REG0_REG_20__SCAN_IN;
  assign n17690 = ~n17684 | ~n17683;
  assign n17686 = ~n17695;
  assign n21666 = P2_REG3_REG_20__SCAN_IN ^ ~n17686;
  assign n17688 = ~n17780 | ~n21666;
  assign n17687 = ~n21356 | ~P2_REG2_REG_20__SCAN_IN;
  assign n17689 = ~n17688 | ~n17687;
  assign n17693 = n21353 | n17692;
  assign n17696 = ~n17711;
  assign n21642 = P2_REG3_REG_21__SCAN_IN ^ ~n17696;
  assign n17698 = ~n17780 | ~n21642;
  assign n17697 = ~n21356 | ~P2_REG2_REG_21__SCAN_IN;
  assign n17702 = ~n17698 | ~n17697;
  assign n17700 = ~n16780 | ~P2_REG1_REG_21__SCAN_IN;
  assign n17699 = ~n21359 | ~P2_REG0_REG_21__SCAN_IN;
  assign n17701 = ~n17700 | ~n17699;
  assign n20948 = ~n25562;
  assign n21411 = n21965 & n20948;
  assign n17707 = n21353 | n17706;
  assign n17710 = ~n16780 | ~P2_REG1_REG_22__SCAN_IN;
  assign n17709 = ~n16781 | ~P2_REG0_REG_22__SCAN_IN;
  assign n17716 = ~n17710 | ~n17709;
  assign n17712 = ~n17722;
  assign n21621 = P2_REG3_REG_22__SCAN_IN ^ ~n17712;
  assign n17714 = ~n17780 | ~n21621;
  assign n17713 = ~n21356 | ~P2_REG2_REG_22__SCAN_IN;
  assign n17715 = ~n17714 | ~n17713;
  assign n17717 = ~n21954 | ~n21586;
  assign n17720 = ~n17718 | ~n13121;
  assign n17719 = ~n21363 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n17721 = ~n17720 | ~n17719;
  assign n17723 = ~n17737;
  assign n21599 = P2_REG3_REG_23__SCAN_IN ^ ~n17723;
  assign n17725 = ~n17780 | ~n21599;
  assign n17724 = ~n21356 | ~P2_REG2_REG_23__SCAN_IN;
  assign n17729 = ~n17725 | ~n17724;
  assign n17727 = ~n16780 | ~P2_REG1_REG_23__SCAN_IN;
  assign n17726 = ~n16781 | ~P2_REG0_REG_23__SCAN_IN;
  assign n17728 = ~n17727 | ~n17726;
  assign n17730 = ~n21598 | ~n25568;
  assign n17731 = n21598 | n25568;
  assign n17733 = n21353 | n18293;
  assign n17736 = ~n16780 | ~P2_REG1_REG_24__SCAN_IN;
  assign n17735 = ~n21359 | ~P2_REG0_REG_24__SCAN_IN;
  assign n17742 = ~n17736 | ~n17735;
  assign n17738 = ~n17746;
  assign n21572 = P2_REG3_REG_24__SCAN_IN ^ ~n17738;
  assign n17740 = ~n17780 | ~n21572;
  assign n17739 = ~n21356 | ~P2_REG2_REG_24__SCAN_IN;
  assign n17741 = ~n17740 | ~n17739;
  assign n21558 = n21932 ^ ~n25571;
  assign n21587 = ~n25571;
  assign n17743 = ~n21932 | ~n21587;
  assign n22166 = ~P1_DATAO_REG_25__SCAN_IN;
  assign n17744 = n21353 | n22166;
  assign n17747 = ~n17758;
  assign n21545 = P2_REG3_REG_25__SCAN_IN ^ ~n17747;
  assign n17749 = ~n17780 | ~n21545;
  assign n17748 = ~n16781 | ~P2_REG0_REG_25__SCAN_IN;
  assign n17753 = ~n17749 | ~n17748;
  assign n17751 = ~n21356 | ~P2_REG2_REG_25__SCAN_IN;
  assign n17750 = ~n16780 | ~P2_REG1_REG_25__SCAN_IN;
  assign n17752 = ~n17751 | ~n17750;
  assign n17754 = ~n21544 | ~n25574;
  assign n22158 = ~P1_DATAO_REG_26__SCAN_IN;
  assign n17755 = n21353 | n22158;
  assign n17757 = ~n21356 | ~P2_REG2_REG_26__SCAN_IN;
  assign n17756 = ~n21359 | ~P2_REG0_REG_26__SCAN_IN;
  assign n17763 = ~n17757 | ~n17756;
  assign n17759 = ~n17768;
  assign n21522 = P2_REG3_REG_26__SCAN_IN ^ ~n17759;
  assign n17761 = ~n17780 | ~n21522;
  assign n17760 = ~n16780 | ~P2_REG1_REG_26__SCAN_IN;
  assign n17762 = ~n17761 | ~n17760;
  assign n21410 = ~n21910 | ~n20881;
  assign n21508 = ~n21921 | ~n21560;
  assign n17764 = n21410 & n21508;
  assign n22151 = ~P1_DATAO_REG_27__SCAN_IN;
  assign n17765 = n21353 | n22151;
  assign n17767 = ~n16780 | ~P2_REG1_REG_27__SCAN_IN;
  assign n17766 = ~n16781 | ~P2_REG0_REG_27__SCAN_IN;
  assign n17772 = ~n17767 | ~n17766;
  assign n17777 = ~n17768 | ~P2_REG3_REG_26__SCAN_IN;
  assign n20807 = P2_REG3_REG_27__SCAN_IN ^ ~n17777;
  assign n17770 = ~n17780 | ~n20807;
  assign n17769 = ~n21356 | ~P2_REG2_REG_27__SCAN_IN;
  assign n17771 = ~n17770 | ~n17769;
  assign n17773 = ~n21323 | ~n19051;
  assign n17775 = ~n23137 | ~n21352;
  assign n22145 = ~P1_DATAO_REG_28__SCAN_IN;
  assign n17774 = n21353 | n22145;
  assign n17776 = ~P2_REG3_REG_27__SCAN_IN;
  assign n17778 = ~n17777 & ~n17776;
  assign n18126 = ~n17778 | ~P2_REG3_REG_28__SCAN_IN;
  assign n17779 = n17778 | P2_REG3_REG_28__SCAN_IN;
  assign n17786 = ~n21478 | ~n17780;
  assign n17782 = ~n16780 | ~P2_REG1_REG_28__SCAN_IN;
  assign n17781 = ~n16781 | ~P2_REG0_REG_28__SCAN_IN;
  assign n17784 = ~n17782 | ~n17781;
  assign n17783 = n21356 & P2_REG2_REG_28__SCAN_IN;
  assign n17785 = ~n17784 & ~n17783;
  assign n18084 = ~n21487 | ~n25583;
  assign n18113 = ~n17787 | ~n18084;
  assign n17789 = n18080 ^ ~n21444;
  assign n21394 = ~n21402 | ~n25194;
  assign n17788 = n21407 | n21456;
  assign n17848 = ~n17789 & ~n25270;
  assign n25218 = ~n25241 | ~n17790;
  assign n17791 = n25137 & n25135;
  assign n25040 = ~n25111 | ~n17792;
  assign n25043 = ~n25150 | ~n25432;
  assign n17794 = n17793 & n25043;
  assign n17796 = n25454 | n25022;
  assign n17797 = n17796 & n25045;
  assign n25052 = n25454 ^ ~n25093;
  assign n17798 = n25052 | n25093;
  assign n25029 = n25467 ^ ~n17800;
  assign n17801 = ~n25467 | ~n25049;
  assign n17802 = ~n25479 | ~n25021;
  assign n17803 = n25489 | n25000;
  assign n17804 = ~n25489 | ~n25000;
  assign n21880 = ~n24394;
  assign n17807 = ~n21880 | ~n21845;
  assign n17808 = ~n24394 | ~n24955;
  assign n17809 = n24473 | n21817;
  assign n17810 = ~n24473 | ~n21817;
  assign n17812 = ~n21830 | ~n24462;
  assign n17813 = ~n22041 | ~n21413;
  assign n17815 = ~n22029 | ~n21818;
  assign n21789 = ~n17816 | ~n17815;
  assign n21758 = n22018 ^ ~n21735;
  assign n17817 = n22008 | n21436;
  assign n17818 = ~n22008 | ~n21436;
  assign n17820 = n21997 | n21734;
  assign n21678 = ~n21986 | ~n25556;
  assign n17821 = n21975 | n25559;
  assign n17822 = ~n21975 | ~n25559;
  assign n20867 = ~n21965;
  assign n17823 = ~n20867 | ~n20948;
  assign n17824 = ~n21965 | ~n25562;
  assign n21617 = n21954 ^ ~n21586;
  assign n17825 = ~n21954 | ~n25565;
  assign n21561 = ~n25568;
  assign n17826 = ~n21598 | ~n21561;
  assign n21943 = ~n21598;
  assign n17827 = ~n21943 | ~n25568;
  assign n17829 = ~n21932 | ~n25571;
  assign n17830 = ~n21544 | ~n21560;
  assign n21517 = ~n21921 | ~n25574;
  assign n17831 = ~n21910 | ~n25577;
  assign n17832 = n21517 & n17831;
  assign n17833 = ~n21521 | ~n20881;
  assign n18118 = ~n21323 | ~n25580;
  assign n17835 = ~n17834 | ~n18118;
  assign n17849 = n17835 ^ ~n21444;
  assign n17836 = n21395 ^ ~n21402;
  assign n17846 = ~n17849 | ~n25248;
  assign n17842 = n18126 | n16777;
  assign n17838 = ~n16780 | ~P2_REG1_REG_29__SCAN_IN;
  assign n17837 = ~n21359 | ~P2_REG0_REG_29__SCAN_IN;
  assign n17840 = ~n17838 | ~n17837;
  assign n17839 = n21356 & P2_REG2_REG_29__SCAN_IN;
  assign n17841 = ~n17840 & ~n17839;
  assign n25586 = ~n17842 | ~n17841;
  assign n21340 = ~n25586;
  assign n17844 = ~n21340 & ~n25092;
  assign n17843 = ~n19051 & ~n25079;
  assign n17845 = ~n17844 & ~n17843;
  assign n17847 = ~n17846 | ~n17845;
  assign n21486 = ~n17849;
  assign n17858 = ~n21486 & ~n25509;
  assign n21722 = ~n21997;
  assign n17852 = ~n24394 & ~n25506;
  assign n25156 = ~n25410;
  assign n17850 = ~n25467 & ~n25454;
  assign n17851 = ~n25479 & ~n25489;
  assign n21829 = n21886 | n24473;
  assign n21802 = n22041 | n21829;
  assign n21771 = ~n22018;
  assign n21620 = ~n21954;
  assign n21497 = ~n21323;
  assign n17854 = ~n17853 | ~n21333;
  assign n17855 = ~n17854 | ~n25503;
  assign n25505 = ~n25441;
  assign n17856 = ~n21333 | ~n25505;
  assign n17857 = ~n21477 | ~n17856;
  assign n17859 = ~n17858 & ~n17857;
  assign n18147 = ~n21483 | ~n17859;
  assign n17865 = ~n18106;
  assign n17861 = ~n25373 | ~n17860;
  assign n18109 = ~n18145;
  assign n17867 = ~n18147 | ~n25553;
  assign n17866 = ~n25551 | ~P2_REG1_REG_28__SCAN_IN;
  assign P2_U3527 = ~n17867 | ~n17866;
  assign n17871 = ~n17872 | ~n25248;
  assign n18088 = ~n25583;
  assign n17869 = ~n18088 & ~n25092;
  assign n17868 = ~n20881 & ~n25079;
  assign n17870 = ~n17869 & ~n17868;
  assign n21495 = ~n17872;
  assign n17877 = ~n21495 & ~n25509;
  assign n21496 = n17873 ^ ~n21323;
  assign n17875 = ~n21496 | ~n25503;
  assign n17874 = ~n21323 | ~n25505;
  assign n17876 = ~n17875 | ~n17874;
  assign n17878 = ~n17877 & ~n17876;
  assign n17880 = ~n22076 | ~n25553;
  assign n17879 = ~n25551 | ~P2_REG1_REG_27__SCAN_IN;
  assign P2_U3526 = ~n17880 | ~n17879;
  assign n23532 = ~P1_ADDR_REG_10__SCAN_IN;
  assign n17883 = ~n23532 | ~P3_ADDR_REG_10__SCAN_IN;
  assign n17884 = ~P3_ADDR_REG_10__SCAN_IN;
  assign n17885 = ~n17884 | ~P1_ADDR_REG_10__SCAN_IN;
  assign n17895 = ~P3_ADDR_REG_11__SCAN_IN;
  assign n17887 = n17895 ^ ~P1_ADDR_REG_11__SCAN_IN;
  assign n17889 = n17894 ^ ~n17887;
  assign n17888 = ~P2_ADDR_REG_11__SCAN_IN;
  assign n17890 = ~n17889;
  assign n17900 = ~n17903;
  assign n17892 = ~P1_ADDR_REG_11__SCAN_IN;
  assign n17893 = ~n17892 | ~P3_ADDR_REG_11__SCAN_IN;
  assign n17896 = ~n17895 | ~P1_ADDR_REG_11__SCAN_IN;
  assign n17898 = P3_ADDR_REG_12__SCAN_IN ^ ~P1_ADDR_REG_12__SCAN_IN;
  assign n17902 = n17905 ^ ~n17898;
  assign n17901 = ~P2_ADDR_REG_12__SCAN_IN;
  assign n23574 = ~P1_ADDR_REG_12__SCAN_IN;
  assign n17904 = ~n23574 | ~P3_ADDR_REG_12__SCAN_IN;
  assign n17906 = ~P3_ADDR_REG_12__SCAN_IN;
  assign n17907 = ~n17906 | ~P1_ADDR_REG_12__SCAN_IN;
  assign n17916 = ~P3_ADDR_REG_13__SCAN_IN;
  assign n17908 = n17916 ^ ~P1_ADDR_REG_13__SCAN_IN;
  assign n17910 = n17915 ^ ~n17908;
  assign n17909 = ~P2_ADDR_REG_13__SCAN_IN;
  assign n17911 = ~n17910;
  assign n17921 = ~n17924;
  assign n17913 = ~P1_ADDR_REG_13__SCAN_IN;
  assign n17914 = ~n17913 | ~P3_ADDR_REG_13__SCAN_IN;
  assign n17917 = ~n17916 | ~P1_ADDR_REG_13__SCAN_IN;
  assign n17919 = P3_ADDR_REG_14__SCAN_IN ^ ~P1_ADDR_REG_14__SCAN_IN;
  assign n17923 = n17927 ^ ~n17919;
  assign n17920 = ~n17923;
  assign n17922 = ~P2_ADDR_REG_14__SCAN_IN;
  assign n23184 = ~n17924 | ~n17923;
  assign n23606 = ~P1_ADDR_REG_14__SCAN_IN;
  assign n17926 = ~P3_ADDR_REG_14__SCAN_IN & ~n23606;
  assign n17928 = ~n23606 | ~P3_ADDR_REG_14__SCAN_IN;
  assign n17929 = P1_ADDR_REG_15__SCAN_IN ^ ~P3_ADDR_REG_15__SCAN_IN;
  assign n17931 = n17934 ^ ~n17929;
  assign n17930 = ~P2_ADDR_REG_15__SCAN_IN;
  assign n17932 = ~n17931;
  assign n17935 = ~P3_ADDR_REG_15__SCAN_IN;
  assign n17933 = ~n17935 | ~P1_ADDR_REG_15__SCAN_IN;
  assign n17936 = P1_ADDR_REG_15__SCAN_IN | n17935;
  assign n17937 = ~P3_ADDR_REG_16__SCAN_IN;
  assign n17938 = n17937 ^ ~P1_ADDR_REG_16__SCAN_IN;
  assign n17939 = ~P2_ADDR_REG_16__SCAN_IN;
  assign n23645 = ~P1_ADDR_REG_16__SCAN_IN;
  assign n17943 = n23645 & P3_ADDR_REG_16__SCAN_IN;
  assign n17941 = ~P3_ADDR_REG_16__SCAN_IN & ~n23645;
  assign n17946 = ~P2_ADDR_REG_17__SCAN_IN;
  assign n17947 = n13355 | n17946;
  assign SUB_1596_U63 = ~n17947 | ~n19060;
  assign n17953 = ~n17948 & ~n24106;
  assign n17951 = n17949 | P1_U3086;
  assign n17950 = ~n24110 | ~P2_DATAO_REG_3__SCAN_IN;
  assign n17952 = ~n17951 | ~n17950;
  assign P1_U3352 = n17953 | n17952;
  assign n17957 = ~n21363 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n17956 = ~n13121 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n17958 = ~n17957 | ~n17956;
  assign n17959 = ~n17958 | ~SI_29_;
  assign n17973 = ~n17962 | ~n17959;
  assign n17960 = ~n17973;
  assign n17964 = ~n21363 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n17963 = ~n13121 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n17965 = ~n17964 | ~n17963;
  assign n17979 = n17965 ^ ~SI_30_;
  assign n17966 = ~n17965 | ~SI_30_;
  assign n17968 = ~n21363 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n17967 = ~n13121 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n17969 = ~n17968 | ~n17967;
  assign n17970 = n17969 ^ ~SI_31_;
  assign n17972 = ~n23114 | ~n14654;
  assign n23118 = ~P2_DATAO_REG_31__SCAN_IN;
  assign n17971 = n15451 | n23118;
  assign n22730 = ~n22753 | ~n23015;
  assign n17976 = ~n17974 | ~n17973;
  assign n17978 = ~n23130 | ~n14654;
  assign n19225 = ~P2_DATAO_REG_29__SCAN_IN;
  assign n17977 = n15451 | n19225;
  assign n23125 = ~P2_DATAO_REG_30__SCAN_IN;
  assign n17981 = n15451 | n23125;
  assign n17983 = ~n22422 | ~n22810;
  assign n17989 = ~n22414 & ~n24241;
  assign n17985 = ~n15251 | ~P1_REG2_REG_31__SCAN_IN;
  assign n17984 = ~n15669 | ~P1_REG1_REG_31__SCAN_IN;
  assign n17987 = n17985 & n17984;
  assign n17986 = ~n13129 | ~P1_REG0_REG_31__SCAN_IN;
  assign n18510 = n17987 & n17986;
  assign n24330 = ~n18510;
  assign n18910 = ~P1_B_REG_SCAN_IN;
  assign n17988 = ~n16818 & ~n18910;
  assign n19086 = ~n24014 & ~n17988;
  assign n22811 = n24330 & n19086;
  assign n17990 = ~n17989 & ~n22811;
  assign n23060 = ~n17991 | ~n17990;
  assign n17993 = ~n23060 | ~n24286;
  assign n17992 = ~n24284 | ~P1_REG1_REG_31__SCAN_IN;
  assign P1_U3559 = ~n17993 | ~n17992;
  assign n18005 = ~n18805 | ~n23331;
  assign n18003 = ~n22515 & ~n23329;
  assign n18001 = ~n22474 | ~n23343;
  assign n17999 = ~n23279 & ~n18062;
  assign n17998 = ~n17997 & ~P1_STATE_REG_SCAN_IN;
  assign n18000 = ~n17999 & ~n17998;
  assign n18002 = ~n18001 | ~n18000;
  assign n18004 = ~n18003 & ~n18002;
  assign n18864 = n19095 ^ ~n24320;
  assign n22953 = ~n24292;
  assign n22624 = ~n22223 | ~n22953;
  assign n18008 = n22341 | n22754;
  assign n18009 = ~n18041 | ~n22731;
  assign n18010 = ~n23015 | ~n23035;
  assign n18044 = ~n22998 | ~n22176;
  assign n18011 = n22998 | n22176;
  assign n18012 = ~n22998 | ~n23016;
  assign n18013 = ~n22702 | ~n22999;
  assign n22680 = ~n22999;
  assign n18014 = ~n22702 | ~n22680;
  assign n22706 = ~n22982;
  assign n18015 = n22295 | n22706;
  assign n22655 = n22664 ^ ~n24289;
  assign n18016 = ~n22952 | ~n24289;
  assign n18048 = n22223 | n24292;
  assign n18017 = ~n22223 | ~n24292;
  assign n22629 = ~n18048 | ~n18017;
  assign n18019 = ~n14515 | ~n24295;
  assign n18052 = ~n22889 | ~n22551;
  assign n18024 = ~n22889;
  assign n18023 = ~n18024 | ~n24301;
  assign n22585 = ~n18052 | ~n18023;
  assign n18025 = ~n18024 | ~n22551;
  assign n18027 = ~n22874 & ~n24304;
  assign n18028 = ~n18027;
  assign n18029 = ~n22535 & ~n24308;
  assign n18056 = n22862 | n24308;
  assign n18030 = ~n22862 | ~n24308;
  assign n22514 = ~n18056 | ~n18030;
  assign n18032 = ~n22514 & ~n18031;
  assign n22509 = ~n22491;
  assign n18034 = ~n22495 | ~n22515;
  assign n18035 = ~n22832 | ~n14111;
  assign n18036 = ~n18805 | ~n22847;
  assign n18037 = ~n22819 | ~n24316;
  assign n18038 = ~n22819 | ~n18062;
  assign n18066 = ~n18039 & ~n23991;
  assign n22771 = n18041 ^ ~n23035;
  assign n18042 = ~n22750;
  assign n18043 = ~n18041 | ~n23035;
  assign n18891 = ~n22295 | ~n22982;
  assign n18892 = n22295 | n22982;
  assign n18047 = ~n22664 | ~n24289;
  assign n18049 = ~n22618 | ~n24295;
  assign n18051 = ~n18050;
  assign n18053 = ~n18052;
  assign n18054 = ~n22874 | ~n22516;
  assign n18055 = ~n22544 | ~n14511;
  assign n18057 = ~n22495 | ~n24311;
  assign n18058 = ~n18805 | ~n14111;
  assign n18061 = ~n24012;
  assign n18065 = n18135 | n18061;
  assign n18064 = ~n18062 & ~n22789;
  assign n18063 = ~n18863 & ~n24014;
  assign n18068 = ~n18141 | ~n24019;
  assign n18067 = n24019 | P1_REG2_REG_28__SCAN_IN;
  assign n18079 = ~n18068 | ~n18067;
  assign n18077 = ~n18135 & ~n23892;
  assign n18136 = n18069 ^ ~n19095;
  assign n18075 = ~n18136 | ~n24026;
  assign n18073 = ~n19092 & ~n23980;
  assign n18071 = ~n18070;
  assign n18072 = ~n23936 & ~n18071;
  assign n18074 = ~n18073 & ~n18072;
  assign n18076 = ~n18075 | ~n18074;
  assign n18078 = ~n18077 & ~n18076;
  assign P1_U3265 = ~n18079 | ~n18078;
  assign n18087 = ~n18080 | ~n21444;
  assign n18082 = ~n23130 | ~n21352;
  assign n22140 = ~P1_DATAO_REG_29__SCAN_IN;
  assign n18081 = n21353 | n22140;
  assign n21447 = n21345 ^ ~n21340;
  assign n18083 = ~n21447 | ~n25246;
  assign n18104 = ~n18087 & ~n18083;
  assign n18085 = ~n18084 | ~n25246;
  assign n18086 = ~n21447 & ~n18085;
  assign n18102 = ~n18087 | ~n18086;
  assign n18123 = ~n21447;
  assign n18089 = ~n18088 & ~n25270;
  assign n18090 = ~n21487 | ~n18089;
  assign n18100 = ~n18123 & ~n18090;
  assign n18098 = ~n25583 | ~n25253;
  assign n18091 = ~P2_B_REG_SCAN_IN;
  assign n18092 = ~n24516 & ~n18091;
  assign n21463 = ~n25092 & ~n18092;
  assign n18094 = ~n16780 | ~P2_REG1_REG_30__SCAN_IN;
  assign n18093 = ~n21356 | ~P2_REG2_REG_30__SCAN_IN;
  assign n18096 = ~n18094 | ~n18093;
  assign n18095 = n16781 & P2_REG0_REG_30__SCAN_IN;
  assign n25589 = n18096 | n18095;
  assign n18097 = ~n21463 | ~n25589;
  assign n18099 = ~n18098 | ~n18097;
  assign n18101 = ~n18100 & ~n18099;
  assign n18103 = ~n18102 | ~n18101;
  assign n18154 = ~n18104 & ~n18103;
  assign n18107 = ~n18105;
  assign n18108 = n18107 & n18106;
  assign n18110 = ~n18109 | ~n18108;
  assign n18112 = ~n18154 | ~n25284;
  assign n18111 = n25284 | P2_REG2_REG_29__SCAN_IN;
  assign n18134 = ~n18112 | ~n18111;
  assign n18117 = ~n21333 | ~n25583;
  assign n18114 = ~n18117;
  assign n18116 = n18114 | n18113;
  assign n18115 = n21445 & n18116;
  assign n18120 = ~n18116;
  assign n18119 = n18118 & n18117;
  assign n18124 = ~n25284 | ~n25248;
  assign n18132 = ~n18150 & ~n21828;
  assign n18151 = n21460 ^ ~n21345;
  assign n21803 = ~n25282 & ~n24449;
  assign n18130 = ~n18151 | ~n25263;
  assign n21459 = ~n21345;
  assign n25189 = ~n25091;
  assign n18128 = ~n21459 & ~n25105;
  assign n18127 = ~n18126 & ~n25267;
  assign n18129 = ~n18128 & ~n18127;
  assign n18131 = ~n18130 | ~n18129;
  assign n18133 = ~n18132 & ~n18131;
  assign P2_U3236 = ~n18134 | ~n18133;
  assign n18140 = ~n18135 & ~n24220;
  assign n18138 = ~n18136 | ~n24216;
  assign n18137 = ~n19095 | ~n24230;
  assign n18139 = ~n18138 | ~n18137;
  assign n18142 = ~n18140 & ~n18139;
  assign n18143 = ~n24284 | ~P1_REG1_REG_28__SCAN_IN;
  assign P1_U3556 = ~n18144 | ~n18143;
  assign n25488 = n18146 | n18145;
  assign n18149 = ~n18147 | ~n25515;
  assign n18148 = ~n25488 | ~P2_REG0_REG_28__SCAN_IN;
  assign P2_U3495 = ~n18149 | ~n18148;
  assign n25477 = ~n25509;
  assign n22038 = ~n25248 & ~n25477;
  assign n18153 = ~n18151 | ~n25503;
  assign n18152 = ~n21345 | ~n25505;
  assign n18156 = ~n18477 | ~n25515;
  assign n18155 = ~n25488 | ~P2_REG0_REG_29__SCAN_IN;
  assign P2_U3496 = ~n18156 | ~n18155;
  assign n18157 = ~n19335;
  assign n18402 = ~n19334;
  assign n26232 = ~n18158 | ~n26245;
  assign n19322 = ~n19315;
  assign n19274 = ~n26287 | ~n26316;
  assign n25707 = ~n26245;
  assign n19329 = ~n26286 | ~n26245;
  assign n25626 = ~n26335;
  assign n18160 = ~n26252 | ~n25626;
  assign n25624 = ~n26229;
  assign n19340 = ~n26229 | ~n26343;
  assign n18162 = ~n26229 | ~n26212;
  assign n25723 = ~n26205;
  assign n18164 = n18176 | SI_5_;
  assign n18163 = n18258 | n25850;
  assign n18167 = ~n18164 | ~n18163;
  assign n18166 = ~n19228 & ~n18165;
  assign n19345 = ~n25723 | ~n26174;
  assign n26181 = ~n19345 | ~n19346;
  assign n26183 = ~n26181;
  assign n18227 = ~n19228;
  assign n18173 = n18227 & n18168;
  assign n18171 = n18176 | n18169;
  assign n18170 = n18258 | n25875;
  assign n18172 = ~n18171 | ~n18170;
  assign n18405 = ~n26138 | ~n26150;
  assign n26160 = ~n18405 | ~n14876;
  assign n19357 = ~n26189 | ~n26150;
  assign n26127 = ~n18174 | ~n19357;
  assign n18180 = n18175 | n19228;
  assign n18178 = n18176 | SI_7_;
  assign n18177 = n18258 | n25893;
  assign n18179 = n18178 & n18177;
  assign n26367 = ~n18180 | ~n18179;
  assign n26106 = n19134 ^ ~n26367;
  assign n25597 = ~n26367;
  assign n18181 = ~n25597 | ~n26165;
  assign n18187 = n18182 | n18351;
  assign n18185 = n18176 | n18183;
  assign n18184 = n18258 | n25916;
  assign n18186 = n18185 & n18184;
  assign n19360 = ~n18187 | ~n18186;
  assign n26375 = ~n19360;
  assign n19371 = ~n26375 & ~n26125;
  assign n19363 = ~n26375 | ~n26125;
  assign n18188 = ~n19363;
  assign n18195 = n18190 | n18351;
  assign n18193 = n18176 | SI_9_;
  assign n18192 = n18258 | n19984;
  assign n18194 = n18193 & n18192;
  assign n18200 = n18196 | n18351;
  assign n18198 = n18176 | SI_10_;
  assign n18197 = n18258 | n19987;
  assign n18199 = n18198 & n18197;
  assign n18201 = ~n26393 | ~n25689;
  assign n18207 = n18203 | n19228;
  assign n18205 = n18176 | SI_11_;
  assign n18204 = n18258 | n19989;
  assign n18206 = n18205 & n18204;
  assign n20681 = ~n18207 | ~n18206;
  assign n18413 = ~n20681 | ~n25611;
  assign n18414 = n20681 | n25611;
  assign n18209 = ~n13122 | ~SI_12_;
  assign n18210 = n18258 | n25988;
  assign n20507 = ~n18211 | ~n18210;
  assign n18418 = n20507 | n25692;
  assign n18417 = ~n20507 | ~n25692;
  assign n18214 = n18176 | SI_13_;
  assign n18213 = n18258 | n19993;
  assign n18215 = n18214 & n18213;
  assign n18217 = ~n20665 | ~n20495;
  assign n20484 = ~n20665;
  assign n18218 = ~n20484 | ~n19552;
  assign n18221 = n18176 | SI_14_;
  assign n18220 = n18258 | n19997;
  assign n18222 = n18221 & n18220;
  assign n18226 = ~n20452 | ~n14570;
  assign n18224 = ~n20656;
  assign n18225 = ~n18224 | ~n19406;
  assign n18232 = ~n18228 | ~n18227;
  assign n18230 = n18176 | SI_15_;
  assign n18229 = n19999 | n18258;
  assign n18231 = n18230 & n18229;
  assign n18233 = ~n20648 | ~n20454;
  assign n19415 = ~n20648;
  assign n18234 = ~n19415 | ~n19646;
  assign n18237 = ~n18236;
  assign n18242 = ~n18237 | ~n18227;
  assign n18240 = ~n20034 | ~n17198;
  assign n18239 = n18176 | n18238;
  assign n18241 = n18240 & n18239;
  assign n20424 = n19413 ^ ~n19795;
  assign n19287 = ~n20424;
  assign n19424 = ~n19413 | ~n19795;
  assign n18245 = ~n20094 | ~n17198;
  assign n18244 = n18176 | SI_17_;
  assign n18246 = n18245 & n18244;
  assign n20406 = n20632 ^ ~n20416;
  assign n18251 = n18176 | n18249;
  assign n18250 = n18258 | n20106;
  assign n18252 = n18251 & n18250;
  assign n19430 = n19427 & n19674;
  assign n18254 = ~n19430;
  assign n18260 = n18176 | n18257;
  assign n18259 = n18258 | n20119;
  assign n18261 = n18260 & n18259;
  assign n19453 = ~n20369 & ~n19446;
  assign n18262 = ~n19453;
  assign n20280 = ~n20369 | ~n19446;
  assign n18265 = n18263 | n13121;
  assign n18264 = ~n13121 | ~SI_22_;
  assign n18266 = ~n18265 | ~n18264;
  assign n18280 = ~n20593 | ~n20310;
  assign n18275 = ~n18280;
  assign n18269 = n18176 | n18268;
  assign n20306 = ~n20349 | ~n19602;
  assign n18272 = n18176 | n18271;
  assign n18274 = ~n18431 | ~n19752;
  assign n20283 = ~n14883 | ~n14881;
  assign n18276 = n20280 & n18279;
  assign n20298 = ~n20593;
  assign n18278 = ~n20298 | ~n20267;
  assign n18277 = n18276 & n18278;
  assign n20254 = ~n20281 | ~n18277;
  assign n18284 = ~n18278;
  assign n18282 = ~n18279;
  assign n18281 = n20282 & n18280;
  assign n20253 = n18284 | n18283;
  assign n18286 = ~SI_23_;
  assign n18287 = n18176 | n18286;
  assign n19568 = ~n20585;
  assign n19466 = ~n19568 | ~n19692;
  assign n20287 = ~n19692;
  assign n19467 = ~n20585 | ~n20287;
  assign n20263 = ~n19466 | ~n19467;
  assign n20228 = n20253 & n20263;
  assign n18290 = ~n18289;
  assign n18295 = ~n18292 | ~P2_DATAO_REG_23__SCAN_IN;
  assign n18294 = ~n18297 | ~n18295;
  assign n18308 = ~n18294 | ~n18293;
  assign n18296 = n18295 & P1_DATAO_REG_24__SCAN_IN;
  assign n18298 = ~n18308 | ~n18306;
  assign n18299 = n18298 ^ ~P2_DATAO_REG_24__SCAN_IN;
  assign n18300 = ~n13122 | ~SI_24_;
  assign n20210 = ~n20266;
  assign n18303 = ~n18436 | ~n20210;
  assign n18305 = ~n20254 | ~n18302;
  assign n18304 = ~n18303;
  assign n20229 = ~n20585 | ~n19692;
  assign n18319 = ~n18308 | ~n18307;
  assign n18318 = n22166 ^ ~P2_DATAO_REG_25__SCAN_IN;
  assign n20793 = n18319 ^ ~n18318;
  assign n20795 = ~SI_25_;
  assign n18309 = n18176 | n20795;
  assign n20221 = n18323 ^ ~P3_REG3_REG_25__SCAN_IN;
  assign n18316 = ~n20221 | ~n16484;
  assign n18312 = ~n16422 | ~P3_REG2_REG_25__SCAN_IN;
  assign n18311 = ~n18368 | ~P3_REG1_REG_25__SCAN_IN;
  assign n18314 = ~n18312 | ~n18311;
  assign n18313 = n18340 & P3_REG0_REG_25__SCAN_IN;
  assign n18315 = ~n18314 & ~n18313;
  assign n19480 = ~n20220 | ~n20235;
  assign n18317 = ~n20220 | ~n26436;
  assign n18320 = ~n23159 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n18334 = P1_DATAO_REG_26__SCAN_IN ^ ~P2_DATAO_REG_26__SCAN_IN;
  assign n20785 = n18335 ^ ~n18334;
  assign n20787 = ~SI_26_;
  assign n20198 = P3_REG3_REG_26__SCAN_IN ^ ~n18339;
  assign n18330 = ~n20198 | ~n16484;
  assign n18325 = ~n18368 | ~P3_REG1_REG_26__SCAN_IN;
  assign n18324 = ~n18380 | ~P3_REG0_REG_26__SCAN_IN;
  assign n18328 = ~n18325 | ~n18324;
  assign n20193 = ~P3_REG2_REG_26__SCAN_IN;
  assign n18327 = ~n18326 & ~n20193;
  assign n18329 = ~n18328 & ~n18327;
  assign n18331 = ~n20560 | ~n20209;
  assign n18332 = ~n20197 | ~n26439;
  assign n18336 = ~n23151 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n18347 = P1_DATAO_REG_27__SCAN_IN ^ ~P2_DATAO_REG_27__SCAN_IN;
  assign n20780 = ~SI_27_;
  assign n18338 = n18176 | n20780;
  assign n20175 = n18355 ^ ~P3_REG3_REG_27__SCAN_IN;
  assign n18346 = ~n20175 | ~n16484;
  assign n18342 = ~n16422 | ~P3_REG2_REG_27__SCAN_IN;
  assign n18341 = ~n18340 | ~P3_REG0_REG_27__SCAN_IN;
  assign n18344 = ~n18342 | ~n18341;
  assign n18343 = n18368 & P3_REG1_REG_27__SCAN_IN;
  assign n18345 = ~n18344 & ~n18343;
  assign n18350 = ~n18348 | ~n18347;
  assign n18349 = ~n23144 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n18360 = P1_DATAO_REG_28__SCAN_IN ^ ~P2_DATAO_REG_28__SCAN_IN;
  assign n18352 = ~SI_28_;
  assign n18353 = n18176 | n18352;
  assign n18356 = ~n16484 | ~n20152;
  assign n18358 = ~n16463 | ~P3_REG1_REG_28__SCAN_IN;
  assign n18357 = ~n18380 | ~P3_REG0_REG_28__SCAN_IN;
  assign n18359 = ~n18358 | ~n18357;
  assign n18362 = ~n18361 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n19223 = P1_DATAO_REG_29__SCAN_IN ^ ~P2_DATAO_REG_29__SCAN_IN;
  assign n20765 = n19224 ^ ~n19223;
  assign n20767 = ~SI_29_;
  assign n18364 = n18176 | n20767;
  assign n18367 = ~n16460 | ~P3_REG2_REG_29__SCAN_IN;
  assign n19231 = ~n16484 | ~n18492;
  assign n18372 = ~n18367 | ~n19231;
  assign n18370 = ~n18368 | ~P3_REG1_REG_29__SCAN_IN;
  assign n18369 = ~n18380 | ~P3_REG0_REG_29__SCAN_IN;
  assign n18371 = ~n18370 | ~n18369;
  assign n19499 = n19503 ^ ~n26448;
  assign n18374 = ~n14256 & ~n20165;
  assign n18373 = ~n18454;
  assign n19252 = n19522 | n19306;
  assign n18375 = ~n18374 & ~n26129;
  assign n18376 = ~n19295 | ~n18375;
  assign n18377 = ~n26445 | ~n26280;
  assign n18378 = ~n14256 & ~n18377;
  assign n18391 = ~n19499 | ~n18378;
  assign n18379 = ~n16422 | ~P3_REG2_REG_30__SCAN_IN;
  assign n18384 = ~n18379 | ~n19231;
  assign n18382 = ~n18368 | ~P3_REG1_REG_30__SCAN_IN;
  assign n18381 = ~n18380 | ~P3_REG0_REG_30__SCAN_IN;
  assign n18383 = ~n18382 | ~n18381;
  assign n19509 = ~n26451;
  assign n19520 = n19364;
  assign n19950 = ~n20773;
  assign n18386 = ~n19950 | ~P3_B_REG_SCAN_IN;
  assign n20130 = ~n18385 | ~n18386;
  assign n18389 = ~n19509 & ~n20130;
  assign n18388 = ~n20165 & ~n26137;
  assign n18390 = ~n18389 & ~n18388;
  assign n18392 = ~n18391 | ~n18390;
  assign n18396 = ~n18393 & ~n18392;
  assign n18394 = ~n19295 & ~n26129;
  assign n18395 = ~n20144 | ~n18394;
  assign n18488 = ~n18396 | ~n18395;
  assign n18397 = ~n19501 & ~n20673;
  assign n18447 = ~n18488 & ~n18397;
  assign n19309 = ~n26273;
  assign n18398 = ~n19309 | ~n19273;
  assign n26248 = ~n18398 | ~n19321;
  assign n18400 = ~n26248 | ~n18399;
  assign n18401 = ~n26233;
  assign n18403 = ~n26227 | ~n18401;
  assign n18404 = ~n26198 | ~n14555;
  assign n26074 = ~n18406 | ~n18405;
  assign n26111 = n19360 ^ ~n26086;
  assign n26075 = n26106 & n26111;
  assign n19373 = ~n26383 | ~n26116;
  assign n18407 = n26075 & n19373;
  assign n18412 = ~n26074 | ~n18407;
  assign n18409 = ~n19373;
  assign n26107 = ~n19134 | ~n25597;
  assign n18408 = ~n19360 | ~n26125;
  assign n19372 = n26383 | n26116;
  assign n19388 = ~n26393 & ~n26085;
  assign n19379 = ~n20681 & ~n26059;
  assign n18415 = ~n19379;
  assign n20493 = ~n18418 | ~n18417;
  assign n19397 = ~n20507 | ~n20517;
  assign n19401 = ~n20665 | ~n19552;
  assign n19400 = ~n20484 | ~n20495;
  assign n19405 = n20656 | n19406;
  assign n20442 = n20648 ^ ~n20454;
  assign n19417 = ~n20648 & ~n19646;
  assign n18420 = ~n19417;
  assign n20435 = ~n19795;
  assign n18422 = ~n19413 | ~n20435;
  assign n19442 = ~n20632 & ~n19771;
  assign n18423 = ~n19442;
  assign n18426 = n19427 | n20398;
  assign n18427 = ~n20363;
  assign n18428 = ~n20369 | ~n20376;
  assign n19459 = ~n18431 & ~n20334;
  assign n18429 = ~n19459;
  assign n19456 = ~n20349 & ~n20354;
  assign n20315 = ~n19456;
  assign n20258 = n18429 & n20315;
  assign n20260 = ~n20593 | ~n20267;
  assign n19462 = ~n20260;
  assign n18430 = n20258 & n20260;
  assign n19461 = ~n20261;
  assign n18433 = n20263 | n19461;
  assign n20259 = ~n19460;
  assign n18432 = ~n20259 & ~n19462;
  assign n18434 = ~n18433 & ~n18432;
  assign n18435 = ~n19466;
  assign n19271 = ~n20245 & ~n20210;
  assign n19473 = ~n19271;
  assign n19270 = ~n18436 & ~n20266;
  assign n19472 = ~n19270;
  assign n18438 = ~n20560 | ~n26439;
  assign n18439 = ~n20197 | ~n20209;
  assign n18440 = ~n20552 | ~n26442;
  assign n18441 = ~n20174 | ~n20186;
  assign n18442 = ~n18455 | ~n20673;
  assign n18445 = n18465 | n18442;
  assign n18444 = n19257 | n18443;
  assign n18452 = n18444 | n18455;
  assign n20684 = ~n20501 | ~n26391;
  assign n18446 = ~n18495 | ~n20684;
  assign n18451 = n18448 ^ ~n18482;
  assign n18450 = n18449 & n18473;
  assign n18481 = ~n18452 | ~n19520;
  assign n18480 = n18481 & n18453;
  assign n18461 = ~n18480 | ~n18482;
  assign n18479 = ~n18482;
  assign n18456 = n18455 | n18454;
  assign n18458 = ~n18456 | ~n19306;
  assign n18459 = ~n18458 | ~n18457;
  assign n18460 = ~n18479 | ~n18459;
  assign n18462 = ~n18461 | ~n18460;
  assign n18463 = ~n26431 | ~P3_REG1_REG_29__SCAN_IN;
  assign P3_U3488 = ~n18464 | ~n18463;
  assign n18466 = ~n18465;
  assign n18472 = ~n18467 | ~n18466;
  assign n18469 = n26303 | n18468;
  assign n18471 = ~n18470 | ~n18469;
  assign n18474 = ~n18472 | ~n18471;
  assign n18475 = ~n26390 | ~P3_REG0_REG_29__SCAN_IN;
  assign P3_U3456 = ~n18476 | ~n18475;
  assign n18478 = ~n25551 | ~P2_REG1_REG_29__SCAN_IN;
  assign n18485 = ~n18480 | ~n18479;
  assign n18483 = ~n18481;
  assign n18484 = ~n18483 | ~n18482;
  assign n18486 = ~n18485 | ~n18484;
  assign n18489 = ~n18487 | ~n18486;
  assign n18491 = ~n18489;
  assign n18490 = n26278 & n26315;
  assign n18493 = ~n19501 & ~n26224;
  assign n20131 = n26152 & n18492;
  assign n18494 = ~n18493 & ~n20131;
  assign n26249 = n26278 | n19306;
  assign n20388 = ~n20501 | ~n26249;
  assign n18496 = ~n18495 | ~n20526;
  assign n18499 = ~n18497 | ~n24251;
  assign n18498 = ~n24240 | ~P1_REG0_REG_28__SCAN_IN;
  assign P1_U3524 = ~n18499 | ~n18498;
  assign n18500 = ~n18854 | ~n23723;
  assign n18506 = n18501 & n18500;
  assign n18502 = ~n18506 | ~n18861;
  assign n18511 = n18502 & n18547;
  assign n18507 = ~n18506;
  assign n18503 = ~n18507 | ~n18860;
  assign n18505 = ~n22414 & ~n18563;
  assign n18504 = ~n18843 & ~n18510;
  assign n18509 = ~n18505 & ~n18504;
  assign n18508 = ~n18506 | ~n18860;
  assign n18522 = ~n18507 | ~n18861;
  assign n18521 = n18735 & n24330;
  assign n18849 = ~n18509 & ~n18521;
  assign n18735 = ~n18779;
  assign n18520 = ~n22421 | ~n18735;
  assign n18517 = ~n18511 | ~n18510;
  assign n18516 = n18512 & P1_REG0_REG_30__SCAN_IN;
  assign n18514 = ~n15251 | ~P1_REG2_REG_30__SCAN_IN;
  assign n18513 = ~n15936 | ~P1_REG1_REG_30__SCAN_IN;
  assign n18515 = ~n18514 | ~n18513;
  assign n24327 = n18516 | n18515;
  assign n18518 = n18517 & n24327;
  assign n18519 = ~n18518 | ~n18563;
  assign n18845 = n18520 & n18519;
  assign n18526 = ~n22421 | ~n18563;
  assign n18523 = ~n18521;
  assign n18524 = ~n18523 | ~n18522;
  assign n18525 = ~n18524 | ~n24327;
  assign n18844 = ~n18526 | ~n18525;
  assign n18532 = ~n18845 | ~n18844;
  assign n18528 = ~n19085 | ~n18735;
  assign n24323 = ~n18863;
  assign n18527 = ~n18563 | ~n24323;
  assign n18836 = n18528 & n18527;
  assign n18530 = ~n19085 | ~n18563;
  assign n18529 = ~n24323 | ~n18735;
  assign n18835 = ~n18530 | ~n18529;
  assign n18531 = ~n18836 | ~n18835;
  assign n18533 = ~n18532 | ~n18531;
  assign n18842 = ~n18849 & ~n18533;
  assign n18534 = ~n18829 | ~n24298;
  assign n18763 = n18535 & n18534;
  assign n18536 = ~n18563 | ~n24298;
  assign n18762 = ~n18537 | ~n18536;
  assign n18761 = ~n18763 | ~n18762;
  assign n18539 = ~n22618 | ~n18563;
  assign n18538 = ~n24295 | ~n18735;
  assign n18757 = n18539 & n18538;
  assign n18541 = ~n22618 | ~n18735;
  assign n18540 = ~n24295 | ~n18563;
  assign n18756 = ~n18541 | ~n18540;
  assign n18755 = ~n18757 | ~n18756;
  assign n18543 = ~n18563 | ~n17352;
  assign n18542 = ~n18829 | ~n17382;
  assign n18559 = n18543 & n18542;
  assign n18552 = ~n18559 | ~n17352;
  assign n18546 = ~n18544 | ~n18545;
  assign n18548 = ~n23993 | ~n18547;
  assign n18550 = ~n18549 | ~n18735;
  assign n18558 = ~n18552 | ~n18551;
  assign n18554 = ~n18563 | ~n17382;
  assign n18553 = ~n18829 | ~n17352;
  assign n18556 = n18554 & n18553;
  assign n18555 = ~n18559;
  assign n18557 = ~n18556 | ~n18555;
  assign n18561 = ~n18558 | ~n18557;
  assign n18560 = ~n18559 | ~n17382;
  assign n18562 = ~n18563 | ~n23254;
  assign n18569 = ~n18829 | ~n23967;
  assign n18566 = n18562 & n18569;
  assign n18565 = ~n18563 | ~n23967;
  assign n18564 = ~n18829 | ~n23254;
  assign n18568 = ~n18565 | ~n18564;
  assign n18567 = ~n18566 | ~n18568;
  assign n18571 = ~n18568;
  assign n18570 = ~n18569 | ~n24000;
  assign n18572 = ~n18571 | ~n18570;
  assign n18574 = ~n18563 | ~n14281;
  assign n18573 = ~n18735 | ~n17357;
  assign n18581 = ~n14281 | ~n18735;
  assign n18576 = n18581 & n18575;
  assign n18578 = ~n18563 | ~n23874;
  assign n18577 = ~n18829 | ~n23903;
  assign n18593 = n18578 & n18577;
  assign n18580 = ~n18563 | ~n23903;
  assign n18579 = ~n18829 | ~n23874;
  assign n18592 = ~n18580 | ~n18579;
  assign n18586 = ~n18593 | ~n18592;
  assign n18582 = ~n18563 | ~n17357;
  assign n18584 = n18582 & n18581;
  assign n18585 = ~n18584 | ~n18583;
  assign n18587 = n18586 & n18585;
  assign n18589 = ~n18563 | ~n14266;
  assign n18588 = ~n18829 | ~n23854;
  assign n18605 = n18589 & n18588;
  assign n18591 = ~n18563 | ~n23854;
  assign n18590 = ~n18829 | ~n14266;
  assign n18604 = ~n18591 | ~n18590;
  assign n18597 = ~n18605 | ~n18604;
  assign n18595 = ~n18592;
  assign n18594 = ~n18593;
  assign n18596 = ~n18595 | ~n18594;
  assign n18598 = n18597 & n18596;
  assign n18611 = ~n18599 | ~n18598;
  assign n18601 = ~n18563 | ~n23875;
  assign n18600 = ~n24190 | ~n18735;
  assign n18616 = n18601 & n18600;
  assign n18603 = ~n18563 | ~n24190;
  assign n18602 = ~n18829 | ~n23875;
  assign n18615 = ~n18603 | ~n18602;
  assign n18609 = ~n18616 | ~n18615;
  assign n18607 = ~n18604;
  assign n18606 = ~n18605;
  assign n18608 = ~n18607 | ~n18606;
  assign n18610 = n18609 & n18608;
  assign n18612 = ~n23818 | ~n18563;
  assign n18614 = ~n23818 | ~n18735;
  assign n18613 = ~n18563 | ~n23853;
  assign n18625 = ~n18614 | ~n18613;
  assign n18620 = ~n18626 | ~n18625;
  assign n18618 = ~n18615;
  assign n18617 = ~n18616;
  assign n18619 = ~n18618 | ~n18617;
  assign n18622 = ~n24213 | ~n18735;
  assign n18621 = ~n18563 | ~n23825;
  assign n18637 = n18622 & n18621;
  assign n18624 = ~n24213 | ~n18563;
  assign n18623 = ~n18735 | ~n23825;
  assign n18636 = ~n18624 | ~n18623;
  assign n18630 = ~n18637 | ~n18636;
  assign n18628 = ~n18625;
  assign n18629 = ~n18628 | ~n18627;
  assign n18631 = n18630 & n18629;
  assign n18633 = ~n24231 | ~n18563;
  assign n18632 = ~n18829 | ~n23801;
  assign n18644 = n18633 & n18632;
  assign n18635 = ~n24231 | ~n18735;
  assign n18634 = ~n18563 | ~n23801;
  assign n18643 = ~n18635 | ~n18634;
  assign n18641 = ~n18644 | ~n18643;
  assign n18639 = ~n18636;
  assign n18638 = ~n18637;
  assign n18640 = ~n18639 | ~n18638;
  assign n18642 = n18641 & n18640;
  assign n18646 = ~n18643;
  assign n18645 = ~n18644;
  assign n18653 = ~n18646 | ~n18645;
  assign n18648 = ~n18649 | ~n18735;
  assign n18647 = ~n18563 | ~n23769;
  assign n18660 = n18648 & n18647;
  assign n18651 = ~n18649 | ~n18563;
  assign n18650 = ~n18735 | ~n23769;
  assign n18659 = ~n18651 | ~n18650;
  assign n18652 = ~n18660 | ~n18659;
  assign n18654 = n18653 & n18652;
  assign n18656 = ~n23051 | ~n18563;
  assign n18655 = ~n18829 | ~n23753;
  assign n18672 = n18656 & n18655;
  assign n18658 = ~n23051 | ~n18829;
  assign n18657 = ~n18563 | ~n23753;
  assign n18671 = ~n18658 | ~n18657;
  assign n18664 = ~n18672 | ~n18671;
  assign n18662 = ~n18659;
  assign n18661 = ~n18660;
  assign n18663 = ~n18662 | ~n18661;
  assign n18665 = n18664 & n18663;
  assign n18668 = ~n18666 | ~n18829;
  assign n18667 = ~n18563 | ~n23034;
  assign n18682 = n18668 & n18667;
  assign n18670 = ~n22257 & ~n13123;
  assign n18669 = ~n18779 & ~n22790;
  assign n18681 = n18670 | n18669;
  assign n18676 = ~n18682 | ~n18681;
  assign n18674 = ~n18671;
  assign n18673 = ~n18672;
  assign n18675 = ~n18674 | ~n18673;
  assign n18678 = ~n22341 | ~n18563;
  assign n18677 = ~n18829 | ~n23017;
  assign n18689 = n18678 & n18677;
  assign n18680 = ~n22341 | ~n18829;
  assign n18679 = ~n18563 | ~n23017;
  assign n18688 = ~n18680 | ~n18679;
  assign n18686 = ~n18689 | ~n18688;
  assign n18684 = ~n18681;
  assign n18683 = ~n18682;
  assign n18685 = ~n18684 | ~n18683;
  assign n18687 = n18686 & n18685;
  assign n18691 = ~n18688;
  assign n18690 = ~n18689;
  assign n18692 = ~n18691 | ~n18690;
  assign n18694 = ~n18041 | ~n18829;
  assign n18693 = ~n18563 | ~n23035;
  assign n18699 = n18694 & n18693;
  assign n18696 = ~n18041 | ~n18563;
  assign n18695 = ~n18829 | ~n23035;
  assign n18698 = ~n18696 | ~n18695;
  assign n18697 = ~n18699 | ~n18698;
  assign n18701 = ~n18698;
  assign n18700 = ~n18699;
  assign n18704 = ~n18702 | ~n18735;
  assign n18703 = n13123 | n22176;
  assign n18709 = n18704 & n18703;
  assign n18706 = ~n22998 & ~n13123;
  assign n18705 = ~n22176 & ~n18779;
  assign n18708 = n18706 | n18705;
  assign n18707 = ~n18709 | ~n18708;
  assign n18711 = ~n18708;
  assign n18710 = ~n18709;
  assign n18712 = ~n18711 | ~n18710;
  assign n18714 = ~n22702 | ~n18829;
  assign n18713 = ~n22999 | ~n18563;
  assign n18720 = n18714 & n18713;
  assign n18716 = ~n22702 | ~n18563;
  assign n18715 = ~n22999 | ~n18829;
  assign n18719 = ~n18716 | ~n18715;
  assign n18717 = ~n18720 | ~n18719;
  assign n18724 = ~n18718 | ~n18717;
  assign n18722 = ~n18719;
  assign n18721 = ~n18720;
  assign n18723 = ~n18722 | ~n18721;
  assign n18726 = ~n22295 | ~n18563;
  assign n18725 = ~n22982 | ~n18829;
  assign n18730 = n18726 & n18725;
  assign n18728 = ~n22295 | ~n18829;
  assign n18727 = ~n22982 | ~n18563;
  assign n18729 = ~n18728 | ~n18727;
  assign n18732 = ~n18731 | ~n18730;
  assign n18734 = ~n22664 | ~n18735;
  assign n18733 = ~n24289 | ~n18563;
  assign n18740 = n18734 & n18733;
  assign n18737 = ~n22664 | ~n18563;
  assign n18736 = ~n24289 | ~n18735;
  assign n18739 = ~n18737 | ~n18736;
  assign n18738 = ~n18740 | ~n18739;
  assign n18742 = ~n18739;
  assign n18741 = ~n18740;
  assign n18743 = ~n18742 | ~n18741;
  assign n18746 = ~n22223 | ~n18563;
  assign n18745 = ~n24292 | ~n18829;
  assign n18751 = n18746 & n18745;
  assign n18748 = ~n22223 | ~n18829;
  assign n18747 = ~n24292 | ~n18563;
  assign n18750 = ~n18748 | ~n18747;
  assign n18749 = n18751 & n18750;
  assign n18753 = ~n18750;
  assign n18752 = ~n18751;
  assign n18754 = ~n18753 | ~n18752;
  assign n18759 = ~n18756;
  assign n18758 = ~n18757;
  assign n18760 = ~n18759 | ~n18758;
  assign n18765 = ~n18762;
  assign n18764 = ~n18763;
  assign n18766 = ~n18765 | ~n18764;
  assign n18768 = n22889 | n13123;
  assign n18767 = ~n24301 | ~n18829;
  assign n18774 = n18768 & n18767;
  assign n18770 = n22889 | n18779;
  assign n18769 = ~n24301 | ~n18563;
  assign n18773 = ~n18770 | ~n18769;
  assign n18771 = ~n18774 | ~n18773;
  assign n18778 = ~n18772 | ~n18771;
  assign n18776 = ~n18773;
  assign n18775 = ~n18774;
  assign n18777 = ~n18776 | ~n18775;
  assign n18788 = n18778 & n18777;
  assign n18781 = n22874 | n18779;
  assign n18780 = ~n24304 | ~n18563;
  assign n18789 = ~n18781 | ~n18780;
  assign n18787 = ~n18788 | ~n18789;
  assign n18783 = ~n22862 | ~n18563;
  assign n18782 = ~n24308 | ~n18829;
  assign n18797 = n18783 & n18782;
  assign n18785 = ~n22862 | ~n18829;
  assign n18784 = ~n24308 | ~n18563;
  assign n18796 = ~n18785 | ~n18784;
  assign n18786 = ~n18797 | ~n18796;
  assign n18791 = ~n18788;
  assign n18790 = ~n18789;
  assign n18795 = ~n18791 | ~n18790;
  assign n18793 = n22874 | n13123;
  assign n18792 = ~n24304 | ~n18829;
  assign n18794 = n18793 & n18792;
  assign n18799 = ~n18796;
  assign n18798 = ~n18797;
  assign n18800 = ~n18799 | ~n18798;
  assign n18802 = ~n22495 | ~n18829;
  assign n18801 = ~n24311 | ~n18563;
  assign n18809 = ~n18802 | ~n18801;
  assign n18804 = ~n18805 | ~n18563;
  assign n18803 = ~n14111 | ~n18829;
  assign n18815 = n18804 & n18803;
  assign n18807 = ~n18805 | ~n18829;
  assign n18806 = ~n14111 | ~n18563;
  assign n18814 = ~n18807 | ~n18806;
  assign n18808 = ~n18815 & ~n18814;
  assign n18812 = ~n22495 | ~n18563;
  assign n18811 = ~n24311 | ~n18829;
  assign n18813 = ~n18812 | ~n18811;
  assign n18816 = ~n18815 | ~n18814;
  assign n18818 = ~n22819 | ~n18829;
  assign n18817 = ~n18563 | ~n24316;
  assign n18824 = n18818 & n18817;
  assign n18820 = ~n22819 | ~n18563;
  assign n18819 = ~n18829 | ~n24316;
  assign n18823 = ~n18820 | ~n18819;
  assign n18821 = ~n18824 | ~n18823;
  assign n18828 = ~n18822 | ~n18821;
  assign n18826 = ~n18823;
  assign n18825 = ~n18824;
  assign n18827 = ~n18826 | ~n18825;
  assign n18834 = ~n18828 | ~n18827;
  assign n18831 = ~n19095 | ~n18829;
  assign n18830 = ~n18563 | ~n24320;
  assign n18838 = n18831 & n18830;
  assign n18833 = ~n19095 | ~n18563;
  assign n18832 = ~n18829 | ~n24320;
  assign n18837 = ~n18833 | ~n18832;
  assign n18840 = ~n18836 & ~n18835;
  assign n18839 = ~n18838 & ~n18837;
  assign n18841 = ~n18840 & ~n18839;
  assign n18847 = ~n18844;
  assign n18846 = ~n18845;
  assign n18848 = ~n18847 | ~n18846;
  assign n18851 = ~n18901 | ~n18848;
  assign n18850 = ~n18849;
  assign n18852 = ~n18851 | ~n18850;
  assign n18855 = ~n18854 | ~n18853;
  assign n18857 = ~n18856 | ~n18855;
  assign n18858 = ~n18857 | ~n23970;
  assign n18862 = n18859 ^ ~n18858;
  assign n19081 = n19085 ^ ~n18863;
  assign n19098 = ~n19081;
  assign n18898 = ~n18865 | ~n22509;
  assign n22521 = ~n22514;
  assign n18867 = ~n18866;
  assign n23910 = n18867 | n23880;
  assign n18870 = ~n18868;
  assign n23990 = n18870 | n18869;
  assign n18875 = ~n23910 | ~n23990;
  assign n23885 = ~n18872 | ~n18871;
  assign n18873 = ~n18544 | ~n24027;
  assign n24121 = ~n18873 | ~n23983;
  assign n18874 = ~n23885 | ~n24121;
  assign n18878 = ~n18875 & ~n18874;
  assign n18879 = ~n18878 | ~n23851;
  assign n18880 = ~n18879 & ~n23831;
  assign n18884 = ~n18881 | ~n23796;
  assign n22786 = ~n18883 | ~n18882;
  assign n18886 = ~n18884 & ~n22786;
  assign n18888 = ~n18886 | ~n18885;
  assign n18889 = ~n18888 & ~n18887;
  assign n18890 = ~n22728 | ~n18889;
  assign n22694 = ~n18892 | ~n18891;
  assign n18894 = ~n18893 | ~n22655;
  assign n18895 = ~n22521 & ~n18894;
  assign n18897 = ~n18896 | ~n22585;
  assign n18903 = n18902 ^ ~n23723;
  assign n18906 = ~n22789 & ~n16818;
  assign n18913 = ~n18907 | ~n18906;
  assign n18911 = ~n18909 & ~n18908;
  assign n18912 = ~n18911 & ~n18910;
  assign n18914 = ~n18913 | ~n18912;
  assign n18917 = n25399 ^ ~n18920;
  assign n18918 = n25252 & n24449;
  assign n18919 = n18917 | n18918;
  assign n18921 = n25410 ^ ~n18920;
  assign n18922 = ~n25214 | ~n24449;
  assign n24366 = n18921 ^ ~n18922;
  assign n18924 = ~n24365 | ~n24366;
  assign n18923 = ~n18921;
  assign n18925 = n25420 ^ ~n18920;
  assign n18926 = n25183 & n24449;
  assign n24422 = ~n18925 | ~n18926;
  assign n24423 = n18926 | n18925;
  assign n24410 = ~n18927 | ~n24423;
  assign n18928 = n25432 ^ ~n18920;
  assign n18929 = n25150 & n24449;
  assign n18933 = n18928 | n18929;
  assign n18931 = ~n18928;
  assign n18930 = ~n18929;
  assign n18932 = n18931 | n18930;
  assign n24411 = n18933 & n18932;
  assign n18935 = ~n25126 | ~n24449;
  assign n24505 = n18936 ^ ~n18935;
  assign n18934 = ~n24505;
  assign n18940 = ~n25022 | ~n24449;
  assign n18941 = ~n18939;
  assign n18942 = n18941 | n18940;
  assign n18944 = n25467 ^ ~n18920;
  assign n18943 = n25049 & n24449;
  assign n24378 = n18944 & n18943;
  assign n24379 = n18944 | n18943;
  assign n18945 = n25479 ^ ~n18920;
  assign n18946 = n25021 & n24449;
  assign n18950 = n18945 | n18946;
  assign n18948 = ~n18945;
  assign n18947 = ~n18946;
  assign n18949 = n18948 | n18947;
  assign n24438 = n18950 & n18949;
  assign n18951 = n25489 ^ ~n18920;
  assign n18952 = ~n25000 | ~n24449;
  assign n24353 = n18951 ^ ~n18952;
  assign n18953 = ~n18951;
  assign n18954 = n18953 | n18952;
  assign n18955 = n25506 ^ ~n18920;
  assign n18956 = n24976 & n24449;
  assign n20974 = n18955 | n18956;
  assign n18959 = ~n20976 | ~n20974;
  assign n18958 = ~n18955;
  assign n18957 = ~n18956;
  assign n20973 = n18958 | n18957;
  assign n18960 = n24394 ^ ~n18920;
  assign n18961 = n24955 & n24449;
  assign n24401 = n18960 | n18961;
  assign n18963 = ~n18960;
  assign n18962 = ~n18961;
  assign n24402 = n18963 | n18962;
  assign n18965 = n24473 ^ ~n18920;
  assign n18964 = n21817 & n24449;
  assign n24467 = n18965 & n18964;
  assign n24466 = n18965 | n18964;
  assign n18966 = n22018 ^ ~n18920;
  assign n18967 = n21735 & n24449;
  assign n18981 = n18966 | n18967;
  assign n18969 = ~n18966;
  assign n18968 = ~n18967;
  assign n18970 = n18969 | n18968;
  assign n20899 = n18981 & n18970;
  assign n20896 = n22029 ^ ~n19033;
  assign n18977 = ~n21818 | ~n24449;
  assign n18971 = n20896 | n18977;
  assign n20903 = ~n20899 | ~n18971;
  assign n18973 = n22041 ^ ~n19033;
  assign n18974 = ~n21413 | ~n24449;
  assign n20819 = n18973 ^ ~n18974;
  assign n18972 = ~n20903 & ~n20819;
  assign n18984 = ~n20818 | ~n18972;
  assign n18980 = ~n20903;
  assign n18976 = ~n18973;
  assign n18975 = ~n18974;
  assign n21017 = ~n18977;
  assign n18979 = ~n20892 | ~n21017;
  assign n20894 = ~n20896;
  assign n18978 = ~n20892 | ~n20894;
  assign n20901 = n18979 & n18978;
  assign n18982 = ~n18980 | ~n20901;
  assign n18983 = n18982 & n18981;
  assign n20918 = ~n18984 | ~n18983;
  assign n18985 = n22008 ^ ~n18920;
  assign n18986 = n21436 & n24449;
  assign n18990 = n18985 | n18986;
  assign n18988 = ~n18985;
  assign n18987 = ~n18986;
  assign n18989 = n18988 | n18987;
  assign n20917 = n18990 & n18989;
  assign n18993 = n21997 ^ ~n19033;
  assign n18992 = ~n21734 | ~n24449;
  assign n20987 = n18993 ^ ~n18992;
  assign n18991 = ~n20987;
  assign n18994 = n18993 | n18992;
  assign n18995 = n21986 ^ ~n18920;
  assign n18996 = n25556 & n24449;
  assign n20851 = n18995 | n18996;
  assign n18998 = ~n18995;
  assign n18997 = ~n18996;
  assign n20850 = n18998 | n18997;
  assign n18999 = n21975 ^ ~n18920;
  assign n19000 = n25559 & n24449;
  assign n20944 = n18999 | n19000;
  assign n19002 = ~n18999;
  assign n19001 = ~n19000;
  assign n20943 = n19002 | n19001;
  assign n19005 = n21965 ^ ~n18920;
  assign n19004 = n25562 & n24449;
  assign n19006 = n21954 ^ ~n18920;
  assign n20961 = ~n25565 | ~n24449;
  assign n19010 = ~n20959 | ~n20961;
  assign n19007 = ~n19006;
  assign n19011 = n21598 ^ ~n18920;
  assign n20834 = ~n19009 | ~n19011;
  assign n20836 = n25568 & n24449;
  assign n19014 = ~n20834 | ~n20836;
  assign n19012 = ~n19011;
  assign n20835 = ~n19010 | ~n19013;
  assign n19015 = n21932 ^ ~n18920;
  assign n19016 = ~n25571 | ~n24449;
  assign n20930 = n19015 ^ ~n19016;
  assign n19017 = ~n19015;
  assign n19018 = n19017 | n19016;
  assign n19021 = n21921 ^ ~n18920;
  assign n19019 = ~n25574 | ~n24449;
  assign n20879 = n19021 ^ ~n19019;
  assign n19020 = ~n19019;
  assign n19022 = ~n19021 | ~n19020;
  assign n19023 = n21910 ^ ~n18920;
  assign n19024 = n25577 & n24449;
  assign n19026 = ~n19023;
  assign n19025 = ~n19024;
  assign n19027 = n19026 | n19025;
  assign n21002 = ~n19029 | ~n19027;
  assign n19028 = ~n21002;
  assign n19031 = n21323 ^ ~n19033;
  assign n19030 = ~n25580 | ~n24449;
  assign n20805 = n19031 ^ ~n19030;
  assign n19032 = n19031 | n19030;
  assign n19034 = ~n25583 | ~n24449;
  assign n19043 = n19034 ^ ~n19033;
  assign n19035 = ~n19043 | ~n21025;
  assign n19037 = ~n21487 & ~n19035;
  assign n19036 = ~n21333 & ~n19043;
  assign n19038 = ~n19037 & ~n19036;
  assign n19041 = ~n19042 & ~n19038;
  assign n19039 = ~n21487 & ~n21025;
  assign n19040 = ~n19039 & ~n24506;
  assign n19046 = ~n21487 | ~n19043;
  assign n19044 = ~n19043 & ~n24508;
  assign n19045 = ~n21333 | ~n19044;
  assign n19047 = ~n19046 | ~n19045;
  assign n19048 = ~n19042 | ~n19047;
  assign n19059 = ~n19049 | ~n19048;
  assign n19050 = ~n21478;
  assign n19055 = ~n19050 & ~n24511;
  assign n19053 = n24484 | n19051;
  assign n19052 = ~P2_REG3_REG_28__SCAN_IN | ~P2_U3088;
  assign n19054 = ~n19053 | ~n19052;
  assign n19057 = ~n19055 & ~n19054;
  assign n19056 = ~n25586 | ~n24455;
  assign n19058 = n19057 & n19056;
  assign P2_U3192 = ~n19059 | ~n19058;
  assign n19063 = ~n19061;
  assign n19062 = ~P3_ADDR_REG_17__SCAN_IN;
  assign n19067 = ~n19065 | ~n13265;
  assign n23685 = ~P1_ADDR_REG_18__SCAN_IN;
  assign n19068 = n23685 ^ ~P3_ADDR_REG_18__SCAN_IN;
  assign n19066 = n19067 ^ ~n19068;
  assign n23197 = ~n23198 & ~P2_ADDR_REG_18__SCAN_IN;
  assign n19070 = ~n19067;
  assign n19069 = ~n19068;
  assign n19072 = ~n19070 | ~n19069;
  assign n19071 = n23685 | P3_ADDR_REG_18__SCAN_IN;
  assign n19075 = ~n19072 | ~n19071;
  assign n19073 = P2_ADDR_REG_19__SCAN_IN ^ ~P1_ADDR_REG_19__SCAN_IN;
  assign n19074 = n19073 ^ ~n14961;
  assign n19076 = n19075 ^ ~n19074;
  assign SUB_1596_U4 = n19077 ^ ~n19076;
  assign n19080 = ~n19078 | ~n18060;
  assign n19079 = ~n19095 | ~n24320;
  assign n19082 = ~n19080 | ~n19079;
  assign n19083 = ~n24012 & ~n24228;
  assign n19091 = ~n22429 | ~n24216;
  assign n19089 = ~n14526 & ~n24241;
  assign n22435 = ~n19086 | ~n24327;
  assign n19087 = ~n23988 | ~n24320;
  assign n19088 = ~n22435 | ~n19087;
  assign n19090 = ~n19089 & ~n19088;
  assign n19093 = ~n19092 | ~n24320;
  assign n19097 = ~n19094 | ~n19093;
  assign n19096 = ~n19095 | ~n22452;
  assign n19099 = ~n24284 | ~P1_REG1_REG_29__SCAN_IN;
  assign P1_U3557 = ~n19100 | ~n19099;
  assign n19104 = ~n19101;
  assign n19103 = ~n19102;
  assign n19105 = ~n19104 | ~n19103;
  assign n19107 = ~n19106 | ~n19105;
  assign n19118 = ~n19107 | ~n23339;
  assign n19116 = ~n14525 & ~n23277;
  assign n19114 = ~n14111 | ~n23322;
  assign n22463 = ~n19108;
  assign n19112 = ~n23311 & ~n22463;
  assign n19110 = ~n23332 | ~n24320;
  assign n19109 = ~P1_U3086 | ~P1_REG3_REG_27__SCAN_IN;
  assign n19111 = ~n19110 | ~n19109;
  assign n19113 = ~n19112 & ~n19111;
  assign n19115 = ~n19114 | ~n19113;
  assign n19117 = ~n19116 & ~n19115;
  assign P1_U3214 = ~n19118 | ~n19117;
  assign n19119 = n19413 ^ ~n17213;
  assign n19668 = ~n19119 | ~n20435;
  assign n19120 = n19119 | n20435;
  assign n19652 = ~n19668 | ~n19120;
  assign n19792 = n20648 ^ ~n17213;
  assign n19121 = n19792 & n19646;
  assign n19161 = ~n19666;
  assign n19122 = n20656 ^ ~n17213;
  assign n19128 = n19122 | n19406;
  assign n19123 = ~n19122;
  assign n19124 = n19123 | n20472;
  assign n19549 = ~n19128 | ~n19124;
  assign n19737 = n20665 ^ ~n19178;
  assign n19125 = ~n19737;
  assign n19157 = ~n19125 | ~n19552;
  assign n19126 = ~n19737 | ~n20495;
  assign n19156 = n20507 ^ ~n17213;
  assign n19127 = n19549 | n19547;
  assign n19644 = n19128 & n19127;
  assign n25672 = ~n19130 | ~n19129;
  assign n19131 = n17213 ^ ~n26351;
  assign n19133 = n19131 | n26205;
  assign n19132 = ~n19131 | ~n26205;
  assign n25671 = n19133 & n19132;
  assign n19136 = n17213 ^ ~n26150;
  assign n25731 = n19136 ^ ~n26189;
  assign n19137 = ~n25603;
  assign n25600 = n19136 | n26138;
  assign n19140 = n19137 | n25600;
  assign n19139 = ~n19138 | ~n26165;
  assign n19141 = n19140 & n19139;
  assign n19142 = n19360 ^ ~n17213;
  assign n25643 = n19142 ^ ~n26086;
  assign n19143 = ~n19142;
  assign n19144 = ~n19143 | ~n26086;
  assign n19146 = n26383 ^ ~n17213;
  assign n19149 = n19146 | n26116;
  assign n19147 = ~n19146;
  assign n19148 = n19147 | n25638;
  assign n19704 = ~n19149 | ~n19148;
  assign n19150 = n26393 ^ ~n17213;
  assign n25615 = n19150 ^ ~n26085;
  assign n19151 = ~n19150;
  assign n19152 = n19151 | n25689;
  assign n25695 = n20681 ^ ~n17213;
  assign n19153 = n25695 | n26059;
  assign n19154 = ~n25695;
  assign n19155 = n19154 | n25611;
  assign n19614 = n19156 | n20517;
  assign n19546 = n19614 & n19157;
  assign n19158 = ~n19549;
  assign n19643 = n19546 & n19158;
  assign n19159 = n19643 & n19666;
  assign n19664 = n19792 | n19646;
  assign n19164 = ~n19161 & ~n19664;
  assign n19670 = n20632 ^ ~n17213;
  assign n19162 = n19670 | n19771;
  assign n19163 = ~n19162 | ~n19668;
  assign n19165 = ~n19164 & ~n19163;
  assign n19167 = ~n19670;
  assign n19168 = n19167 | n20416;
  assign n19169 = n19427 ^ ~n17213;
  assign n19765 = n19169 | n20398;
  assign n19170 = ~n19169;
  assign n19579 = n20369 ^ ~n19178;
  assign n19171 = n20349 ^ ~n19178;
  assign n19719 = n19171 | n19602;
  assign n19172 = n18431 ^ ~n17213;
  assign n19596 = n19172 | n20334;
  assign n19173 = ~n19172;
  assign n19175 = ~n19174 & ~n13231;
  assign n19563 = n20585 ^ ~n19178;
  assign n19179 = n18436 ^ ~n17213;
  assign n19183 = n19179 | n20266;
  assign n19180 = ~n19179;
  assign n19181 = n19180 | n20210;
  assign n19688 = n19183 & n19181;
  assign n19182 = ~n19563 | ~n19692;
  assign n19184 = ~n19183;
  assign n19186 = n20220 ^ ~n17213;
  assign n19189 = ~n19186 | ~n20235;
  assign n19187 = ~n19186;
  assign n19188 = ~n19187 | ~n26436;
  assign n19629 = ~n19189 | ~n19188;
  assign n19190 = ~n19189;
  assign n19191 = n20197 ^ ~n17213;
  assign n19194 = ~n19191 | ~n20209;
  assign n19192 = ~n19191;
  assign n19193 = ~n19192 | ~n26439;
  assign n19195 = ~n19194;
  assign n19201 = n20174 ^ ~n19178;
  assign n19198 = n19201 | n26442;
  assign n19196 = ~n19201;
  assign n19197 = n19196 | n20186;
  assign n19532 = ~n19198 | ~n19197;
  assign n19215 = n20141 ^ ~n17213;
  assign n19199 = n19198 & n25732;
  assign n19203 = ~n19215;
  assign n19200 = ~n20186 | ~n25732;
  assign n19202 = ~n19201 & ~n19200;
  assign n19214 = ~n19203 | ~n19202;
  assign n19212 = ~n14256 & ~n25725;
  assign n19210 = ~n26442 | ~n25706;
  assign n25654 = ~n25734;
  assign n19204 = ~n20152;
  assign n19208 = ~n25654 & ~n19204;
  assign n20147 = ~n26448;
  assign n19206 = n25666 | n20147;
  assign n19205 = ~P3_REG3_REG_28__SCAN_IN | ~P3_U3151;
  assign n19207 = ~n19206 | ~n19205;
  assign n19209 = ~n19208 & ~n19207;
  assign n19211 = ~n19210 | ~n19209;
  assign n19213 = ~n19212 & ~n19211;
  assign n25684 = ~n25732;
  assign n19216 = ~n19215 & ~n25684;
  assign n19218 = ~n19217 | ~n19216;
  assign P3_U3160 = ~n19219 | ~n19218;
  assign n19220 = ~n24240 | ~P1_REG0_REG_29__SCAN_IN;
  assign n19221 = ~n19503 & ~n20147;
  assign n19227 = ~n19224 | ~n19223;
  assign n19226 = ~n19225 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n19240 = P1_DATAO_REG_30__SCAN_IN ^ ~P2_DATAO_REG_30__SCAN_IN;
  assign n20760 = ~SI_30_;
  assign n19229 = n18176 | n20760;
  assign n19238 = ~n20539;
  assign n19232 = ~n16422 | ~P3_REG2_REG_31__SCAN_IN;
  assign n19236 = ~n19232 | ~n19231;
  assign n19234 = ~n16463 | ~P3_REG1_REG_31__SCAN_IN;
  assign n19233 = ~n18380 | ~P3_REG0_REG_31__SCAN_IN;
  assign n19235 = ~n19234 | ~n19233;
  assign n19237 = ~n20129 & ~n19509;
  assign n19255 = ~n19503 | ~n20147;
  assign n19239 = ~n19255 | ~n20119;
  assign n19246 = ~n19248 & ~n19239;
  assign n19241 = ~n23125 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n19244 = ~n19242 | ~n19241;
  assign n19243 = P1_DATAO_REG_31__SCAN_IN ^ ~P2_DATAO_REG_31__SCAN_IN;
  assign n19245 = ~n13121 | ~SI_31_;
  assign n19516 = ~n19269 | ~n26455;
  assign n19247 = ~n19255;
  assign n19249 = ~n19247 & ~n26455;
  assign n19256 = ~n19248;
  assign n19250 = ~n19249 | ~n19256;
  assign n19251 = ~n19250 | ~n19257;
  assign n19263 = ~n19253 & ~n19252;
  assign n19511 = n20539 | n19509;
  assign n19265 = ~n19511 | ~n26455;
  assign n19254 = ~n19265 | ~n20119;
  assign n19261 = ~n19254 & ~n19269;
  assign n19258 = ~n19256 | ~n19255;
  assign n19259 = ~n19258 | ~n19257;
  assign n19260 = ~n19259 & ~n19265;
  assign n19262 = ~n19261 & ~n19260;
  assign n19264 = ~n19263 | ~n19262;
  assign n19266 = ~n19265;
  assign n19267 = ~n19266 & ~n19269;
  assign n19268 = ~n19267 & ~n20119;
  assign n19514 = n26455 ^ n19269;
  assign n19299 = ~n19514;
  assign n20292 = ~n20261 | ~n20260;
  assign n20362 = n20369 ^ ~n19446;
  assign n20477 = n20665 ^ ~n20495;
  assign n20500 = ~n20493;
  assign n19272 = ~n18399 | ~n14555;
  assign n19278 = ~n19272 & ~n26233;
  assign n19275 = ~n19304 | ~n14005;
  assign n26305 = ~n19275 | ~n19274;
  assign n19276 = ~n19273 | ~n26305;
  assign n19277 = ~n19276 & ~n26181;
  assign n19280 = ~n19279 & ~n26109;
  assign n19281 = ~n19280 | ~n26053;
  assign n26081 = n26383 ^ ~n25638;
  assign n26078 = ~n26081;
  assign n19282 = ~n19281 & ~n26078;
  assign n19283 = ~n19282 | ~n20524;
  assign n19284 = ~n20500 & ~n19283;
  assign n19285 = ~n20477 | ~n19284;
  assign n19286 = ~n14570 & ~n19285;
  assign n19289 = ~n18424 | ~n19288;
  assign n19290 = ~n20292 & ~n13901;
  assign n19291 = ~n19465 | ~n19290;
  assign n19292 = ~n19291 & ~n20330;
  assign n19293 = ~n19292 | ~n13190;
  assign n19294 = ~n20141 & ~n13269;
  assign n19296 = n20539 ^ ~n26451;
  assign n19298 = ~n19297 | ~n19296;
  assign n19302 = n19300 ^ ~n20119;
  assign n19303 = ~n19302 | ~n19301;
  assign n19307 = ~n19313 & ~n19305;
  assign n19311 = ~n19307 & ~n19306;
  assign n19310 = ~n19309 & ~n19308;
  assign n19320 = ~n19311 & ~n19310;
  assign n19318 = ~n19312 & ~n19834;
  assign n19316 = ~n19314 | ~n19834;
  assign n19317 = ~n19316 & ~n19315;
  assign n19319 = ~n19318 & ~n19317;
  assign n19326 = ~n19320 & ~n19319;
  assign n19324 = ~n19321 | ~n19834;
  assign n19323 = ~n19322 | ~n19520;
  assign n19325 = ~n19324 | ~n19323;
  assign n19328 = ~n19327 | ~n19520;
  assign n19332 = ~n19328 & ~n19334;
  assign n19330 = ~n19329 | ~n19834;
  assign n19331 = ~n19330 & ~n19335;
  assign n19337 = ~n19334 & ~n19520;
  assign n19336 = ~n19335 & ~n19834;
  assign n19339 = ~n19338;
  assign n19343 = ~n19339 & ~n19520;
  assign n19341 = ~n19340;
  assign n19342 = ~n19341 & ~n19834;
  assign n19355 = ~n19344 & ~n26181;
  assign n19348 = ~n19345 | ~n19834;
  assign n19347 = ~n19346 | ~n19520;
  assign n19353 = ~n19348 | ~n19347;
  assign n19350 = ~n26138 | ~n19834;
  assign n19349 = ~n26359 | ~n19520;
  assign n19356 = ~n19350 | ~n19349;
  assign n19351 = ~n26138 | ~n26359;
  assign n19352 = ~n19356 | ~n19351;
  assign n19354 = ~n19353 | ~n19352;
  assign n19358 = ~n19356;
  assign n19359 = ~n19358 | ~n19357;
  assign n19362 = ~n19360 & ~n19834;
  assign n19361 = ~n26086 & ~n19520;
  assign n19370 = n19362 | n19361;
  assign n19369 = ~n19370 | ~n19363;
  assign n19365 = ~n26165 | ~n26367;
  assign n19367 = ~n19365 | ~n19520;
  assign n19366 = ~n26107 | ~n19834;
  assign n19368 = ~n19367 | ~n19366;
  assign n19375 = ~n19372 | ~n19834;
  assign n19374 = ~n19373 | ~n19520;
  assign n19376 = ~n19375 | ~n19374;
  assign n20674 = ~n20507;
  assign n19396 = ~n20674 | ~n25692;
  assign n25691 = ~n20681;
  assign n19377 = ~n25691 & ~n25611;
  assign n19378 = ~n19377 & ~n19520;
  assign n19382 = ~n19396 | ~n19378;
  assign n19380 = ~n19379 & ~n19834;
  assign n19381 = ~n19397 | ~n19380;
  assign n19385 = ~n19382 | ~n19381;
  assign n19383 = n26053 & n19385;
  assign n19395 = ~n19384 | ~n19383;
  assign n19394 = ~n19385;
  assign n19386 = ~n26393;
  assign n19387 = ~n19386 & ~n25689;
  assign n19390 = ~n19387 & ~n19834;
  assign n19389 = ~n19388 & ~n19520;
  assign n19392 = ~n19390 & ~n19389;
  assign n19393 = ~n19392 & ~n19391;
  assign n19399 = ~n19396 | ~n19520;
  assign n19398 = ~n19397 | ~n19834;
  assign n19403 = ~n19400 | ~n19834;
  assign n19402 = ~n19401 | ~n19520;
  assign n19404 = ~n19403 | ~n19402;
  assign n19409 = ~n19405 | ~n19834;
  assign n19407 = ~n20656 | ~n19406;
  assign n19408 = ~n19407 | ~n19520;
  assign n19410 = ~n19409 | ~n19408;
  assign n20640 = ~n19413;
  assign n19412 = ~n20640 | ~n19520;
  assign n19411 = ~n20435 | ~n19834;
  assign n19425 = n19412 & n19411;
  assign n19414 = ~n19413 & ~n19795;
  assign n19421 = ~n19425 & ~n19414;
  assign n19416 = ~n19415 & ~n20454;
  assign n19419 = ~n19416 & ~n19834;
  assign n19418 = ~n19417 & ~n19520;
  assign n19420 = ~n19419 & ~n19418;
  assign n19422 = ~n19421 & ~n19420;
  assign n19426 = ~n19425 | ~n19424;
  assign n19429 = n19427 | n19520;
  assign n19428 = ~n20398 | ~n19520;
  assign n19433 = ~n19431 & ~n19430;
  assign n19440 = ~n19431;
  assign n19432 = ~n19440 & ~n20398;
  assign n19437 = ~n19432 & ~n19520;
  assign n19443 = ~n19433;
  assign n19434 = ~n20632;
  assign n19435 = ~n19434 & ~n20416;
  assign n19436 = ~n19443 | ~n19435;
  assign n19439 = ~n19437 | ~n19436;
  assign n19438 = ~n19452 & ~n20369;
  assign n20624 = ~n19427;
  assign n19445 = ~n19441 & ~n19834;
  assign n19444 = ~n19443 | ~n19442;
  assign n19448 = ~n19445 | ~n19444;
  assign n19447 = ~n19452 & ~n19446;
  assign n19451 = ~n19450 & ~n19449;
  assign n19454 = ~n19452;
  assign n20609 = ~n20349;
  assign n19455 = ~n20609 & ~n19602;
  assign n19458 = ~n19455 & ~n19520;
  assign n19457 = ~n19456 & ~n19834;
  assign n19464 = ~n19461 & ~n19520;
  assign n19463 = ~n19462 & ~n19834;
  assign n19469 = ~n19466 | ~n19520;
  assign n19468 = ~n19467 | ~n19834;
  assign n19470 = ~n19469 | ~n19468;
  assign n19477 = ~n19471 | ~n20233;
  assign n19475 = ~n19472 | ~n19834;
  assign n19474 = ~n19473 | ~n19520;
  assign n19476 = ~n19475 | ~n19474;
  assign n19478 = ~n19477 | ~n19476;
  assign n19482 = ~n19479 | ~n19520;
  assign n19481 = ~n19480 | ~n19834;
  assign n19483 = ~n20560 | ~n19520;
  assign n19486 = ~n19483 | ~n26439;
  assign n19484 = ~n20197 | ~n19834;
  assign n19485 = ~n19484 | ~n20209;
  assign n19487 = ~n20552 | ~n19520;
  assign n19490 = ~n19487 | ~n26442;
  assign n19488 = ~n20174 | ~n19834;
  assign n19489 = ~n19488 | ~n20186;
  assign n19491 = ~n19490 | ~n19489;
  assign n20155 = ~n20141;
  assign n19498 = ~n19492 | ~n20155;
  assign n19496 = ~n19493 | ~n19520;
  assign n19495 = ~n19494 | ~n19834;
  assign n19497 = ~n19496 | ~n19495;
  assign n19500 = ~n19498 | ~n19497;
  assign n19508 = ~n19500 | ~n19499;
  assign n19502 = ~n19501 | ~n19520;
  assign n19506 = ~n19502 | ~n26448;
  assign n19504 = ~n19503 | ~n19834;
  assign n19505 = ~n19504 | ~n20147;
  assign n19507 = ~n19506 | ~n19505;
  assign n19512 = ~n20539 | ~n19509;
  assign n19515 = ~n20535 | ~n20129;
  assign n19518 = ~n19515 | ~n19834;
  assign n19517 = ~n19516 | ~n19520;
  assign n19519 = ~n19518 | ~n19517;
  assign n19521 = n19520 ^ ~n20119;
  assign n19832 = ~n19835;
  assign n19523 = n20078 & n19950;
  assign n19525 = ~n19524 | ~n19523;
  assign n19529 = n19525 & P3_B_REG_SCAN_IN;
  assign n19527 = ~n19832 | ~n19526;
  assign n19528 = ~n19529 | ~n19527;
  assign n19530 = ~n19529;
  assign n19531 = ~n19530 | ~P3_U3151;
  assign n19534 = n19533 ^ ~n19532;
  assign n19544 = ~n19534 | ~n25732;
  assign n19542 = ~n20552 & ~n25725;
  assign n19538 = ~n20209 & ~n25724;
  assign n19536 = n25666 | n20165;
  assign n19535 = ~P3_REG3_REG_27__SCAN_IN | ~P3_U3151;
  assign n19537 = ~n19536 | ~n19535;
  assign n19540 = ~n19538 & ~n19537;
  assign n19539 = ~n20175 | ~n25734;
  assign n19541 = ~n19540 | ~n19539;
  assign n19543 = ~n19542 & ~n19541;
  assign P3_U3154 = ~n19544 | ~n19543;
  assign n19548 = ~n19545 | ~n19546;
  assign n19550 = n19548 & n19547;
  assign n19551 = n19550 ^ ~n19549;
  assign n19561 = ~n19551 | ~n25732;
  assign n19559 = ~n20656 & ~n25725;
  assign n19557 = ~n25734 | ~n20463;
  assign n19553 = ~n25706 | ~n19552;
  assign n26035 = ~P3_REG3_REG_14__SCAN_IN | ~P3_U3151;
  assign n19555 = ~n19553 | ~n26035;
  assign n19554 = ~n25666 & ~n20454;
  assign n19556 = ~n19555 & ~n19554;
  assign n19558 = ~n19557 | ~n19556;
  assign n19560 = ~n19559 & ~n19558;
  assign P3_U3155 = ~n19561 | ~n19560;
  assign n19562 = ~n19565;
  assign n19685 = ~n19562 & ~n19563;
  assign n19564 = ~n19563;
  assign n19566 = ~n19565 & ~n19564;
  assign n19684 = ~n19685 & ~n19566;
  assign n19567 = n19684 ^ ~n20287;
  assign n19578 = ~n19567 | ~n25732;
  assign n19576 = ~n19568 & ~n25725;
  assign n19572 = ~n20210 & ~n25666;
  assign n19570 = ~n20267 | ~n25706;
  assign n19569 = ~P3_REG3_REG_23__SCAN_IN | ~P3_U3151;
  assign n19571 = ~n19570 | ~n19569;
  assign n19574 = ~n19572 & ~n19571;
  assign n19573 = ~n20273 | ~n25734;
  assign n19575 = ~n19574 | ~n19573;
  assign n19577 = ~n19576 & ~n19575;
  assign P3_U3156 = ~n19578 | ~n19577;
  assign n19580 = n19579 ^ ~n20376;
  assign n19582 = n19581 ^ ~n19580;
  assign n19593 = ~n19582 | ~n25732;
  assign n20616 = ~n20369;
  assign n19591 = ~n20616 & ~n25725;
  assign n19586 = ~n20354 & ~n25666;
  assign n19584 = ~n19674 | ~n25706;
  assign n20120 = P3_STATE_REG_SCAN_IN | n19583;
  assign n19585 = ~n19584 | ~n20120;
  assign n19589 = ~n19586 & ~n19585;
  assign n20359 = ~n19587;
  assign n19588 = ~n25734 | ~n20359;
  assign n19590 = ~n19589 | ~n19588;
  assign n19592 = ~n19591 & ~n19590;
  assign P3_U3159 = ~n19593 | ~n19592;
  assign n19595 = ~n19594;
  assign n19600 = ~n19595 | ~n19597;
  assign n19598 = ~n19597 | ~n19596;
  assign n19599 = ~n13167 | ~n19598;
  assign n19601 = ~n19600 | ~n19599;
  assign n19612 = ~n19601 | ~n25732;
  assign n19610 = ~n20601 & ~n25725;
  assign n19606 = ~n20310 & ~n25666;
  assign n19604 = ~n19602 | ~n25706;
  assign n19603 = ~P3_REG3_REG_21__SCAN_IN | ~P3_U3151;
  assign n19605 = ~n19604 | ~n19603;
  assign n19608 = ~n19606 & ~n19605;
  assign n19607 = ~n25734 | ~n20321;
  assign n19609 = ~n19608 | ~n19607;
  assign n19611 = ~n19610 & ~n19609;
  assign P3_U3163 = ~n19612 | ~n19611;
  assign n19736 = ~n19545 | ~n19614;
  assign n19613 = ~n19736;
  assign n19618 = ~n19613 | ~n19735;
  assign n19616 = ~n19545;
  assign n19615 = ~n19735 | ~n19614;
  assign n19617 = ~n19616 | ~n19615;
  assign n19619 = ~n19618 | ~n19617;
  assign n19628 = ~n19619 | ~n25732;
  assign n19626 = ~n20674 & ~n25725;
  assign n19624 = ~n25734 | ~n20508;
  assign n19620 = ~n25706 | ~n26059;
  assign n25990 = ~P3_U3151 | ~P3_REG3_REG_12__SCAN_IN;
  assign n19622 = ~n19620 | ~n25990;
  assign n19621 = ~n25666 & ~n20495;
  assign n19623 = ~n19622 & ~n19621;
  assign n19625 = ~n19624 | ~n19623;
  assign n19627 = ~n19626 & ~n19625;
  assign P3_U3164 = ~n19628 | ~n19627;
  assign n19631 = n19630 ^ ~n19629;
  assign n19642 = ~n19631 | ~n25732;
  assign n20568 = ~n20220;
  assign n19640 = ~n20568 & ~n25725;
  assign n19632 = ~n20221;
  assign n19636 = ~n19632 & ~n25654;
  assign n19634 = ~n20266 | ~n25706;
  assign n19633 = ~P3_REG3_REG_25__SCAN_IN | ~P3_U3151;
  assign n19635 = ~n19634 | ~n19633;
  assign n19638 = ~n19636 & ~n19635;
  assign n19637 = ~n26439 | ~n25728;
  assign n19639 = ~n19638 | ~n19637;
  assign n19641 = ~n19640 & ~n19639;
  assign P3_U3165 = ~n19642 | ~n19641;
  assign n19645 = ~n19545 | ~n19643;
  assign n19647 = ~n19645 | ~n19644;
  assign n19665 = ~n19647;
  assign n19648 = ~n19665 | ~n19646;
  assign n19649 = ~n19647 | ~n20454;
  assign n19793 = ~n19648 | ~n19649;
  assign n19651 = ~n19793 & ~n19792;
  assign n19650 = ~n19649;
  assign n19653 = ~n19651 & ~n19650;
  assign n19654 = n19653 ^ ~n19652;
  assign n19663 = ~n19654 | ~n25732;
  assign n19661 = ~n20640 & ~n25725;
  assign n19659 = ~n25734 | ~n20425;
  assign n19655 = ~n19771 | ~n25728;
  assign n20022 = ~P3_REG3_REG_16__SCAN_IN | ~P3_U3151;
  assign n19657 = ~n19655 | ~n20022;
  assign n19656 = ~n25724 & ~n20454;
  assign n19658 = ~n19657 & ~n19656;
  assign n19660 = ~n19659 | ~n19658;
  assign n19662 = ~n19661 & ~n19660;
  assign P3_U3166 = ~n19663 | ~n19662;
  assign n19667 = ~n19665 | ~n19664;
  assign n19669 = ~n19667 | ~n19666;
  assign n19672 = ~n19669 | ~n19668;
  assign n19671 = n19670 ^ ~n20416;
  assign n19673 = n19672 ^ ~n19671;
  assign n19683 = ~n19673 | ~n25732;
  assign n19681 = ~n20632 & ~n25725;
  assign n19679 = ~n25734 | ~n20407;
  assign n19675 = ~n19674 | ~n25728;
  assign n20050 = ~P3_REG3_REG_17__SCAN_IN | ~P3_U3151;
  assign n19677 = ~n19675 | ~n20050;
  assign n19676 = ~n20435 & ~n25724;
  assign n19678 = ~n19677 & ~n19676;
  assign n19680 = ~n19679 | ~n19678;
  assign n19682 = ~n19681 & ~n19680;
  assign P3_U3168 = ~n19683 | ~n19682;
  assign n19687 = ~n19684 | ~n20287;
  assign n19686 = ~n19685;
  assign n19689 = ~n19687 | ~n19686;
  assign n19690 = n19689 ^ ~n19688;
  assign n19702 = ~n19690 | ~n25732;
  assign n19700 = ~n18436 & ~n25725;
  assign n19698 = ~n26436 | ~n25728;
  assign n19691 = ~n20246;
  assign n19696 = ~n19691 & ~n25654;
  assign n19694 = ~n19692 | ~n25706;
  assign n19693 = ~P3_REG3_REG_24__SCAN_IN | ~P3_U3151;
  assign n19695 = ~n19694 | ~n19693;
  assign n19697 = ~n19696 & ~n19695;
  assign n19699 = ~n19698 | ~n19697;
  assign n19701 = ~n19700 & ~n19699;
  assign P3_U3169 = ~n19702 | ~n19701;
  assign n19717 = ~n25734 | ~n26094;
  assign n19715 = ~n26383 & ~n25725;
  assign n19713 = ~n25724 & ~n26125;
  assign n19705 = ~n19704 | ~n19703;
  assign n19707 = ~n19706 | ~n19705;
  assign n19711 = ~n25732 | ~n19707;
  assign n25924 = ~n19708 & ~P3_STATE_REG_SCAN_IN;
  assign n19709 = ~n25689 & ~n25666;
  assign n19710 = ~n25924 & ~n19709;
  assign n19712 = ~n19711 | ~n19710;
  assign n19714 = n19713 | n19712;
  assign n19716 = ~n19715 & ~n19714;
  assign P3_U3171 = ~n19717 | ~n19716;
  assign n19718 = ~n13301;
  assign n19723 = ~n19718 | ~n19719;
  assign n19720 = ~n14882 | ~n19719;
  assign n19722 = ~n19721 | ~n19720;
  assign n19724 = ~n19723 | ~n19722;
  assign n19734 = ~n19724 | ~n25732;
  assign n19732 = ~n20609 & ~n25725;
  assign n19726 = ~n19752 | ~n25728;
  assign n19725 = ~P3_REG3_REG_20__SCAN_IN | ~P3_U3151;
  assign n19728 = ~n19726 | ~n19725;
  assign n19727 = ~n20376 & ~n25724;
  assign n19730 = ~n19728 & ~n19727;
  assign n19729 = ~n25734 | ~n20342;
  assign n19731 = ~n19730 | ~n19729;
  assign n19733 = ~n19732 & ~n19731;
  assign P3_U3173 = ~n19734 | ~n19733;
  assign n19739 = n19736 & n19735;
  assign n19738 = n19737 ^ ~n20495;
  assign n19740 = n19739 ^ ~n19738;
  assign n19749 = ~n19740 | ~n25732;
  assign n19747 = ~n20665 & ~n25725;
  assign n19745 = ~n25734 | ~n20485;
  assign n19741 = ~n25706 | ~n25692;
  assign n26016 = ~P3_REG3_REG_13__SCAN_IN | ~P3_U3151;
  assign n19743 = ~n19741 | ~n26016;
  assign n19742 = ~n25666 & ~n20472;
  assign n19744 = ~n19743 & ~n19742;
  assign n19746 = ~n19745 | ~n19744;
  assign n19748 = ~n19747 & ~n19746;
  assign P3_U3174 = ~n19749 | ~n19748;
  assign n19751 = n19750 ^ ~n20310;
  assign n19762 = ~n19751 | ~n25732;
  assign n19760 = ~n20593 & ~n25725;
  assign n19756 = ~n20287 & ~n25666;
  assign n19754 = ~n19752 | ~n25706;
  assign n19753 = ~P3_REG3_REG_22__SCAN_IN | ~P3_U3151;
  assign n19755 = ~n19754 | ~n19753;
  assign n19758 = ~n19756 & ~n19755;
  assign n19757 = ~n20299 | ~n25734;
  assign n19759 = ~n19758 | ~n19757;
  assign n19761 = ~n19760 & ~n19759;
  assign P3_U3175 = ~n19762 | ~n19761;
  assign n19764 = ~n19763;
  assign n19769 = ~n19764 | ~n19766;
  assign n19767 = ~n19766 | ~n19765;
  assign n19768 = ~n13389 | ~n19767;
  assign n19770 = ~n19769 | ~n19768;
  assign n19780 = ~n19770 | ~n25732;
  assign n19778 = ~n20624 & ~n25725;
  assign n19774 = ~n20376 & ~n25666;
  assign n19772 = ~n25706 | ~n19771;
  assign n20086 = ~P3_REG3_REG_18__SCAN_IN | ~P3_U3151;
  assign n19773 = ~n19772 | ~n20086;
  assign n19776 = ~n19774 & ~n19773;
  assign n19775 = ~n25734 | ~n20381;
  assign n19777 = ~n19776 | ~n19775;
  assign n19779 = ~n19778 & ~n19777;
  assign P3_U3178 = ~n19780 | ~n19779;
  assign n19791 = ~n19781 | ~n25732;
  assign n19789 = ~n20560 & ~n25725;
  assign n19787 = ~n20186 & ~n25666;
  assign n19783 = ~n26436 | ~n25706;
  assign n19782 = ~P3_REG3_REG_26__SCAN_IN | ~P3_U3151;
  assign n19785 = n19783 & n19782;
  assign n19784 = ~n20198 | ~n25734;
  assign n19786 = ~n19785 | ~n19784;
  assign n19788 = n19787 | n19786;
  assign n19790 = ~n19789 & ~n19788;
  assign P3_U3180 = ~n19791 | ~n19790;
  assign n19794 = n19793 ^ ~n19792;
  assign n19804 = ~n19794 | ~n25732;
  assign n19802 = ~n20648 & ~n25725;
  assign n19800 = ~n25734 | ~n20444;
  assign n19796 = ~n25728 | ~n19795;
  assign n19956 = ~P3_REG3_REG_15__SCAN_IN | ~P3_U3151;
  assign n19798 = ~n19796 | ~n19956;
  assign n19797 = ~n25724 & ~n20472;
  assign n19799 = ~n19798 & ~n19797;
  assign n19801 = ~n19800 | ~n19799;
  assign n19803 = ~n19802 & ~n19801;
  assign P3_U3181 = ~n19804 | ~n19803;
  assign n19805 = ~P3_REG1_REG_0__SCAN_IN;
  assign n25742 = P3_IR_REG_0__SCAN_IN | n19805;
  assign n19807 = ~n19806 | ~P3_REG1_REG_0__SCAN_IN;
  assign n25778 = ~n19967;
  assign n19808 = ~n25778 | ~P3_REG1_REG_2__SCAN_IN;
  assign n19970 = ~n25811;
  assign n19810 = ~n19809 | ~n19970;
  assign n25820 = n19972 ^ ~P3_REG1_REG_4__SCAN_IN;
  assign n25832 = ~n19972;
  assign n19812 = ~n25832 | ~P3_REG1_REG_4__SCAN_IN;
  assign n19974 = ~n25850;
  assign n19814 = ~n19813 | ~n19974;
  assign n25859 = P3_REG1_REG_6__SCAN_IN ^ n25875;
  assign n19815 = ~n25875 | ~P3_REG1_REG_6__SCAN_IN;
  assign n19979 = ~n25893;
  assign n19817 = ~n19816 | ~n19979;
  assign n25903 = n25916 ^ P3_REG1_REG_8__SCAN_IN;
  assign n19818 = ~n25916 | ~P3_REG1_REG_8__SCAN_IN;
  assign n25923 = ~n19984;
  assign n19820 = ~n19819 | ~n25923;
  assign n25942 = n19987 ^ ~P3_REG1_REG_10__SCAN_IN;
  assign n25955 = ~n19987;
  assign n19821 = ~n25955 | ~P3_REG1_REG_10__SCAN_IN;
  assign n25966 = ~n19989;
  assign n19823 = ~n19822 | ~n25966;
  assign n25986 = ~n19824 | ~n19823;
  assign n19825 = ~P3_REG1_REG_12__SCAN_IN;
  assign n25985 = n25988 ^ ~n19825;
  assign n19826 = ~n25988 | ~P3_REG1_REG_12__SCAN_IN;
  assign n26017 = ~n19993;
  assign n19828 = ~n19827 | ~n26017;
  assign n26026 = n19997 ^ ~P3_REG1_REG_14__SCAN_IN;
  assign n19830 = ~n26036 | ~P3_REG1_REG_14__SCAN_IN;
  assign n19837 = P3_REG1_REG_15__SCAN_IN ^ n20006;
  assign n19833 = n19832 | n19831;
  assign n19955 = ~n19833 | ~P3_STATE_REG_SCAN_IN;
  assign n19836 = ~n19835 | ~n19834;
  assign n19953 = ~n19836 | ~n18258;
  assign n20002 = ~n19955 & ~n19953;
  assign n20078 = ~n19868;
  assign n25741 = ~n20002 | ~n20078;
  assign n19963 = ~n19837 & ~n25741;
  assign n19839 = ~n19847 | ~P3_REG1_REG_1__SCAN_IN;
  assign n19838 = n19847 | n13874;
  assign n19841 = ~n13286 | ~n25773;
  assign n19885 = ~n19868;
  assign n19843 = ~n19885 | ~P3_REG1_REG_0__SCAN_IN;
  assign n26300 = ~P3_REG2_REG_0__SCAN_IN;
  assign n19842 = n19847 | n26300;
  assign n25751 = ~n19843 | ~n19842;
  assign n25750 = ~P3_IR_REG_0__SCAN_IN;
  assign n25789 = ~n19845 | ~n19844;
  assign n19849 = ~n19885 | ~P3_REG1_REG_2__SCAN_IN;
  assign n19846 = ~P3_REG2_REG_2__SCAN_IN;
  assign n19848 = n19847 | n19846;
  assign n19850 = n19849 & n19848;
  assign n19853 = ~n19850 | ~n19967;
  assign n19851 = ~n19850;
  assign n19852 = ~n19851 | ~n25778;
  assign n25790 = n19853 & n19852;
  assign n19854 = ~n25789 | ~n25790;
  assign n25807 = ~n19854 | ~n19853;
  assign n19856 = ~n19885 | ~P3_REG1_REG_3__SCAN_IN;
  assign n19855 = n20078 | n13965;
  assign n19857 = n19856 & n19855;
  assign n19860 = ~n19857 | ~n25811;
  assign n19858 = ~n19857;
  assign n19859 = ~n19858 | ~n19970;
  assign n25806 = n19859 & n19860;
  assign n25809 = ~n25807 | ~n25806;
  assign n25829 = ~n25809 | ~n19860;
  assign n19862 = ~n19885 | ~P3_REG1_REG_4__SCAN_IN;
  assign n26216 = ~P3_REG2_REG_4__SCAN_IN;
  assign n19861 = n20078 | n26216;
  assign n19863 = n19862 & n19861;
  assign n19866 = ~n19863 | ~n19972;
  assign n19864 = ~n19863;
  assign n19865 = ~n19864 | ~n25832;
  assign n25830 = n19866 & n19865;
  assign n19867 = ~n25829 | ~n25830;
  assign n19870 = ~n20078 | ~n13743;
  assign n19869 = n20078 | P3_REG2_REG_5__SCAN_IN;
  assign n19871 = ~n19870 | ~n19869;
  assign n25846 = n19871 & n25850;
  assign n19873 = ~n20078 | ~P3_REG1_REG_5__SCAN_IN;
  assign n26178 = ~P3_REG2_REG_5__SCAN_IN;
  assign n19872 = n19885 | n26178;
  assign n19874 = ~n19873 | ~n19872;
  assign n25845 = ~n19874 | ~n19974;
  assign n19876 = ~n19885 | ~P3_REG1_REG_6__SCAN_IN;
  assign n26155 = ~P3_REG2_REG_6__SCAN_IN;
  assign n19875 = n20078 | n26155;
  assign n19877 = ~n19876 | ~n19875;
  assign n25870 = n19877 & n25875;
  assign n19878 = ~P3_REG1_REG_6__SCAN_IN;
  assign n19880 = ~n19885 | ~n19878;
  assign n19879 = n19885 | P3_REG2_REG_6__SCAN_IN;
  assign n19882 = ~n19880 | ~n19879;
  assign n19881 = ~n25875;
  assign n25869 = ~n19882 | ~n19881;
  assign n25889 = ~n19883 | ~n25869;
  assign n19887 = ~n20078 | ~P3_REG1_REG_7__SCAN_IN;
  assign n19884 = ~P3_REG2_REG_7__SCAN_IN;
  assign n19886 = n19885 | n19884;
  assign n19888 = n19887 & n19886;
  assign n19891 = ~n19888 | ~n25893;
  assign n19889 = ~n19888;
  assign n19890 = ~n19889 | ~n19979;
  assign n25888 = n19891 & n19890;
  assign n25891 = ~n25889 | ~n25888;
  assign n25913 = ~n25891 | ~n19891;
  assign n19894 = ~n19885 | ~P3_REG1_REG_8__SCAN_IN;
  assign n19892 = ~P3_REG2_REG_8__SCAN_IN;
  assign n19893 = n20078 | n19892;
  assign n19896 = n19894 & n19893;
  assign n19895 = ~n25916;
  assign n19899 = ~n19896 | ~n19895;
  assign n19897 = ~n19896;
  assign n19898 = ~n19897 | ~n25916;
  assign n25914 = n19899 & n19898;
  assign n19900 = ~n25913 | ~n25914;
  assign n19901 = ~P3_REG1_REG_9__SCAN_IN;
  assign n19903 = ~n20078 | ~n19901;
  assign n19902 = n20078 | P3_REG2_REG_9__SCAN_IN;
  assign n19904 = ~n19903 | ~n19902;
  assign n25931 = n19904 & n19984;
  assign n19906 = ~n20078 | ~P3_REG1_REG_9__SCAN_IN;
  assign n26093 = ~P3_REG2_REG_9__SCAN_IN;
  assign n19905 = n20078 | n26093;
  assign n19907 = ~n19906 | ~n19905;
  assign n25930 = ~n19907 | ~n25923;
  assign n19909 = ~n20078 | ~P3_REG1_REG_10__SCAN_IN;
  assign n26066 = ~P3_REG2_REG_10__SCAN_IN;
  assign n19908 = n20078 | n26066;
  assign n19910 = n19909 & n19908;
  assign n19913 = ~n19910 | ~n19987;
  assign n19911 = ~n19910;
  assign n19912 = ~n19911 | ~n25955;
  assign n25948 = n19913 & n19912;
  assign n19916 = ~n20078 | ~P3_REG1_REG_11__SCAN_IN;
  assign n19914 = ~P3_REG2_REG_11__SCAN_IN;
  assign n19915 = n20078 | n19914;
  assign n19917 = ~n19916 | ~n19915;
  assign n25973 = n19917 ^ ~n19989;
  assign n19920 = ~n25974 | ~n25973;
  assign n19918 = ~n19917;
  assign n19919 = ~n19918 | ~n19989;
  assign n19921 = ~n25985;
  assign n19923 = ~n20078 | ~n19921;
  assign n20504 = ~P3_REG2_REG_12__SCAN_IN;
  assign n25982 = n25988 ^ ~n20504;
  assign n19922 = n20078 | n25982;
  assign n25996 = ~n19923 | ~n19922;
  assign n19925 = ~n20078 | ~P3_REG1_REG_12__SCAN_IN;
  assign n19924 = n20078 | n20504;
  assign n19926 = ~n19925 | ~n19924;
  assign n19927 = ~n19926 | ~n25988;
  assign n19929 = ~n20078 | ~P3_REG1_REG_13__SCAN_IN;
  assign n26007 = ~P3_REG2_REG_13__SCAN_IN;
  assign n19928 = n20078 | n26007;
  assign n19930 = ~n19929 | ~n19928;
  assign n26011 = n19930 ^ ~n19993;
  assign n19931 = ~n19930;
  assign n19932 = ~n19931 | ~n19993;
  assign n26029 = n19997 ^ ~P3_REG2_REG_14__SCAN_IN;
  assign n19934 = n26029 | n20078;
  assign n19933 = n26026 | n19868;
  assign n26042 = n19934 & n19933;
  assign n19937 = ~n20078 | ~P3_REG1_REG_14__SCAN_IN;
  assign n19935 = ~P3_REG2_REG_14__SCAN_IN;
  assign n19936 = n20078 | n19935;
  assign n19938 = ~n19937 | ~n19936;
  assign n19939 = ~n19938 | ~n26036;
  assign n20010 = ~n19940 | ~n19999;
  assign n20030 = ~n19999;
  assign n19942 = ~n19941 | ~n20030;
  assign n19945 = ~n20078 | ~P3_REG1_REG_15__SCAN_IN;
  assign n19943 = ~P3_REG2_REG_15__SCAN_IN;
  assign n19944 = n20078 | n19943;
  assign n19946 = ~n19945 | ~n19944;
  assign n19948 = ~n19947 | ~n19946;
  assign n19949 = ~n13380 | ~n19948;
  assign n19961 = ~n19949 | ~n26013;
  assign n19952 = ~n20002 | ~n20773;
  assign n19951 = ~P3_U3897 | ~n19950;
  assign n25894 = ~n19952 | ~n19951;
  assign n26037 = ~n25894;
  assign n19959 = ~n26037 & ~n20030;
  assign n19954 = ~n19953;
  assign n26033 = ~n19955 & ~n19954;
  assign n19957 = ~n26033 | ~P3_ADDR_REG_15__SCAN_IN;
  assign n19958 = ~n19957 | ~n19956;
  assign n19960 = ~n19959 & ~n19958;
  assign n19962 = ~n19961 | ~n19960;
  assign n20005 = ~n19963 & ~n19962;
  assign n25746 = ~P3_IR_REG_0__SCAN_IN & ~n26300;
  assign n19965 = ~n19964 & ~n26300;
  assign n19966 = ~n19965;
  assign n25782 = n19967 ^ ~P3_REG2_REG_2__SCAN_IN;
  assign n19969 = ~n25783 | ~n25782;
  assign n19968 = ~n25778 | ~P3_REG2_REG_2__SCAN_IN;
  assign n25822 = n19972 ^ ~P3_REG2_REG_4__SCAN_IN;
  assign n19973 = ~n25832 | ~P3_REG2_REG_4__SCAN_IN;
  assign n19976 = ~n19975 | ~n19974;
  assign n25862 = P3_REG2_REG_6__SCAN_IN ^ n25875;
  assign n19978 = ~n25875 | ~P3_REG2_REG_6__SCAN_IN;
  assign n19982 = ~n25882 | ~P3_REG2_REG_7__SCAN_IN;
  assign n19981 = ~n19980 | ~n19979;
  assign n25907 = ~n19982 | ~n19981;
  assign n25906 = P3_REG2_REG_8__SCAN_IN ^ n25916;
  assign n19983 = ~n25916 | ~P3_REG2_REG_8__SCAN_IN;
  assign n19986 = ~n19985 | ~n25923;
  assign n25946 = n19987 ^ ~P3_REG2_REG_10__SCAN_IN;
  assign n19988 = ~n25955 | ~P3_REG2_REG_10__SCAN_IN;
  assign n19991 = ~n19990 | ~n25966;
  assign n19992 = ~n25988 | ~P3_REG2_REG_12__SCAN_IN;
  assign n26008 = n19994 ^ ~n19993;
  assign n19996 = ~n26008 | ~P3_REG2_REG_13__SCAN_IN;
  assign n19995 = ~n19994 | ~n26017;
  assign n19998 = ~n26030 | ~P3_REG2_REG_14__SCAN_IN;
  assign n20003 = n20029 ^ ~P3_REG2_REG_15__SCAN_IN;
  assign n20001 = ~n20000;
  assign n20004 = ~n20003 | ~n26031;
  assign P3_U3197 = ~n20005 | ~n20004;
  assign n20038 = n20034 ^ ~P3_REG1_REG_16__SCAN_IN;
  assign n20008 = ~n20007 | ~n20030;
  assign n20009 = n20038 ^ n20039;
  assign n20028 = ~n20009 & ~n25741;
  assign n20013 = ~n20078 | ~P3_REG1_REG_16__SCAN_IN;
  assign n20011 = ~P3_REG2_REG_16__SCAN_IN;
  assign n20012 = n20078 | n20011;
  assign n20014 = ~n20013 | ~n20012;
  assign n20046 = ~n20014 | ~n20059;
  assign n20015 = ~P3_REG1_REG_16__SCAN_IN;
  assign n20017 = ~n20078 | ~n20015;
  assign n20016 = n20078 | P3_REG2_REG_16__SCAN_IN;
  assign n20018 = ~n20017 | ~n20016;
  assign n20045 = ~n20018 | ~n20034;
  assign n20019 = ~n20046 | ~n20045;
  assign n20020 = n13186 ^ ~n20019;
  assign n20026 = ~n20020 | ~n26013;
  assign n20021 = ~n26033 | ~P3_ADDR_REG_16__SCAN_IN;
  assign n20024 = ~n20022 | ~n20021;
  assign n20023 = ~n26037 & ~n20059;
  assign n20025 = ~n20024 & ~n20023;
  assign n20027 = ~n20026 | ~n20025;
  assign n20037 = ~n20028 & ~n20027;
  assign n20032 = ~n20031 | ~n20030;
  assign n20058 = ~n20033 | ~n20032;
  assign n20057 = n20034 ^ ~P3_REG2_REG_16__SCAN_IN;
  assign n20035 = n20058 ^ ~n20057;
  assign n20036 = ~n20035 | ~n26031;
  assign P3_U3198 = ~n20037 | ~n20036;
  assign n20040 = ~n20059 | ~P3_REG1_REG_16__SCAN_IN;
  assign n20041 = P3_REG1_REG_17__SCAN_IN ^ n20065;
  assign n20056 = ~n20041 & ~n25741;
  assign n20044 = ~n20078 | ~P3_REG1_REG_17__SCAN_IN;
  assign n20042 = ~P3_REG2_REG_17__SCAN_IN;
  assign n20043 = n20078 | n20042;
  assign n20071 = n20044 & n20043;
  assign n20069 = n20071 ^ ~n20094;
  assign n20047 = ~n13186 | ~n20045;
  assign n20070 = ~n20047 | ~n20046;
  assign n20048 = n20069 ^ n20070;
  assign n20054 = ~n20048 | ~n26013;
  assign n20049 = ~n26033 | ~P3_ADDR_REG_17__SCAN_IN;
  assign n20052 = ~n20050 | ~n20049;
  assign n20051 = ~n26037 & ~n20094;
  assign n20053 = ~n20052 & ~n20051;
  assign n20055 = ~n20054 | ~n20053;
  assign n20064 = ~n20056 & ~n20055;
  assign n20061 = ~n20058 | ~n20057;
  assign n20060 = ~n20059 | ~P3_REG2_REG_16__SCAN_IN;
  assign n20063 = ~n20062 | ~n26031;
  assign P3_U3199 = ~n20064 | ~n20063;
  assign n20104 = P3_REG1_REG_18__SCAN_IN ^ n20106;
  assign n20067 = ~n20066 | ~n20094;
  assign n20068 = n20104 ^ n20105;
  assign n20093 = ~n20068 & ~n25741;
  assign n20074 = ~n20070 | ~n20069;
  assign n20072 = ~n20071;
  assign n20073 = ~n20094 | ~n20072;
  assign n20075 = ~n20106;
  assign n20077 = ~n20076 | ~n20106;
  assign n20080 = ~n19868 | ~P3_REG2_REG_18__SCAN_IN;
  assign n20079 = ~n20078 | ~P3_REG1_REG_18__SCAN_IN;
  assign n20081 = ~n20080 | ~n20079;
  assign n20084 = ~n20110;
  assign n20083 = ~n20082 | ~n20081;
  assign n20085 = ~n20084 | ~n20083;
  assign n20091 = ~n20085 | ~n26013;
  assign n20089 = ~n26037 & ~n20106;
  assign n20087 = ~n26033 | ~P3_ADDR_REG_18__SCAN_IN;
  assign n20088 = ~n20087 | ~n20086;
  assign n20090 = ~n20089 & ~n20088;
  assign n20092 = ~n20091 | ~n20090;
  assign n20100 = ~n20093 & ~n20092;
  assign n20096 = ~n20095 | ~n20094;
  assign n20101 = P3_REG2_REG_18__SCAN_IN ^ n20106;
  assign n20098 = n20102 ^ ~n20101;
  assign n20099 = ~n20098 | ~n26031;
  assign P3_U3200 = ~n20100 | ~n20099;
  assign n20103 = ~n20106 | ~P3_REG2_REG_18__SCAN_IN;
  assign n20111 = n20119 ^ ~n20366;
  assign n20107 = ~n20106 | ~P3_REG1_REG_18__SCAN_IN;
  assign n20113 = n20119 ^ ~P3_REG1_REG_19__SCAN_IN;
  assign n20109 = ~n20108;
  assign n20112 = ~n20111;
  assign n20115 = ~n19868 | ~n20112;
  assign n20114 = ~n20078 | ~n20113;
  assign n20116 = ~n20115 | ~n20114;
  assign n20118 = n20117 ^ ~n20116;
  assign n20125 = ~n20118 | ~n26013;
  assign n20123 = ~n26037 & ~n20119;
  assign n20121 = ~n26033 | ~P3_ADDR_REG_19__SCAN_IN;
  assign n20122 = ~n20121 | ~n20120;
  assign n20124 = ~n20123 & ~n20122;
  assign n20126 = ~n20125 | ~n20124;
  assign n20136 = ~n20535 | ~n26297;
  assign n20132 = ~n20540;
  assign n20133 = ~n20132 & ~n20131;
  assign n20138 = ~n20133 | ~n20481;
  assign n20134 = n20481 | P3_REG2_REG_31__SCAN_IN;
  assign n20135 = ~n20138 | ~n20134;
  assign P3_U3202 = ~n20136 | ~n20135;
  assign n20140 = ~n20539 | ~n26297;
  assign n20137 = n20481 | P3_REG2_REG_30__SCAN_IN;
  assign n20139 = ~n20138 | ~n20137;
  assign P3_U3203 = ~n20140 | ~n20139;
  assign n20143 = ~n20142 & ~n20141;
  assign n20146 = ~n20143 & ~n26129;
  assign n20145 = ~n20144;
  assign n20151 = ~n20146 | ~n20145;
  assign n20149 = ~n20186 & ~n26137;
  assign n20148 = ~n26126 & ~n20147;
  assign n20150 = ~n20149 & ~n20148;
  assign n20545 = ~n20151 | ~n20150;
  assign n20153 = ~n26152 | ~n20152;
  assign n20154 = ~n20481 | ~n20153;
  assign n20157 = ~n20545 & ~n20154;
  assign n20156 = ~n20546 | ~n20388;
  assign n20159 = ~n20157 | ~n20156;
  assign n20158 = n20481 | P3_REG2_REG_28__SCAN_IN;
  assign n20162 = ~n20159 | ~n20158;
  assign n20161 = ~n20160 | ~n26297;
  assign P3_U3205 = ~n20162 | ~n20161;
  assign n20173 = n20164 ^ ~n20163;
  assign n20169 = ~n20173 | ~n26282;
  assign n20167 = ~n20209 & ~n26137;
  assign n20166 = ~n26126 & ~n20165;
  assign n20168 = ~n20167 & ~n20166;
  assign n20170 = ~n20169 | ~n20168;
  assign n20172 = ~n20556 | ~n20481;
  assign n20171 = n20481 | P3_REG2_REG_27__SCAN_IN;
  assign n20181 = ~n20172 | ~n20171;
  assign n20551 = ~n20173;
  assign n26228 = ~n26249;
  assign n26274 = ~n20481 | ~n26228;
  assign n20179 = ~n20551 & ~n26274;
  assign n20177 = ~n20174 | ~n26297;
  assign n20176 = ~n20175 | ~n26152;
  assign n20178 = ~n20177 | ~n20176;
  assign n20180 = ~n20179 & ~n20178;
  assign P3_U3206 = ~n20181 | ~n20180;
  assign n20183 = n20182 ^ n20184;
  assign n20192 = ~n20183 & ~n26129;
  assign n20196 = n20185 ^ ~n20184;
  assign n20190 = ~n20196 | ~n26282;
  assign n20188 = ~n20186 & ~n26126;
  assign n20187 = ~n20235 & ~n26137;
  assign n20189 = ~n20188 & ~n20187;
  assign n20191 = ~n20190 | ~n20189;
  assign n20564 = ~n20192 & ~n20191;
  assign n20195 = ~n20564 | ~n20481;
  assign n20194 = ~n26270 | ~n20193;
  assign n20204 = ~n20195 | ~n20194;
  assign n20559 = ~n20196;
  assign n20202 = ~n20559 & ~n26274;
  assign n20200 = ~n20197 | ~n26297;
  assign n20199 = ~n20198 | ~n26152;
  assign n20201 = ~n20200 | ~n20199;
  assign n20203 = ~n20202 & ~n20201;
  assign P3_U3207 = ~n20204 | ~n20203;
  assign n20216 = ~n20206 & ~n26129;
  assign n20219 = n20207 ^ ~n20208;
  assign n20214 = ~n20219 | ~n26282;
  assign n20212 = ~n20209 & ~n26126;
  assign n20211 = ~n20210 & ~n26137;
  assign n20213 = ~n20212 & ~n20211;
  assign n20215 = ~n20214 | ~n20213;
  assign n20572 = ~n20216 & ~n20215;
  assign n20218 = ~n20572 | ~n20481;
  assign n20217 = n20481 | P3_REG2_REG_25__SCAN_IN;
  assign n20227 = ~n20218 | ~n20217;
  assign n20567 = ~n20219;
  assign n20225 = ~n20567 & ~n26274;
  assign n20223 = ~n20220 | ~n26297;
  assign n20222 = ~n20221 | ~n26152;
  assign n20224 = ~n20223 | ~n20222;
  assign n20226 = ~n20225 & ~n20224;
  assign P3_U3208 = ~n20227 | ~n20226;
  assign n20230 = ~n20254 | ~n20228;
  assign n20231 = ~n20230 | ~n20229;
  assign n20232 = n20233 ^ n20231;
  assign n20241 = ~n20232 & ~n26129;
  assign n20244 = n20234 ^ ~n20233;
  assign n20239 = ~n20244 | ~n26282;
  assign n20237 = ~n20235 & ~n26126;
  assign n20236 = ~n20287 & ~n26137;
  assign n20238 = ~n20237 & ~n20236;
  assign n20240 = ~n20239 | ~n20238;
  assign n20579 = ~n20241 & ~n20240;
  assign n20243 = ~n20579 | ~n20481;
  assign n20242 = n20481 | P3_REG2_REG_24__SCAN_IN;
  assign n20252 = ~n20243 | ~n20242;
  assign n20575 = ~n20244;
  assign n20250 = ~n20575 & ~n26274;
  assign n20248 = ~n20245 | ~n26297;
  assign n20247 = ~n20246 | ~n26152;
  assign n20249 = ~n20248 | ~n20247;
  assign n20251 = ~n20250 & ~n20249;
  assign P3_U3209 = ~n20252 | ~n20251;
  assign n20255 = n20254 & n20253;
  assign n20256 = n20255 ^ ~n19465;
  assign n20270 = ~n20256 | ~n26280;
  assign n20262 = ~n20293 | ~n20260;
  assign n20264 = ~n20262 | ~n20261;
  assign n20265 = ~n20264 | ~n20263;
  assign n20582 = ~n13934 | ~n20265;
  assign n20269 = ~n20266 | ~n18385;
  assign n20268 = ~n20267 | ~n26288;
  assign n20272 = ~n20589 & ~n26270;
  assign n20271 = ~n20481 & ~P3_REG2_REG_23__SCAN_IN;
  assign n20279 = n20272 | n20271;
  assign n20277 = ~n20582 & ~n26274;
  assign n20275 = ~n20585 | ~n26297;
  assign n20274 = ~n20273 | ~n26152;
  assign n20276 = ~n20275 | ~n20274;
  assign n20278 = ~n20277 & ~n20276;
  assign P3_U3210 = ~n20279 | ~n20278;
  assign n20328 = ~n20281 | ~n20280;
  assign n20284 = ~n20328 | ~n20282;
  assign n20285 = ~n20284 | ~n20283;
  assign n20286 = n20292 ^ n20285;
  assign n20291 = ~n20286 | ~n26280;
  assign n20289 = ~n20287 & ~n26126;
  assign n20288 = ~n20334 & ~n26137;
  assign n20290 = ~n20289 & ~n20288;
  assign n20295 = ~n20291 | ~n20290;
  assign n20592 = n20293 ^ ~n20292;
  assign n20294 = ~n20592 & ~n20501;
  assign n20597 = ~n20295 & ~n20294;
  assign n20297 = ~n20597 | ~n20481;
  assign n20296 = n20481 | P3_REG2_REG_22__SCAN_IN;
  assign n20305 = ~n20297 | ~n20296;
  assign n20303 = ~n20592 & ~n26274;
  assign n20301 = ~n20298 | ~n26297;
  assign n20300 = ~n20299 | ~n26152;
  assign n20302 = ~n20301 | ~n20300;
  assign n20304 = ~n20303 & ~n20302;
  assign P3_U3211 = ~n20305 | ~n20304;
  assign n20307 = ~n20328 | ~n20330;
  assign n20308 = ~n20307 | ~n20306;
  assign n20309 = n20308 ^ ~n13190;
  assign n20314 = ~n20309 | ~n26280;
  assign n20312 = ~n20310 & ~n26126;
  assign n20311 = ~n20354 & ~n26137;
  assign n20313 = ~n20312 & ~n20311;
  assign n20318 = ~n20314 | ~n20313;
  assign n20316 = ~n20333 | ~n20315;
  assign n20600 = n20316 ^ ~n13190;
  assign n20317 = ~n20600 & ~n20501;
  assign n20605 = ~n20318 & ~n20317;
  assign n20320 = ~n20605 | ~n20481;
  assign n20319 = n20481 | P3_REG2_REG_21__SCAN_IN;
  assign n20327 = ~n20320 | ~n20319;
  assign n20325 = ~n20600 & ~n26274;
  assign n20323 = ~n18431 | ~n26297;
  assign n20322 = ~n20321 | ~n26152;
  assign n20324 = ~n20323 | ~n20322;
  assign n20326 = ~n20325 & ~n20324;
  assign P3_U3212 = ~n20327 | ~n20326;
  assign n20329 = n20328 ^ ~n20330;
  assign n20340 = ~n20329 & ~n26129;
  assign n20332 = ~n20331 | ~n20330;
  assign n20341 = n20333 & n20332;
  assign n20338 = ~n20341 | ~n26282;
  assign n20336 = ~n20334 & ~n26126;
  assign n20335 = ~n20376 & ~n26137;
  assign n20337 = ~n20336 & ~n20335;
  assign n20339 = ~n20338 | ~n20337;
  assign n20613 = ~n20340 & ~n20339;
  assign n20608 = ~n20341;
  assign n20345 = ~n20608 & ~n26249;
  assign n20343 = ~n20342 | ~n26152;
  assign n20344 = ~n20343 | ~n20481;
  assign n20346 = ~n20345 & ~n20344;
  assign n20348 = ~n20613 | ~n20346;
  assign n20347 = n20481 | P3_REG2_REG_20__SCAN_IN;
  assign n20351 = ~n20348 | ~n20347;
  assign n20350 = ~n20349 | ~n26297;
  assign P3_U3213 = ~n20351 | ~n20350;
  assign n20353 = n20352 ^ n20362;
  assign n20358 = ~n20353 | ~n26280;
  assign n20356 = ~n20354 & ~n26126;
  assign n20355 = ~n20398 & ~n26137;
  assign n20357 = ~n20356 & ~n20355;
  assign n20618 = ~n20358 | ~n20357;
  assign n20360 = ~n20359 | ~n26152;
  assign n20361 = ~n20360 | ~n20481;
  assign n20365 = ~n20618 & ~n20361;
  assign n20619 = n20363 ^ n20362;
  assign n20364 = ~n20619 | ~n20388;
  assign n20368 = ~n20365 | ~n20364;
  assign n20367 = ~n26270 | ~n20366;
  assign n20371 = ~n20368 | ~n20367;
  assign n20370 = ~n20369 | ~n26297;
  assign P3_U3214 = ~n20371 | ~n20370;
  assign n20373 = n20372 | n20385;
  assign n20375 = ~n20374 | ~n20373;
  assign n20380 = ~n20375 | ~n26280;
  assign n20378 = ~n20376 & ~n26126;
  assign n20377 = ~n20416 & ~n26137;
  assign n20379 = ~n20378 & ~n20377;
  assign n20626 = ~n20380 | ~n20379;
  assign n20382 = ~n20381 | ~n26152;
  assign n20383 = ~n20382 | ~n20481;
  assign n20390 = ~n20626 & ~n20383;
  assign n20386 = ~n20384 | ~n20385;
  assign n20389 = ~n20627 | ~n20388;
  assign n20393 = ~n20390 | ~n20389;
  assign n20392 = ~n26270 | ~n20391;
  assign n20395 = ~n20393 | ~n20392;
  assign n20394 = ~n19427 | ~n26297;
  assign P3_U3215 = ~n20395 | ~n20394;
  assign n20397 = n20396 ^ ~n14709;
  assign n20402 = ~n20397 | ~n26280;
  assign n20400 = ~n20398 & ~n26126;
  assign n20399 = ~n20435 & ~n26137;
  assign n20401 = ~n20400 & ~n20399;
  assign n20634 = ~n20402 | ~n20401;
  assign n20404 = ~n20634 & ~n26270;
  assign n20403 = ~n20481 & ~P3_REG2_REG_17__SCAN_IN;
  assign n20413 = n20404 | n20403;
  assign n20635 = n20405 ^ ~n20406;
  assign n20411 = n20635 & n20526;
  assign n20409 = n20632 | n26224;
  assign n20408 = ~n20407 | ~n26152;
  assign n20410 = ~n20409 | ~n20408;
  assign n20412 = ~n20411 & ~n20410;
  assign P3_U3216 = ~n20413 | ~n20412;
  assign n20415 = n20414 ^ ~n20424;
  assign n20420 = ~n20415 | ~n26280;
  assign n20418 = ~n20416 & ~n26126;
  assign n20417 = ~n20454 & ~n26137;
  assign n20419 = ~n20418 & ~n20417;
  assign n20642 = ~n20420 | ~n20419;
  assign n20422 = ~n20642 & ~n26270;
  assign n20421 = ~n20481 & ~P3_REG2_REG_16__SCAN_IN;
  assign n20432 = ~n20422 & ~n20421;
  assign n20643 = n20423 ^ ~n20424;
  assign n20430 = ~n20643 | ~n20526;
  assign n20428 = ~n20640 & ~n26224;
  assign n20426 = ~n20425;
  assign n20427 = ~n20426 & ~n20528;
  assign n20429 = ~n20428 & ~n20427;
  assign n20431 = ~n20430 | ~n20429;
  assign P3_U3217 = n20432 | n20431;
  assign n20434 = n20433 ^ ~n20442;
  assign n20439 = ~n20434 | ~n26280;
  assign n20437 = ~n20435 & ~n26126;
  assign n20436 = ~n20472 & ~n26137;
  assign n20438 = ~n20437 & ~n20436;
  assign n20650 = ~n20439 | ~n20438;
  assign n20441 = ~n20650 & ~n26270;
  assign n20440 = ~n20481 & ~P3_REG2_REG_15__SCAN_IN;
  assign n20451 = ~n20441 & ~n20440;
  assign n20651 = n20443 ^ ~n20442;
  assign n20449 = ~n20651 | ~n20526;
  assign n20447 = ~n20648 & ~n26224;
  assign n20445 = ~n20444;
  assign n20446 = ~n20528 & ~n20445;
  assign n20448 = ~n20447 & ~n20446;
  assign n20450 = ~n20449 | ~n20448;
  assign P3_U3218 = n20451 | n20450;
  assign n20453 = n20452 ^ ~n20461;
  assign n20458 = ~n20453 | ~n26280;
  assign n20456 = ~n20454 & ~n26126;
  assign n20455 = ~n20495 & ~n26137;
  assign n20457 = ~n20456 & ~n20455;
  assign n20658 = ~n20458 | ~n20457;
  assign n20460 = ~n20658 & ~n26270;
  assign n20459 = ~n20481 & ~P3_REG2_REG_14__SCAN_IN;
  assign n20469 = n20460 | n20459;
  assign n20659 = n20462 ^ ~n20461;
  assign n20467 = n20659 & n20526;
  assign n20465 = n20656 | n26224;
  assign n20464 = ~n26152 | ~n20463;
  assign n20466 = ~n20465 | ~n20464;
  assign n20468 = ~n20467 & ~n20466;
  assign P3_U3219 = ~n20469 | ~n20468;
  assign n20471 = n20470 ^ ~n20477;
  assign n20476 = ~n20471 | ~n26280;
  assign n20474 = ~n26126 & ~n20472;
  assign n20473 = ~n20517 & ~n26137;
  assign n20475 = ~n20474 & ~n20473;
  assign n20480 = ~n20476 | ~n20475;
  assign n20664 = n20478 ^ n20477;
  assign n20479 = ~n20664 & ~n20501;
  assign n20669 = ~n20480 & ~n20479;
  assign n20483 = ~n20669 | ~n20481;
  assign n20482 = ~n26270 | ~n26007;
  assign n20491 = ~n20483 | ~n20482;
  assign n20489 = ~n20664 & ~n26274;
  assign n20487 = ~n20484 | ~n26297;
  assign n20486 = ~n26152 | ~n20485;
  assign n20488 = ~n20487 | ~n20486;
  assign n20490 = ~n20489 & ~n20488;
  assign P3_U3220 = ~n20491 | ~n20490;
  assign n20494 = n20492 ^ ~n20493;
  assign n20499 = ~n20494 | ~n26280;
  assign n20497 = ~n26126 & ~n20495;
  assign n20496 = ~n25611 & ~n26137;
  assign n20498 = ~n20497 & ~n20496;
  assign n20503 = ~n20499 | ~n20498;
  assign n20502 = ~n20672 & ~n20501;
  assign n20678 = ~n20503 & ~n20502;
  assign n20506 = ~n20678 | ~n20481;
  assign n20505 = ~n26270 | ~n20504;
  assign n20514 = ~n20506 | ~n20505;
  assign n20512 = ~n20672 & ~n26274;
  assign n20510 = ~n20507 | ~n26297;
  assign n20509 = ~n26152 | ~n20508;
  assign n20511 = ~n20510 | ~n20509;
  assign n20513 = ~n20512 & ~n20511;
  assign P3_U3221 = ~n20514 | ~n20513;
  assign n20516 = n20515 ^ ~n20524;
  assign n20521 = ~n20516 | ~n26280;
  assign n20519 = ~n26126 & ~n20517;
  assign n20518 = ~n25689 & ~n26137;
  assign n20520 = ~n20519 & ~n20518;
  assign n20683 = ~n20521 | ~n20520;
  assign n20523 = ~n20683 & ~n26270;
  assign n20522 = ~n20481 & ~P3_REG2_REG_11__SCAN_IN;
  assign n20534 = ~n20523 & ~n20522;
  assign n20685 = n20525 ^ ~n20524;
  assign n20532 = ~n20685 | ~n20526;
  assign n20530 = ~n20681 & ~n26224;
  assign n20527 = ~n25699;
  assign n20529 = ~n20528 & ~n20527;
  assign n20531 = ~n20530 & ~n20529;
  assign n20533 = ~n20532 | ~n20531;
  assign P3_U3222 = n20534 | n20533;
  assign n20536 = ~n20535 | ~n26315;
  assign n20690 = ~n20536 | ~n20540;
  assign n20538 = ~n20690 | ~n26433;
  assign n20537 = ~n26431 | ~P3_REG1_REG_31__SCAN_IN;
  assign P3_U3490 = ~n20538 | ~n20537;
  assign n20541 = ~n20539 | ~n26315;
  assign n20693 = ~n20541 | ~n20540;
  assign n20543 = ~n20693 | ~n26433;
  assign n20542 = ~n26431 | ~P3_REG1_REG_30__SCAN_IN;
  assign P3_U3489 = ~n20543 | ~n20542;
  assign n20544 = ~n14256 & ~n20673;
  assign n20548 = ~n20545 & ~n20544;
  assign n20547 = ~n20546 | ~n20684;
  assign n20696 = ~n20548 | ~n20547;
  assign n20550 = ~n20696 | ~n26433;
  assign n20549 = ~n26431 | ~P3_REG1_REG_28__SCAN_IN;
  assign P3_U3487 = ~n20550 | ~n20549;
  assign n20554 = ~n20551 & ~n26391;
  assign n20553 = ~n20552 & ~n20673;
  assign n20555 = ~n20554 & ~n20553;
  assign n20699 = ~n20556 | ~n20555;
  assign n20558 = ~n20699 | ~n26433;
  assign n20557 = ~n26431 | ~P3_REG1_REG_27__SCAN_IN;
  assign P3_U3486 = ~n20558 | ~n20557;
  assign n20562 = ~n20559 & ~n26391;
  assign n20561 = ~n20560 & ~n20673;
  assign n20563 = ~n20562 & ~n20561;
  assign n20702 = ~n20564 | ~n20563;
  assign n20566 = ~n20702 | ~n26433;
  assign n20565 = ~n26431 | ~P3_REG1_REG_26__SCAN_IN;
  assign P3_U3485 = ~n20566 | ~n20565;
  assign n20570 = ~n20567 & ~n26391;
  assign n20569 = ~n20568 & ~n20673;
  assign n20571 = ~n20570 & ~n20569;
  assign n20705 = ~n20572 | ~n20571;
  assign n20574 = ~n20705 | ~n26433;
  assign n20573 = ~n26431 | ~P3_REG1_REG_25__SCAN_IN;
  assign P3_U3484 = ~n20574 | ~n20573;
  assign n20577 = ~n20575 & ~n26391;
  assign n20576 = ~n18436 & ~n20673;
  assign n20578 = ~n20577 & ~n20576;
  assign n20708 = ~n20579 | ~n20578;
  assign n20581 = ~n20708 | ~n26433;
  assign n20580 = ~n26431 | ~P3_REG1_REG_24__SCAN_IN;
  assign P3_U3483 = ~n20581 | ~n20580;
  assign n20584 = ~n20582;
  assign n20583 = ~n26391;
  assign n20587 = ~n20584 | ~n20583;
  assign n20586 = ~n20585 | ~n26315;
  assign n20588 = ~n20587 | ~n20586;
  assign n20591 = ~n13193 | ~n26433;
  assign n20590 = ~n26431 | ~P3_REG1_REG_23__SCAN_IN;
  assign P3_U3482 = ~n20591 | ~n20590;
  assign n20595 = ~n20592 & ~n26391;
  assign n20594 = ~n20593 & ~n20673;
  assign n20596 = ~n20595 & ~n20594;
  assign n20713 = ~n20597 | ~n20596;
  assign n20599 = ~n20713 | ~n26433;
  assign n20598 = ~n26431 | ~P3_REG1_REG_22__SCAN_IN;
  assign P3_U3481 = ~n20599 | ~n20598;
  assign n20603 = ~n20600 & ~n26391;
  assign n20602 = ~n20601 & ~n20673;
  assign n20604 = ~n20603 & ~n20602;
  assign n20716 = ~n20605 | ~n20604;
  assign n20607 = ~n20716 | ~n26433;
  assign n20606 = ~n26431 | ~P3_REG1_REG_21__SCAN_IN;
  assign P3_U3480 = ~n20607 | ~n20606;
  assign n20611 = ~n20608 & ~n26391;
  assign n20610 = ~n20609 & ~n20673;
  assign n20612 = ~n20611 & ~n20610;
  assign n20719 = ~n20613 | ~n20612;
  assign n20615 = ~n20719 | ~n26433;
  assign n20614 = ~n26431 | ~P3_REG1_REG_20__SCAN_IN;
  assign P3_U3479 = ~n20615 | ~n20614;
  assign n20617 = ~n20616 & ~n20673;
  assign n20621 = ~n20618 & ~n20617;
  assign n20620 = ~n20619 | ~n20684;
  assign n20722 = ~n20621 | ~n20620;
  assign n20623 = ~n20722 | ~n26433;
  assign n20622 = ~n26431 | ~P3_REG1_REG_19__SCAN_IN;
  assign P3_U3478 = ~n20623 | ~n20622;
  assign n20625 = ~n20624 & ~n20673;
  assign n20629 = ~n20626 & ~n20625;
  assign n20628 = ~n20627 | ~n20684;
  assign n20725 = ~n20629 | ~n20628;
  assign n20631 = ~n20725 | ~n26433;
  assign n20630 = ~n26431 | ~P3_REG1_REG_18__SCAN_IN;
  assign P3_U3477 = ~n20631 | ~n20630;
  assign n20633 = ~n20632 & ~n20673;
  assign n20637 = ~n20634 & ~n20633;
  assign n20636 = ~n20635 | ~n20684;
  assign n20728 = ~n20637 | ~n20636;
  assign n20639 = ~n20728 | ~n26433;
  assign n20638 = ~n26431 | ~P3_REG1_REG_17__SCAN_IN;
  assign P3_U3476 = ~n20639 | ~n20638;
  assign n20641 = ~n20640 & ~n20673;
  assign n20645 = ~n20642 & ~n20641;
  assign n20644 = ~n20643 | ~n20684;
  assign n20731 = ~n20645 | ~n20644;
  assign n20647 = ~n20731 | ~n26433;
  assign n20646 = ~n26431 | ~P3_REG1_REG_16__SCAN_IN;
  assign P3_U3475 = ~n20647 | ~n20646;
  assign n20649 = ~n20648 & ~n20673;
  assign n20653 = ~n20650 & ~n20649;
  assign n20652 = ~n20651 | ~n20684;
  assign n20734 = ~n20653 | ~n20652;
  assign n20655 = ~n20734 | ~n26433;
  assign n20654 = ~n26431 | ~P3_REG1_REG_15__SCAN_IN;
  assign P3_U3474 = ~n20655 | ~n20654;
  assign n20657 = ~n20656 & ~n20673;
  assign n20661 = ~n20658 & ~n20657;
  assign n20660 = ~n20659 | ~n20684;
  assign n20737 = ~n20661 | ~n20660;
  assign n20663 = ~n20737 | ~n26433;
  assign n20662 = ~n26431 | ~P3_REG1_REG_14__SCAN_IN;
  assign P3_U3473 = ~n20663 | ~n20662;
  assign n20667 = ~n20664 & ~n26391;
  assign n20666 = ~n20665 & ~n20673;
  assign n20668 = ~n20667 & ~n20666;
  assign n20740 = ~n20669 | ~n20668;
  assign n20671 = ~n20740 | ~n26433;
  assign n20670 = ~n26431 | ~P3_REG1_REG_13__SCAN_IN;
  assign P3_U3472 = ~n20671 | ~n20670;
  assign n20676 = ~n20672 & ~n26391;
  assign n20675 = ~n20674 & ~n20673;
  assign n20677 = ~n20676 & ~n20675;
  assign n20743 = ~n20678 | ~n20677;
  assign n20680 = ~n20743 | ~n26433;
  assign n20679 = ~n26431 | ~P3_REG1_REG_12__SCAN_IN;
  assign P3_U3471 = ~n20680 | ~n20679;
  assign n20682 = ~n20681 & ~n20673;
  assign n20687 = ~n20683 & ~n20682;
  assign n20686 = ~n20685 | ~n20684;
  assign n20746 = ~n20687 | ~n20686;
  assign n20689 = ~n20746 | ~n26433;
  assign n20688 = ~n26431 | ~P3_REG1_REG_11__SCAN_IN;
  assign P3_U3470 = ~n20689 | ~n20688;
  assign n20692 = ~n20690 | ~n26398;
  assign n20691 = ~n26390 | ~P3_REG0_REG_31__SCAN_IN;
  assign P3_U3458 = ~n20692 | ~n20691;
  assign n20695 = ~n20693 | ~n26398;
  assign n20694 = ~n26390 | ~P3_REG0_REG_30__SCAN_IN;
  assign P3_U3457 = ~n20695 | ~n20694;
  assign n20698 = ~n20696 | ~n26398;
  assign n20697 = ~n26390 | ~P3_REG0_REG_28__SCAN_IN;
  assign P3_U3455 = ~n20698 | ~n20697;
  assign n20701 = ~n20699 | ~n26398;
  assign n20700 = ~n26390 | ~P3_REG0_REG_27__SCAN_IN;
  assign P3_U3454 = ~n20701 | ~n20700;
  assign n20704 = ~n20702 | ~n26398;
  assign n20703 = ~n26390 | ~P3_REG0_REG_26__SCAN_IN;
  assign P3_U3453 = ~n20704 | ~n20703;
  assign n20707 = ~n20705 | ~n26398;
  assign n20706 = ~n26390 | ~P3_REG0_REG_25__SCAN_IN;
  assign P3_U3452 = ~n20707 | ~n20706;
  assign n20710 = ~n20708 | ~n26398;
  assign n20709 = ~n26390 | ~P3_REG0_REG_24__SCAN_IN;
  assign P3_U3451 = ~n20710 | ~n20709;
  assign n20712 = ~n13193 | ~n26398;
  assign n20711 = ~n26390 | ~P3_REG0_REG_23__SCAN_IN;
  assign P3_U3450 = ~n20712 | ~n20711;
  assign n20715 = ~n20713 | ~n26398;
  assign n20714 = ~n26390 | ~P3_REG0_REG_22__SCAN_IN;
  assign P3_U3449 = ~n20715 | ~n20714;
  assign n20718 = ~n20716 | ~n26398;
  assign n20717 = ~n26390 | ~P3_REG0_REG_21__SCAN_IN;
  assign P3_U3448 = ~n20718 | ~n20717;
  assign n20721 = ~n20719 | ~n26398;
  assign n20720 = ~n26390 | ~P3_REG0_REG_20__SCAN_IN;
  assign P3_U3447 = ~n20721 | ~n20720;
  assign n20724 = ~n20722 | ~n26398;
  assign n20723 = ~n26390 | ~P3_REG0_REG_19__SCAN_IN;
  assign P3_U3446 = ~n20724 | ~n20723;
  assign n20727 = ~n20725 | ~n26398;
  assign n20726 = ~n26390 | ~P3_REG0_REG_18__SCAN_IN;
  assign P3_U3444 = ~n20727 | ~n20726;
  assign n20730 = ~n20728 | ~n26398;
  assign n20729 = ~n26390 | ~P3_REG0_REG_17__SCAN_IN;
  assign P3_U3441 = ~n20730 | ~n20729;
  assign n20733 = ~n20731 | ~n26398;
  assign n20732 = ~n26390 | ~P3_REG0_REG_16__SCAN_IN;
  assign P3_U3438 = ~n20733 | ~n20732;
  assign n20736 = ~n20734 | ~n26398;
  assign n20735 = ~n26390 | ~P3_REG0_REG_15__SCAN_IN;
  assign P3_U3435 = ~n20736 | ~n20735;
  assign n20739 = ~n20737 | ~n26398;
  assign n20738 = ~n26390 | ~P3_REG0_REG_14__SCAN_IN;
  assign P3_U3432 = ~n20739 | ~n20738;
  assign n20742 = ~n20740 | ~n26398;
  assign n20741 = ~n26390 | ~P3_REG0_REG_13__SCAN_IN;
  assign P3_U3429 = ~n20742 | ~n20741;
  assign n20745 = ~n20743 | ~n26398;
  assign n20744 = ~n26390 | ~P3_REG0_REG_12__SCAN_IN;
  assign P3_U3426 = ~n20745 | ~n20744;
  assign n20748 = ~n20746 | ~n26398;
  assign n20747 = ~n26390 | ~P3_REG0_REG_11__SCAN_IN;
  assign P3_U3423 = ~n20748 | ~n20747;
  assign n20757 = n20749 | n20792;
  assign n20750 = ~n16337 & ~P3_IR_REG_30__SCAN_IN;
  assign n20751 = ~n20750 | ~P3_STATE_REG_SCAN_IN;
  assign n20755 = ~n20752 & ~n20751;
  assign n20753 = ~SI_31_;
  assign n20754 = ~n20796 & ~n20753;
  assign n20756 = ~n20755 & ~n20754;
  assign P3_U3264 = ~n20757 | ~n20756;
  assign n20764 = n20758 | n20792;
  assign n20762 = ~n20759 & ~P3_U3151;
  assign n20761 = ~n20796 & ~n20760;
  assign n20763 = ~n20762 & ~n20761;
  assign P3_U3265 = ~n20764 | ~n20763;
  assign n20771 = n20765 | n20792;
  assign n20769 = ~n20766 & ~P3_U3151;
  assign n20768 = ~n20796 & ~n20767;
  assign n20770 = ~n20769 & ~n20768;
  assign P3_U3266 = ~n20771 | ~n20770;
  assign n20778 = ~n20772 & ~n20792;
  assign n20776 = n20773 | P3_U3151;
  assign n20775 = ~n20774 | ~SI_28_;
  assign n20777 = ~n20776 | ~n20775;
  assign P3_U3267 = n20778 | n20777;
  assign n20784 = n20779 | n20792;
  assign n20782 = ~n20078 & ~P3_U3151;
  assign n20781 = ~n20796 & ~n20780;
  assign n20783 = ~n20782 & ~n20781;
  assign P3_U3268 = ~n20784 | ~n20783;
  assign n20791 = n20785 | n20792;
  assign n20789 = ~n20786 & ~P3_U3151;
  assign n20788 = ~n20796 & ~n20787;
  assign n20790 = ~n20789 & ~n20788;
  assign P3_U3269 = ~n20791 | ~n20790;
  assign n20800 = n20793 | n20792;
  assign n20798 = ~n20794 & ~P3_U3151;
  assign n20797 = ~n20796 & ~n20795;
  assign n20799 = ~n20798 & ~n20797;
  assign P3_U3270 = ~n20800 | ~n20799;
  assign n20804 = ~n20801 | ~P3_U3151;
  assign n20803 = ~n20802 | ~P3_STATE_REG_SCAN_IN;
  assign P3_U3271 = ~n20804 | ~n20803;
  assign n20817 = ~n20806 | ~n24506;
  assign n20815 = ~n21497 & ~n21025;
  assign n20813 = ~n25583 | ~n24455;
  assign n21498 = ~n20807;
  assign n20811 = ~n24511 & ~n21498;
  assign n20809 = ~n24500 | ~n25577;
  assign n20808 = ~P2_REG3_REG_27__SCAN_IN | ~P2_U3088;
  assign n20810 = ~n20809 | ~n20808;
  assign n20812 = ~n20811 & ~n20810;
  assign n20814 = ~n20813 | ~n20812;
  assign n20816 = ~n20815 & ~n20814;
  assign P2_U3186 = ~n20817 | ~n20816;
  assign n20820 = ~n20818;
  assign n20902 = ~n20820 & ~n20819;
  assign n20822 = ~n20902;
  assign n20821 = ~n20820 | ~n20819;
  assign n20823 = ~n20822 | ~n20821;
  assign n20833 = ~n20823 | ~n24506;
  assign n20825 = ~n24484 & ~n24389;
  assign n24811 = ~P2_STATE_REG_SCAN_IN & ~n20824;
  assign n20827 = ~n20825 & ~n24811;
  assign n20826 = ~n24455 | ~n21818;
  assign n20829 = n20827 & n20826;
  assign n20828 = ~n24475 | ~n21831;
  assign n20831 = ~n20829 | ~n20828;
  assign n20830 = ~n21025 & ~n21830;
  assign n20832 = ~n20831 & ~n20830;
  assign P2_U3187 = ~n20833 | ~n20832;
  assign n20837 = ~n20834 | ~n20835;
  assign n20838 = n20837 ^ ~n20836;
  assign n20848 = ~n20838 | ~n24506;
  assign n20846 = ~n21598 & ~n21025;
  assign n20840 = ~n24455 | ~n25571;
  assign n20839 = ~P2_REG3_REG_23__SCAN_IN | ~P2_U3088;
  assign n20842 = ~n20840 | ~n20839;
  assign n20841 = ~n24484 & ~n21586;
  assign n20844 = ~n20842 & ~n20841;
  assign n20843 = ~n24475 | ~n21599;
  assign n20845 = ~n20844 | ~n20843;
  assign n20847 = ~n20846 & ~n20845;
  assign P2_U3188 = ~n20848 | ~n20847;
  assign n20852 = ~n20851 | ~n20850;
  assign n20853 = n20849 ^ ~n20852;
  assign n20862 = ~n20853 | ~n24506;
  assign n20860 = ~n14434 & ~n21025;
  assign n20854 = ~n24455 | ~n25559;
  assign n24915 = ~P2_REG3_REG_19__SCAN_IN | ~P2_U3088;
  assign n20856 = ~n20854 | ~n24915;
  assign n20855 = ~n24484 & ~n13885;
  assign n20858 = ~n20856 & ~n20855;
  assign n20857 = ~n24475 | ~n21695;
  assign n20859 = ~n20858 | ~n20857;
  assign n20861 = ~n20860 & ~n20859;
  assign P2_U3191 = ~n20862 | ~n20861;
  assign n20864 = ~n13388 | ~n20863;
  assign n20866 = n20865 ^ ~n20864;
  assign n20877 = ~n20866 | ~n24506;
  assign n20875 = ~n20867 & ~n21025;
  assign n20869 = ~n24455 | ~n25565;
  assign n20868 = ~P2_REG3_REG_21__SCAN_IN | ~P2_U3088;
  assign n20871 = ~n20869 | ~n20868;
  assign n20870 = ~n24484 & ~n21684;
  assign n20873 = ~n20871 & ~n20870;
  assign n20872 = ~n24475 | ~n21642;
  assign n20874 = ~n20873 | ~n20872;
  assign n20876 = ~n20875 & ~n20874;
  assign P2_U3195 = ~n20877 | ~n20876;
  assign n20880 = n20879 ^ n20878;
  assign n20891 = ~n20880 | ~n24506;
  assign n20889 = ~n21544 & ~n21025;
  assign n20885 = ~n24499 & ~n20881;
  assign n20883 = ~n24500 | ~n25571;
  assign n20882 = ~P2_REG3_REG_25__SCAN_IN | ~P2_U3088;
  assign n20884 = ~n20883 | ~n20882;
  assign n20887 = ~n20885 & ~n20884;
  assign n20886 = ~n24475 | ~n21545;
  assign n20888 = ~n20887 | ~n20886;
  assign n20890 = ~n20889 & ~n20888;
  assign P2_U3197 = ~n20891 | ~n20890;
  assign n20893 = ~n20892;
  assign n20895 = ~n20902 & ~n20893;
  assign n21016 = ~n20895 | ~n20894;
  assign n20897 = ~n20895;
  assign n21015 = ~n20897 | ~n20896;
  assign n20898 = ~n21015 | ~n21017;
  assign n20900 = n21016 & n20898;
  assign n20906 = ~n20900 & ~n20899;
  assign n20904 = ~n20902 & ~n20901;
  assign n20905 = ~n20904 & ~n20903;
  assign n20907 = n20906 | n20905;
  assign n20916 = ~n20907 | ~n24506;
  assign n20914 = ~n21771 & ~n21025;
  assign n20908 = ~n24455 | ~n21436;
  assign n24854 = ~P2_REG3_REG_16__SCAN_IN | ~P2_U3088;
  assign n20910 = ~n20908 | ~n24854;
  assign n20909 = ~n24484 & ~n21760;
  assign n20912 = ~n20910 & ~n20909;
  assign n20911 = ~n24475 | ~n21778;
  assign n20913 = ~n20912 | ~n20911;
  assign n20915 = ~n20914 & ~n20913;
  assign P2_U3198 = ~n20916 | ~n20915;
  assign n20919 = n20918 | n20917;
  assign n20929 = ~n20920 | ~n24506;
  assign n20927 = ~n14436 & ~n21025;
  assign n20921 = ~n24455 | ~n21734;
  assign n24879 = ~P2_REG3_REG_17__SCAN_IN | ~P2_U3088;
  assign n20923 = ~n20921 | ~n24879;
  assign n20922 = ~n24484 & ~n21791;
  assign n20925 = ~n20923 & ~n20922;
  assign n20924 = ~n24475 | ~n21745;
  assign n20926 = ~n20925 | ~n20924;
  assign n20928 = ~n20927 & ~n20926;
  assign P2_U3200 = ~n20929 | ~n20928;
  assign n20941 = ~n20931 | ~n24506;
  assign n20939 = ~n13986 & ~n21025;
  assign n20935 = ~n24499 & ~n21560;
  assign n20933 = ~n24500 | ~n25568;
  assign n20932 = ~P2_REG3_REG_24__SCAN_IN | ~P2_U3088;
  assign n20934 = ~n20933 | ~n20932;
  assign n20937 = ~n20935 & ~n20934;
  assign n20936 = ~n24475 | ~n21572;
  assign n20938 = ~n20937 | ~n20936;
  assign n20940 = ~n20939 & ~n20938;
  assign P2_U3201 = ~n20941 | ~n20940;
  assign n20945 = ~n20944 | ~n20943;
  assign n20946 = n20942 ^ ~n20945;
  assign n20958 = ~n20946 | ~n24506;
  assign n20947 = ~n21975;
  assign n20956 = ~n20947 & ~n21025;
  assign n20952 = ~n24499 & ~n20948;
  assign n20950 = ~n24500 | ~n25556;
  assign n20949 = ~P2_REG3_REG_20__SCAN_IN | ~P2_U3088;
  assign n20951 = ~n20950 | ~n20949;
  assign n20954 = ~n20952 & ~n20951;
  assign n20953 = ~n24475 | ~n21666;
  assign n20955 = ~n20954 | ~n20953;
  assign n20957 = ~n20956 & ~n20955;
  assign P2_U3205 = ~n20958 | ~n20957;
  assign n20962 = n20961 ^ n20960;
  assign n20972 = ~n20962 | ~n24506;
  assign n20970 = ~n21620 & ~n21025;
  assign n20966 = ~n24499 & ~n21561;
  assign n20964 = ~n24500 | ~n25562;
  assign n20963 = ~P2_REG3_REG_22__SCAN_IN | ~P2_U3088;
  assign n20965 = ~n20964 | ~n20963;
  assign n20968 = ~n20966 & ~n20965;
  assign n20967 = ~n24475 | ~n21621;
  assign n20969 = ~n20968 | ~n20967;
  assign n20971 = ~n20970 & ~n20969;
  assign P2_U3207 = ~n20972 | ~n20971;
  assign n20975 = ~n20974 | ~n20973;
  assign n20977 = n20976 ^ ~n20975;
  assign n20982 = ~n20977 | ~n24506;
  assign n20980 = ~n24499 & ~n21845;
  assign n20978 = ~n24500 | ~n25000;
  assign n24739 = ~P2_REG3_REG_11__SCAN_IN | ~P2_U3088;
  assign n20979 = ~n20978 | ~n24739;
  assign n20981 = ~n20980 & ~n20979;
  assign n20984 = ~n20982 | ~n20981;
  assign n20983 = ~n24511 & ~n24941;
  assign n20986 = ~n20984 & ~n20983;
  assign n20985 = ~n24508 | ~n25506;
  assign P2_U3208 = ~n20986 | ~n20985;
  assign n20989 = n20988 ^ n20987;
  assign n20999 = ~n20989 | ~n24506;
  assign n20997 = ~n21722 & ~n21025;
  assign n20990 = ~n24455 | ~n25556;
  assign n24895 = ~P2_REG3_REG_18__SCAN_IN | ~P2_U3088;
  assign n20992 = ~n20990 | ~n24895;
  assign n20991 = ~n24484 & ~n21759;
  assign n20995 = ~n20992 & ~n20991;
  assign n20993 = ~n21723;
  assign n20994 = ~n24475 | ~n20993;
  assign n20996 = ~n20995 | ~n20994;
  assign n20998 = ~n20997 & ~n20996;
  assign P2_U3210 = ~n20999 | ~n20998;
  assign n21003 = ~n21001 | ~n21002;
  assign n21004 = ~n21000 | ~n21003;
  assign n21014 = ~n21004 | ~n24506;
  assign n21012 = ~n21521 & ~n21025;
  assign n21006 = ~n24455 | ~n25580;
  assign n21005 = ~P2_REG3_REG_26__SCAN_IN | ~P2_U3088;
  assign n21008 = ~n21006 | ~n21005;
  assign n21007 = ~n24484 & ~n21560;
  assign n21010 = ~n21008 & ~n21007;
  assign n21009 = ~n24475 | ~n21522;
  assign n21011 = ~n21010 | ~n21009;
  assign n21013 = ~n21012 & ~n21011;
  assign P2_U3212 = ~n21014 | ~n21013;
  assign n21018 = ~n21016 | ~n21015;
  assign n21019 = n21018 ^ ~n21017;
  assign n21029 = ~n21019 | ~n24506;
  assign n21022 = ~n24499 & ~n21791;
  assign n21020 = ~n24500 | ~n21413;
  assign n24831 = ~P2_REG3_REG_15__SCAN_IN | ~P2_U3088;
  assign n21021 = ~n21020 | ~n24831;
  assign n21024 = ~n21022 & ~n21021;
  assign n21023 = ~n24475 | ~n21805;
  assign n21027 = ~n21024 | ~n21023;
  assign n21026 = ~n21025 & ~n21804;
  assign n21028 = ~n21027 & ~n21026;
  assign P2_U3213 = ~n21029 | ~n21028;
  assign n24334 = n21031 | n21339;
  assign n21033 = n21032 | n21456;
  assign n21034 = ~n24334 | ~n21033;
  assign n21392 = n21394 | n21417;
  assign n21159 = ~n21365 | ~n21407;
  assign n21369 = ~n21058;
  assign n21038 = ~n13124 | ~n21818;
  assign n21036 = n21035 & n21038;
  assign n21041 = ~n21037 | ~n21036;
  assign n21039 = ~n21038;
  assign n21040 = n21039 | n21377;
  assign n21220 = ~n21041 | ~n21040;
  assign n21046 = ~n21219 | ~n21220;
  assign n21212 = ~n22041 | ~n21377;
  assign n21211 = ~n13124 | ~n21413;
  assign n21044 = n21212 & n21211;
  assign n21043 = ~n22041 | ~n13124;
  assign n21042 = ~n21369 | ~n21413;
  assign n21210 = ~n21043 | ~n21042;
  assign n21045 = ~n21044 | ~n21210;
  assign n21047 = ~n13124 | ~n25254;
  assign n21055 = ~n21047 | ~n14816;
  assign n21049 = ~n21395;
  assign n21048 = n17029 | n21402;
  assign n21054 = n21049 & n21048;
  assign n21051 = n21055 | n21054;
  assign n21050 = n14877 | n14816;
  assign n21053 = n21051 & n21050;
  assign n21052 = ~n21377 | ~n25254;
  assign n21057 = ~n21053 | ~n21052;
  assign n21056 = ~n21055 | ~n21054;
  assign n21065 = ~n21057 | ~n21056;
  assign n21060 = ~n21309 | ~n25389;
  assign n21059 = ~n13124 | ~n25274;
  assign n21063 = ~n21309 | ~n25274;
  assign n21062 = n14877 | n21061;
  assign n21064 = ~n21071 | ~n21070;
  assign n21075 = ~n21065 | ~n21064;
  assign n21067 = ~n21309 | ~n25252;
  assign n21066 = ~n13124 | ~n25399;
  assign n21077 = n21067 & n21066;
  assign n21069 = ~n21309 | ~n25399;
  assign n21068 = ~n13124 | ~n25252;
  assign n21076 = ~n21069 | ~n21068;
  assign n21073 = n21077 & n21076;
  assign n21079 = ~n21076;
  assign n21078 = ~n21077;
  assign n21080 = ~n21079 | ~n21078;
  assign n21082 = ~n25410 | ~n21377;
  assign n21081 = ~n13124 | ~n25214;
  assign n21087 = n21082 & n21081;
  assign n21084 = ~n25410 | ~n13124;
  assign n21083 = ~n21309 | ~n25214;
  assign n21086 = ~n21084 | ~n21083;
  assign n21085 = ~n21087 | ~n21086;
  assign n21089 = ~n21086;
  assign n21088 = ~n21087;
  assign n21096 = ~n21089 | ~n21088;
  assign n21092 = ~n21309 | ~n25183;
  assign n21091 = n14877 | n21090;
  assign n21099 = n21092 & n21091;
  assign n21094 = ~n21369 | ~n25420;
  assign n21093 = ~n13124 | ~n25183;
  assign n21098 = ~n21094 | ~n21093;
  assign n21095 = ~n21099 | ~n21098;
  assign n21097 = n21096 & n21095;
  assign n21101 = ~n21098;
  assign n21100 = ~n21099;
  assign n21107 = ~n21101 | ~n21100;
  assign n21103 = ~n21369 | ~n25432;
  assign n21102 = ~n13124 | ~n25150;
  assign n21115 = n21103 & n21102;
  assign n21105 = ~n21369 | ~n25150;
  assign n21104 = ~n13124 | ~n25432;
  assign n21114 = ~n21105 | ~n21104;
  assign n21106 = ~n21115 | ~n21114;
  assign n21108 = n21107 & n21106;
  assign n21121 = ~n21109 | ~n21108;
  assign n21111 = ~n21369 | ~n25126;
  assign n21110 = ~n25090 | ~n13124;
  assign n21127 = n21111 & n21110;
  assign n21113 = ~n21369 | ~n25090;
  assign n21112 = ~n13124 | ~n25126;
  assign n21126 = ~n21113 | ~n21112;
  assign n21119 = ~n21127 | ~n21126;
  assign n21117 = ~n21114;
  assign n21116 = ~n21115;
  assign n21118 = ~n21117 | ~n21116;
  assign n21120 = n21119 & n21118;
  assign n21140 = ~n21121 | ~n21120;
  assign n21123 = ~n25454 | ~n21159;
  assign n21122 = ~n13124 | ~n25022;
  assign n21145 = n21123 & n21122;
  assign n21125 = ~n25454 | ~n13124;
  assign n21124 = ~n21309 | ~n25022;
  assign n21144 = ~n21125 | ~n21124;
  assign n21131 = ~n21145 | ~n21144;
  assign n21129 = ~n21126;
  assign n21128 = ~n21127;
  assign n21130 = ~n21129 | ~n21128;
  assign n21138 = n21131 & n21130;
  assign n21133 = ~n25467 | ~n21377;
  assign n21132 = ~n13124 | ~n25049;
  assign n21142 = ~n21133 | ~n21132;
  assign n21137 = ~n21142;
  assign n21135 = ~n25467 | ~n13124;
  assign n21134 = ~n21377 | ~n25049;
  assign n21143 = n21135 & n21134;
  assign n21136 = ~n21143;
  assign n21141 = ~n21137 | ~n21136;
  assign n21139 = n21138 & n21141;
  assign n21149 = ~n21143 | ~n21142;
  assign n21147 = ~n21144;
  assign n21146 = ~n21145;
  assign n21148 = ~n21147 | ~n21146;
  assign n21151 = ~n25479 | ~n13124;
  assign n21150 = ~n21369 | ~n25021;
  assign n21171 = n21151 & n21150;
  assign n21153 = ~n25479 | ~n21377;
  assign n21152 = ~n13124 | ~n25021;
  assign n21170 = ~n21153 | ~n21152;
  assign n21154 = ~n21171 | ~n21170;
  assign n21156 = ~n25506 | ~n13124;
  assign n21155 = ~n21369 | ~n24976;
  assign n21186 = n21156 & n21155;
  assign n21158 = ~n25506 | ~n21377;
  assign n21157 = ~n13124 | ~n24976;
  assign n21185 = ~n21158 | ~n21157;
  assign n21167 = ~n21186 | ~n21185;
  assign n21161 = ~n25489 | ~n13124;
  assign n21341 = ~n21058 | ~n21339;
  assign n21160 = ~n21341 | ~n25000;
  assign n21174 = ~n21161 | ~n21160;
  assign n21165 = ~n21174;
  assign n21163 = ~n25489 | ~n21377;
  assign n21162 = ~n13124 | ~n25000;
  assign n21175 = n21163 & n21162;
  assign n21164 = ~n21175;
  assign n21166 = ~n21165 | ~n21164;
  assign n21169 = n21167 & n21166;
  assign n21179 = ~n21169;
  assign n21173 = ~n21170;
  assign n21172 = ~n21171;
  assign n21177 = ~n21173 | ~n21172;
  assign n21176 = ~n21175 | ~n21174;
  assign n21178 = n21177 & n21176;
  assign n21180 = n21179 | n21178;
  assign n21182 = ~n24394 | ~n21377;
  assign n21181 = ~n13124 | ~n24955;
  assign n21197 = n21182 & n21181;
  assign n21184 = ~n24394 | ~n13124;
  assign n21183 = ~n21341 | ~n24955;
  assign n21196 = ~n21184 | ~n21183;
  assign n21190 = ~n21197 | ~n21196;
  assign n21188 = ~n21185;
  assign n21187 = ~n21186;
  assign n21189 = ~n21188 | ~n21187;
  assign n21191 = n21190 & n21189;
  assign n21193 = ~n24473 | ~n13124;
  assign n21192 = ~n21369 | ~n21817;
  assign n21205 = n21193 & n21192;
  assign n21195 = ~n24473 | ~n21377;
  assign n21194 = ~n13124 | ~n21817;
  assign n21204 = ~n21195 | ~n21194;
  assign n21201 = ~n21205 | ~n21204;
  assign n21199 = ~n21196;
  assign n21198 = ~n21197;
  assign n21200 = ~n21199 | ~n21198;
  assign n21202 = n21201 & n21200;
  assign n21209 = ~n21203 | ~n21202;
  assign n21207 = ~n21204;
  assign n21206 = ~n21205;
  assign n21208 = ~n21207 | ~n21206;
  assign n21216 = ~n21209 | ~n21208;
  assign n21214 = ~n21210;
  assign n21213 = ~n21212 | ~n21211;
  assign n21215 = ~n21214 | ~n21213;
  assign n21217 = ~n21216 | ~n21215;
  assign n21222 = ~n21219;
  assign n21221 = ~n21220;
  assign n21230 = ~n21222 | ~n21221;
  assign n21224 = ~n22018 | ~n21377;
  assign n21223 = ~n13124 | ~n21735;
  assign n21229 = ~n21224 | ~n21223;
  assign n21226 = ~n22018 | ~n13124;
  assign n21225 = ~n21369 | ~n21735;
  assign n21227 = ~n21226 | ~n21225;
  assign n21231 = ~n21229;
  assign n21232 = n21231 & n21230;
  assign n21233 = ~n21228 | ~n21232;
  assign n21242 = ~n21234 | ~n21233;
  assign n21236 = ~n22008 | ~n21377;
  assign n21235 = ~n21436 | ~n13124;
  assign n21241 = n21236 & n21235;
  assign n21238 = ~n22008 | ~n13124;
  assign n21237 = ~n21309 | ~n21436;
  assign n21239 = ~n21238 | ~n21237;
  assign n21243 = ~n21242 | ~n21241;
  assign n21245 = ~n21997 | ~n21369;
  assign n21244 = ~n21734 | ~n13124;
  assign n21249 = n21245 & n21244;
  assign n21247 = ~n21997 | ~n13124;
  assign n21246 = ~n21377 | ~n21734;
  assign n21248 = ~n21247 | ~n21246;
  assign n21251 = ~n21250 | ~n21249;
  assign n21254 = ~n21986 | ~n21377;
  assign n21253 = ~n13124 | ~n25556;
  assign n21260 = ~n21254 | ~n21253;
  assign n21258 = ~n21259 | ~n21260;
  assign n21256 = ~n21986 | ~n13124;
  assign n21255 = ~n21309 | ~n25556;
  assign n21257 = ~n21256 | ~n21255;
  assign n21264 = ~n21258 | ~n21257;
  assign n21262 = ~n21259;
  assign n21261 = ~n21260;
  assign n21263 = ~n21262 | ~n21261;
  assign n21270 = ~n21264 | ~n21263;
  assign n21266 = ~n21975 | ~n13124;
  assign n21265 = ~n21309 | ~n25559;
  assign n21268 = ~n21975 | ~n21377;
  assign n21267 = ~n13124 | ~n25559;
  assign n21269 = ~n21268 | ~n21267;
  assign n21272 = ~n21965 | ~n21377;
  assign n21271 = ~n13124 | ~n25562;
  assign n21281 = n21272 & n21271;
  assign n21274 = ~n21965 | ~n13124;
  assign n21273 = ~n21377 | ~n25562;
  assign n21280 = ~n21274 | ~n21273;
  assign n21275 = ~n21281 | ~n21280;
  assign n21277 = ~n21954 | ~n21377;
  assign n21276 = ~n13124 | ~n25565;
  assign n21285 = n21277 & n21276;
  assign n21279 = ~n21954 | ~n13124;
  assign n21278 = ~n21377 | ~n25565;
  assign n21284 = ~n21279 | ~n21278;
  assign n21283 = ~n21285 & ~n21284;
  assign n21282 = ~n21281 & ~n21280;
  assign n21286 = ~n21285 | ~n21284;
  assign n21288 = n21598 | n14877;
  assign n21287 = ~n21341 | ~n25568;
  assign n21293 = n21288 & n21287;
  assign n21290 = n21598 | n21058;
  assign n21289 = ~n13124 | ~n25568;
  assign n21292 = ~n21290 | ~n21289;
  assign n21291 = ~n21293 | ~n21292;
  assign n21295 = ~n21292;
  assign n21294 = ~n21293;
  assign n21296 = ~n21295 | ~n21294;
  assign n21299 = ~n13986 & ~n21058;
  assign n21298 = ~n21587 & ~n14877;
  assign n21303 = ~n21299 & ~n21298;
  assign n21302 = ~n13986 & ~n14877;
  assign n21300 = ~n21341;
  assign n21301 = ~n21300 & ~n21587;
  assign n21305 = ~n21921 | ~n21377;
  assign n21304 = ~n13124 | ~n25574;
  assign n21315 = n21305 & n21304;
  assign n21307 = ~n21921 | ~n13124;
  assign n21306 = ~n21369 | ~n25574;
  assign n21314 = ~n21307 | ~n21306;
  assign n21308 = ~n21315 | ~n21314;
  assign n21311 = ~n21910 | ~n13124;
  assign n21310 = ~n21309 | ~n25577;
  assign n21327 = n21311 & n21310;
  assign n21313 = ~n21910 | ~n21369;
  assign n21312 = ~n13124 | ~n25577;
  assign n21326 = ~n21313 | ~n21312;
  assign n21319 = ~n21327 | ~n21326;
  assign n21317 = ~n21314;
  assign n21316 = ~n21315;
  assign n21318 = ~n21317 | ~n21316;
  assign n21320 = ~n21319 | ~n21318;
  assign n21322 = ~n21323 | ~n21369;
  assign n21321 = ~n13124 | ~n25580;
  assign n21332 = n21322 & n21321;
  assign n21325 = ~n21323 | ~n13124;
  assign n21324 = ~n21341 | ~n25580;
  assign n21331 = ~n21325 | ~n21324;
  assign n21329 = ~n21332 | ~n21331;
  assign n21330 = ~n21329 | ~n21328;
  assign n21335 = ~n21333 | ~n13124;
  assign n21334 = ~n25583 | ~n21341;
  assign n21349 = n21335 & n21334;
  assign n21337 = n21487 | n21058;
  assign n21336 = ~n25583 | ~n13124;
  assign n21348 = ~n21337 | ~n21336;
  assign n21338 = ~n21349 & ~n21348;
  assign n21344 = ~n21345 | ~n13124;
  assign n21342 = ~n21340 | ~n21339;
  assign n21343 = ~n21342 | ~n21341;
  assign n21373 = n21344 & n21343;
  assign n21347 = ~n21345 | ~n21309;
  assign n21346 = ~n25586 | ~n13124;
  assign n21372 = ~n21347 | ~n21346;
  assign n21351 = ~n21373 | ~n21372;
  assign n21350 = ~n21349 | ~n21348;
  assign n21355 = ~n23114 | ~n21352;
  assign n22127 = ~P1_DATAO_REG_31__SCAN_IN;
  assign n21354 = n21353 | n22127;
  assign n21358 = ~n16780 | ~P2_REG1_REG_31__SCAN_IN;
  assign n21357 = ~n21356 | ~P2_REG2_REG_31__SCAN_IN;
  assign n21361 = ~n21358 | ~n21357;
  assign n21360 = n21359 & P2_REG0_REG_31__SCAN_IN;
  assign n25593 = n21361 | n21360;
  assign n21376 = n21462 | n25593;
  assign n21362 = ~n21462 | ~n25593;
  assign n21450 = ~n21376 | ~n21362;
  assign n21364 = ~n21363 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n21368 = ~n21469 | ~n13124;
  assign n21385 = ~n21309 | ~n25593;
  assign n21366 = ~n21385 | ~n21365;
  assign n21367 = ~n21366 | ~n25589;
  assign n21382 = n21368 & n21367;
  assign n21370 = ~n13124 | ~n25589;
  assign n21381 = ~n21371 | ~n21370;
  assign n21375 = ~n21382 & ~n21381;
  assign n21374 = ~n21373 & ~n21372;
  assign n21388 = ~n21376;
  assign n21379 = ~n21462 | ~n21377;
  assign n21378 = ~n13124 | ~n25593;
  assign n21380 = ~n21379 | ~n21378;
  assign n21384 = ~n21381;
  assign n21383 = ~n21382;
  assign n21386 = ~n21462 | ~n13124;
  assign n21387 = ~n21386 | ~n21385;
  assign n21389 = ~n21388 & ~n21387;
  assign n21390 = ~n17029 & ~n21456;
  assign n21391 = ~n21390 | ~n21417;
  assign n21393 = ~n21392 | ~n21391;
  assign n21399 = ~n21394;
  assign n21397 = ~n21395 | ~n25194;
  assign n21396 = ~n21417 | ~n21456;
  assign n21398 = ~n21397 | ~n21396;
  assign n24518 = ~n24516;
  assign n21400 = ~n25253 | ~n24518;
  assign n21406 = ~n21401 & ~n21400;
  assign n21404 = n21403 | n21402;
  assign n21405 = ~n21404 | ~P2_B_REG_SCAN_IN;
  assign n21519 = ~n21410 | ~n21409;
  assign n21442 = ~n21519 & ~n21556;
  assign n21639 = ~n14384 | ~n21412;
  assign n21679 = n21986 ^ ~n21709;
  assign n21827 = n22041 ^ ~n21413;
  assign n21869 = ~n21415 | ~n21414;
  assign n21429 = ~n21869 & ~n24997;
  assign n24969 = n25489 ^ ~n24434;
  assign n21428 = ~n24947 & ~n24969;
  assign n21416 = n25254 | n24454;
  assign n21419 = ~n25142 | ~n25279;
  assign n21418 = ~n25245 | ~n21417;
  assign n21420 = ~n21419 & ~n21418;
  assign n21421 = ~n25076 | ~n21420;
  assign n25122 = n25104 ^ ~n25150;
  assign n21422 = ~n21421 & ~n25122;
  assign n21423 = ~n21422 | ~n25174;
  assign n21425 = ~n21423 & ~n25136;
  assign n21424 = ~n25052;
  assign n21426 = ~n21425 | ~n21424;
  assign n21427 = ~n21426 & ~n25029;
  assign n21844 = ~n21431 | ~n21430;
  assign n21433 = ~n21432 & ~n21844;
  assign n21434 = n21789 & n21433;
  assign n21435 = n21827 & n21434;
  assign n21743 = n22008 ^ ~n21436;
  assign n21438 = ~n21707 | ~n21437;
  assign n21439 = n21679 | n21438;
  assign n21443 = ~n21442 | ~n21441;
  assign n21540 = n21921 ^ ~n21560;
  assign n21585 = n21598 ^ ~n25568;
  assign n21448 = ~n21446 | ~n14257;
  assign n21452 = ~n21450 | ~n21449;
  assign n21451 = n13990 ^ ~n25589;
  assign n21453 = ~n21455 & ~n17029;
  assign n21458 = ~n21457 & ~P2_B_REG_SCAN_IN;
  assign n21894 = n21461 ^ ~n21462;
  assign n21468 = ~n21894 | ~n25263;
  assign n21895 = ~n21462;
  assign n21466 = ~n21895 & ~n25105;
  assign n21902 = n21463 & n25593;
  assign n21472 = ~n25284 | ~n21902;
  assign n21464 = ~n25282 | ~P2_REG2_REG_31__SCAN_IN;
  assign n21465 = ~n21472 | ~n21464;
  assign n21467 = ~n21466 & ~n21465;
  assign P2_U3234 = ~n21468 | ~n21467;
  assign n21901 = n21470 ^ n21469;
  assign n21476 = ~n21901 | ~n25263;
  assign n21474 = ~n13990 & ~n25105;
  assign n21471 = ~n25282 | ~P2_REG2_REG_30__SCAN_IN;
  assign n21473 = ~n21472 | ~n21471;
  assign n21475 = ~n21474 & ~n21473;
  assign P2_U3235 = ~n21476 | ~n21475;
  assign n21481 = ~n21477 & ~n25194;
  assign n21479 = ~n21478 | ~n25233;
  assign n21480 = ~n21479 | ~n25284;
  assign n21482 = ~n21481 & ~n21480;
  assign n21485 = ~n21483 | ~n21482;
  assign n21484 = n25284 | P2_REG2_REG_28__SCAN_IN;
  assign n21491 = ~n21485 | ~n21484;
  assign n21489 = ~n21486 & ~n25099;
  assign n21488 = ~n21487 & ~n25105;
  assign n21490 = ~n21489 & ~n21488;
  assign P2_U3237 = ~n21491 | ~n21490;
  assign n21494 = ~n21492 | ~n25284;
  assign n21493 = n25284 | P2_REG2_REG_27__SCAN_IN;
  assign n21506 = ~n21494 | ~n21493;
  assign n21504 = ~n21495 & ~n25099;
  assign n21502 = ~n21496 | ~n21803;
  assign n21500 = ~n21497 & ~n25105;
  assign n21499 = ~n25267 & ~n21498;
  assign n21501 = ~n21500 & ~n21499;
  assign n21503 = ~n21502 | ~n21501;
  assign n21505 = ~n21504 & ~n21503;
  assign P2_U3238 = ~n21506 | ~n21505;
  assign n21509 = ~n21507 | ~n21508;
  assign n21510 = n21509 ^ ~n21519;
  assign n21514 = ~n21510 & ~n25270;
  assign n21512 = ~n25580 | ~n25273;
  assign n21511 = ~n25574 | ~n25253;
  assign n21513 = ~n21512 | ~n21511;
  assign n21516 = ~n21916 | ~n25284;
  assign n21515 = n25284 | P2_REG2_REG_26__SCAN_IN;
  assign n21531 = ~n21516 | ~n21515;
  assign n21520 = ~n21518 | ~n21517;
  assign n21908 = n21520 ^ ~n21519;
  assign n21529 = ~n21908 & ~n21828;
  assign n21909 = n13136 ^ ~n21521;
  assign n21527 = ~n21909 | ~n25263;
  assign n21525 = ~n21521 & ~n25105;
  assign n21523 = ~n21522;
  assign n21524 = ~n25267 & ~n21523;
  assign n21526 = ~n21525 & ~n21524;
  assign n21528 = ~n21527 | ~n21526;
  assign n21530 = ~n21529 & ~n21528;
  assign P2_U3239 = ~n21531 | ~n21530;
  assign n21533 = n21532 ^ ~n21540;
  assign n21537 = ~n21533 & ~n25270;
  assign n21535 = ~n25571 | ~n25253;
  assign n21534 = ~n25577 | ~n25273;
  assign n21536 = ~n21535 | ~n21534;
  assign n21927 = ~n21537 & ~n21536;
  assign n21539 = ~n21927 | ~n25284;
  assign n21538 = n25284 | P2_REG2_REG_25__SCAN_IN;
  assign n21554 = ~n21539 | ~n21538;
  assign n21919 = n21541 ^ ~n21540;
  assign n21552 = ~n21919 & ~n21828;
  assign n21543 = ~n21542 | ~n21921;
  assign n21920 = n13136 & n21543;
  assign n21550 = ~n21920 | ~n25263;
  assign n21548 = ~n21544 & ~n25105;
  assign n21546 = ~n21545;
  assign n21547 = ~n25267 & ~n21546;
  assign n21549 = ~n21548 & ~n21547;
  assign n21551 = ~n21550 | ~n21549;
  assign n21553 = ~n21552 & ~n21551;
  assign P2_U3240 = ~n21554 | ~n21553;
  assign n21557 = n21555 ^ ~n21556;
  assign n21567 = ~n21557 & ~n25270;
  assign n21570 = n21559 ^ ~n21558;
  assign n21565 = ~n21570 | ~n25248;
  assign n21563 = ~n21560 & ~n25092;
  assign n21562 = ~n21561 & ~n25079;
  assign n21564 = ~n21563 & ~n21562;
  assign n21566 = ~n21565 | ~n21564;
  assign n21938 = ~n21567 & ~n21566;
  assign n21569 = ~n21938 | ~n25284;
  assign n21568 = n25284 | P2_REG2_REG_24__SCAN_IN;
  assign n21581 = ~n21569 | ~n21568;
  assign n21930 = ~n21570;
  assign n21579 = ~n21930 & ~n25099;
  assign n21571 = ~n21943 & ~n21597;
  assign n21931 = n21571 ^ ~n21932;
  assign n21577 = ~n21931 | ~n25263;
  assign n21575 = ~n13986 & ~n25105;
  assign n21573 = ~n21572;
  assign n21574 = ~n25267 & ~n21573;
  assign n21576 = ~n21575 & ~n21574;
  assign n21578 = ~n21577 | ~n21576;
  assign n21580 = ~n21579 & ~n21578;
  assign P2_U3241 = ~n21581 | ~n21580;
  assign n21583 = n21582 ^ ~n21585;
  assign n21593 = ~n21583 & ~n25270;
  assign n21596 = n21584 ^ n21585;
  assign n21591 = ~n21596 | ~n25248;
  assign n21589 = ~n21586 & ~n25079;
  assign n21588 = ~n21587 & ~n25092;
  assign n21590 = ~n21589 & ~n21588;
  assign n21592 = ~n21591 | ~n21590;
  assign n21949 = ~n21593 & ~n21592;
  assign n21595 = ~n21949 | ~n25284;
  assign n21594 = n25284 | P2_REG2_REG_23__SCAN_IN;
  assign n21608 = ~n21595 | ~n21594;
  assign n21941 = ~n21596;
  assign n21606 = ~n21941 & ~n25099;
  assign n21942 = n21598 ^ ~n21597;
  assign n21604 = ~n21942 | ~n25263;
  assign n21602 = ~n21598 & ~n25105;
  assign n21600 = ~n21599;
  assign n21601 = ~n25267 & ~n21600;
  assign n21603 = ~n21602 & ~n21601;
  assign n21605 = ~n21604 | ~n21603;
  assign n21607 = ~n21606 & ~n21605;
  assign P2_U3242 = ~n21608 | ~n21607;
  assign n21610 = n21609 ^ n21617;
  assign n21614 = ~n21610 & ~n25270;
  assign n21612 = ~n25562 | ~n25253;
  assign n21611 = ~n25568 | ~n25273;
  assign n21613 = ~n21612 | ~n21611;
  assign n21960 = ~n21614 & ~n21613;
  assign n21616 = ~n21960 | ~n25284;
  assign n21615 = n25284 | P2_REG2_REG_22__SCAN_IN;
  assign n21630 = ~n21616 | ~n21615;
  assign n21952 = n21618 ^ ~n21617;
  assign n21628 = ~n21952 & ~n21828;
  assign n21953 = n21619 ^ ~n21954;
  assign n21626 = ~n21953 | ~n25263;
  assign n21624 = ~n21620 & ~n25105;
  assign n21622 = ~n21621;
  assign n21623 = ~n25267 & ~n21622;
  assign n21625 = ~n21624 & ~n21623;
  assign n21627 = ~n21626 | ~n21625;
  assign n21629 = ~n21628 & ~n21627;
  assign P2_U3243 = ~n21630 | ~n21629;
  assign n21632 = n21631 ^ ~n21639;
  assign n21636 = ~n21632 & ~n25270;
  assign n21634 = ~n25565 | ~n25273;
  assign n21633 = ~n25559 | ~n25253;
  assign n21635 = ~n21634 | ~n21633;
  assign n21971 = ~n21636 & ~n21635;
  assign n21638 = ~n21971 | ~n25284;
  assign n21637 = n25284 | P2_REG2_REG_21__SCAN_IN;
  assign n21651 = ~n21638 | ~n21637;
  assign n21963 = n21640 ^ ~n21639;
  assign n21649 = n21963 | n21828;
  assign n21641 = ~n21664;
  assign n21964 = n21641 ^ ~n21965;
  assign n21647 = ~n21964 | ~n25263;
  assign n21645 = ~n21965 | ~n25264;
  assign n21643 = ~n21642;
  assign n21644 = n25267 | n21643;
  assign n21646 = n21645 & n21644;
  assign n21648 = n21647 & n21646;
  assign n21650 = n21649 & n21648;
  assign P2_U3244 = ~n21651 | ~n21650;
  assign n21653 = n21660 ^ n21652;
  assign n21657 = ~n21653 & ~n25270;
  assign n21655 = ~n25556 | ~n25253;
  assign n21654 = ~n25562 | ~n25273;
  assign n21656 = ~n21655 | ~n21654;
  assign n21981 = ~n21657 & ~n21656;
  assign n21659 = n21981 & n25284;
  assign n21658 = ~n25284 & ~P2_REG2_REG_20__SCAN_IN;
  assign n21675 = ~n21659 & ~n21658;
  assign n21974 = n21661 ^ ~n21660;
  assign n21673 = n21974 | n21828;
  assign n21663 = ~n21975 | ~n21662;
  assign n21665 = n21663 & n25503;
  assign n21977 = ~n21665 | ~n21664;
  assign n21777 = ~n25284 | ~n17029;
  assign n21671 = ~n21977 & ~n21777;
  assign n21669 = ~n21975 | ~n25264;
  assign n21667 = ~n21666;
  assign n21668 = n25267 | n21667;
  assign n21670 = ~n21669 | ~n21668;
  assign n21672 = ~n21671 & ~n21670;
  assign n21674 = ~n21673 | ~n21672;
  assign P2_U3245 = n21675 | n21674;
  assign n21677 = n21676 ^ n21679;
  assign n21690 = ~n21677 & ~n25270;
  assign n21683 = ~n13256 | ~n21678;
  assign n21680 = ~n21679;
  assign n21682 = ~n21681 | ~n21680;
  assign n21688 = ~n21694 | ~n25248;
  assign n21686 = ~n13885 & ~n25079;
  assign n21685 = ~n21684 & ~n25092;
  assign n21687 = ~n21686 & ~n21685;
  assign n21689 = ~n21688 | ~n21687;
  assign n21992 = ~n21690 & ~n21689;
  assign n21693 = ~n21992 | ~n25284;
  assign n21691 = ~P2_REG2_REG_19__SCAN_IN;
  assign n21692 = ~n25282 | ~n21691;
  assign n21704 = ~n21693 | ~n21692;
  assign n21984 = ~n21694;
  assign n21702 = ~n21984 & ~n25099;
  assign n21985 = n21720 ^ n21986;
  assign n21700 = ~n21985 | ~n21803;
  assign n21698 = ~n14434 & ~n25105;
  assign n21696 = ~n21695;
  assign n21697 = ~n25267 & ~n21696;
  assign n21699 = ~n21698 & ~n21697;
  assign n21701 = ~n21700 | ~n21699;
  assign n21703 = ~n21702 & ~n21701;
  assign P2_U3246 = ~n21704 | ~n21703;
  assign n21706 = n21705 ^ ~n21707;
  assign n21715 = ~n21706 & ~n25270;
  assign n21719 = n21708 ^ ~n21707;
  assign n21713 = ~n21719 | ~n25248;
  assign n21711 = ~n21759 & ~n25079;
  assign n21710 = ~n21709 & ~n25092;
  assign n21712 = ~n21711 & ~n21710;
  assign n21714 = ~n21713 | ~n21712;
  assign n22003 = ~n21715 & ~n21714;
  assign n21718 = ~n22003 | ~n25284;
  assign n21716 = ~P2_REG2_REG_18__SCAN_IN;
  assign n21717 = ~n25282 | ~n21716;
  assign n21731 = ~n21718 | ~n21717;
  assign n21995 = ~n21719;
  assign n21729 = ~n21995 & ~n25099;
  assign n21721 = ~n21722 & ~n13386;
  assign n21996 = ~n13987 & ~n21721;
  assign n21727 = ~n21996 | ~n25263;
  assign n21725 = ~n21722 & ~n25105;
  assign n21724 = ~n25267 & ~n21723;
  assign n21726 = ~n21725 & ~n21724;
  assign n21728 = ~n21727 | ~n21726;
  assign n21730 = ~n21729 & ~n21728;
  assign P2_U3247 = ~n21731 | ~n21730;
  assign n21733 = n21732 ^ ~n21743;
  assign n21739 = ~n21733 & ~n25270;
  assign n21737 = ~n21734 | ~n25273;
  assign n21736 = ~n21735 | ~n25253;
  assign n21738 = ~n21737 | ~n21736;
  assign n22014 = ~n21739 & ~n21738;
  assign n21742 = ~n22014 | ~n25284;
  assign n21740 = ~P2_REG2_REG_17__SCAN_IN;
  assign n21741 = ~n25282 | ~n21740;
  assign n21754 = ~n21742 | ~n21741;
  assign n22006 = n21744 ^ n21743;
  assign n21752 = ~n22006 & ~n21828;
  assign n22007 = n21774 ^ n22008;
  assign n21750 = ~n22007 | ~n25263;
  assign n21748 = ~n14436 & ~n25105;
  assign n21746 = ~n21745;
  assign n21747 = ~n25267 & ~n21746;
  assign n21749 = ~n21748 & ~n21747;
  assign n21751 = ~n21750 | ~n21749;
  assign n21753 = ~n21752 & ~n21751;
  assign P2_U3248 = ~n21754 | ~n21753;
  assign n21756 = n21755 ^ ~n21758;
  assign n21766 = ~n21756 & ~n25270;
  assign n21770 = n21758 ^ n21757;
  assign n21764 = ~n21770 | ~n25248;
  assign n21762 = ~n21759 & ~n25092;
  assign n21761 = ~n21760 & ~n25079;
  assign n21763 = ~n21762 & ~n21761;
  assign n21765 = ~n21764 | ~n21763;
  assign n22024 = ~n21766 & ~n21765;
  assign n21769 = ~n22024 | ~n25284;
  assign n21767 = ~P2_REG2_REG_16__SCAN_IN;
  assign n21768 = ~n25282 | ~n21767;
  assign n21786 = ~n21769 | ~n21768;
  assign n22017 = ~n21770;
  assign n21784 = ~n22017 & ~n25099;
  assign n21773 = n21772 | n21771;
  assign n21776 = ~n21773 | ~n25503;
  assign n21775 = ~n21774;
  assign n22020 = n21776 | n21775;
  assign n21782 = ~n22020 & ~n21777;
  assign n21780 = ~n25264 | ~n22018;
  assign n21779 = ~n25233 | ~n21778;
  assign n21781 = ~n21780 | ~n21779;
  assign n21783 = n21782 | n21781;
  assign n21785 = ~n21784 & ~n21783;
  assign P2_U3249 = ~n21786 | ~n21785;
  assign n21788 = n21787 ^ ~n21789;
  assign n21797 = ~n21788 & ~n25270;
  assign n21801 = n21790 ^ ~n21789;
  assign n21795 = ~n21801 | ~n25248;
  assign n21793 = ~n21791 & ~n25092;
  assign n21792 = ~n24462 & ~n25079;
  assign n21794 = ~n21793 & ~n21792;
  assign n21796 = ~n21795 | ~n21794;
  assign n22035 = ~n21797 & ~n21796;
  assign n21800 = ~n22035 | ~n25284;
  assign n21798 = ~P2_REG2_REG_15__SCAN_IN;
  assign n21799 = ~n25282 | ~n21798;
  assign n21814 = ~n21800 | ~n21799;
  assign n22027 = ~n21801;
  assign n21812 = ~n22027 & ~n25099;
  assign n22028 = n21802 ^ ~n21804;
  assign n21810 = ~n22028 | ~n21803;
  assign n21808 = ~n25105 & ~n21804;
  assign n21806 = ~n21805;
  assign n21807 = ~n25267 & ~n21806;
  assign n21809 = ~n21808 & ~n21807;
  assign n21811 = ~n21810 | ~n21809;
  assign n21813 = ~n21812 & ~n21811;
  assign P2_U3250 = ~n21814 | ~n21813;
  assign n21816 = n21815 ^ n21827;
  assign n21822 = ~n21816 & ~n25270;
  assign n21820 = ~n21817 | ~n25253;
  assign n21819 = ~n21818 | ~n25273;
  assign n21821 = ~n21820 | ~n21819;
  assign n22047 = ~n21822 & ~n21821;
  assign n21825 = ~n22047 | ~n25284;
  assign n21823 = ~P2_REG2_REG_14__SCAN_IN;
  assign n21824 = ~n25282 | ~n21823;
  assign n21840 = ~n21825 | ~n21824;
  assign n22039 = n21827 ^ n21826;
  assign n21838 = ~n22039 & ~n21828;
  assign n22040 = n21830 ^ ~n21829;
  assign n21836 = ~n22040 | ~n25263;
  assign n21834 = ~n21830 & ~n25105;
  assign n21832 = ~n21831;
  assign n21833 = ~n25267 & ~n21832;
  assign n21835 = ~n21834 & ~n21833;
  assign n21837 = ~n21836 | ~n21835;
  assign n21839 = ~n21838 & ~n21837;
  assign P2_U3251 = ~n21840 | ~n21839;
  assign n21842 = n21841 ^ ~n21844;
  assign n21851 = ~n21842 & ~n25270;
  assign n21858 = n21843 ^ n21844;
  assign n21849 = ~n21858 | ~n25248;
  assign n21847 = ~n21845 & ~n25079;
  assign n21846 = ~n24462 & ~n25092;
  assign n21848 = ~n21847 & ~n21846;
  assign n21850 = ~n21849 | ~n21848;
  assign n22057 = ~n21851 & ~n21850;
  assign n21852 = ~n24474;
  assign n21853 = ~n25267 & ~n21852;
  assign n21854 = ~n25282 & ~n21853;
  assign n21857 = ~n22057 | ~n21854;
  assign n21855 = ~P2_REG2_REG_13__SCAN_IN;
  assign n21856 = ~n25282 | ~n21855;
  assign n21865 = ~n21857 | ~n21856;
  assign n22050 = ~n21858;
  assign n21863 = ~n22050 & ~n25099;
  assign n21859 = ~n24473;
  assign n22051 = n21859 ^ ~n21886;
  assign n21861 = ~n22051 | ~n25263;
  assign n21860 = n25105 | n21859;
  assign n21862 = ~n21861 | ~n21860;
  assign n21864 = ~n21863 & ~n21862;
  assign P2_U3252 = ~n21865 | ~n21864;
  assign n21867 = n21866 ^ ~n21869;
  assign n21875 = ~n21867 & ~n25270;
  assign n21879 = n21869 ^ n21868;
  assign n21873 = ~n21879 | ~n25248;
  assign n21871 = ~n24349 & ~n25079;
  assign n21870 = ~n24389 & ~n25092;
  assign n21872 = ~n21871 & ~n21870;
  assign n21874 = ~n21873 | ~n21872;
  assign n22067 = ~n21875 & ~n21874;
  assign n21878 = ~n22067 | ~n25284;
  assign n21876 = ~P2_REG2_REG_12__SCAN_IN;
  assign n21877 = ~n25282 | ~n21876;
  assign n21893 = ~n21878 | ~n21877;
  assign n22060 = ~n21879;
  assign n21891 = ~n22060 & ~n25099;
  assign n21883 = ~n25105 & ~n21880;
  assign n21881 = ~n24395;
  assign n21882 = ~n25267 & ~n21881;
  assign n21889 = ~n21883 & ~n21882;
  assign n21884 = ~n25506;
  assign n21885 = ~n24982 | ~n21884;
  assign n21887 = ~n21885 | ~n24394;
  assign n22061 = n21887 & n21886;
  assign n21888 = ~n25263 | ~n22061;
  assign n21890 = ~n21889 | ~n21888;
  assign n21892 = ~n21891 & ~n21890;
  assign P2_U3253 = ~n21893 | ~n21892;
  assign n21898 = ~n21894 | ~n25503;
  assign n21896 = ~n21895 & ~n25441;
  assign n21897 = ~n21896 & ~n21902;
  assign n22070 = ~n21898 | ~n21897;
  assign n21900 = ~n22070 | ~n25553;
  assign n21899 = ~n25551 | ~P2_REG1_REG_31__SCAN_IN;
  assign P2_U3530 = ~n21900 | ~n21899;
  assign n21905 = ~n21901 | ~n25503;
  assign n21903 = ~n13990 & ~n25441;
  assign n21904 = ~n21903 & ~n21902;
  assign n22073 = ~n21905 | ~n21904;
  assign n21907 = ~n22073 | ~n25553;
  assign n21906 = ~n25551 | ~P2_REG1_REG_30__SCAN_IN;
  assign P2_U3529 = ~n21907 | ~n21906;
  assign n21914 = ~n21908 & ~n22038;
  assign n21912 = ~n21909 | ~n25503;
  assign n21911 = ~n21910 | ~n25505;
  assign n21913 = ~n21912 | ~n21911;
  assign n21915 = ~n21914 & ~n21913;
  assign n22079 = ~n21916 | ~n21915;
  assign n21918 = ~n22079 | ~n25553;
  assign n21917 = ~n25551 | ~P2_REG1_REG_26__SCAN_IN;
  assign P2_U3525 = ~n21918 | ~n21917;
  assign n21925 = ~n21919 & ~n22038;
  assign n21923 = ~n21920 | ~n25503;
  assign n21922 = ~n21921 | ~n25505;
  assign n21924 = ~n21923 | ~n21922;
  assign n21926 = ~n21925 & ~n21924;
  assign n22082 = ~n21927 | ~n21926;
  assign n21929 = ~n22082 | ~n25553;
  assign n21928 = ~n25551 | ~P2_REG1_REG_25__SCAN_IN;
  assign P2_U3524 = ~n21929 | ~n21928;
  assign n21936 = ~n21930 & ~n25509;
  assign n21934 = ~n21931 | ~n25503;
  assign n21933 = ~n21932 | ~n25505;
  assign n21935 = ~n21934 | ~n21933;
  assign n21937 = ~n21936 & ~n21935;
  assign n22085 = ~n21938 | ~n21937;
  assign n21940 = ~n22085 | ~n25553;
  assign n21939 = ~n25551 | ~P2_REG1_REG_24__SCAN_IN;
  assign P2_U3523 = ~n21940 | ~n21939;
  assign n21947 = ~n21941 & ~n25509;
  assign n21945 = ~n21942 | ~n25503;
  assign n21944 = ~n21943 | ~n25505;
  assign n21946 = ~n21945 | ~n21944;
  assign n21948 = ~n21947 & ~n21946;
  assign n22088 = ~n21949 | ~n21948;
  assign n21951 = ~n22088 | ~n25553;
  assign n21950 = ~n25551 | ~P2_REG1_REG_23__SCAN_IN;
  assign P2_U3522 = ~n21951 | ~n21950;
  assign n21958 = ~n21952 & ~n22038;
  assign n21956 = ~n21953 | ~n25503;
  assign n21955 = ~n21954 | ~n25505;
  assign n21957 = ~n21956 | ~n21955;
  assign n21959 = ~n21958 & ~n21957;
  assign n22091 = ~n21960 | ~n21959;
  assign n21962 = ~n22091 | ~n25553;
  assign n21961 = ~n25551 | ~P2_REG1_REG_22__SCAN_IN;
  assign P2_U3521 = ~n21962 | ~n21961;
  assign n21969 = ~n21963 & ~n22038;
  assign n21967 = ~n21964 | ~n25503;
  assign n21966 = ~n21965 | ~n25505;
  assign n21968 = ~n21967 | ~n21966;
  assign n21970 = ~n21969 & ~n21968;
  assign n22094 = ~n21971 | ~n21970;
  assign n21973 = ~n22094 | ~n25553;
  assign n21972 = ~n25551 | ~P2_REG1_REG_21__SCAN_IN;
  assign P2_U3520 = ~n21973 | ~n21972;
  assign n21979 = ~n21974 & ~n22038;
  assign n21976 = ~n21975 | ~n25505;
  assign n21978 = ~n21977 | ~n21976;
  assign n21980 = ~n21979 & ~n21978;
  assign n22097 = ~n21981 | ~n21980;
  assign n21983 = ~n22097 | ~n25553;
  assign n21982 = ~n25551 | ~P2_REG1_REG_20__SCAN_IN;
  assign P2_U3519 = ~n21983 | ~n21982;
  assign n21990 = ~n21984 & ~n25509;
  assign n21988 = ~n21985 | ~n25503;
  assign n21987 = ~n21986 | ~n25505;
  assign n21989 = ~n21988 | ~n21987;
  assign n21991 = ~n21990 & ~n21989;
  assign n22100 = ~n21992 | ~n21991;
  assign n21994 = ~n22100 | ~n25553;
  assign n21993 = ~n25551 | ~P2_REG1_REG_19__SCAN_IN;
  assign P2_U3518 = ~n21994 | ~n21993;
  assign n22001 = ~n21995 & ~n25509;
  assign n21999 = ~n21996 | ~n25503;
  assign n21998 = ~n21997 | ~n25505;
  assign n22000 = ~n21999 | ~n21998;
  assign n22002 = ~n22001 & ~n22000;
  assign n22103 = ~n22003 | ~n22002;
  assign n22005 = ~n22103 | ~n25553;
  assign n22004 = ~n25551 | ~P2_REG1_REG_18__SCAN_IN;
  assign P2_U3517 = ~n22005 | ~n22004;
  assign n22012 = ~n22006 & ~n22038;
  assign n22010 = ~n22007 | ~n25503;
  assign n22009 = ~n22008 | ~n25505;
  assign n22011 = ~n22010 | ~n22009;
  assign n22013 = ~n22012 & ~n22011;
  assign n22106 = ~n22014 | ~n22013;
  assign n22016 = ~n22106 | ~n25553;
  assign n22015 = ~n25551 | ~P2_REG1_REG_17__SCAN_IN;
  assign P2_U3516 = ~n22016 | ~n22015;
  assign n22022 = ~n22017 & ~n25509;
  assign n22019 = ~n22018 | ~n25505;
  assign n22021 = ~n22020 | ~n22019;
  assign n22023 = ~n22022 & ~n22021;
  assign n22109 = ~n22024 | ~n22023;
  assign n22026 = ~n22109 | ~n25553;
  assign n22025 = ~n25551 | ~P2_REG1_REG_16__SCAN_IN;
  assign P2_U3515 = ~n22026 | ~n22025;
  assign n22033 = ~n22027 & ~n25509;
  assign n22031 = ~n22028 | ~n25503;
  assign n22030 = ~n22029 | ~n25505;
  assign n22032 = ~n22031 | ~n22030;
  assign n22034 = ~n22033 & ~n22032;
  assign n22112 = ~n22035 | ~n22034;
  assign n22037 = ~n22112 | ~n25553;
  assign n22036 = ~n25551 | ~P2_REG1_REG_15__SCAN_IN;
  assign P2_U3514 = ~n22037 | ~n22036;
  assign n22045 = ~n22039 & ~n22038;
  assign n22043 = ~n22040 | ~n25503;
  assign n22042 = ~n22041 | ~n25505;
  assign n22044 = ~n22043 | ~n22042;
  assign n22046 = ~n22045 & ~n22044;
  assign n22115 = ~n22047 | ~n22046;
  assign n22049 = ~n22115 | ~n25553;
  assign n22048 = ~n25551 | ~P2_REG1_REG_14__SCAN_IN;
  assign P2_U3513 = ~n22049 | ~n22048;
  assign n22055 = ~n22050 & ~n25509;
  assign n22053 = ~n22051 | ~n25503;
  assign n22052 = ~n24473 | ~n25505;
  assign n22054 = ~n22053 | ~n22052;
  assign n22056 = ~n22055 & ~n22054;
  assign n22118 = ~n22057 | ~n22056;
  assign n22059 = ~n22118 | ~n25553;
  assign n22058 = ~n25551 | ~P2_REG1_REG_13__SCAN_IN;
  assign P2_U3512 = ~n22059 | ~n22058;
  assign n22065 = ~n22060 & ~n25509;
  assign n22063 = ~n22061 | ~n25503;
  assign n22062 = ~n24394 | ~n25505;
  assign n22064 = ~n22063 | ~n22062;
  assign n22066 = ~n22065 & ~n22064;
  assign n22121 = ~n22067 | ~n22066;
  assign n22069 = ~n22121 | ~n25553;
  assign n22068 = ~n25551 | ~P2_REG1_REG_12__SCAN_IN;
  assign P2_U3511 = ~n22069 | ~n22068;
  assign n22072 = ~n22070 | ~n25515;
  assign n22071 = ~n25488 | ~P2_REG0_REG_31__SCAN_IN;
  assign P2_U3498 = ~n22072 | ~n22071;
  assign n22075 = ~n22073 | ~n25515;
  assign n22074 = ~n25488 | ~P2_REG0_REG_30__SCAN_IN;
  assign P2_U3497 = ~n22075 | ~n22074;
  assign n22078 = ~n22076 | ~n25515;
  assign n22077 = ~n25488 | ~P2_REG0_REG_27__SCAN_IN;
  assign P2_U3494 = ~n22078 | ~n22077;
  assign n22081 = ~n22079 | ~n25515;
  assign n22080 = ~n25488 | ~P2_REG0_REG_26__SCAN_IN;
  assign P2_U3493 = ~n22081 | ~n22080;
  assign n22084 = ~n22082 | ~n25515;
  assign n22083 = ~n25488 | ~P2_REG0_REG_25__SCAN_IN;
  assign P2_U3492 = ~n22084 | ~n22083;
  assign n22087 = ~n22085 | ~n25515;
  assign n22086 = ~n25488 | ~P2_REG0_REG_24__SCAN_IN;
  assign P2_U3491 = ~n22087 | ~n22086;
  assign n22090 = ~n22088 | ~n25515;
  assign n22089 = ~n25488 | ~P2_REG0_REG_23__SCAN_IN;
  assign P2_U3490 = ~n22090 | ~n22089;
  assign n22093 = ~n22091 | ~n25515;
  assign n22092 = ~n25488 | ~P2_REG0_REG_22__SCAN_IN;
  assign P2_U3489 = ~n22093 | ~n22092;
  assign n22096 = ~n22094 | ~n25515;
  assign n22095 = ~n25488 | ~P2_REG0_REG_21__SCAN_IN;
  assign P2_U3488 = ~n22096 | ~n22095;
  assign n22099 = ~n22097 | ~n25515;
  assign n22098 = ~n25488 | ~P2_REG0_REG_20__SCAN_IN;
  assign P2_U3487 = ~n22099 | ~n22098;
  assign n22102 = ~n22100 | ~n25515;
  assign n22101 = ~n25488 | ~P2_REG0_REG_19__SCAN_IN;
  assign P2_U3486 = ~n22102 | ~n22101;
  assign n22105 = ~n22103 | ~n25515;
  assign n22104 = ~n25488 | ~P2_REG0_REG_18__SCAN_IN;
  assign P2_U3484 = ~n22105 | ~n22104;
  assign n22108 = ~n22106 | ~n25515;
  assign n22107 = ~n25488 | ~P2_REG0_REG_17__SCAN_IN;
  assign P2_U3481 = ~n22108 | ~n22107;
  assign n22111 = ~n22109 | ~n25515;
  assign n22110 = ~n25488 | ~P2_REG0_REG_16__SCAN_IN;
  assign P2_U3478 = ~n22111 | ~n22110;
  assign n22114 = ~n22112 | ~n25515;
  assign n22113 = ~n25488 | ~P2_REG0_REG_15__SCAN_IN;
  assign P2_U3475 = ~n22114 | ~n22113;
  assign n22117 = ~n22115 | ~n25515;
  assign n22116 = ~n25488 | ~P2_REG0_REG_14__SCAN_IN;
  assign P2_U3472 = ~n22117 | ~n22116;
  assign n22120 = ~n22118 | ~n25515;
  assign n22119 = ~n25488 | ~P2_REG0_REG_13__SCAN_IN;
  assign P2_U3469 = ~n22120 | ~n22119;
  assign n22123 = ~n22121 | ~n25515;
  assign n22122 = ~n25488 | ~P2_REG0_REG_12__SCAN_IN;
  assign P2_U3466 = ~n22123 | ~n22122;
  assign n22131 = ~n23114 | ~n22164;
  assign n22125 = ~P2_U3088 & ~n17032;
  assign n22126 = ~n22125 | ~n22124;
  assign n22129 = ~n16583 & ~n22126;
  assign n22128 = ~n25337 & ~n22127;
  assign n22130 = ~n22129 & ~n22128;
  assign P2_U3296 = ~n22131 | ~n22130;
  assign n23123 = ~n22132;
  assign n22138 = ~n23123 | ~n22164;
  assign n22136 = ~n22133 & ~P2_U3088;
  assign n22134 = ~P1_DATAO_REG_30__SCAN_IN;
  assign n22135 = ~n25337 & ~n22134;
  assign n22137 = ~n22136 & ~n22135;
  assign P2_U3297 = ~n22138 | ~n22137;
  assign n22144 = ~n23130 | ~n22164;
  assign n22142 = ~n22139 & ~P2_U3088;
  assign n22141 = ~n25337 & ~n22140;
  assign n22143 = ~n22142 & ~n22141;
  assign P2_U3298 = ~n22144 | ~n22143;
  assign n22149 = ~n23137 | ~n22164;
  assign n24519 = n17049 | P2_U3088;
  assign n22147 = ~n24519;
  assign n22146 = ~n25337 & ~n22145;
  assign n22148 = ~n22147 & ~n22146;
  assign P2_U3299 = ~n22149 | ~n22148;
  assign n23143 = ~n22150;
  assign n22155 = ~n23143 | ~n22164;
  assign n22153 = ~n24516 & ~P2_U3088;
  assign n22152 = ~n25337 & ~n22151;
  assign n22154 = ~n22153 & ~n22152;
  assign P2_U3300 = ~n22155 | ~n22154;
  assign n22162 = ~n23149 | ~n22164;
  assign n22157 = ~n22156;
  assign n22160 = ~n22157 & ~P2_U3088;
  assign n22159 = ~n25337 & ~n22158;
  assign n22161 = ~n22160 & ~n22159;
  assign P2_U3301 = ~n22162 | ~n22161;
  assign n23157 = ~n22163;
  assign n22170 = ~n23157 | ~n22164;
  assign n22168 = ~n22165 & ~P2_U3088;
  assign n22167 = ~n25337 & ~n22166;
  assign n22169 = ~n22168 & ~n22167;
  assign P2_U3302 = ~n22170 | ~n22169;
  assign n22173 = ~n22172 | ~n22171;
  assign n22175 = ~n22174 | ~n22173;
  assign n22185 = ~n22175 | ~n23339;
  assign n22183 = ~n23015 & ~n23277;
  assign n22181 = ~n23343 | ~n22756;
  assign n22177 = ~n23279 & ~n22176;
  assign n23608 = P1_U3086 & P1_REG3_REG_14__SCAN_IN;
  assign n22179 = ~n22177 & ~n23608;
  assign n22178 = ~n23322 | ~n23017;
  assign n22180 = n22179 & n22178;
  assign n22182 = ~n22181 | ~n22180;
  assign n22184 = ~n22183 & ~n22182;
  assign P1_U3215 = ~n22185 | ~n22184;
  assign n22188 = n22186 ^ ~n22187;
  assign n22198 = ~n22188 | ~n23339;
  assign n22196 = ~n22874 & ~n23277;
  assign n22192 = ~n22550 & ~n23311;
  assign n22190 = ~n24301 | ~n23322;
  assign n22189 = ~P1_U3086 | ~P1_REG3_REG_23__SCAN_IN;
  assign n22191 = ~n22190 | ~n22189;
  assign n22194 = ~n22192 & ~n22191;
  assign n22193 = ~n24308 | ~n23332;
  assign n22195 = ~n22194 | ~n22193;
  assign n22197 = ~n22196 & ~n22195;
  assign P1_U3216 = ~n22198 | ~n22197;
  assign n22201 = ~n23307 & ~n23308;
  assign n22369 = ~n22201 & ~n22200;
  assign n22370 = n22203 | n22202;
  assign n22204 = ~n22367 | ~n22370;
  assign n22205 = n22369 ^ ~n22204;
  assign n22217 = ~n22205 | ~n23339;
  assign n22215 = ~n23277 & ~n24242;
  assign n22206 = ~P1_REG3_REG_10__SCAN_IN;
  assign n23534 = ~P1_STATE_REG_SCAN_IN & ~n22206;
  assign n22208 = ~n22207 & ~n23279;
  assign n22213 = ~n23534 & ~n22208;
  assign n22211 = ~n23241 & ~n23329;
  assign n23732 = ~n22209;
  assign n22210 = ~n23311 & ~n23732;
  assign n22212 = ~n22211 & ~n22210;
  assign n22214 = ~n22213 | ~n22212;
  assign n22216 = ~n22215 & ~n22214;
  assign P1_U3217 = ~n22217 | ~n22216;
  assign n22220 = ~n22219 & ~n22218;
  assign n22222 = ~n22220 & ~n23309;
  assign n22232 = ~n22222 | ~n22221;
  assign n22936 = ~n22223;
  assign n22230 = ~n22936 & ~n23277;
  assign n22228 = ~n23343 | ~n22635;
  assign n22226 = ~n22589 & ~n23279;
  assign n22224 = ~n23322 | ~n24289;
  assign n23731 = ~P1_REG3_REG_19__SCAN_IN | ~P1_U3086;
  assign n22225 = ~n22224 | ~n23731;
  assign n22227 = ~n22226 & ~n22225;
  assign n22229 = ~n22228 | ~n22227;
  assign n22231 = ~n22230 & ~n22229;
  assign P1_U3219 = ~n22232 | ~n22231;
  assign n22235 = ~n22233 & ~n22349;
  assign n22236 = n22235 ^ n22234;
  assign n22246 = ~n22236 | ~n23339;
  assign n22244 = ~n22905 & ~n23277;
  assign n22240 = ~n22551 & ~n23279;
  assign n22238 = ~n24295 | ~n23322;
  assign n22237 = ~P1_U3086 | ~P1_REG3_REG_21__SCAN_IN;
  assign n22239 = ~n22238 | ~n22237;
  assign n22242 = ~n22240 & ~n22239;
  assign n22241 = ~n23343 | ~n22590;
  assign n22243 = ~n22242 | ~n22241;
  assign n22245 = ~n22244 & ~n22243;
  assign P1_U3223 = ~n22246 | ~n22245;
  assign n22249 = ~n22248 | ~n22247;
  assign n22251 = n22250 ^ ~n22249;
  assign n22263 = ~n22251 | ~n23339;
  assign n22261 = ~n23343 | ~n22252;
  assign n22254 = ~n23279 & ~n22754;
  assign n23576 = ~P1_STATE_REG_SCAN_IN & ~n22253;
  assign n22256 = ~n22254 & ~n23576;
  assign n22255 = ~n23322 | ~n23753;
  assign n22259 = ~n22256 | ~n22255;
  assign n22258 = ~n22257 & ~n23277;
  assign n22260 = ~n22259 & ~n22258;
  assign n22262 = n22261 & n22260;
  assign P1_U3224 = ~n22263 | ~n22262;
  assign n22266 = n22264 ^ ~n22265;
  assign n22276 = ~n22266 | ~n23339;
  assign n22274 = ~n13598 & ~n23277;
  assign n22272 = n22847 | n23279;
  assign n22270 = ~n22496 & ~n23311;
  assign n22268 = ~n24308 | ~n23322;
  assign n22267 = ~P1_U3086 | ~P1_REG3_REG_25__SCAN_IN;
  assign n22269 = ~n22268 | ~n22267;
  assign n22271 = ~n22270 & ~n22269;
  assign n22273 = ~n22272 | ~n22271;
  assign n22275 = ~n22274 & ~n22273;
  assign P1_U3225 = ~n22276 | ~n22275;
  assign n22278 = n22277;
  assign n22280 = n22278 ^ ~n22279;
  assign n22289 = ~n22280 | ~n23339;
  assign n22287 = ~n13617 & ~n23277;
  assign n22285 = ~n23343 | ~n22708;
  assign n22281 = ~n23279 & ~n22706;
  assign n23647 = P1_U3086 & P1_REG3_REG_16__SCAN_IN;
  assign n22283 = ~n22281 & ~n23647;
  assign n22282 = ~n23322 | ~n23016;
  assign n22284 = n22283 & n22282;
  assign n22286 = ~n22285 | ~n22284;
  assign n22288 = ~n22287 & ~n22286;
  assign P1_U3226 = ~n22289 | ~n22288;
  assign n22292 = ~n22291 | ~n22290;
  assign n22294 = n22293 ^ ~n22292;
  assign n22305 = ~n22294 | ~n23339;
  assign n22966 = ~n22295;
  assign n22303 = ~n22966 & ~n23277;
  assign n22681 = ~n22296;
  assign n22301 = ~n23343 | ~n22681;
  assign n22634 = ~n24289;
  assign n22299 = ~n22634 & ~n23279;
  assign n22297 = ~n23322 | ~n22999;
  assign n23668 = ~P1_U3086 | ~P1_REG3_REG_17__SCAN_IN;
  assign n22298 = ~n22297 | ~n23668;
  assign n22300 = ~n22299 & ~n22298;
  assign n22302 = ~n22301 | ~n22300;
  assign n22304 = ~n22303 & ~n22302;
  assign P1_U3228 = ~n22305 | ~n22304;
  assign n22308 = n22306 ^ ~n22307;
  assign n22318 = ~n22308 | ~n23339;
  assign n22316 = ~n22535 & ~n23277;
  assign n22314 = ~n24311 | ~n23332;
  assign n22312 = ~n22516 & ~n23329;
  assign n22310 = ~n22527 | ~n23343;
  assign n22309 = ~P1_U3086 | ~P1_REG3_REG_24__SCAN_IN;
  assign n22311 = ~n22310 | ~n22309;
  assign n22313 = ~n22312 & ~n22311;
  assign n22315 = ~n22314 | ~n22313;
  assign n22317 = ~n22316 & ~n22315;
  assign P1_U3229 = ~n22318 | ~n22317;
  assign n22321 = n22320 ^ n22319;
  assign n22331 = ~n22321 | ~n23339;
  assign n22329 = ~n14515 & ~n23277;
  assign n22327 = ~n23343 | ~n22612;
  assign n22325 = ~n23329 & ~n22953;
  assign n22323 = ~n23332 | ~n24298;
  assign n22322 = ~P1_U3086 | ~P1_REG3_REG_20__SCAN_IN;
  assign n22324 = ~n22323 | ~n22322;
  assign n22326 = ~n22325 & ~n22324;
  assign n22328 = ~n22327 | ~n22326;
  assign n22330 = ~n22329 & ~n22328;
  assign P1_U3233 = ~n22331 | ~n22330;
  assign n22335 = ~n22333 & ~n22332;
  assign n22336 = n22335 ^ n22334;
  assign n22347 = ~n22336 | ~n23339;
  assign n22345 = ~n23311 & ~n22337;
  assign n22340 = ~n23329 & ~n22790;
  assign n22338 = ~n23332 | ~n23035;
  assign n23590 = ~P1_U3086 | ~P1_REG3_REG_13__SCAN_IN;
  assign n22339 = ~n22338 | ~n23590;
  assign n22343 = ~n22340 & ~n22339;
  assign n22342 = ~n22341 | ~n23331;
  assign n22344 = ~n22343 | ~n22342;
  assign n22346 = ~n22345 & ~n22344;
  assign P1_U3234 = ~n22347 | ~n22346;
  assign n22350 = ~n22348;
  assign n22352 = n22350 | n22349;
  assign n22354 = ~n22352 | ~n22351;
  assign n22353 = n22352 | n22351;
  assign n22355 = ~n22354 | ~n22353;
  assign n22366 = ~n22355 | ~n23339;
  assign n22364 = ~n22889 & ~n23277;
  assign n22362 = ~n24304 | ~n23332;
  assign n22572 = ~n22356;
  assign n22360 = ~n23311 & ~n22572;
  assign n22358 = ~n23322 | ~n24298;
  assign n22357 = ~P1_U3086 | ~P1_REG3_REG_22__SCAN_IN;
  assign n22359 = ~n22358 | ~n22357;
  assign n22361 = ~n22360 & ~n22359;
  assign n22363 = ~n22362 | ~n22361;
  assign n22365 = ~n22364 & ~n22363;
  assign P1_U3235 = ~n22366 | ~n22365;
  assign n22368 = ~n22367;
  assign n22373 = ~n22369 & ~n22368;
  assign n22372 = ~n22371 | ~n22370;
  assign n22374 = ~n22373 & ~n22372;
  assign n22375 = n22374 | n13392;
  assign n22385 = ~n22375 | ~n23339;
  assign n22800 = ~n22376;
  assign n22383 = ~n23311 & ~n22800;
  assign n22379 = ~n23329 & ~n14344;
  assign n22377 = ~n23332 | ~n23034;
  assign n23557 = ~P1_REG3_REG_11__SCAN_IN | ~P1_U3086;
  assign n22378 = ~n22377 | ~n23557;
  assign n22381 = ~n22379 & ~n22378;
  assign n22380 = ~n23331 | ~n23051;
  assign n22382 = ~n22381 | ~n22380;
  assign n22384 = ~n22383 & ~n22382;
  assign P1_U3236 = ~n22385 | ~n22384;
  assign n22388 = n22386 ^ ~n22387;
  assign n22398 = ~n22388 | ~n23339;
  assign n22396 = ~n22664 | ~n23331;
  assign n22394 = ~n23311 & ~n22389;
  assign n22390 = ~n23329 & ~n22706;
  assign n23687 = P1_U3086 & P1_REG3_REG_18__SCAN_IN;
  assign n22392 = ~n22390 & ~n23687;
  assign n22391 = ~n23332 | ~n24292;
  assign n22393 = ~n22392 | ~n22391;
  assign n22395 = ~n22394 & ~n22393;
  assign n22397 = n22396 & n22395;
  assign P1_U3238 = ~n22398 | ~n22397;
  assign n22402 = ~n22400 | ~n22399;
  assign n22403 = n22402 ^ ~n22401;
  assign n22412 = ~n22403 | ~n23339;
  assign n22410 = ~n22998 & ~n23277;
  assign n22408 = ~n23343 | ~n22732;
  assign n22406 = ~n23329 & ~n22731;
  assign n22404 = ~n23332 | ~n22999;
  assign n23635 = ~P1_U3086 | ~P1_REG3_REG_15__SCAN_IN;
  assign n22405 = ~n22404 | ~n23635;
  assign n22407 = ~n22406 & ~n22405;
  assign n22409 = ~n22408 | ~n22407;
  assign n22411 = ~n22410 & ~n22409;
  assign P1_U3241 = ~n22412 | ~n22411;
  assign n22420 = ~n22413 | ~n24026;
  assign n22418 = ~n22414 & ~n23980;
  assign n22415 = ~n22811;
  assign n22424 = n24021 | n22415;
  assign n22416 = ~n24021 | ~P1_REG2_REG_31__SCAN_IN;
  assign n22417 = ~n22424 | ~n22416;
  assign n22419 = ~n22418 & ~n22417;
  assign P1_U3263 = ~n22420 | ~n22419;
  assign n22809 = n22422 ^ ~n22421;
  assign n22428 = ~n22809 | ~n24026;
  assign n22426 = ~n22810 & ~n23980;
  assign n22423 = ~n24021 | ~P1_REG2_REG_30__SCAN_IN;
  assign n22425 = ~n22424 | ~n22423;
  assign n22427 = ~n22426 & ~n22425;
  assign P1_U3264 = ~n22428 | ~n22427;
  assign n22444 = ~n22429 | ~n24026;
  assign n22442 = ~n14526 & ~n23980;
  assign n22431 = ~n22436;
  assign n22430 = ~n23936 | ~P1_REG2_REG_29__SCAN_IN;
  assign n22434 = ~n22431 & ~n22430;
  assign n22433 = ~n23936 & ~n22432;
  assign n22438 = n22434 | n22433;
  assign n22437 = ~n22436 & ~n22435;
  assign n22440 = ~n22438 & ~n22437;
  assign n22439 = ~n22713 | ~n24320;
  assign n22441 = ~n22440 | ~n22439;
  assign n22443 = ~n22442 & ~n22441;
  assign n22445 = ~n22444 | ~n22443;
  assign n22449 = ~n22446 & ~n22445;
  assign n22448 = ~n22447 | ~n22772;
  assign P1_U3356 = ~n22449 | ~n22448;
  assign n22451 = ~n22817;
  assign n22456 = ~n22451 | ~n24012;
  assign n22454 = ~n22847 & ~n22789;
  assign n22453 = ~n22452 & ~n24014;
  assign n22455 = ~n22454 & ~n22453;
  assign n22460 = ~n22456 | ~n22455;
  assign n22459 = ~n22458 & ~n23991;
  assign n22462 = ~n22824 | ~n24019;
  assign n22461 = n24019 | P1_REG2_REG_27__SCAN_IN;
  assign n22471 = ~n22462 | ~n22461;
  assign n22469 = ~n22817 & ~n23892;
  assign n22818 = n22830 ^ ~n14525;
  assign n22467 = ~n22818 | ~n24026;
  assign n22465 = ~n14525 & ~n23980;
  assign n22464 = ~n23936 & ~n22463;
  assign n22466 = ~n22465 & ~n22464;
  assign n22468 = ~n22467 | ~n22466;
  assign n22470 = ~n22469 & ~n22468;
  assign P1_U3266 = ~n22471 | ~n22470;
  assign n22828 = n22472 ^ ~n22488;
  assign n22487 = ~n22828 & ~n22752;
  assign n22829 = ~n22494 & ~n22832;
  assign n22473 = ~n22829 & ~n23944;
  assign n22485 = ~n22473 | ~n22830;
  assign n22483 = ~n22832 & ~n23980;
  assign n22481 = ~n24311 | ~n22713;
  assign n22475 = ~n22474;
  assign n22479 = ~n22475 & ~n23936;
  assign n22477 = ~n22761 | ~n24316;
  assign n22476 = ~n24021 | ~P1_REG2_REG_26__SCAN_IN;
  assign n22478 = ~n22477 | ~n22476;
  assign n22480 = ~n22479 & ~n22478;
  assign n22482 = ~n22481 | ~n22480;
  assign n22484 = ~n22483 & ~n22482;
  assign n22486 = ~n22485 | ~n22484;
  assign n22490 = ~n22487 & ~n22486;
  assign n22489 = ~n22841 | ~n22772;
  assign P1_U3267 = ~n22490 | ~n22489;
  assign n22508 = ~n22845 & ~n22752;
  assign n22493 = n22492 & n22495;
  assign n22846 = ~n22494 & ~n22493;
  assign n22506 = ~n22846 | ~n24026;
  assign n24025 = ~n23980;
  assign n22504 = ~n22495 | ~n24025;
  assign n22502 = n22847 | n22707;
  assign n22500 = ~n22496 & ~n23936;
  assign n22498 = ~n24308 | ~n22713;
  assign n22497 = ~n24021 | ~P1_REG2_REG_25__SCAN_IN;
  assign n22499 = ~n22498 | ~n22497;
  assign n22501 = ~n22500 & ~n22499;
  assign n22503 = n22502 & n22501;
  assign n22505 = n22504 & n22503;
  assign n22507 = ~n22506 | ~n22505;
  assign n22512 = ~n22508 & ~n22507;
  assign n22856 = n22510 ^ ~n22509;
  assign n22511 = ~n22856 | ~n22772;
  assign P1_U3268 = ~n22512 | ~n22511;
  assign n22534 = n22513 ^ ~n22514;
  assign n22520 = ~n22534 | ~n24012;
  assign n22518 = ~n22515 & ~n24014;
  assign n22517 = ~n22516 & ~n22789;
  assign n22519 = ~n22518 & ~n22517;
  assign n22525 = ~n22520 | ~n22519;
  assign n22523 = n22522 ^ ~n22521;
  assign n22524 = ~n22523 & ~n23991;
  assign n22868 = ~n22525 & ~n22524;
  assign n22526 = n22548 ^ ~n22535;
  assign n22864 = ~n22526 | ~n24216;
  assign n22530 = ~n22864 & ~n23723;
  assign n22528 = ~n22527 | ~n24022;
  assign n22529 = ~n22528 | ~n24019;
  assign n22531 = ~n22530 & ~n22529;
  assign n22533 = ~n22868 | ~n22531;
  assign n22532 = n24019 | P1_REG2_REG_24__SCAN_IN;
  assign n22539 = ~n22533 | ~n22532;
  assign n22861 = ~n22534;
  assign n22537 = ~n22861 & ~n23892;
  assign n22536 = ~n22535 & ~n23980;
  assign n22538 = ~n22537 & ~n22536;
  assign P1_U3269 = ~n22539 | ~n22538;
  assign n22540 = ~n22871 | ~n23914;
  assign n22542 = ~n22540 | ~n24019;
  assign n22541 = n24019 | P1_REG2_REG_23__SCAN_IN;
  assign n22563 = ~n22542 | ~n22541;
  assign n22547 = ~n22543;
  assign n22546 = ~n22545 & ~n22544;
  assign n22872 = ~n22547 & ~n22546;
  assign n22561 = ~n22872 & ~n22568;
  assign n22549 = ~n22570 & ~n22874;
  assign n22873 = ~n13596 & ~n22549;
  assign n22559 = ~n22873 | ~n24026;
  assign n22557 = ~n22874 & ~n23980;
  assign n22553 = ~n22550 & ~n23936;
  assign n22552 = ~n22551 & ~n22755;
  assign n22555 = ~n22553 & ~n22552;
  assign n22554 = ~n24308 | ~n22761;
  assign n22556 = ~n22555 | ~n22554;
  assign n22558 = ~n22557 & ~n22556;
  assign n22560 = ~n22559 | ~n22558;
  assign n22562 = ~n22561 & ~n22560;
  assign P1_U3270 = ~n22563 | ~n22562;
  assign n22567 = ~n22564;
  assign n22566 = ~n22565 & ~n22585;
  assign n22887 = ~n22567 & ~n22566;
  assign n22584 = ~n22887 & ~n22568;
  assign n22571 = ~n22569 & ~n22889;
  assign n22888 = ~n22571 & ~n22570;
  assign n22582 = ~n22888 | ~n24026;
  assign n22580 = ~n22889 & ~n23980;
  assign n22578 = ~n24304 | ~n22761;
  assign n22576 = ~n22572 & ~n23936;
  assign n22574 = ~n22713 | ~n24298;
  assign n22573 = ~n24021 | ~P1_REG2_REG_22__SCAN_IN;
  assign n22575 = ~n22574 | ~n22573;
  assign n22577 = ~n22576 & ~n22575;
  assign n22579 = ~n22578 | ~n22577;
  assign n22581 = ~n22580 & ~n22579;
  assign n22583 = ~n22582 | ~n22581;
  assign n22587 = ~n22584 & ~n22583;
  assign n22898 = n13217 ^ ~n22585;
  assign n22586 = ~n22898 | ~n13493;
  assign P1_U3271 = ~n22587 | ~n22586;
  assign n22903 = n22588 ^ n22604;
  assign n22602 = ~n22903 & ~n22752;
  assign n22600 = ~n22904 | ~n24026;
  assign n22598 = ~n22905 & ~n23980;
  assign n22596 = ~n24301 | ~n22761;
  assign n22594 = ~n22589 & ~n22755;
  assign n22592 = ~n24021 | ~P1_REG2_REG_21__SCAN_IN;
  assign n22591 = ~n24022 | ~n22590;
  assign n22593 = ~n22592 | ~n22591;
  assign n22595 = ~n22594 & ~n22593;
  assign n22597 = ~n22596 | ~n22595;
  assign n22599 = ~n22598 & ~n22597;
  assign n22601 = ~n22600 | ~n22599;
  assign n22606 = ~n22602 & ~n22601;
  assign n22914 = n22603 ^ n22604;
  assign n22605 = ~n22914 | ~n22772;
  assign P1_U3272 = ~n22606 | ~n22605;
  assign n22919 = n22607 ^ ~n22625;
  assign n22623 = ~n22919 & ~n22752;
  assign n22616 = ~n14515 & ~n23980;
  assign n22609 = ~n22761 | ~n24298;
  assign n22608 = ~n24021 | ~P1_REG2_REG_20__SCAN_IN;
  assign n22611 = ~n22609 | ~n22608;
  assign n22610 = ~n22953 & ~n22755;
  assign n22614 = ~n22611 & ~n22610;
  assign n22613 = ~n22612 | ~n24022;
  assign n22615 = ~n22614 | ~n22613;
  assign n22621 = ~n22616 & ~n22615;
  assign n22619 = ~n22618 | ~n22617;
  assign n22924 = n13321 & n22619;
  assign n22620 = ~n22924 | ~n24026;
  assign n22622 = ~n22621 | ~n22620;
  assign n22628 = ~n22623 & ~n22622;
  assign n22626 = n22649 & n22624;
  assign n22929 = n22626 ^ ~n22625;
  assign n22627 = ~n22929 | ~n22772;
  assign P1_U3273 = ~n22628 | ~n22627;
  assign n22631 = n22630 & n22629;
  assign n22934 = ~n22632 & ~n22631;
  assign n22647 = ~n22934 & ~n22752;
  assign n22935 = n22633 ^ ~n22936;
  assign n22645 = ~n22935 | ~n24026;
  assign n22643 = ~n22936 & ~n23980;
  assign n22639 = ~n22634 & ~n22755;
  assign n22637 = ~n24021 | ~P1_REG2_REG_19__SCAN_IN;
  assign n22636 = ~n22635 | ~n24022;
  assign n22638 = ~n22637 | ~n22636;
  assign n22641 = ~n22639 & ~n22638;
  assign n22640 = ~n24295 | ~n22761;
  assign n22642 = ~n22641 | ~n22640;
  assign n22644 = ~n22643 & ~n22642;
  assign n22646 = ~n22645 | ~n22644;
  assign n22651 = ~n22647 & ~n22646;
  assign n22945 = ~n22649 | ~n22648;
  assign n22650 = ~n22945 | ~n22772;
  assign P1_U3274 = ~n22651 | ~n22650;
  assign n22663 = n22652 ^ n22655;
  assign n22654 = ~n22663 | ~n24012;
  assign n22653 = ~n22982 | ~n23988;
  assign n22659 = ~n22654 | ~n22653;
  assign n22657 = n22656 ^ ~n22655;
  assign n22658 = ~n22657 & ~n23991;
  assign n22961 = ~n22659 & ~n22658;
  assign n22662 = ~n22961 | ~n24019;
  assign n22661 = ~n24021 | ~n22660;
  assign n22675 = ~n22662 | ~n22661;
  assign n22950 = ~n22663;
  assign n22673 = ~n22950 & ~n23892;
  assign n22951 = n22678 ^ ~n22664;
  assign n22671 = ~n22951 | ~n24026;
  assign n22669 = ~n22952 & ~n23980;
  assign n22667 = ~n22761 | ~n24292;
  assign n22666 = ~n22665 | ~n24022;
  assign n22668 = ~n22667 | ~n22666;
  assign n22670 = ~n22669 & ~n22668;
  assign n22672 = ~n22671 | ~n22670;
  assign n22674 = ~n22673 & ~n22672;
  assign P1_U3275 = ~n22675 | ~n22674;
  assign n22964 = n22676 ^ ~n22694;
  assign n22693 = ~n22964 & ~n22752;
  assign n22677 = ~n22705;
  assign n22679 = ~n22677 & ~n22966;
  assign n22965 = ~n22679 & ~n22678;
  assign n22691 = ~n22965 | ~n24026;
  assign n22689 = ~n22966 & ~n23980;
  assign n22685 = ~n22755 & ~n22680;
  assign n22683 = ~n24021 | ~P1_REG2_REG_17__SCAN_IN;
  assign n22682 = ~n24022 | ~n22681;
  assign n22684 = ~n22683 | ~n22682;
  assign n22687 = ~n22685 & ~n22684;
  assign n22686 = ~n24289 | ~n22761;
  assign n22688 = ~n22687 | ~n22686;
  assign n22690 = ~n22689 & ~n22688;
  assign n22692 = ~n22691 | ~n22690;
  assign n22697 = ~n22693 & ~n22692;
  assign n22975 = n22695 ^ ~n22694;
  assign n22696 = ~n22975 | ~n22772;
  assign P1_U3276 = ~n22697 | ~n22696;
  assign n22701 = ~n22698;
  assign n22700 = ~n22699 & ~n22723;
  assign n22980 = ~n22701 & ~n22700;
  assign n22721 = ~n22980 & ~n22752;
  assign n22704 = ~n22703 | ~n22702;
  assign n22981 = n22705 & n22704;
  assign n22719 = ~n22981 | ~n24026;
  assign n22717 = ~n13617 & ~n23980;
  assign n22712 = ~n22707 & ~n22706;
  assign n22710 = ~n24021 | ~P1_REG2_REG_16__SCAN_IN;
  assign n22709 = ~n24022 | ~n22708;
  assign n22711 = ~n22710 | ~n22709;
  assign n22715 = ~n22712 & ~n22711;
  assign n22714 = ~n22713 | ~n23016;
  assign n22716 = ~n22715 | ~n22714;
  assign n22718 = ~n22717 & ~n22716;
  assign n22720 = ~n22719 | ~n22718;
  assign n22727 = ~n22721 & ~n22720;
  assign n22724 = ~n22722 | ~n22723;
  assign n22991 = ~n14271 | ~n22724;
  assign n22726 = ~n22991 | ~n22772;
  assign P1_U3277 = ~n22727 | ~n22726;
  assign n22996 = n22729 ^ ~n22728;
  assign n22744 = ~n22996 & ~n22752;
  assign n22997 = n22730 ^ ~n22998;
  assign n22742 = ~n22997 | ~n24026;
  assign n22740 = ~n22998 & ~n23980;
  assign n22736 = ~n22755 & ~n22731;
  assign n22734 = ~n24021 | ~P1_REG2_REG_15__SCAN_IN;
  assign n22733 = ~n24022 | ~n22732;
  assign n22735 = ~n22734 | ~n22733;
  assign n22738 = ~n22736 & ~n22735;
  assign n22737 = ~n22761 | ~n22999;
  assign n22739 = ~n22738 | ~n22737;
  assign n22741 = ~n22740 & ~n22739;
  assign n22743 = ~n22742 | ~n22741;
  assign n22748 = ~n22744 & ~n22743;
  assign n23008 = n22745 ^ ~n22746;
  assign n22747 = ~n23008 | ~n22772;
  assign P1_U3278 = ~n22748 | ~n22747;
  assign n22751 = ~n22749 | ~n22750;
  assign n23013 = n22751 ^ ~n22771;
  assign n22769 = ~n23013 & ~n22752;
  assign n23014 = n22753 ^ ~n18041;
  assign n22767 = ~n23014 | ~n24026;
  assign n22765 = ~n23015 & ~n23980;
  assign n22760 = ~n22755 & ~n22754;
  assign n22758 = ~n24021 | ~P1_REG2_REG_14__SCAN_IN;
  assign n22757 = ~n24022 | ~n22756;
  assign n22759 = ~n22758 | ~n22757;
  assign n22763 = ~n22760 & ~n22759;
  assign n22762 = ~n22761 | ~n23016;
  assign n22764 = ~n22763 | ~n22762;
  assign n22766 = ~n22765 & ~n22764;
  assign n22768 = ~n22767 | ~n22766;
  assign n22774 = ~n22769 & ~n22768;
  assign n23026 = n22770 ^ n22771;
  assign n22773 = ~n23026 | ~n22772;
  assign P1_U3279 = ~n22774 | ~n22773;
  assign n23780 = ~n22775 | ~n22776;
  assign n22779 = ~n23780;
  assign n22778 = ~n22777;
  assign n23746 = n22779 | n22778;
  assign n23745 = ~n23740;
  assign n23748 = ~n23746 | ~n23745;
  assign n22781 = ~n23748 | ~n22780;
  assign n23049 = n22786 ^ n22781;
  assign n22796 = ~n23049 & ~n18061;
  assign n22785 = n22784 & n22783;
  assign n22787 = ~n22782 | ~n22785;
  assign n22788 = n22787 ^ ~n22786;
  assign n22794 = ~n22788 | ~n24011;
  assign n22792 = ~n14344 & ~n22789;
  assign n22791 = ~n22790 & ~n24014;
  assign n22793 = ~n22792 & ~n22791;
  assign n22795 = ~n22794 | ~n22793;
  assign n23057 = ~n22796 & ~n22795;
  assign n22799 = ~n23057 | ~n24019;
  assign n22797 = ~P1_REG2_REG_11__SCAN_IN;
  assign n22798 = ~n24021 | ~n22797;
  assign n22808 = ~n22799 | ~n22798;
  assign n22806 = ~n23049 & ~n23892;
  assign n23050 = n23051 ^ n23751;
  assign n22804 = ~n23050 | ~n24026;
  assign n22802 = ~n14521 & ~n23980;
  assign n22801 = ~n23936 & ~n22800;
  assign n22803 = ~n22802 & ~n22801;
  assign n22805 = ~n22804 | ~n22803;
  assign n22807 = ~n22806 & ~n22805;
  assign P1_U3282 = ~n22808 | ~n22807;
  assign n22814 = ~n22809 | ~n24216;
  assign n22812 = ~n22810 & ~n24241;
  assign n22813 = ~n22812 & ~n22811;
  assign n23063 = ~n22814 | ~n22813;
  assign n22816 = ~n23063 | ~n24286;
  assign n22815 = ~n24284 | ~P1_REG1_REG_30__SCAN_IN;
  assign P1_U3558 = ~n22816 | ~n22815;
  assign n22823 = ~n22817 & ~n24220;
  assign n22821 = ~n22818 | ~n24216;
  assign n22820 = ~n22819 | ~n24230;
  assign n22822 = ~n22821 | ~n22820;
  assign n22825 = ~n22823 & ~n22822;
  assign n23066 = ~n22825 | ~n22824;
  assign n22827 = ~n23066 | ~n24286;
  assign n22826 = ~n24284 | ~P1_REG1_REG_27__SCAN_IN;
  assign P1_U3555 = ~n22827 | ~n22826;
  assign n22840 = ~n22828 & ~n19083;
  assign n24201 = ~n24216;
  assign n22831 = ~n22829 & ~n24201;
  assign n22838 = ~n22831 | ~n22830;
  assign n22836 = ~n22832 & ~n24241;
  assign n22834 = ~n24311 | ~n23988;
  assign n23953 = ~n24014;
  assign n22833 = ~n23953 | ~n24316;
  assign n22835 = ~n22834 | ~n22833;
  assign n22837 = ~n22836 & ~n22835;
  assign n22839 = ~n22838 | ~n22837;
  assign n22842 = ~n22840 & ~n22839;
  assign n22844 = ~n23069 | ~n24286;
  assign n22843 = ~n24284 | ~P1_REG1_REG_26__SCAN_IN;
  assign P1_U3554 = ~n22844 | ~n22843;
  assign n22855 = ~n22845 & ~n19083;
  assign n22853 = ~n22846 | ~n24216;
  assign n22851 = ~n13598 & ~n24241;
  assign n22849 = n22847 | n24014;
  assign n22848 = ~n24308 | ~n23988;
  assign n22850 = ~n22849 | ~n22848;
  assign n22852 = ~n22851 & ~n22850;
  assign n22854 = ~n22853 | ~n22852;
  assign n22858 = ~n22855 & ~n22854;
  assign n22857 = ~n22856 | ~n24011;
  assign n23072 = ~n22858 | ~n22857;
  assign n22860 = ~n23072 | ~n24286;
  assign n22859 = ~n24284 | ~P1_REG1_REG_25__SCAN_IN;
  assign P1_U3553 = ~n22860 | ~n22859;
  assign n22866 = ~n22861 & ~n24220;
  assign n22863 = ~n22862 | ~n24230;
  assign n22865 = ~n22864 | ~n22863;
  assign n22867 = ~n22866 & ~n22865;
  assign n23075 = ~n22868 | ~n22867;
  assign n22870 = ~n23075 | ~n24286;
  assign n22869 = ~n24284 | ~P1_REG1_REG_24__SCAN_IN;
  assign P1_U3552 = ~n22870 | ~n22869;
  assign n24247 = ~n19083;
  assign n22884 = ~n22871 | ~n24247;
  assign n22882 = ~n22872 & ~n23991;
  assign n22880 = ~n22873 | ~n24216;
  assign n22878 = ~n22874 & ~n24241;
  assign n22876 = ~n24308 | ~n23953;
  assign n22875 = ~n24301 | ~n23988;
  assign n22877 = ~n22876 | ~n22875;
  assign n22879 = ~n22878 & ~n22877;
  assign n22881 = ~n22880 | ~n22879;
  assign n22883 = ~n22882 & ~n22881;
  assign n23078 = ~n22884 | ~n22883;
  assign n22886 = ~n23078 | ~n24286;
  assign n22885 = ~n24284 | ~P1_REG1_REG_23__SCAN_IN;
  assign P1_U3551 = ~n22886 | ~n22885;
  assign n22897 = ~n22887 & ~n23991;
  assign n22895 = ~n22888 | ~n24216;
  assign n22893 = ~n22889 & ~n24241;
  assign n22891 = ~n24304 | ~n23953;
  assign n22890 = ~n23988 | ~n24298;
  assign n22892 = ~n22891 | ~n22890;
  assign n22894 = ~n22893 & ~n22892;
  assign n22896 = ~n22895 | ~n22894;
  assign n22900 = ~n22897 & ~n22896;
  assign n22899 = ~n22898 | ~n24247;
  assign n23081 = ~n22900 | ~n22899;
  assign n22902 = ~n23081 | ~n24286;
  assign n22901 = ~n24284 | ~P1_REG1_REG_22__SCAN_IN;
  assign P1_U3550 = ~n22902 | ~n22901;
  assign n22913 = ~n22903 & ~n19083;
  assign n22911 = ~n22904 | ~n24216;
  assign n22909 = ~n22905 & ~n24241;
  assign n22907 = ~n24301 | ~n23953;
  assign n22906 = ~n24295 | ~n23988;
  assign n22908 = ~n22907 | ~n22906;
  assign n22910 = ~n22909 & ~n22908;
  assign n22912 = ~n22911 | ~n22910;
  assign n22916 = ~n22913 & ~n22912;
  assign n22915 = ~n22914 | ~n24011;
  assign n23084 = ~n22916 | ~n22915;
  assign n22918 = ~n23084 | ~n24286;
  assign n22917 = ~n24284 | ~P1_REG1_REG_21__SCAN_IN;
  assign P1_U3549 = ~n22918 | ~n22917;
  assign n22928 = ~n22919 & ~n19083;
  assign n22923 = ~n14515 & ~n24241;
  assign n22921 = ~n24292 | ~n23988;
  assign n22920 = ~n23953 | ~n24298;
  assign n22922 = ~n22921 | ~n22920;
  assign n22926 = ~n22923 & ~n22922;
  assign n22925 = ~n22924 | ~n24216;
  assign n22927 = ~n22926 | ~n22925;
  assign n22931 = ~n22928 & ~n22927;
  assign n22930 = ~n22929 | ~n24011;
  assign n23087 = ~n22931 | ~n22930;
  assign n22933 = ~n23087 | ~n24286;
  assign n22932 = ~n24284 | ~P1_REG1_REG_20__SCAN_IN;
  assign P1_U3548 = ~n22933 | ~n22932;
  assign n22944 = ~n22934 & ~n19083;
  assign n22942 = ~n22935 | ~n24216;
  assign n22940 = ~n22936 & ~n24241;
  assign n22938 = ~n24295 | ~n23953;
  assign n22937 = ~n24289 | ~n23988;
  assign n22939 = ~n22938 | ~n22937;
  assign n22941 = ~n22940 & ~n22939;
  assign n22943 = ~n22942 | ~n22941;
  assign n22947 = ~n22944 & ~n22943;
  assign n22946 = ~n22945 | ~n24011;
  assign n23090 = ~n22947 | ~n22946;
  assign n22949 = ~n23090 | ~n24286;
  assign n22948 = ~n24284 | ~P1_REG1_REG_19__SCAN_IN;
  assign P1_U3547 = ~n22949 | ~n22948;
  assign n22959 = ~n22950 & ~n24220;
  assign n22957 = ~n22951 | ~n24216;
  assign n22955 = ~n22952 & ~n24241;
  assign n22954 = ~n22953 & ~n24014;
  assign n22956 = ~n22955 & ~n22954;
  assign n22958 = ~n22957 | ~n22956;
  assign n22960 = ~n22959 & ~n22958;
  assign n23093 = ~n22961 | ~n22960;
  assign n22963 = ~n23093 | ~n24286;
  assign n22962 = ~n24284 | ~P1_REG1_REG_18__SCAN_IN;
  assign P1_U3546 = ~n22963 | ~n22962;
  assign n22974 = ~n22964 & ~n19083;
  assign n22972 = ~n22965 | ~n24216;
  assign n22970 = ~n22966 & ~n24241;
  assign n22968 = ~n24289 | ~n23953;
  assign n22967 = ~n22999 | ~n23988;
  assign n22969 = ~n22968 | ~n22967;
  assign n22971 = ~n22970 & ~n22969;
  assign n22973 = ~n22972 | ~n22971;
  assign n22977 = ~n22974 & ~n22973;
  assign n22976 = ~n22975 | ~n24011;
  assign n23096 = ~n22977 | ~n22976;
  assign n22979 = ~n23096 | ~n24286;
  assign n22978 = ~n24284 | ~P1_REG1_REG_17__SCAN_IN;
  assign P1_U3545 = ~n22979 | ~n22978;
  assign n22990 = ~n22980 & ~n19083;
  assign n22988 = ~n22981 | ~n24216;
  assign n22986 = ~n13617 & ~n24241;
  assign n22984 = ~n22982 | ~n23953;
  assign n22983 = ~n23016 | ~n23988;
  assign n22985 = ~n22984 | ~n22983;
  assign n22987 = ~n22986 & ~n22985;
  assign n22989 = ~n22988 | ~n22987;
  assign n22993 = ~n22990 & ~n22989;
  assign n22992 = ~n22991 | ~n24011;
  assign n23099 = ~n22993 | ~n22992;
  assign n22995 = ~n23099 | ~n24286;
  assign n22994 = ~n24284 | ~P1_REG1_REG_16__SCAN_IN;
  assign P1_U3544 = ~n22995 | ~n22994;
  assign n23007 = ~n22996 & ~n19083;
  assign n23005 = ~n22997 | ~n24216;
  assign n23003 = ~n22998 & ~n24241;
  assign n23001 = ~n22999 | ~n23953;
  assign n23000 = ~n23035 | ~n23988;
  assign n23002 = ~n23001 | ~n23000;
  assign n23004 = ~n23003 & ~n23002;
  assign n23006 = ~n23005 | ~n23004;
  assign n23010 = ~n23007 & ~n23006;
  assign n23009 = ~n23008 | ~n24011;
  assign n23102 = ~n23010 | ~n23009;
  assign n23012 = ~n23102 | ~n24286;
  assign n23011 = ~n24284 | ~P1_REG1_REG_15__SCAN_IN;
  assign P1_U3543 = ~n23012 | ~n23011;
  assign n23025 = ~n23013 & ~n19083;
  assign n23023 = ~n23014 | ~n24216;
  assign n23021 = ~n23015 & ~n24241;
  assign n23019 = ~n23016 | ~n23953;
  assign n23018 = ~n23017 | ~n23988;
  assign n23020 = ~n23019 | ~n23018;
  assign n23022 = ~n23021 & ~n23020;
  assign n23024 = ~n23023 | ~n23022;
  assign n23028 = ~n23025 & ~n23024;
  assign n23027 = ~n23026 | ~n24011;
  assign n23105 = ~n23028 | ~n23027;
  assign n23030 = ~n23105 | ~n24286;
  assign n23029 = ~n24284 | ~P1_REG1_REG_14__SCAN_IN;
  assign P1_U3542 = ~n23030 | ~n23029;
  assign n23043 = ~n23031 & ~n19083;
  assign n23041 = ~n23032 | ~n24216;
  assign n23039 = ~n23033 & ~n24241;
  assign n23037 = ~n23034 | ~n23988;
  assign n23036 = ~n23035 | ~n23953;
  assign n23038 = ~n23037 | ~n23036;
  assign n23040 = ~n23039 & ~n23038;
  assign n23042 = ~n23041 | ~n23040;
  assign n23046 = ~n23043 & ~n23042;
  assign n23045 = ~n23044 | ~n24011;
  assign n23108 = ~n23046 | ~n23045;
  assign n23048 = ~n23108 | ~n24286;
  assign n23047 = ~n24284 | ~P1_REG1_REG_13__SCAN_IN;
  assign P1_U3541 = ~n23048 | ~n23047;
  assign n23055 = ~n23049 & ~n24220;
  assign n23053 = ~n23050 | ~n24216;
  assign n23052 = ~n23051 | ~n24230;
  assign n23054 = ~n23053 | ~n23052;
  assign n23056 = ~n23055 & ~n23054;
  assign n23111 = ~n23057 | ~n23056;
  assign n23059 = ~n23111 | ~n24286;
  assign n23058 = ~n24284 | ~P1_REG1_REG_11__SCAN_IN;
  assign P1_U3539 = ~n23059 | ~n23058;
  assign n23062 = ~n23060 | ~n24251;
  assign n23061 = ~n24240 | ~P1_REG0_REG_31__SCAN_IN;
  assign P1_U3527 = ~n23062 | ~n23061;
  assign n23065 = ~n23063 | ~n24251;
  assign n23064 = ~n24240 | ~P1_REG0_REG_30__SCAN_IN;
  assign P1_U3526 = ~n23065 | ~n23064;
  assign n23068 = ~n23066 | ~n24251;
  assign n23067 = ~n24240 | ~P1_REG0_REG_27__SCAN_IN;
  assign P1_U3523 = ~n23068 | ~n23067;
  assign n23071 = ~n23069 | ~n24251;
  assign n23070 = ~n24240 | ~P1_REG0_REG_26__SCAN_IN;
  assign P1_U3522 = ~n23071 | ~n23070;
  assign n23074 = ~n23072 | ~n24251;
  assign n23073 = ~n24240 | ~P1_REG0_REG_25__SCAN_IN;
  assign P1_U3521 = ~n23074 | ~n23073;
  assign n23077 = ~n23075 | ~n24251;
  assign n23076 = ~n24240 | ~P1_REG0_REG_24__SCAN_IN;
  assign P1_U3520 = ~n23077 | ~n23076;
  assign n23080 = ~n23078 | ~n24251;
  assign n23079 = ~n24240 | ~P1_REG0_REG_23__SCAN_IN;
  assign P1_U3519 = ~n23080 | ~n23079;
  assign n23083 = ~n23081 | ~n24251;
  assign n23082 = ~n24240 | ~P1_REG0_REG_22__SCAN_IN;
  assign P1_U3518 = ~n23083 | ~n23082;
  assign n23086 = ~n23084 | ~n24251;
  assign n23085 = ~n24240 | ~P1_REG0_REG_21__SCAN_IN;
  assign P1_U3517 = ~n23086 | ~n23085;
  assign n23089 = ~n23087 | ~n24251;
  assign n23088 = ~n24240 | ~P1_REG0_REG_20__SCAN_IN;
  assign P1_U3516 = ~n23089 | ~n23088;
  assign n23092 = ~n23090 | ~n24251;
  assign n23091 = ~n24240 | ~P1_REG0_REG_19__SCAN_IN;
  assign P1_U3515 = ~n23092 | ~n23091;
  assign n23095 = ~n23093 | ~n24251;
  assign n23094 = ~n24240 | ~P1_REG0_REG_18__SCAN_IN;
  assign P1_U3513 = ~n23095 | ~n23094;
  assign n23098 = ~n23096 | ~n24251;
  assign n23097 = ~n24240 | ~P1_REG0_REG_17__SCAN_IN;
  assign P1_U3510 = ~n23098 | ~n23097;
  assign n23101 = ~n23099 | ~n24251;
  assign n23100 = ~n24240 | ~P1_REG0_REG_16__SCAN_IN;
  assign P1_U3507 = ~n23101 | ~n23100;
  assign n23104 = ~n23102 | ~n24251;
  assign n23103 = ~n24240 | ~P1_REG0_REG_15__SCAN_IN;
  assign P1_U3504 = ~n23104 | ~n23103;
  assign n23107 = ~n23105 | ~n24251;
  assign n23106 = ~n24240 | ~P1_REG0_REG_14__SCAN_IN;
  assign P1_U3501 = ~n23107 | ~n23106;
  assign n23110 = ~n23108 | ~n24251;
  assign n23109 = ~n24240 | ~P1_REG0_REG_13__SCAN_IN;
  assign P1_U3498 = ~n23110 | ~n23109;
  assign n23113 = ~n23111 | ~n24251;
  assign n23112 = ~n24240 | ~P1_REG0_REG_11__SCAN_IN;
  assign P1_U3492 = ~n23113 | ~n23112;
  assign n23122 = ~n23114 | ~n23156;
  assign n23115 = ~n15904 & ~P1_IR_REG_30__SCAN_IN;
  assign n23116 = ~n23115 | ~P1_STATE_REG_SCAN_IN;
  assign n23120 = ~n23117 & ~n23116;
  assign n23119 = ~n24085 & ~n23118;
  assign n23121 = ~n23120 & ~n23119;
  assign P1_U3324 = ~n23122 | ~n23121;
  assign n23129 = ~n23123 | ~n23156;
  assign n23127 = ~n23124 & ~P1_U3086;
  assign n23126 = ~n24085 & ~n23125;
  assign n23128 = ~n23127 & ~n23126;
  assign P1_U3325 = ~n23129 | ~n23128;
  assign n23131 = ~n23130;
  assign n23136 = ~n23131 & ~n24106;
  assign n23134 = n23132 | P1_U3086;
  assign n23133 = ~n24110 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n23135 = ~n23134 | ~n23133;
  assign P1_U3326 = n23136 | n23135;
  assign n23138 = ~n23137;
  assign n23142 = ~n23138 & ~n24106;
  assign n23140 = n23351 | P1_U3086;
  assign n23139 = ~n24110 | ~P2_DATAO_REG_28__SCAN_IN;
  assign n23141 = ~n23140 | ~n23139;
  assign P1_U3327 = n23142 | n23141;
  assign n23148 = ~n23143 | ~n23156;
  assign n23146 = ~n16818 & ~P1_U3086;
  assign n23145 = ~n24085 & ~n23144;
  assign n23147 = ~n23146 & ~n23145;
  assign P1_U3328 = ~n23148 | ~n23147;
  assign n23155 = ~n23149 | ~n23156;
  assign n23150 = ~n15865;
  assign n23153 = ~n23150 & ~P1_U3086;
  assign n23152 = ~n24085 & ~n23151;
  assign n23154 = ~n23153 & ~n23152;
  assign P1_U3329 = ~n23155 | ~n23154;
  assign n23163 = ~n23157 | ~n23156;
  assign n23158 = ~n15901;
  assign n23161 = ~n23158 & ~P1_U3086;
  assign n23160 = ~n24085 & ~n23159;
  assign n23162 = ~n23161 & ~n23160;
  assign P1_U3330 = ~n23163 | ~n23162;
  assign n23165 = ~n23164;
  assign n23170 = ~n23165 | ~n23166;
  assign n23168 = ~n23167 | ~n23166;
  assign n23169 = ~n23168 | ~P2_ADDR_REG_11__SCAN_IN;
  assign SUB_1596_U69 = ~n23170 | ~n23169;
  assign n23172 = ~n23171;
  assign n23177 = ~n23172 | ~n23173;
  assign n23175 = ~n23174 | ~n23173;
  assign n23176 = ~n23175 | ~P2_ADDR_REG_12__SCAN_IN;
  assign SUB_1596_U68 = ~n23177 | ~n23176;
  assign n23179 = ~n23178;
  assign n23182 = ~n23181 | ~P2_ADDR_REG_13__SCAN_IN;
  assign SUB_1596_U67 = ~n23183 | ~n23182;
  assign n23186 = ~n23185 | ~n23184;
  assign SUB_1596_U66 = n23186 ^ ~P2_ADDR_REG_14__SCAN_IN;
  assign SUB_1596_U65 = n23188 ^ ~P2_ADDR_REG_15__SCAN_IN;
  assign n23190 = ~n23189;
  assign n23195 = ~n23190 | ~n23191;
  assign n23193 = ~n23192 | ~n23191;
  assign n23194 = ~n23193 | ~P2_ADDR_REG_16__SCAN_IN;
  assign SUB_1596_U64 = ~n23195 | ~n23194;
  assign n23196 = ~n13184;
  assign n23200 = ~n23197 | ~n23196;
  assign n23199 = n13184 | n23198;
  assign n23202 = ~n23343 | ~n23815;
  assign n23201 = ~n23322 | ~n23875;
  assign n23209 = ~n23202 | ~n23201;
  assign n23205 = ~n23204 & ~n23203;
  assign n23206 = ~n23205 & ~n23309;
  assign n23208 = n23207 & n23206;
  assign n23214 = ~n23209 & ~n23208;
  assign n24203 = ~n23818;
  assign n23212 = ~n23277 & ~n24203;
  assign n23210 = ~n23332 | ~n23825;
  assign n23471 = ~P1_REG3_REG_7__SCAN_IN | ~P1_U3086;
  assign n23211 = ~n23210 | ~n23471;
  assign n23213 = ~n23212 & ~n23211;
  assign P1_U3213 = ~n23214 | ~n23213;
  assign n23216 = ~n23988 | ~n23254;
  assign n23215 = ~n23953 | ~n23874;
  assign n23927 = ~n23216 | ~n23215;
  assign n23218 = ~n23217 | ~n23927;
  assign n23229 = ~n23219 | ~n23218;
  assign n23223 = n23221 & n23220;
  assign n23224 = ~n23223 & ~n23222;
  assign n23227 = ~n23224 & ~n23309;
  assign n23226 = n23225;
  assign n23228 = n23227 & n23226;
  assign n23233 = ~n23229 & ~n23228;
  assign n23231 = ~n23277 & ~n24155;
  assign n23230 = ~P1_REG3_REG_3__SCAN_IN & ~n23311;
  assign n23232 = ~n23231 & ~n23230;
  assign P1_U3218 = ~n23233 | ~n23232;
  assign n23236 = ~n23329 & ~n23234;
  assign n23491 = ~P1_STATE_REG_SCAN_IN & ~n23235;
  assign n23249 = ~n23236 & ~n23491;
  assign n23239 = n23238 ^ ~n23237;
  assign n23245 = ~n23239 | ~n23339;
  assign n23240 = ~n24213;
  assign n23243 = ~n23277 & ~n23240;
  assign n23242 = ~n23279 & ~n23241;
  assign n23244 = ~n23243 & ~n23242;
  assign n23247 = ~n23245 | ~n23244;
  assign n23246 = ~n23805 & ~n23311;
  assign n23248 = ~n23247 & ~n23246;
  assign P1_U3221 = ~n23249 | ~n23248;
  assign n23251 = n23250;
  assign n23253 = n23252 ^ ~n23251;
  assign n23262 = ~n23253 | ~n23339;
  assign n23256 = ~n23332 | ~n23254;
  assign n23255 = ~n23322 | ~n23993;
  assign n23260 = ~n23256 | ~n23255;
  assign n23258 = ~P1_REG3_REG_1__SCAN_IN | ~n23319;
  assign n23257 = ~n23331 | ~n17352;
  assign n23259 = ~n23258 | ~n23257;
  assign n23261 = ~n23260 & ~n23259;
  assign P1_U3222 = ~n23262 | ~n23261;
  assign n23263 = ~n23322 | ~n23874;
  assign n23429 = ~P1_REG3_REG_5__SCAN_IN | ~P1_U3086;
  assign n23285 = ~n23263 | ~n23429;
  assign n23270 = ~n23226 | ~n23264;
  assign n23268 = ~n15167 | ~n23265;
  assign n23267 = ~n15823 | ~n23266;
  assign n23269 = n23268 & n23267;
  assign n23291 = ~n23270 | ~n23269;
  assign n23273 = ~n23291 | ~n23293;
  assign n23272 = ~n23271;
  assign n23290 = ~n23226 | ~n23272;
  assign n23275 = ~n23273 | ~n23290;
  assign n23276 = n23275 ^ ~n23274;
  assign n23283 = ~n23276 | ~n23339;
  assign n23281 = ~n23277 & ~n23872;
  assign n23280 = ~n23279 & ~n23278;
  assign n23282 = ~n23281 & ~n23280;
  assign n23284 = ~n23283 | ~n23282;
  assign n23287 = ~n23285 & ~n23284;
  assign n23286 = ~n23867 | ~n23343;
  assign P1_U3227 = ~n23287 | ~n23286;
  assign n23289 = ~n23331 | ~n23903;
  assign n23288 = ~n23332 | ~n23854;
  assign n23296 = ~n23289 | ~n23288;
  assign n23292 = ~n23291 | ~n23290;
  assign n23294 = n23293 ^ ~n23292;
  assign n23295 = ~n23294 & ~n23309;
  assign n23301 = ~n23296 & ~n23295;
  assign n23297 = ~n23322 | ~n17357;
  assign n23408 = ~P1_REG3_REG_4__SCAN_IN | ~P1_U3086;
  assign n23299 = ~n23297 | ~n23408;
  assign n23298 = ~n23919 & ~n23311;
  assign n23300 = ~n23299 & ~n23298;
  assign P1_U3230 = ~n23301 | ~n23300;
  assign n23302 = ~n23322 | ~n23825;
  assign n23519 = ~P1_REG3_REG_9__SCAN_IN | ~P1_U3086;
  assign n23306 = ~n23302 | ~n23519;
  assign n23304 = ~n23331 | ~n24231;
  assign n23303 = ~n23332 | ~n23769;
  assign n23305 = ~n23304 | ~n23303;
  assign n23315 = ~n23306 & ~n23305;
  assign n23310 = n23308 ^ n23307;
  assign n23313 = ~n23310 & ~n23309;
  assign n23312 = ~n23311 & ~n23789;
  assign n23314 = ~n23313 & ~n23312;
  assign P1_U3231 = ~n23315 | ~n23314;
  assign n23318 = n23317 ^ ~n23316;
  assign n23328 = ~n23318 | ~n23339;
  assign n23321 = ~P1_REG3_REG_2__SCAN_IN | ~n23319;
  assign n23320 = ~n23332 | ~n17357;
  assign n23326 = ~n23321 | ~n23320;
  assign n23324 = ~n23331 | ~n23967;
  assign n23323 = ~n23322 | ~n17382;
  assign n23325 = ~n23324 | ~n23323;
  assign n23327 = ~n23326 & ~n23325;
  assign P1_U3237 = ~n23328 | ~n23327;
  assign n23330 = ~n23329 & ~n23906;
  assign n23454 = ~P1_STATE_REG_SCAN_IN & ~n13538;
  assign n23349 = ~n23330 & ~n23454;
  assign n23334 = ~n23331 | ~n24190;
  assign n23333 = ~n23332 | ~n23853;
  assign n23347 = ~n23334 | ~n23333;
  assign n23335 = ~n23337;
  assign n23338 = ~n13147 | ~n23337;
  assign n23340 = ~n23336 | ~n23338;
  assign n23341 = ~n23340 | ~n23339;
  assign n23345 = n23342 | n23341;
  assign n23344 = ~n23343 | ~n23842;
  assign n23346 = ~n23345 | ~n23344;
  assign n23348 = ~n23347 & ~n23346;
  assign P1_U3239 = ~n23349 | ~n23348;
  assign n23358 = ~n23684 & ~n23350;
  assign n23352 = ~P1_REG2_REG_0__SCAN_IN & ~n16818;
  assign n23393 = ~n23352 & ~n23351;
  assign n23353 = ~n14946 | ~n16818;
  assign n23354 = ~n23393 | ~n23353;
  assign n23355 = P1_IR_REG_0__SCAN_IN ^ n23354;
  assign n23357 = ~n23356 & ~n23355;
  assign n23360 = ~n23358 & ~n23357;
  assign n23359 = ~P1_REG3_REG_0__SCAN_IN | ~P1_U3086;
  assign P1_U3243 = ~n23360 | ~n23359;
  assign n23362 = ~P1_ADDR_REG_1__SCAN_IN | ~n23729;
  assign n23361 = ~P1_REG3_REG_1__SCAN_IN | ~P1_U3086;
  assign n23370 = ~n23362 | ~n23361;
  assign n23365 = n23364 ^ ~n23363;
  assign n23368 = ~n23720 | ~n23365;
  assign n23367 = ~n23688 | ~n23366;
  assign n23369 = ~n23368 | ~n23367;
  assign n23377 = ~n23370 & ~n23369;
  assign n23373 = ~n23372 | ~n23371;
  assign n23375 = n23374 & n23373;
  assign n23376 = ~n23722 | ~n23375;
  assign P1_U3244 = ~n23377 | ~n23376;
  assign n23379 = ~P1_ADDR_REG_2__SCAN_IN | ~n23729;
  assign n23378 = ~P1_REG3_REG_2__SCAN_IN | ~P1_U3086;
  assign n23387 = ~n23379 | ~n23378;
  assign n23385 = ~n23688 | ~n23380;
  assign n23383 = n23382 ^ n23381;
  assign n23384 = ~n23722 | ~n23383;
  assign n23386 = ~n23385 | ~n23384;
  assign n23406 = ~n23387 & ~n23386;
  assign n23388 = ~n23391 | ~n16818;
  assign n23398 = ~n23389 & ~n23388;
  assign n24307 = ~n24319;
  assign n23392 = ~n23391 | ~n23390;
  assign n23395 = ~n16818 & ~n23392;
  assign n23394 = ~P1_IR_REG_0__SCAN_IN & ~n23393;
  assign n23396 = ~n23395 & ~n23394;
  assign n23397 = ~n24307 | ~n23396;
  assign n23425 = ~n23398 & ~n23397;
  assign n23403 = ~n23720 | ~n23399;
  assign n23402 = ~n23401 & ~n23400;
  assign n23404 = ~n23403 & ~n23402;
  assign n23405 = ~n23425 & ~n23404;
  assign P1_U3245 = ~n23406 | ~n23405;
  assign n23407 = ~P1_ADDR_REG_4__SCAN_IN | ~n23729;
  assign n23423 = ~n23408 | ~n23407;
  assign n23445 = n24101 ^ ~P1_REG2_REG_4__SCAN_IN;
  assign n23412 = ~n23410 | ~n23409;
  assign n23411 = ~n23416 | ~P1_REG2_REG_3__SCAN_IN;
  assign n23446 = ~n23412 | ~n23411;
  assign n23413 = n23445 ^ n23446;
  assign n23421 = ~n23413 | ~n23720;
  assign n23418 = ~n23415 | ~n23414;
  assign n23417 = ~n23416 | ~P1_REG1_REG_3__SCAN_IN;
  assign n23431 = ~n23418 | ~n23417;
  assign n23430 = n24101 ^ ~P1_REG1_REG_4__SCAN_IN;
  assign n23419 = n23431 ^ n23430;
  assign n23420 = ~n23722 | ~n23419;
  assign n23422 = ~n23421 | ~n23420;
  assign n23427 = ~n23423 & ~n23422;
  assign n23424 = ~n23724 & ~n24101;
  assign n23426 = ~n23425 & ~n23424;
  assign P1_U3247 = ~n23427 | ~n23426;
  assign n23428 = ~P1_ADDR_REG_5__SCAN_IN | ~n23729;
  assign n23443 = ~n23429 | ~n23428;
  assign n23457 = ~n23444;
  assign n23441 = ~n23688 | ~n23457;
  assign n23432 = ~P1_REG1_REG_4__SCAN_IN;
  assign n23433 = n24101 | n23432;
  assign n23434 = ~P1_REG1_REG_5__SCAN_IN;
  assign n23463 = ~n23444 | ~n23434;
  assign n23435 = n23444 | n23434;
  assign n23436 = ~n23463 | ~n23435;
  assign n23438 = ~n23437 | ~n23436;
  assign n23439 = ~n23464 | ~n23438;
  assign n23440 = ~n23722 | ~n23439;
  assign n23442 = ~n23441 | ~n23440;
  assign n23452 = ~n23443 & ~n23442;
  assign n23455 = n23444 ^ ~P1_REG2_REG_5__SCAN_IN;
  assign n23449 = ~n23446 | ~n23445;
  assign n23447 = ~n24101;
  assign n23448 = ~n23447 | ~P1_REG2_REG_4__SCAN_IN;
  assign n23456 = ~n23449 | ~n23448;
  assign n23450 = n23455 ^ n23456;
  assign n23451 = ~n23720 | ~n23450;
  assign P1_U3248 = ~n23452 | ~n23451;
  assign n23453 = n23729 & P1_ADDR_REG_6__SCAN_IN;
  assign n23469 = ~n23454 & ~n23453;
  assign n23474 = ~n24096;
  assign n23462 = ~n23688 | ~n23474;
  assign n23472 = n24096 ^ ~P1_REG2_REG_6__SCAN_IN;
  assign n23459 = ~n23456 | ~n23455;
  assign n23458 = ~n23457 | ~P1_REG2_REG_5__SCAN_IN;
  assign n23473 = ~n23459 | ~n23458;
  assign n23460 = n23472 ^ n23473;
  assign n23461 = ~n23460 | ~n23720;
  assign n23467 = ~n23462 | ~n23461;
  assign n23484 = ~P1_REG1_REG_6__SCAN_IN;
  assign n23482 = n24096 ^ ~n23484;
  assign n23465 = n23483 ^ ~n23482;
  assign n23466 = ~n23501 & ~n23465;
  assign n23468 = ~n23467 & ~n23466;
  assign P1_U3249 = ~n23469 | ~n23468;
  assign n23470 = ~P1_ADDR_REG_7__SCAN_IN | ~n23729;
  assign n23481 = ~n23471 | ~n23470;
  assign n23476 = ~n23473 | ~n23472;
  assign n23475 = ~n23474 | ~P1_REG2_REG_6__SCAN_IN;
  assign n23508 = ~n23476 | ~n23475;
  assign n23506 = P1_REG2_REG_7__SCAN_IN ^ n23486;
  assign n23477 = n23508 ^ ~n23506;
  assign n23479 = ~n23720 | ~n23477;
  assign n23509 = ~n23486;
  assign n23478 = ~n23688 | ~n23509;
  assign n23480 = ~n23479 | ~n23478;
  assign n23489 = ~n23481 & ~n23480;
  assign n23485 = n24096 | n23484;
  assign n23492 = n23486 ^ ~P1_REG1_REG_7__SCAN_IN;
  assign n23487 = n23493 ^ n23492;
  assign n23488 = ~n23722 | ~n23487;
  assign P1_U3250 = ~n23489 | ~n23488;
  assign n23490 = P1_ADDR_REG_8__SCAN_IN & n23729;
  assign n23505 = n23491 | n23490;
  assign n23494 = ~n23509 | ~P1_REG1_REG_7__SCAN_IN;
  assign n23495 = ~P1_REG1_REG_8__SCAN_IN;
  assign n23515 = ~n24091 | ~n23495;
  assign n23496 = n24091 | n23495;
  assign n23497 = n23515 & n23496;
  assign n23498 = ~n23497;
  assign n23499 = ~n13403 | ~n23498;
  assign n23500 = n23516 & n23499;
  assign n23503 = n23501 | n23500;
  assign n23502 = n23724 | n24091;
  assign n23504 = ~n23503 | ~n23502;
  assign n23514 = ~n23505 & ~n23504;
  assign n23520 = n24091 ^ ~P1_REG2_REG_8__SCAN_IN;
  assign n23507 = ~n23506;
  assign n23511 = ~n23508 | ~n23507;
  assign n23510 = ~n23509 | ~P1_REG2_REG_7__SCAN_IN;
  assign n23521 = ~n23511 | ~n23510;
  assign n23512 = n23520 ^ n23521;
  assign n23513 = ~n23720 | ~n23512;
  assign P1_U3251 = ~n23514 | ~n23513;
  assign n23540 = P1_REG1_REG_9__SCAN_IN ^ ~n24088;
  assign n23517 = n23541 ^ ~n23540;
  assign n23531 = ~n23517 | ~n23722;
  assign n23518 = ~P1_ADDR_REG_9__SCAN_IN | ~n23729;
  assign n23529 = ~n23519 | ~n23518;
  assign n23536 = P1_REG2_REG_9__SCAN_IN ^ n24088;
  assign n23524 = ~n23521 | ~n23520;
  assign n23522 = ~n24091;
  assign n23523 = ~n23522 | ~P1_REG2_REG_8__SCAN_IN;
  assign n23535 = ~n23524 | ~n23523;
  assign n23525 = n23536 ^ n23535;
  assign n23527 = ~n23525 | ~n23720;
  assign n23526 = ~n23688 | ~n24088;
  assign n23528 = ~n23527 | ~n23526;
  assign n23530 = ~n23529 & ~n23528;
  assign P1_U3252 = ~n23531 | ~n23530;
  assign n23533 = ~n23532 & ~n23684;
  assign n23551 = ~n23534 & ~n23533;
  assign n23547 = ~n24081;
  assign n23559 = P1_REG2_REG_10__SCAN_IN ^ ~n23547;
  assign n23538 = ~P1_REG2_REG_9__SCAN_IN | ~n24088;
  assign n23537 = ~n23536 | ~n23535;
  assign n23558 = ~n23538 | ~n23537;
  assign n23539 = n23559 ^ n23558;
  assign n23546 = ~n23539 | ~n23720;
  assign n23553 = P1_REG1_REG_10__SCAN_IN ^ ~n23547;
  assign n23543 = ~P1_REG1_REG_9__SCAN_IN & ~n24088;
  assign n23542 = ~n23541 & ~n23540;
  assign n23544 = n23553 ^ n23552;
  assign n23545 = ~n23544 | ~n23722;
  assign n23549 = ~n23546 | ~n23545;
  assign n23548 = ~n23724 & ~n23547;
  assign n23550 = ~n23549 & ~n23548;
  assign P1_U3253 = ~n23551 | ~n23550;
  assign n23582 = P1_REG1_REG_11__SCAN_IN ^ ~n24075;
  assign n23554 = ~P1_REG1_REG_10__SCAN_IN | ~n24081;
  assign n23555 = n23582 ^ ~n23583;
  assign n23568 = ~n23555 | ~n23722;
  assign n23556 = ~P1_ADDR_REG_11__SCAN_IN | ~n23729;
  assign n23566 = ~n23557 | ~n23556;
  assign n23570 = P1_REG2_REG_11__SCAN_IN ^ n24075;
  assign n23561 = ~P1_REG2_REG_10__SCAN_IN | ~n24081;
  assign n23560 = ~n23559 | ~n23558;
  assign n23569 = ~n23561 | ~n23560;
  assign n23562 = n23570 ^ n23569;
  assign n23564 = ~n23562 | ~n23720;
  assign n23563 = ~n23688 | ~n24075;
  assign n23565 = ~n23564 | ~n23563;
  assign n23567 = ~n23566 & ~n23565;
  assign P1_U3254 = ~n23568 | ~n23567;
  assign n23579 = ~n24069;
  assign n23591 = P1_REG2_REG_12__SCAN_IN ^ n23579;
  assign n23572 = ~P1_REG2_REG_11__SCAN_IN | ~n24075;
  assign n23571 = ~n23570 | ~n23569;
  assign n23592 = ~n23572 | ~n23571;
  assign n23573 = n23591 ^ ~n23592;
  assign n23578 = ~n23573 | ~n23720;
  assign n23575 = ~n23574 & ~n23684;
  assign n23577 = ~n23576 & ~n23575;
  assign n23581 = ~n23578 | ~n23577;
  assign n23580 = ~n23724 & ~n23579;
  assign n23588 = ~n23581 & ~n23580;
  assign n23584 = ~P1_REG1_REG_11__SCAN_IN & ~n24075;
  assign n23598 = ~P1_REG1_REG_12__SCAN_IN & ~n24069;
  assign n23597 = P1_REG1_REG_12__SCAN_IN & n24069;
  assign n23585 = ~n23598 & ~n23597;
  assign n23586 = n23596 ^ n23585;
  assign n23587 = ~n23586 | ~n23722;
  assign P1_U3255 = ~n23588 | ~n23587;
  assign n23589 = ~P1_ADDR_REG_13__SCAN_IN | ~n23729;
  assign n23603 = ~n23590 | ~n23589;
  assign n23613 = P1_REG2_REG_13__SCAN_IN ^ n24062;
  assign n23594 = ~P1_REG2_REG_12__SCAN_IN & ~n24069;
  assign n23593 = ~n23592 & ~n23591;
  assign n23612 = ~n23594 & ~n23593;
  assign n23595 = n23613 ^ n23612;
  assign n23601 = ~n23595 | ~n23720;
  assign n23622 = P1_REG1_REG_13__SCAN_IN ^ n24062;
  assign n23599 = n23623 ^ n23622;
  assign n23600 = ~n23599 | ~n23722;
  assign n23602 = ~n23601 | ~n23600;
  assign n23605 = ~n23603 & ~n23602;
  assign n23604 = ~n23688 | ~n24062;
  assign P1_U3256 = ~n23605 | ~n23604;
  assign n23607 = ~n23606 & ~n23684;
  assign n23610 = ~n23608 & ~n23607;
  assign n23609 = ~n23688 | ~n24056;
  assign n23621 = ~n23610 | ~n23609;
  assign n23611 = ~n24056;
  assign n23617 = P1_REG2_REG_14__SCAN_IN ^ ~n23611;
  assign n23615 = ~P1_REG2_REG_13__SCAN_IN | ~n24062;
  assign n23614 = ~n23613 | ~n23612;
  assign n23616 = ~n23615 | ~n23614;
  assign n23636 = ~n23617 | ~n23616;
  assign n23619 = ~n23720 | ~n23636;
  assign n23618 = ~n23617 & ~n23616;
  assign n23620 = ~n23619 & ~n23618;
  assign n23628 = ~n23621 & ~n23620;
  assign n23631 = ~P1_REG1_REG_14__SCAN_IN & ~n24056;
  assign n23630 = P1_REG1_REG_14__SCAN_IN & n24056;
  assign n23625 = ~n23631 & ~n23630;
  assign n23624 = ~P1_REG1_REG_13__SCAN_IN | ~n24062;
  assign n23626 = n23625 ^ n23629;
  assign n23627 = ~n23626 | ~n23722;
  assign P1_U3257 = ~n23628 | ~n23627;
  assign n23633 = n23657 ^ ~P1_REG1_REG_15__SCAN_IN;
  assign n23644 = ~n23633 | ~n23722;
  assign n23634 = ~P1_ADDR_REG_15__SCAN_IN | ~n23729;
  assign n23642 = ~n23635 | ~n23634;
  assign n23637 = ~P1_REG2_REG_14__SCAN_IN | ~n24056;
  assign n23648 = ~n23637 | ~n23636;
  assign n23649 = n23648 ^ ~n23656;
  assign n23638 = n23649 ^ ~P1_REG2_REG_15__SCAN_IN;
  assign n23640 = ~n23638 | ~n23720;
  assign n23639 = ~n23688 | ~n23656;
  assign n23641 = ~n23640 | ~n23639;
  assign n23643 = ~n23642 & ~n23641;
  assign P1_U3258 = ~n23644 | ~n23643;
  assign n23646 = ~n23645 & ~n23684;
  assign n23666 = ~n23647 & ~n23646;
  assign n24047 = ~n23678;
  assign n23670 = P1_REG2_REG_16__SCAN_IN ^ ~n24047;
  assign n23651 = ~n23656 & ~n23648;
  assign n23650 = ~P1_REG2_REG_15__SCAN_IN & ~n23649;
  assign n23669 = ~n23651 & ~n23650;
  assign n23652 = n23670 ^ n23669;
  assign n23654 = ~n23652 | ~n23720;
  assign n23653 = ~n23688 | ~n23678;
  assign n23664 = ~n23654 | ~n23653;
  assign n23659 = P1_REG1_REG_16__SCAN_IN ^ ~n24047;
  assign n23658 = ~n23656 & ~n23655;
  assign n23679 = ~n23659 | ~n23660;
  assign n23662 = ~n23679 | ~n23722;
  assign n23661 = ~n23660 & ~n23659;
  assign n23663 = ~n23662 & ~n23661;
  assign n23665 = ~n23664 & ~n23663;
  assign P1_U3259 = ~n23666 | ~n23665;
  assign n23667 = ~P1_ADDR_REG_17__SCAN_IN | ~n23729;
  assign n23677 = ~n23668 | ~n23667;
  assign n23692 = P1_REG2_REG_17__SCAN_IN ^ n24044;
  assign n23672 = ~P1_REG2_REG_16__SCAN_IN | ~n23678;
  assign n23671 = ~n23670 | ~n23669;
  assign n23691 = ~n23672 | ~n23671;
  assign n23673 = n23692 ^ n23691;
  assign n23675 = ~n23673 | ~n23720;
  assign n23674 = ~n23688 | ~n24044;
  assign n23676 = ~n23675 | ~n23674;
  assign n23683 = ~n23677 & ~n23676;
  assign n23701 = P1_REG1_REG_17__SCAN_IN ^ n24044;
  assign n23680 = ~P1_REG1_REG_16__SCAN_IN | ~n23678;
  assign n23700 = ~n23680 | ~n23679;
  assign n23681 = n23701 ^ n23700;
  assign n23682 = ~n23681 | ~n23722;
  assign P1_U3260 = ~n23683 | ~n23682;
  assign n23686 = ~n23685 & ~n23684;
  assign n23690 = ~n23687 & ~n23686;
  assign n23689 = ~n23688 | ~n23711;
  assign n23699 = ~n23690 | ~n23689;
  assign n24036 = ~n23711;
  assign n23694 = ~P1_REG2_REG_17__SCAN_IN | ~n24044;
  assign n23693 = ~n23692 | ~n23691;
  assign n23710 = ~n23694 | ~n23693;
  assign n23695 = n24036 ^ ~n23710;
  assign n23713 = ~P1_REG2_REG_18__SCAN_IN | ~n23695;
  assign n23697 = ~n23720 | ~n23713;
  assign n23696 = ~n23695 & ~P1_REG2_REG_18__SCAN_IN;
  assign n23698 = ~n23697 & ~n23696;
  assign n23705 = ~n23699 & ~n23698;
  assign n23702 = ~P1_REG1_REG_17__SCAN_IN | ~n24044;
  assign n23703 = P1_REG1_REG_18__SCAN_IN ^ n23707;
  assign n23704 = ~n23703 | ~n23722;
  assign P1_U3261 = ~n23705 | ~n23704;
  assign n23709 = ~n23711 | ~n23706;
  assign n23717 = ~n23721 | ~n23722;
  assign n23712 = ~n23711 | ~n23710;
  assign n23714 = ~n23713 | ~n23712;
  assign n23718 = P1_REG2_REG_19__SCAN_IN ^ n23714;
  assign n23715 = ~n23720 | ~n23718;
  assign n23716 = n23715 & n23905;
  assign n23728 = ~n23717 | ~n23716;
  assign n23719 = ~n23718;
  assign n23727 = ~n23720 | ~n23719;
  assign n23725 = n23724 & n23723;
  assign n23730 = ~n23729 | ~P1_ADDR_REG_19__SCAN_IN;
  assign n23734 = ~n23980 & ~n24242;
  assign n23733 = ~n23936 & ~n23732;
  assign n23736 = ~n23734 & ~n23733;
  assign n23735 = ~P1_REG2_REG_10__SCAN_IN | ~n24021;
  assign n23761 = ~n23736 | ~n23735;
  assign n23738 = ~n23737;
  assign n23774 = ~n23738 | ~n23777;
  assign n23741 = ~n23774 | ~n23739;
  assign n23742 = n23741 ^ ~n23740;
  assign n23744 = ~n23742 | ~n24011;
  assign n23743 = ~n23988 | ~n23801;
  assign n24246 = ~n23744 | ~n23743;
  assign n23747 = n23746 | n23745;
  assign n24248 = ~n23748 | ~n23747;
  assign n23757 = ~n24248 | ~n24012;
  assign n23750 = n23749 | n24242;
  assign n23752 = n23750 & n24216;
  assign n23755 = ~n23752 | ~n23751;
  assign n23754 = ~n23953 | ~n23753;
  assign n24244 = ~n23755 | ~n23754;
  assign n23756 = ~n24244 | ~n23905;
  assign n23758 = ~n23757 | ~n23756;
  assign n23759 = ~n24246 & ~n23758;
  assign n23760 = ~n24021 & ~n23759;
  assign n23764 = ~n23761 & ~n23760;
  assign n23762 = ~n23892;
  assign n23763 = ~n24248 | ~n23762;
  assign P1_U3283 = ~n23764 | ~n23763;
  assign n23766 = n23765 ^ ~n13914;
  assign n24235 = ~n23766 & ~n24201;
  assign n23768 = ~n24235 | ~n23905;
  assign n23767 = ~n24231 | ~n23966;
  assign n23787 = ~n23768 | ~n23767;
  assign n23771 = ~n23988 | ~n23825;
  assign n23770 = ~n23953 | ~n23769;
  assign n23784 = ~n23771 | ~n23770;
  assign n23773 = ~n23737 | ~n23772;
  assign n23775 = ~n23774 | ~n23773;
  assign n23782 = ~n23775 | ~n24011;
  assign n23778 = ~n22775 | ~n23776;
  assign n23779 = ~n23778 | ~n23777;
  assign n24229 = ~n23780 | ~n23779;
  assign n23781 = ~n24229 | ~n24012;
  assign n23783 = ~n23782 | ~n23781;
  assign n24237 = ~n23784 & ~n23783;
  assign n24009 = ~n23970;
  assign n23785 = ~n24229 | ~n24009;
  assign n23786 = ~n24237 | ~n23785;
  assign n23788 = ~n23787 & ~n23786;
  assign n23791 = ~n24021 & ~n23788;
  assign n23790 = ~n23936 & ~n23789;
  assign n23793 = ~n23791 & ~n23790;
  assign n23792 = ~P1_REG2_REG_9__SCAN_IN | ~n24021;
  assign P1_U3284 = ~n23793 | ~n23792;
  assign n23795 = n23794 ^ ~n23796;
  assign n23800 = ~n23795 & ~n23991;
  assign n23810 = n13396 ^ ~n23796;
  assign n23798 = ~n23810 | ~n24012;
  assign n23797 = ~n23988 | ~n23853;
  assign n23799 = ~n23798 | ~n23797;
  assign n24225 = ~n23800 & ~n23799;
  assign n24214 = ~n23953 | ~n23801;
  assign n23802 = ~n24225 | ~n24214;
  assign n23809 = ~n23802 | ~n24019;
  assign n23804 = ~n24025 | ~n24213;
  assign n23803 = ~n24021 | ~P1_REG2_REG_8__SCAN_IN;
  assign n23807 = ~n23804 | ~n23803;
  assign n23806 = ~n23805 & ~n23936;
  assign n23808 = ~n23807 & ~n23806;
  assign n23812 = ~n23809 | ~n23808;
  assign n24221 = ~n23810;
  assign n23811 = ~n24221 & ~n23892;
  assign n23814 = ~n23812 & ~n23811;
  assign n24217 = n23820 ^ n24213;
  assign n23813 = ~n24217 | ~n24026;
  assign P1_U3285 = ~n23814 | ~n23813;
  assign n23817 = ~n24022 | ~n23815;
  assign n23816 = ~n24021 | ~P1_REG2_REG_7__SCAN_IN;
  assign n23822 = ~n23817 | ~n23816;
  assign n23819 = ~n13407 | ~n23818;
  assign n24202 = ~n23820 | ~n23819;
  assign n23821 = ~n24202 & ~n23944;
  assign n23841 = ~n23822 & ~n23821;
  assign n23824 = n23823 ^ ~n23831;
  assign n23835 = ~n23824 | ~n24011;
  assign n23827 = ~n23988 | ~n23875;
  assign n23826 = ~n23953 | ~n23825;
  assign n23833 = ~n23827 | ~n23826;
  assign n23830 = n23829 & n23828;
  assign n24206 = n23831 ^ n23830;
  assign n23832 = ~n24206 & ~n18061;
  assign n23834 = ~n23833 & ~n23832;
  assign n24208 = ~n23835 | ~n23834;
  assign n23836 = ~n24203 & ~n23931;
  assign n23837 = ~n24208 & ~n23836;
  assign n23839 = ~n24021 & ~n23837;
  assign n23838 = ~n24206 & ~n23892;
  assign n23840 = ~n23839 & ~n23838;
  assign P1_U3286 = ~n23841 | ~n23840;
  assign n23844 = ~n24022 | ~n23842;
  assign n23843 = ~n24021 | ~P1_REG2_REG_6__SCAN_IN;
  assign n23847 = ~n23844 | ~n23843;
  assign n23846 = ~n23980 & ~n23845;
  assign n23866 = ~n23847 & ~n23846;
  assign n24189 = n23848 ^ ~n24190;
  assign n23862 = ~n24189 | ~n24026;
  assign n23850 = n23851 ^ n23849;
  assign n23860 = ~n23850 | ~n24011;
  assign n24195 = n23852 ^ ~n23851;
  assign n23858 = ~n24195 & ~n18061;
  assign n23856 = ~n23953 | ~n23853;
  assign n23855 = ~n23988 | ~n23854;
  assign n23857 = ~n23856 | ~n23855;
  assign n23859 = ~n23858 & ~n23857;
  assign n24194 = ~n23860 | ~n23859;
  assign n23861 = ~n24194 | ~n24019;
  assign n23864 = ~n23862 | ~n23861;
  assign n23863 = ~n24195 & ~n23892;
  assign n23865 = ~n23864 & ~n23863;
  assign P1_U3287 = ~n23866 | ~n23865;
  assign n23869 = ~n24022 | ~n23867;
  assign n23868 = ~n24021 | ~P1_REG2_REG_5__SCAN_IN;
  assign n23871 = ~n23869 | ~n23868;
  assign n23870 = ~n23980 & ~n23872;
  assign n23896 = ~n23871 & ~n23870;
  assign n24177 = n23873 ^ ~n23872;
  assign n23891 = ~n24026 | ~n24177;
  assign n23877 = ~n23988 | ~n23874;
  assign n23876 = ~n23953 | ~n23875;
  assign n23884 = ~n23877 | ~n23876;
  assign n23879 = ~n23910;
  assign n23912 = ~n23878 | ~n23879;
  assign n23881 = ~n23880;
  assign n23882 = ~n23912 | ~n23881;
  assign n24183 = n23882 ^ ~n23885;
  assign n23883 = ~n24183 & ~n18061;
  assign n23889 = ~n23884 & ~n23883;
  assign n23887 = n23886 ^ n23885;
  assign n23888 = ~n23887 | ~n24011;
  assign n24182 = ~n23889 | ~n23888;
  assign n23890 = ~n24182 | ~n24019;
  assign n23894 = ~n23891 | ~n23890;
  assign n23893 = ~n24183 & ~n23892;
  assign n23895 = ~n23894 & ~n23893;
  assign P1_U3288 = ~n23896 | ~n23895;
  assign n23899 = ~n23898 | ~n23897;
  assign n23900 = n23910 ^ n23899;
  assign n23902 = ~n23900 | ~n24011;
  assign n23901 = ~n23988 | ~n17357;
  assign n24174 = ~n23902 | ~n23901;
  assign n23904 = n23942 ^ ~n23903;
  assign n24169 = ~n23904 & ~n24201;
  assign n23909 = ~n24169 | ~n23905;
  assign n24167 = ~n23906 & ~n24014;
  assign n23907 = ~n23931 & ~n24165;
  assign n23908 = ~n24167 & ~n23907;
  assign n23916 = n23909 & n23908;
  assign n23911 = ~n23878;
  assign n23913 = ~n23911 | ~n23910;
  assign n24170 = ~n23913 | ~n23912;
  assign n23915 = ~n24170 | ~n23914;
  assign n23917 = ~n23916 | ~n23915;
  assign n23918 = ~n24174 & ~n23917;
  assign n23921 = ~n24021 & ~n23918;
  assign n23920 = ~n23936 & ~n23919;
  assign n23923 = ~n23921 & ~n23920;
  assign n23922 = ~P1_REG2_REG_4__SCAN_IN | ~n24021;
  assign P1_U3289 = ~n23923 | ~n23922;
  assign n23930 = ~n23925 | ~n24011;
  assign n23928 = ~n18061 & ~n24158;
  assign n23929 = ~n23928 & ~n23927;
  assign n24160 = ~n23930 | ~n23929;
  assign n23932 = ~n24155 & ~n23931;
  assign n23935 = ~n24160 & ~n23932;
  assign n23933 = ~n24158;
  assign n23934 = ~n23933 | ~n24009;
  assign n23938 = ~n23935 | ~n23934;
  assign n23937 = ~n23936 & ~P1_REG3_REG_3__SCAN_IN;
  assign n23939 = ~n23938 & ~n23937;
  assign n23946 = ~n24021 & ~n23939;
  assign n23943 = ~n14517 | ~n14281;
  assign n24154 = ~n23943 | ~n23942;
  assign n23945 = ~n23944 & ~n24154;
  assign n23948 = ~n23946 & ~n23945;
  assign n23947 = ~P1_REG2_REG_3__SCAN_IN | ~n24021;
  assign P1_U3290 = ~n23948 | ~n23947;
  assign n23951 = n23950 | n23958;
  assign n23952 = ~n23949 | ~n23951;
  assign n23962 = ~n23952 | ~n24011;
  assign n23955 = ~n23988 | ~n17382;
  assign n23954 = ~n23953 | ~n17357;
  assign n23960 = ~n23955 | ~n23954;
  assign n23956 = ~n23983;
  assign n23984 = ~n23990 & ~n23956;
  assign n23957 = ~n23984 & ~n18869;
  assign n24147 = n23958 ^ n23957;
  assign n23959 = ~n18061 & ~n24147;
  assign n23961 = ~n23960 & ~n23959;
  assign n24149 = ~n23962 | ~n23961;
  assign n23964 = ~n23967 | ~n23963;
  assign n24143 = ~n14517 | ~n23964;
  assign n23965 = ~n24143 & ~n24001;
  assign n23974 = ~n24149 & ~n23965;
  assign n23969 = ~n24022 | ~P1_REG3_REG_2__SCAN_IN;
  assign n23968 = ~n23967 | ~n23966;
  assign n23972 = ~n23969 | ~n23968;
  assign n23971 = ~n24147 & ~n23970;
  assign n23973 = ~n23972 & ~n23971;
  assign n23975 = ~n23974 | ~n23973;
  assign n23977 = ~n24019 | ~n23975;
  assign n23976 = ~n24021 | ~P1_REG2_REG_2__SCAN_IN;
  assign P1_U3291 = ~n23977 | ~n23976;
  assign n23979 = ~n24022 | ~P1_REG3_REG_1__SCAN_IN;
  assign n23978 = ~n24021 | ~P1_REG2_REG_1__SCAN_IN;
  assign n23982 = ~n23979 | ~n23978;
  assign n23981 = ~n23980 & ~n24131;
  assign n24008 = ~n23982 & ~n23981;
  assign n23986 = ~n23990;
  assign n23985 = ~n23986 & ~n23983;
  assign n23997 = ~n23985 & ~n23984;
  assign n24130 = ~n23997;
  assign n24005 = ~n24130 | ~n24009;
  assign n23987 = ~n23986 & ~n18544;
  assign n23989 = ~n23987 & ~n23991;
  assign n23996 = ~n23989 & ~n23988;
  assign n23992 = n23990 ^ ~n24027;
  assign n23994 = ~n23992 & ~n23991;
  assign n23995 = ~n23994 & ~n23993;
  assign n23999 = ~n23996 & ~n23995;
  assign n23998 = ~n23997 & ~n18061;
  assign n24140 = ~n23999 & ~n23998;
  assign n24133 = ~n24000 & ~n24014;
  assign n24134 = n17352 ^ ~n24122;
  assign n24002 = ~n24134 & ~n24001;
  assign n24003 = ~n24133 & ~n24002;
  assign n24004 = n24140 & n24003;
  assign n24006 = ~n24005 | ~n24004;
  assign n24007 = ~n24006 | ~n24019;
  assign P1_U3292 = ~n24008 | ~n24007;
  assign n24010 = ~n24121;
  assign n24018 = ~n24010 | ~n24009;
  assign n24013 = ~n24012 & ~n24011;
  assign n24017 = ~n24013 & ~n24121;
  assign n24016 = ~n24015 & ~n24014;
  assign n24127 = ~n24017 & ~n24016;
  assign n24020 = ~n24018 | ~n24127;
  assign n24032 = ~n24020 | ~n24019;
  assign n24024 = ~n24021 | ~P1_REG2_REG_0__SCAN_IN;
  assign n24023 = ~n24022 | ~P1_REG3_REG_0__SCAN_IN;
  assign n24030 = ~n24024 | ~n24023;
  assign n24028 = ~n24026 & ~n24025;
  assign n24029 = ~n24028 & ~n24027;
  assign n24031 = ~n24030 & ~n24029;
  assign P1_U3293 = ~n24032 | ~n24031;
  assign n24035 = ~n24033;
  assign n24116 = ~n24035 | ~n24034;
  assign P1_U3294 = P1_D_REG_31__SCAN_IN & n24116;
  assign P1_U3295 = P1_D_REG_30__SCAN_IN & n24116;
  assign P1_U3296 = P1_D_REG_29__SCAN_IN & n24116;
  assign P1_U3297 = P1_D_REG_28__SCAN_IN & n24116;
  assign P1_U3298 = P1_D_REG_27__SCAN_IN & n24116;
  assign P1_U3299 = P1_D_REG_26__SCAN_IN & n24116;
  assign P1_U3300 = P1_D_REG_25__SCAN_IN & n24116;
  assign P1_U3301 = P1_D_REG_24__SCAN_IN & n24116;
  assign P1_U3302 = P1_D_REG_23__SCAN_IN & n24116;
  assign P1_U3303 = P1_D_REG_22__SCAN_IN & n24116;
  assign P1_U3304 = P1_D_REG_21__SCAN_IN & n24116;
  assign P1_U3305 = P1_D_REG_20__SCAN_IN & n24116;
  assign P1_U3306 = P1_D_REG_19__SCAN_IN & n24116;
  assign P1_U3307 = P1_D_REG_18__SCAN_IN & n24116;
  assign P1_U3308 = P1_D_REG_17__SCAN_IN & n24116;
  assign P1_U3309 = P1_D_REG_16__SCAN_IN & n24116;
  assign P1_U3310 = P1_D_REG_15__SCAN_IN & n24116;
  assign P1_U3311 = P1_D_REG_14__SCAN_IN & n24116;
  assign P1_U3312 = P1_D_REG_13__SCAN_IN & n24116;
  assign P1_U3313 = P1_D_REG_12__SCAN_IN & n24116;
  assign P1_U3314 = P1_D_REG_11__SCAN_IN & n24116;
  assign P1_U3315 = P1_D_REG_10__SCAN_IN & n24116;
  assign P1_U3316 = P1_D_REG_9__SCAN_IN & n24116;
  assign P1_U3317 = P1_D_REG_8__SCAN_IN & n24116;
  assign P1_U3318 = P1_D_REG_7__SCAN_IN & n24116;
  assign P1_U3319 = P1_D_REG_6__SCAN_IN & n24116;
  assign P1_U3320 = P1_D_REG_5__SCAN_IN & n24116;
  assign P1_U3321 = P1_D_REG_4__SCAN_IN & n24116;
  assign P1_U3322 = P1_D_REG_3__SCAN_IN & n24116;
  assign P1_U3323 = P1_D_REG_2__SCAN_IN & n24116;
  assign n24038 = ~n25290 & ~n24106;
  assign n24037 = ~n24036 & ~P1_U3086;
  assign n24040 = ~n24038 & ~n24037;
  assign n24039 = ~n24110 | ~P2_DATAO_REG_18__SCAN_IN;
  assign P1_U3337 = ~n24040 | ~n24039;
  assign n24043 = ~n25296 & ~n24106;
  assign n24042 = ~n24085 & ~n24041;
  assign n24046 = ~n24043 & ~n24042;
  assign n24045 = ~n24044 | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3338 = ~n24046 | ~n24045;
  assign n24049 = ~n25302 & ~n24106;
  assign n24048 = ~n24047 & ~P1_U3086;
  assign n24051 = ~n24049 & ~n24048;
  assign n24050 = ~n24110 | ~P2_DATAO_REG_16__SCAN_IN;
  assign P1_U3339 = ~n24051 | ~n24050;
  assign n24055 = ~n24052 & ~n24106;
  assign n24054 = ~n24085 & ~n24053;
  assign n24058 = ~n24055 & ~n24054;
  assign n24057 = ~n24056 | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3341 = ~n24058 | ~n24057;
  assign n24061 = ~n25311 & ~n24106;
  assign n24060 = ~n24085 & ~n24059;
  assign n24064 = ~n24061 & ~n24060;
  assign n24063 = ~n24062 | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3342 = ~n24064 | ~n24063;
  assign n24068 = ~n24065 & ~n24106;
  assign n24067 = ~n24085 & ~n24066;
  assign n24071 = ~n24068 & ~n24067;
  assign n24070 = ~n24069 | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3343 = ~n24071 | ~n24070;
  assign n24074 = ~n25320 & ~n24106;
  assign n24073 = ~n24085 & ~n24072;
  assign n24077 = ~n24074 & ~n24073;
  assign n24076 = ~n24075 | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3344 = ~n24077 | ~n24076;
  assign n24080 = ~n25325 & ~n24106;
  assign n24079 = ~n24085 & ~n24078;
  assign n24083 = ~n24080 & ~n24079;
  assign n24082 = ~n24081 | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3345 = ~n24083 | ~n24082;
  assign n24087 = ~n25330 & ~n24106;
  assign n24086 = ~n24085 & ~n24084;
  assign n24090 = ~n24087 & ~n24086;
  assign n24089 = ~n24088 | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3346 = ~n24090 | ~n24089;
  assign n24093 = ~n25335 & ~n24106;
  assign n24092 = ~n24091 & ~P1_U3086;
  assign n24095 = ~n24093 & ~n24092;
  assign n24094 = ~n24110 | ~P2_DATAO_REG_8__SCAN_IN;
  assign P1_U3347 = ~n24095 | ~n24094;
  assign n24098 = ~n25348 & ~n24106;
  assign n24097 = ~n24096 & ~P1_U3086;
  assign n24100 = ~n24098 & ~n24097;
  assign n24099 = ~n24110 | ~P2_DATAO_REG_6__SCAN_IN;
  assign P1_U3349 = ~n24100 | ~n24099;
  assign n24103 = ~n25354 & ~n24106;
  assign n24102 = ~n24101 & ~P1_U3086;
  assign n24105 = ~n24103 & ~n24102;
  assign n24104 = ~n24110 | ~P2_DATAO_REG_4__SCAN_IN;
  assign P1_U3351 = ~n24105 | ~n24104;
  assign n24109 = ~n25361 & ~n24106;
  assign n24108 = ~n24107 & ~P1_U3086;
  assign n24112 = ~n24109 & ~n24108;
  assign n24111 = ~n24110 | ~P2_DATAO_REG_2__SCAN_IN;
  assign P1_U3353 = ~n24112 | ~n24111;
  assign n24115 = ~P1_D_REG_0__SCAN_IN | ~n24116;
  assign n24118 = ~n24116;
  assign n24114 = ~n24118 | ~n24113;
  assign P1_U3445 = ~n24115 | ~n24114;
  assign n24120 = ~P1_D_REG_1__SCAN_IN | ~n24116;
  assign n24119 = ~n24118 | ~n24117;
  assign P1_U3446 = ~n24120 | ~n24119;
  assign n24129 = ~P1_REG0_REG_0__SCAN_IN | ~n24240;
  assign n24125 = n24121 | n24220;
  assign n24124 = ~n24123 | ~n24122;
  assign n24126 = n24125 & n24124;
  assign n24254 = ~n24127 | ~n24126;
  assign n24128 = ~n24251 | ~n24254;
  assign P1_U3459 = ~n24129 | ~n24128;
  assign n24142 = ~P1_REG0_REG_1__SCAN_IN | ~n24240;
  assign n24138 = ~n24130 | ~n24228;
  assign n24132 = ~n24241 & ~n24131;
  assign n24136 = n24133 | n24132;
  assign n24135 = ~n24134 & ~n24201;
  assign n24137 = ~n24136 & ~n24135;
  assign n24139 = n24138 & n24137;
  assign n24257 = ~n24140 | ~n24139;
  assign n24141 = ~n24251 | ~n24257;
  assign P1_U3462 = ~n24142 | ~n24141;
  assign n24153 = ~P1_REG0_REG_2__SCAN_IN | ~n24240;
  assign n24146 = ~n24143 & ~n24201;
  assign n24145 = ~n24144 & ~n24241;
  assign n24151 = ~n24146 & ~n24145;
  assign n24148 = ~n24147 & ~n24220;
  assign n24150 = ~n24149 & ~n24148;
  assign n24260 = ~n24151 | ~n24150;
  assign n24152 = ~n24251 | ~n24260;
  assign P1_U3465 = ~n24153 | ~n24152;
  assign n24164 = ~P1_REG0_REG_3__SCAN_IN | ~n24240;
  assign n24157 = ~n24154 & ~n24201;
  assign n24156 = ~n24155 & ~n24241;
  assign n24162 = ~n24157 & ~n24156;
  assign n24159 = ~n24158 & ~n24220;
  assign n24161 = ~n24160 & ~n24159;
  assign n24263 = ~n24162 | ~n24161;
  assign n24163 = ~n24251 | ~n24263;
  assign P1_U3468 = ~n24164 | ~n24163;
  assign n24176 = ~P1_REG0_REG_4__SCAN_IN | ~n24240;
  assign n24166 = ~n24241 & ~n24165;
  assign n24168 = n24167 | n24166;
  assign n24172 = ~n24169 & ~n24168;
  assign n24171 = ~n24170 | ~n24247;
  assign n24173 = ~n24172 | ~n24171;
  assign n24266 = n24174 | n24173;
  assign n24175 = ~n24251 | ~n24266;
  assign P1_U3471 = ~n24176 | ~n24175;
  assign n24188 = ~P1_REG0_REG_5__SCAN_IN | ~n24240;
  assign n24180 = ~n24177 | ~n24216;
  assign n24179 = ~n24230 | ~n14266;
  assign n24181 = ~n24180 | ~n24179;
  assign n24186 = ~n24182 & ~n24181;
  assign n24184 = ~n24183;
  assign n24185 = ~n24184 | ~n24228;
  assign n24269 = ~n24186 | ~n24185;
  assign n24187 = ~n24251 | ~n24269;
  assign P1_U3474 = ~n24188 | ~n24187;
  assign n24200 = ~P1_REG0_REG_6__SCAN_IN | ~n24240;
  assign n24192 = ~n24189 | ~n24216;
  assign n24191 = ~n24190 | ~n24230;
  assign n24193 = ~n24192 | ~n24191;
  assign n24198 = ~n24194 & ~n24193;
  assign n24196 = ~n24195;
  assign n24197 = ~n24196 | ~n24228;
  assign n24272 = ~n24198 | ~n24197;
  assign n24199 = ~n24251 | ~n24272;
  assign P1_U3477 = ~n24200 | ~n24199;
  assign n24212 = ~P1_REG0_REG_7__SCAN_IN | ~n24240;
  assign n24205 = ~n24202 & ~n24201;
  assign n24204 = ~n24203 & ~n24241;
  assign n24210 = ~n24205 & ~n24204;
  assign n24207 = ~n24206 & ~n24220;
  assign n24209 = ~n24208 & ~n24207;
  assign n24275 = ~n24210 | ~n24209;
  assign n24211 = ~n24251 | ~n24275;
  assign P1_U3480 = ~n24212 | ~n24211;
  assign n24227 = ~P1_REG0_REG_8__SCAN_IN | ~n24240;
  assign n24215 = ~n24213 | ~n24230;
  assign n24219 = n24215 & n24214;
  assign n24218 = ~n24217 | ~n24216;
  assign n24223 = ~n24219 | ~n24218;
  assign n24222 = ~n24221 & ~n24220;
  assign n24224 = ~n24223 & ~n24222;
  assign n24278 = ~n24225 | ~n24224;
  assign n24226 = ~n24251 | ~n24278;
  assign P1_U3483 = ~n24227 | ~n24226;
  assign n24239 = ~P1_REG0_REG_9__SCAN_IN | ~n24240;
  assign n24233 = ~n24229 | ~n24228;
  assign n24232 = ~n24231 | ~n24230;
  assign n24234 = ~n24233 | ~n24232;
  assign n24236 = ~n24235 & ~n24234;
  assign n24281 = ~n24237 | ~n24236;
  assign n24238 = ~n24251 | ~n24281;
  assign P1_U3486 = ~n24239 | ~n24238;
  assign n24253 = ~P1_REG0_REG_10__SCAN_IN | ~n24240;
  assign n24243 = ~n24242 & ~n24241;
  assign n24245 = n24244 | n24243;
  assign n24250 = ~n24246 & ~n24245;
  assign n24249 = ~n24248 | ~n24247;
  assign n24285 = ~n24250 | ~n24249;
  assign n24252 = ~n24251 | ~n24285;
  assign P1_U3489 = ~n24253 | ~n24252;
  assign n24256 = ~P1_REG1_REG_0__SCAN_IN | ~n24284;
  assign n24255 = ~n24286 | ~n24254;
  assign P1_U3528 = ~n24256 | ~n24255;
  assign n24259 = ~P1_REG1_REG_1__SCAN_IN | ~n24284;
  assign n24258 = ~n24286 | ~n24257;
  assign P1_U3529 = ~n24259 | ~n24258;
  assign n24262 = ~P1_REG1_REG_2__SCAN_IN | ~n24284;
  assign n24261 = ~n24286 | ~n24260;
  assign P1_U3530 = ~n24262 | ~n24261;
  assign n24265 = ~P1_REG1_REG_3__SCAN_IN | ~n24284;
  assign n24264 = ~n24286 | ~n24263;
  assign P1_U3531 = ~n24265 | ~n24264;
  assign n24268 = ~P1_REG1_REG_4__SCAN_IN | ~n24284;
  assign n24267 = ~n24286 | ~n24266;
  assign P1_U3532 = ~n24268 | ~n24267;
  assign n24271 = ~P1_REG1_REG_5__SCAN_IN | ~n24284;
  assign n24270 = ~n24286 | ~n24269;
  assign P1_U3533 = ~n24271 | ~n24270;
  assign n24274 = ~P1_REG1_REG_6__SCAN_IN | ~n24284;
  assign n24273 = ~n24286 | ~n24272;
  assign P1_U3534 = ~n24274 | ~n24273;
  assign n24277 = ~P1_REG1_REG_7__SCAN_IN | ~n24284;
  assign n24276 = ~n24286 | ~n24275;
  assign P1_U3535 = ~n24277 | ~n24276;
  assign n24280 = ~P1_REG1_REG_8__SCAN_IN | ~n24284;
  assign n24279 = ~n24286 | ~n24278;
  assign P1_U3536 = ~n24280 | ~n24279;
  assign n24283 = ~P1_REG1_REG_9__SCAN_IN | ~n24284;
  assign n24282 = ~n24286 | ~n24281;
  assign P1_U3537 = ~n24283 | ~n24282;
  assign n24288 = ~P1_REG1_REG_10__SCAN_IN | ~n24284;
  assign n24287 = ~n24286 | ~n24285;
  assign P1_U3538 = ~n24288 | ~n24287;
  assign n24291 = ~n24319 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n24290 = ~n24289 | ~P1_U4016;
  assign P1_U3578 = ~n24291 | ~n24290;
  assign n24294 = ~n24319 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n24293 = ~n24292 | ~n24307;
  assign P1_U3579 = ~n24294 | ~n24293;
  assign n24297 = ~n24319 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n24296 = ~n24295 | ~n24307;
  assign P1_U3580 = ~n24297 | ~n24296;
  assign n24300 = ~n24319 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n24299 = ~P1_U4016 | ~n24298;
  assign P1_U3581 = ~n24300 | ~n24299;
  assign n24303 = ~n24319 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n24302 = ~n24301 | ~n24307;
  assign P1_U3582 = ~n24303 | ~n24302;
  assign n24306 = ~n24319 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n24305 = ~n24304 | ~n24307;
  assign P1_U3583 = ~n24306 | ~n24305;
  assign n24310 = ~n24319 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n24309 = ~n24308 | ~n24307;
  assign P1_U3584 = ~n24310 | ~n24309;
  assign n24313 = ~n24319 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n24312 = ~n24311 | ~P1_U4016;
  assign P1_U3585 = ~n24313 | ~n24312;
  assign n24315 = ~n24319 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n24314 = ~n14111 | ~P1_U4016;
  assign P1_U3586 = ~n24315 | ~n24314;
  assign n24318 = ~n24319 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n24317 = ~P1_U4016 | ~n24316;
  assign P1_U3587 = ~n24318 | ~n24317;
  assign n24322 = ~n24319 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n24321 = ~P1_U4016 | ~n24320;
  assign P1_U3588 = ~n24322 | ~n24321;
  assign n24326 = ~n24319 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n24325 = ~P1_U4016 | ~n24323;
  assign P1_U3589 = ~n24326 | ~n24325;
  assign n24329 = ~n24319 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n24328 = ~P1_U4016 | ~n24327;
  assign P1_U3590 = ~n24329 | ~n24328;
  assign n24332 = ~n24319 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n24331 = ~P1_U4016 | ~n24330;
  assign P1_U3591 = ~n24332 | ~n24331;
  assign n24335 = ~n24334 | ~n24333;
  assign n24913 = ~P2_U3088 & ~n24521;
  assign P2_U3087 = ~n24913 & ~P2_U3947;
  assign n24337 = ~n24455 | ~n25049;
  assign n24657 = ~P2_REG3_REG_7__SCAN_IN | ~P2_U3088;
  assign n24339 = ~n24337 | ~n24657;
  assign n24338 = ~n24484 & ~n13779;
  assign n24348 = ~n24339 & ~n24338;
  assign n24342 = n24340 ^ n24341;
  assign n24344 = ~n24342 | ~n24506;
  assign n24343 = ~n24508 | ~n25454;
  assign n24346 = ~n24344 | ~n24343;
  assign n24345 = ~n24511 & ~n25059;
  assign n24347 = ~n24346 & ~n24345;
  assign P2_U3185 = ~n24348 | ~n24347;
  assign n24352 = ~n24499 & ~n24349;
  assign n24350 = ~n24500 | ~n25021;
  assign n24717 = ~P2_REG3_REG_10__SCAN_IN | ~P2_U3088;
  assign n24351 = ~n24350 | ~n24717;
  assign n24361 = ~n24352 & ~n24351;
  assign n24355 = n24354 ^ ~n24353;
  assign n24359 = ~n24355 & ~n24471;
  assign n24357 = ~n24508 | ~n25489;
  assign n24356 = ~n24475 | ~n24964;
  assign n24358 = ~n24357 | ~n24356;
  assign n24360 = ~n24359 & ~n24358;
  assign P2_U3189 = ~n24361 | ~n24360;
  assign n24364 = ~n24499 & ~n14079;
  assign n24362 = ~n24500 | ~n25252;
  assign n24575 = ~P2_REG3_REG_3__SCAN_IN | ~P2_U3088;
  assign n24363 = ~n24362 | ~n24575;
  assign n24373 = ~n24364 & ~n24363;
  assign n24369 = ~n24508 | ~n25410;
  assign n24367 = n24365 ^ n24366;
  assign n24368 = ~n24506 | ~n24367;
  assign n24371 = ~n24369 | ~n24368;
  assign n24370 = ~P2_REG3_REG_3__SCAN_IN & ~n24511;
  assign n24372 = ~n24371 & ~n24370;
  assign P2_U3190 = ~n24373 | ~n24372;
  assign n24374 = ~n24455 | ~n25021;
  assign n24682 = ~P2_REG3_REG_8__SCAN_IN | ~P2_U3088;
  assign n24376 = ~n24374 | ~n24682;
  assign n24375 = ~n24484 & ~n25093;
  assign n24388 = ~n24376 & ~n24375;
  assign n24380 = ~n24378;
  assign n24381 = ~n24380 | ~n24379;
  assign n24382 = n24377 ^ ~n24381;
  assign n24384 = ~n24382 | ~n24506;
  assign n24383 = ~n24508 | ~n25467;
  assign n24386 = ~n24384 | ~n24383;
  assign n24385 = ~n24511 & ~n25033;
  assign n24387 = ~n24386 & ~n24385;
  assign P2_U3193 = ~n24388 | ~n24387;
  assign n24391 = ~n24499 & ~n24389;
  assign n24774 = ~P2_STATE_REG_SCAN_IN & ~n24390;
  assign n24393 = ~n24391 & ~n24774;
  assign n24392 = ~n24500 | ~n24976;
  assign n24399 = ~n24393 | ~n24392;
  assign n24397 = ~n24508 | ~n24394;
  assign n24396 = ~n24475 | ~n24395;
  assign n24398 = ~n24397 | ~n24396;
  assign n24406 = ~n24399 & ~n24398;
  assign n24403 = ~n24402 | ~n24401;
  assign n24404 = n24400 ^ ~n24403;
  assign n24405 = ~n24404 | ~n24506;
  assign P2_U3196 = ~n24406 | ~n24405;
  assign n24409 = ~n24499 & ~n13779;
  assign n24407 = ~n24500 | ~n25183;
  assign n24622 = ~P2_REG3_REG_5__SCAN_IN | ~P2_U3088;
  assign n24408 = ~n24407 | ~n24622;
  assign n24418 = ~n24409 & ~n24408;
  assign n24412 = n24410 ^ n24411;
  assign n24416 = ~n24412 & ~n24471;
  assign n24414 = ~n24508 | ~n25432;
  assign n24413 = ~n24475 | ~n25106;
  assign n24415 = ~n24414 | ~n24413;
  assign n24417 = ~n24416 & ~n24415;
  assign P2_U3199 = ~n24418 | ~n24417;
  assign n25080 = ~n25150;
  assign n24421 = ~n24499 & ~n25080;
  assign n24419 = ~n24500 | ~n25214;
  assign n24596 = ~P2_REG3_REG_4__SCAN_IN | ~P2_U3088;
  assign n24420 = ~n24419 | ~n24596;
  assign n24433 = ~n24421 & ~n24420;
  assign n24428 = ~n24508 | ~n25420;
  assign n24425 = ~n24423 | ~n24422;
  assign n24426 = n24425 ^ n24424;
  assign n24427 = ~n24506 | ~n24426;
  assign n24431 = ~n24428 | ~n24427;
  assign n24430 = ~n24511 & ~n24429;
  assign n24432 = ~n24431 & ~n24430;
  assign P2_U3202 = ~n24433 | ~n24432;
  assign n24437 = ~n24499 & ~n24434;
  assign n24435 = ~n24500 | ~n25049;
  assign n24697 = ~P2_REG3_REG_9__SCAN_IN | ~P2_U3088;
  assign n24436 = ~n24435 | ~n24697;
  assign n24448 = ~n24437 & ~n24436;
  assign n24441 = n24439 | n24438;
  assign n24442 = ~n24441 | ~n24440;
  assign n24444 = ~n24442 | ~n24506;
  assign n24443 = ~n24508 | ~n25479;
  assign n24446 = ~n24444 | ~n24443;
  assign n24445 = ~n24511 & ~n25009;
  assign n24447 = ~n24446 & ~n24445;
  assign P2_U3203 = ~n24448 | ~n24447;
  assign n24450 = ~n25254 | ~n24449;
  assign n24451 = ~n24450 | ~n14816;
  assign n24453 = n24452 & n24451;
  assign n24461 = ~n24506 | ~n24453;
  assign n24457 = ~n24508 | ~n24454;
  assign n24456 = ~n24455 | ~n25274;
  assign n24459 = ~n24457 | ~n24456;
  assign n25266 = ~P2_REG3_REG_0__SCAN_IN;
  assign n24458 = ~n24487 & ~n25266;
  assign n24460 = ~n24459 & ~n24458;
  assign P2_U3204 = ~n24461 | ~n24460;
  assign n24465 = ~n24499 & ~n24462;
  assign n24463 = ~n24500 | ~n24955;
  assign n24784 = ~P2_REG3_REG_13__SCAN_IN | ~P2_U3088;
  assign n24464 = ~n24463 | ~n24784;
  assign n24481 = ~n24465 & ~n24464;
  assign n24468 = ~n24466;
  assign n24469 = ~n24468 & ~n24467;
  assign n24472 = n24470 ^ ~n24469;
  assign n24479 = ~n24472 & ~n24471;
  assign n24477 = ~n24508 | ~n24473;
  assign n24476 = ~n24475 | ~n24474;
  assign n24478 = ~n24477 | ~n24476;
  assign n24480 = ~n24479 & ~n24478;
  assign P2_U3206 = ~n24481 | ~n24480;
  assign n24486 = ~n24499 & ~n24482;
  assign n24483 = ~n25274;
  assign n24485 = ~n24484 & ~n24483;
  assign n24498 = ~n24486 & ~n24485;
  assign n24496 = ~n24487 & ~n16613;
  assign n24494 = ~n24508 | ~n25399;
  assign n24490 = n24489 | n24488;
  assign n24492 = ~n24491 | ~n24490;
  assign n24493 = ~n24506 | ~n24492;
  assign n24495 = ~n24494 | ~n24493;
  assign n24497 = ~n24496 & ~n24495;
  assign P2_U3209 = ~n24498 | ~n24497;
  assign n24503 = ~n24499 & ~n25093;
  assign n24501 = ~n24500 | ~n25150;
  assign n24637 = ~P2_REG3_REG_6__SCAN_IN | ~P2_U3088;
  assign n24502 = ~n24501 | ~n24637;
  assign n24515 = ~n24503 & ~n24502;
  assign n24507 = n24504 ^ n24505;
  assign n24510 = ~n24507 | ~n24506;
  assign n24509 = ~n24508 | ~n25090;
  assign n24513 = ~n24510 | ~n24509;
  assign n24512 = ~n24511 & ~n25073;
  assign n24514 = ~n24513 & ~n24512;
  assign P2_U3211 = ~n24515 | ~n24514;
  assign n24896 = ~n24521 | ~n17049;
  assign n24517 = ~n24519 & ~n24516;
  assign n24933 = ~n24521 | ~n24517;
  assign n24523 = ~n24933 & ~P2_REG2_REG_0__SCAN_IN;
  assign n24520 = ~n24519 & ~n24518;
  assign n24925 = ~n24521 | ~n24520;
  assign n24522 = ~n24925 & ~P2_REG1_REG_0__SCAN_IN;
  assign n24524 = ~n24523 & ~n24522;
  assign n24525 = ~n24916 | ~n24524;
  assign n24533 = ~n24525 | ~P2_IR_REG_0__SCAN_IN;
  assign n25283 = ~P2_REG2_REG_0__SCAN_IN;
  assign n24535 = ~n24933 & ~n25283;
  assign n24526 = ~P2_REG1_REG_0__SCAN_IN;
  assign n24545 = ~n24925 & ~n24526;
  assign n24527 = ~n24535 & ~n24545;
  assign n24531 = ~P2_IR_REG_0__SCAN_IN & ~n24527;
  assign n24529 = ~n24913 | ~P2_ADDR_REG_0__SCAN_IN;
  assign n24528 = ~P2_REG3_REG_0__SCAN_IN | ~P2_U3088;
  assign n24530 = ~n24529 | ~n24528;
  assign n24532 = ~n24531 & ~n24530;
  assign P2_U3214 = ~n24533 | ~n24532;
  assign n24559 = P2_REG2_REG_1__SCAN_IN ^ n24565;
  assign n24534 = ~n24559 & ~n14091;
  assign n24539 = ~n24535 | ~n24534;
  assign n24744 = ~n24933;
  assign n24536 = ~n24559;
  assign n24558 = P2_IR_REG_0__SCAN_IN & P2_REG2_REG_0__SCAN_IN;
  assign n24537 = ~n24536 & ~n24558;
  assign n24538 = ~n24744 | ~n24537;
  assign n24543 = ~n24539 | ~n24538;
  assign n24541 = ~n24913 | ~P2_ADDR_REG_1__SCAN_IN;
  assign n24540 = ~P2_REG3_REG_1__SCAN_IN | ~P2_U3088;
  assign n24542 = ~n24541 | ~n24540;
  assign n24553 = ~n24543 & ~n24542;
  assign n24564 = P2_REG1_REG_1__SCAN_IN ^ n24565;
  assign n24544 = ~n24564 & ~n14091;
  assign n24549 = ~n24545 | ~n24544;
  assign n24771 = ~n24925;
  assign n24546 = ~n24564;
  assign n24563 = P2_IR_REG_0__SCAN_IN & P2_REG1_REG_0__SCAN_IN;
  assign n24547 = ~n24546 & ~n24563;
  assign n24548 = ~n24771 | ~n24547;
  assign n24551 = ~n24549 | ~n24548;
  assign n24550 = ~n24916 & ~n14424;
  assign n24552 = ~n24551 & ~n24550;
  assign P2_U3215 = ~n24553 | ~n24552;
  assign n24555 = ~n24913 | ~P2_ADDR_REG_2__SCAN_IN;
  assign n24554 = ~P2_REG3_REG_2__SCAN_IN | ~P2_U3088;
  assign n24557 = ~n24555 | ~n24554;
  assign n24556 = ~n24916 & ~n13793;
  assign n24573 = ~n24557 & ~n24556;
  assign n24561 = ~n24559 | ~n24558;
  assign n24560 = ~n24565 | ~P2_REG2_REG_1__SCAN_IN;
  assign n24579 = ~n24561 | ~n24560;
  assign n24580 = P2_REG2_REG_2__SCAN_IN ^ n24586;
  assign n24562 = n24579 ^ ~n24580;
  assign n24571 = ~n24933 & ~n24562;
  assign n24567 = ~n24564 | ~n24563;
  assign n24566 = ~n24565 | ~P2_REG1_REG_1__SCAN_IN;
  assign n24585 = ~n24567 | ~n24566;
  assign n24568 = ~P2_REG1_REG_2__SCAN_IN;
  assign n24584 = n24586 ^ ~n24568;
  assign n24569 = n24585 ^ ~n24584;
  assign n24570 = ~n24925 & ~n24569;
  assign n24572 = ~n24571 & ~n24570;
  assign P2_U3216 = ~n24573 | ~n24572;
  assign n24574 = ~P2_ADDR_REG_3__SCAN_IN | ~n24913;
  assign n24578 = ~n24575 | ~n24574;
  assign n24577 = ~n24916 & ~n24576;
  assign n24594 = ~n24578 & ~n24577;
  assign n24582 = ~n24580 | ~n24579;
  assign n24581 = ~n24586 | ~P2_REG2_REG_2__SCAN_IN;
  assign n24600 = ~n24582 | ~n24581;
  assign n24599 = P2_REG2_REG_3__SCAN_IN ^ n24606;
  assign n24583 = n24600 ^ ~n24599;
  assign n24592 = ~n24933 & ~n24583;
  assign n24588 = ~n24585 | ~n24584;
  assign n24587 = ~n24586 | ~P2_REG1_REG_2__SCAN_IN;
  assign n24605 = ~n24588 | ~n24587;
  assign n24589 = ~P2_REG1_REG_3__SCAN_IN;
  assign n24604 = n24606 ^ ~n24589;
  assign n24590 = n24605 ^ ~n24604;
  assign n24591 = ~n24925 & ~n24590;
  assign n24593 = ~n24592 & ~n24591;
  assign P2_U3217 = ~n24594 | ~n24593;
  assign n24595 = ~P2_ADDR_REG_4__SCAN_IN | ~n24913;
  assign n24598 = ~n24596 | ~n24595;
  assign n25355 = ~n24627;
  assign n24597 = ~n24916 & ~n25355;
  assign n24614 = ~n24598 & ~n24597;
  assign n24602 = ~n24600 | ~n24599;
  assign n24601 = ~n24606 | ~P2_REG2_REG_3__SCAN_IN;
  assign n24626 = ~n24602 | ~n24601;
  assign n24625 = P2_REG2_REG_4__SCAN_IN ^ n24627;
  assign n24603 = n24626 ^ ~n24625;
  assign n24612 = ~n24933 & ~n24603;
  assign n24608 = ~n24605 | ~n24604;
  assign n24607 = ~n24606 | ~P2_REG1_REG_3__SCAN_IN;
  assign n24616 = ~n24608 | ~n24607;
  assign n24609 = ~P2_REG1_REG_4__SCAN_IN;
  assign n24615 = n24627 ^ ~n24609;
  assign n24610 = n24616 ^ ~n24615;
  assign n24611 = ~n24925 & ~n24610;
  assign n24613 = ~n24612 & ~n24611;
  assign P2_U3218 = ~n24614 | ~n24613;
  assign n24618 = ~n24616 | ~n24615;
  assign n24617 = ~n24627 | ~P2_REG1_REG_4__SCAN_IN;
  assign n24646 = ~n24618 | ~n24617;
  assign n24619 = ~P2_REG1_REG_5__SCAN_IN;
  assign n24645 = n24647 ^ ~n24619;
  assign n24620 = n24646 ^ ~n24645;
  assign n24624 = ~n24925 & ~n24620;
  assign n24621 = ~P2_ADDR_REG_5__SCAN_IN | ~n24913;
  assign n24623 = ~n24622 | ~n24621;
  assign n24635 = ~n24624 & ~n24623;
  assign n24629 = ~n24626 | ~n24625;
  assign n24628 = ~n24627 | ~P2_REG2_REG_4__SCAN_IN;
  assign n24641 = ~n24629 | ~n24628;
  assign n24640 = P2_REG2_REG_5__SCAN_IN ^ n24647;
  assign n24630 = n24641 ^ ~n24640;
  assign n24633 = ~n24933 & ~n24630;
  assign n24632 = ~n24916 & ~n24631;
  assign n24634 = ~n24633 & ~n24632;
  assign P2_U3219 = ~n24635 | ~n24634;
  assign n24636 = ~P2_ADDR_REG_6__SCAN_IN | ~n24913;
  assign n24639 = ~n24637 | ~n24636;
  assign n25349 = ~n24668;
  assign n24638 = ~n24916 & ~n25349;
  assign n24655 = ~n24639 & ~n24638;
  assign n24643 = ~n24641 | ~n24640;
  assign n24642 = ~n24647 | ~P2_REG2_REG_5__SCAN_IN;
  assign n24667 = ~n24643 | ~n24642;
  assign n24666 = P2_REG2_REG_6__SCAN_IN ^ n24668;
  assign n24644 = n24667 ^ ~n24666;
  assign n24653 = ~n24933 & ~n24644;
  assign n24649 = ~n24646 | ~n24645;
  assign n24648 = ~n24647 | ~P2_REG1_REG_5__SCAN_IN;
  assign n24661 = ~n24649 | ~n24648;
  assign n24650 = ~P2_REG1_REG_6__SCAN_IN;
  assign n24660 = n24668 ^ ~n24650;
  assign n24651 = n24661 ^ ~n24660;
  assign n24652 = ~n24925 & ~n24651;
  assign n24654 = ~n24653 & ~n24652;
  assign P2_U3220 = ~n24655 | ~n24654;
  assign n24656 = ~P2_ADDR_REG_7__SCAN_IN | ~n24913;
  assign n24659 = ~n24657 | ~n24656;
  assign n25343 = ~n24687;
  assign n24658 = ~n24916 & ~n25343;
  assign n24675 = ~n24659 & ~n24658;
  assign n24663 = ~n24661 | ~n24660;
  assign n24662 = ~n24668 | ~P2_REG1_REG_6__SCAN_IN;
  assign n24686 = ~n24663 | ~n24662;
  assign n24664 = ~P2_REG1_REG_7__SCAN_IN;
  assign n24685 = n24687 ^ ~n24664;
  assign n24665 = n24686 ^ ~n24685;
  assign n24673 = ~n24925 & ~n24665;
  assign n24670 = ~n24667 | ~n24666;
  assign n24669 = ~n24668 | ~P2_REG2_REG_6__SCAN_IN;
  assign n24677 = ~n24670 | ~n24669;
  assign n24676 = P2_REG2_REG_7__SCAN_IN ^ n24687;
  assign n24671 = n24677 ^ ~n24676;
  assign n24672 = ~n24933 & ~n24671;
  assign n24674 = ~n24673 & ~n24672;
  assign P2_U3221 = ~n24675 | ~n24674;
  assign n24679 = ~n24677 | ~n24676;
  assign n24678 = ~n24687 | ~P2_REG2_REG_7__SCAN_IN;
  assign n24698 = ~n24679 | ~n24678;
  assign n24699 = P2_REG2_REG_8__SCAN_IN ^ n24707;
  assign n24680 = n24698 ^ ~n24699;
  assign n24684 = ~n24933 & ~n24680;
  assign n24681 = ~P2_ADDR_REG_8__SCAN_IN | ~n24913;
  assign n24683 = ~n24682 | ~n24681;
  assign n24695 = ~n24684 & ~n24683;
  assign n24689 = ~n24686 | ~n24685;
  assign n24688 = ~n24687 | ~P2_REG1_REG_7__SCAN_IN;
  assign n24708 = ~n24689 | ~n24688;
  assign n24690 = ~P2_REG1_REG_8__SCAN_IN;
  assign n24709 = n24707 ^ ~n24690;
  assign n24691 = n24708 ^ ~n24709;
  assign n24693 = ~n24925 & ~n24691;
  assign n25340 = ~n24707 | ~P2_STATE_REG_SCAN_IN;
  assign n24692 = ~n24896 & ~n25340;
  assign n24694 = ~n24693 & ~n24692;
  assign P2_U3222 = ~n24695 | ~n24694;
  assign n24712 = ~n24725;
  assign n25331 = ~n24712 & ~P2_U3088;
  assign n24696 = ~n24875 | ~n25331;
  assign n24706 = ~n24697 | ~n24696;
  assign n24704 = ~P2_ADDR_REG_9__SCAN_IN | ~n24913;
  assign n24701 = ~n24707 | ~P2_REG2_REG_8__SCAN_IN;
  assign n24700 = ~n24699 | ~n24698;
  assign n24727 = ~n24701 | ~n24700;
  assign n24726 = P2_REG2_REG_9__SCAN_IN ^ n24712;
  assign n24702 = n24727 ^ ~n24726;
  assign n24703 = ~n24702 | ~n24744;
  assign n24705 = ~n24704 | ~n24703;
  assign n24715 = ~n24706 & ~n24705;
  assign n24711 = ~n24707 | ~P2_REG1_REG_8__SCAN_IN;
  assign n24710 = ~n24709 | ~n24708;
  assign n24720 = ~n24711 | ~n24710;
  assign n24719 = P2_REG1_REG_9__SCAN_IN ^ n24712;
  assign n24713 = n24720 ^ ~n24719;
  assign n24714 = ~n24713 | ~n24771;
  assign P2_U3223 = ~n24715 | ~n24714;
  assign n24716 = ~P2_ADDR_REG_10__SCAN_IN | ~n24913;
  assign n24734 = ~n24717 | ~n24716;
  assign n24718 = ~P2_REG1_REG_10__SCAN_IN;
  assign n24753 = n24751 ^ ~n24718;
  assign n24722 = ~P2_REG1_REG_9__SCAN_IN & ~n24725;
  assign n24721 = ~n24720 & ~n24719;
  assign n24752 = ~n24722 & ~n24721;
  assign n24723 = n24753 ^ n24752;
  assign n24732 = ~n24723 | ~n24771;
  assign n24724 = ~P2_REG2_REG_10__SCAN_IN;
  assign n24740 = n24751 ^ ~n24724;
  assign n24729 = ~P2_REG2_REG_9__SCAN_IN & ~n24725;
  assign n24728 = ~n24727 & ~n24726;
  assign n24730 = n24740 ^ n24741;
  assign n24731 = ~n24730 | ~n24744;
  assign n24733 = ~n24732 | ~n24731;
  assign n24737 = ~n24734 & ~n24733;
  assign n24735 = ~n24751;
  assign n25326 = ~n24735 & ~P2_U3088;
  assign n24736 = ~n24875 | ~n25326;
  assign P2_U3224 = ~n24737 | ~n24736;
  assign n24750 = ~n24765;
  assign n25321 = ~n24750 & ~P2_U3088;
  assign n24738 = ~n24875 | ~n25321;
  assign n24749 = ~n24739 | ~n24738;
  assign n24761 = P2_REG2_REG_11__SCAN_IN ^ n24750;
  assign n24743 = ~n24751 | ~P2_REG2_REG_10__SCAN_IN;
  assign n24742 = ~n24741 | ~n24740;
  assign n24760 = ~n24743 | ~n24742;
  assign n24745 = n24761 ^ ~n24760;
  assign n24747 = ~n24745 | ~n24744;
  assign n24746 = ~P2_ADDR_REG_11__SCAN_IN | ~n24913;
  assign n24748 = ~n24747 | ~n24746;
  assign n24758 = ~n24749 & ~n24748;
  assign n24767 = P2_REG1_REG_11__SCAN_IN ^ ~n24750;
  assign n24755 = ~n24751 | ~P2_REG1_REG_10__SCAN_IN;
  assign n24754 = ~n24753 | ~n24752;
  assign n24766 = ~n24755 | ~n24754;
  assign n24756 = n24767 ^ n24766;
  assign n24757 = ~n24756 | ~n24771;
  assign P2_U3225 = ~n24758 | ~n24757;
  assign n24794 = n24779 | P2_REG2_REG_12__SCAN_IN;
  assign n24759 = ~n24779 | ~P2_REG2_REG_12__SCAN_IN;
  assign n24795 = ~n24794 | ~n24759;
  assign n24763 = ~P2_REG2_REG_11__SCAN_IN & ~n24765;
  assign n24762 = ~n24761 & ~n24760;
  assign n24764 = n24795 ^ n24796;
  assign n24778 = ~n24764 & ~n24933;
  assign n24769 = ~P2_REG1_REG_11__SCAN_IN | ~n24765;
  assign n24768 = ~n24767 | ~n24766;
  assign n24787 = ~n24769 | ~n24768;
  assign n24785 = n24779 | P2_REG1_REG_12__SCAN_IN;
  assign n24770 = ~n24779 | ~P2_REG1_REG_12__SCAN_IN;
  assign n24786 = ~n24785 | ~n24770;
  assign n24772 = n24787 ^ ~n24786;
  assign n24776 = ~n24772 | ~n24771;
  assign n24773 = P2_ADDR_REG_12__SCAN_IN & n24913;
  assign n24775 = ~n24774 & ~n24773;
  assign n24777 = ~n24776 | ~n24775;
  assign n24782 = ~n24778 & ~n24777;
  assign n24780 = ~n24779;
  assign n25316 = ~n24780 & ~P2_U3088;
  assign n24781 = ~n24875 | ~n25316;
  assign P2_U3226 = ~n24782 | ~n24781;
  assign n24783 = ~P2_ADDR_REG_13__SCAN_IN | ~n24913;
  assign n24806 = ~n24784 | ~n24783;
  assign n24792 = P2_REG1_REG_13__SCAN_IN ^ n24817;
  assign n24789 = ~n24785;
  assign n24788 = ~n24787 & ~n24786;
  assign n24791 = ~n24789 & ~n24788;
  assign n24790 = ~n24792 & ~n24791;
  assign n24793 = ~n24790 & ~n24925;
  assign n24818 = ~n24792 | ~n24791;
  assign n24804 = ~n24793 | ~n24818;
  assign n24798 = ~n24794;
  assign n24797 = ~n24796 & ~n24795;
  assign n24801 = ~n24798 & ~n24797;
  assign n24800 = P2_REG2_REG_13__SCAN_IN ^ n24817;
  assign n24799 = ~n24801 & ~n24800;
  assign n24802 = ~n24799 & ~n24933;
  assign n24812 = ~n24801 | ~n24800;
  assign n24803 = ~n24802 | ~n24812;
  assign n24805 = ~n24804 | ~n24803;
  assign n24809 = ~n24806 & ~n24805;
  assign n24807 = ~n24817;
  assign n25312 = ~n24807 & ~P2_U3088;
  assign n24808 = ~n24875 | ~n25312;
  assign P2_U3227 = ~n24809 | ~n24808;
  assign n24810 = P2_ADDR_REG_14__SCAN_IN & n24913;
  assign n24829 = ~n24811 & ~n24810;
  assign n24813 = ~P2_REG2_REG_13__SCAN_IN | ~n24817;
  assign n24838 = ~n24813 | ~n24812;
  assign n24841 = ~P2_REG2_REG_14__SCAN_IN | ~n24832;
  assign n24839 = P2_REG2_REG_14__SCAN_IN | n24832;
  assign n24814 = ~n24841 | ~n24839;
  assign n24815 = n24838 ^ n24814;
  assign n24827 = ~n24815 & ~n24933;
  assign n24816 = ~n24832;
  assign n25307 = ~n24816 & ~P2_U3088;
  assign n24825 = ~n24875 | ~n25307;
  assign n24822 = P2_REG1_REG_14__SCAN_IN ^ n24832;
  assign n24819 = ~P2_REG1_REG_13__SCAN_IN | ~n24817;
  assign n24821 = ~n24819 | ~n24818;
  assign n24820 = ~n24822 & ~n24821;
  assign n24823 = ~n24820 & ~n24925;
  assign n24833 = ~n24822 | ~n24821;
  assign n24824 = ~n24823 | ~n24833;
  assign n24826 = ~n24825 | ~n24824;
  assign n24828 = ~n24827 & ~n24826;
  assign P2_U3228 = ~n24829 | ~n24828;
  assign n24830 = ~P2_ADDR_REG_15__SCAN_IN | ~n24913;
  assign n24849 = ~n24831 | ~n24830;
  assign n24834 = ~P2_REG1_REG_14__SCAN_IN | ~n24832;
  assign n24855 = ~n24834 | ~n24833;
  assign n24836 = n24842 ^ ~n24855;
  assign n24835 = ~P2_REG1_REG_15__SCAN_IN & ~n24836;
  assign n24837 = ~n24835 & ~n24925;
  assign n24856 = ~P2_REG1_REG_15__SCAN_IN | ~n24836;
  assign n24847 = ~n24837 | ~n24856;
  assign n24840 = ~n24839 | ~n24838;
  assign n24862 = ~n24841 | ~n24840;
  assign n24844 = n24842 ^ ~n24862;
  assign n24843 = ~P2_REG2_REG_15__SCAN_IN & ~n24844;
  assign n24845 = ~n24843 & ~n24933;
  assign n24864 = ~P2_REG2_REG_15__SCAN_IN | ~n24844;
  assign n24846 = ~n24845 | ~n24864;
  assign n24848 = ~n24847 | ~n24846;
  assign n24852 = ~n24849 & ~n24848;
  assign n24850 = ~n24916;
  assign n24851 = ~n24850 | ~n24863;
  assign P2_U3229 = ~n24852 | ~n24851;
  assign n24853 = ~P2_ADDR_REG_16__SCAN_IN | ~n24913;
  assign n24873 = ~n24854 | ~n24853;
  assign n24874 = ~n24886;
  assign n24860 = P2_REG1_REG_16__SCAN_IN ^ ~n24874;
  assign n24857 = ~n24863 | ~n24855;
  assign n24859 = ~n24857 | ~n24856;
  assign n24858 = ~n24860 & ~n24859;
  assign n24861 = ~n24858 & ~n24925;
  assign n24882 = ~n24860 | ~n24859;
  assign n24871 = ~n24861 | ~n24882;
  assign n24868 = P2_REG2_REG_16__SCAN_IN ^ ~n24874;
  assign n24865 = ~n24863 | ~n24862;
  assign n24867 = ~n24865 | ~n24864;
  assign n24866 = ~n24868 & ~n24867;
  assign n24869 = ~n24866 & ~n24933;
  assign n24887 = ~n24868 | ~n24867;
  assign n24870 = ~n24869 | ~n24887;
  assign n24872 = ~n24871 | ~n24870;
  assign n24877 = ~n24873 & ~n24872;
  assign n25303 = ~n24874 & ~P2_U3088;
  assign n24876 = ~n24875 | ~n25303;
  assign P2_U3230 = ~n24877 | ~n24876;
  assign n24878 = ~P2_ADDR_REG_17__SCAN_IN | ~n24913;
  assign n24881 = ~n24879 | ~n24878;
  assign n25300 = ~n24903 | ~P2_STATE_REG_SCAN_IN;
  assign n24880 = ~n24896 & ~n25300;
  assign n24893 = ~n24881 & ~n24880;
  assign n24885 = ~n24903;
  assign n24905 = P2_REG1_REG_17__SCAN_IN ^ ~n24885;
  assign n24883 = ~P2_REG1_REG_16__SCAN_IN | ~n24886;
  assign n24904 = ~n24883 | ~n24882;
  assign n24884 = n24905 ^ ~n24904;
  assign n24891 = ~n24884 & ~n24925;
  assign n24900 = P2_REG2_REG_17__SCAN_IN ^ ~n24885;
  assign n24888 = ~P2_REG2_REG_16__SCAN_IN | ~n24886;
  assign n24899 = ~n24888 | ~n24887;
  assign n24889 = n24900 ^ ~n24899;
  assign n24890 = ~n24889 & ~n24933;
  assign n24892 = ~n24891 & ~n24890;
  assign P2_U3231 = ~n24893 | ~n24892;
  assign n24894 = ~P2_ADDR_REG_18__SCAN_IN | ~n24913;
  assign n24898 = ~n24895 | ~n24894;
  assign n25294 = ~n24928 | ~P2_STATE_REG_SCAN_IN;
  assign n24897 = ~n24896 & ~n25294;
  assign n24912 = ~n24898 & ~n24897;
  assign n24901 = ~P2_REG2_REG_17__SCAN_IN | ~n24903;
  assign n24929 = n24928 ^ ~n24927;
  assign n24902 = P2_REG2_REG_18__SCAN_IN ^ n24929;
  assign n24910 = ~n24902 & ~n24933;
  assign n24907 = ~P2_REG1_REG_17__SCAN_IN | ~n24903;
  assign n24906 = ~n24905 | ~n24904;
  assign n24920 = ~n24907 | ~n24906;
  assign n24919 = n24928 ^ n24920;
  assign n24908 = n24919 ^ ~P2_REG1_REG_18__SCAN_IN;
  assign n24909 = ~n24908 & ~n24925;
  assign n24911 = ~n24910 & ~n24909;
  assign P2_U3232 = ~n24912 | ~n24911;
  assign n24914 = ~P2_ADDR_REG_19__SCAN_IN | ~n24913;
  assign n24918 = ~n24915 | ~n24914;
  assign n24917 = ~n24916 & ~n17029;
  assign n24938 = ~n24918 & ~n24917;
  assign n24922 = ~P2_REG1_REG_18__SCAN_IN | ~n24919;
  assign n24921 = ~n24928 | ~n24920;
  assign n24924 = ~n24922 | ~n24921;
  assign n24923 = P2_REG1_REG_19__SCAN_IN ^ n25194;
  assign n24926 = n24924 ^ ~n24923;
  assign n24936 = ~n24926 & ~n24925;
  assign n24931 = ~n24928 & ~n24927;
  assign n24930 = ~P2_REG2_REG_18__SCAN_IN & ~n24929;
  assign n24932 = ~n24931 & ~n24930;
  assign n24935 = ~n24934 & ~n24933;
  assign n24937 = ~n24936 & ~n24935;
  assign P2_U3233 = ~n24938 | ~n24937;
  assign n24940 = ~n25264 | ~n25506;
  assign n24939 = ~n25282 | ~P2_REG2_REG_11__SCAN_IN;
  assign n24943 = ~n24940 | ~n24939;
  assign n24942 = ~n24941 & ~n25267;
  assign n24963 = ~n24943 & ~n24942;
  assign n25504 = n24982 ^ ~n25506;
  assign n24946 = ~n25263 | ~n25504;
  assign n25510 = n24944 ^ ~n24947;
  assign n24952 = ~n25510;
  assign n25226 = ~n25099;
  assign n24945 = ~n24952 | ~n25226;
  assign n24961 = ~n24946 | ~n24945;
  assign n24949 = ~n24948 | ~n24947;
  assign n24951 = ~n24950 | ~n24949;
  assign n24954 = ~n24951 | ~n25246;
  assign n24953 = ~n24952 | ~n25248;
  assign n24959 = ~n24954 | ~n24953;
  assign n24957 = ~n24955 | ~n25273;
  assign n24956 = ~n25000 | ~n25253;
  assign n24958 = ~n24957 | ~n24956;
  assign n25514 = ~n24959 & ~n24958;
  assign n24960 = ~n25282 & ~n25514;
  assign n24962 = ~n24961 & ~n24960;
  assign P2_U3254 = ~n24963 | ~n24962;
  assign n24966 = ~n25233 | ~n24964;
  assign n24965 = ~n25282 | ~P2_REG2_REG_10__SCAN_IN;
  assign n24981 = ~n24966 | ~n24965;
  assign n24968 = n24967 ^ ~n24969;
  assign n24975 = ~n24968 | ~n25246;
  assign n25492 = n24970 ^ ~n24969;
  assign n25271 = ~n25248;
  assign n24973 = ~n25492 & ~n25271;
  assign n24972 = ~n24971 & ~n25079;
  assign n24974 = ~n24973 & ~n24972;
  assign n25498 = ~n24975 | ~n24974;
  assign n24977 = ~n25489 | ~n25189;
  assign n25490 = ~n24976 | ~n25273;
  assign n24978 = ~n24977 | ~n25490;
  assign n24979 = ~n25498 & ~n24978;
  assign n24980 = ~n25282 & ~n24979;
  assign n24989 = ~n24981 & ~n24980;
  assign n25068 = ~n25263;
  assign n24985 = ~n24982;
  assign n24990 = ~n25479;
  assign n24983 = ~n25017 | ~n24990;
  assign n24984 = ~n24983 | ~n25489;
  assign n25496 = ~n24985 | ~n24984;
  assign n24987 = ~n25068 & ~n25496;
  assign n24986 = ~n25492 & ~n25099;
  assign n24988 = ~n24987 & ~n24986;
  assign P2_U3255 = ~n24989 | ~n24988;
  assign n24991 = n25017 ^ ~n24990;
  assign n25495 = ~n25503;
  assign n25483 = ~n24991 & ~n25495;
  assign n24993 = ~n25483 | ~n17029;
  assign n24992 = ~n25479 | ~n25189;
  assign n25007 = ~n24993 | ~n24992;
  assign n24995 = n24994 ^ ~n24997;
  assign n24999 = ~n24995 | ~n25246;
  assign n25478 = n24997 ^ n24996;
  assign n24998 = ~n25478 | ~n25248;
  assign n25004 = ~n24999 | ~n24998;
  assign n25002 = ~n25000 | ~n25273;
  assign n25001 = ~n25049 | ~n25253;
  assign n25003 = ~n25002 | ~n25001;
  assign n25485 = ~n25004 & ~n25003;
  assign n25005 = ~n25478 | ~n25277;
  assign n25006 = ~n25485 | ~n25005;
  assign n25008 = ~n25007 & ~n25006;
  assign n25011 = ~n25282 & ~n25008;
  assign n25010 = ~n25267 & ~n25009;
  assign n25013 = ~n25011 & ~n25010;
  assign n25012 = ~P2_REG2_REG_9__SCAN_IN | ~n25282;
  assign P2_U3256 = ~n25013 | ~n25012;
  assign n25015 = ~n25264 | ~n25467;
  assign n25014 = ~n25282 | ~P2_REG2_REG_8__SCAN_IN;
  assign n25020 = ~n25015 | ~n25014;
  assign n25060 = ~n25454;
  assign n25016 = ~n25067 | ~n25060;
  assign n25018 = n25016 & n25467;
  assign n25466 = n25018 | n25017;
  assign n25019 = ~n25068 & ~n25466;
  assign n25039 = ~n25020 & ~n25019;
  assign n25024 = ~n25021 | ~n25273;
  assign n25023 = ~n25022 | ~n25253;
  assign n25027 = ~n25024 | ~n25023;
  assign n25470 = n25025 ^ ~n25029;
  assign n25026 = ~n25470 & ~n25271;
  assign n25032 = ~n25027 & ~n25026;
  assign n25030 = n25028 ^ ~n25029;
  assign n25031 = ~n25030 | ~n25246;
  assign n25472 = ~n25032 | ~n25031;
  assign n25034 = ~n25033 & ~n25267;
  assign n25035 = ~n25472 & ~n25034;
  assign n25037 = ~n25282 & ~n25035;
  assign n25036 = ~n25099 & ~n25470;
  assign n25038 = ~n25037 & ~n25036;
  assign P2_U3257 = ~n25039 | ~n25038;
  assign n25041 = ~n25040;
  assign n25044 = ~n25042 | ~n13274;
  assign n25084 = ~n25044 | ~n25043;
  assign n25047 = ~n25084 & ~n25076;
  assign n25046 = ~n25045;
  assign n25048 = ~n25047 & ~n25046;
  assign n25056 = n25048 ^ ~n25052;
  assign n25453 = ~n25056;
  assign n25050 = ~n25453 | ~n25277;
  assign n25455 = ~n25049 | ~n25273;
  assign n25065 = ~n25050 | ~n25455;
  assign n25053 = n25051 ^ ~n25052;
  assign n25055 = ~n25053 | ~n25246;
  assign n25054 = ~n25126 | ~n25253;
  assign n25058 = ~n25055 | ~n25054;
  assign n25057 = ~n25056 & ~n25271;
  assign n25463 = ~n25058 & ~n25057;
  assign n25062 = ~n25267 & ~n25059;
  assign n25061 = ~n25060 & ~n25091;
  assign n25063 = ~n25062 & ~n25061;
  assign n25064 = ~n25463 | ~n25063;
  assign n25066 = ~n25065 & ~n25064;
  assign n25070 = ~n25282 & ~n25066;
  assign n25457 = n25454 ^ n25067;
  assign n25069 = ~n25068 & ~n25457;
  assign n25072 = ~n25070 & ~n25069;
  assign n25071 = ~P2_REG2_REG_7__SCAN_IN | ~n25282;
  assign P2_U3258 = ~n25072 | ~n25071;
  assign n25075 = P2_REG2_REG_6__SCAN_IN & n25282;
  assign n25074 = ~n25267 & ~n25073;
  assign n25103 = ~n25075 & ~n25074;
  assign n25078 = n25077 ^ ~n25076;
  assign n25082 = ~n25078 & ~n25270;
  assign n25081 = ~n25080 & ~n25079;
  assign n25087 = ~n25082 & ~n25081;
  assign n25446 = n25084 ^ ~n25083;
  assign n25085 = ~n25446;
  assign n25086 = ~n25085 | ~n25248;
  assign n25448 = ~n25087 | ~n25086;
  assign n25089 = n25088 ^ ~n25090;
  assign n25445 = ~n25089 & ~n25495;
  assign n25096 = ~n25445 | ~n17029;
  assign n25094 = ~n13983 & ~n25091;
  assign n25442 = ~n25093 & ~n25092;
  assign n25095 = ~n25094 & ~n25442;
  assign n25097 = ~n25096 | ~n25095;
  assign n25098 = ~n25448 & ~n25097;
  assign n25101 = ~n25282 & ~n25098;
  assign n25100 = ~n25099 & ~n25446;
  assign n25102 = ~n25101 & ~n25100;
  assign P2_U3259 = ~n25103 | ~n25102;
  assign n25110 = ~n25105 & ~n25104;
  assign n25108 = ~n25233 | ~n25106;
  assign n25107 = ~n25282 | ~P2_REG2_REG_5__SCAN_IN;
  assign n25109 = ~n25108 | ~n25107;
  assign n25134 = ~n25110 & ~n25109;
  assign n25431 = n13142 ^ ~n25432;
  assign n25117 = ~n25263 | ~n25431;
  assign n25112 = ~n25111;
  assign n25113 = ~n25112 & ~n25142;
  assign n25115 = ~n25139 | ~n25114;
  assign n25429 = n25115 ^ ~n25122;
  assign n25116 = ~n25226 | ~n25429;
  assign n25132 = ~n25117 | ~n25116;
  assign n25143 = n25118 | n25119;
  assign n25144 = ~n25143 | ~n25142;
  assign n25121 = ~n25144 | ~n25120;
  assign n25123 = n25122 ^ n25121;
  assign n25125 = ~n25123 | ~n25246;
  assign n25124 = ~n25429 | ~n25248;
  assign n25130 = ~n25125 | ~n25124;
  assign n25128 = ~n25126 | ~n25273;
  assign n25127 = ~n25183 | ~n25253;
  assign n25129 = ~n25128 | ~n25127;
  assign n25438 = ~n25130 & ~n25129;
  assign n25131 = ~n25282 & ~n25438;
  assign n25133 = ~n25132 & ~n25131;
  assign P2_U3260 = ~n25134 | ~n25133;
  assign n25171 = n25219 & n25135;
  assign n25177 = ~n25136;
  assign n25173 = ~n25171 & ~n25177;
  assign n25138 = ~n25137 | ~n25142;
  assign n25141 = ~n25173 & ~n25138;
  assign n25140 = ~n25139;
  assign n25419 = ~n25141 & ~n25140;
  assign n25147 = ~n25419;
  assign n25167 = ~n25147 | ~n25277;
  assign n25145 = n25143 | n25142;
  assign n25146 = ~n25145 | ~n25144;
  assign n25149 = ~n25146 | ~n25246;
  assign n25148 = ~n25147 | ~n25248;
  assign n25154 = ~n25149 | ~n25148;
  assign n25152 = ~n25150 | ~n25273;
  assign n25151 = ~n25214 | ~n25253;
  assign n25153 = ~n25152 | ~n25151;
  assign n25426 = ~n25154 & ~n25153;
  assign n25159 = ~n13142 & ~n25495;
  assign n25192 = ~n25155;
  assign n25157 = ~n25192 | ~n25156;
  assign n25158 = ~n25157 | ~n25420;
  assign n25422 = ~n25159 | ~n25158;
  assign n25164 = ~n25422 & ~n25194;
  assign n25162 = ~n25233 | ~n25160;
  assign n25161 = ~n25189 | ~n25420;
  assign n25163 = ~n25162 | ~n25161;
  assign n25165 = ~n25164 & ~n25163;
  assign n25166 = n25426 & n25165;
  assign n25168 = ~n25167 | ~n25166;
  assign n25170 = ~n25284 | ~n25168;
  assign n25169 = ~n25282 | ~P2_REG2_REG_4__SCAN_IN;
  assign P2_U3261 = ~n25170 | ~n25169;
  assign n25172 = n25171 & n25177;
  assign n25409 = ~n25173 & ~n25172;
  assign n25180 = ~n25409;
  assign n25199 = ~n25180 | ~n25277;
  assign n25211 = ~n25209 | ~n25174;
  assign n25176 = ~n25211 | ~n25175;
  assign n25178 = ~n25177 & ~n25176;
  assign n25179 = n25118 | n25178;
  assign n25182 = ~n25179 | ~n25246;
  assign n25181 = ~n25180 | ~n25248;
  assign n25187 = ~n25182 | ~n25181;
  assign n25185 = ~n25183 | ~n25273;
  assign n25184 = ~n25252 | ~n25253;
  assign n25186 = ~n25185 | ~n25184;
  assign n25416 = ~n25187 & ~n25186;
  assign n25191 = ~n25233 | ~n25188;
  assign n25190 = ~n25410 | ~n25189;
  assign n25196 = ~n25191 | ~n25190;
  assign n25193 = n25192 ^ ~n25410;
  assign n25412 = ~n25193 | ~n25503;
  assign n25195 = ~n25412 & ~n25194;
  assign n25197 = ~n25196 & ~n25195;
  assign n25198 = n25416 & n25197;
  assign n25200 = ~n25199 | ~n25198;
  assign n25202 = ~n25284 | ~n25200;
  assign n25201 = ~n25282 | ~P2_REG2_REG_3__SCAN_IN;
  assign P2_U3262 = ~n25202 | ~n25201;
  assign n25203 = ~P2_REG2_REG_2__SCAN_IN;
  assign n25205 = ~n25284 & ~n25203;
  assign n25204 = ~n25267 & ~n16613;
  assign n25232 = ~n25205 & ~n25204;
  assign n25208 = ~n25264 | ~n25399;
  assign n25398 = n25206 ^ n25399;
  assign n25207 = ~n25263 | ~n25398;
  assign n25230 = ~n25208 | ~n25207;
  assign n25210 = ~n25209;
  assign n25212 = ~n25210 | ~n25217;
  assign n25213 = ~n25212 | ~n25211;
  assign n25225 = ~n25213 | ~n25246;
  assign n25216 = ~n25214 | ~n25273;
  assign n25215 = ~n25274 | ~n25253;
  assign n25223 = ~n25216 | ~n25215;
  assign n25220 = n25218 | n25217;
  assign n25404 = ~n25220 | ~n25219;
  assign n25221 = ~n25404;
  assign n25222 = ~n25221 & ~n25271;
  assign n25224 = ~n25223 & ~n25222;
  assign n25403 = ~n25225 | ~n25224;
  assign n25228 = ~n25403 | ~n25284;
  assign n25227 = ~n25226 | ~n25404;
  assign n25229 = ~n25228 | ~n25227;
  assign n25231 = ~n25230 & ~n25229;
  assign P2_U3263 = ~n25232 | ~n25231;
  assign n25235 = ~n25282 | ~P2_REG2_REG_1__SCAN_IN;
  assign n25234 = ~n25233 | ~P2_REG3_REG_1__SCAN_IN;
  assign n25239 = ~n25235 | ~n25234;
  assign n25237 = ~n25264 | ~n25389;
  assign n25388 = n25389 ^ ~n14816;
  assign n25236 = ~n25263 | ~n25388;
  assign n25238 = ~n25237 | ~n25236;
  assign n25262 = ~n25239 & ~n25238;
  assign n25242 = ~n25241;
  assign n25387 = ~n25243 & ~n25242;
  assign n25249 = ~n25387;
  assign n25259 = ~n25249 | ~n25277;
  assign n25247 = n25245 ^ ~n25244;
  assign n25251 = ~n25247 | ~n25246;
  assign n25250 = ~n25249 | ~n25248;
  assign n25258 = ~n25251 | ~n25250;
  assign n25256 = ~n25252 | ~n25273;
  assign n25255 = ~n25254 | ~n25253;
  assign n25257 = ~n25256 | ~n25255;
  assign n25395 = ~n25258 & ~n25257;
  assign n25260 = ~n25259 | ~n25395;
  assign n25261 = ~n25260 | ~n25284;
  assign P2_U3264 = ~n25262 | ~n25261;
  assign n25265 = ~n25264 & ~n25263;
  assign n25269 = ~n25265 & ~n14816;
  assign n25268 = ~n25267 & ~n25266;
  assign n25288 = ~n25269 & ~n25268;
  assign n25382 = ~n25279;
  assign n25272 = ~n25271 | ~n25270;
  assign n25276 = ~n25382 | ~n25272;
  assign n25275 = ~n25274 | ~n25273;
  assign n25381 = ~n25276 | ~n25275;
  assign n25278 = ~n25277;
  assign n25280 = ~n25279 & ~n25278;
  assign n25281 = ~n25381 & ~n25280;
  assign n25286 = ~n25282 & ~n25281;
  assign n25285 = ~n25284 & ~n25283;
  assign n25287 = ~n25286 & ~n25285;
  assign P2_U3265 = ~n25288 | ~n25287;
  assign P2_U3266 = P2_D_REG_31__SCAN_IN & n25368;
  assign P2_U3267 = P2_D_REG_30__SCAN_IN & n25368;
  assign P2_U3268 = P2_D_REG_29__SCAN_IN & n25368;
  assign P2_U3269 = P2_D_REG_28__SCAN_IN & n25368;
  assign n25375 = ~n25368;
  assign n25369 = ~n25375;
  assign P2_U3270 = P2_D_REG_27__SCAN_IN & n25369;
  assign P2_U3271 = P2_D_REG_26__SCAN_IN & n25368;
  assign P2_U3272 = P2_D_REG_25__SCAN_IN & n25368;
  assign P2_U3273 = P2_D_REG_24__SCAN_IN & n25368;
  assign P2_U3274 = P2_D_REG_23__SCAN_IN & n25368;
  assign P2_U3275 = P2_D_REG_22__SCAN_IN & n25368;
  assign P2_U3276 = P2_D_REG_21__SCAN_IN & n25368;
  assign P2_U3277 = P2_D_REG_20__SCAN_IN & n25368;
  assign P2_U3278 = P2_D_REG_19__SCAN_IN & n25368;
  assign P2_U3279 = P2_D_REG_18__SCAN_IN & n25368;
  assign P2_U3280 = P2_D_REG_17__SCAN_IN & n25368;
  assign P2_U3281 = P2_D_REG_16__SCAN_IN & n25369;
  assign P2_U3282 = P2_D_REG_15__SCAN_IN & n25369;
  assign P2_U3283 = P2_D_REG_14__SCAN_IN & n25368;
  assign P2_U3284 = P2_D_REG_13__SCAN_IN & n25368;
  assign P2_U3285 = P2_D_REG_12__SCAN_IN & n25368;
  assign P2_U3286 = P2_D_REG_11__SCAN_IN & n25368;
  assign P2_U3287 = P2_D_REG_10__SCAN_IN & n25368;
  assign P2_U3288 = P2_D_REG_9__SCAN_IN & n25368;
  assign P2_U3289 = P2_D_REG_8__SCAN_IN & n25368;
  assign P2_U3290 = P2_D_REG_7__SCAN_IN & n25368;
  assign P2_U3291 = P2_D_REG_6__SCAN_IN & n25368;
  assign P2_U3292 = P2_D_REG_5__SCAN_IN & n25368;
  assign P2_U3293 = P2_D_REG_4__SCAN_IN & n25368;
  assign P2_U3294 = P2_D_REG_3__SCAN_IN & n25368;
  assign P2_U3295 = P2_D_REG_2__SCAN_IN & n25368;
  assign n25293 = ~n25290 & ~n25360;
  assign n25292 = ~n25337 & ~n25291;
  assign n25295 = ~n25293 & ~n25292;
  assign P2_U3309 = ~n25295 | ~n25294;
  assign n25299 = ~n25296 & ~n25360;
  assign n25298 = ~n25337 & ~n25297;
  assign n25301 = ~n25299 & ~n25298;
  assign P2_U3310 = ~n25301 | ~n25300;
  assign n25304 = ~n25302 & ~n25360;
  assign n25306 = ~n25304 & ~n25303;
  assign n25305 = ~n25365 | ~P1_DATAO_REG_16__SCAN_IN;
  assign P2_U3311 = ~n25306 | ~n25305;
  assign n25308 = ~n24052 & ~n25360;
  assign n25310 = ~n25308 & ~n25307;
  assign n25309 = ~n25365 | ~P1_DATAO_REG_14__SCAN_IN;
  assign P2_U3313 = ~n25310 | ~n25309;
  assign n25313 = ~n25311 & ~n25360;
  assign n25315 = ~n25313 & ~n25312;
  assign n25314 = ~n25365 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P2_U3314 = ~n25315 | ~n25314;
  assign n25317 = ~n24065 & ~n25360;
  assign n25319 = ~n25317 & ~n25316;
  assign n25318 = ~n25365 | ~P1_DATAO_REG_12__SCAN_IN;
  assign P2_U3315 = ~n25319 | ~n25318;
  assign n25322 = ~n25320 & ~n25360;
  assign n25324 = ~n25322 & ~n25321;
  assign n25323 = ~n25365 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P2_U3316 = ~n25324 | ~n25323;
  assign n25327 = ~n25325 & ~n25360;
  assign n25329 = ~n25327 & ~n25326;
  assign n25328 = ~n25365 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P2_U3317 = ~n25329 | ~n25328;
  assign n25332 = ~n25330 & ~n25360;
  assign n25334 = ~n25332 & ~n25331;
  assign n25333 = ~n25365 | ~P1_DATAO_REG_9__SCAN_IN;
  assign P2_U3318 = ~n25334 | ~n25333;
  assign n25339 = ~n25335 & ~n25360;
  assign n25338 = ~n25337 & ~n25336;
  assign n25341 = ~n25339 & ~n25338;
  assign P2_U3319 = ~n25341 | ~n25340;
  assign n25345 = ~n25342 & ~n25360;
  assign n25344 = ~n25343 & ~P2_U3088;
  assign n25347 = ~n25345 & ~n25344;
  assign n25346 = ~n25365 | ~P1_DATAO_REG_7__SCAN_IN;
  assign P2_U3320 = ~n25347 | ~n25346;
  assign n25351 = ~n25348 & ~n25360;
  assign n25350 = ~n25349 & ~P2_U3088;
  assign n25353 = ~n25351 & ~n25350;
  assign n25352 = ~n25365 | ~P1_DATAO_REG_6__SCAN_IN;
  assign P2_U3321 = ~n25353 | ~n25352;
  assign n25357 = ~n25354 & ~n25360;
  assign n25356 = ~n25355 & ~P2_U3088;
  assign n25359 = ~n25357 & ~n25356;
  assign n25358 = ~n25365 | ~P1_DATAO_REG_4__SCAN_IN;
  assign P2_U3323 = ~n25359 | ~n25358;
  assign n25364 = ~n25361 & ~n25360;
  assign n25363 = ~n13793 & ~P2_U3088;
  assign n25367 = ~n25364 & ~n25363;
  assign n25366 = ~n25365 | ~P1_DATAO_REG_2__SCAN_IN;
  assign P2_U3325 = ~n25367 | ~n25366;
  assign n25372 = ~P2_D_REG_0__SCAN_IN | ~n25368;
  assign n25371 = n25370 | n25369;
  assign P2_U3416 = ~n25372 | ~n25371;
  assign n25377 = n25374 & n25373;
  assign n25376 = ~P2_D_REG_1__SCAN_IN & ~n25375;
  assign P2_U3417 = ~n25377 & ~n25376;
  assign n25386 = ~P2_REG0_REG_0__SCAN_IN | ~n25488;
  assign n25379 = ~n25378;
  assign n25380 = ~n25379 & ~n14816;
  assign n25384 = ~n25381 & ~n25380;
  assign n25383 = ~n25382 | ~n25477;
  assign n25518 = ~n25384 | ~n25383;
  assign n25385 = ~n25515 | ~n25518;
  assign P2_U3430 = ~n25386 | ~n25385;
  assign n25397 = ~P2_REG0_REG_1__SCAN_IN | ~n25488;
  assign n25393 = ~n25387 & ~n25509;
  assign n25391 = ~n25388 | ~n25503;
  assign n25390 = ~n25505 | ~n25389;
  assign n25392 = ~n25391 | ~n25390;
  assign n25394 = ~n25393 & ~n25392;
  assign n25521 = ~n25395 | ~n25394;
  assign n25396 = ~n25515 | ~n25521;
  assign P2_U3433 = ~n25397 | ~n25396;
  assign n25408 = ~P2_REG0_REG_2__SCAN_IN | ~n25488;
  assign n25401 = ~n25398 | ~n25503;
  assign n25400 = ~n25399 | ~n25505;
  assign n25402 = ~n25401 | ~n25400;
  assign n25406 = ~n25403 & ~n25402;
  assign n25405 = ~n25404 | ~n25477;
  assign n25524 = ~n25406 | ~n25405;
  assign n25407 = ~n25515 | ~n25524;
  assign P2_U3436 = ~n25408 | ~n25407;
  assign n25418 = ~P2_REG0_REG_3__SCAN_IN | ~n25488;
  assign n25414 = ~n25409 & ~n25509;
  assign n25411 = ~n25410 | ~n25505;
  assign n25413 = ~n25412 | ~n25411;
  assign n25415 = ~n25414 & ~n25413;
  assign n25527 = ~n25416 | ~n25415;
  assign n25417 = ~n25515 | ~n25527;
  assign P2_U3439 = ~n25418 | ~n25417;
  assign n25428 = ~P2_REG0_REG_4__SCAN_IN | ~n25488;
  assign n25424 = ~n25419 & ~n25509;
  assign n25421 = ~n25505 | ~n25420;
  assign n25423 = ~n25422 | ~n25421;
  assign n25425 = ~n25424 & ~n25423;
  assign n25530 = ~n25426 | ~n25425;
  assign n25427 = ~n25515 | ~n25530;
  assign P2_U3442 = ~n25428 | ~n25427;
  assign n25440 = ~P2_REG0_REG_5__SCAN_IN | ~n25488;
  assign n25430 = ~n25429;
  assign n25436 = ~n25430 & ~n25509;
  assign n25434 = ~n25431 | ~n25503;
  assign n25433 = ~n25505 | ~n25432;
  assign n25435 = ~n25434 | ~n25433;
  assign n25437 = ~n25436 & ~n25435;
  assign n25533 = ~n25438 | ~n25437;
  assign n25439 = ~n25515 | ~n25533;
  assign P2_U3445 = ~n25440 | ~n25439;
  assign n25452 = ~P2_REG0_REG_6__SCAN_IN | ~n25488;
  assign n25443 = ~n13983 & ~n25441;
  assign n25444 = n25443 | n25442;
  assign n25450 = ~n25445 & ~n25444;
  assign n25447 = ~n25446 & ~n25509;
  assign n25449 = ~n25448 & ~n25447;
  assign n25536 = ~n25450 | ~n25449;
  assign n25451 = ~n25515 | ~n25536;
  assign P2_U3448 = ~n25452 | ~n25451;
  assign n25465 = ~P2_REG0_REG_7__SCAN_IN | ~n25488;
  assign n25461 = ~n25453 | ~n25477;
  assign n25456 = ~n25454 | ~n25505;
  assign n25459 = ~n25456 | ~n25455;
  assign n25458 = ~n25457 & ~n25495;
  assign n25460 = ~n25459 & ~n25458;
  assign n25462 = n25461 & n25460;
  assign n25539 = ~n25463 | ~n25462;
  assign n25464 = ~n25515 | ~n25539;
  assign P2_U3451 = ~n25465 | ~n25464;
  assign n25476 = ~P2_REG0_REG_8__SCAN_IN | ~n25488;
  assign n25469 = ~n25466 & ~n25495;
  assign n25468 = n25467 & n25505;
  assign n25474 = ~n25469 & ~n25468;
  assign n25471 = ~n25470 & ~n25509;
  assign n25473 = ~n25472 & ~n25471;
  assign n25542 = ~n25474 | ~n25473;
  assign n25475 = ~n25515 | ~n25542;
  assign P2_U3454 = ~n25476 | ~n25475;
  assign n25487 = ~P2_REG0_REG_9__SCAN_IN | ~n25488;
  assign n25481 = ~n25478 | ~n25477;
  assign n25480 = ~n25479 | ~n25505;
  assign n25482 = ~n25481 | ~n25480;
  assign n25484 = ~n25483 & ~n25482;
  assign n25545 = ~n25485 | ~n25484;
  assign n25486 = ~n25515 | ~n25545;
  assign P2_U3457 = ~n25487 | ~n25486;
  assign n25502 = ~P2_REG0_REG_10__SCAN_IN | ~n25488;
  assign n25491 = ~n25489 | ~n25505;
  assign n25494 = ~n25491 | ~n25490;
  assign n25493 = ~n25492 & ~n25509;
  assign n25500 = ~n25494 & ~n25493;
  assign n25497 = ~n25496 & ~n25495;
  assign n25499 = ~n25498 & ~n25497;
  assign n25548 = ~n25500 | ~n25499;
  assign n25501 = ~n25515 | ~n25548;
  assign P2_U3460 = ~n25502 | ~n25501;
  assign n25517 = ~P2_REG0_REG_11__SCAN_IN | ~n25488;
  assign n25508 = ~n25504 | ~n25503;
  assign n25507 = ~n25506 | ~n25505;
  assign n25512 = ~n25508 | ~n25507;
  assign n25511 = ~n25510 & ~n25509;
  assign n25513 = ~n25512 & ~n25511;
  assign n25552 = ~n25514 | ~n25513;
  assign n25516 = ~n25515 | ~n25552;
  assign P2_U3463 = ~n25517 | ~n25516;
  assign n25520 = ~P2_REG1_REG_0__SCAN_IN | ~n25551;
  assign n25519 = ~n25553 | ~n25518;
  assign P2_U3499 = ~n25520 | ~n25519;
  assign n25523 = ~P2_REG1_REG_1__SCAN_IN | ~n25551;
  assign n25522 = ~n25553 | ~n25521;
  assign P2_U3500 = ~n25523 | ~n25522;
  assign n25526 = ~P2_REG1_REG_2__SCAN_IN | ~n25551;
  assign n25525 = ~n25553 | ~n25524;
  assign P2_U3501 = ~n25526 | ~n25525;
  assign n25529 = ~P2_REG1_REG_3__SCAN_IN | ~n25551;
  assign n25528 = ~n25553 | ~n25527;
  assign P2_U3502 = ~n25529 | ~n25528;
  assign n25532 = ~P2_REG1_REG_4__SCAN_IN | ~n25551;
  assign n25531 = ~n25553 | ~n25530;
  assign P2_U3503 = ~n25532 | ~n25531;
  assign n25535 = ~P2_REG1_REG_5__SCAN_IN | ~n25551;
  assign n25534 = ~n25553 | ~n25533;
  assign P2_U3504 = ~n25535 | ~n25534;
  assign n25538 = ~P2_REG1_REG_6__SCAN_IN | ~n25551;
  assign n25537 = ~n25553 | ~n25536;
  assign P2_U3505 = ~n25538 | ~n25537;
  assign n25541 = ~P2_REG1_REG_7__SCAN_IN | ~n25551;
  assign n25540 = ~n25553 | ~n25539;
  assign P2_U3506 = ~n25541 | ~n25540;
  assign n25544 = ~P2_REG1_REG_8__SCAN_IN | ~n25551;
  assign n25543 = ~n25553 | ~n25542;
  assign P2_U3507 = ~n25544 | ~n25543;
  assign n25547 = ~P2_REG1_REG_9__SCAN_IN | ~n25551;
  assign n25546 = ~n25553 | ~n25545;
  assign P2_U3508 = ~n25547 | ~n25546;
  assign n25550 = ~P2_REG1_REG_10__SCAN_IN | ~n25551;
  assign n25549 = ~n25553 | ~n25548;
  assign P2_U3509 = ~n25550 | ~n25549;
  assign n25555 = ~P2_REG1_REG_11__SCAN_IN | ~n25551;
  assign n25554 = ~n25553 | ~n25552;
  assign P2_U3510 = ~n25555 | ~n25554;
  assign n25558 = ~P2_DATAO_REG_19__SCAN_IN | ~n25592;
  assign n25557 = ~P2_U3947 | ~n25556;
  assign P2_U3550 = ~n25558 | ~n25557;
  assign n25561 = ~P2_DATAO_REG_20__SCAN_IN | ~n25592;
  assign n25560 = ~P2_U3947 | ~n25559;
  assign P2_U3551 = ~n25561 | ~n25560;
  assign n25564 = ~P2_DATAO_REG_21__SCAN_IN | ~n25592;
  assign n25563 = ~P2_U3947 | ~n25562;
  assign P2_U3552 = ~n25564 | ~n25563;
  assign n25567 = ~P2_DATAO_REG_22__SCAN_IN | ~n25592;
  assign n25566 = ~P2_U3947 | ~n25565;
  assign P2_U3553 = ~n25567 | ~n25566;
  assign n25570 = ~P2_DATAO_REG_23__SCAN_IN | ~n25592;
  assign n25569 = ~P2_U3947 | ~n25568;
  assign P2_U3554 = ~n25570 | ~n25569;
  assign n25573 = ~P2_DATAO_REG_24__SCAN_IN | ~n25592;
  assign n25572 = ~P2_U3947 | ~n25571;
  assign P2_U3555 = ~n25573 | ~n25572;
  assign n25576 = ~P2_DATAO_REG_25__SCAN_IN | ~n25592;
  assign n25575 = ~P2_U3947 | ~n25574;
  assign P2_U3556 = ~n25576 | ~n25575;
  assign n25579 = ~P2_DATAO_REG_26__SCAN_IN | ~n25592;
  assign n25578 = ~P2_U3947 | ~n25577;
  assign P2_U3557 = ~n25579 | ~n25578;
  assign n25582 = ~P2_DATAO_REG_27__SCAN_IN | ~n25592;
  assign n25581 = ~P2_U3947 | ~n25580;
  assign P2_U3558 = ~n25582 | ~n25581;
  assign n25585 = ~P2_DATAO_REG_28__SCAN_IN | ~n25592;
  assign n25584 = ~P2_U3947 | ~n25583;
  assign P2_U3559 = ~n25585 | ~n25584;
  assign n25588 = ~P2_DATAO_REG_29__SCAN_IN | ~n25592;
  assign n25587 = ~P2_U3947 | ~n25586;
  assign P2_U3560 = ~n25588 | ~n25587;
  assign n25591 = ~P2_DATAO_REG_30__SCAN_IN | ~n25592;
  assign n25590 = ~P2_U3947 | ~n25589;
  assign P2_U3561 = ~n25591 | ~n25590;
  assign n25595 = ~P2_DATAO_REG_31__SCAN_IN | ~n25592;
  assign n25594 = ~P2_U3947 | ~n25593;
  assign P2_U3562 = ~n25595 | ~n25594;
  assign P3_U3150 = ~P3_U3897 & ~n26033;
  assign n25596 = ~n25724 & ~n26138;
  assign n25880 = P3_U3151 & P3_REG3_REG_7__SCAN_IN;
  assign n25610 = ~n25596 & ~n25880;
  assign n25599 = ~n25728 | ~n26086;
  assign n25708 = ~n25725;
  assign n25598 = ~n25708 | ~n25597;
  assign n25608 = ~n25599 | ~n25598;
  assign n25601 = ~n25730 | ~n25731;
  assign n25602 = ~n25601 | ~n25600;
  assign n25604 = n25603 ^ n25602;
  assign n25606 = ~n25604 | ~n25732;
  assign n25605 = ~n25734 | ~n26141;
  assign n25607 = ~n25606 | ~n25605;
  assign n25609 = ~n25608 & ~n25607;
  assign P3_U3153 = ~n25610 | ~n25609;
  assign n25613 = ~n26393 & ~n25725;
  assign n25612 = ~n25666 & ~n25611;
  assign n25623 = ~n25613 & ~n25612;
  assign n25614 = ~n25706 | ~n26116;
  assign n25954 = ~P3_REG3_REG_10__SCAN_IN | ~P3_U3151;
  assign n25621 = ~n25614 | ~n25954;
  assign n25617 = n25616 ^ n25615;
  assign n25619 = ~n25617 | ~n25732;
  assign n25618 = ~n25734 | ~n26067;
  assign n25620 = ~n25619 | ~n25618;
  assign n25622 = ~n25621 & ~n25620;
  assign P3_U3157 = ~n25623 | ~n25622;
  assign n25625 = ~n25666 & ~n25624;
  assign n25798 = ~P3_STATE_REG_SCAN_IN & ~n16443;
  assign n25637 = ~n25625 & ~n25798;
  assign n25628 = ~n25706 | ~n26286;
  assign n25627 = ~n25708 | ~n25626;
  assign n25635 = ~n25628 | ~n25627;
  assign n25631 = n25629 ^ n25630;
  assign n25633 = ~n25631 | ~n25732;
  assign n25632 = ~n25734 | ~n16443;
  assign n25634 = ~n25633 | ~n25632;
  assign n25636 = ~n25635 & ~n25634;
  assign P3_U3158 = ~n25637 | ~n25636;
  assign n25640 = ~n26375 & ~n25725;
  assign n25639 = ~n25666 & ~n25638;
  assign n25650 = ~n25640 & ~n25639;
  assign n25641 = ~n25706 | ~n26165;
  assign n25902 = ~P3_REG3_REG_8__SCAN_IN | ~P3_U3151;
  assign n25648 = ~n25641 | ~n25902;
  assign n25644 = n25643 ^ n25642;
  assign n25646 = ~n25644 | ~n25732;
  assign n25645 = ~n25734 | ~n26101;
  assign n25647 = ~n25646 | ~n25645;
  assign n25649 = ~n25648 & ~n25647;
  assign P3_U3161 = ~n25650 | ~n25649;
  assign n25653 = ~n25706 | ~n26287;
  assign n25652 = ~n25708 | ~n25651;
  assign n25658 = ~n25653 | ~n25652;
  assign n25720 = ~P3_STATE_REG_SCAN_IN | ~n25654;
  assign n25656 = ~P3_REG3_REG_1__SCAN_IN | ~n25720;
  assign n25655 = ~n25728 | ~n26286;
  assign n25657 = ~n25656 | ~n25655;
  assign n25665 = ~n25658 & ~n25657;
  assign n25662 = n25660 | n25659;
  assign n25663 = ~n25662 | ~n25661;
  assign n25664 = ~n25663 | ~n25732;
  assign P3_U3162 = ~n25665 | ~n25664;
  assign n25668 = ~n25666 & ~n26138;
  assign n25837 = ~n25667 & ~P3_STATE_REG_SCAN_IN;
  assign n25681 = ~n25668 & ~n25837;
  assign n25670 = ~n25706 | ~n26229;
  assign n25669 = ~n25708 | ~n26174;
  assign n25679 = ~n25670 | ~n25669;
  assign n25674 = n25672 | n25671;
  assign n25675 = ~n25674 | ~n25673;
  assign n25677 = ~n25675 | ~n25732;
  assign n25676 = ~n25734 | ~n26175;
  assign n25678 = ~n25677 | ~n25676;
  assign n25680 = ~n25679 & ~n25678;
  assign P3_U3167 = ~n25681 | ~n25680;
  assign n25682 = ~n25708 | ~n26316;
  assign n25686 = ~n25683 | ~n25682;
  assign n25685 = ~n25684 & ~n26305;
  assign n25688 = ~n25686 & ~n25685;
  assign n25687 = ~P3_REG3_REG_0__SCAN_IN | ~n25720;
  assign P3_U3172 = ~n25688 | ~n25687;
  assign n25690 = ~n25724 & ~n25689;
  assign n25967 = P3_U3151 & P3_REG3_REG_11__SCAN_IN;
  assign n25705 = ~n25690 & ~n25967;
  assign n25694 = ~n25691 | ~n25708;
  assign n25693 = ~n25728 | ~n25692;
  assign n25703 = ~n25694 | ~n25693;
  assign n25696 = n25695 ^ ~n26059;
  assign n25698 = n25697 ^ ~n25696;
  assign n25701 = ~n25698 | ~n25732;
  assign n25700 = ~n25734 | ~n25699;
  assign n25702 = ~n25701 | ~n25700;
  assign n25704 = ~n25703 & ~n25702;
  assign P3_U3176 = ~n25705 | ~n25704;
  assign n25709 = ~n25708 | ~n25707;
  assign n25719 = ~n25710 | ~n25709;
  assign n25713 = n25712 | n25711;
  assign n25715 = ~n25714 | ~n25713;
  assign n25717 = ~n25715 | ~n25732;
  assign n25716 = ~n25728 | ~n26252;
  assign n25718 = ~n25717 | ~n25716;
  assign n25722 = ~n25719 & ~n25718;
  assign n25721 = ~P3_REG3_REG_2__SCAN_IN | ~n25720;
  assign P3_U3177 = ~n25722 | ~n25721;
  assign n25727 = ~n25724 & ~n25723;
  assign n25726 = ~n25725 & ~n26359;
  assign n25740 = ~n25727 & ~n25726;
  assign n25729 = ~n25728 | ~n26165;
  assign n25858 = ~P3_REG3_REG_6__SCAN_IN | ~P3_U3151;
  assign n25738 = ~n25729 | ~n25858;
  assign n25733 = n25731 ^ n25730;
  assign n25736 = ~n25733 | ~n25732;
  assign n25735 = ~n25734 | ~n26151;
  assign n25737 = ~n25736 | ~n25735;
  assign n25739 = ~n25738 & ~n25737;
  assign P3_U3179 = ~n25740 | ~n25739;
  assign n25753 = ~n25771;
  assign n25743 = ~n25753 | ~n25742;
  assign n25745 = ~n26027 | ~n25743;
  assign n25744 = ~n26033 | ~P3_ADDR_REG_0__SCAN_IN;
  assign n25749 = ~n25745 | ~n25744;
  assign n26010 = ~n26031;
  assign n25747 = ~n25771 & ~n25746;
  assign n25748 = ~n26010 & ~n25747;
  assign n25760 = ~n25749 & ~n25748;
  assign n25752 = ~n25751 | ~n25750;
  assign n25754 = ~n25753 | ~n25752;
  assign n25756 = ~n25754 | ~n26013;
  assign n25755 = ~P3_REG3_REG_0__SCAN_IN | ~P3_U3151;
  assign n25758 = ~n25756 | ~n25755;
  assign n25757 = n25894 & P3_IR_REG_0__SCAN_IN;
  assign n25759 = ~n25758 & ~n25757;
  assign P3_U3182 = ~n25760 | ~n25759;
  assign n25762 = ~P3_ADDR_REG_1__SCAN_IN | ~n26033;
  assign n25761 = ~P3_REG3_REG_1__SCAN_IN | ~P3_U3151;
  assign n25770 = ~n25762 | ~n25761;
  assign n25764 = n25763 ^ ~P3_REG2_REG_1__SCAN_IN;
  assign n25768 = ~n25764 | ~n26031;
  assign n25766 = n25765 ^ P3_REG1_REG_1__SCAN_IN;
  assign n25767 = ~n26027 | ~n25766;
  assign n25769 = ~n25768 | ~n25767;
  assign n25777 = ~n25770 & ~n25769;
  assign n25772 = n25771 ^ n13224;
  assign n26044 = ~n26013;
  assign n25775 = ~n25772 & ~n26044;
  assign n25774 = ~n26037 & ~n25773;
  assign n25776 = ~n25775 & ~n25774;
  assign P3_U3183 = ~n25777 | ~n25776;
  assign n25788 = ~n26037 & ~n25778;
  assign n25781 = n25780 ^ ~n25779;
  assign n25786 = ~n26027 | ~n25781;
  assign n25784 = n25783 ^ ~n25782;
  assign n25785 = ~n25784 | ~n26031;
  assign n25787 = ~n25786 | ~n25785;
  assign n25797 = ~n25788 & ~n25787;
  assign n25791 = n25789 ^ n25790;
  assign n25795 = ~n25791 & ~n26044;
  assign n25793 = ~P3_ADDR_REG_2__SCAN_IN | ~n26033;
  assign n25792 = ~P3_REG3_REG_2__SCAN_IN | ~P3_U3151;
  assign n25794 = ~n25793 | ~n25792;
  assign n25796 = ~n25795 & ~n25794;
  assign P3_U3184 = ~n25797 | ~n25796;
  assign n25799 = n26033 & P3_ADDR_REG_3__SCAN_IN;
  assign n25817 = ~n25799 & ~n25798;
  assign n25801 = n25800 ^ ~P3_REG2_REG_3__SCAN_IN;
  assign n25805 = ~n25801 | ~n26031;
  assign n25803 = n25802 ^ ~P3_REG1_REG_3__SCAN_IN;
  assign n25804 = ~n26027 | ~n25803;
  assign n25815 = ~n25805 | ~n25804;
  assign n25808 = n25807 | n25806;
  assign n25810 = ~n25809 | ~n25808;
  assign n25813 = ~n25810 | ~n26013;
  assign n25812 = ~n25894 | ~n25811;
  assign n25814 = ~n25813 | ~n25812;
  assign n25816 = ~n25815 & ~n25814;
  assign P3_U3185 = ~n25817 | ~n25816;
  assign n25818 = ~n26033 | ~P3_ADDR_REG_4__SCAN_IN;
  assign n25828 = ~n25819 | ~n25818;
  assign n25826 = ~n26027 | ~n25821;
  assign n25824 = n25823 ^ ~n25822;
  assign n25825 = ~n25824 | ~n26031;
  assign n25827 = ~n25826 | ~n25825;
  assign n25836 = ~n25828 & ~n25827;
  assign n25831 = n25829 ^ n25830;
  assign n25834 = ~n25831 & ~n26044;
  assign n25833 = ~n26037 & ~n25832;
  assign n25835 = ~n25834 & ~n25833;
  assign P3_U3186 = ~n25836 | ~n25835;
  assign n25838 = n26033 & P3_ADDR_REG_5__SCAN_IN;
  assign n25856 = ~n25838 & ~n25837;
  assign n25840 = n25839 ^ ~P3_REG1_REG_5__SCAN_IN;
  assign n25844 = ~n25840 | ~n26027;
  assign n25842 = n25841 ^ ~P3_REG2_REG_5__SCAN_IN;
  assign n25843 = ~n25842 | ~n26031;
  assign n25854 = ~n25844 | ~n25843;
  assign n25847 = ~n14236 & ~n25846;
  assign n25849 = n25848 ^ ~n25847;
  assign n25852 = ~n25849 | ~n26013;
  assign n25851 = ~n25894 | ~n25850;
  assign n25853 = ~n25852 | ~n25851;
  assign n25855 = ~n25854 & ~n25853;
  assign P3_U3187 = ~n25856 | ~n25855;
  assign n25857 = ~n26033 | ~P3_ADDR_REG_6__SCAN_IN;
  assign n25868 = ~n25858 | ~n25857;
  assign n25861 = n25860 ^ ~n25859;
  assign n25866 = ~n25861 | ~n26027;
  assign n25864 = n25863 ^ ~n25862;
  assign n25865 = ~n25864 | ~n26031;
  assign n25867 = ~n25866 | ~n25865;
  assign n25879 = ~n25868 & ~n25867;
  assign n25871 = ~n25869;
  assign n25872 = ~n25871 & ~n25870;
  assign n25874 = n25873 ^ ~n25872;
  assign n25877 = ~n25874 & ~n26044;
  assign n25876 = ~n26037 & ~n25875;
  assign n25878 = ~n25877 & ~n25876;
  assign P3_U3188 = ~n25879 | ~n25878;
  assign n25881 = n26033 & P3_ADDR_REG_7__SCAN_IN;
  assign n25900 = ~n25881 & ~n25880;
  assign n25883 = n25882 ^ ~P3_REG2_REG_7__SCAN_IN;
  assign n25887 = ~n25883 | ~n26031;
  assign n25885 = n25884 ^ ~P3_REG1_REG_7__SCAN_IN;
  assign n25886 = ~n25885 | ~n26027;
  assign n25898 = ~n25887 | ~n25886;
  assign n25890 = n25889 | n25888;
  assign n25892 = ~n25891 | ~n25890;
  assign n25896 = ~n25892 | ~n26013;
  assign n25895 = ~n25894 | ~n25893;
  assign n25897 = ~n25896 | ~n25895;
  assign n25899 = ~n25898 & ~n25897;
  assign P3_U3189 = ~n25900 | ~n25899;
  assign n25901 = ~n26033 | ~P3_ADDR_REG_8__SCAN_IN;
  assign n25912 = ~n25902 | ~n25901;
  assign n25905 = n25904 ^ ~n25903;
  assign n25910 = ~n25905 | ~n26027;
  assign n25908 = n25907 ^ ~n25906;
  assign n25909 = ~n25908 | ~n26031;
  assign n25911 = ~n25910 | ~n25909;
  assign n25920 = ~n25912 & ~n25911;
  assign n25915 = n25913 ^ n25914;
  assign n25918 = ~n25915 & ~n26044;
  assign n25917 = ~n26037 & ~n25916;
  assign n25919 = ~n25918 & ~n25917;
  assign P3_U3190 = ~n25920 | ~n25919;
  assign n25922 = n25921 ^ ~P3_REG2_REG_9__SCAN_IN;
  assign n25941 = ~n25922 | ~n26031;
  assign n25925 = ~n26037 & ~n25923;
  assign n25927 = ~n25925 & ~n25924;
  assign n25926 = ~n26033 | ~P3_ADDR_REG_9__SCAN_IN;
  assign n25939 = ~n25927 | ~n25926;
  assign n25929 = n25928 ^ ~P3_REG1_REG_9__SCAN_IN;
  assign n25937 = ~n25929 | ~n26027;
  assign n25932 = ~n25930;
  assign n25933 = ~n25932 & ~n25931;
  assign n25935 = n25934 ^ ~n25933;
  assign n25936 = ~n25935 | ~n26013;
  assign n25938 = ~n25937 | ~n25936;
  assign n25940 = ~n25939 & ~n25938;
  assign P3_U3191 = ~n25941 | ~n25940;
  assign n25944 = n25943 ^ ~n25942;
  assign n25963 = ~n25944 | ~n26027;
  assign n25947 = n25946 ^ n25945;
  assign n25961 = ~n26010 & ~n25947;
  assign n25951 = n25949 | n25948;
  assign n25952 = ~n25951 | ~n25950;
  assign n25959 = ~n25952 | ~n26013;
  assign n25953 = ~n26033 | ~P3_ADDR_REG_10__SCAN_IN;
  assign n25957 = ~n25954 | ~n25953;
  assign n25956 = ~n26037 & ~n25955;
  assign n25958 = ~n25957 & ~n25956;
  assign n25960 = ~n25959 | ~n25958;
  assign n25962 = ~n25961 & ~n25960;
  assign P3_U3192 = ~n25963 | ~n25962;
  assign n25965 = n25964 ^ ~P3_REG2_REG_11__SCAN_IN;
  assign n25981 = ~n25965 | ~n26031;
  assign n25968 = ~n26037 & ~n25966;
  assign n25970 = ~n25968 & ~n25967;
  assign n25969 = ~n26033 | ~P3_ADDR_REG_11__SCAN_IN;
  assign n25979 = ~n25970 | ~n25969;
  assign n25972 = n25971 ^ ~P3_REG1_REG_11__SCAN_IN;
  assign n25977 = ~n25972 | ~n26027;
  assign n25975 = n25974 ^ ~n25973;
  assign n25976 = ~n25975 | ~n26013;
  assign n25978 = ~n25977 | ~n25976;
  assign n25980 = ~n25979 & ~n25978;
  assign P3_U3193 = ~n25981 | ~n25980;
  assign n25984 = n25983 ^ ~n25982;
  assign n26004 = ~n25984 | ~n26031;
  assign n25987 = n25986 ^ ~n25985;
  assign n25994 = ~n25987 | ~n26027;
  assign n25992 = ~n26037 & ~n25988;
  assign n25989 = ~n26033 | ~P3_ADDR_REG_12__SCAN_IN;
  assign n25991 = ~n25990 | ~n25989;
  assign n25993 = ~n25992 & ~n25991;
  assign n26002 = ~n25994 | ~n25993;
  assign n26000 = ~n25995;
  assign n25998 = ~n25997 | ~n25996;
  assign n25999 = ~n25998 | ~n26013;
  assign n26001 = ~n26000 & ~n25999;
  assign n26003 = ~n26002 & ~n26001;
  assign P3_U3194 = ~n26004 | ~n26003;
  assign n26006 = n26005 ^ ~P3_REG1_REG_13__SCAN_IN;
  assign n26025 = ~n26006 | ~n26027;
  assign n26009 = n26008 ^ ~n26007;
  assign n26023 = ~n26010 & ~n26009;
  assign n26014 = n26012 ^ ~n26011;
  assign n26021 = ~n26014 | ~n26013;
  assign n26015 = ~n26033 | ~P3_ADDR_REG_13__SCAN_IN;
  assign n26019 = ~n26016 | ~n26015;
  assign n26018 = ~n26037 & ~n26017;
  assign n26020 = ~n26019 & ~n26018;
  assign n26022 = ~n26021 | ~n26020;
  assign n26024 = ~n26023 & ~n26022;
  assign P3_U3195 = ~n26025 | ~n26024;
  assign n26051 = ~n26028 | ~n26027;
  assign n26032 = n26030 ^ ~n26029;
  assign n26041 = ~n26032 | ~n26031;
  assign n26034 = ~n26033 | ~P3_ADDR_REG_14__SCAN_IN;
  assign n26039 = ~n26035 | ~n26034;
  assign n26038 = ~n26037 & ~n26036;
  assign n26040 = ~n26039 & ~n26038;
  assign n26049 = ~n26041 | ~n26040;
  assign n26045 = ~n26043 & ~n26042;
  assign n26047 = ~n26045 & ~n26044;
  assign n26048 = n26047 & n26046;
  assign n26050 = ~n26049 & ~n26048;
  assign P3_U3196 = ~n26051 | ~n26050;
  assign n26392 = n26052 ^ ~n14741;
  assign n26056 = ~n26392;
  assign n26064 = ~n26056 | ~n26228;
  assign n26055 = n26054 ^ ~n26053;
  assign n26058 = ~n26055 | ~n26280;
  assign n26057 = ~n26056 | ~n26282;
  assign n26063 = ~n26058 | ~n26057;
  assign n26061 = ~n26059 | ~n18385;
  assign n26060 = ~n26288 | ~n26116;
  assign n26062 = ~n26061 | ~n26060;
  assign n26397 = ~n26063 & ~n26062;
  assign n26065 = ~n26064 | ~n26397;
  assign n26073 = ~n26065 | ~n20481;
  assign n26071 = ~n26393 & ~n26224;
  assign n26069 = n20481 | n26066;
  assign n26068 = ~n26152 | ~n26067;
  assign n26070 = ~n26069 | ~n26068;
  assign n26072 = ~n26071 & ~n26070;
  assign P3_U3223 = ~n26073 | ~n26072;
  assign n26077 = ~n26074 | ~n26075;
  assign n26079 = ~n26077 | ~n26076;
  assign n26382 = n26079 ^ ~n26078;
  assign n26080 = ~n26382;
  assign n26091 = ~n26080 | ~n26228;
  assign n26084 = ~n26080 | ~n26282;
  assign n26082 = n13382 ^ ~n26081;
  assign n26083 = ~n26082 | ~n26280;
  assign n26090 = ~n26084 | ~n26083;
  assign n26088 = ~n26085 | ~n18385;
  assign n26087 = ~n26288 | ~n26086;
  assign n26089 = ~n26088 | ~n26087;
  assign n26387 = ~n26090 & ~n26089;
  assign n26092 = ~n26091 | ~n26387;
  assign n26100 = ~n26092 | ~n20481;
  assign n26098 = ~n26224 & ~n26383;
  assign n26096 = n20481 | n26093;
  assign n26095 = ~n26152 | ~n26094;
  assign n26097 = ~n26096 | ~n26095;
  assign n26099 = ~n26098 & ~n26097;
  assign P3_U3224 = ~n26100 | ~n26099;
  assign n26103 = ~n26270 | ~P3_REG2_REG_8__SCAN_IN;
  assign n26102 = ~n26152 | ~n26101;
  assign n26105 = ~n26103 | ~n26102;
  assign n26104 = ~n26224 & ~n26375;
  assign n26124 = ~n26105 & ~n26104;
  assign n26108 = ~n26074 | ~n26106;
  assign n26110 = ~n26108 | ~n26107;
  assign n26374 = n26110 ^ ~n26109;
  assign n26113 = ~n26374;
  assign n26121 = ~n26113 | ~n26228;
  assign n26115 = ~n26112 | ~n26280;
  assign n26114 = ~n26113 | ~n26282;
  assign n26120 = ~n26115 | ~n26114;
  assign n26118 = ~n26165 | ~n26288;
  assign n26117 = ~n18385 | ~n26116;
  assign n26119 = ~n26118 | ~n26117;
  assign n26379 = ~n26120 & ~n26119;
  assign n26122 = ~n26121 | ~n26379;
  assign n26123 = ~n26122 | ~n20481;
  assign P3_U3225 = ~n26124 | ~n26123;
  assign n26136 = ~n26126 & ~n26125;
  assign n26128 = ~n13906 & ~n26127;
  assign n26131 = ~n26129 & ~n26128;
  assign n26134 = ~n26131 | ~n26130;
  assign n26366 = n26074 ^ ~n13906;
  assign n26132 = ~n26366;
  assign n26133 = ~n26132 | ~n26282;
  assign n26135 = ~n26134 | ~n26133;
  assign n26139 = ~n26138 & ~n26137;
  assign n26371 = ~n26140 & ~n26139;
  assign n26142 = ~n26152 | ~n26141;
  assign n26144 = ~n26371 | ~n26142;
  assign n26143 = ~n26249 & ~n26366;
  assign n26145 = ~n26144 & ~n26143;
  assign n26147 = ~n26270 & ~n26145;
  assign n26146 = ~n26224 & ~n26367;
  assign n26149 = ~n26147 & ~n26146;
  assign n26148 = ~P3_REG2_REG_7__SCAN_IN | ~n26270;
  assign P3_U3226 = ~n26149 | ~n26148;
  assign n26154 = ~n26297 | ~n26150;
  assign n26153 = ~n26152 | ~n26151;
  assign n26157 = ~n26154 | ~n26153;
  assign n26156 = ~n20481 & ~n26155;
  assign n26173 = ~n26157 & ~n26156;
  assign n26358 = n26158 ^ n26160;
  assign n26159 = ~n26358;
  assign n26170 = ~n26159 | ~n26228;
  assign n26164 = ~n26159 | ~n26282;
  assign n26162 = n26161 ^ n26160;
  assign n26163 = ~n26162 | ~n26280;
  assign n26169 = ~n26164 | ~n26163;
  assign n26167 = ~n26165 | ~n18385;
  assign n26166 = ~n26288 | ~n26205;
  assign n26168 = ~n26167 | ~n26166;
  assign n26363 = ~n26169 & ~n26168;
  assign n26171 = ~n26170 | ~n26363;
  assign n26172 = ~n26171 | ~n20481;
  assign P3_U3227 = ~n26173 | ~n26172;
  assign n26177 = ~n26297 | ~n26174;
  assign n26176 = ~n26152 | ~n26175;
  assign n26180 = ~n26177 | ~n26176;
  assign n26179 = ~n20481 & ~n26178;
  assign n26197 = ~n26180 & ~n26179;
  assign n26350 = n26182 ^ ~n26181;
  assign n26186 = ~n26350;
  assign n26194 = ~n26186 | ~n26228;
  assign n26185 = n26184 ^ ~n26183;
  assign n26188 = ~n26185 | ~n26280;
  assign n26187 = ~n26186 | ~n26282;
  assign n26193 = ~n26188 | ~n26187;
  assign n26191 = ~n18385 | ~n26189;
  assign n26190 = ~n26288 | ~n26229;
  assign n26192 = ~n26191 | ~n26190;
  assign n26355 = ~n26193 & ~n26192;
  assign n26195 = ~n26194 | ~n26355;
  assign n26196 = ~n26195 | ~n20481;
  assign P3_U3228 = ~n26197 | ~n26196;
  assign n26342 = n26199 ^ ~n26198;
  assign n26202 = ~n26342;
  assign n26210 = ~n26202 | ~n26228;
  assign n26201 = n26200 ^ ~n14555;
  assign n26204 = ~n26201 | ~n26280;
  assign n26203 = ~n26202 | ~n26282;
  assign n26209 = ~n26204 | ~n26203;
  assign n26207 = ~n18385 | ~n26205;
  assign n26206 = ~n26288 | ~n26252;
  assign n26208 = ~n26207 | ~n26206;
  assign n26347 = ~n26209 & ~n26208;
  assign n26211 = ~n26210 | ~n26347;
  assign n26221 = ~n26211 | ~n20481;
  assign n26215 = ~n26297 | ~n26212;
  assign n26214 = ~n26152 | ~n26213;
  assign n26219 = ~n26215 | ~n26214;
  assign n26218 = ~n20481 & ~n26216;
  assign n26220 = ~n26219 & ~n26218;
  assign P3_U3229 = ~n26221 | ~n26220;
  assign n26223 = ~P3_REG2_REG_3__SCAN_IN | ~n26270;
  assign n26222 = ~n26152 | ~n16443;
  assign n26226 = ~n26223 | ~n26222;
  assign n26225 = ~n26224 & ~n26335;
  assign n26244 = ~n26226 & ~n26225;
  assign n26334 = n26227 ^ ~n26233;
  assign n26236 = ~n26334;
  assign n26241 = ~n26236 | ~n26228;
  assign n26231 = ~n18385 | ~n26229;
  assign n26230 = ~n26288 | ~n26286;
  assign n26240 = ~n26231 | ~n26230;
  assign n26235 = n26234 ^ ~n26233;
  assign n26238 = ~n26235 | ~n26280;
  assign n26237 = ~n26236 | ~n26282;
  assign n26239 = ~n26238 | ~n26237;
  assign n26339 = ~n26240 & ~n26239;
  assign n26242 = ~n26241 | ~n26339;
  assign n26243 = ~n26242 | ~n20481;
  assign P3_U3230 = ~n26244 | ~n26243;
  assign n26247 = ~n26152 | ~P3_REG3_REG_2__SCAN_IN;
  assign n26328 = ~n26245 & ~n20673;
  assign n26246 = ~n26328 | ~n26278;
  assign n26251 = ~n26247 | ~n26246;
  assign n26327 = n26248 ^ ~n26258;
  assign n26250 = ~n26327 & ~n26249;
  assign n26266 = ~n26251 & ~n26250;
  assign n26254 = ~n18385 | ~n26252;
  assign n26265 = ~n26254 | ~n26253;
  assign n26257 = ~n26255;
  assign n26259 = ~n26257 | ~n26256;
  assign n26260 = n26258 ^ ~n26259;
  assign n26263 = ~n26260 | ~n26280;
  assign n26261 = ~n26327;
  assign n26262 = ~n26261 | ~n26282;
  assign n26264 = ~n26263 | ~n26262;
  assign n26331 = ~n26265 & ~n26264;
  assign n26267 = ~n26266 | ~n26331;
  assign n26269 = ~n20481 | ~n26267;
  assign n26268 = ~n26270 | ~P3_REG2_REG_2__SCAN_IN;
  assign P3_U3231 = ~n26269 | ~n26268;
  assign n26272 = ~n26152 | ~P3_REG3_REG_1__SCAN_IN;
  assign n26271 = ~n26270 | ~P3_REG2_REG_1__SCAN_IN;
  assign n26276 = ~n26272 | ~n26271;
  assign n26320 = n26273 ^ ~n19273;
  assign n26275 = ~n26320 & ~n26274;
  assign n26296 = ~n26276 & ~n26275;
  assign n26321 = ~n26277 & ~n20673;
  assign n26293 = ~n26321 | ~n26278;
  assign n26281 = n19273 ^ ~n26279;
  assign n26285 = ~n26281 | ~n26280;
  assign n26283 = ~n26320;
  assign n26284 = ~n26283 | ~n26282;
  assign n26292 = ~n26285 | ~n26284;
  assign n26290 = ~n18385 | ~n26286;
  assign n26289 = ~n26288 | ~n26287;
  assign n26291 = ~n26290 | ~n26289;
  assign n26324 = ~n26292 & ~n26291;
  assign n26294 = ~n26293 | ~n26324;
  assign n26295 = ~n26294 | ~n20481;
  assign P3_U3232 = ~n26296 | ~n26295;
  assign n26299 = ~n26297 | ~n26316;
  assign n26298 = ~n26152 | ~P3_REG3_REG_0__SCAN_IN;
  assign n26302 = ~n26299 | ~n26298;
  assign n26301 = ~n26300 & ~n20481;
  assign n26309 = ~n26302 & ~n26301;
  assign n26304 = n26303 | n26315;
  assign n26307 = n26305 | n26304;
  assign n26317 = ~n26307 | ~n26306;
  assign n26308 = ~n26317 | ~n20481;
  assign P3_U3233 = ~n26309 | ~n26308;
  assign n26314 = ~n26311 & ~n26310;
  assign n26313 = ~n26312 & ~P3_D_REG_1__SCAN_IN;
  assign P3_U3377 = ~n26314 & ~n26313;
  assign n26319 = ~P3_REG0_REG_0__SCAN_IN | ~n26390;
  assign n26401 = n26317 | n14879;
  assign n26318 = ~n26398 | ~n26401;
  assign P3_U3390 = ~n26319 | ~n26318;
  assign n26326 = ~P3_REG0_REG_1__SCAN_IN | ~n26390;
  assign n26322 = ~n26320 & ~n26391;
  assign n26323 = ~n26322 & ~n26321;
  assign n26404 = ~n26324 | ~n26323;
  assign n26325 = ~n26398 | ~n26404;
  assign P3_U3393 = ~n26326 | ~n26325;
  assign n26333 = ~P3_REG0_REG_2__SCAN_IN | ~n26390;
  assign n26329 = ~n26327 & ~n26391;
  assign n26330 = ~n26329 & ~n26328;
  assign n26407 = ~n26331 | ~n26330;
  assign n26332 = ~n26398 | ~n26407;
  assign P3_U3396 = ~n26333 | ~n26332;
  assign n26341 = ~P3_REG0_REG_3__SCAN_IN | ~n26390;
  assign n26337 = ~n26334 & ~n26391;
  assign n26336 = ~n26335 & ~n20673;
  assign n26338 = ~n26337 & ~n26336;
  assign n26410 = ~n26339 | ~n26338;
  assign n26340 = ~n26398 | ~n26410;
  assign P3_U3399 = ~n26341 | ~n26340;
  assign n26349 = ~P3_REG0_REG_4__SCAN_IN | ~n26390;
  assign n26345 = ~n26342 & ~n26391;
  assign n26344 = ~n26343 & ~n20673;
  assign n26346 = ~n26345 & ~n26344;
  assign n26413 = ~n26347 | ~n26346;
  assign n26348 = ~n26398 | ~n26413;
  assign P3_U3402 = ~n26349 | ~n26348;
  assign n26357 = ~P3_REG0_REG_5__SCAN_IN | ~n26390;
  assign n26353 = ~n26350 & ~n26391;
  assign n26352 = ~n26351 & ~n20673;
  assign n26354 = ~n26353 & ~n26352;
  assign n26416 = ~n26355 | ~n26354;
  assign n26356 = ~n26398 | ~n26416;
  assign P3_U3405 = ~n26357 | ~n26356;
  assign n26365 = ~P3_REG0_REG_6__SCAN_IN | ~n26390;
  assign n26361 = ~n26358 & ~n26391;
  assign n26360 = ~n26359 & ~n20673;
  assign n26362 = ~n26361 & ~n26360;
  assign n26419 = ~n26363 | ~n26362;
  assign n26364 = ~n26398 | ~n26419;
  assign P3_U3408 = ~n26365 | ~n26364;
  assign n26373 = ~P3_REG0_REG_7__SCAN_IN | ~n26390;
  assign n26369 = ~n26366 & ~n26391;
  assign n26368 = ~n26367 & ~n20673;
  assign n26370 = ~n26369 & ~n26368;
  assign n26422 = ~n26371 | ~n26370;
  assign n26372 = ~n26398 | ~n26422;
  assign P3_U3411 = ~n26373 | ~n26372;
  assign n26381 = ~P3_REG0_REG_8__SCAN_IN | ~n26390;
  assign n26377 = ~n26374 & ~n26391;
  assign n26376 = ~n26375 & ~n20673;
  assign n26378 = ~n26377 & ~n26376;
  assign n26425 = ~n26379 | ~n26378;
  assign n26380 = ~n26398 | ~n26425;
  assign P3_U3414 = ~n26381 | ~n26380;
  assign n26389 = ~P3_REG0_REG_9__SCAN_IN | ~n26390;
  assign n26385 = ~n26382 & ~n26391;
  assign n26384 = ~n26383 & ~n20673;
  assign n26386 = ~n26385 & ~n26384;
  assign n26428 = ~n26387 | ~n26386;
  assign n26388 = ~n26398 | ~n26428;
  assign P3_U3417 = ~n26389 | ~n26388;
  assign n26400 = ~P3_REG0_REG_10__SCAN_IN | ~n26390;
  assign n26395 = ~n26392 & ~n26391;
  assign n26394 = ~n26393 & ~n20673;
  assign n26396 = ~n26395 & ~n26394;
  assign n26432 = ~n26397 | ~n26396;
  assign n26399 = ~n26398 | ~n26432;
  assign P3_U3420 = ~n26400 | ~n26399;
  assign n26403 = ~P3_REG1_REG_0__SCAN_IN | ~n26431;
  assign n26402 = ~n26433 | ~n26401;
  assign P3_U3459 = ~n26403 | ~n26402;
  assign n26406 = ~P3_REG1_REG_1__SCAN_IN | ~n26431;
  assign n26405 = ~n26433 | ~n26404;
  assign P3_U3460 = ~n26406 | ~n26405;
  assign n26409 = ~P3_REG1_REG_2__SCAN_IN | ~n26431;
  assign n26408 = ~n26433 | ~n26407;
  assign P3_U3461 = ~n26409 | ~n26408;
  assign n26412 = ~P3_REG1_REG_3__SCAN_IN | ~n26431;
  assign n26411 = ~n26433 | ~n26410;
  assign P3_U3462 = ~n26412 | ~n26411;
  assign n26415 = ~P3_REG1_REG_4__SCAN_IN | ~n26431;
  assign n26414 = ~n26433 | ~n26413;
  assign P3_U3463 = ~n26415 | ~n26414;
  assign n26418 = ~P3_REG1_REG_5__SCAN_IN | ~n26431;
  assign n26417 = ~n26433 | ~n26416;
  assign P3_U3464 = ~n26418 | ~n26417;
  assign n26421 = ~P3_REG1_REG_6__SCAN_IN | ~n26431;
  assign n26420 = ~n26433 | ~n26419;
  assign P3_U3465 = ~n26421 | ~n26420;
  assign n26424 = ~P3_REG1_REG_7__SCAN_IN | ~n26431;
  assign n26423 = ~n26433 | ~n26422;
  assign P3_U3466 = ~n26424 | ~n26423;
  assign n26427 = ~P3_REG1_REG_8__SCAN_IN | ~n26431;
  assign n26426 = ~n26433 | ~n26425;
  assign P3_U3467 = ~n26427 | ~n26426;
  assign n26430 = ~P3_REG1_REG_9__SCAN_IN | ~n26431;
  assign n26429 = ~n26433 | ~n26428;
  assign P3_U3468 = ~n26430 | ~n26429;
  assign n26435 = ~P3_REG1_REG_10__SCAN_IN | ~n26431;
  assign n26434 = ~n26433 | ~n26432;
  assign P3_U3469 = ~n26435 | ~n26434;
  assign n26438 = ~P3_DATAO_REG_25__SCAN_IN | ~n26454;
  assign n26437 = ~P3_U3897 | ~n26436;
  assign P3_U3516 = ~n26438 | ~n26437;
  assign n26441 = ~P3_DATAO_REG_26__SCAN_IN | ~n26454;
  assign n26440 = ~P3_U3897 | ~n26439;
  assign P3_U3517 = ~n26441 | ~n26440;
  assign n26444 = ~P3_DATAO_REG_27__SCAN_IN | ~n26454;
  assign n26443 = ~P3_U3897 | ~n26442;
  assign P3_U3518 = ~n26444 | ~n26443;
  assign n26447 = ~P3_DATAO_REG_28__SCAN_IN | ~n26454;
  assign n26446 = ~P3_U3897 | ~n26445;
  assign P3_U3519 = ~n26447 | ~n26446;
  assign n26450 = ~P3_DATAO_REG_29__SCAN_IN | ~n26454;
  assign n26449 = ~P3_U3897 | ~n26448;
  assign P3_U3520 = ~n26450 | ~n26449;
  assign n26453 = ~P3_DATAO_REG_30__SCAN_IN | ~n26454;
  assign n26452 = ~P3_U3897 | ~n26451;
  assign P3_U3521 = ~n26453 | ~n26452;
  assign n26457 = ~P3_DATAO_REG_31__SCAN_IN | ~n26454;
  assign n26456 = ~P3_U3897 | ~n26455;
  assign P3_U3522 = ~n26457 | ~n26456;
  assign n13665 = n18154 & n13239;
  assign n20481 = ~n26270;
endmodule


