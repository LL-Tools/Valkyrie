

module b17_C_AntiSAT_k_128_6 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14207, n14208, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148;

  AOI21_X1 U11080 ( .B1(n14090), .B2(n14088), .A(n14089), .ZN(n14477) );
  OAI21_X1 U11081 ( .B1(n12536), .B2(n19366), .A(n9799), .ZN(n10116) );
  CLKBUF_X1 U11082 ( .A(n12508), .Z(n12538) );
  OR2_X1 U11083 ( .A1(n16054), .A2(n14187), .ZN(n16045) );
  XNOR2_X1 U11084 ( .A(n14400), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14398) );
  CLKBUF_X2 U11085 ( .A(n12139), .Z(n9668) );
  AND2_X1 U11086 ( .A1(n12076), .A2(n15636), .ZN(n12150) );
  INV_X1 U11087 ( .A(n11236), .ZN(n11235) );
  CLKBUF_X1 U11088 ( .A(n11212), .Z(n13178) );
  INV_X1 U11090 ( .A(n9695), .ZN(n13834) );
  CLKBUF_X2 U11091 ( .A(n10586), .Z(n13971) );
  CLKBUF_X2 U11093 ( .A(n11111), .Z(n11627) );
  CLKBUF_X2 U11094 ( .A(n12842), .Z(n15814) );
  CLKBUF_X3 U11095 ( .A(n15669), .Z(n9649) );
  CLKBUF_X3 U11096 ( .A(n12838), .Z(n9644) );
  CLKBUF_X1 U11097 ( .A(n12842), .Z(n9642) );
  INV_X2 U11098 ( .A(n15827), .ZN(n17247) );
  CLKBUF_X1 U11099 ( .A(n10394), .Z(n19411) );
  NAND2_X1 U11100 ( .A1(n10963), .A2(n10964), .ZN(n20285) );
  INV_X1 U11101 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18901) );
  NAND2_X1 U11102 ( .A1(n10394), .A2(n10584), .ZN(n12243) );
  INV_X1 U11103 ( .A(n11845), .ZN(n11139) );
  INV_X1 U11104 ( .A(n11031), .ZN(n11814) );
  BUF_X2 U11105 ( .A(n11849), .Z(n11904) );
  AND2_X1 U11106 ( .A1(n10916), .A2(n10911), .ZN(n11003) );
  AND2_X1 U11107 ( .A1(n10916), .A2(n13177), .ZN(n11021) );
  AND2_X1 U11108 ( .A1(n10911), .A2(n10912), .ZN(n10977) );
  AND2_X1 U11109 ( .A1(n10914), .A2(n10902), .ZN(n10903) );
  AND2_X1 U11110 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U11111 ( .A1(n10908), .A2(n13177), .ZN(n11810) );
  AND2_X1 U11112 ( .A1(n13056), .A2(n15646), .ZN(n13875) );
  CLKBUF_X1 U11113 ( .A(n20291), .Z(n9636) );
  NOR2_X1 U11114 ( .A1(n20241), .A2(n20243), .ZN(n20291) );
  CLKBUF_X1 U11115 ( .A(n20290), .Z(n9637) );
  NOR2_X1 U11116 ( .A1(n20243), .A2(n20242), .ZN(n20290) );
  INV_X1 U11118 ( .A(n10952), .ZN(n11839) );
  AND2_X2 U11119 ( .A1(n10916), .A2(n10915), .ZN(n11130) );
  AND3_X1 U11120 ( .A1(n10962), .A2(n10961), .A3(n10960), .ZN(n10963) );
  NAND2_X1 U11121 ( .A1(n12343), .A2(n9690), .ZN(n12339) );
  OR2_X1 U11122 ( .A1(n10633), .A2(n10632), .ZN(n12115) );
  INV_X1 U11123 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10383) );
  CLKBUF_X2 U11125 ( .A(n9920), .Z(n12440) );
  NOR2_X1 U11126 ( .A1(n12279), .A2(n12280), .ZN(n12278) );
  AND2_X1 U11127 ( .A1(n12077), .A2(n15636), .ZN(n12151) );
  AND2_X1 U11128 ( .A1(n10149), .A2(n10147), .ZN(n12153) );
  NOR2_X1 U11129 ( .A1(n17012), .A2(n12740), .ZN(n12816) );
  NAND2_X1 U11130 ( .A1(n18742), .A2(n18249), .ZN(n18140) );
  CLKBUF_X3 U11131 ( .A(n12843), .Z(n9657) );
  AND2_X2 U11132 ( .A1(n11067), .A2(n20272), .ZN(n14073) );
  NAND2_X2 U11133 ( .A1(n13352), .A2(n20246), .ZN(n20954) );
  BUF_X1 U11134 ( .A(n11067), .Z(n20262) );
  NAND2_X1 U11135 ( .A1(n12336), .A2(n12385), .ZN(n12384) );
  OR2_X1 U11136 ( .A1(n10580), .A2(n13008), .ZN(n10511) );
  OAI21_X1 U11137 ( .B1(n12932), .B2(n12931), .A(n12930), .ZN(n12934) );
  NAND2_X2 U11138 ( .A1(n12716), .A2(n10585), .ZN(n12452) );
  NAND2_X1 U11139 ( .A1(n10444), .A2(n10443), .ZN(n12039) );
  OAI21_X1 U11140 ( .B1(n15161), .B2(n10155), .A(n9869), .ZN(n15147) );
  NOR2_X1 U11141 ( .A1(n16804), .A2(n16979), .ZN(n16798) );
  INV_X1 U11142 ( .A(n18749), .ZN(n18249) );
  AND2_X1 U11143 ( .A1(n14459), .A2(n13346), .ZN(n20140) );
  NAND2_X1 U11144 ( .A1(n13383), .A2(n11211), .ZN(n13306) );
  NAND2_X1 U11146 ( .A1(n13765), .A2(n10106), .ZN(n14978) );
  INV_X2 U11147 ( .A(n10406), .ZN(n10598) );
  NAND2_X1 U11148 ( .A1(n12039), .A2(n12040), .ZN(n9915) );
  INV_X1 U11149 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9640) );
  INV_X1 U11150 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20870) );
  NAND2_X1 U11151 ( .A1(n9915), .A2(n9797), .ZN(n15624) );
  AND4_X1 U11152 ( .A1(n12065), .A2(n12064), .A3(n12066), .A4(n12063), .ZN(
        n9638) );
  AND4_X1 U11153 ( .A1(n10928), .A2(n10927), .A3(n10926), .A4(n10925), .ZN(
        n9639) );
  XNOR2_X1 U11154 ( .A(n11182), .B(n11196), .ZN(n13369) );
  NOR2_X2 U11155 ( .A1(n12337), .A2(n12339), .ZN(n12363) );
  NAND2_X2 U11156 ( .A1(n10090), .A2(n13054), .ZN(n12447) );
  AND2_X2 U11157 ( .A1(n12111), .A2(n12133), .ZN(n12127) );
  NOR3_X4 U11158 ( .A1(n13557), .A2(n15566), .A3(n10176), .ZN(n15550) );
  AND2_X4 U11159 ( .A1(n12252), .A2(n15620), .ZN(n9666) );
  AND2_X2 U11160 ( .A1(n12252), .A2(n15620), .ZN(n9667) );
  INV_X2 U11162 ( .A(n10397), .ZN(n10398) );
  AND2_X1 U11163 ( .A1(n10586), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10357) );
  AOI21_X2 U11164 ( .B1(n12127), .B2(n13455), .A(n12126), .ZN(n12131) );
  XNOR2_X2 U11165 ( .A(n13907), .B(n10228), .ZN(n14956) );
  NAND2_X2 U11166 ( .A1(n14960), .A2(n13893), .ZN(n13907) );
  AND2_X4 U11167 ( .A1(n15632), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9641) );
  NOR2_X1 U11168 ( .A1(n12741), .A2(n12742), .ZN(n12842) );
  INV_X2 U11169 ( .A(n12452), .ZN(n10162) );
  INV_X2 U11170 ( .A(n16641), .ZN(n16979) );
  NOR2_X1 U11171 ( .A1(n19608), .A2(n19814), .ZN(n19650) );
  AND2_X1 U11172 ( .A1(n15445), .A2(n10175), .ZN(n14907) );
  OAI21_X1 U11173 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n16434), .A(n16618), 
        .ZN(n17939) );
  AND2_X1 U11174 ( .A1(n11233), .A2(n11232), .ZN(n13370) );
  NOR2_X1 U11175 ( .A1(n17403), .A2(n17577), .ZN(n17399) );
  INV_X2 U11176 ( .A(n17985), .ZN(n18716) );
  NAND2_X1 U11177 ( .A1(n11153), .A2(n14430), .ZN(n11184) );
  NOR2_X1 U11178 ( .A1(n13073), .A2(n10164), .ZN(n13658) );
  NAND3_X1 U11179 ( .A1(n20006), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19868), 
        .ZN(n19376) );
  NAND2_X1 U11180 ( .A1(n17898), .A2(n15881), .ZN(n15884) );
  NAND2_X1 U11181 ( .A1(n9724), .A2(n10066), .ZN(n12871) );
  NAND4_X1 U11182 ( .A1(n11042), .A2(n12970), .A3(n12969), .A4(n14305), .ZN(
        n13242) );
  OR2_X1 U11183 ( .A1(n17447), .A2(n15866), .ZN(n15886) );
  AND2_X1 U11184 ( .A1(n11049), .A2(n11064), .ZN(n11963) );
  INV_X1 U11185 ( .A(n12952), .ZN(n12970) );
  AND4_X2 U11186 ( .A1(n10421), .A2(n12468), .A3(n9733), .A4(n9671), .ZN(n9920) );
  BUF_X2 U11187 ( .A(n11040), .Z(n20292) );
  INV_X4 U11188 ( .A(n17404), .ZN(n18307) );
  AND3_X2 U11189 ( .A1(n9728), .A2(n10126), .A3(n15801), .ZN(n15870) );
  INV_X4 U11190 ( .A(n19378), .ZN(n12215) );
  CLKBUF_X1 U11191 ( .A(n11139), .Z(n11876) );
  INV_X2 U11192 ( .A(n11923), .ZN(n9643) );
  CLKBUF_X2 U11193 ( .A(n11003), .Z(n11925) );
  INV_X2 U11194 ( .A(n11810), .ZN(n11111) );
  INV_X1 U11195 ( .A(n11849), .ZN(n11676) );
  BUF_X2 U11196 ( .A(n10957), .Z(n11926) );
  CLKBUF_X1 U11197 ( .A(n11129), .Z(n11884) );
  INV_X2 U11198 ( .A(n11700), .ZN(n9658) );
  AND2_X2 U11199 ( .A1(n10911), .A2(n10913), .ZN(n10957) );
  NAND2_X1 U11200 ( .A1(n13177), .A2(n10912), .ZN(n11700) );
  OAI21_X1 U11201 ( .B1(n12564), .B2(n16324), .A(n12551), .ZN(n12552) );
  AOI21_X1 U11202 ( .B1(n12539), .B2(n12537), .A(n12538), .ZN(n12555) );
  XNOR2_X1 U11203 ( .A(n9899), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14666) );
  AND3_X1 U11204 ( .A1(n9944), .A2(n9943), .A3(n9945), .ZN(n15419) );
  OR2_X1 U11205 ( .A1(n9714), .A2(n14463), .ZN(n9899) );
  NOR2_X1 U11206 ( .A1(n14471), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14463) );
  AOI211_X1 U11207 ( .C1(n16138), .C2(n14510), .A(n14509), .B(n14508), .ZN(
        n14511) );
  NAND2_X1 U11208 ( .A1(n15148), .A2(n10000), .ZN(n10005) );
  INV_X1 U11209 ( .A(n9924), .ZN(n15214) );
  NAND2_X1 U11210 ( .A1(n14504), .A2(n10030), .ZN(n14471) );
  AOI211_X1 U11211 ( .C1(n16138), .C2(n14502), .A(n14501), .B(n14500), .ZN(
        n14503) );
  NAND2_X1 U11212 ( .A1(n9786), .A2(n9785), .ZN(n15251) );
  OR2_X1 U11213 ( .A1(n14480), .A2(n14512), .ZN(n14485) );
  AND2_X1 U11214 ( .A1(n14453), .A2(n14454), .ZN(n10030) );
  NAND2_X1 U11215 ( .A1(n14505), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14504) );
  AOI21_X1 U11216 ( .B1(n15256), .B2(n9678), .A(n9925), .ZN(n9924) );
  AOI21_X1 U11217 ( .B1(n16490), .B2(n18070), .A(n10118), .ZN(n16492) );
  NAND2_X1 U11218 ( .A1(n9870), .A2(n15263), .ZN(n15161) );
  AND2_X2 U11219 ( .A1(n14087), .A2(n11900), .ZN(n14089) );
  OAI21_X1 U11220 ( .B1(n14110), .B2(n14111), .A(n14099), .ZN(n14499) );
  AND2_X1 U11221 ( .A1(n9862), .A2(n10119), .ZN(n16490) );
  OR2_X1 U11222 ( .A1(n10200), .A2(n9735), .ZN(n9789) );
  NOR2_X1 U11223 ( .A1(n12507), .A2(n9800), .ZN(n9799) );
  AND2_X1 U11224 ( .A1(n9981), .A2(n10159), .ZN(n9871) );
  NAND2_X1 U11226 ( .A1(n9856), .A2(n16444), .ZN(n15965) );
  OR2_X1 U11227 ( .A1(n9984), .A2(n9983), .ZN(n9872) );
  XNOR2_X1 U11228 ( .A(n12446), .B(n12445), .ZN(n16279) );
  INV_X1 U11229 ( .A(n9983), .ZN(n9982) );
  AND2_X1 U11230 ( .A1(n15603), .A2(n12298), .ZN(n9984) );
  AND2_X1 U11231 ( .A1(n16341), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10202) );
  OR2_X1 U11232 ( .A1(n12304), .A2(n9754), .ZN(n9983) );
  XNOR2_X1 U11233 ( .A(n12202), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16341) );
  NAND2_X1 U11234 ( .A1(n12200), .A2(n12433), .ZN(n12202) );
  OR2_X1 U11235 ( .A1(n13848), .A2(n13870), .ZN(n10094) );
  NAND2_X1 U11236 ( .A1(n9793), .A2(n9987), .ZN(n13649) );
  NAND2_X1 U11237 ( .A1(n12189), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13654) );
  NAND2_X1 U11238 ( .A1(n10038), .A2(n10037), .ZN(n10036) );
  NOR2_X1 U11239 ( .A1(n17608), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17607) );
  NAND2_X1 U11240 ( .A1(n9846), .A2(n9845), .ZN(n17608) );
  OAI21_X1 U11241 ( .B1(n12295), .B2(n12433), .A(n19142), .ZN(n13651) );
  XNOR2_X1 U11242 ( .A(n12163), .B(n12162), .ZN(n12295) );
  NAND2_X1 U11243 ( .A1(n12455), .A2(n10861), .ZN(n15308) );
  INV_X1 U11244 ( .A(n12558), .ZN(n15033) );
  NOR2_X2 U11245 ( .A1(n9694), .A2(n14903), .ZN(n14904) );
  AND2_X1 U11246 ( .A1(n12414), .A2(n9711), .ZN(n9880) );
  AND2_X1 U11247 ( .A1(n14569), .A2(n14571), .ZN(n16086) );
  OR2_X1 U11248 ( .A1(n10003), .A2(n12574), .ZN(n9996) );
  AND2_X2 U11249 ( .A1(n13639), .A2(n13638), .ZN(n13765) );
  OR2_X1 U11250 ( .A1(n15020), .A2(n15019), .ZN(n15022) );
  OR2_X1 U11251 ( .A1(n12420), .A2(n15365), .ZN(n15121) );
  NAND2_X1 U11252 ( .A1(n17684), .A2(n9843), .ZN(n9847) );
  AND2_X1 U11253 ( .A1(n9716), .A2(n12103), .ZN(n9976) );
  NOR2_X1 U11254 ( .A1(n19789), .A2(n19788), .ZN(n19851) );
  NAND2_X1 U11255 ( .A1(n11306), .A2(n11305), .ZN(n13432) );
  OR2_X1 U11256 ( .A1(n14886), .A2(n9942), .ZN(n12420) );
  CLKBUF_X1 U11257 ( .A(n14889), .Z(n14909) );
  AND2_X1 U11258 ( .A1(n15915), .A2(n9844), .ZN(n9843) );
  OR2_X1 U11259 ( .A1(n13479), .A2(n13480), .ZN(n13486) );
  OAI22_X1 U11260 ( .A1(n17943), .A2(n18127), .B1(n17850), .B2(n18125), .ZN(
        n17841) );
  OAI21_X1 U11261 ( .B1(n14403), .B2(n14429), .A(n14405), .ZN(n14406) );
  NAND2_X1 U11262 ( .A1(n12047), .A2(n19175), .ZN(n12134) );
  AND2_X1 U11263 ( .A1(n12059), .A2(n12058), .ZN(n12064) );
  NAND2_X1 U11264 ( .A1(n10149), .A2(n10148), .ZN(n12135) );
  AND2_X1 U11265 ( .A1(n13203), .A2(n13012), .ZN(n13125) );
  NAND2_X1 U11266 ( .A1(n9926), .A2(n15166), .ZN(n9925) );
  NOR2_X1 U11267 ( .A1(n10494), .A2(n13119), .ZN(n13194) );
  NAND2_X1 U11268 ( .A1(n12888), .A2(n12887), .ZN(n12932) );
  OR2_X1 U11269 ( .A1(n12732), .A2(n12731), .ZN(n12888) );
  OR2_X2 U11270 ( .A1(n18720), .A2(n18925), .ZN(n16618) );
  XNOR2_X1 U11271 ( .A(n12726), .B(n12886), .ZN(n12732) );
  NAND2_X2 U11272 ( .A1(n20161), .A2(n20292), .ZN(n16075) );
  OAI21_X2 U11273 ( .B1(n15624), .B2(n12940), .A(n12687), .ZN(n12726) );
  NOR2_X1 U11274 ( .A1(n16783), .A2(n17129), .ZN(n17117) );
  NAND2_X1 U11275 ( .A1(n12948), .A2(n20868), .ZN(n11233) );
  XNOR2_X1 U11276 ( .A(n11103), .B(n11102), .ZN(n11187) );
  XNOR2_X1 U11277 ( .A(n13178), .B(n20406), .ZN(n12948) );
  NAND2_X1 U11278 ( .A1(n9798), .A2(n9914), .ZN(n9797) );
  OR2_X1 U11279 ( .A1(n11184), .A2(n11183), .ZN(n11185) );
  XNOR2_X1 U11280 ( .A(n11184), .B(n11175), .ZN(n11195) );
  NOR2_X1 U11281 ( .A1(n17439), .A2(n21109), .ZN(n17434) );
  NAND2_X1 U11282 ( .A1(n10480), .A2(n10479), .ZN(n12038) );
  CLKBUF_X1 U11283 ( .A(n13347), .Z(n20667) );
  NOR2_X2 U11284 ( .A1(n18140), .A2(n18065), .ZN(n18006) );
  OAI22_X1 U11285 ( .A1(n15607), .A2(n10721), .B1(n9942), .B2(n10720), .ZN(
        n16370) );
  NAND2_X1 U11286 ( .A1(n17316), .A2(n17404), .ZN(n17458) );
  OR2_X1 U11287 ( .A1(n13587), .A2(n13588), .ZN(n13604) );
  INV_X1 U11288 ( .A(n18745), .ZN(n18065) );
  NAND2_X1 U11289 ( .A1(n11178), .A2(n11177), .ZN(n20301) );
  AOI21_X2 U11290 ( .B1(n15981), .B2(n15980), .A(n18925), .ZN(n17316) );
  XNOR2_X1 U11291 ( .A(n15884), .B(n15883), .ZN(n17882) );
  NAND2_X1 U11292 ( .A1(n20369), .A2(n11176), .ZN(n11179) );
  CLKBUF_X1 U11293 ( .A(n11204), .Z(n20368) );
  NOR2_X2 U11294 ( .A1(n13428), .A2(n10041), .ZN(n16235) );
  AND2_X1 U11295 ( .A1(n11106), .A2(n11104), .ZN(n11176) );
  OR2_X1 U11296 ( .A1(n10656), .A2(n10653), .ZN(n13072) );
  AOI21_X1 U11297 ( .B1(n13077), .B2(n9697), .A(n10652), .ZN(n10656) );
  NOR2_X1 U11298 ( .A1(n12313), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U11299 ( .A1(n10463), .A2(n10462), .ZN(n12041) );
  AOI21_X1 U11300 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n10442), .A(n10441), 
        .ZN(n10443) );
  NOR2_X1 U11301 ( .A1(n19276), .A2(n16417), .ZN(n19185) );
  NAND2_X1 U11302 ( .A1(n11060), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11074) );
  INV_X2 U11303 ( .A(n17570), .ZN(n9646) );
  NAND2_X1 U11304 ( .A1(n16498), .A2(n16495), .ZN(n17849) );
  NAND2_X1 U11305 ( .A1(n13699), .A2(n17510), .ZN(n16617) );
  NAND2_X1 U11306 ( .A1(n13686), .A2(n9886), .ZN(n17510) );
  OR2_X1 U11307 ( .A1(n10673), .A2(n10672), .ZN(n13461) );
  AND2_X1 U11308 ( .A1(n12714), .A2(n12712), .ZN(n10637) );
  NAND2_X1 U11309 ( .A1(n10420), .A2(n10419), .ZN(n10435) );
  AND3_X1 U11310 ( .A1(n10692), .A2(n10691), .A3(n10690), .ZN(n13615) );
  NAND2_X1 U11311 ( .A1(n10616), .A2(n10615), .ZN(n12714) );
  CLKBUF_X1 U11312 ( .A(n13113), .Z(n14055) );
  NAND2_X1 U11313 ( .A1(n12465), .A2(n10433), .ZN(n10415) );
  NOR2_X1 U11314 ( .A1(n15864), .A2(n13696), .ZN(n13686) );
  NOR2_X1 U11315 ( .A1(n20954), .A2(n13238), .ZN(n11052) );
  NAND2_X1 U11316 ( .A1(n11148), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14430) );
  NOR2_X1 U11317 ( .A1(n17454), .A2(n15868), .ZN(n15878) );
  NAND2_X1 U11318 ( .A1(n13673), .A2(n18301), .ZN(n18744) );
  OR2_X1 U11319 ( .A1(n11145), .A2(n11144), .ZN(n13270) );
  CLKBUF_X1 U11320 ( .A(n11050), .Z(n12972) );
  AND2_X1 U11321 ( .A1(n11048), .A2(n20292), .ZN(n11064) );
  NOR4_X1 U11322 ( .A1(n13683), .A2(n13672), .A3(n13685), .A4(n13677), .ZN(
        n13688) );
  OR2_X1 U11323 ( .A1(n18289), .A2(n18307), .ZN(n13696) );
  AND2_X1 U11324 ( .A1(n12015), .A2(n11066), .ZN(n12869) );
  NAND2_X1 U11325 ( .A1(n9671), .A2(n9680), .ZN(n10418) );
  CLKBUF_X1 U11326 ( .A(n10410), .Z(n16418) );
  OR2_X1 U11327 ( .A1(n17459), .A2(n15870), .ZN(n15868) );
  INV_X1 U11328 ( .A(n12243), .ZN(n10378) );
  AND2_X1 U11330 ( .A1(n10598), .A2(n19632), .ZN(n10619) );
  CLKBUF_X3 U11331 ( .A(n10393), .Z(n9660) );
  NAND3_X1 U11332 ( .A1(n12825), .A2(n12824), .A3(n12823), .ZN(n17317) );
  INV_X1 U11333 ( .A(n20246), .ZN(n11043) );
  INV_X1 U11334 ( .A(n12221), .ZN(n10421) );
  OR2_X2 U11335 ( .A1(n10719), .A2(n10718), .ZN(n12433) );
  OR2_X2 U11336 ( .A1(n16566), .A2(n16512), .ZN(n16568) );
  INV_X1 U11337 ( .A(n12237), .ZN(n12467) );
  AND4_X1 U11338 ( .A1(n10920), .A2(n10919), .A3(n10918), .A4(n10917), .ZN(
        n10921) );
  AND4_X1 U11339 ( .A1(n10938), .A2(n10062), .A3(n10942), .A4(n10941), .ZN(
        n10061) );
  AND4_X1 U11340 ( .A1(n10956), .A2(n10955), .A3(n10954), .A4(n10953), .ZN(
        n10964) );
  NAND2_X1 U11342 ( .A1(n10338), .A2(n10337), .ZN(n10401) );
  AND4_X1 U11343 ( .A1(n11011), .A2(n11010), .A3(n11009), .A4(n11008), .ZN(
        n11018) );
  NOR2_X1 U11344 ( .A1(n11007), .A2(n11006), .ZN(n11019) );
  AND2_X1 U11345 ( .A1(n10940), .A2(n10943), .ZN(n10062) );
  AND4_X1 U11346 ( .A1(n10981), .A2(n10980), .A3(n10979), .A4(n10978), .ZN(
        n10982) );
  OR2_X1 U11347 ( .A1(n11697), .A2(n10985), .ZN(n10987) );
  INV_X2 U11348 ( .A(n11090), .ZN(n11883) );
  INV_X2 U11349 ( .A(n20923), .ZN(n9647) );
  AND2_X1 U11350 ( .A1(n11023), .A2(n11022), .ZN(n11026) );
  NAND2_X2 U11351 ( .A1(n18939), .A2(n18807), .ZN(n18855) );
  NAND4_X1 U11352 ( .A1(n10219), .A2(n10299), .A3(n10298), .A4(n10297), .ZN(
        n10300) );
  NAND2_X1 U11353 ( .A1(n10331), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10338) );
  NAND2_X1 U11354 ( .A1(n9703), .A2(n10310), .ZN(n10311) );
  NAND2_X1 U11355 ( .A1(n10294), .A2(n10293), .ZN(n10301) );
  AND2_X1 U11356 ( .A1(n10309), .A2(n10308), .ZN(n10310) );
  CLKBUF_X3 U11357 ( .A(n12839), .Z(n17269) );
  AND2_X1 U11358 ( .A1(n10292), .A2(n10291), .ZN(n10293) );
  AND2_X2 U11359 ( .A1(n13964), .A2(n10383), .ZN(n13837) );
  AND2_X2 U11360 ( .A1(n10903), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11028) );
  NAND2_X2 U11361 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19995), .ZN(n19994) );
  NAND2_X2 U11362 ( .A1(n19995), .A2(n19951), .ZN(n19997) );
  AND2_X2 U11363 ( .A1(n13971), .A2(n10383), .ZN(n13838) );
  AND2_X2 U11364 ( .A1(n9663), .A2(n10383), .ZN(n10663) );
  INV_X1 U11365 ( .A(n11700), .ZN(n10968) );
  BUF_X2 U11366 ( .A(n10591), .Z(n13972) );
  NAND2_X1 U11367 ( .A1(n12965), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11031) );
  CLKBUF_X3 U11368 ( .A(n10318), .Z(n13968) );
  INV_X4 U11369 ( .A(n15803), .ZN(n9648) );
  OR2_X1 U11370 ( .A1(n12741), .A2(n18739), .ZN(n10212) );
  OR2_X1 U11371 ( .A1(n12745), .A2(n17012), .ZN(n9706) );
  INV_X2 U11372 ( .A(n16606), .ZN(n16608) );
  INV_X2 U11373 ( .A(n18940), .ZN(n18939) );
  INV_X4 U11374 ( .A(n10230), .ZN(n9650) );
  AND2_X2 U11375 ( .A1(n18751), .A2(n18540), .ZN(n18541) );
  INV_X1 U11376 ( .A(n13055), .ZN(n9662) );
  NAND2_X1 U11377 ( .A1(n18909), .A2(n18901), .ZN(n17012) );
  NAND2_X1 U11378 ( .A1(n18883), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12744) );
  NAND2_X1 U11379 ( .A1(n18883), .A2(n18891), .ZN(n12740) );
  NAND2_X1 U11380 ( .A1(n18901), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12742) );
  AND2_X1 U11381 ( .A1(n10914), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10915) );
  NAND2_X1 U11382 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18731) );
  NAND2_X1 U11383 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18739) );
  NOR2_X2 U11384 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15632) );
  NOR2_X1 U11385 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10288) );
  NAND3_X1 U11386 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13055) );
  AND2_X1 U11387 ( .A1(n12076), .A2(n12060), .ZN(n19859) );
  AND2_X1 U11388 ( .A1(n12077), .A2(n12060), .ZN(n12141) );
  NOR2_X1 U11389 ( .A1(n14975), .A2(n14974), .ZN(n14973) );
  AND2_X1 U11390 ( .A1(n9700), .A2(n12073), .ZN(n12140) );
  NAND2_X2 U11391 ( .A1(n14277), .A2(n14278), .ZN(n14271) );
  NOR2_X4 U11392 ( .A1(n14194), .A2(n10190), .ZN(n14277) );
  NOR2_X1 U11393 ( .A1(n12941), .A2(n12057), .ZN(n12076) );
  OR2_X1 U11394 ( .A1(n18739), .A2(n12740), .ZN(n15803) );
  AND2_X1 U11395 ( .A1(n13056), .A2(n15646), .ZN(n9651) );
  AND2_X1 U11396 ( .A1(n13056), .A2(n15646), .ZN(n9652) );
  AND2_X1 U11397 ( .A1(n13056), .A2(n15646), .ZN(n9655) );
  AND3_X2 U11398 ( .A1(n15620), .A2(n15646), .A3(n13713), .ZN(n10318) );
  AND2_X2 U11399 ( .A1(n13056), .A2(n15646), .ZN(n9656) );
  NOR2_X2 U11400 ( .A1(n14133), .A2(n14120), .ZN(n10050) );
  NAND2_X2 U11401 ( .A1(n10326), .A2(n10325), .ZN(n10397) );
  NAND2_X1 U11402 ( .A1(n18891), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12741) );
  NOR2_X1 U11403 ( .A1(n18929), .A2(n16618), .ZN(n9653) );
  XNOR2_X2 U11404 ( .A(n12044), .B(n12043), .ZN(n12068) );
  NAND2_X2 U11405 ( .A1(n9953), .A2(n10455), .ZN(n12044) );
  NOR2_X2 U11406 ( .A1(n14257), .A2(n14342), .ZN(n14154) );
  INV_X1 U11407 ( .A(n10431), .ZN(n10432) );
  AND2_X2 U11408 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12252) );
  NAND2_X2 U11409 ( .A1(n14193), .A2(n14196), .ZN(n14194) );
  AOI21_X4 U11410 ( .B1(n14208), .B2(n11473), .A(n11472), .ZN(n14193) );
  OR2_X2 U11411 ( .A1(n12941), .A2(n19191), .ZN(n12075) );
  NAND2_X4 U11412 ( .A1(n9878), .A2(n9876), .ZN(n12941) );
  NOR2_X1 U11413 ( .A1(n12742), .A2(n12745), .ZN(n12843) );
  INV_X1 U11414 ( .A(n11845), .ZN(n9659) );
  INV_X2 U11415 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15620) );
  OAI21_X2 U11416 ( .B1(n10094), .B2(n14973), .A(n10093), .ZN(n13889) );
  NOR2_X2 U11417 ( .A1(n14956), .A2(n14955), .ZN(n14954) );
  INV_X2 U11418 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15646) );
  AND2_X1 U11419 ( .A1(n13907), .A2(n10228), .ZN(n13908) );
  NAND2_X2 U11420 ( .A1(n12198), .A2(n15602), .ZN(n15297) );
  NOR2_X2 U11421 ( .A1(n13534), .A2(n13540), .ZN(n13539) );
  INV_X4 U11422 ( .A(n12060), .ZN(n15636) );
  OR2_X2 U11423 ( .A1(n13927), .A2(n13926), .ZN(n13930) );
  NAND2_X1 U11424 ( .A1(n10336), .A2(n10383), .ZN(n10337) );
  AND2_X1 U11425 ( .A1(n10407), .A2(n10398), .ZN(n12468) );
  AND4_X1 U11426 ( .A1(n12237), .A2(n10407), .A3(n10397), .A4(n10401), .ZN(
        n10405) );
  OAI222_X1 U11427 ( .A1(n16075), .A2(n14507), .B1(n14253), .B2(n20161), .C1(
        n14252), .C2(n16076), .ZN(P1_U2846) );
  OAI21_X2 U11428 ( .B1(n14125), .B2(n14123), .A(n14124), .ZN(n14507) );
  AOI21_X1 U11429 ( .B1(n10461), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10474), .ZN(n10476) );
  NAND2_X4 U11430 ( .A1(n9974), .A2(n9972), .ZN(n19378) );
  INV_X4 U11431 ( .A(n10583), .ZN(n10406) );
  XNOR2_X2 U11433 ( .A(n14077), .B(n14089), .ZN(n14078) );
  INV_X2 U11434 ( .A(n13055), .ZN(n9663) );
  INV_X1 U11435 ( .A(n9662), .ZN(n9664) );
  NAND2_X2 U11436 ( .A1(n13209), .A2(n13210), .ZN(n13379) );
  NAND2_X2 U11437 ( .A1(n15206), .A2(n12486), .ZN(n15185) );
  NAND2_X4 U11438 ( .A1(n9788), .A2(n9787), .ZN(n15206) );
  NOR2_X2 U11439 ( .A1(n13379), .A2(n10102), .ZN(n13639) );
  BUF_X4 U11440 ( .A(n10431), .Z(n10473) );
  OAI21_X2 U11441 ( .B1(n14945), .B2(n13943), .A(n14940), .ZN(n14935) );
  NOR2_X2 U11442 ( .A1(n14947), .A2(n14946), .ZN(n14945) );
  NOR2_X2 U11443 ( .A1(n14978), .A2(n14980), .ZN(n13847) );
  AND2_X2 U11444 ( .A1(n10350), .A2(n10349), .ZN(n10412) );
  NAND2_X1 U11445 ( .A1(n12944), .A2(n12943), .ZN(n12995) );
  AND2_X1 U11446 ( .A1(n12941), .A2(n12053), .ZN(n19429) );
  NOR2_X2 U11447 ( .A1(n12078), .A2(n19175), .ZN(n12145) );
  AND2_X2 U11448 ( .A1(n13968), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10601) );
  INV_X1 U11449 ( .A(n13242), .ZN(n9816) );
  NAND2_X1 U11450 ( .A1(n10435), .A2(n9719), .ZN(n10145) );
  NAND2_X1 U11451 ( .A1(n10417), .A2(n10397), .ZN(n10413) );
  OR2_X1 U11452 ( .A1(n16291), .A2(n12404), .ZN(n12421) );
  NAND2_X1 U11453 ( .A1(n12456), .A2(n12468), .ZN(n13054) );
  NAND2_X1 U11454 ( .A1(n12271), .A2(n19274), .ZN(n12477) );
  AND2_X1 U11455 ( .A1(n9918), .A2(n9916), .ZN(n12097) );
  AOI21_X1 U11456 ( .B1(n9721), .B2(n9919), .A(n10406), .ZN(n9918) );
  INV_X1 U11457 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11502) );
  NAND2_X1 U11458 ( .A1(n12871), .A2(n10065), .ZN(n10063) );
  OAI21_X1 U11459 ( .B1(n11060), .B2(n12871), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11054) );
  NAND3_X1 U11460 ( .A1(n9897), .A2(n9896), .A3(n11059), .ZN(n10198) );
  NAND2_X1 U11461 ( .A1(n11060), .A2(n9898), .ZN(n9897) );
  OAI22_X1 U11462 ( .A1(n10568), .A2(n10560), .B1(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20023), .ZN(n10566) );
  NOR2_X1 U11463 ( .A1(n10153), .A2(n12132), .ZN(n10151) );
  NAND2_X1 U11464 ( .A1(n12457), .A2(n19378), .ZN(n10416) );
  AND2_X1 U11465 ( .A1(n14111), .A2(n9745), .ZN(n10197) );
  NAND2_X1 U11466 ( .A1(n12949), .A2(n14012), .ZN(n13113) );
  NAND2_X1 U11467 ( .A1(n10068), .A2(n14565), .ZN(n9911) );
  NAND2_X1 U11468 ( .A1(n14043), .A2(n14073), .ZN(n14047) );
  NAND2_X1 U11469 ( .A1(n14612), .A2(n14439), .ZN(n14596) );
  NAND2_X1 U11470 ( .A1(n14628), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9826) );
  INV_X1 U11471 ( .A(n14047), .ZN(n14050) );
  INV_X1 U11472 ( .A(n13429), .ZN(n10045) );
  NAND2_X1 U11473 ( .A1(n14053), .A2(n14043), .ZN(n14048) );
  NAND2_X1 U11475 ( .A1(n9704), .A2(n13221), .ZN(n10999) );
  AND2_X1 U11476 ( .A1(n12013), .A2(n12012), .ZN(n12987) );
  OR2_X2 U11477 ( .A1(n11039), .A2(n11038), .ZN(n11067) );
  OAI21_X1 U11478 ( .B1(n20955), .B2(n16262), .A(n13184), .ZN(n20245) );
  INV_X1 U11479 ( .A(n15956), .ZN(n13184) );
  NOR2_X1 U11480 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n12412), .ZN(n12401) );
  NAND2_X1 U11481 ( .A1(n12291), .A2(n10137), .ZN(n12306) );
  INV_X1 U11482 ( .A(n14876), .ZN(n10169) );
  INV_X1 U11483 ( .A(n14990), .ZN(n10107) );
  NAND2_X1 U11484 ( .A1(n12215), .A2(n10406), .ZN(n12224) );
  NAND2_X1 U11485 ( .A1(n12204), .A2(n12502), .ZN(n15179) );
  NAND2_X1 U11486 ( .A1(n12184), .A2(n12183), .ZN(n12190) );
  INV_X1 U11487 ( .A(n13611), .ZN(n9988) );
  INV_X1 U11488 ( .A(n10866), .ZN(n12273) );
  AND2_X1 U11489 ( .A1(n10232), .A2(n19422), .ZN(n10150) );
  INV_X1 U11490 ( .A(n12072), .ZN(n12073) );
  NOR2_X1 U11491 ( .A1(n12741), .A2(n12743), .ZN(n15796) );
  NOR2_X1 U11492 ( .A1(n17510), .A2(n18281), .ZN(n13704) );
  AND2_X1 U11493 ( .A1(n18943), .A2(n16617), .ZN(n13694) );
  NOR2_X1 U11494 ( .A1(n13694), .A2(n13704), .ZN(n15743) );
  NAND2_X1 U11495 ( .A1(n17858), .A2(n15892), .ZN(n10129) );
  NAND2_X1 U11496 ( .A1(n17920), .A2(n15873), .ZN(n15876) );
  XNOR2_X1 U11497 ( .A(n15870), .B(n17459), .ZN(n15872) );
  OR2_X2 U11498 ( .A1(n12306), .A2(n9660), .ZN(n12435) );
  NAND2_X1 U11499 ( .A1(n12278), .A2(n12273), .ZN(n12290) );
  AND2_X1 U11500 ( .A1(n12568), .A2(n12544), .ZN(n12546) );
  INV_X1 U11501 ( .A(n12578), .ZN(n12426) );
  NAND2_X1 U11502 ( .A1(n12329), .A2(n9921), .ZN(n9870) );
  NOR2_X1 U11503 ( .A1(n15262), .A2(n9922), .ZN(n9921) );
  INV_X1 U11504 ( .A(n12328), .ZN(n9922) );
  INV_X1 U11505 ( .A(n12127), .ZN(n13454) );
  OAI22_X1 U11506 ( .A1(n10448), .A2(n10447), .B1(n9920), .B2(n10446), .ZN(
        n10451) );
  OAI21_X1 U11507 ( .B1(n10213), .B2(n13704), .A(n9889), .ZN(n15981) );
  NOR2_X1 U11508 ( .A1(n9891), .A2(n9890), .ZN(n9889) );
  AND2_X1 U11509 ( .A1(n17618), .A2(n9770), .ZN(n9845) );
  NAND2_X1 U11510 ( .A1(n9839), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9846) );
  INV_X1 U11511 ( .A(n18281), .ZN(n18929) );
  NOR2_X1 U11512 ( .A1(n17849), .A2(n17945), .ZN(n9852) );
  NAND2_X1 U11513 ( .A1(n17731), .A2(n17849), .ZN(n17684) );
  NAND2_X1 U11514 ( .A1(n17732), .A2(n18056), .ZN(n17731) );
  NAND2_X1 U11515 ( .A1(n18281), .A2(n18006), .ZN(n17985) );
  AND2_X1 U11516 ( .A1(n9683), .A2(n13130), .ZN(n10096) );
  NAND2_X1 U11517 ( .A1(n10167), .A2(n9698), .ZN(n9800) );
  NOR2_X1 U11518 ( .A1(n14938), .A2(n15589), .ZN(n9958) );
  INV_X1 U11519 ( .A(n15589), .ZN(n19369) );
  NOR2_X1 U11520 ( .A1(n9821), .A2(n9819), .ZN(n9818) );
  NAND2_X1 U11521 ( .A1(n20246), .A2(n9820), .ZN(n9819) );
  INV_X1 U11522 ( .A(n12865), .ZN(n9820) );
  INV_X1 U11523 ( .A(n11275), .ZN(n11276) );
  INV_X1 U11524 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11907) );
  INV_X1 U11525 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11919) );
  AND2_X1 U11526 ( .A1(n11327), .A2(n11326), .ZN(n11338) );
  INV_X1 U11527 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11688) );
  INV_X1 U11528 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11692) );
  INV_X1 U11529 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11693) );
  OAI21_X1 U11530 ( .B1(n10952), .B2(n11903), .A(n10969), .ZN(n10179) );
  NOR2_X1 U11531 ( .A1(n10974), .A2(n10973), .ZN(n10984) );
  AND2_X1 U11532 ( .A1(n12309), .A2(n12300), .ZN(n10137) );
  AND2_X1 U11533 ( .A1(n10137), .A2(n10136), .ZN(n10135) );
  INV_X1 U11534 ( .A(n12305), .ZN(n10136) );
  AOI21_X1 U11535 ( .B1(n13058), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10423), 
        .ZN(n10424) );
  NAND2_X1 U11536 ( .A1(n10461), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10425) );
  AND2_X1 U11537 ( .A1(n16419), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10423) );
  NAND2_X1 U11538 ( .A1(n10421), .A2(n12468), .ZN(n10445) );
  NOR2_X1 U11539 ( .A1(n10583), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10585) );
  NOR2_X1 U11540 ( .A1(n15636), .A2(n12728), .ZN(n10148) );
  NAND2_X1 U11541 ( .A1(n10559), .A2(n10558), .ZN(n10568) );
  INV_X1 U11542 ( .A(n12206), .ZN(n10570) );
  OR2_X1 U11543 ( .A1(n12768), .A2(n12769), .ZN(n12764) );
  NOR2_X1 U11544 ( .A1(n11047), .A2(n11965), .ZN(n12015) );
  NAND2_X1 U11545 ( .A1(n14825), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11896) );
  NOR2_X1 U11546 ( .A1(n9687), .A2(n10182), .ZN(n10181) );
  INV_X1 U11547 ( .A(n10234), .ZN(n10182) );
  INV_X1 U11548 ( .A(n11896), .ZN(n11938) );
  NAND2_X1 U11549 ( .A1(n9775), .A2(n11516), .ZN(n10193) );
  CLKBUF_X1 U11551 ( .A(n11138), .Z(n11880) );
  NOR2_X2 U11552 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13340) );
  INV_X1 U11553 ( .A(n13537), .ZN(n11336) );
  OR2_X1 U11554 ( .A1(n20292), .A2(n20870), .ZN(n11936) );
  INV_X1 U11555 ( .A(n13340), .ZN(n11935) );
  NOR2_X1 U11556 ( .A1(n10058), .A2(n10059), .ZN(n9824) );
  INV_X1 U11557 ( .A(n14171), .ZN(n10054) );
  NAND2_X1 U11558 ( .A1(n10070), .A2(n9777), .ZN(n10069) );
  NOR2_X1 U11559 ( .A1(n14573), .A2(n9717), .ZN(n10037) );
  INV_X1 U11560 ( .A(n14570), .ZN(n10038) );
  INV_X1 U11561 ( .A(n14048), .ZN(n14034) );
  AND4_X1 U11562 ( .A1(n11115), .A2(n11114), .A3(n11113), .A4(n11112), .ZN(
        n11124) );
  NAND2_X1 U11563 ( .A1(n13286), .A2(n13285), .ZN(n13287) );
  OR2_X1 U11564 ( .A1(n13284), .A2(n13283), .ZN(n13285) );
  OAI21_X1 U11565 ( .B1(n11063), .B2(n11044), .A(n11043), .ZN(n11053) );
  AND2_X1 U11566 ( .A1(n12985), .A2(n12984), .ZN(n13234) );
  AND2_X1 U11567 ( .A1(n11213), .A2(n20857), .ZN(n20542) );
  INV_X1 U11568 ( .A(n12417), .ZN(n12429) );
  OR2_X1 U11569 ( .A1(n12415), .A2(n12416), .ZN(n12417) );
  NOR2_X1 U11570 ( .A1(n15145), .A2(n10026), .ZN(n10025) );
  INV_X1 U11571 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10026) );
  AND2_X1 U11572 ( .A1(n12291), .A2(n12300), .ZN(n12311) );
  NAND2_X1 U11573 ( .A1(n13892), .A2(n13891), .ZN(n13893) );
  INV_X1 U11574 ( .A(n13889), .ZN(n13892) );
  NOR2_X1 U11575 ( .A1(n10239), .A2(n10016), .ZN(n10015) );
  INV_X1 U11576 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U11577 ( .A1(n15298), .A2(n16374), .ZN(n10206) );
  INV_X1 U11578 ( .A(n15298), .ZN(n10205) );
  OR2_X1 U11579 ( .A1(n10649), .A2(n10648), .ZN(n12118) );
  NAND2_X1 U11580 ( .A1(n12429), .A2(n12428), .ZN(n12434) );
  INV_X1 U11581 ( .A(n15113), .ZN(n10004) );
  NOR2_X1 U11582 ( .A1(n12574), .A2(n9999), .ZN(n9998) );
  INV_X1 U11583 ( .A(n10000), .ZN(n9999) );
  INV_X1 U11584 ( .A(n14880), .ZN(n10089) );
  OR2_X1 U11585 ( .A1(n10076), .A2(n10075), .ZN(n10074) );
  INV_X1 U11586 ( .A(n14993), .ZN(n10075) );
  NOR2_X1 U11587 ( .A1(n9934), .A2(n15164), .ZN(n9932) );
  NOR2_X1 U11588 ( .A1(n15163), .A2(n9938), .ZN(n9937) );
  INV_X1 U11589 ( .A(n15254), .ZN(n9938) );
  NOR2_X1 U11590 ( .A1(n13211), .A2(n10086), .ZN(n10085) );
  INV_X1 U11591 ( .A(n13124), .ZN(n10086) );
  INV_X1 U11592 ( .A(n12187), .ZN(n12186) );
  NOR2_X1 U11593 ( .A1(n10406), .A2(n10408), .ZN(n10409) );
  NAND2_X1 U11594 ( .A1(n10416), .A2(n10415), .ZN(n10436) );
  INV_X1 U11595 ( .A(n13008), .ZN(n13924) );
  AND2_X1 U11596 ( .A1(n10585), .A2(n10584), .ZN(n10825) );
  INV_X1 U11597 ( .A(n10656), .ZN(n10163) );
  NAND2_X1 U11598 ( .A1(n10399), .A2(n10398), .ZN(n10400) );
  AND2_X1 U11599 ( .A1(n12467), .A2(n19422), .ZN(n10395) );
  NAND2_X1 U11600 ( .A1(n15636), .A2(n12728), .ZN(n12072) );
  AND3_X1 U11601 ( .A1(n10290), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10289), .ZN(n10294) );
  AOI22_X1 U11602 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10299) );
  NOR2_X1 U11603 ( .A1(n12209), .A2(n10864), .ZN(n12229) );
  AOI21_X1 U11604 ( .B1(n18539), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12763), .ZN(n12769) );
  AND2_X1 U11605 ( .A1(n13691), .A2(n13690), .ZN(n12763) );
  NOR2_X1 U11606 ( .A1(n12742), .A2(n12740), .ZN(n12838) );
  NOR2_X1 U11607 ( .A1(n12744), .A2(n12743), .ZN(n15669) );
  INV_X1 U11608 ( .A(n17619), .ZN(n9839) );
  AND2_X1 U11609 ( .A1(n9675), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9960) );
  NAND2_X1 U11610 ( .A1(n16500), .A2(n16461), .ZN(n16444) );
  NAND2_X1 U11611 ( .A1(n17986), .A2(n9809), .ZN(n15922) );
  NOR2_X1 U11612 ( .A1(n17948), .A2(n9810), .ZN(n9809) );
  NAND2_X1 U11613 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9810) );
  OAI21_X1 U11614 ( .B1(n15905), .B2(n15907), .A(n17849), .ZN(n15911) );
  NOR2_X1 U11615 ( .A1(n17875), .A2(n15855), .ZN(n15858) );
  NOR2_X1 U11616 ( .A1(n17906), .A2(n15846), .ZN(n15847) );
  XNOR2_X1 U11617 ( .A(n15840), .B(n9814), .ZN(n15843) );
  INV_X1 U11618 ( .A(n17459), .ZN(n9814) );
  AND2_X1 U11619 ( .A1(n13997), .A2(n13996), .ZN(n14299) );
  AND2_X1 U11620 ( .A1(n13427), .A2(n13426), .ZN(n13429) );
  INV_X1 U11621 ( .A(n20057), .ZN(n13235) );
  INV_X1 U11622 ( .A(n20241), .ZN(n20242) );
  INV_X1 U11623 ( .A(n11936), .ZN(n11942) );
  AND2_X1 U11624 ( .A1(n20870), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11941) );
  AND2_X1 U11625 ( .A1(n10196), .A2(n10197), .ZN(n10195) );
  INV_X1 U11626 ( .A(n14100), .ZN(n10196) );
  NAND2_X1 U11627 ( .A1(n11748), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11804) );
  NAND2_X1 U11628 ( .A1(n11618), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11663) );
  OR2_X1 U11629 ( .A1(n13231), .A2(n20057), .ZN(n13036) );
  NOR2_X1 U11630 ( .A1(n14456), .A2(n14678), .ZN(n9830) );
  NAND2_X1 U11631 ( .A1(n10050), .A2(n10048), .ZN(n14085) );
  NOR2_X1 U11632 ( .A1(n10049), .A2(n14102), .ZN(n10048) );
  INV_X1 U11633 ( .A(n14086), .ZN(n10049) );
  AND2_X1 U11634 ( .A1(n10050), .A2(n10047), .ZN(n14101) );
  INV_X1 U11635 ( .A(n14102), .ZN(n10047) );
  NAND2_X1 U11636 ( .A1(n14504), .A2(n14453), .ZN(n14455) );
  INV_X1 U11637 ( .A(n14512), .ZN(n10035) );
  NAND2_X1 U11638 ( .A1(n10033), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14518) );
  OR2_X1 U11639 ( .A1(n9823), .A2(n14601), .ZN(n10033) );
  NAND2_X1 U11640 ( .A1(n9702), .A2(n14299), .ZN(n14298) );
  NAND2_X1 U11641 ( .A1(n9825), .A2(n9828), .ZN(n14623) );
  NAND2_X1 U11642 ( .A1(n9829), .A2(n16228), .ZN(n9828) );
  NAND2_X1 U11643 ( .A1(n16235), .A2(n13547), .ZN(n13587) );
  NAND2_X1 U11644 ( .A1(n12014), .A2(n14043), .ZN(n11041) );
  OR2_X2 U11645 ( .A1(n11187), .A2(n11188), .ZN(n11236) );
  INV_X1 U11646 ( .A(n11020), .ZN(n10055) );
  NOR2_X1 U11647 ( .A1(n20250), .A2(n20413), .ZN(n20598) );
  NAND2_X1 U11648 ( .A1(n20868), .A2(n20245), .ZN(n20413) );
  INV_X1 U11649 ( .A(n20445), .ZN(n20694) );
  NAND2_X1 U11650 ( .A1(n10995), .A2(n9709), .ZN(n9903) );
  NOR2_X1 U11651 ( .A1(n13368), .A2(n13370), .ZN(n20735) );
  AND2_X1 U11652 ( .A1(n10574), .A2(n10573), .ZN(n12235) );
  XNOR2_X1 U11653 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U11654 ( .A1(n10141), .A2(n10140), .ZN(n12207) );
  NAND2_X1 U11655 ( .A1(n12221), .A2(n12225), .ZN(n10140) );
  OR2_X1 U11656 ( .A1(n12118), .A2(n12221), .ZN(n10141) );
  AOI21_X1 U11657 ( .B1(n9661), .B2(n12402), .A(n12401), .ZN(n12403) );
  INV_X1 U11658 ( .A(n18983), .ZN(n10023) );
  AND2_X1 U11659 ( .A1(n16384), .A2(n19274), .ZN(n12613) );
  NAND2_X1 U11660 ( .A1(n13380), .A2(n13444), .ZN(n10105) );
  NOR2_X1 U11661 ( .A1(n10105), .A2(n10104), .ZN(n10103) );
  INV_X1 U11662 ( .A(n13477), .ZN(n10104) );
  NAND2_X1 U11663 ( .A1(n12997), .A2(n12995), .ZN(n10099) );
  OR2_X1 U11664 ( .A1(n12944), .A2(n12943), .ZN(n12945) );
  NAND2_X1 U11665 ( .A1(n9758), .A2(n15047), .ZN(n10168) );
  AND2_X1 U11666 ( .A1(n9743), .A2(n14984), .ZN(n10106) );
  AND2_X1 U11667 ( .A1(n10829), .A2(n10828), .ZN(n14921) );
  AND2_X1 U11668 ( .A1(n9660), .A2(n19422), .ZN(n12716) );
  INV_X1 U11669 ( .A(n12224), .ZN(n10392) );
  OR2_X1 U11670 ( .A1(n10275), .A2(n10274), .ZN(n10277) );
  NAND2_X1 U11671 ( .A1(n15297), .A2(n9701), .ZN(n9785) );
  AND2_X1 U11672 ( .A1(n10490), .A2(n10489), .ZN(n13149) );
  NAND2_X1 U11673 ( .A1(n10084), .A2(n10082), .ZN(n13148) );
  INV_X1 U11674 ( .A(n10083), .ZN(n10082) );
  NAND2_X1 U11675 ( .A1(n9955), .A2(n10207), .ZN(n9954) );
  INV_X1 U11676 ( .A(n9956), .ZN(n9955) );
  NAND2_X1 U11677 ( .A1(n15152), .A2(n10156), .ZN(n10155) );
  AND2_X1 U11678 ( .A1(n10154), .A2(n15153), .ZN(n9869) );
  INV_X1 U11679 ( .A(n12368), .ZN(n10156) );
  NOR2_X1 U11680 ( .A1(n15171), .A2(n9950), .ZN(n9949) );
  INV_X1 U11681 ( .A(n15167), .ZN(n9950) );
  NAND2_X1 U11682 ( .A1(n9673), .A2(n15170), .ZN(n9951) );
  NOR2_X1 U11683 ( .A1(n9673), .A2(n9948), .ZN(n9947) );
  INV_X1 U11684 ( .A(n9949), .ZN(n9948) );
  OAI22_X1 U11685 ( .A1(n9951), .A2(n9949), .B1(n9673), .B2(n15170), .ZN(n9946) );
  INV_X1 U11686 ( .A(n9932), .ZN(n9930) );
  AOI21_X1 U11687 ( .B1(n9932), .B2(n9929), .A(n9928), .ZN(n9927) );
  INV_X1 U11688 ( .A(n15234), .ZN(n9928) );
  INV_X1 U11689 ( .A(n9937), .ZN(n9929) );
  NAND2_X1 U11690 ( .A1(n9935), .A2(n15242), .ZN(n9934) );
  OR2_X1 U11691 ( .A1(n15163), .A2(n9936), .ZN(n9935) );
  NAND2_X1 U11692 ( .A1(n15162), .A2(n15254), .ZN(n9936) );
  NAND2_X1 U11693 ( .A1(n15256), .A2(n9937), .ZN(n9933) );
  NAND2_X1 U11694 ( .A1(n9872), .A2(n9871), .ZN(n12329) );
  NOR2_X1 U11695 ( .A1(n10160), .A2(n15275), .ZN(n10159) );
  NAND2_X1 U11696 ( .A1(n13125), .A2(n13124), .ZN(n13212) );
  INV_X1 U11697 ( .A(n13652), .ZN(n9794) );
  CLKBUF_X1 U11698 ( .A(n10577), .Z(n10578) );
  AND2_X1 U11699 ( .A1(n9991), .A2(n12287), .ZN(n9990) );
  OR2_X1 U11700 ( .A1(n12286), .A2(n9992), .ZN(n9991) );
  NAND2_X1 U11701 ( .A1(n13529), .A2(n12433), .ZN(n9992) );
  INV_X1 U11702 ( .A(n13529), .ZN(n9995) );
  INV_X1 U11703 ( .A(n12109), .ZN(n12107) );
  NAND2_X1 U11704 ( .A1(n13972), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12253) );
  AND2_X1 U11705 ( .A1(n10375), .A2(n12215), .ZN(n10377) );
  AND2_X1 U11706 ( .A1(n10398), .A2(n12237), .ZN(n10375) );
  NAND2_X1 U11707 ( .A1(n19630), .A2(n20037), .ZN(n19572) );
  NAND2_X1 U11708 ( .A1(n20019), .A2(n20026), .ZN(n19662) );
  NAND2_X1 U11709 ( .A1(n20019), .A2(n20028), .ZN(n20007) );
  OR2_X1 U11710 ( .A1(n19630), .A2(n19629), .ZN(n19815) );
  OR2_X1 U11711 ( .A1(n19630), .A2(n20037), .ZN(n19789) );
  NAND2_X1 U11712 ( .A1(n16676), .A2(n10223), .ZN(n16666) );
  INV_X1 U11713 ( .A(n15648), .ZN(n17252) );
  NOR2_X1 U11714 ( .A1(n9849), .A2(n9848), .ZN(n10126) );
  OAI22_X1 U11715 ( .A1(n18717), .A2(n15741), .B1(n13684), .B2(n12837), .ZN(
        n15979) );
  NOR2_X1 U11716 ( .A1(n13687), .A2(n9887), .ZN(n9886) );
  NAND2_X1 U11717 ( .A1(n18301), .A2(n9888), .ZN(n9887) );
  NOR2_X1 U11718 ( .A1(n18925), .A2(n9891), .ZN(n17511) );
  OR2_X1 U11719 ( .A1(n17728), .A2(n17727), .ZN(n17704) );
  AND2_X1 U11720 ( .A1(n9864), .A2(n15905), .ZN(n17755) );
  NOR2_X1 U11721 ( .A1(n16436), .A2(n9963), .ZN(n9962) );
  INV_X1 U11722 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9963) );
  NAND2_X1 U11723 ( .A1(n16435), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16436) );
  INV_X1 U11724 ( .A(n17828), .ZN(n16435) );
  INV_X1 U11725 ( .A(n17742), .ZN(n16819) );
  NOR2_X2 U11726 ( .A1(n17888), .A2(n17887), .ZN(n17878) );
  NAND2_X1 U11727 ( .A1(n17909), .A2(n15877), .ZN(n17899) );
  NAND2_X1 U11728 ( .A1(n16445), .A2(n16447), .ZN(n10125) );
  AOI21_X1 U11729 ( .B1(n17849), .B2(n16448), .A(n9766), .ZN(n10124) );
  AND2_X1 U11730 ( .A1(n10123), .A2(n10121), .ZN(n10120) );
  NOR2_X1 U11731 ( .A1(n10122), .A2(n16489), .ZN(n10121) );
  OR2_X1 U11732 ( .A1(n17833), .A2(n18887), .ZN(n10123) );
  NOR2_X1 U11733 ( .A1(n17849), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10122) );
  NAND2_X1 U11734 ( .A1(n15965), .A2(n16460), .ZN(n16445) );
  NOR2_X1 U11735 ( .A1(n17607), .A2(n15919), .ZN(n15920) );
  OR2_X1 U11736 ( .A1(n15918), .A2(n15917), .ZN(n15919) );
  INV_X1 U11737 ( .A(n15922), .ZN(n17951) );
  NOR2_X1 U11738 ( .A1(n17641), .A2(n18077), .ZN(n17981) );
  NOR2_X1 U11739 ( .A1(n18075), .A2(n17641), .ZN(n17986) );
  NAND2_X1 U11740 ( .A1(n9863), .A2(n15905), .ZN(n9864) );
  AND2_X1 U11741 ( .A1(n18125), .A2(n17833), .ZN(n9863) );
  OAI21_X1 U11742 ( .B1(n17882), .B2(n9838), .A(n9836), .ZN(n17870) );
  AND2_X1 U11743 ( .A1(n9837), .A2(n17872), .ZN(n9836) );
  OR2_X1 U11744 ( .A1(n18739), .A2(n12744), .ZN(n10230) );
  NOR2_X2 U11745 ( .A1(n12751), .A2(n12750), .ZN(n18281) );
  INV_X1 U11746 ( .A(n11195), .ZN(n11196) );
  CLKBUF_X1 U11747 ( .A(n13161), .Z(n13162) );
  AND2_X1 U11748 ( .A1(n10010), .A2(n19145), .ZN(n10285) );
  OR2_X1 U11749 ( .A1(n14861), .A2(n10011), .ZN(n10010) );
  INV_X1 U11750 ( .A(n10012), .ZN(n10011) );
  CLKBUF_X1 U11751 ( .A(n10267), .Z(n19145) );
  INV_X1 U11752 ( .A(n20037), .ZN(n19629) );
  OR2_X1 U11753 ( .A1(n12546), .A2(n12545), .ZN(n14938) );
  OR2_X1 U11754 ( .A1(n10759), .A2(n10758), .ZN(n13130) );
  INV_X1 U11755 ( .A(n15025), .ZN(n15012) );
  OR2_X1 U11756 ( .A1(n15015), .A2(n12711), .ZN(n15025) );
  NOR2_X1 U11757 ( .A1(n14945), .A2(n10112), .ZN(n15040) );
  OR2_X1 U11758 ( .A1(n15336), .A2(n19215), .ZN(n10110) );
  AND2_X1 U11759 ( .A1(n13982), .A2(n19377), .ZN(n19208) );
  INV_X1 U11760 ( .A(n19216), .ZN(n19269) );
  OR2_X1 U11761 ( .A1(n18958), .A2(n10598), .ZN(n16325) );
  XNOR2_X1 U11762 ( .A(n9865), .B(n9707), .ZN(n10114) );
  XNOR2_X1 U11763 ( .A(n12546), .B(n12439), .ZN(n15315) );
  AND2_X1 U11764 ( .A1(n12563), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10072) );
  XNOR2_X1 U11765 ( .A(n12580), .B(n12579), .ZN(n15334) );
  AND2_X1 U11766 ( .A1(n15394), .A2(n12504), .ZN(n15366) );
  INV_X1 U11767 ( .A(n16371), .ZN(n19364) );
  INV_X1 U11768 ( .A(n15597), .ZN(n19361) );
  INV_X1 U11769 ( .A(n12039), .ZN(n9798) );
  OR2_X1 U11770 ( .A1(n12477), .A2(n12448), .ZN(n15589) );
  OR2_X1 U11771 ( .A1(n12477), .A2(n20045), .ZN(n15597) );
  INV_X1 U11772 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20035) );
  INV_X1 U11773 ( .A(n20028), .ZN(n20026) );
  OR2_X1 U11774 ( .A1(n19789), .A2(n19662), .ZN(n19696) );
  INV_X1 U11775 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19926) );
  NAND2_X1 U11776 ( .A1(n9967), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9966) );
  OR2_X1 U11777 ( .A1(n16668), .A2(n17026), .ZN(n9967) );
  OR2_X1 U11778 ( .A1(n16682), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9965) );
  XNOR2_X1 U11779 ( .A(n16666), .B(n9969), .ZN(n9968) );
  INV_X1 U11780 ( .A(n16667), .ZN(n9969) );
  NAND2_X1 U11781 ( .A1(n18766), .A2(n16640), .ZN(n17018) );
  NAND2_X1 U11782 ( .A1(n17027), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17014) );
  INV_X1 U11783 ( .A(n16997), .ZN(n17025) );
  NOR2_X1 U11784 ( .A1(n9885), .A2(n9884), .ZN(n9883) );
  AOI211_X1 U11785 ( .C1(n17035), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n12791), .B(n12790), .ZN(n12792) );
  INV_X1 U11786 ( .A(n12794), .ZN(n9884) );
  NAND2_X1 U11787 ( .A1(n17356), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17355) );
  INV_X1 U11788 ( .A(n17466), .ZN(n17463) );
  NOR2_X2 U11789 ( .A1(n17704), .A2(n17706), .ZN(n17686) );
  INV_X1 U11790 ( .A(n9805), .ZN(n17962) );
  NAND2_X1 U11791 ( .A1(n17672), .A2(n10113), .ZN(n17645) );
  AND2_X1 U11792 ( .A1(n12069), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U11793 ( .A1(n10914), .A2(n20868), .ZN(n10065) );
  INV_X1 U11794 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11033) );
  INV_X1 U11795 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11903) );
  INV_X1 U11796 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11672) );
  NOR2_X1 U11797 ( .A1(n10901), .A2(n20868), .ZN(n9898) );
  INV_X1 U11798 ( .A(n14481), .ZN(n10056) );
  INV_X1 U11799 ( .A(n11338), .ZN(n11339) );
  NAND2_X1 U11800 ( .A1(n11268), .A2(n11267), .ZN(n11275) );
  NOR2_X1 U11801 ( .A1(n12960), .A2(n11052), .ZN(n11073) );
  AND2_X1 U11802 ( .A1(n13238), .A2(n14434), .ZN(n11148) );
  NAND2_X1 U11803 ( .A1(n13226), .A2(n9902), .ZN(n12952) );
  NAND2_X1 U11804 ( .A1(n13113), .A2(n11045), .ZN(n12954) );
  AND2_X1 U11805 ( .A1(n11047), .A2(n20246), .ZN(n11217) );
  INV_X1 U11806 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11701) );
  INV_X1 U11807 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11694) );
  INV_X1 U11808 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11695) );
  OR2_X1 U11809 ( .A1(n10952), .A2(n11033), .ZN(n11034) );
  NOR2_X1 U11810 ( .A1(n10901), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10902) );
  AOI21_X1 U11811 ( .B1(n10351), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n10357), .ZN(n10358) );
  NAND2_X1 U11812 ( .A1(n10005), .A2(n9880), .ZN(n12422) );
  INV_X1 U11813 ( .A(n12413), .ZN(n12414) );
  OAI21_X1 U11814 ( .B1(n12575), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15120), .ZN(n12413) );
  NOR2_X1 U11815 ( .A1(n10002), .A2(n10001), .ZN(n10000) );
  INV_X1 U11816 ( .A(n12394), .ZN(n10002) );
  INV_X1 U11817 ( .A(n9748), .ZN(n10001) );
  NAND2_X1 U11818 ( .A1(n9873), .A2(n10218), .ZN(n10152) );
  NOR2_X1 U11819 ( .A1(n12138), .A2(n9874), .ZN(n9873) );
  AOI22_X1 U11820 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12141), .B1(
        n12151), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12096) );
  AND2_X1 U11821 ( .A1(n12153), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12100) );
  AOI22_X1 U11822 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19859), .B1(
        n12141), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12080) );
  NOR2_X1 U11823 ( .A1(n12135), .A2(n12046), .ZN(n12050) );
  NAND2_X1 U11824 ( .A1(n10139), .A2(n10138), .ZN(n12280) );
  NAND2_X1 U11825 ( .A1(n9660), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10138) );
  NAND2_X1 U11826 ( .A1(n12207), .A2(n10869), .ZN(n10139) );
  NAND2_X1 U11827 ( .A1(n10412), .A2(n10393), .ZN(n12242) );
  INV_X1 U11828 ( .A(n12074), .ZN(n12069) );
  AND2_X1 U11829 ( .A1(n10586), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10369) );
  NAND2_X1 U11830 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10127) );
  NOR2_X1 U11831 ( .A1(n12744), .A2(n17012), .ZN(n15795) );
  NAND2_X1 U11832 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12745) );
  NAND2_X1 U11833 ( .A1(n17464), .A2(n15985), .ZN(n15840) );
  INV_X1 U11834 ( .A(n14272), .ZN(n10185) );
  INV_X1 U11835 ( .A(n14743), .ZN(n9910) );
  INV_X1 U11836 ( .A(n10036), .ZN(n9907) );
  NOR2_X1 U11837 ( .A1(n9913), .A2(n9910), .ZN(n9909) );
  OR2_X1 U11838 ( .A1(n16112), .A2(n14444), .ZN(n14569) );
  OAI21_X1 U11839 ( .B1(n11182), .B2(n13352), .A(n13032), .ZN(n13282) );
  INV_X1 U11840 ( .A(n20369), .ZN(n11178) );
  NAND2_X1 U11841 ( .A1(n11217), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U11842 ( .A1(n11179), .A2(n11078), .ZN(n11079) );
  OAI211_X1 U11843 ( .C1(n20249), .C2(n13040), .A(n11056), .B(n11055), .ZN(
        n11080) );
  OR2_X1 U11844 ( .A1(n11054), .A2(n12964), .ZN(n11056) );
  OR2_X1 U11845 ( .A1(n11231), .A2(n11230), .ZN(n13499) );
  NOR2_X1 U11846 ( .A1(n11217), .A2(n20868), .ZN(n11989) );
  AND2_X1 U11847 ( .A1(n11955), .A2(n11954), .ZN(n11966) );
  OR2_X1 U11848 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20240), .ZN(
        n11954) );
  OR2_X1 U11849 ( .A1(n11956), .A2(n11953), .ZN(n11955) );
  NAND2_X1 U11850 ( .A1(n11969), .A2(n11043), .ZN(n11020) );
  NAND2_X1 U11851 ( .A1(n11216), .A2(n11215), .ZN(n20406) );
  OR2_X1 U11852 ( .A1(n11054), .A2(n10052), .ZN(n11216) );
  OAI21_X1 U11853 ( .B1(n11845), .B2(n11693), .A(n9901), .ZN(n9900) );
  OAI22_X1 U11854 ( .A1(n11906), .A2(n11692), .B1(n11904), .B2(n11688), .ZN(
        n11012) );
  NAND2_X1 U11855 ( .A1(n11129), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n9901) );
  OAI21_X1 U11856 ( .B1(n11849), .B2(n11386), .A(n9834), .ZN(n10909) );
  NAND2_X1 U11857 ( .A1(n11129), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n9834) );
  AND2_X1 U11858 ( .A1(n11129), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10929) );
  AND2_X1 U11859 ( .A1(n10959), .A2(n10958), .ZN(n10961) );
  NAND3_X1 U11860 ( .A1(n9705), .A2(n10983), .A3(n10982), .ZN(n11040) );
  INV_X1 U11861 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20592) );
  AND2_X1 U11862 ( .A1(n10563), .A2(n10562), .ZN(n10572) );
  INV_X1 U11863 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U11864 ( .A1(n12363), .A2(n14997), .ZN(n12365) );
  NAND2_X1 U11865 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  AND2_X1 U11866 ( .A1(n12324), .A2(n10130), .ZN(n12357) );
  NOR2_X1 U11867 ( .A1(n9765), .A2(n10131), .ZN(n10130) );
  INV_X1 U11868 ( .A(n10872), .ZN(n10131) );
  NAND2_X1 U11869 ( .A1(n12291), .A2(n9682), .ZN(n12313) );
  NAND2_X1 U11870 ( .A1(n13869), .A2(n14965), .ZN(n10093) );
  AND2_X1 U11871 ( .A1(n10172), .A2(n10846), .ZN(n10171) );
  INV_X1 U11872 ( .A(n14890), .ZN(n10172) );
  INV_X1 U11873 ( .A(n14889), .ZN(n10170) );
  AND2_X1 U11874 ( .A1(n13786), .A2(n15018), .ZN(n10108) );
  OR2_X1 U11875 ( .A1(n10709), .A2(n10708), .ZN(n12181) );
  OR2_X1 U11876 ( .A1(n10597), .A2(n10596), .ZN(n12159) );
  AND2_X1 U11877 ( .A1(n9676), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10027) );
  NAND2_X1 U11878 ( .A1(n10250), .A2(n9676), .ZN(n10258) );
  NOR2_X1 U11879 ( .A1(n16331), .A2(n10029), .ZN(n10028) );
  INV_X1 U11880 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U11881 ( .A1(n10084), .A2(n10081), .ZN(n13119) );
  NOR2_X1 U11882 ( .A1(n10481), .A2(n10077), .ZN(n10081) );
  INV_X1 U11883 ( .A(n13149), .ZN(n10078) );
  INV_X1 U11884 ( .A(n12118), .ZN(n12106) );
  XNOR2_X1 U11885 ( .A(n12434), .B(n10879), .ZN(n12430) );
  NOR2_X1 U11886 ( .A1(n10208), .A2(n15329), .ZN(n10207) );
  INV_X1 U11887 ( .A(n10209), .ZN(n10208) );
  NOR2_X1 U11888 ( .A1(n15323), .A2(n15348), .ZN(n10209) );
  NAND2_X1 U11889 ( .A1(n9782), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9956) );
  OR2_X1 U11890 ( .A1(n10157), .A2(n12383), .ZN(n10154) );
  OR2_X1 U11891 ( .A1(n14911), .A2(n9942), .ZN(n12389) );
  AND2_X1 U11892 ( .A1(n15508), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10211) );
  INV_X1 U11893 ( .A(n12319), .ZN(n10160) );
  NOR2_X1 U11894 ( .A1(n12433), .A2(n15604), .ZN(n9941) );
  INV_X1 U11895 ( .A(n12199), .ZN(n12200) );
  OAI21_X1 U11896 ( .B1(n10473), .B2(n13613), .A(n10472), .ZN(n10478) );
  NAND2_X1 U11897 ( .A1(n10461), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10463) );
  NAND2_X1 U11898 ( .A1(n9952), .A2(n10436), .ZN(n10448) );
  NAND2_X1 U11899 ( .A1(n10435), .A2(n10421), .ZN(n9952) );
  NOR2_X1 U11900 ( .A1(n10445), .A2(n10418), .ZN(n12691) );
  NAND2_X1 U11901 ( .A1(n10092), .A2(n10091), .ZN(n10422) );
  AND2_X1 U11902 ( .A1(n12062), .A2(n12068), .ZN(n9919) );
  AND2_X1 U11903 ( .A1(n12060), .A2(n12062), .ZN(n12061) );
  NAND2_X1 U11904 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18909), .ZN(
        n12743) );
  OR2_X1 U11905 ( .A1(n12742), .A2(n12744), .ZN(n12841) );
  INV_X1 U11906 ( .A(n15798), .ZN(n9849) );
  NAND2_X1 U11907 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n15792) );
  OR2_X1 U11908 ( .A1(n18739), .A2(n12745), .ZN(n15827) );
  XOR2_X1 U11909 ( .A(n17444), .B(n15886), .Z(n15887) );
  NOR2_X1 U11910 ( .A1(n17884), .A2(n15851), .ZN(n15853) );
  NAND2_X1 U11911 ( .A1(n15743), .A2(n9893), .ZN(n9892) );
  NAND2_X1 U11912 ( .A1(n13689), .A2(n18281), .ZN(n9893) );
  AOI211_X1 U11913 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n12781), .B(n12780), .ZN(n12782) );
  INV_X1 U11914 ( .A(n13231), .ZN(n13224) );
  AND2_X1 U11915 ( .A1(n14024), .A2(n14023), .ZN(n14275) );
  NOR2_X1 U11916 ( .A1(n11474), .A2(n14606), .ZN(n11497) );
  OR2_X1 U11917 ( .A1(n20949), .A2(n13342), .ZN(n14232) );
  NAND2_X1 U11918 ( .A1(n10040), .A2(n10045), .ZN(n10044) );
  NAND2_X1 U11919 ( .A1(n11248), .A2(n11247), .ZN(n13305) );
  AOI21_X1 U11920 ( .B1(n14464), .B2(n13340), .A(n11940), .ZN(n14077) );
  NAND2_X1 U11921 ( .A1(n11899), .A2(n11898), .ZN(n14090) );
  OR2_X1 U11922 ( .A1(n11804), .A2(n14506), .ZN(n11805) );
  AOI21_X1 U11923 ( .B1(n14502), .B2(n13340), .A(n11829), .ZN(n14111) );
  AND2_X1 U11924 ( .A1(n11747), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11748) );
  INV_X1 U11925 ( .A(n11746), .ZN(n11747) );
  AND2_X1 U11926 ( .A1(n11774), .A2(n11773), .ZN(n14136) );
  OR2_X1 U11927 ( .A1(n14514), .A2(n11935), .ZN(n11774) );
  CLKBUF_X1 U11928 ( .A(n14257), .Z(n14258) );
  NOR2_X1 U11929 ( .A1(n11617), .A2(n14550), .ZN(n11618) );
  OR2_X1 U11930 ( .A1(n16006), .A2(n11935), .ZN(n11640) );
  NOR2_X1 U11931 ( .A1(n11578), .A2(n14562), .ZN(n11579) );
  NAND2_X1 U11932 ( .A1(n11538), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11558) );
  NAND2_X1 U11933 ( .A1(n10191), .A2(n14368), .ZN(n10190) );
  INV_X1 U11934 ( .A(n10193), .ZN(n10191) );
  NOR2_X1 U11935 ( .A1(n11517), .A2(n16057), .ZN(n11538) );
  NAND2_X1 U11936 ( .A1(n11497), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11517) );
  INV_X1 U11937 ( .A(n14194), .ZN(n10192) );
  CLKBUF_X1 U11938 ( .A(n14194), .Z(n14195) );
  NAND2_X1 U11939 ( .A1(n11449), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11474) );
  AND2_X1 U11940 ( .A1(n11406), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11407) );
  NAND2_X1 U11941 ( .A1(n11407), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11429) );
  NOR2_X1 U11942 ( .A1(n11384), .A2(n11383), .ZN(n11406) );
  AND2_X1 U11943 ( .A1(n11405), .A2(n13600), .ZN(n10194) );
  NAND2_X1 U11944 ( .A1(n11365), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11384) );
  INV_X1 U11945 ( .A(n11364), .ZN(n11365) );
  NAND2_X1 U11946 ( .A1(n11344), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11364) );
  AND2_X1 U11947 ( .A1(n11328), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11344) );
  AOI21_X1 U11948 ( .B1(n14410), .B2(n11513), .A(n11335), .ZN(n13537) );
  CLKBUF_X1 U11949 ( .A(n13534), .Z(n13535) );
  AND2_X1 U11950 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11300), .ZN(
        n11301) );
  CLKBUF_X1 U11951 ( .A(n13421), .Z(n13422) );
  NAND2_X1 U11952 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11240) );
  NOR2_X1 U11953 ( .A1(n11240), .A2(n11239), .ZN(n11300) );
  INV_X1 U11954 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11239) );
  AOI21_X1 U11955 ( .B1(n11193), .B2(n11298), .A(n10189), .ZN(n10188) );
  INV_X1 U11956 ( .A(n11211), .ZN(n10189) );
  AND2_X1 U11957 ( .A1(n14479), .A2(n14696), .ZN(n14480) );
  AOI22_X1 U11958 ( .A1(n14450), .A2(n9824), .B1(n9823), .B2(n10057), .ZN(
        n9822) );
  NOR2_X1 U11959 ( .A1(n14153), .A2(n14142), .ZN(n14141) );
  OR2_X1 U11960 ( .A1(n14726), .A2(n14151), .ZN(n14153) );
  NAND2_X1 U11961 ( .A1(n14724), .A2(n14723), .ZN(n14726) );
  NAND2_X1 U11962 ( .A1(n14450), .A2(n14601), .ZN(n14532) );
  OAI21_X1 U11963 ( .B1(n9906), .B2(n14596), .A(n9904), .ZN(n14531) );
  INV_X1 U11964 ( .A(n9905), .ZN(n9904) );
  NAND2_X1 U11965 ( .A1(n9907), .A2(n9909), .ZN(n9906) );
  OAI21_X1 U11966 ( .B1(n9911), .B2(n9910), .A(n14449), .ZN(n9905) );
  AND2_X1 U11967 ( .A1(n16044), .A2(n9772), .ZN(n14268) );
  INV_X1 U11968 ( .A(n14265), .ZN(n10053) );
  NAND2_X1 U11969 ( .A1(n16044), .A2(n9759), .ZN(n14266) );
  NAND2_X1 U11970 ( .A1(n16044), .A2(n9757), .ZN(n14274) );
  AND2_X1 U11971 ( .A1(n13252), .A2(n14785), .ZN(n16171) );
  NAND2_X1 U11972 ( .A1(n16113), .A2(n9908), .ZN(n9912) );
  NOR2_X1 U11973 ( .A1(n10036), .A2(n9913), .ZN(n9908) );
  AND2_X1 U11974 ( .A1(n16044), .A2(n14279), .ZN(n14281) );
  NAND2_X1 U11975 ( .A1(n16113), .A2(n10071), .ZN(n16087) );
  NOR2_X1 U11976 ( .A1(n14570), .A2(n14573), .ZN(n10071) );
  OR2_X1 U11977 ( .A1(n16112), .A2(n14445), .ZN(n14571) );
  AND2_X1 U11978 ( .A1(n14011), .A2(n14010), .ZN(n16052) );
  NAND2_X1 U11979 ( .A1(n10046), .A2(n9744), .ZN(n14213) );
  INV_X1 U11980 ( .A(n14298), .ZN(n10046) );
  NAND2_X1 U11981 ( .A1(n16112), .A2(n14437), .ZN(n14628) );
  NAND2_X1 U11982 ( .A1(n16121), .A2(n14426), .ZN(n9827) );
  AND2_X1 U11983 ( .A1(n13585), .A2(n13584), .ZN(n13588) );
  AND2_X1 U11984 ( .A1(n13545), .A2(n13544), .ZN(n16234) );
  NAND2_X1 U11985 ( .A1(n13439), .A2(n10045), .ZN(n10041) );
  NAND2_X1 U11986 ( .A1(n16255), .A2(n20868), .ZN(n13040) );
  AND2_X1 U11987 ( .A1(n14783), .A2(n14788), .ZN(n16197) );
  INV_X1 U11988 ( .A(n20229), .ZN(n16175) );
  NOR2_X1 U11989 ( .A1(n11063), .A2(n11020), .ZN(n12722) );
  AND2_X2 U11990 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12963) );
  AND4_X1 U11991 ( .A1(n12989), .A2(n12988), .A3(n12987), .A4(n13020), .ZN(
        n15939) );
  OR2_X1 U11992 ( .A1(n9665), .A2(n20244), .ZN(n20405) );
  AND2_X1 U11993 ( .A1(n20372), .A2(n20797), .ZN(n20374) );
  AOI21_X1 U11994 ( .B1(n19145), .B2(n14862), .A(n14852), .ZN(n10012) );
  OR2_X1 U11995 ( .A1(n12599), .A2(n15107), .ZN(n12597) );
  NAND2_X1 U11996 ( .A1(n10877), .A2(n10876), .ZN(n12415) );
  NAND2_X1 U11997 ( .A1(n12336), .A2(n10142), .ZN(n12412) );
  NOR2_X1 U11998 ( .A1(n12391), .A2(n10143), .ZN(n10142) );
  NAND2_X1 U11999 ( .A1(n12385), .A2(n9692), .ZN(n10143) );
  AND2_X1 U12000 ( .A1(n12324), .A2(n10132), .ZN(n12349) );
  NOR2_X1 U12001 ( .A1(n9765), .A2(n10133), .ZN(n10132) );
  NAND2_X1 U12002 ( .A1(n10873), .A2(n10872), .ZN(n10133) );
  NAND2_X1 U12003 ( .A1(n12349), .A2(n13648), .ZN(n12346) );
  INV_X1 U12004 ( .A(n10511), .ZN(n12441) );
  AND2_X1 U12005 ( .A1(n12603), .A2(n12567), .ZN(n12568) );
  INV_X1 U12006 ( .A(n12556), .ZN(n14867) );
  NAND2_X1 U12007 ( .A1(n13930), .A2(n13928), .ZN(n14947) );
  NAND2_X1 U12008 ( .A1(n14959), .A2(n14961), .ZN(n14960) );
  NAND2_X1 U12009 ( .A1(n10170), .A2(n10171), .ZN(n15062) );
  XNOR2_X1 U12010 ( .A(n13847), .B(n13868), .ZN(n14975) );
  AND2_X1 U12011 ( .A1(n9685), .A2(n9776), .ZN(n10175) );
  BUF_X1 U12012 ( .A(n13847), .Z(n14979) );
  NAND2_X1 U12013 ( .A1(n15445), .A2(n9685), .ZN(n15422) );
  AND2_X1 U12014 ( .A1(n10832), .A2(n10831), .ZN(n15093) );
  INV_X1 U12015 ( .A(n14921), .ZN(n10830) );
  NAND2_X1 U12016 ( .A1(n10103), .A2(n13484), .ZN(n10102) );
  OR3_X1 U12017 ( .A1(n13557), .A2(n15566), .A3(n15581), .ZN(n15568) );
  OR2_X1 U12018 ( .A1(n13557), .A2(n15581), .ZN(n15584) );
  INV_X1 U12019 ( .A(n18956), .ZN(n19274) );
  OR2_X1 U12020 ( .A1(n12997), .A2(n12996), .ZN(n10100) );
  AND2_X1 U12021 ( .A1(n19239), .A2(n12717), .ZN(n13982) );
  NAND2_X1 U12022 ( .A1(n10613), .A2(n10825), .ZN(n10616) );
  OAI211_X1 U12023 ( .C1(n12452), .C2(n10440), .A(n10618), .B(n10617), .ZN(
        n12712) );
  INV_X1 U12024 ( .A(n12234), .ZN(n19281) );
  INV_X1 U12025 ( .A(n12595), .ZN(n19377) );
  XNOR2_X1 U12026 ( .A(n10241), .B(n21100), .ZN(n12529) );
  NAND2_X1 U12027 ( .A1(n10283), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10241) );
  AND2_X1 U12028 ( .A1(n10279), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10283) );
  NOR2_X1 U12029 ( .A1(n10277), .A2(n15105), .ZN(n10280) );
  AND2_X1 U12030 ( .A1(n9689), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10024) );
  AND2_X1 U12031 ( .A1(n9686), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10014) );
  NOR2_X1 U12032 ( .A1(n15022), .A2(n15006), .ZN(n15008) );
  AND2_X1 U12033 ( .A1(n10211), .A2(n12487), .ZN(n10210) );
  NAND2_X1 U12034 ( .A1(n10264), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10265) );
  AND2_X1 U12035 ( .A1(n10245), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10264) );
  NOR2_X1 U12036 ( .A1(n13486), .A2(n13485), .ZN(n13644) );
  INV_X1 U12037 ( .A(n13445), .ZN(n10087) );
  NAND2_X1 U12038 ( .A1(n10248), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10262) );
  NAND2_X1 U12039 ( .A1(n13125), .A2(n9677), .ZN(n13446) );
  NAND2_X1 U12040 ( .A1(n15287), .A2(n12319), .ZN(n15273) );
  AND2_X1 U12041 ( .A1(n13194), .A2(n13202), .ZN(n13203) );
  NAND2_X1 U12042 ( .A1(n10250), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10256) );
  NAND2_X1 U12043 ( .A1(n15297), .A2(n10206), .ZN(n10203) );
  NAND2_X1 U12044 ( .A1(n10205), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10204) );
  NOR2_X1 U12045 ( .A1(n13525), .A2(n10018), .ZN(n10017) );
  NOR2_X1 U12046 ( .A1(n10083), .A2(n13149), .ZN(n10080) );
  NAND2_X1 U12047 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U12048 ( .A1(n16279), .A2(n19369), .ZN(n10167) );
  NOR2_X1 U12049 ( .A1(n9868), .A2(n9867), .ZN(n9866) );
  INV_X1 U12050 ( .A(n12541), .ZN(n9867) );
  INV_X1 U12051 ( .A(n12521), .ZN(n9868) );
  NAND2_X1 U12052 ( .A1(n12542), .A2(n12540), .ZN(n12519) );
  OR3_X1 U12053 ( .A1(n12431), .A2(n9942), .A3(n12506), .ZN(n12521) );
  NOR2_X1 U12054 ( .A1(n14864), .A2(n9942), .ZN(n12578) );
  NOR2_X1 U12055 ( .A1(n12601), .A2(n9942), .ZN(n12575) );
  NAND2_X1 U12056 ( .A1(n9997), .A2(n9996), .ZN(n12577) );
  AND2_X1 U12057 ( .A1(n9711), .A2(n15120), .ZN(n10003) );
  NAND2_X1 U12058 ( .A1(n14904), .A2(n9769), .ZN(n14953) );
  INV_X1 U12059 ( .A(n14950), .ZN(n10088) );
  NOR2_X1 U12060 ( .A1(n14953), .A2(n12602), .ZN(n12603) );
  OAI21_X1 U12061 ( .B1(n16291), .B2(n9942), .A(n15348), .ZN(n12405) );
  NAND2_X1 U12062 ( .A1(n14904), .A2(n9760), .ZN(n14951) );
  NAND2_X1 U12063 ( .A1(n10005), .A2(n15133), .ZN(n15123) );
  AND2_X1 U12064 ( .A1(n14904), .A2(n14887), .ZN(n14969) );
  OR2_X1 U12065 ( .A1(n15006), .A2(n14985), .ZN(n10073) );
  OR2_X1 U12066 ( .A1(n15581), .A2(n15551), .ZN(n10176) );
  INV_X1 U12067 ( .A(n9789), .ZN(n9786) );
  CLKBUF_X1 U12068 ( .A(n13557), .Z(n15582) );
  NAND2_X1 U12069 ( .A1(n9940), .A2(n19131), .ZN(n12303) );
  AOI21_X1 U12070 ( .B1(n9669), .B2(n9994), .A(n9691), .ZN(n9987) );
  NAND2_X1 U12071 ( .A1(n12127), .A2(n9669), .ZN(n9793) );
  NAND2_X1 U12072 ( .A1(n13608), .A2(n13656), .ZN(n9796) );
  NAND2_X1 U12073 ( .A1(n10163), .A2(n9720), .ZN(n10164) );
  INV_X1 U12074 ( .A(n13615), .ZN(n10165) );
  OR2_X1 U12075 ( .A1(n12726), .A2(n12886), .ZN(n12887) );
  NAND2_X1 U12076 ( .A1(n10163), .A2(n13461), .ZN(n10166) );
  NAND2_X1 U12077 ( .A1(n12686), .A2(n19632), .ZN(n12938) );
  AND2_X1 U12078 ( .A1(n12060), .A2(n12054), .ZN(n12052) );
  NAND2_X1 U12079 ( .A1(n9975), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9974) );
  NAND2_X1 U12080 ( .A1(n9973), .A2(n10383), .ZN(n9972) );
  NAND2_X1 U12081 ( .A1(n10384), .A2(n10383), .ZN(n10391) );
  NAND2_X1 U12082 ( .A1(n10389), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10390) );
  NAND2_X2 U12083 ( .A1(n10312), .A2(n10311), .ZN(n10407) );
  NAND2_X1 U12084 ( .A1(n10220), .A2(n10221), .ZN(n10312) );
  OAI21_X1 U12085 ( .B1(n10324), .B2(n10323), .A(n10383), .ZN(n10325) );
  NAND2_X1 U12086 ( .A1(n10317), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10326) );
  NAND2_X2 U12087 ( .A1(n10301), .A2(n10300), .ZN(n12237) );
  NAND2_X1 U12088 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19868), .ZN(n19401) );
  CLKBUF_X1 U12089 ( .A(n10584), .Z(n10869) );
  NOR2_X2 U12090 ( .A1(n19377), .A2(n19376), .ZN(n19416) );
  NOR2_X2 U12091 ( .A1(n19375), .A2(n19376), .ZN(n19415) );
  AND2_X1 U12092 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19858), .ZN(
        n12935) );
  OR2_X1 U12093 ( .A1(n20019), .A2(n20026), .ZN(n19814) );
  INV_X1 U12094 ( .A(n19401), .ZN(n19421) );
  AND2_X1 U12095 ( .A1(n10576), .A2(n10575), .ZN(n16384) );
  NOR2_X1 U12096 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16419) );
  NOR2_X1 U12097 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18909), .ZN(
        n13690) );
  AOI21_X1 U12098 ( .B1(n12769), .B2(n12768), .A(n12767), .ZN(n15894) );
  AND2_X1 U12099 ( .A1(n12770), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12772) );
  INV_X1 U12100 ( .A(n15743), .ZN(n18710) );
  AOI22_X1 U12101 ( .A1(n16432), .A2(n18716), .B1(n18714), .B2(n16499), .ZN(
        n18720) );
  AND2_X1 U12102 ( .A1(n16709), .A2(n16641), .ZN(n16694) );
  NOR2_X1 U12103 ( .A1(n16694), .A2(n16695), .ZN(n16693) );
  AND2_X1 U12104 ( .A1(n16733), .A2(n16641), .ZN(n16720) );
  OR2_X1 U12105 ( .A1(n16765), .A2(n17679), .ZN(n16763) );
  AND2_X1 U12106 ( .A1(n16784), .A2(n16641), .ZN(n16774) );
  NOR2_X1 U12107 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16806), .ZN(n16794) );
  NAND2_X1 U12108 ( .A1(n16641), .A2(n9747), .ZN(n9971) );
  NOR2_X1 U12109 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16831), .ZN(n16816) );
  NOR2_X1 U12110 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16852), .ZN(n16840) );
  INV_X1 U12111 ( .A(n12793), .ZN(n9885) );
  AOI211_X1 U12112 ( .C1(n15834), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12822), .B(n12821), .ZN(n12823) );
  AND2_X1 U12113 ( .A1(n13694), .A2(n18928), .ZN(n17473) );
  NOR2_X1 U12114 ( .A1(n16439), .A2(n17933), .ZN(n16452) );
  AND2_X1 U12115 ( .A1(n17686), .A2(n9736), .ZN(n17609) );
  INV_X1 U12116 ( .A(n17624), .ZN(n9959) );
  NAND2_X1 U12117 ( .A1(n17686), .A2(n9960), .ZN(n17623) );
  NOR3_X1 U12118 ( .A1(n16647), .A2(n17676), .A3(n17662), .ZN(n17621) );
  NOR2_X1 U12119 ( .A1(n18082), .A2(n18125), .ZN(n17772) );
  INV_X1 U12120 ( .A(n9811), .ZN(n17846) );
  AND2_X1 U12121 ( .A1(n15862), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9812) );
  NAND2_X1 U12122 ( .A1(n17878), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16919) );
  XNOR2_X1 U12123 ( .A(n15843), .B(n18222), .ZN(n17918) );
  NAND2_X1 U12124 ( .A1(n15920), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17597) );
  NAND2_X1 U12125 ( .A1(n9847), .A2(n9842), .ZN(n9841) );
  AND2_X1 U12126 ( .A1(n10113), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9842) );
  AND2_X1 U12127 ( .A1(n15916), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10113) );
  INV_X1 U12128 ( .A(n17736), .ZN(n18043) );
  NAND2_X1 U12129 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17772), .ZN(
        n18077) );
  AND2_X1 U12130 ( .A1(n9813), .A2(n18067), .ZN(n17771) );
  INV_X1 U12131 ( .A(n13696), .ZN(n15746) );
  INV_X1 U12132 ( .A(n9892), .ZN(n18729) );
  INV_X1 U12133 ( .A(n10129), .ZN(n10128) );
  NOR2_X1 U12134 ( .A1(n15901), .A2(n15865), .ZN(n16499) );
  XNOR2_X1 U12135 ( .A(n15853), .B(n15854), .ZN(n17876) );
  NOR2_X1 U12136 ( .A1(n17876), .A2(n18186), .ZN(n17875) );
  NOR2_X1 U12137 ( .A1(n17894), .A2(n15849), .ZN(n17886) );
  NOR2_X1 U12138 ( .A1(n17886), .A2(n17885), .ZN(n17884) );
  INV_X1 U12139 ( .A(n15882), .ZN(n15883) );
  XNOR2_X1 U12140 ( .A(n15847), .B(n18209), .ZN(n17896) );
  NOR2_X1 U12141 ( .A1(n17896), .A2(n17895), .ZN(n17894) );
  XNOR2_X1 U12142 ( .A(n15876), .B(n15875), .ZN(n17910) );
  NAND2_X1 U12143 ( .A1(n17910), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17909) );
  NAND2_X1 U12144 ( .A1(n15871), .A2(n17929), .ZN(n17921) );
  XNOR2_X1 U12145 ( .A(n15870), .B(n9850), .ZN(n17930) );
  NAND2_X1 U12146 ( .A1(n17930), .A2(n9674), .ZN(n17929) );
  INV_X1 U12147 ( .A(n15985), .ZN(n17937) );
  INV_X1 U12148 ( .A(n18718), .ZN(n18742) );
  NOR2_X1 U12149 ( .A1(n9892), .A2(n15747), .ZN(n10213) );
  INV_X1 U12150 ( .A(n18372), .ZN(n18621) );
  NOR2_X1 U12151 ( .A1(n12814), .A2(n12813), .ZN(n18293) );
  INV_X1 U12152 ( .A(n19377), .ZN(n19375) );
  OR2_X1 U12153 ( .A1(n12864), .A2(n20057), .ZN(n12858) );
  INV_X1 U12154 ( .A(n20143), .ZN(n20117) );
  NAND2_X1 U12155 ( .A1(n13359), .A2(n13356), .ZN(n20102) );
  AND2_X1 U12156 ( .A1(n13359), .A2(n13358), .ZN(n20145) );
  AND2_X1 U12157 ( .A1(n13359), .A2(n13354), .ZN(n20143) );
  INV_X1 U12158 ( .A(n16076), .ZN(n20156) );
  AND2_X1 U12159 ( .A1(n13021), .A2(n13235), .ZN(n20161) );
  NAND2_X1 U12160 ( .A1(n20161), .A2(n9821), .ZN(n16076) );
  AND2_X1 U12161 ( .A1(n12033), .A2(n20242), .ZN(n14378) );
  INV_X1 U12162 ( .A(n14304), .ZN(n14377) );
  OR2_X1 U12163 ( .A1(n13156), .A2(n13155), .ZN(n14394) );
  AND2_X1 U12164 ( .A1(n12899), .A2(n12898), .ZN(n20167) );
  XNOR2_X1 U12165 ( .A(n13338), .B(n13337), .ZN(n14459) );
  OR2_X1 U12166 ( .A1(n13336), .A2(n14466), .ZN(n13338) );
  OAI21_X1 U12167 ( .B1(n9775), .B2(n9696), .A(n9672), .ZN(n14579) );
  AOI21_X1 U12168 ( .B1(n14293), .B2(n14292), .A(n14291), .ZN(n16108) );
  AND2_X1 U12169 ( .A1(n13028), .A2(n20797), .ZN(n16140) );
  INV_X1 U12170 ( .A(n20063), .ZN(n16141) );
  INV_X1 U12171 ( .A(n16140), .ZN(n20243) );
  OR2_X2 U12172 ( .A1(n13036), .A2(n15947), .ZN(n20063) );
  INV_X1 U12173 ( .A(n16144), .ZN(n16128) );
  MUX2_X1 U12174 ( .A(n14074), .B(n14073), .S(n14085), .Z(n14057) );
  NAND2_X1 U12175 ( .A1(n9832), .A2(n9831), .ZN(n14457) );
  XNOR2_X1 U12176 ( .A(n14076), .B(n14075), .ZN(n14663) );
  AOI22_X1 U12177 ( .A1(n14085), .A2(n14073), .B1(n14101), .B2(n14072), .ZN(
        n14076) );
  NAND2_X1 U12178 ( .A1(n14455), .A2(n14670), .ZN(n14470) );
  INV_X1 U12179 ( .A(n14455), .ZN(n14495) );
  XNOR2_X1 U12180 ( .A(n10031), .B(n14452), .ZN(n14711) );
  AOI21_X1 U12181 ( .B1(n16112), .B2(n14717), .A(n9746), .ZN(n10034) );
  NAND2_X1 U12182 ( .A1(n14518), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10032) );
  AND2_X1 U12183 ( .A1(n13256), .A2(n13241), .ZN(n16249) );
  NAND2_X1 U12184 ( .A1(n11946), .A2(n11041), .ZN(n13240) );
  AND2_X1 U12185 ( .A1(n16197), .A2(n20229), .ZN(n14798) );
  INV_X1 U12186 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20696) );
  CLKBUF_X1 U12187 ( .A(n12948), .Z(n20541) );
  OR2_X1 U12188 ( .A1(n13371), .A2(n13372), .ZN(n20637) );
  INV_X1 U12189 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20240) );
  OAI21_X1 U12190 ( .B1(n13185), .B2(n16270), .A(n20413), .ZN(n20239) );
  NOR2_X1 U12191 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16255) );
  OR2_X1 U12192 ( .A1(n20371), .A2(n20365), .ZN(n20409) );
  INV_X1 U12193 ( .A(n20409), .ZN(n20432) );
  INV_X1 U12194 ( .A(n20501), .ZN(n20462) );
  OAI211_X1 U12195 ( .C1(n20562), .C2(n20669), .A(n20598), .B(n20546), .ZN(
        n20564) );
  INV_X1 U12196 ( .A(n20629), .ZN(n20587) );
  NAND2_X1 U12197 ( .A1(n20631), .A2(n20694), .ZN(n20629) );
  OAI22_X1 U12198 ( .A1(n20602), .A2(n20601), .B1(n20600), .B2(n20730), .ZN(
        n20625) );
  INV_X1 U12199 ( .A(n20640), .ZN(n20657) );
  OAI211_X1 U12200 ( .C1(n20688), .C2(n20669), .A(n20742), .B(n20668), .ZN(
        n20690) );
  AND2_X1 U12201 ( .A1(n20735), .A2(n20661), .ZN(n20724) );
  INV_X1 U12202 ( .A(n20802), .ZN(n20733) );
  INV_X1 U12203 ( .A(n20814), .ZN(n20749) );
  INV_X1 U12204 ( .A(n20821), .ZN(n20755) );
  INV_X1 U12205 ( .A(n20828), .ZN(n20761) );
  INV_X1 U12206 ( .A(n20835), .ZN(n20767) );
  INV_X1 U12207 ( .A(n20842), .ZN(n20773) );
  INV_X1 U12208 ( .A(n20849), .ZN(n20779) );
  OAI211_X1 U12209 ( .C1(n20786), .C2(n20743), .A(n20742), .B(n20741), .ZN(
        n20789) );
  INV_X1 U12210 ( .A(n20858), .ZN(n20787) );
  OR2_X1 U12211 ( .A1(n15953), .A2(n20868), .ZN(n20057) );
  AND2_X1 U12212 ( .A1(n12597), .A2(n19145), .ZN(n14861) );
  INV_X1 U12213 ( .A(n10013), .ZN(n14860) );
  NOR2_X1 U12214 ( .A1(n16286), .A2(n16288), .ZN(n16287) );
  OAI21_X1 U12215 ( .B1(n16303), .B2(n10007), .A(n10006), .ZN(n14874) );
  NAND2_X1 U12216 ( .A1(n10008), .A2(n15136), .ZN(n10007) );
  NAND2_X1 U12217 ( .A1(n19162), .A2(n10008), .ZN(n10006) );
  INV_X1 U12218 ( .A(n15128), .ZN(n10008) );
  NOR2_X1 U12219 ( .A1(n16303), .A2(n16305), .ZN(n16304) );
  NAND2_X1 U12220 ( .A1(n19162), .A2(n15156), .ZN(n10020) );
  NAND2_X1 U12221 ( .A1(n19000), .A2(n10023), .ZN(n10022) );
  NOR2_X1 U12222 ( .A1(n19000), .A2(n19162), .ZN(n18982) );
  NOR2_X1 U12223 ( .A1(n18982), .A2(n18983), .ZN(n18981) );
  OR2_X1 U12224 ( .A1(n18952), .A2(n10887), .ZN(n19188) );
  AND2_X1 U12225 ( .A1(n10882), .A2(n10881), .ZN(n19153) );
  INV_X1 U12226 ( .A(n19174), .ZN(n19190) );
  INV_X1 U12227 ( .A(n19153), .ZN(n19194) );
  INV_X1 U12228 ( .A(n19097), .ZN(n19198) );
  OR2_X1 U12229 ( .A1(n10811), .A2(n10810), .ZN(n13477) );
  OR2_X1 U12230 ( .A1(n10732), .A2(n10731), .ZN(n13201) );
  AND2_X1 U12231 ( .A1(n13982), .A2(n19375), .ZN(n19209) );
  OR2_X1 U12232 ( .A1(n19207), .A2(n13982), .ZN(n19241) );
  INV_X1 U12233 ( .A(n19215), .ZN(n19265) );
  INV_X1 U12234 ( .A(n19280), .ZN(n19345) );
  NAND2_X1 U12236 ( .A1(n9789), .A2(n10210), .ZN(n9788) );
  NAND2_X1 U12237 ( .A1(n15297), .A2(n9722), .ZN(n9787) );
  NAND2_X1 U12238 ( .A1(n18958), .A2(n12513), .ZN(n16359) );
  AND2_X1 U12239 ( .A1(n10084), .A2(n10480), .ZN(n13004) );
  INV_X1 U12240 ( .A(n16351), .ZN(n19359) );
  INV_X1 U12241 ( .A(n16325), .ZN(n19352) );
  AND2_X1 U12242 ( .A1(n16359), .A2(n12927), .ZN(n16351) );
  INV_X1 U12243 ( .A(n16359), .ZN(n19349) );
  NAND2_X1 U12244 ( .A1(n15148), .A2(n12394), .ZN(n15135) );
  NOR2_X1 U12245 ( .A1(n15438), .A2(n12503), .ZN(n15394) );
  INV_X1 U12246 ( .A(n9946), .ZN(n9945) );
  OR2_X1 U12247 ( .A1(n15213), .A2(n9951), .ZN(n9944) );
  OR2_X1 U12248 ( .A1(n15497), .A2(n12501), .ZN(n15438) );
  OAI21_X1 U12249 ( .B1(n15256), .B2(n9930), .A(n9927), .ZN(n15224) );
  NAND2_X1 U12250 ( .A1(n9933), .A2(n9931), .ZN(n15236) );
  INV_X1 U12251 ( .A(n9934), .ZN(n9931) );
  OAI21_X1 U12252 ( .B1(n15256), .B2(n15162), .A(n15254), .ZN(n15244) );
  NAND2_X1 U12253 ( .A1(n12329), .A2(n12328), .ZN(n9923) );
  CLKBUF_X1 U12254 ( .A(n15600), .Z(n15601) );
  OR2_X1 U12255 ( .A1(n12477), .A2(n12459), .ZN(n16371) );
  NAND2_X1 U12256 ( .A1(n9989), .A2(n9990), .ZN(n13610) );
  NAND2_X1 U12257 ( .A1(n13454), .A2(n9993), .ZN(n9989) );
  NAND2_X1 U12258 ( .A1(n12127), .A2(n9942), .ZN(n9792) );
  INV_X1 U12259 ( .A(n9915), .ZN(n12045) );
  NAND2_X1 U12260 ( .A1(n15458), .A2(n12478), .ZN(n19370) );
  OR2_X1 U12261 ( .A1(n12726), .A2(n12689), .ZN(n20037) );
  INV_X1 U12262 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20033) );
  INV_X1 U12263 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20023) );
  XNOR2_X1 U12264 ( .A(n12932), .B(n12894), .ZN(n20019) );
  XNOR2_X1 U12265 ( .A(n12930), .B(n12931), .ZN(n12894) );
  INV_X1 U12266 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15978) );
  INV_X1 U12267 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16424) );
  NAND2_X1 U12268 ( .A1(n12888), .A2(n12733), .ZN(n20028) );
  INV_X1 U12269 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16397) );
  OAI21_X1 U12270 ( .B1(n19389), .B2(n19384), .A(n19383), .ZN(n19426) );
  OAI211_X1 U12271 ( .C1(n19475), .C2(n19460), .A(n19459), .B(n19868), .ZN(
        n19478) );
  OAI21_X1 U12272 ( .B1(n19523), .B2(n19522), .A(n19521), .ZN(n19541) );
  NOR2_X1 U12273 ( .A1(n19572), .A2(n19788), .ZN(n19558) );
  NOR2_X1 U12274 ( .A1(n19608), .A2(n19788), .ZN(n19590) );
  OAI21_X1 U12275 ( .B1(n19655), .B2(n19635), .A(n19868), .ZN(n19657) );
  OAI21_X1 U12276 ( .B1(n19701), .B2(n19716), .A(n19868), .ZN(n19719) );
  INV_X1 U12277 ( .A(n19696), .ZN(n19718) );
  OAI21_X1 U12278 ( .B1(n19774), .B2(n19632), .A(n19757), .ZN(n19777) );
  NOR2_X1 U12279 ( .A1(n19753), .A2(n19752), .ZN(n19775) );
  OAI22_X1 U12280 ( .A1(n19406), .A2(n19419), .B1(n19405), .B2(n19417), .ZN(
        n19800) );
  INV_X1 U12281 ( .A(n19879), .ZN(n19829) );
  INV_X1 U12282 ( .A(n19897), .ZN(n19841) );
  OAI21_X1 U12283 ( .B1(n19826), .B2(n19825), .A(n19824), .ZN(n19853) );
  OAI22_X1 U12284 ( .A1(n19420), .A2(n19419), .B1(n19418), .B2(n19417), .ZN(
        n19852) );
  AND2_X1 U12285 ( .A1(n10583), .A2(n19421), .ZN(n19874) );
  INV_X1 U12286 ( .A(n19803), .ZN(n19900) );
  AND2_X1 U12287 ( .A1(n10869), .A2(n19421), .ZN(n19898) );
  NOR2_X1 U12288 ( .A1(n19815), .A2(n19814), .ZN(n19901) );
  NOR2_X2 U12289 ( .A1(n19789), .A2(n19814), .ZN(n19917) );
  INV_X1 U12290 ( .A(n19852), .ZN(n19922) );
  INV_X1 U12291 ( .A(n19901), .ZN(n19921) );
  OR2_X1 U12292 ( .A1(n19932), .A2(n20035), .ZN(n18956) );
  AND2_X1 U12293 ( .A1(n16394), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16421) );
  XNOR2_X1 U12294 ( .A(n18929), .B(n18277), .ZN(n18943) );
  OAI21_X1 U12295 ( .B1(n18710), .B2(n10213), .A(n17511), .ZN(n18944) );
  INV_X1 U12296 ( .A(n18771), .ZN(n18925) );
  INV_X1 U12297 ( .A(n17018), .ZN(n16983) );
  NOR2_X1 U12298 ( .A1(n16754), .A2(n17665), .ZN(n16753) );
  AND2_X1 U12299 ( .A1(n16763), .A2(n16641), .ZN(n16754) );
  AND2_X1 U12300 ( .A1(n9971), .A2(n9970), .ZN(n16804) );
  INV_X1 U12301 ( .A(n17730), .ZN(n9970) );
  INV_X1 U12302 ( .A(n9971), .ZN(n16805) );
  NOR2_X1 U12303 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16960), .ZN(n16942) );
  NAND2_X1 U12304 ( .A1(n17278), .A2(n17149), .ZN(n17174) );
  AND2_X1 U12305 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17282), .ZN(n17278) );
  INV_X1 U12306 ( .A(n17148), .ZN(n17282) );
  INV_X1 U12307 ( .A(n17326), .ZN(n17321) );
  NOR2_X1 U12308 ( .A1(n17335), .A2(n17537), .ZN(n17329) );
  NAND2_X1 U12309 ( .A1(n17339), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n17335) );
  NOR2_X1 U12310 ( .A1(n17345), .A2(n17533), .ZN(n17339) );
  INV_X1 U12311 ( .A(n17349), .ZN(n17346) );
  NAND2_X1 U12312 ( .A1(n17346), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17345) );
  NOR2_X1 U12313 ( .A1(n17404), .A2(n17355), .ZN(n17350) );
  NOR2_X1 U12314 ( .A1(n17395), .A2(n9881), .ZN(n17356) );
  NAND2_X1 U12315 ( .A1(n9781), .A2(n9882), .ZN(n9881) );
  INV_X1 U12316 ( .A(n17360), .ZN(n9882) );
  NOR2_X1 U12317 ( .A1(n17518), .A2(n17388), .ZN(n17382) );
  NOR3_X1 U12318 ( .A1(n17404), .A2(n17395), .A3(n17516), .ZN(n17384) );
  NAND2_X1 U12319 ( .A1(n17399), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17395) );
  INV_X1 U12320 ( .A(n17367), .ZN(n17393) );
  INV_X1 U12321 ( .A(n17387), .ZN(n17394) );
  NAND4_X1 U12322 ( .A1(n17434), .A2(P3_EAX_REG_13__SCAN_IN), .A3(
        P3_EAX_REG_12__SCAN_IN), .A4(n17315), .ZN(n17403) );
  INV_X1 U12323 ( .A(n17458), .ZN(n17435) );
  OR2_X1 U12324 ( .A1(n17468), .A2(n9894), .ZN(n17439) );
  INV_X1 U12325 ( .A(n17440), .ZN(n9895) );
  NOR2_X1 U12326 ( .A1(n15770), .A2(n15769), .ZN(n17450) );
  INV_X1 U12327 ( .A(n15869), .ZN(n17454) );
  NOR2_X1 U12328 ( .A1(n15780), .A2(n15779), .ZN(n17459) );
  NAND2_X1 U12329 ( .A1(n15984), .A2(n17316), .ZN(n17460) );
  INV_X1 U12330 ( .A(n15870), .ZN(n17464) );
  NAND2_X1 U12331 ( .A1(n17316), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n17468) );
  INV_X1 U12332 ( .A(n17460), .ZN(n17465) );
  NOR2_X1 U12333 ( .A1(n15983), .A2(n15982), .ZN(n17466) );
  NOR2_X1 U12334 ( .A1(n18281), .A2(n17564), .ZN(n17565) );
  INV_X1 U12335 ( .A(n17510), .ZN(n17512) );
  NAND2_X1 U12337 ( .A1(n16451), .A2(n9859), .ZN(n9858) );
  NAND2_X1 U12338 ( .A1(n16487), .A2(n17774), .ZN(n9859) );
  NOR2_X1 U12339 ( .A1(n17589), .A2(n17590), .ZN(n16469) );
  NAND2_X1 U12340 ( .A1(n17986), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17629) );
  NOR3_X1 U12341 ( .A1(n9808), .A2(n17948), .A3(n9844), .ZN(n17628) );
  INV_X1 U12342 ( .A(n17986), .ZN(n9808) );
  INV_X1 U12343 ( .A(n17743), .ZN(n9961) );
  INV_X1 U12344 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17727) );
  NAND4_X1 U12345 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17828) );
  NAND2_X1 U12346 ( .A1(n16966), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17888) );
  INV_X1 U12347 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17927) );
  OAI21_X1 U12348 ( .B1(n16447), .B2(n16446), .A(n10120), .ZN(n10119) );
  NAND2_X1 U12349 ( .A1(n10125), .A2(n10124), .ZN(n9862) );
  AND2_X1 U12350 ( .A1(n16491), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10118) );
  NAND2_X1 U12351 ( .A1(n17595), .A2(n21110), .ZN(n15964) );
  NOR2_X1 U12352 ( .A1(n15886), .A2(n17444), .ZN(n16495) );
  NOR2_X1 U12353 ( .A1(n17966), .A2(n18172), .ZN(n9802) );
  OR2_X1 U12354 ( .A1(n17952), .A2(n9806), .ZN(n9805) );
  INV_X1 U12355 ( .A(n9807), .ZN(n9806) );
  AOI21_X1 U12356 ( .B1(n17953), .B2(n17954), .A(n17971), .ZN(n9807) );
  INV_X1 U12357 ( .A(n18166), .ZN(n18126) );
  NAND2_X1 U12358 ( .A1(n17684), .A2(n15915), .ZN(n17635) );
  INV_X1 U12359 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18930) );
  NAND2_X1 U12360 ( .A1(n17771), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18075) );
  INV_X1 U12361 ( .A(n18236), .ZN(n18151) );
  NAND2_X1 U12362 ( .A1(n15905), .A2(n18125), .ZN(n18167) );
  NOR2_X1 U12363 ( .A1(n18713), .A2(n18242), .ZN(n18196) );
  NOR2_X1 U12364 ( .A1(n18943), .A2(n15741), .ZN(n18718) );
  INV_X1 U12365 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18755) );
  INV_X1 U12366 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18905) );
  AND2_X1 U12367 ( .A1(n12031), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20241)
         );
  CLKBUF_X1 U12368 ( .A(n16597), .Z(n16603) );
  NAND2_X1 U12369 ( .A1(n10287), .A2(n10286), .ZN(n10893) );
  CLKBUF_X1 U12370 ( .A(n13208), .Z(n13129) );
  AND2_X1 U12371 ( .A1(n10110), .A2(n15045), .ZN(n10109) );
  INV_X1 U12372 ( .A(n12533), .ZN(n12534) );
  OAI21_X1 U12373 ( .B1(n12532), .B2(n19376), .A(n12531), .ZN(n12533) );
  OAI21_X1 U12374 ( .B1(n15334), .B2(n16324), .A(n9985), .ZN(P2_U2986) );
  NOR2_X1 U12375 ( .A1(n9715), .A2(n9986), .ZN(n9985) );
  INV_X1 U12376 ( .A(n12581), .ZN(n9986) );
  INV_X1 U12377 ( .A(n10114), .ZN(n10117) );
  INV_X1 U12378 ( .A(n10116), .ZN(n10115) );
  AOI21_X1 U12379 ( .B1(n15317), .B2(n19361), .A(n15316), .ZN(n15318) );
  NAND2_X1 U12380 ( .A1(n9723), .A2(n9681), .ZN(P2_U3017) );
  NOR2_X1 U12381 ( .A1(n9725), .A2(n9958), .ZN(n9957) );
  AOI21_X1 U12382 ( .B1(n15332), .B2(n16361), .A(n15331), .ZN(n15333) );
  AOI21_X1 U12383 ( .B1(n9968), .B2(n17006), .A(n9964), .ZN(n16669) );
  NAND2_X1 U12384 ( .A1(n9966), .A2(n9965), .ZN(n9964) );
  INV_X1 U12385 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16994) );
  NAND2_X1 U12386 ( .A1(n9861), .A2(n9857), .ZN(P3_U2799) );
  AOI21_X1 U12387 ( .B1(n9860), .B2(n9653), .A(n9858), .ZN(n9857) );
  NAND2_X1 U12388 ( .A1(n16490), .A2(n17748), .ZN(n9861) );
  INV_X1 U12389 ( .A(n16485), .ZN(n9860) );
  NAND2_X1 U12390 ( .A1(n17686), .A2(n9675), .ZN(n17652) );
  NAND2_X1 U12391 ( .A1(n9803), .A2(n9801), .ZN(P3_U2836) );
  OAI21_X1 U12392 ( .B1(n9805), .B2(n18242), .A(n9804), .ZN(n9803) );
  AOI211_X1 U12393 ( .C1(n17964), .C2(n17965), .A(n9802), .B(n17963), .ZN(
        n9801) );
  NOR2_X1 U12394 ( .A1(n18252), .A2(n17961), .ZN(n9804) );
  AND2_X1 U12395 ( .A1(n9990), .A2(n9988), .ZN(n9669) );
  NOR2_X1 U12396 ( .A1(n15179), .A2(n15409), .ZN(n9670) );
  NAND2_X1 U12397 ( .A1(n9670), .A2(n9780), .ZN(n15131) );
  AND2_X1 U12398 ( .A1(n12711), .A2(n12237), .ZN(n9671) );
  INV_X4 U12399 ( .A(n12841), .ZN(n17263) );
  INV_X1 U12400 ( .A(n10201), .ZN(n10200) );
  NAND2_X1 U12401 ( .A1(n10202), .A2(n10205), .ZN(n10201) );
  NAND2_X1 U12402 ( .A1(n10264), .A2(n9686), .ZN(n10244) );
  NAND2_X1 U12403 ( .A1(n10242), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10243) );
  OR2_X1 U12404 ( .A1(n19422), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10235) );
  OR2_X1 U12405 ( .A1(n17012), .A2(n12741), .ZN(n15648) );
  INV_X2 U12406 ( .A(n14449), .ZN(n14601) );
  INV_X1 U12407 ( .A(n10059), .ZN(n10070) );
  OR2_X1 U12408 ( .A1(n14194), .A2(n10193), .ZN(n9672) );
  INV_X4 U12409 ( .A(n14601), .ZN(n16112) );
  AND2_X1 U12410 ( .A1(n15173), .A2(n15172), .ZN(n9673) );
  AND2_X1 U12411 ( .A1(n9666), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10675) );
  OR2_X1 U12412 ( .A1(n15179), .A2(n9954), .ZN(n12537) );
  NAND2_X1 U12413 ( .A1(n10180), .A2(n10183), .ZN(n14165) );
  NAND2_X1 U12414 ( .A1(n14904), .A2(n9756), .ZN(n14879) );
  AND2_X1 U12415 ( .A1(n15985), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n9674) );
  NAND2_X1 U12416 ( .A1(n10059), .A2(n14696), .ZN(n10058) );
  AND2_X2 U12417 ( .A1(n10288), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10351) );
  AND2_X1 U12418 ( .A1(n12941), .A2(n12061), .ZN(n12152) );
  AND2_X1 U12419 ( .A1(n17658), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9675) );
  AND2_X1 U12420 ( .A1(n10028), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9676) );
  INV_X1 U12421 ( .A(n17317), .ZN(n18301) );
  AND2_X1 U12422 ( .A1(n10085), .A2(n13377), .ZN(n9677) );
  AND2_X1 U12423 ( .A1(n10013), .A2(n19145), .ZN(n14851) );
  AND2_X1 U12424 ( .A1(n10201), .A2(n9785), .ZN(n16340) );
  INV_X1 U12425 ( .A(n10199), .ZN(n15141) );
  NAND2_X1 U12426 ( .A1(n12129), .A2(n12128), .ZN(n13608) );
  AND2_X1 U12427 ( .A1(n9927), .A2(n15165), .ZN(n9678) );
  NOR2_X1 U12428 ( .A1(n14964), .A2(n14965), .ZN(n9679) );
  AND2_X1 U12429 ( .A1(n9661), .A2(n10394), .ZN(n9680) );
  AND2_X1 U12430 ( .A1(n9667), .A2(n10383), .ZN(n10694) );
  NAND2_X1 U12431 ( .A1(n10170), .A2(n9758), .ZN(n10174) );
  AND2_X1 U12432 ( .A1(n12565), .A2(n9957), .ZN(n9681) );
  AND2_X1 U12433 ( .A1(n10135), .A2(n10871), .ZN(n9682) );
  AND2_X1 U12434 ( .A1(n13009), .A2(n13011), .ZN(n9683) );
  OAI21_X1 U12435 ( .B1(n10431), .B2(n12277), .A(n10430), .ZN(n10452) );
  AND2_X1 U12436 ( .A1(n13765), .A2(n9743), .ZN(n14983) );
  NOR2_X1 U12437 ( .A1(n10243), .A2(n10240), .ZN(n10268) );
  NOR2_X1 U12438 ( .A1(n13379), .A2(n10105), .ZN(n13476) );
  NAND2_X1 U12439 ( .A1(n15509), .A2(n9741), .ZN(n14920) );
  INV_X1 U12440 ( .A(n10253), .ZN(n10019) );
  AND4_X1 U12441 ( .A1(n10019), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n9684) );
  AND2_X1 U12442 ( .A1(n10838), .A2(n15085), .ZN(n9685) );
  AND2_X1 U12443 ( .A1(n10015), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9686) );
  OR2_X1 U12444 ( .A1(n10184), .A2(n14262), .ZN(n9687) );
  AOI21_X1 U12445 ( .B1(n13693), .B2(n15894), .A(n13692), .ZN(n18712) );
  INV_X1 U12446 ( .A(n18712), .ZN(n9891) );
  NOR2_X1 U12447 ( .A1(n16304), .A2(n19162), .ZN(n9688) );
  AND2_X1 U12448 ( .A1(n10025), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9689) );
  AND2_X1 U12449 ( .A1(n12342), .A2(n9764), .ZN(n9690) );
  AND2_X1 U12450 ( .A1(n19152), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9691) );
  NAND2_X1 U12451 ( .A1(n10483), .A2(n10482), .ZN(n10084) );
  AND2_X1 U12452 ( .A1(n14962), .A2(n10144), .ZN(n9692) );
  AND2_X1 U12453 ( .A1(n9780), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9693) );
  INV_X2 U12454 ( .A(n11027), .ZN(n11869) );
  AND2_X2 U12455 ( .A1(n13875), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10602) );
  OR3_X1 U12456 ( .A1(n15022), .A2(n10074), .A3(n10073), .ZN(n9694) );
  INV_X1 U12457 ( .A(n10619), .ZN(n10722) );
  NAND2_X1 U12459 ( .A1(n10146), .A2(n10145), .ZN(n10461) );
  NAND2_X1 U12460 ( .A1(n12330), .A2(n12435), .ZN(n12324) );
  OR4_X1 U12461 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9695) );
  AND2_X1 U12462 ( .A1(n10192), .A2(n11516), .ZN(n9696) );
  INV_X2 U12463 ( .A(n13435), .ZN(n14008) );
  AND2_X1 U12464 ( .A1(n9980), .A2(n9979), .ZN(n15300) );
  OR2_X1 U12465 ( .A1(n10637), .A2(n10636), .ZN(n9697) );
  OR4_X1 U12466 ( .A1(n15324), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15310), .A4(n12506), .ZN(n9698) );
  INV_X1 U12467 ( .A(n14565), .ZN(n9913) );
  AND2_X1 U12468 ( .A1(n11066), .A2(n11965), .ZN(n11046) );
  NOR2_X1 U12469 ( .A1(n14271), .A2(n9687), .ZN(n14256) );
  NAND2_X1 U12470 ( .A1(n9670), .A2(n9693), .ZN(n15124) );
  INV_X1 U12471 ( .A(n12827), .ZN(n17190) );
  AND4_X1 U12472 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(
        n9699) );
  AND2_X1 U12473 ( .A1(n12941), .A2(n15624), .ZN(n9700) );
  INV_X1 U12474 ( .A(n12728), .ZN(n19175) );
  AND2_X1 U12475 ( .A1(n10206), .A2(n16341), .ZN(n9701) );
  NOR2_X1 U12476 ( .A1(n14271), .A2(n14272), .ZN(n14164) );
  AND2_X1 U12477 ( .A1(n14224), .A2(n14223), .ZN(n9702) );
  NAND2_X1 U12478 ( .A1(n14623), .A2(n14438), .ZN(n14612) );
  AND3_X1 U12479 ( .A1(n10307), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10306), .ZN(n9703) );
  NAND2_X1 U12480 ( .A1(n11047), .A2(n11040), .ZN(n9704) );
  AND3_X1 U12481 ( .A1(n10984), .A2(n10178), .A3(n10177), .ZN(n9705) );
  AND2_X1 U12482 ( .A1(n12941), .A2(n12052), .ZN(n12154) );
  NAND2_X1 U12483 ( .A1(n9827), .A2(n14428), .ZN(n14627) );
  XNOR2_X1 U12484 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12437), .ZN(
        n9707) );
  INV_X1 U12485 ( .A(n15624), .ZN(n19191) );
  NAND2_X1 U12486 ( .A1(n14532), .A2(n14493), .ZN(n14479) );
  AND4_X1 U12487 ( .A1(n10931), .A2(n10933), .A3(n10930), .A4(n10932), .ZN(
        n9708) );
  AND2_X1 U12488 ( .A1(n10946), .A2(n11965), .ZN(n11969) );
  NAND2_X1 U12489 ( .A1(n12186), .A2(n12185), .ZN(n12199) );
  AND3_X1 U12490 ( .A1(n10997), .A2(n10994), .A3(n10996), .ZN(n9709) );
  AND3_X1 U12491 ( .A1(n10945), .A2(n10939), .A3(n10944), .ZN(n9710) );
  AND2_X1 U12492 ( .A1(n15133), .A2(n10004), .ZN(n9711) );
  OR3_X1 U12493 ( .A1(n15324), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15310), .ZN(n9712) );
  NAND2_X1 U12494 ( .A1(n10584), .A2(n10412), .ZN(n10417) );
  INV_X1 U12495 ( .A(n20272), .ZN(n9902) );
  AND4_X1 U12496 ( .A1(n12082), .A2(n12081), .A3(n12080), .A4(n12079), .ZN(
        n9713) );
  NAND2_X1 U12497 ( .A1(n10203), .A2(n10204), .ZN(n16339) );
  AND2_X1 U12498 ( .A1(n14455), .A2(n9830), .ZN(n9714) );
  NAND2_X1 U12499 ( .A1(n10128), .A2(n18162), .ZN(n15905) );
  INV_X1 U12500 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13713) );
  NOR2_X1 U12501 ( .A1(n15320), .A2(n16325), .ZN(n9715) );
  AND2_X1 U12502 ( .A1(n10351), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10680) );
  XNOR2_X1 U12503 ( .A(n12455), .B(n12454), .ZN(n16277) );
  NAND2_X1 U12504 ( .A1(n9670), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10199) );
  AND2_X1 U12505 ( .A1(n12098), .A2(n12097), .ZN(n9716) );
  AND2_X1 U12506 ( .A1(n10059), .A2(n14446), .ZN(n9717) );
  OR2_X1 U12507 ( .A1(n14889), .A2(n14890), .ZN(n9718) );
  AND2_X1 U12508 ( .A1(n10421), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9719) );
  AND2_X1 U12509 ( .A1(n13461), .A2(n10165), .ZN(n9720) );
  INV_X1 U12510 ( .A(n9994), .ZN(n9993) );
  OR2_X1 U12511 ( .A1(n12286), .A2(n9995), .ZN(n9994) );
  AND2_X1 U12512 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9721) );
  AND2_X1 U12513 ( .A1(n9701), .A2(n10210), .ZN(n9722) );
  OR2_X1 U12514 ( .A1(n12564), .A2(n15597), .ZN(n9723) );
  NAND2_X1 U12515 ( .A1(n9912), .A2(n9911), .ZN(n14537) );
  AND3_X1 U12516 ( .A1(n11073), .A2(n12954), .A3(n11053), .ZN(n9724) );
  AND2_X1 U12517 ( .A1(n14137), .A2(n10195), .ZN(n14087) );
  INV_X1 U12518 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11523) );
  INV_X1 U12519 ( .A(n12075), .ZN(n10149) );
  INV_X1 U12520 ( .A(n9851), .ZN(n16500) );
  NAND2_X1 U12521 ( .A1(n15920), .A2(n9852), .ZN(n9851) );
  OR2_X1 U12522 ( .A1(n12562), .A2(n10072), .ZN(n9725) );
  INV_X1 U12523 ( .A(n10050), .ZN(n14119) );
  NAND3_X1 U12524 ( .A1(n14493), .A2(n14532), .A3(n10056), .ZN(n9726) );
  INV_X1 U12525 ( .A(n10058), .ZN(n10057) );
  OR2_X1 U12526 ( .A1(n12094), .A2(n12093), .ZN(n9727) );
  INV_X1 U12527 ( .A(n10134), .ZN(n12353) );
  NAND2_X1 U12528 ( .A1(n12324), .A2(n10872), .ZN(n10134) );
  INV_X1 U12529 ( .A(n13439), .ZN(n10042) );
  INV_X1 U12530 ( .A(n10068), .ZN(n10067) );
  NAND2_X1 U12531 ( .A1(n16086), .A2(n10069), .ZN(n10068) );
  NOR2_X1 U12532 ( .A1(n14889), .A2(n10168), .ZN(n12606) );
  AND3_X1 U12533 ( .A1(n15794), .A2(n15793), .A3(n15792), .ZN(n9728) );
  AND2_X1 U12534 ( .A1(n17595), .A2(n9854), .ZN(n9729) );
  AND3_X1 U12535 ( .A1(n12096), .A2(n9727), .A3(n12095), .ZN(n9730) );
  AND3_X1 U12536 ( .A1(n13029), .A2(n12869), .A3(n9818), .ZN(n9731) );
  AND2_X1 U12537 ( .A1(n15799), .A2(n10127), .ZN(n9732) );
  AND3_X1 U12538 ( .A1(n9661), .A2(n10394), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n9733) );
  AND2_X1 U12539 ( .A1(n10891), .A2(n10890), .ZN(n9734) );
  NOR2_X1 U12540 ( .A1(n12202), .A2(n12481), .ZN(n9735) );
  AND2_X1 U12541 ( .A1(n9960), .A2(n9959), .ZN(n9736) );
  AND2_X1 U12542 ( .A1(n10425), .A2(n10424), .ZN(n10453) );
  AND2_X1 U12543 ( .A1(n10407), .A2(n12215), .ZN(n9737) );
  AND2_X1 U12544 ( .A1(n9677), .A2(n10087), .ZN(n9738) );
  AND2_X1 U12545 ( .A1(n16819), .A2(n9961), .ZN(n9739) );
  INV_X1 U12546 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10910) );
  INV_X1 U12547 ( .A(n12302), .ZN(n12196) );
  NAND2_X1 U12548 ( .A1(n12199), .A2(n12188), .ZN(n12302) );
  NAND2_X1 U12549 ( .A1(n17684), .A2(n17671), .ZN(n17672) );
  INV_X1 U12550 ( .A(n17672), .ZN(n9840) );
  AND3_X1 U12551 ( .A1(n13029), .A2(n12869), .A3(n20292), .ZN(n12014) );
  NOR2_X1 U12552 ( .A1(n12762), .A2(n12761), .ZN(n18277) );
  INV_X1 U12553 ( .A(n18277), .ZN(n9888) );
  NOR2_X1 U12554 ( .A1(n10262), .A2(n15257), .ZN(n10247) );
  NAND2_X1 U12555 ( .A1(n13578), .A2(n13600), .ZN(n13599) );
  NAND2_X1 U12556 ( .A1(n13421), .A2(n13432), .ZN(n13431) );
  NOR2_X1 U12557 ( .A1(n10255), .A2(n15302), .ZN(n10250) );
  NAND2_X1 U12558 ( .A1(n12291), .A2(n10135), .ZN(n9740) );
  AND2_X1 U12559 ( .A1(n12293), .A2(n12292), .ZN(n12291) );
  AND2_X1 U12560 ( .A1(n15489), .A2(n15510), .ZN(n9741) );
  NOR2_X1 U12561 ( .A1(n15094), .A2(n15093), .ZN(n15095) );
  AND2_X1 U12562 ( .A1(n10247), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10245) );
  AND2_X1 U12563 ( .A1(n13765), .A2(n15018), .ZN(n14999) );
  NAND2_X1 U12564 ( .A1(n13765), .A2(n10108), .ZN(n14989) );
  AND2_X1 U12565 ( .A1(n10250), .A2(n10028), .ZN(n10249) );
  NAND2_X1 U12566 ( .A1(n9792), .A2(n13529), .ZN(n13451) );
  INV_X1 U12567 ( .A(n14601), .ZN(n10059) );
  NOR3_X1 U12568 ( .A1(n15022), .A2(n15006), .A3(n10076), .ZN(n14992) );
  OR3_X1 U12569 ( .A1(n15022), .A2(n10074), .A3(n15006), .ZN(n9742) );
  OAI22_X1 U12570 ( .A1(n12529), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19926), 
        .B2(n12444), .ZN(n10267) );
  INV_X1 U12571 ( .A(n17932), .ZN(n17943) );
  NOR2_X2 U12572 ( .A1(n18929), .A2(n16618), .ZN(n17932) );
  NOR2_X1 U12573 ( .A1(n14897), .A2(n19162), .ZN(n16303) );
  AND2_X1 U12574 ( .A1(n17686), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10229) );
  XNOR2_X1 U12575 ( .A(n13889), .B(n13891), .ZN(n14959) );
  NOR2_X1 U12576 ( .A1(n10253), .A2(n13525), .ZN(n10251) );
  NOR2_X1 U12577 ( .A1(n13848), .A2(n14973), .ZN(n14964) );
  NAND2_X1 U12578 ( .A1(n15445), .A2(n15085), .ZN(n15084) );
  OR2_X1 U12579 ( .A1(n17846), .A2(n15863), .ZN(n9813) );
  AND2_X1 U12580 ( .A1(n10108), .A2(n10107), .ZN(n9743) );
  NOR2_X1 U12581 ( .A1(n14294), .A2(n14212), .ZN(n9744) );
  AND2_X1 U12582 ( .A1(n14125), .A2(n14136), .ZN(n9745) );
  AND2_X1 U12583 ( .A1(n12893), .A2(n12892), .ZN(n12930) );
  AND2_X1 U12584 ( .A1(n14601), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9746) );
  NAND2_X1 U12585 ( .A1(n16643), .A2(n16980), .ZN(n9747) );
  INV_X1 U12586 ( .A(n13011), .ZN(n13126) );
  NAND2_X1 U12587 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9748) );
  INV_X1 U12588 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10901) );
  INV_X1 U12589 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10051) );
  INV_X1 U12590 ( .A(n13484), .ZN(n13626) );
  OR2_X1 U12591 ( .A1(n10824), .A2(n10823), .ZN(n13484) );
  INV_X1 U12592 ( .A(n10184), .ZN(n10183) );
  NAND2_X1 U12593 ( .A1(n10185), .A2(n14166), .ZN(n10184) );
  AND2_X1 U12594 ( .A1(n10250), .A2(n10027), .ZN(n10248) );
  INV_X2 U12595 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20868) );
  NAND2_X1 U12596 ( .A1(n9796), .A2(n13607), .ZN(n9795) );
  AND2_X1 U12597 ( .A1(n15509), .A2(n15510), .ZN(n9749) );
  AND2_X1 U12598 ( .A1(n12299), .A2(n12298), .ZN(n9750) );
  AND2_X1 U12599 ( .A1(n14601), .A2(n10056), .ZN(n9751) );
  AND2_X1 U12600 ( .A1(n10009), .A2(n10012), .ZN(n9752) );
  OR2_X1 U12601 ( .A1(n19131), .A2(n15604), .ZN(n9753) );
  NAND2_X1 U12602 ( .A1(n16335), .A2(n16333), .ZN(n9754) );
  AND2_X1 U12603 ( .A1(n9741), .A2(n10830), .ZN(n9755) );
  INV_X1 U12604 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13525) );
  OR2_X1 U12605 ( .A1(n10481), .A2(n10079), .ZN(n10083) );
  NAND2_X1 U12606 ( .A1(n15903), .A2(n18771), .ZN(n18242) );
  AND2_X2 U12607 ( .A1(n12692), .A2(n19274), .ZN(n14998) );
  NAND2_X1 U12608 ( .A1(n16370), .A2(n16369), .ZN(n13556) );
  OR2_X1 U12609 ( .A1(n13073), .A2(n10166), .ZN(n13459) );
  AND4_X1 U12610 ( .A1(n10400), .A2(n12466), .A3(n10395), .A4(n10413), .ZN(
        n12456) );
  NOR2_X1 U12611 ( .A1(n13379), .A2(n13378), .ZN(n13442) );
  NAND2_X1 U12612 ( .A1(n10268), .A2(n9689), .ZN(n10271) );
  NAND2_X1 U12613 ( .A1(n10100), .A2(n12995), .ZN(n13010) );
  AND2_X1 U12614 ( .A1(n10264), .A2(n10014), .ZN(n10242) );
  INV_X1 U12615 ( .A(n20267), .ZN(n13226) );
  AND2_X1 U12616 ( .A1(n14968), .A2(n14887), .ZN(n9756) );
  AND2_X1 U12617 ( .A1(n14275), .A2(n14279), .ZN(n9757) );
  AND2_X1 U12618 ( .A1(n10171), .A2(n10169), .ZN(n9758) );
  AND2_X1 U12619 ( .A1(n9757), .A2(n10054), .ZN(n9759) );
  AND2_X1 U12620 ( .A1(n10089), .A2(n9756), .ZN(n9760) );
  AND2_X1 U12621 ( .A1(n10280), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10279) );
  AND2_X1 U12622 ( .A1(n10268), .A2(n10025), .ZN(n9761) );
  NAND2_X1 U12623 ( .A1(n10084), .A2(n10080), .ZN(n9762) );
  AND2_X1 U12624 ( .A1(n13125), .A2(n10085), .ZN(n9763) );
  INV_X1 U12625 ( .A(n19366), .ZN(n16361) );
  BUF_X1 U12626 ( .A(n10422), .Z(n13058) );
  OR2_X1 U12627 ( .A1(n10869), .A2(n10874), .ZN(n9764) );
  AND2_X1 U12628 ( .A1(n9661), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n9765) );
  XNOR2_X1 U12629 ( .A(n13282), .B(n13284), .ZN(n13281) );
  NAND2_X1 U12630 ( .A1(n10101), .A2(n10103), .ZN(n13627) );
  AND2_X1 U12631 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17833), .ZN(
        n9766) );
  INV_X1 U12632 ( .A(n10267), .ZN(n19162) );
  XNOR2_X1 U12633 ( .A(n10637), .B(n10621), .ZN(n13076) );
  AND2_X1 U12634 ( .A1(n10044), .A2(n10043), .ZN(n9767) );
  AND3_X1 U12635 ( .A1(n10095), .A2(n9683), .A3(n10097), .ZN(n13128) );
  NAND2_X1 U12636 ( .A1(n11066), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11298) );
  AND2_X1 U12637 ( .A1(n10022), .A2(n19145), .ZN(n9768) );
  AND2_X1 U12638 ( .A1(n9760), .A2(n10088), .ZN(n9769) );
  NAND2_X1 U12639 ( .A1(n10268), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10269) );
  INV_X1 U12640 ( .A(n13379), .ZN(n10101) );
  OR2_X1 U12641 ( .A1(n17849), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9770) );
  AND2_X1 U12642 ( .A1(n10264), .A2(n10015), .ZN(n9771) );
  AND2_X1 U12643 ( .A1(n9759), .A2(n10053), .ZN(n9772) );
  INV_X1 U12644 ( .A(n10867), .ZN(n12132) );
  OR2_X1 U12645 ( .A1(n10689), .A2(n10688), .ZN(n10867) );
  AND2_X1 U12646 ( .A1(n15156), .A2(n10023), .ZN(n9773) );
  AND2_X1 U12647 ( .A1(n10044), .A2(n10042), .ZN(n9774) );
  INV_X1 U12648 ( .A(n12161), .ZN(n10153) );
  INV_X1 U12649 ( .A(n15701), .ZN(n17046) );
  INV_X1 U12650 ( .A(n18794), .ZN(n9890) );
  AND2_X1 U12651 ( .A1(n11537), .A2(n11536), .ZN(n9775) );
  NAND2_X1 U12652 ( .A1(n10840), .A2(n10839), .ZN(n9776) );
  OR2_X1 U12653 ( .A1(n13387), .A2(n13301), .ZN(n13428) );
  INV_X1 U12654 ( .A(n13428), .ZN(n10040) );
  INV_X1 U12655 ( .A(n12433), .ZN(n9942) );
  OR2_X1 U12656 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9777) );
  AND2_X1 U12657 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .ZN(n9778) );
  AND2_X1 U12658 ( .A1(n9962), .A2(n17878), .ZN(n9779) );
  AND2_X1 U12659 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16966) );
  INV_X1 U12660 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9850) );
  INV_X1 U12661 ( .A(n20292), .ZN(n9821) );
  AND2_X1 U12662 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n9780) );
  AND4_X1 U12663 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n9781)
         );
  INV_X1 U12664 ( .A(n9855), .ZN(n9854) );
  NAND2_X1 U12665 ( .A1(n21110), .A2(n16472), .ZN(n9855) );
  AND2_X1 U12666 ( .A1(n9693), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9782) );
  AND2_X1 U12667 ( .A1(n10207), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9783) );
  INV_X1 U12668 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9844) );
  NOR2_X1 U12669 ( .A1(n20042), .A2(n19550), .ZN(n9784) );
  INV_X1 U12670 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20042) );
  NAND2_X2 U12671 ( .A1(n18946), .A2(n18932), .ZN(n18236) );
  INV_X1 U12672 ( .A(n17574), .ZN(n17573) );
  AOI22_X2 U12673 ( .A1(DATAI_19_), .A2(n9636), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n9637), .ZN(n20833) );
  AOI22_X2 U12674 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n9637), .B1(DATAI_17_), 
        .B2(n9636), .ZN(n20819) );
  AOI22_X2 U12675 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n9637), .B1(DATAI_20_), 
        .B2(n9636), .ZN(n20840) );
  AOI22_X2 U12676 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9637), .B1(DATAI_29_), 
        .B2(n9636), .ZN(n20777) );
  AOI22_X2 U12677 ( .A1(DATAI_16_), .A2(n9636), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n9637), .ZN(n20812) );
  AOI22_X2 U12678 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9637), .B1(DATAI_26_), 
        .B2(n9636), .ZN(n20759) );
  AOI22_X2 U12679 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n9637), .B1(DATAI_23_), 
        .B2(n9636), .ZN(n20866) );
  AOI21_X1 U12680 ( .B1(n10285), .B2(n10284), .A(n19929), .ZN(n10286) );
  NOR3_X2 U12681 ( .A1(n18616), .A2(n18539), .A3(n18397), .ZN(n18367) );
  AOI22_X2 U12682 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n9637), .B1(DATAI_22_), 
        .B2(n9636), .ZN(n20854) );
  NOR3_X2 U12683 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18616), .A3(
        n18490), .ZN(n18459) );
  NOR2_X2 U12684 ( .A1(n18878), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18616) );
  NOR2_X2 U12685 ( .A1(n18285), .A2(n18306), .ZN(n18669) );
  NAND2_X2 U12686 ( .A1(n9790), .A2(n12084), .ZN(n12110) );
  NAND2_X1 U12687 ( .A1(n9791), .A2(n10598), .ZN(n9790) );
  NAND3_X1 U12688 ( .A1(n9713), .A2(n12067), .A3(n9638), .ZN(n9791) );
  NOR2_X2 U12689 ( .A1(n9795), .A2(n9794), .ZN(n13655) );
  AND2_X2 U12691 ( .A1(n15111), .A2(n9783), .ZN(n12508) );
  NOR2_X2 U12692 ( .A1(n15179), .A2(n9956), .ZN(n15111) );
  AOI21_X1 U12693 ( .B1(n15862), .B2(n15861), .A(n15860), .ZN(n17847) );
  AOI22_X1 U12694 ( .A1(n15860), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n15861), .B2(n9812), .ZN(n9811) );
  INV_X1 U12695 ( .A(n9813), .ZN(n18127) );
  NAND3_X1 U12696 ( .A1(n15789), .A2(n15791), .A3(n15790), .ZN(n15985) );
  INV_X2 U12697 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18891) );
  INV_X2 U12698 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18909) );
  NAND3_X2 U12699 ( .A1(n11041), .A2(n11946), .A3(n9815), .ZN(n11060) );
  NOR2_X1 U12700 ( .A1(n9816), .A2(n9731), .ZN(n9815) );
  NAND3_X2 U12701 ( .A1(n10055), .A2(n9817), .A3(n13352), .ZN(n11946) );
  INV_X1 U12702 ( .A(n11063), .ZN(n9817) );
  NAND4_X1 U12703 ( .A1(n13029), .A2(n12869), .A3(n20292), .A4(n20246), .ZN(
        n12723) );
  INV_X1 U12704 ( .A(n14493), .ZN(n9823) );
  NAND2_X1 U12705 ( .A1(n10060), .A2(n9822), .ZN(n14505) );
  NAND3_X1 U12706 ( .A1(n9827), .A2(n9826), .A3(n14428), .ZN(n9825) );
  INV_X1 U12707 ( .A(n14628), .ZN(n9829) );
  NAND2_X1 U12708 ( .A1(n14463), .A2(n9833), .ZN(n9832) );
  NAND2_X1 U12709 ( .A1(n9714), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9831) );
  INV_X1 U12710 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9833) );
  INV_X2 U12711 ( .A(n11129), .ZN(n11917) );
  AND2_X2 U12712 ( .A1(n10911), .A2(n10908), .ZN(n11129) );
  AND2_X2 U12713 ( .A1(n10052), .A2(n10910), .ZN(n10908) );
  AND2_X2 U12714 ( .A1(n10051), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10911) );
  OAI21_X1 U12715 ( .B1(n20328), .B2(n14429), .A(n13034), .ZN(n13048) );
  XNOR2_X2 U12716 ( .A(n11202), .B(n11201), .ZN(n20328) );
  NAND2_X2 U12717 ( .A1(n11147), .A2(n11146), .ZN(n11202) );
  NAND3_X1 U12718 ( .A1(n10946), .A2(n11965), .A3(n20267), .ZN(n10967) );
  NAND2_X2 U12719 ( .A1(n10921), .A2(n9699), .ZN(n20267) );
  NAND2_X1 U12720 ( .A1(n15885), .A2(n18192), .ZN(n9837) );
  NAND2_X1 U12721 ( .A1(n9835), .A2(n15885), .ZN(n17871) );
  NAND2_X1 U12722 ( .A1(n17882), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9835) );
  INV_X1 U12723 ( .A(n15885), .ZN(n9838) );
  NOR2_X2 U12724 ( .A1(n9841), .A2(n9840), .ZN(n17619) );
  INV_X1 U12725 ( .A(n9847), .ZN(n17634) );
  NAND2_X1 U12726 ( .A1(n9847), .A2(n17849), .ZN(n17618) );
  NAND3_X1 U12727 ( .A1(n15797), .A2(n15800), .A3(n9732), .ZN(n9848) );
  NAND2_X1 U12728 ( .A1(n17595), .A2(n9853), .ZN(n9856) );
  NOR2_X1 U12729 ( .A1(n9855), .A2(n17833), .ZN(n9853) );
  NAND3_X1 U12730 ( .A1(n9864), .A2(n15905), .A3(n18043), .ZN(n15910) );
  INV_X1 U12731 ( .A(n9864), .ZN(n17848) );
  OAI21_X2 U12732 ( .B1(n12519), .B2(n12520), .A(n9866), .ZN(n9865) );
  NAND4_X1 U12733 ( .A1(n10152), .A2(n10151), .A3(n12110), .A4(n12109), .ZN(
        n12187) );
  AND2_X2 U12734 ( .A1(n9977), .A2(n12121), .ZN(n12109) );
  NAND4_X1 U12735 ( .A1(n12158), .A2(n12155), .A3(n12156), .A4(n12157), .ZN(
        n9874) );
  INV_X1 U12736 ( .A(n10467), .ZN(n9879) );
  NAND2_X1 U12737 ( .A1(n9875), .A2(n12038), .ZN(n9878) );
  NAND2_X1 U12738 ( .A1(n10468), .A2(n10467), .ZN(n9875) );
  NAND2_X1 U12739 ( .A1(n10468), .A2(n10467), .ZN(n10483) );
  NAND2_X1 U12740 ( .A1(n9877), .A2(n10468), .ZN(n9876) );
  NOR2_X1 U12741 ( .A1(n12038), .A2(n9879), .ZN(n9877) );
  NAND3_X1 U12742 ( .A1(n12199), .A2(n12188), .A3(n9942), .ZN(n9940) );
  NAND2_X2 U12743 ( .A1(n12792), .A2(n9883), .ZN(n17404) );
  NAND4_X1 U12744 ( .A1(n9895), .A2(n9778), .A3(P3_EAX_REG_0__SCAN_IN), .A4(
        P3_EAX_REG_2__SCAN_IN), .ZN(n9894) );
  INV_X2 U12745 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18883) );
  NAND2_X1 U12746 ( .A1(n12871), .A2(n9898), .ZN(n9896) );
  NOR2_X2 U12747 ( .A1(n11012), .A2(n9900), .ZN(n11017) );
  OR2_X2 U12748 ( .A1(n9903), .A2(n10998), .ZN(n20272) );
  OAI21_X1 U12749 ( .B1(n14596), .B2(n10036), .A(n10067), .ZN(n14566) );
  NAND2_X1 U12750 ( .A1(n12056), .A2(n9915), .ZN(n9953) );
  INV_X1 U12751 ( .A(n12040), .ZN(n9914) );
  NAND2_X1 U12752 ( .A1(n9700), .A2(n9917), .ZN(n9916) );
  AND2_X1 U12753 ( .A1(n9919), .A2(n12941), .ZN(n19487) );
  NAND2_X1 U12754 ( .A1(n9700), .A2(n12069), .ZN(n12142) );
  XNOR2_X1 U12755 ( .A(n9923), .B(n15265), .ZN(n15543) );
  NAND3_X1 U12756 ( .A1(n9927), .A2(n9930), .A3(n15165), .ZN(n9926) );
  NAND2_X1 U12757 ( .A1(n9939), .A2(n9753), .ZN(n12304) );
  NAND3_X1 U12758 ( .A1(n12199), .A2(n9941), .A3(n12188), .ZN(n9939) );
  NAND2_X1 U12759 ( .A1(n15213), .A2(n9947), .ZN(n9943) );
  AOI21_X1 U12760 ( .B1(n15213), .B2(n9949), .A(n9951), .ZN(n15187) );
  NAND2_X1 U12761 ( .A1(n15213), .A2(n15167), .ZN(n15212) );
  NAND2_X1 U12762 ( .A1(n15251), .A2(n10211), .ZN(n15227) );
  NAND2_X1 U12763 ( .A1(n15251), .A2(n15508), .ZN(n15245) );
  NAND3_X1 U12764 ( .A1(n17878), .A2(n9962), .A3(n16819), .ZN(n17739) );
  NAND3_X1 U12765 ( .A1(n17878), .A2(n9962), .A3(n9739), .ZN(n17728) );
  NAND4_X1 U12766 ( .A1(n10373), .A2(n10372), .A3(n10370), .A4(n10371), .ZN(
        n9973) );
  NAND4_X1 U12767 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n9975) );
  NAND4_X1 U12768 ( .A1(n9976), .A2(n12104), .A3(n9730), .A4(n12105), .ZN(
        n9977) );
  NAND2_X1 U12769 ( .A1(n9978), .A2(n9982), .ZN(n9981) );
  INV_X1 U12770 ( .A(n12299), .ZN(n9978) );
  INV_X1 U12771 ( .A(n12304), .ZN(n9979) );
  NAND2_X1 U12772 ( .A1(n9980), .A2(n9982), .ZN(n15287) );
  NAND2_X1 U12773 ( .A1(n9984), .A2(n12299), .ZN(n9980) );
  NAND2_X1 U12774 ( .A1(n15148), .A2(n9998), .ZN(n9997) );
  NAND2_X1 U12775 ( .A1(n14861), .A2(n19145), .ZN(n10009) );
  OR2_X1 U12776 ( .A1(n14861), .A2(n14862), .ZN(n10013) );
  NAND2_X1 U12777 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10018) );
  NAND3_X1 U12778 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n10017), .A3(
        n10019), .ZN(n10255) );
  NAND3_X1 U12779 ( .A1(n10019), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U12780 ( .A1(n19000), .A2(n9773), .ZN(n10021) );
  NAND2_X1 U12781 ( .A1(n10021), .A2(n10020), .ZN(n14915) );
  NAND2_X1 U12782 ( .A1(n10268), .A2(n10024), .ZN(n10275) );
  NAND3_X1 U12783 ( .A1(n10035), .A2(n10034), .A3(n10032), .ZN(n10031) );
  NAND2_X1 U12784 ( .A1(n11337), .A2(n10039), .ZN(n14403) );
  OR2_X1 U12785 ( .A1(n11297), .A2(n11296), .ZN(n10039) );
  NAND2_X1 U12786 ( .A1(n13428), .A2(n13429), .ZN(n10043) );
  NOR2_X2 U12787 ( .A1(n13604), .A2(n13603), .ZN(n14224) );
  INV_X2 U12788 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10052) );
  NAND3_X1 U12789 ( .A1(n14493), .A2(n14532), .A3(n9751), .ZN(n10060) );
  NAND4_X1 U12790 ( .A1(n11066), .A2(n11040), .A3(n11965), .A4(n11047), .ZN(
        n11050) );
  NAND2_X2 U12791 ( .A1(n9708), .A2(n9639), .ZN(n11047) );
  NAND2_X2 U12792 ( .A1(n10061), .A2(n9710), .ZN(n11965) );
  INV_X2 U12793 ( .A(n20285), .ZN(n11066) );
  NAND2_X1 U12794 ( .A1(n11060), .A2(n10065), .ZN(n10064) );
  NAND3_X1 U12795 ( .A1(n10064), .A2(n11062), .A3(n10063), .ZN(n11106) );
  NAND2_X1 U12796 ( .A1(n11070), .A2(n12972), .ZN(n10066) );
  AND3_X4 U12797 ( .A1(n9640), .A2(n15620), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10586) );
  INV_X1 U12798 ( .A(n15001), .ZN(n10076) );
  NAND3_X1 U12799 ( .A1(n10078), .A2(n13003), .A3(n13118), .ZN(n10077) );
  INV_X1 U12800 ( .A(n13003), .ZN(n10079) );
  NAND2_X1 U12801 ( .A1(n13125), .A2(n9738), .ZN(n13479) );
  NAND2_X1 U12802 ( .A1(n10422), .A2(n10406), .ZN(n10090) );
  NAND2_X1 U12803 ( .A1(n10222), .A2(n10224), .ZN(n10091) );
  INV_X1 U12804 ( .A(n10577), .ZN(n10092) );
  AND3_X2 U12805 ( .A1(n13713), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10591) );
  CLKBUF_X1 U12806 ( .A(n10099), .Z(n10095) );
  NAND2_X1 U12807 ( .A1(n12996), .A2(n12995), .ZN(n10098) );
  NAND3_X1 U12808 ( .A1(n10099), .A2(n10096), .A3(n10098), .ZN(n13208) );
  CLKBUF_X1 U12809 ( .A(n10098), .Z(n10097) );
  NAND3_X1 U12810 ( .A1(n10095), .A2(n13009), .A3(n10097), .ZN(n13127) );
  NAND2_X1 U12811 ( .A1(n10111), .A2(n10109), .ZN(P2_U2892) );
  NAND2_X1 U12812 ( .A1(n15040), .A2(n19269), .ZN(n10111) );
  AND2_X1 U12813 ( .A1(n14947), .A2(n14946), .ZN(n10112) );
  NAND2_X1 U12814 ( .A1(n10114), .A2(n19355), .ZN(n12535) );
  OAI21_X1 U12815 ( .B1(n10117), .B2(n15597), .A(n10115), .ZN(P2_U3015) );
  NOR2_X2 U12816 ( .A1(n15920), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17595) );
  NAND2_X2 U12817 ( .A1(n10129), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18125) );
  NAND2_X2 U12818 ( .A1(n12346), .A2(n12435), .ZN(n12343) );
  NOR3_X2 U12819 ( .A1(n12384), .A2(n12391), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n12408) );
  OR2_X2 U12820 ( .A1(n12384), .A2(n12391), .ZN(n12395) );
  NAND3_X1 U12821 ( .A1(n10415), .A2(n10416), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10146) );
  NOR2_X1 U12822 ( .A1(n15636), .A2(n19175), .ZN(n10147) );
  NAND4_X1 U12823 ( .A1(n10150), .A2(n9737), .A3(n10413), .A4(n12243), .ZN(
        n10414) );
  AND2_X1 U12825 ( .A1(n10152), .A2(n12161), .ZN(n12162) );
  NAND2_X1 U12826 ( .A1(n12110), .A2(n12109), .ZN(n12133) );
  AND3_X2 U12827 ( .A1(n12110), .A2(n12109), .A3(n10867), .ZN(n12163) );
  INV_X1 U12828 ( .A(n15152), .ZN(n10157) );
  NAND2_X1 U12829 ( .A1(n10158), .A2(n12383), .ZN(n15155) );
  OR2_X1 U12830 ( .A1(n15161), .A2(n12368), .ZN(n10158) );
  NAND2_X1 U12831 ( .A1(n10620), .A2(n10161), .ZN(n10636) );
  NAND2_X1 U12832 ( .A1(n10162), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10161) );
  NOR2_X1 U12833 ( .A1(n13072), .A2(n13071), .ZN(n13073) );
  NOR2_X1 U12834 ( .A1(n13073), .A2(n10656), .ZN(n13460) );
  INV_X1 U12835 ( .A(n10174), .ZN(n15048) );
  INV_X1 U12836 ( .A(n15047), .ZN(n10173) );
  NAND2_X1 U12837 ( .A1(n15509), .A2(n9755), .ZN(n15094) );
  NAND2_X1 U12838 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10177) );
  INV_X1 U12839 ( .A(n10179), .ZN(n10178) );
  INV_X1 U12840 ( .A(n14271), .ZN(n10180) );
  NAND2_X1 U12841 ( .A1(n10180), .A2(n10181), .ZN(n14257) );
  NAND3_X1 U12842 ( .A1(n13421), .A2(n13432), .A3(n11336), .ZN(n13534) );
  NOR2_X2 U12843 ( .A1(n13304), .A2(n13423), .ZN(n13421) );
  NAND2_X1 U12844 ( .A1(n13368), .A2(n11193), .ZN(n10186) );
  NAND2_X1 U12845 ( .A1(n10186), .A2(n10188), .ZN(n13386) );
  INV_X1 U12846 ( .A(n13386), .ZN(n10187) );
  NAND2_X1 U12847 ( .A1(n10187), .A2(n11210), .ZN(n13383) );
  NAND2_X1 U12849 ( .A1(n14137), .A2(n10197), .ZN(n14099) );
  AND2_X1 U12850 ( .A1(n14137), .A2(n9745), .ZN(n14110) );
  AND2_X1 U12851 ( .A1(n14137), .A2(n14136), .ZN(n14123) );
  NOR2_X4 U12852 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13177) );
  XNOR2_X2 U12853 ( .A(n10198), .B(n11074), .ZN(n20369) );
  AND2_X1 U12855 ( .A1(n15111), .A2(n10209), .ZN(n12566) );
  NAND2_X1 U12856 ( .A1(n15111), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15104) );
  INV_X1 U12857 ( .A(n13208), .ZN(n13209) );
  INV_X4 U12858 ( .A(n12253), .ZN(n13839) );
  AOI21_X1 U12859 ( .B1(n9667), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U12860 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U12861 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9667), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U12862 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10340) );
  INV_X2 U12863 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10914) );
  NAND2_X1 U12864 ( .A1(n13927), .A2(n13926), .ZN(n13928) );
  AND3_X1 U12865 ( .A1(n11963), .A2(n13029), .A3(n11964), .ZN(n13035) );
  NOR2_X1 U12866 ( .A1(n12075), .A2(n12074), .ZN(n12139) );
  AOI22_X1 U12867 ( .A1(n11003), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10957), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11023) );
  NOR2_X1 U12868 ( .A1(n12134), .A2(n12099), .ZN(n12101) );
  NOR2_X1 U12869 ( .A1(n12134), .A2(n12048), .ZN(n12049) );
  AOI22_X1 U12870 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12152), .B1(
        n19429), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U12871 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9655), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10305) );
  AOI21_X1 U12872 ( .B1(n14461), .B2(n16140), .A(n14460), .ZN(n14462) );
  NAND2_X1 U12873 ( .A1(n14461), .A2(n12020), .ZN(n12037) );
  INV_X2 U12874 ( .A(n13156), .ZN(n14389) );
  AND2_X1 U12875 ( .A1(n15323), .A2(n15329), .ZN(n10214) );
  NAND2_X1 U12876 ( .A1(n17939), .A2(n17782), .ZN(n17648) );
  INV_X1 U12877 ( .A(n17648), .ZN(n17689) );
  NOR2_X1 U12878 ( .A1(n20541), .A2(n20252), .ZN(n10215) );
  NAND2_X2 U12879 ( .A1(n14389), .A2(n13155), .ZN(n14396) );
  AND2_X1 U12880 ( .A1(n10892), .A2(n9734), .ZN(n10216) );
  AND4_X1 U12881 ( .A1(n12174), .A2(n12173), .A3(n12172), .A4(n12171), .ZN(
        n10217) );
  AND4_X1 U12882 ( .A1(n12149), .A2(n12148), .A3(n12147), .A4(n12146), .ZN(
        n10218) );
  AND2_X1 U12883 ( .A1(n10296), .A2(n10295), .ZN(n10219) );
  AND3_X1 U12884 ( .A1(n10303), .A2(n10383), .A3(n10302), .ZN(n10220) );
  AND2_X1 U12885 ( .A1(n10305), .A2(n10304), .ZN(n10221) );
  AND3_X1 U12886 ( .A1(n9660), .A2(n19411), .A3(n19422), .ZN(n10222) );
  OR2_X1 U12887 ( .A1(n16677), .A2(n16664), .ZN(n10223) );
  INV_X1 U12888 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10240) );
  INV_X1 U12889 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17808) );
  AND2_X1 U12890 ( .A1(n12468), .A2(n10392), .ZN(n10224) );
  OR2_X1 U12891 ( .A1(n14055), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10225) );
  OR3_X1 U12892 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17666), .ZN(n10226) );
  INV_X1 U12893 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11383) );
  INV_X1 U12894 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16042) );
  AOI22_X1 U12895 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10297) );
  INV_X1 U12896 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10239) );
  OR2_X1 U12897 ( .A1(n14055), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10227) );
  INV_X1 U12898 ( .A(n13370), .ZN(n11234) );
  AND2_X1 U12899 ( .A1(n13906), .A2(n13924), .ZN(n10228) );
  INV_X1 U12900 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10561) );
  INV_X1 U12901 ( .A(n10977), .ZN(n11091) );
  OR2_X1 U12902 ( .A1(n10772), .A2(n10771), .ZN(n13210) );
  OR2_X1 U12903 ( .A1(n18958), .A2(n10406), .ZN(n16324) );
  INV_X1 U12904 ( .A(n16324), .ZN(n19355) );
  INV_X1 U12905 ( .A(n12115), .ZN(n12112) );
  INV_X1 U12906 ( .A(n10957), .ZN(n11697) );
  AND2_X1 U12907 ( .A1(n12615), .A2(n19926), .ZN(n19348) );
  INV_X1 U12908 ( .A(n19348), .ZN(n19129) );
  OR2_X1 U12909 ( .A1(n10797), .A2(n10796), .ZN(n13444) );
  AND2_X1 U12910 ( .A1(n12242), .A2(n12237), .ZN(n10231) );
  NAND2_X1 U12911 ( .A1(n10412), .A2(n12237), .ZN(n10232) );
  AND3_X1 U12912 ( .A1(n20662), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10233) );
  INV_X1 U12913 ( .A(n10401), .ZN(n12711) );
  AND2_X1 U12914 ( .A1(n11662), .A2(n11661), .ZN(n10234) );
  INV_X1 U12915 ( .A(n14256), .ZN(n14264) );
  INV_X1 U12916 ( .A(n14207), .ZN(n11411) );
  AND2_X1 U12917 ( .A1(n12556), .A2(n10856), .ZN(n10236) );
  AND4_X1 U12918 ( .A1(n12179), .A2(n12178), .A3(n12177), .A4(n12176), .ZN(
        n10237) );
  NAND2_X1 U12919 ( .A1(n13651), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10238) );
  INV_X1 U12920 ( .A(n11021), .ZN(n11090) );
  INV_X1 U12921 ( .A(n11130), .ZN(n11082) );
  NAND2_X1 U12922 ( .A1(n12154), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12098) );
  OAI22_X1 U12923 ( .A1(n19700), .A2(n12070), .B1(n12942), .B2(n12142), .ZN(
        n12071) );
  OR2_X1 U12924 ( .A1(n11989), .A2(n11978), .ZN(n12000) );
  INV_X1 U12925 ( .A(n10407), .ZN(n10408) );
  INV_X1 U12926 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11811) );
  AOI21_X1 U12927 ( .B1(n9659), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A(n10929), .ZN(n10933) );
  NAND2_X1 U12928 ( .A1(n13226), .A2(n10965), .ZN(n10966) );
  AND2_X1 U12929 ( .A1(n20696), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11967) );
  OR3_X1 U12930 ( .A1(n11956), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n20240), .ZN(n11999) );
  INV_X1 U12931 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11731) );
  OR2_X1 U12932 ( .A1(n11325), .A2(n11324), .ZN(n14419) );
  OR2_X1 U12933 ( .A1(n11293), .A2(n11292), .ZN(n14412) );
  NAND2_X1 U12934 ( .A1(n11202), .A2(n11201), .ZN(n11153) );
  OR2_X1 U12935 ( .A1(n10566), .A2(n10565), .ZN(n10563) );
  AOI22_X1 U12936 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9666), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10345) );
  NAND2_X1 U12937 ( .A1(n12083), .A2(n10406), .ZN(n12084) );
  AOI22_X1 U12938 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10290) );
  INV_X1 U12939 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11905) );
  INV_X1 U12940 ( .A(n14155), .ZN(n11745) );
  OR2_X1 U12942 ( .A1(n11171), .A2(n11170), .ZN(n13269) );
  OR2_X1 U12943 ( .A1(n16112), .A2(n16214), .ZN(n14438) );
  OR2_X1 U12944 ( .A1(n11266), .A2(n11265), .ZN(n13503) );
  INV_X1 U12945 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12964) );
  OR2_X1 U12946 ( .A1(n10952), .A2(n10951), .ZN(n10953) );
  AND2_X1 U12947 ( .A1(n14979), .A2(n13868), .ZN(n13848) );
  NOR2_X1 U12948 ( .A1(n13008), .A2(n12942), .ZN(n12943) );
  INV_X1 U12949 ( .A(n13890), .ZN(n13891) );
  AOI22_X1 U12950 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10368) );
  INV_X1 U12951 ( .A(n11663), .ZN(n11664) );
  INV_X1 U12952 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11684) );
  OR2_X1 U12953 ( .A1(n15989), .A2(n11935), .ZN(n11714) );
  NAND2_X1 U12954 ( .A1(n21148), .A2(n11411), .ZN(n14208) );
  INV_X1 U12955 ( .A(n14222), .ZN(n11405) );
  NAND2_X1 U12956 ( .A1(n11340), .A2(n11339), .ZN(n14409) );
  AND2_X1 U12957 ( .A1(n14007), .A2(n14006), .ZN(n14198) );
  INV_X1 U12958 ( .A(n11047), .ZN(n13238) );
  NOR2_X1 U12959 ( .A1(n11994), .A2(n14429), .ZN(n11998) );
  AND2_X1 U12960 ( .A1(n20632), .A2(n10895), .ZN(n20249) );
  INV_X1 U12961 ( .A(n11994), .ZN(n12003) );
  AND2_X1 U12962 ( .A1(n10572), .A2(n10564), .ZN(n12209) );
  INV_X1 U12963 ( .A(n10248), .ZN(n10260) );
  NAND2_X1 U12964 ( .A1(n12060), .A2(n12727), .ZN(n12893) );
  INV_X1 U12965 ( .A(n13869), .ZN(n13870) );
  NAND2_X1 U12966 ( .A1(n12423), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12424) );
  INV_X1 U12967 ( .A(n17636), .ZN(n16652) );
  NAND2_X1 U12968 ( .A1(n17833), .A2(n18073), .ZN(n15908) );
  NOR2_X1 U12969 ( .A1(n13685), .A2(n13684), .ZN(n13689) );
  AND2_X1 U12970 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15850), .ZN(
        n15851) );
  INV_X1 U12971 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n21083) );
  INV_X1 U12972 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n20994) );
  NOR2_X1 U12973 ( .A1(n11863), .A2(n14489), .ZN(n11864) );
  AND2_X1 U12974 ( .A1(n11664), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11665) );
  INV_X1 U12975 ( .A(n13385), .ZN(n11210) );
  OAI22_X1 U12976 ( .A1(n11031), .A2(n11695), .B1(n11002), .B2(n11684), .ZN(
        n11007) );
  OR2_X1 U12977 ( .A1(n14475), .A2(n11935), .ZN(n11899) );
  INV_X1 U12978 ( .A(n11273), .ZN(n11274) );
  INV_X1 U12979 ( .A(n11298), .ZN(n11513) );
  AND2_X1 U12980 ( .A1(n14728), .A2(n14640), .ZN(n14687) );
  AND2_X1 U12981 ( .A1(n14802), .A2(n14639), .ZN(n14728) );
  AND2_X1 U12982 ( .A1(n13438), .A2(n13437), .ZN(n13439) );
  NAND2_X1 U12983 ( .A1(n11965), .A2(n20262), .ZN(n14429) );
  OAI21_X1 U12984 ( .B1(n11994), .B2(n11699), .A(n11152), .ZN(n11201) );
  AND3_X1 U12985 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20868), .A3(n20245), 
        .ZN(n20293) );
  AND2_X1 U12986 ( .A1(n12360), .A2(n12359), .ZN(n19053) );
  INV_X1 U12987 ( .A(n12441), .ZN(n10557) );
  NAND2_X1 U12988 ( .A1(n10412), .A2(n10402), .ZN(n13008) );
  INV_X1 U12989 ( .A(n15060), .ZN(n10846) );
  OAI211_X1 U12990 ( .C1(n12506), .C2(n15312), .A(n15311), .B(n9712), .ZN(
        n15313) );
  OR2_X1 U12991 ( .A1(n19370), .A2(n19362), .ZN(n15565) );
  XNOR2_X1 U12992 ( .A(n12042), .B(n12041), .ZN(n12043) );
  NAND2_X1 U12993 ( .A1(n12235), .A2(n19281), .ZN(n12236) );
  NOR2_X1 U12994 ( .A1(n18944), .A2(n18277), .ZN(n16640) );
  INV_X2 U12995 ( .A(n15648), .ZN(n15804) );
  NAND2_X1 U12996 ( .A1(n15911), .A2(n15908), .ZN(n15909) );
  NAND2_X1 U12997 ( .A1(n18729), .A2(n15747), .ZN(n18749) );
  NAND3_X1 U12998 ( .A1(n12784), .A2(n12783), .A3(n12782), .ZN(n15864) );
  INV_X1 U12999 ( .A(n14073), .ZN(n12949) );
  NAND2_X1 U13000 ( .A1(n11665), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11746) );
  NOR2_X1 U13001 ( .A1(n13349), .A2(n11043), .ZN(n13359) );
  OR2_X1 U13002 ( .A1(n11805), .A2(n14498), .ZN(n11863) );
  OR2_X1 U13003 ( .A1(n11558), .A2(n16042), .ZN(n11578) );
  INV_X1 U13004 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16057) );
  INV_X1 U13005 ( .A(n11429), .ZN(n11449) );
  AND2_X1 U13006 ( .A1(n11301), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11328) );
  AND2_X1 U13007 ( .A1(n12011), .A2(n12010), .ZN(n13231) );
  AND2_X1 U13008 ( .A1(n20507), .A2(n20506), .ZN(n20533) );
  INV_X1 U13009 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20662) );
  NOR2_X1 U13010 ( .A1(n20414), .A2(n20413), .ZN(n20742) );
  AOI21_X1 U13011 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20696), .A(n20413), 
        .ZN(n20806) );
  XNOR2_X1 U13012 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12865) );
  NAND2_X1 U13013 ( .A1(n12224), .A2(n12221), .ZN(n12466) );
  INV_X1 U13014 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19087) );
  INV_X1 U13015 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15302) );
  OR2_X1 U13016 ( .A1(n10745), .A2(n10744), .ZN(n13011) );
  OR2_X1 U13017 ( .A1(n12477), .A2(n16393), .ZN(n15458) );
  NAND2_X1 U13018 ( .A1(n12238), .A2(n12236), .ZN(n16394) );
  NAND2_X1 U13019 ( .A1(n19630), .A2(n19629), .ZN(n19608) );
  OR3_X1 U13020 ( .A1(n12150), .A2(n19744), .A3(n20035), .ZN(n19727) );
  OR2_X1 U13021 ( .A1(n20019), .A2(n20028), .ZN(n19788) );
  OR2_X1 U13022 ( .A1(n12701), .A2(n12700), .ZN(n16402) );
  NOR2_X1 U13023 ( .A1(n17581), .A2(n16687), .ZN(n16686) );
  NOR2_X1 U13024 ( .A1(n17690), .A2(n16774), .ZN(n16773) );
  NOR2_X1 U13025 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16882), .ZN(n16869) );
  NAND4_X1 U13026 ( .A1(n16640), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n18929), 
        .A4(n16639), .ZN(n16997) );
  NOR2_X1 U13027 ( .A1(n16813), .A2(n17174), .ZN(n17150) );
  INV_X1 U13028 ( .A(n17934), .ZN(n17877) );
  NOR2_X1 U13029 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17833), .ZN(
        n17721) );
  INV_X1 U13030 ( .A(n17832), .ZN(n17822) );
  INV_X1 U13031 ( .A(n17849), .ZN(n17833) );
  INV_X1 U13032 ( .A(n15874), .ZN(n15875) );
  INV_X1 U13033 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18539) );
  INV_X1 U13034 ( .A(n13683), .ZN(n18289) );
  OR2_X1 U13035 ( .A1(n13036), .A2(n12723), .ZN(n12857) );
  NAND2_X1 U13036 ( .A1(n11579), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11617) );
  NOR2_X2 U13037 ( .A1(n14459), .A2(n13345), .ZN(n20119) );
  INV_X1 U13038 ( .A(n20111), .ZN(n20139) );
  INV_X1 U13039 ( .A(n14074), .ZN(n14075) );
  INV_X1 U13040 ( .A(n20161), .ZN(n14296) );
  NOR2_X1 U13041 ( .A1(n14304), .A2(n19420), .ZN(n12034) );
  NAND2_X1 U13042 ( .A1(n12019), .A2(n13235), .ZN(n13156) );
  AND2_X1 U13043 ( .A1(n11863), .A2(n11806), .ZN(n14502) );
  AND2_X1 U13044 ( .A1(n14289), .A2(n14290), .ZN(n14291) );
  AND2_X1 U13045 ( .A1(n16144), .A2(n13049), .ZN(n16138) );
  AND2_X1 U13046 ( .A1(n13236), .A2(n13235), .ZN(n13256) );
  INV_X1 U13047 ( .A(n14798), .ZN(n16221) );
  NOR2_X1 U13048 ( .A1(n16197), .A2(n13293), .ZN(n20223) );
  AND2_X1 U13049 ( .A1(n13290), .A2(n14783), .ZN(n13293) );
  NOR2_X1 U13050 ( .A1(n20669), .A2(n13231), .ZN(n15956) );
  OAI22_X1 U13051 ( .A1(n20259), .A2(n20258), .B1(n20600), .B2(n20408), .ZN(
        n20297) );
  INV_X1 U13052 ( .A(n20364), .ZN(n20323) );
  OAI22_X1 U13053 ( .A1(n20337), .A2(n20336), .B1(n20600), .B2(n20472), .ZN(
        n20360) );
  OR2_X1 U13054 ( .A1(n9665), .A2(n20328), .ZN(n20445) );
  NAND2_X1 U13055 ( .A1(n13371), .A2(n13368), .ZN(n20371) );
  OAI221_X1 U13056 ( .B1(n20431), .B2(n20669), .C1(n20431), .C2(n20415), .A(
        n20742), .ZN(n20433) );
  OAI22_X1 U13057 ( .A1(n20474), .A2(n20473), .B1(n20472), .B2(n20731), .ZN(
        n20497) );
  NOR2_X1 U13058 ( .A1(n13368), .A2(n11234), .ZN(n20502) );
  INV_X1 U13059 ( .A(n20540), .ZN(n20563) );
  INV_X1 U13060 ( .A(n20405), .ZN(n20661) );
  AND2_X1 U13061 ( .A1(n9665), .A2(n20328), .ZN(n20734) );
  OAI22_X1 U13062 ( .A1(n20673), .A2(n20672), .B1(n20731), .B2(n20671), .ZN(
        n20689) );
  INV_X1 U13063 ( .A(n20637), .ZN(n20631) );
  AND2_X1 U13064 ( .A1(n20735), .A2(n20734), .ZN(n20861) );
  AND2_X1 U13065 ( .A1(n9665), .A2(n20244), .ZN(n20630) );
  INV_X1 U13066 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20867) );
  AND2_X1 U13067 ( .A1(n19145), .A2(n19178), .ZN(n16280) );
  INV_X1 U13068 ( .A(n16281), .ZN(n10287) );
  NAND2_X1 U13069 ( .A1(n16272), .A2(n10885), .ZN(n19183) );
  INV_X1 U13070 ( .A(n19188), .ZN(n19170) );
  OR2_X1 U13071 ( .A1(n10785), .A2(n10784), .ZN(n13380) );
  AND2_X1 U13072 ( .A1(n19239), .A2(n12716), .ZN(n19207) );
  INV_X1 U13073 ( .A(n19239), .ZN(n19264) );
  INV_X1 U13074 ( .A(n19276), .ZN(n12683) );
  AND2_X1 U13075 ( .A1(n15251), .A2(n15549), .ZN(n15285) );
  AND2_X1 U13076 ( .A1(n16375), .A2(n12499), .ZN(n15592) );
  NOR2_X1 U13077 ( .A1(n15610), .A2(n15617), .ZN(n16375) );
  INV_X1 U13078 ( .A(n19754), .ZN(n19868) );
  OAI21_X1 U13079 ( .B1(n19389), .B2(n19388), .A(n19387), .ZN(n19425) );
  NOR2_X1 U13080 ( .A1(n19572), .A2(n20007), .ZN(n19507) );
  AND2_X1 U13081 ( .A1(n19520), .A2(n19515), .ZN(n19539) );
  OR3_X1 U13082 ( .A1(n19579), .A2(n19754), .A3(n19578), .ZN(n19597) );
  NOR2_X1 U13083 ( .A1(n19814), .A2(n19572), .ZN(n19625) );
  NAND2_X1 U13084 ( .A1(n19639), .A2(n19638), .ZN(n19656) );
  INV_X1 U13085 ( .A(n19684), .ZN(n19685) );
  AND2_X1 U13086 ( .A1(n19727), .A2(n19725), .ZN(n19745) );
  NOR2_X1 U13087 ( .A1(n19815), .A2(n19788), .ZN(n19805) );
  INV_X1 U13088 ( .A(n19891), .ZN(n19837) );
  AND2_X1 U13089 ( .A1(n12935), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19913) );
  INV_X1 U13090 ( .A(n18944), .ZN(n18945) );
  NOR2_X1 U13091 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16769), .ZN(n16755) );
  NOR2_X1 U13092 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16787), .ZN(n16775) );
  NOR3_X1 U13093 ( .A1(n17018), .A2(n18838), .A3(n16803), .ZN(n16800) );
  NOR2_X1 U13094 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16887), .ZN(n16886) );
  NOR2_X1 U13095 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16936), .ZN(n16903) );
  INV_X1 U13096 ( .A(n17014), .ZN(n16940) );
  NOR4_X2 U13097 ( .A1(n18151), .A2(n18945), .A3(n17006), .A4(n18769), .ZN(
        n16999) );
  NOR2_X1 U13098 ( .A1(n16756), .A2(n17104), .ZN(n17086) );
  AND3_X1 U13099 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(n17278), .ZN(n17245) );
  NOR2_X1 U13100 ( .A1(n17291), .A2(n17295), .ZN(n17290) );
  NAND4_X1 U13101 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .A3(n17314), .A4(n17301), .ZN(n17295) );
  INV_X1 U13102 ( .A(n17377), .ZN(n17373) );
  INV_X1 U13103 ( .A(n17509), .ZN(n17491) );
  INV_X1 U13104 ( .A(n17573), .ZN(n17564) );
  INV_X1 U13105 ( .A(n17787), .ZN(n17799) );
  INV_X1 U13106 ( .A(n17851), .ZN(n17748) );
  NOR2_X1 U13107 ( .A1(n16618), .A2(n18281), .ZN(n17883) );
  INV_X1 U13108 ( .A(n18172), .ZN(n18070) );
  AOI21_X1 U13109 ( .B1(n18042), .B2(n18090), .A(n18242), .ZN(n18150) );
  NAND3_X1 U13110 ( .A1(n15837), .A2(n15836), .A3(n15835), .ZN(n16498) );
  INV_X1 U13111 ( .A(n18242), .ZN(n18248) );
  INV_X1 U13112 ( .A(n18211), .ZN(n18244) );
  NAND2_X1 U13113 ( .A1(n18932), .A2(n18275), .ZN(n18372) );
  NOR2_X1 U13114 ( .A1(n18878), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n18897) );
  INV_X1 U13115 ( .A(n18463), .ZN(n18456) );
  NOR2_X1 U13116 ( .A1(n18775), .A2(n18930), .ZN(n18771) );
  INV_X1 U13117 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18807) );
  NAND2_X1 U13118 ( .A1(n12858), .A2(n12857), .ZN(n20949) );
  INV_X1 U13119 ( .A(n20948), .ZN(n20960) );
  INV_X1 U13120 ( .A(n20932), .ZN(n20948) );
  INV_X1 U13121 ( .A(n20145), .ZN(n20128) );
  INV_X1 U13122 ( .A(n20119), .ZN(n20104) );
  INV_X1 U13123 ( .A(n20140), .ZN(n20098) );
  INV_X1 U13124 ( .A(n20167), .ZN(n20187) );
  AND2_X1 U13125 ( .A1(n13088), .A2(n13087), .ZN(n13110) );
  OAI21_X1 U13126 ( .B1(n14291), .B2(n14211), .A(n14210), .ZN(n14611) );
  INV_X1 U13127 ( .A(n16138), .ZN(n16135) );
  NAND2_X1 U13128 ( .A1(n20063), .A2(n13037), .ZN(n16144) );
  NAND2_X1 U13129 ( .A1(n13256), .A2(n13243), .ZN(n16200) );
  INV_X1 U13130 ( .A(n16249), .ZN(n20230) );
  INV_X1 U13131 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20663) );
  OR2_X1 U13132 ( .A1(n20371), .A2(n20405), .ZN(n20327) );
  OR2_X1 U13133 ( .A1(n20371), .A2(n20445), .ZN(n20364) );
  OR2_X1 U13134 ( .A1(n20371), .A2(n20329), .ZN(n20399) );
  NAND2_X1 U13135 ( .A1(n20502), .A2(n20661), .ZN(n20466) );
  NAND2_X1 U13136 ( .A1(n20502), .A2(n20694), .ZN(n20501) );
  NAND2_X1 U13137 ( .A1(n20502), .A2(n20734), .ZN(n20529) );
  NAND2_X1 U13138 ( .A1(n20631), .A2(n20661), .ZN(n20591) );
  NAND2_X1 U13139 ( .A1(n20631), .A2(n20734), .ZN(n20640) );
  NAND2_X1 U13140 ( .A1(n20631), .A2(n20630), .ZN(n20693) );
  NAND2_X1 U13141 ( .A1(n20735), .A2(n20694), .ZN(n20792) );
  NAND2_X1 U13142 ( .A1(n20735), .A2(n20630), .ZN(n20865) );
  INV_X1 U13143 ( .A(n20938), .ZN(n20872) );
  OR2_X1 U13144 ( .A1(n10579), .A2(n10883), .ZN(n19174) );
  INV_X1 U13145 ( .A(n19183), .ZN(n19156) );
  INV_X1 U13146 ( .A(n19185), .ZN(n19154) );
  INV_X1 U13147 ( .A(n14998), .ZN(n15015) );
  INV_X1 U13148 ( .A(n14998), .ZN(n15004) );
  XNOR2_X1 U13149 ( .A(n12997), .B(n12996), .ZN(n19630) );
  NAND2_X1 U13150 ( .A1(n19239), .A2(n12710), .ZN(n19216) );
  AND2_X1 U13151 ( .A1(n12709), .A2(n19274), .ZN(n19239) );
  INV_X1 U13152 ( .A(n19241), .ZN(n19273) );
  NOR2_X1 U13153 ( .A1(n19313), .A2(n19345), .ZN(n19331) );
  INV_X1 U13154 ( .A(n19313), .ZN(n19347) );
  OR2_X1 U13155 ( .A1(n12618), .A2(n10598), .ZN(n19276) );
  INV_X1 U13156 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16331) );
  INV_X1 U13157 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16358) );
  OR2_X1 U13158 ( .A1(n15285), .A2(n15284), .ZN(n15579) );
  OR2_X1 U13159 ( .A1(n12477), .A2(n20046), .ZN(n19366) );
  OR2_X1 U13160 ( .A1(n19662), .A2(n19572), .ZN(n19454) );
  INV_X1 U13161 ( .A(n19507), .ZN(n19503) );
  INV_X1 U13162 ( .A(n19558), .ZN(n19571) );
  INV_X1 U13163 ( .A(n19590), .ZN(n19600) );
  INV_X1 U13164 ( .A(n19625), .ZN(n19621) );
  INV_X1 U13165 ( .A(n19650), .ZN(n19660) );
  OR2_X1 U13166 ( .A1(n19815), .A2(n19662), .ZN(n19684) );
  OR2_X1 U13167 ( .A1(n19815), .A2(n20007), .ZN(n19749) );
  INV_X1 U13168 ( .A(n19805), .ZN(n19813) );
  INV_X1 U13169 ( .A(n19851), .ZN(n19849) );
  INV_X1 U13170 ( .A(n19800), .ZN(n19905) );
  INV_X1 U13171 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16638) );
  INV_X1 U13172 ( .A(n17026), .ZN(n17017) );
  INV_X1 U13173 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17887) );
  INV_X1 U13174 ( .A(n16999), .ZN(n17027) );
  NOR3_X1 U13175 ( .A1(n16723), .A2(n17075), .A3(n17081), .ZN(n17080) );
  NOR2_X1 U13176 ( .A1(n17134), .A2(n17133), .ZN(n17147) );
  AND2_X1 U13177 ( .A1(n17314), .A2(n17404), .ZN(n17311) );
  AND4_X1 U13178 ( .A1(n18771), .A2(n18929), .A3(n9888), .A4(n15979), .ZN(
        n17314) );
  NOR2_X1 U13179 ( .A1(n15759), .A2(n15758), .ZN(n17444) );
  NAND2_X1 U13180 ( .A1(n17491), .A2(n9888), .ZN(n17489) );
  NAND2_X1 U13181 ( .A1(n17511), .A2(n17473), .ZN(n17509) );
  NAND2_X1 U13182 ( .A1(n17841), .A2(n18043), .ZN(n17751) );
  NAND2_X1 U13183 ( .A1(n16498), .A2(n17883), .ZN(n17851) );
  NAND2_X1 U13184 ( .A1(n18621), .A2(n18330), .ZN(n18373) );
  NAND2_X1 U13185 ( .A1(n16498), .A2(n18196), .ZN(n18172) );
  INV_X1 U13186 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18263) );
  INV_X1 U13187 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18932) );
  INV_X1 U13188 ( .A(n18874), .ZN(n21145) );
  INV_X1 U13189 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18804) );
  NAND2_X1 U13190 ( .A1(n12037), .A2(n12036), .ZN(P1_U2873) );
  INV_X1 U13191 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10259) );
  INV_X1 U13192 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15257) );
  INV_X1 U13193 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15196) );
  INV_X1 U13194 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15145) );
  INV_X1 U13195 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15125) );
  INV_X1 U13196 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10274) );
  INV_X1 U13197 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15105) );
  INV_X1 U13198 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n21100) );
  INV_X1 U13199 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12444) );
  OAI21_X1 U13200 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10242), .A(
        n10243), .ZN(n18991) );
  AOI21_X1 U13201 ( .B1(n15196), .B2(n10244), .A(n10242), .ZN(n19003) );
  AOI21_X1 U13202 ( .B1(n10265), .B2(n10239), .A(n9771), .ZN(n19028) );
  INV_X1 U13203 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19036) );
  INV_X1 U13204 ( .A(n10245), .ZN(n10246) );
  AOI21_X1 U13205 ( .B1(n19036), .B2(n10246), .A(n10264), .ZN(n19044) );
  AOI21_X1 U13206 ( .B1(n15257), .B2(n10262), .A(n10247), .ZN(n19064) );
  AOI21_X1 U13207 ( .B1(n19087), .B2(n10258), .A(n10248), .ZN(n19090) );
  AOI21_X1 U13208 ( .B1(n16331), .B2(n10256), .A(n10249), .ZN(n19110) );
  AOI21_X1 U13209 ( .B1(n15302), .B2(n10255), .A(n10250), .ZN(n19120) );
  AOI21_X1 U13210 ( .B1(n16358), .B2(n10254), .A(n9684), .ZN(n19147) );
  AOI21_X1 U13211 ( .B1(n13525), .B2(n10253), .A(n10251), .ZN(n13523) );
  INV_X1 U13212 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13721) );
  INV_X1 U13213 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U13214 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13721), .B1(n10252), 
        .B2(n19926), .ZN(n13720) );
  INV_X1 U13215 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U13216 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12277), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19926), .ZN(n13719) );
  NOR2_X1 U13217 ( .A1(n13720), .A2(n13719), .ZN(n13718) );
  OAI21_X1 U13218 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n10253), .ZN(n13740) );
  NAND2_X1 U13219 ( .A1(n13718), .A2(n13740), .ZN(n13521) );
  NOR2_X1 U13220 ( .A1(n13523), .A2(n13521), .ZN(n19161) );
  OAI21_X1 U13221 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10251), .A(
        n10254), .ZN(n19358) );
  NAND2_X1 U13222 ( .A1(n19161), .A2(n19358), .ZN(n19144) );
  NOR2_X1 U13223 ( .A1(n19147), .A2(n19144), .ZN(n19134) );
  OAI21_X1 U13224 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9684), .A(
        n10255), .ZN(n19135) );
  NAND2_X1 U13225 ( .A1(n19134), .A2(n19135), .ZN(n19119) );
  NOR2_X1 U13226 ( .A1(n19120), .A2(n19119), .ZN(n13552) );
  OAI21_X1 U13227 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10250), .A(
        n10256), .ZN(n16345) );
  NAND2_X1 U13228 ( .A1(n13552), .A2(n16345), .ZN(n19109) );
  NOR2_X1 U13229 ( .A1(n19110), .A2(n19109), .ZN(n19100) );
  OR2_X1 U13230 ( .A1(n10249), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10257) );
  NAND2_X1 U13231 ( .A1(n10258), .A2(n10257), .ZN(n19102) );
  NAND2_X1 U13232 ( .A1(n19100), .A2(n19102), .ZN(n19089) );
  NOR2_X1 U13233 ( .A1(n19090), .A2(n19089), .ZN(n19078) );
  NAND2_X1 U13234 ( .A1(n10260), .A2(n10259), .ZN(n10261) );
  NAND2_X1 U13235 ( .A1(n10262), .A2(n10261), .ZN(n19079) );
  NAND2_X1 U13236 ( .A1(n19078), .A2(n19079), .ZN(n19062) );
  NOR2_X1 U13237 ( .A1(n19064), .A2(n19062), .ZN(n19050) );
  NOR2_X1 U13238 ( .A1(n10247), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10263) );
  OR2_X1 U13239 ( .A1(n10245), .A2(n10263), .ZN(n19051) );
  NAND2_X1 U13240 ( .A1(n19050), .A2(n19051), .ZN(n19043) );
  NOR2_X1 U13241 ( .A1(n19044), .A2(n19043), .ZN(n14923) );
  OR2_X1 U13242 ( .A1(n10264), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10266) );
  NAND2_X1 U13243 ( .A1(n10266), .A2(n10265), .ZN(n15226) );
  NAND2_X1 U13244 ( .A1(n14923), .A2(n15226), .ZN(n19029) );
  NOR2_X1 U13245 ( .A1(n19028), .A2(n19029), .ZN(n19013) );
  OAI21_X1 U13246 ( .B1(n9771), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n10244), .ZN(n19014) );
  NAND2_X1 U13247 ( .A1(n19013), .A2(n19014), .ZN(n19001) );
  OAI21_X1 U13248 ( .B1(n19003), .B2(n19001), .A(n10267), .ZN(n18990) );
  AND2_X1 U13249 ( .A1(n18991), .A2(n18990), .ZN(n19000) );
  AOI21_X1 U13250 ( .B1(n10243), .B2(n10240), .A(n10268), .ZN(n18983) );
  OAI21_X1 U13251 ( .B1(n10268), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n10269), .ZN(n15156) );
  INV_X1 U13252 ( .A(n15156), .ZN(n14916) );
  NOR2_X1 U13253 ( .A1(n19162), .A2(n14915), .ZN(n14898) );
  AND2_X1 U13254 ( .A1(n10269), .A2(n15145), .ZN(n10270) );
  NOR2_X1 U13255 ( .A1(n9761), .A2(n10270), .ZN(n15143) );
  NOR2_X1 U13256 ( .A1(n14898), .A2(n15143), .ZN(n14897) );
  OR2_X1 U13257 ( .A1(n9761), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10272) );
  NAND2_X1 U13258 ( .A1(n10271), .A2(n10272), .ZN(n15136) );
  INV_X1 U13259 ( .A(n15136), .ZN(n16305) );
  INV_X1 U13260 ( .A(n10275), .ZN(n10273) );
  AOI21_X1 U13261 ( .B1(n15125), .B2(n10271), .A(n10273), .ZN(n15128) );
  NOR2_X1 U13262 ( .A1(n14874), .A2(n19162), .ZN(n16286) );
  NAND2_X1 U13263 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  NAND2_X1 U13264 ( .A1(n10277), .A2(n10276), .ZN(n15116) );
  INV_X1 U13265 ( .A(n15116), .ZN(n16288) );
  NOR2_X1 U13266 ( .A1(n19162), .A2(n16287), .ZN(n12599) );
  AND2_X1 U13267 ( .A1(n10277), .A2(n15105), .ZN(n10278) );
  NOR2_X1 U13268 ( .A1(n10280), .A2(n10278), .ZN(n15107) );
  NOR2_X1 U13269 ( .A1(n10280), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10281) );
  OR2_X1 U13270 ( .A1(n10279), .A2(n10281), .ZN(n12572) );
  INV_X1 U13271 ( .A(n12572), .ZN(n14862) );
  NOR2_X1 U13272 ( .A1(n10279), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10282) );
  OR2_X1 U13273 ( .A1(n10283), .A2(n10282), .ZN(n12548) );
  INV_X1 U13274 ( .A(n12548), .ZN(n14852) );
  XNOR2_X1 U13275 ( .A(n10283), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12516) );
  INV_X1 U13276 ( .A(n12516), .ZN(n10284) );
  NOR2_X1 U13277 ( .A1(n10285), .A2(n10284), .ZN(n16281) );
  INV_X1 U13278 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19695) );
  NAND4_X1 U13279 ( .A1(n20035), .A2(n19926), .A3(n19695), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19929) );
  AOI22_X1 U13280 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10289) );
  AND2_X2 U13281 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U13282 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10292) );
  AND2_X4 U13283 ( .A1(n15632), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13854) );
  AOI22_X1 U13284 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U13285 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10295) );
  AOI22_X1 U13286 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13875), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13287 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13288 ( .A1(n10591), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10351), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13289 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13290 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13291 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13292 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U13293 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U13294 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13295 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10313) );
  NAND4_X1 U13296 ( .A1(n10316), .A2(n10315), .A3(n10314), .A4(n10313), .ZN(
        n10317) );
  AOI22_X1 U13297 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13298 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9666), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10319) );
  NAND2_X1 U13299 ( .A1(n10320), .A2(n10319), .ZN(n10324) );
  AOI22_X1 U13300 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13301 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U13302 ( .A1(n10322), .A2(n10321), .ZN(n10323) );
  AOI22_X1 U13303 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10351), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13304 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13305 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9666), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U13306 ( .A1(n10591), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10327) );
  NAND4_X1 U13307 ( .A1(n10330), .A2(n10329), .A3(n10328), .A4(n10327), .ZN(
        n10331) );
  AOI22_X1 U13308 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9655), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13309 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13310 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10351), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13311 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9662), .B1(n9666), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10332) );
  NAND4_X1 U13312 ( .A1(n10335), .A2(n10334), .A3(n10333), .A4(n10332), .ZN(
        n10336) );
  AOI22_X1 U13313 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13314 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13315 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10339) );
  NAND4_X1 U13316 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  NAND2_X1 U13317 ( .A1(n10343), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10350) );
  AOI22_X1 U13318 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13319 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13320 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10344) );
  NAND4_X1 U13321 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10348) );
  NAND2_X1 U13322 ( .A1(n10348), .A2(n10383), .ZN(n10349) );
  AOI22_X1 U13323 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13875), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U13324 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9666), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13325 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13326 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10352) );
  NAND4_X1 U13327 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        n10356) );
  NAND2_X1 U13328 ( .A1(n10356), .A2(n10383), .ZN(n10364) );
  AOI22_X1 U13329 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13330 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13875), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13331 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10359) );
  NAND4_X1 U13332 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10362) );
  NAND2_X1 U13333 ( .A1(n10362), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10363) );
  AND2_X2 U13334 ( .A1(n10364), .A2(n10363), .ZN(n10393) );
  INV_X1 U13335 ( .A(n12242), .ZN(n10396) );
  NAND2_X1 U13336 ( .A1(n10405), .A2(n10396), .ZN(n10410) );
  INV_X1 U13337 ( .A(n10410), .ZN(n10374) );
  AOI22_X1 U13338 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13339 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13340 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U13341 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10373) );
  AOI21_X2 U13342 ( .B1(n10351), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n10369), .ZN(n10372) );
  AOI22_X1 U13343 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13875), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13344 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9666), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10370) );
  NAND2_X1 U13345 ( .A1(n10374), .A2(n19378), .ZN(n10580) );
  AND2_X1 U13346 ( .A1(n10408), .A2(n10401), .ZN(n10376) );
  NAND3_X2 U13347 ( .A1(n10378), .A2(n10377), .A3(n10376), .ZN(n12704) );
  NAND2_X1 U13348 ( .A1(n10580), .A2(n12704), .ZN(n10577) );
  AOI22_X1 U13349 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n9666), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13350 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9655), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13351 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13352 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10379) );
  NAND4_X1 U13353 ( .A1(n10382), .A2(n10381), .A3(n10380), .A4(n10379), .ZN(
        n10384) );
  AOI22_X1 U13354 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9666), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13355 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13356 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13357 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10586), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10385) );
  NAND4_X1 U13358 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10389) );
  NAND2_X2 U13359 ( .A1(n10391), .A2(n10390), .ZN(n10583) );
  NAND2_X2 U13360 ( .A1(n10583), .A2(n19378), .ZN(n12221) );
  NAND2_X1 U13361 ( .A1(n10396), .A2(n12215), .ZN(n10399) );
  INV_X1 U13362 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16374) );
  AOI22_X1 U13363 ( .A1(n12440), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10404) );
  AND2_X1 U13364 ( .A1(n10583), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U13365 ( .A1(n12441), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10403) );
  OAI211_X1 U13366 ( .C1(n10473), .C2(n16374), .A(n10404), .B(n10403), .ZN(
        n13196) );
  INV_X1 U13367 ( .A(n13196), .ZN(n10494) );
  NAND2_X1 U13368 ( .A1(n10405), .A2(n10378), .ZN(n12213) );
  NAND2_X1 U13369 ( .A1(n12213), .A2(n10409), .ZN(n10411) );
  NAND2_X1 U13370 ( .A1(n10411), .A2(n16418), .ZN(n12457) );
  NAND2_X1 U13371 ( .A1(n10414), .A2(n12704), .ZN(n12465) );
  AND2_X1 U13372 ( .A1(n10417), .A2(n10406), .ZN(n10433) );
  NAND2_X1 U13373 ( .A1(n12243), .A2(n10231), .ZN(n12241) );
  NAND2_X1 U13374 ( .A1(n10417), .A2(n12467), .ZN(n12246) );
  NAND3_X1 U13375 ( .A1(n12241), .A2(n12246), .A3(n19422), .ZN(n12463) );
  NAND2_X1 U13376 ( .A1(n12463), .A2(n10397), .ZN(n10420) );
  NAND2_X1 U13377 ( .A1(n10418), .A2(n10398), .ZN(n10419) );
  INV_X1 U13378 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10428) );
  NAND2_X1 U13379 ( .A1(n9920), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U13380 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10426) );
  OAI211_X1 U13381 ( .C1(n10511), .C2(n10428), .A(n10427), .B(n10426), .ZN(
        n10429) );
  INV_X1 U13382 ( .A(n10429), .ZN(n10430) );
  XNOR2_X1 U13383 ( .A(n10453), .B(n10452), .ZN(n12056) );
  NAND2_X1 U13384 ( .A1(n10432), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10444) );
  INV_X1 U13385 ( .A(n10433), .ZN(n10434) );
  NAND2_X1 U13386 ( .A1(n10435), .A2(n10434), .ZN(n12475) );
  NAND2_X1 U13387 ( .A1(n12475), .A2(n10436), .ZN(n10442) );
  INV_X1 U13388 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10440) );
  NAND2_X1 U13389 ( .A1(n9920), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10439) );
  AND2_X1 U13390 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10437) );
  NOR2_X1 U13391 ( .A1(n16419), .A2(n10437), .ZN(n10438) );
  OAI211_X1 U13392 ( .C1(n10511), .C2(n10440), .A(n10439), .B(n10438), .ZN(
        n10441) );
  INV_X1 U13393 ( .A(n10445), .ZN(n10447) );
  AND2_X1 U13394 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10446) );
  INV_X1 U13395 ( .A(n13054), .ZN(n10449) );
  AOI22_X1 U13396 ( .A1(n10449), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16419), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10450) );
  NAND2_X1 U13397 ( .A1(n10451), .A2(n10450), .ZN(n12040) );
  INV_X1 U13398 ( .A(n10452), .ZN(n10454) );
  NAND2_X1 U13399 ( .A1(n10454), .A2(n10453), .ZN(n10455) );
  INV_X1 U13400 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21118) );
  INV_X1 U13401 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U13402 ( .A1(n9920), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10457) );
  NAND2_X1 U13403 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10456) );
  OAI211_X1 U13404 ( .C1(n10511), .C2(n10458), .A(n10457), .B(n10456), .ZN(
        n10459) );
  INV_X1 U13405 ( .A(n10459), .ZN(n10460) );
  OAI21_X2 U13406 ( .B1(n10473), .B2(n21118), .A(n10460), .ZN(n12042) );
  AOI21_X1 U13407 ( .B1(n19926), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U13408 ( .A1(n12042), .A2(n12041), .ZN(n10464) );
  NAND2_X1 U13409 ( .A1(n12044), .A2(n10464), .ZN(n10468) );
  INV_X1 U13410 ( .A(n12042), .ZN(n10466) );
  INV_X1 U13411 ( .A(n12041), .ZN(n10465) );
  NAND2_X1 U13412 ( .A1(n10466), .A2(n10465), .ZN(n10467) );
  INV_X1 U13413 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13613) );
  INV_X1 U13414 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10658) );
  NAND2_X1 U13415 ( .A1(n9920), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U13416 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10469) );
  OAI211_X1 U13417 ( .C1(n10511), .C2(n10658), .A(n10470), .B(n10469), .ZN(
        n10471) );
  INV_X1 U13418 ( .A(n10471), .ZN(n10472) );
  INV_X1 U13419 ( .A(n10478), .ZN(n10475) );
  AND2_X1 U13420 ( .A1(n16419), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10474) );
  NAND2_X1 U13421 ( .A1(n10475), .A2(n10476), .ZN(n10480) );
  INV_X1 U13422 ( .A(n10476), .ZN(n10477) );
  NAND2_X1 U13423 ( .A1(n10478), .A2(n10477), .ZN(n10479) );
  INV_X1 U13424 ( .A(n12038), .ZN(n10482) );
  INV_X1 U13425 ( .A(n10480), .ZN(n10481) );
  INV_X1 U13426 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10674) );
  INV_X1 U13427 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13656) );
  OR2_X1 U13428 ( .A1(n10473), .A2(n13656), .ZN(n10485) );
  AOI22_X1 U13429 ( .A1(n12440), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10484) );
  OAI211_X1 U13430 ( .C1(n10511), .C2(n10674), .A(n10485), .B(n10484), .ZN(
        n13003) );
  INV_X1 U13431 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13662) );
  OR2_X1 U13432 ( .A1(n10473), .A2(n13662), .ZN(n10490) );
  INV_X1 U13433 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13659) );
  NAND2_X1 U13434 ( .A1(n12440), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10487) );
  NAND2_X1 U13435 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10486) );
  OAI211_X1 U13436 ( .C1(n10511), .C2(n13659), .A(n10487), .B(n10486), .ZN(
        n10488) );
  INV_X1 U13437 ( .A(n10488), .ZN(n10489) );
  INV_X1 U13438 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n10493) );
  INV_X1 U13439 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15604) );
  OR2_X1 U13440 ( .A1(n10473), .A2(n15604), .ZN(n10492) );
  AOI22_X1 U13441 ( .A1(n12440), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10491) );
  OAI211_X1 U13442 ( .C1(n10511), .C2(n10493), .A(n10492), .B(n10491), .ZN(
        n13118) );
  INV_X1 U13443 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U13444 ( .A1(n12440), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10496) );
  NAND2_X1 U13445 ( .A1(n12441), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10495) );
  OAI211_X1 U13446 ( .C1(n10473), .C2(n12481), .A(n10496), .B(n10495), .ZN(
        n13202) );
  INV_X1 U13447 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15591) );
  OR2_X1 U13448 ( .A1(n10473), .A2(n15591), .ZN(n10501) );
  INV_X1 U13449 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n10748) );
  NAND2_X1 U13450 ( .A1(n12440), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10498) );
  NAND2_X1 U13451 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10497) );
  OAI211_X1 U13452 ( .C1(n10511), .C2(n10748), .A(n10498), .B(n10497), .ZN(
        n10499) );
  INV_X1 U13453 ( .A(n10499), .ZN(n10500) );
  NAND2_X1 U13454 ( .A1(n10501), .A2(n10500), .ZN(n13012) );
  INV_X1 U13455 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19961) );
  INV_X1 U13456 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15546) );
  OR2_X1 U13457 ( .A1(n10473), .A2(n15546), .ZN(n10503) );
  AOI22_X1 U13458 ( .A1(n12440), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10502) );
  OAI211_X1 U13459 ( .C1(n10511), .C2(n19961), .A(n10503), .B(n10502), .ZN(
        n13124) );
  INV_X1 U13460 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n15278) );
  NAND2_X1 U13461 ( .A1(n12440), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10505) );
  NAND2_X1 U13462 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10504) );
  OAI211_X1 U13463 ( .C1(n10511), .C2(n15278), .A(n10505), .B(n10504), .ZN(
        n10506) );
  AOI21_X1 U13464 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10506), .ZN(n13211) );
  INV_X1 U13465 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19964) );
  INV_X1 U13466 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15521) );
  OR2_X1 U13467 ( .A1(n10473), .A2(n15521), .ZN(n10508) );
  AOI22_X1 U13468 ( .A1(n12440), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10507) );
  OAI211_X1 U13469 ( .C1(n10511), .C2(n19964), .A(n10508), .B(n10507), .ZN(
        n13377) );
  INV_X1 U13470 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19966) );
  NAND2_X1 U13471 ( .A1(n12440), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10510) );
  NAND2_X1 U13472 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10509) );
  OAI211_X1 U13473 ( .C1(n10511), .C2(n19966), .A(n10510), .B(n10509), .ZN(
        n10512) );
  AOI21_X1 U13474 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10512), .ZN(n13445) );
  INV_X1 U13475 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U13476 ( .A1(n12440), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10514) );
  NAND2_X1 U13477 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10513) );
  OAI211_X1 U13478 ( .C1(n10557), .C2(n10814), .A(n10514), .B(n10513), .ZN(
        n10515) );
  AOI21_X1 U13479 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10515), .ZN(n13480) );
  INV_X1 U13480 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n21116) );
  NAND2_X1 U13481 ( .A1(n12440), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10517) );
  NAND2_X1 U13482 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10516) );
  OAI211_X1 U13483 ( .C1(n10557), .C2(n21116), .A(n10517), .B(n10516), .ZN(
        n10518) );
  AOI21_X1 U13484 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10518), .ZN(n13485) );
  INV_X1 U13485 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19970) );
  INV_X1 U13486 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15478) );
  OR2_X1 U13487 ( .A1(n10473), .A2(n15478), .ZN(n10520) );
  AOI22_X1 U13488 ( .A1(n12440), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10519) );
  OAI211_X1 U13489 ( .C1(n10557), .C2(n19970), .A(n10520), .B(n10519), .ZN(
        n13643) );
  NAND2_X1 U13490 ( .A1(n13644), .A2(n13643), .ZN(n15020) );
  INV_X1 U13491 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19972) );
  NAND2_X1 U13492 ( .A1(n12440), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10522) );
  NAND2_X1 U13493 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10521) );
  OAI211_X1 U13494 ( .C1(n10557), .C2(n19972), .A(n10522), .B(n10521), .ZN(
        n10523) );
  AOI21_X1 U13495 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10523), .ZN(n15019) );
  INV_X1 U13496 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n10834) );
  NAND2_X1 U13497 ( .A1(n12440), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10525) );
  NAND2_X1 U13498 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10524) );
  OAI211_X1 U13499 ( .C1(n10557), .C2(n10834), .A(n10525), .B(n10524), .ZN(
        n10526) );
  AOI21_X1 U13500 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10526), .ZN(n15006) );
  INV_X1 U13501 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19975) );
  INV_X1 U13502 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15432) );
  OR2_X1 U13503 ( .A1(n10473), .A2(n15432), .ZN(n10528) );
  AOI22_X1 U13504 ( .A1(n12440), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10527) );
  OAI211_X1 U13505 ( .C1(n10557), .C2(n19975), .A(n10528), .B(n10527), .ZN(
        n15001) );
  INV_X1 U13506 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15188) );
  INV_X1 U13507 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15425) );
  OR2_X1 U13508 ( .A1(n10473), .A2(n15425), .ZN(n10530) );
  AOI22_X1 U13509 ( .A1(n12440), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10529) );
  OAI211_X1 U13510 ( .C1(n10557), .C2(n15188), .A(n10530), .B(n10529), .ZN(
        n14993) );
  INV_X1 U13511 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U13512 ( .A1(n12440), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10532) );
  NAND2_X1 U13513 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10531) );
  OAI211_X1 U13514 ( .C1(n10557), .C2(n10533), .A(n10532), .B(n10531), .ZN(
        n10534) );
  AOI21_X1 U13515 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10534), .ZN(n14985) );
  INV_X1 U13516 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19979) );
  NAND2_X1 U13517 ( .A1(n12440), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10536) );
  NAND2_X1 U13518 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10535) );
  OAI211_X1 U13519 ( .C1(n10557), .C2(n19979), .A(n10536), .B(n10535), .ZN(
        n10537) );
  AOI21_X1 U13520 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10537), .ZN(n14903) );
  INV_X1 U13521 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19981) );
  INV_X1 U13522 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12491) );
  OR2_X1 U13523 ( .A1(n10473), .A2(n12491), .ZN(n10539) );
  AOI22_X1 U13524 ( .A1(n12440), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10538) );
  OAI211_X1 U13525 ( .C1(n10557), .C2(n19981), .A(n10539), .B(n10538), .ZN(
        n14887) );
  INV_X1 U13526 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19983) );
  INV_X1 U13527 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12399) );
  OR2_X1 U13528 ( .A1(n10473), .A2(n12399), .ZN(n10541) );
  AOI22_X1 U13529 ( .A1(n12440), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10540) );
  OAI211_X1 U13530 ( .C1(n10557), .C2(n19983), .A(n10541), .B(n10540), .ZN(
        n14968) );
  INV_X1 U13531 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19985) );
  NAND2_X1 U13532 ( .A1(n12440), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10543) );
  NAND2_X1 U13533 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10542) );
  OAI211_X1 U13534 ( .C1(n10557), .C2(n19985), .A(n10543), .B(n10542), .ZN(
        n10544) );
  AOI21_X1 U13535 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10544), .ZN(n14880) );
  INV_X1 U13536 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n10850) );
  NAND2_X1 U13537 ( .A1(n12440), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10546) );
  NAND2_X1 U13538 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10545) );
  OAI211_X1 U13539 ( .C1(n10557), .C2(n10850), .A(n10546), .B(n10545), .ZN(
        n10547) );
  AOI21_X1 U13540 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10547), .ZN(n14950) );
  INV_X1 U13541 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19989) );
  NAND2_X1 U13542 ( .A1(n12440), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10549) );
  NAND2_X1 U13543 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10548) );
  OAI211_X1 U13544 ( .C1(n10557), .C2(n19989), .A(n10549), .B(n10548), .ZN(
        n10550) );
  AOI21_X1 U13545 ( .B1(n9654), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10550), .ZN(n12602) );
  INV_X1 U13546 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19990) );
  INV_X1 U13547 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15329) );
  OR2_X1 U13548 ( .A1(n10473), .A2(n15329), .ZN(n10552) );
  AOI22_X1 U13549 ( .A1(n12440), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10551) );
  OAI211_X1 U13550 ( .C1(n10557), .C2(n19990), .A(n10552), .B(n10551), .ZN(
        n12567) );
  INV_X1 U13551 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19992) );
  INV_X1 U13552 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12539) );
  OR2_X1 U13553 ( .A1(n10473), .A2(n12539), .ZN(n10554) );
  AOI22_X1 U13554 ( .A1(n12440), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10553) );
  OAI211_X1 U13555 ( .C1(n10557), .C2(n19992), .A(n10554), .B(n10553), .ZN(
        n12544) );
  INV_X1 U13556 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n10859) );
  INV_X1 U13557 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12506) );
  OR2_X1 U13558 ( .A1(n10473), .A2(n12506), .ZN(n10556) );
  AOI22_X1 U13559 ( .A1(n12440), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10555) );
  OAI211_X1 U13560 ( .C1(n10557), .C2(n10859), .A(n10556), .B(n10555), .ZN(
        n12439) );
  NAND2_X1 U13561 ( .A1(n20042), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12206) );
  NAND2_X1 U13562 ( .A1(n12214), .A2(n10570), .ZN(n10559) );
  NAND2_X1 U13563 ( .A1(n20033), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10558) );
  NOR2_X1 U13564 ( .A1(n9640), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10560) );
  MUX2_X1 U13565 ( .A(n10561), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n10383), .Z(n10565) );
  NAND2_X1 U13566 ( .A1(n10561), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10562) );
  NOR2_X1 U13567 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15978), .ZN(
        n10564) );
  XNOR2_X1 U13568 ( .A(n10566), .B(n10565), .ZN(n10864) );
  XNOR2_X1 U13569 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10567) );
  XNOR2_X1 U13570 ( .A(n10568), .B(n10567), .ZN(n12225) );
  INV_X1 U13571 ( .A(n12225), .ZN(n10569) );
  NAND2_X1 U13572 ( .A1(n12229), .A2(n10569), .ZN(n12257) );
  XNOR2_X1 U13573 ( .A(n12214), .B(n10570), .ZN(n12216) );
  OR2_X1 U13574 ( .A1(n12257), .A2(n12216), .ZN(n10576) );
  NAND2_X1 U13575 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15978), .ZN(
        n10571) );
  NAND2_X1 U13576 ( .A1(n10572), .A2(n10571), .ZN(n10574) );
  NAND2_X1 U13577 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16397), .ZN(
        n10573) );
  INV_X1 U13578 ( .A(n12235), .ZN(n10575) );
  NAND2_X1 U13579 ( .A1(n16424), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19932) );
  AND2_X1 U13580 ( .A1(n12613), .A2(n10578), .ZN(n18952) );
  AND2_X1 U13581 ( .A1(n18952), .A2(n10421), .ZN(n10882) );
  INV_X1 U13582 ( .A(n10882), .ZN(n10579) );
  NAND2_X1 U13583 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19924) );
  NAND2_X1 U13584 ( .A1(n19924), .A2(n19695), .ZN(n10883) );
  INV_X1 U13585 ( .A(n10580), .ZN(n10581) );
  NAND2_X1 U13586 ( .A1(n12613), .A2(n10581), .ZN(n12618) );
  NOR2_X1 U13587 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n18955) );
  AOI211_X1 U13588 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n18955), .ZN(n19938) );
  INV_X1 U13589 ( .A(n19938), .ZN(n10582) );
  INV_X1 U13590 ( .A(n19924), .ZN(n19943) );
  NOR2_X1 U13591 ( .A1(n10582), .A2(n19943), .ZN(n16385) );
  NAND2_X1 U13592 ( .A1(n19695), .A2(n16385), .ZN(n16417) );
  AND2_X2 U13593 ( .A1(n9662), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10693) );
  AOI22_X1 U13594 ( .A1(n10694), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10590) );
  AOI22_X1 U13595 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10675), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13596 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10588) );
  AND2_X2 U13597 ( .A1(n9652), .A2(n10383), .ZN(n10623) );
  AND2_X2 U13598 ( .A1(n13971), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10638) );
  AOI22_X1 U13599 ( .A1(n10623), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10587) );
  NAND4_X1 U13600 ( .A1(n10590), .A2(n10589), .A3(n10588), .A4(n10587), .ZN(
        n10597) );
  AND2_X1 U13601 ( .A1(n9641), .A2(n10383), .ZN(n10643) );
  AOI22_X1 U13602 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13834), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13603 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10594) );
  AND2_X2 U13604 ( .A1(n13854), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13835) );
  AOI22_X1 U13605 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10593) );
  AND2_X2 U13606 ( .A1(n13972), .A2(n10383), .ZN(n13836) );
  CLKBUF_X3 U13607 ( .A(n10351), .Z(n13964) );
  AOI22_X1 U13608 ( .A1(n13836), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10592) );
  NAND4_X1 U13609 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n10596) );
  AOI22_X1 U13610 ( .A1(n10162), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n10825), 
        .B2(n12159), .ZN(n10600) );
  AOI22_X1 U13611 ( .A1(n10857), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12449), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U13612 ( .A1(n10600), .A2(n10599), .ZN(n13657) );
  AOI22_X1 U13613 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13614 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13615 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13616 ( .A1(n13836), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10603) );
  NAND4_X1 U13617 ( .A1(n10606), .A2(n10605), .A3(n10604), .A4(n10603), .ZN(
        n10612) );
  AOI22_X1 U13618 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13834), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13619 ( .A1(n10694), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13620 ( .A1(n13838), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13621 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13839), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10607) );
  NAND4_X1 U13622 ( .A1(n10610), .A2(n10609), .A3(n10608), .A4(n10607), .ZN(
        n10611) );
  NOR2_X1 U13623 ( .A1(n10612), .A2(n10611), .ZN(n12881) );
  INV_X1 U13624 ( .A(n12881), .ZN(n10613) );
  MUX2_X1 U13625 ( .A(n19422), .B(n20042), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10614) );
  INV_X1 U13626 ( .A(n10417), .ZN(n12710) );
  NAND2_X1 U13627 ( .A1(n12710), .A2(n10619), .ZN(n10650) );
  AND2_X1 U13628 ( .A1(n10614), .A2(n10650), .ZN(n10615) );
  AOI21_X1 U13629 ( .B1(n10598), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10618) );
  NAND2_X1 U13630 ( .A1(n12711), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10617) );
  INV_X2 U13631 ( .A(n10235), .ZN(n10857) );
  AOI22_X1 U13632 ( .A1(n10857), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10619), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10620) );
  INV_X1 U13633 ( .A(n10636), .ZN(n10621) );
  NAND2_X1 U13634 ( .A1(n10417), .A2(n19422), .ZN(n10622) );
  MUX2_X1 U13635 ( .A(n10622), .B(n20033), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10635) );
  AOI22_X1 U13636 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10694), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13637 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13638 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13639 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10624) );
  NAND4_X1 U13640 ( .A1(n10627), .A2(n10626), .A3(n10625), .A4(n10624), .ZN(
        n10633) );
  AOI22_X1 U13641 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n13834), .ZN(n10631) );
  AOI22_X1 U13642 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10630) );
  AOI22_X1 U13643 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U13644 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10628) );
  NAND4_X1 U13645 ( .A1(n10631), .A2(n10630), .A3(n10629), .A4(n10628), .ZN(
        n10632) );
  NAND2_X1 U13646 ( .A1(n10825), .A2(n12115), .ZN(n10634) );
  AND2_X1 U13647 ( .A1(n10635), .A2(n10634), .ZN(n13078) );
  NAND2_X1 U13648 ( .A1(n13076), .A2(n13078), .ZN(n13077) );
  AOI22_X1 U13649 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10694), .B1(
        n10675), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U13650 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10693), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U13651 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10640) );
  AOI22_X1 U13652 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10639) );
  NAND4_X1 U13653 ( .A1(n10642), .A2(n10641), .A3(n10640), .A4(n10639), .ZN(
        n10649) );
  AOI22_X1 U13654 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U13655 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U13656 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13836), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U13657 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n13834), .ZN(n10644) );
  NAND4_X1 U13658 ( .A1(n10647), .A2(n10646), .A3(n10645), .A4(n10644), .ZN(
        n10648) );
  NAND2_X1 U13659 ( .A1(n10825), .A2(n12118), .ZN(n10651) );
  OAI211_X1 U13660 ( .C1(n20023), .C2(n19632), .A(n10651), .B(n10650), .ZN(
        n10652) );
  AND3_X1 U13661 ( .A1(n13077), .A2(n9697), .A3(n10652), .ZN(n10653) );
  OR2_X1 U13662 ( .A1(n12452), .A2(n10458), .ZN(n10655) );
  AOI22_X1 U13663 ( .A1(n10857), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12449), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10654) );
  NAND2_X1 U13664 ( .A1(n10655), .A2(n10654), .ZN(n13071) );
  INV_X2 U13665 ( .A(n10722), .ZN(n12449) );
  AOI22_X1 U13666 ( .A1(n12449), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10657) );
  OAI21_X1 U13667 ( .B1(n12452), .B2(n10658), .A(n10657), .ZN(n10673) );
  AOI22_X1 U13668 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10643), .B1(
        n13835), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13669 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n13834), .ZN(n10661) );
  AOI22_X1 U13670 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10638), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13671 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13836), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10659) );
  NAND4_X1 U13672 ( .A1(n10662), .A2(n10661), .A3(n10660), .A4(n10659), .ZN(
        n10669) );
  AOI22_X1 U13673 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10694), .B1(
        n10675), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13674 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10693), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13675 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13676 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10623), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10664) );
  NAND4_X1 U13677 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10668) );
  NOR2_X1 U13678 ( .A1(n10669), .A2(n10668), .ZN(n10865) );
  INV_X1 U13679 ( .A(n10865), .ZN(n12083) );
  NAND2_X1 U13680 ( .A1(n10825), .A2(n12083), .ZN(n10671) );
  NAND2_X1 U13681 ( .A1(n10857), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10670) );
  NAND2_X1 U13682 ( .A1(n10671), .A2(n10670), .ZN(n10672) );
  OR2_X1 U13683 ( .A1(n12452), .A2(n10674), .ZN(n10692) );
  AOI22_X1 U13684 ( .A1(n10857), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12449), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13685 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10694), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13686 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13687 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13688 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10676) );
  NAND4_X1 U13689 ( .A1(n10679), .A2(n10678), .A3(n10677), .A4(n10676), .ZN(
        n10689) );
  AOI22_X1 U13690 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n13834), .ZN(n10687) );
  AOI22_X1 U13691 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13692 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10685) );
  INV_X1 U13693 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21126) );
  INV_X1 U13694 ( .A(n10680), .ZN(n10682) );
  INV_X1 U13695 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10681) );
  OAI22_X1 U13696 ( .A1(n21126), .A2(n12253), .B1(n10682), .B2(n10681), .ZN(
        n10683) );
  INV_X1 U13697 ( .A(n10683), .ZN(n10684) );
  NAND4_X1 U13698 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n10688) );
  NAND2_X1 U13699 ( .A1(n10825), .A2(n10867), .ZN(n10690) );
  INV_X1 U13700 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10698) );
  INV_X1 U13701 ( .A(n10693), .ZN(n10697) );
  INV_X1 U13702 ( .A(n10694), .ZN(n10696) );
  INV_X1 U13703 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10695) );
  OAI22_X1 U13704 ( .A1(n10698), .A2(n10697), .B1(n10696), .B2(n10695), .ZN(
        n10699) );
  INV_X1 U13705 ( .A(n10699), .ZN(n10703) );
  AOI22_X1 U13706 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13707 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13708 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10700) );
  NAND4_X1 U13709 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n10709) );
  AOI22_X1 U13710 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n13834), .ZN(n10707) );
  AOI22_X1 U13711 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n13839), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13712 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13713 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10704) );
  NAND4_X1 U13714 ( .A1(n10707), .A2(n10706), .A3(n10705), .A4(n10704), .ZN(
        n10708) );
  AOI22_X1 U13715 ( .A1(n13657), .A2(n13658), .B1(n10825), .B2(n12181), .ZN(
        n15607) );
  INV_X1 U13716 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19333) );
  OAI222_X1 U13717 ( .A1(n15604), .A2(n10722), .B1(n10235), .B2(n19333), .C1(
        n12452), .C2(n10493), .ZN(n15606) );
  INV_X1 U13718 ( .A(n15606), .ZN(n10721) );
  AOI22_X1 U13719 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10694), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13720 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13721 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13722 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10710) );
  NAND4_X1 U13723 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n10719) );
  AOI22_X1 U13724 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n13834), .ZN(n10717) );
  AOI22_X1 U13725 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n13839), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13726 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13727 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10714) );
  NAND4_X1 U13728 ( .A1(n10717), .A2(n10716), .A3(n10715), .A4(n10714), .ZN(
        n10718) );
  INV_X1 U13729 ( .A(n10825), .ZN(n10720) );
  INV_X1 U13730 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19330) );
  INV_X1 U13731 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20984) );
  OAI222_X1 U13732 ( .A1(n16374), .A2(n10722), .B1(n10235), .B2(n19330), .C1(
        n12452), .C2(n20984), .ZN(n16369) );
  INV_X1 U13733 ( .A(n13556), .ZN(n10735) );
  INV_X1 U13734 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13561) );
  AOI22_X1 U13735 ( .A1(n10857), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12449), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13736 ( .A1(n10694), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13737 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10675), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13738 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13739 ( .A1(n10623), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10723) );
  NAND4_X1 U13740 ( .A1(n10726), .A2(n10725), .A3(n10724), .A4(n10723), .ZN(
        n10732) );
  AOI22_X1 U13741 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13834), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13742 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13743 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13744 ( .A1(n13836), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10727) );
  NAND4_X1 U13745 ( .A1(n10730), .A2(n10729), .A3(n10728), .A4(n10727), .ZN(
        n10731) );
  NAND2_X1 U13746 ( .A1(n10825), .A2(n13201), .ZN(n10733) );
  OAI211_X1 U13747 ( .C1(n12452), .C2(n13561), .A(n10734), .B(n10733), .ZN(
        n13555) );
  NAND2_X1 U13748 ( .A1(n10735), .A2(n13555), .ZN(n13557) );
  AOI22_X1 U13749 ( .A1(n10857), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12449), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13750 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10693), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U13751 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U13752 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U13753 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10736) );
  NAND4_X1 U13754 ( .A1(n10739), .A2(n10738), .A3(n10737), .A4(n10736), .ZN(
        n10745) );
  AOI22_X1 U13755 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n13834), .ZN(n10743) );
  AOI22_X1 U13756 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13757 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13758 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10740) );
  NAND4_X1 U13759 ( .A1(n10743), .A2(n10742), .A3(n10741), .A4(n10740), .ZN(
        n10744) );
  NAND2_X1 U13760 ( .A1(n10825), .A2(n13011), .ZN(n10746) );
  OAI211_X1 U13761 ( .C1(n12452), .C2(n10748), .A(n10747), .B(n10746), .ZN(
        n10749) );
  INV_X1 U13762 ( .A(n10749), .ZN(n15581) );
  AOI22_X1 U13763 ( .A1(n10857), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13764 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10693), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U13765 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10675), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U13766 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U13767 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10623), .B1(
        n13836), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10750) );
  NAND4_X1 U13768 ( .A1(n10753), .A2(n10752), .A3(n10751), .A4(n10750), .ZN(
        n10759) );
  AOI22_X1 U13769 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13770 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13771 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U13772 ( .A1(n10680), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n13834), .ZN(n10754) );
  NAND4_X1 U13773 ( .A1(n10757), .A2(n10756), .A3(n10755), .A4(n10754), .ZN(
        n10758) );
  NAND2_X1 U13774 ( .A1(n10825), .A2(n13130), .ZN(n10760) );
  OAI211_X1 U13775 ( .C1(n12452), .C2(n19961), .A(n10761), .B(n10760), .ZN(
        n10762) );
  INV_X1 U13776 ( .A(n10762), .ZN(n15566) );
  AOI22_X1 U13777 ( .A1(n10857), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13778 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10693), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13779 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U13780 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13781 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10763) );
  NAND4_X1 U13782 ( .A1(n10766), .A2(n10765), .A3(n10764), .A4(n10763), .ZN(
        n10772) );
  AOI22_X1 U13783 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n13834), .ZN(n10770) );
  AOI22_X1 U13784 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13785 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U13786 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10767) );
  NAND4_X1 U13787 ( .A1(n10770), .A2(n10769), .A3(n10768), .A4(n10767), .ZN(
        n10771) );
  NAND2_X1 U13788 ( .A1(n10825), .A2(n13210), .ZN(n10773) );
  OAI211_X1 U13789 ( .C1(n12452), .C2(n15278), .A(n10774), .B(n10773), .ZN(
        n10775) );
  INV_X1 U13790 ( .A(n10775), .ZN(n15551) );
  AOI22_X1 U13791 ( .A1(n10857), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13792 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10779) );
  AOI22_X1 U13793 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10693), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13794 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13795 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10623), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10776) );
  NAND4_X1 U13796 ( .A1(n10779), .A2(n10778), .A3(n10777), .A4(n10776), .ZN(
        n10785) );
  AOI22_X1 U13797 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13811), .B1(
        n13839), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13798 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n13834), .ZN(n10782) );
  AOI22_X1 U13799 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10638), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10781) );
  AOI22_X1 U13800 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13836), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10780) );
  NAND4_X1 U13801 ( .A1(n10783), .A2(n10782), .A3(n10781), .A4(n10780), .ZN(
        n10784) );
  NAND2_X1 U13802 ( .A1(n10825), .A2(n13380), .ZN(n10786) );
  OAI211_X1 U13803 ( .C1(n12452), .C2(n19964), .A(n10787), .B(n10786), .ZN(
        n15535) );
  AND2_X2 U13804 ( .A1(n15550), .A2(n15535), .ZN(n15533) );
  AOI22_X1 U13805 ( .A1(n10857), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U13806 ( .A1(n10694), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13807 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10675), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13808 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13809 ( .A1(n10623), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10788) );
  NAND4_X1 U13810 ( .A1(n10791), .A2(n10790), .A3(n10789), .A4(n10788), .ZN(
        n10797) );
  AOI22_X1 U13811 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13834), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13812 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13813 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13814 ( .A1(n13836), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10792) );
  NAND4_X1 U13815 ( .A1(n10795), .A2(n10794), .A3(n10793), .A4(n10792), .ZN(
        n10796) );
  NAND2_X1 U13816 ( .A1(n10825), .A2(n13444), .ZN(n10798) );
  OAI211_X1 U13817 ( .C1(n12452), .C2(n19966), .A(n10799), .B(n10798), .ZN(
        n15519) );
  AND2_X2 U13818 ( .A1(n15533), .A2(n15519), .ZN(n15509) );
  AOI22_X1 U13819 ( .A1(n10857), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13820 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10693), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13821 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10675), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13822 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13823 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10623), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10800) );
  NAND4_X1 U13824 ( .A1(n10803), .A2(n10802), .A3(n10801), .A4(n10800), .ZN(
        n10811) );
  AOI22_X1 U13825 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13826 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13827 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10807) );
  INV_X1 U13828 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10804) );
  INV_X1 U13829 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12169) );
  OAI22_X1 U13830 ( .A1(n12253), .A2(n10804), .B1(n12169), .B2(n9695), .ZN(
        n10805) );
  INV_X1 U13831 ( .A(n10805), .ZN(n10806) );
  NAND4_X1 U13832 ( .A1(n10809), .A2(n10808), .A3(n10807), .A4(n10806), .ZN(
        n10810) );
  NAND2_X1 U13833 ( .A1(n10825), .A2(n13477), .ZN(n10812) );
  OAI211_X1 U13834 ( .C1(n12452), .C2(n10814), .A(n10813), .B(n10812), .ZN(
        n15510) );
  AOI22_X1 U13835 ( .A1(n10857), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13836 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10693), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13837 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U13838 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U13839 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10815) );
  NAND4_X1 U13840 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(
        n10824) );
  AOI22_X1 U13841 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n13834), .ZN(n10822) );
  AOI22_X1 U13842 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13843 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13844 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10819) );
  NAND4_X1 U13845 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        n10823) );
  NAND2_X1 U13846 ( .A1(n10825), .A2(n13484), .ZN(n10826) );
  OAI211_X1 U13847 ( .C1(n12452), .C2(n21116), .A(n10827), .B(n10826), .ZN(
        n15489) );
  NAND2_X1 U13848 ( .A1(n10162), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13849 ( .A1(n10857), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10828) );
  NAND2_X1 U13850 ( .A1(n10162), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13851 ( .A1(n10857), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U13852 ( .A1(n10857), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10833) );
  OAI21_X1 U13853 ( .B1(n12452), .B2(n10834), .A(n10833), .ZN(n15443) );
  AND2_X2 U13854 ( .A1(n15095), .A2(n15443), .ZN(n15445) );
  AOI22_X1 U13855 ( .A1(n10857), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10835) );
  OAI21_X1 U13856 ( .B1(n12452), .B2(n19975), .A(n10835), .ZN(n15085) );
  NAND2_X1 U13857 ( .A1(n10162), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U13858 ( .A1(n10857), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10836) );
  AND2_X1 U13859 ( .A1(n10837), .A2(n10836), .ZN(n15420) );
  INV_X1 U13860 ( .A(n15420), .ZN(n10838) );
  NAND2_X1 U13861 ( .A1(n10162), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13862 ( .A1(n10857), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13863 ( .A1(n10857), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10841) );
  OAI21_X1 U13864 ( .B1(n12452), .B2(n19979), .A(n10841), .ZN(n14906) );
  NAND2_X1 U13865 ( .A1(n14907), .A2(n14906), .ZN(n14889) );
  NAND2_X1 U13866 ( .A1(n10162), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13867 ( .A1(n10857), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10842) );
  AND2_X1 U13868 ( .A1(n10843), .A2(n10842), .ZN(n14890) );
  NAND2_X1 U13869 ( .A1(n10162), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13870 ( .A1(n10857), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10844) );
  AND2_X1 U13871 ( .A1(n10845), .A2(n10844), .ZN(n15060) );
  NAND2_X1 U13872 ( .A1(n10162), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U13873 ( .A1(n10857), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10847) );
  AND2_X1 U13874 ( .A1(n10848), .A2(n10847), .ZN(n14876) );
  AOI22_X1 U13875 ( .A1(n10857), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10849) );
  OAI21_X1 U13876 ( .B1(n12452), .B2(n10850), .A(n10849), .ZN(n15047) );
  AOI22_X1 U13877 ( .A1(n10857), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10851) );
  OAI21_X1 U13878 ( .B1(n12452), .B2(n19989), .A(n10851), .ZN(n12607) );
  NAND2_X1 U13879 ( .A1(n12606), .A2(n12607), .ZN(n12605) );
  NAND2_X1 U13880 ( .A1(n10162), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13881 ( .A1(n10857), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10852) );
  AND2_X1 U13882 ( .A1(n10853), .A2(n10852), .ZN(n14865) );
  NOR2_X2 U13883 ( .A1(n12605), .A2(n14865), .ZN(n12556) );
  NAND2_X1 U13884 ( .A1(n10162), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13885 ( .A1(n10857), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10854) );
  AND2_X1 U13886 ( .A1(n10855), .A2(n10854), .ZN(n12557) );
  INV_X1 U13887 ( .A(n12557), .ZN(n10856) );
  AOI22_X1 U13888 ( .A1(n10857), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10858) );
  OAI21_X1 U13889 ( .B1(n12452), .B2(n10859), .A(n10858), .ZN(n10860) );
  NAND2_X1 U13890 ( .A1(n10236), .A2(n10860), .ZN(n12455) );
  OR2_X1 U13891 ( .A1(n10236), .A2(n10860), .ZN(n10861) );
  OAI22_X1 U13892 ( .A1(n15315), .A2(n19174), .B1(n19154), .B2(n15308), .ZN(
        n10862) );
  INV_X1 U13893 ( .A(n10862), .ZN(n10892) );
  INV_X1 U13894 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12693) );
  INV_X1 U13895 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12734) );
  NAND2_X1 U13896 ( .A1(n12693), .A2(n12734), .ZN(n10863) );
  MUX2_X1 U13897 ( .A(n12112), .B(n10863), .S(n9661), .Z(n12279) );
  MUX2_X1 U13898 ( .A(n10865), .B(n10864), .S(n12221), .Z(n12210) );
  MUX2_X1 U13899 ( .A(n12210), .B(P2_EBX_REG_3__SCAN_IN), .S(n9661), .Z(n10866) );
  MUX2_X1 U13900 ( .A(n12209), .B(n12132), .S(n10421), .Z(n10868) );
  MUX2_X1 U13901 ( .A(n10868), .B(P2_EBX_REG_4__SCAN_IN), .S(n9660), .Z(n12288) );
  NOR2_X2 U13902 ( .A1(n12290), .A2(n12288), .ZN(n12293) );
  INV_X1 U13903 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13153) );
  MUX2_X1 U13904 ( .A(n12159), .B(n13153), .S(n9661), .Z(n12292) );
  INV_X1 U13905 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19130) );
  MUX2_X1 U13906 ( .A(n12181), .B(n19130), .S(n9661), .Z(n12300) );
  INV_X1 U13907 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13199) );
  MUX2_X1 U13908 ( .A(n12433), .B(n13199), .S(n9660), .Z(n12309) );
  INV_X1 U13909 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13216) );
  INV_X1 U13910 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10870) );
  NOR2_X1 U13911 ( .A1(n10869), .A2(n10870), .ZN(n12305) );
  INV_X1 U13912 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10871) );
  NAND2_X1 U13913 ( .A1(n13216), .A2(n12320), .ZN(n12330) );
  NAND2_X1 U13914 ( .A1(n9661), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10872) );
  OAI21_X1 U13915 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n9661), .ZN(n10873) );
  INV_X1 U13916 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n13648) );
  NAND2_X1 U13917 ( .A1(n9660), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12342) );
  INV_X1 U13918 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10874) );
  INV_X1 U13919 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10875) );
  NOR2_X1 U13920 ( .A1(n10869), .A2(n10875), .ZN(n12337) );
  INV_X1 U13921 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n14997) );
  OR2_X2 U13922 ( .A1(n12365), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12387) );
  NAND2_X2 U13923 ( .A1(n12387), .A2(n12435), .ZN(n12336) );
  NAND2_X1 U13924 ( .A1(n9661), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12385) );
  INV_X1 U13925 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n14893) );
  NOR2_X1 U13926 ( .A1(n10869), .A2(n14893), .ZN(n12391) );
  INV_X1 U13927 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14962) );
  INV_X1 U13928 ( .A(n12401), .ZN(n12406) );
  NAND2_X1 U13929 ( .A1(n12435), .A2(n12406), .ZN(n10877) );
  NAND2_X1 U13930 ( .A1(n9660), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10876) );
  INV_X1 U13931 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10878) );
  NOR2_X1 U13932 ( .A1(n10869), .A2(n10878), .ZN(n12416) );
  NAND2_X1 U13933 ( .A1(n9660), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12428) );
  NAND2_X1 U13934 ( .A1(n9661), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10879) );
  INV_X1 U13935 ( .A(n12430), .ZN(n12431) );
  INV_X1 U13936 ( .A(n10883), .ZN(n10880) );
  INV_X1 U13937 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16273) );
  NOR2_X1 U13938 ( .A1(n10880), .A2(n16273), .ZN(n10881) );
  NAND2_X1 U13939 ( .A1(n12683), .A2(n16417), .ZN(n16272) );
  NAND2_X1 U13940 ( .A1(n10883), .A2(n16273), .ZN(n10884) );
  OR2_X1 U13941 ( .A1(n12618), .A2(n10884), .ZN(n10885) );
  NOR2_X1 U13942 ( .A1(n19632), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19602) );
  INV_X1 U13943 ( .A(n19602), .ZN(n19923) );
  NOR2_X1 U13944 ( .A1(n19932), .A2(n19923), .ZN(n16413) );
  NAND2_X1 U13945 ( .A1(n16424), .A2(n19632), .ZN(n20008) );
  NOR2_X1 U13946 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20008), .ZN(n12615) );
  NAND2_X1 U13947 ( .A1(n19129), .A2(n19929), .ZN(n10886) );
  OR2_X1 U13948 ( .A1(n16413), .A2(n10886), .ZN(n10887) );
  AOI22_X1 U13949 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19183), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19170), .ZN(n10888) );
  OAI21_X1 U13950 ( .B1(n12431), .B2(n19194), .A(n10888), .ZN(n10889) );
  INV_X1 U13951 ( .A(n10889), .ZN(n10891) );
  NAND2_X1 U13952 ( .A1(n19188), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19097) );
  NAND2_X1 U13953 ( .A1(n19198), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10890) );
  NAND2_X1 U13954 ( .A1(n10893), .A2(n10216), .ZN(P2_U2825) );
  NAND2_X1 U13955 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11057) );
  INV_X1 U13956 ( .A(n11057), .ZN(n10894) );
  NAND2_X1 U13957 ( .A1(n10894), .A2(n20663), .ZN(n20632) );
  NAND2_X1 U13958 ( .A1(n11057), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10895) );
  AND2_X2 U13959 ( .A1(n10912), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12965) );
  NAND2_X2 U13960 ( .A1(n12965), .A2(n10914), .ZN(n11155) );
  INV_X1 U13961 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10899) );
  INV_X1 U13962 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10896) );
  AND2_X2 U13963 ( .A1(n10896), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10916) );
  NAND2_X1 U13964 ( .A1(n11003), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10898) );
  NAND2_X1 U13965 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10897) );
  OAI211_X1 U13966 ( .C1(n11155), .C2(n10899), .A(n10898), .B(n10897), .ZN(
        n10900) );
  INV_X1 U13967 ( .A(n10900), .ZN(n10907) );
  NAND2_X2 U13968 ( .A1(n10903), .A2(n12964), .ZN(n11002) );
  AOI22_X1 U13969 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13970 ( .A1(n11814), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10905) );
  AND2_X2 U13971 ( .A1(n12963), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13165) );
  NAND2_X2 U13972 ( .A1(n13165), .A2(n10052), .ZN(n10952) );
  NAND2_X1 U13973 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10904) );
  INV_X1 U13974 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11565) );
  NAND2_X4 U13975 ( .A1(n12963), .A2(n10908), .ZN(n11849) );
  INV_X1 U13976 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11386) );
  INV_X1 U13977 ( .A(n10909), .ZN(n10920) );
  NAND2_X4 U13978 ( .A1(n10916), .A2(n12963), .ZN(n11906) );
  AOI22_X1 U13980 ( .A1(n11138), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10919) );
  NOR2_X2 U13981 ( .A1(n10910), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10913) );
  AOI22_X1 U13982 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10918) );
  NAND2_X4 U13983 ( .A1(n10913), .A2(n13177), .ZN(n11845) );
  AOI22_X1 U13984 ( .A1(n11139), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11130), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13985 ( .A1(n11814), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10928) );
  INV_X2 U13986 ( .A(n11002), .ZN(n11923) );
  AOI22_X1 U13987 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10957), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10927) );
  NAND2_X1 U13988 ( .A1(n11021), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10923) );
  NAND2_X1 U13989 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10922) );
  OAI211_X1 U13990 ( .C1(n11155), .C2(n11811), .A(n10923), .B(n10922), .ZN(
        n10924) );
  INV_X1 U13991 ( .A(n10924), .ZN(n10926) );
  NAND2_X1 U13992 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10925) );
  AOI22_X1 U13993 ( .A1(n11003), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13994 ( .A1(n11130), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10931) );
  INV_X4 U13995 ( .A(n11849), .ZN(n11881) );
  AOI22_X1 U13996 ( .A1(n11138), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11881), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10930) );
  INV_X1 U13997 ( .A(n11047), .ZN(n10946) );
  AOI22_X1 U13998 ( .A1(n11814), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11923), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13999 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10940) );
  INV_X1 U14000 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10936) );
  NAND2_X1 U14001 ( .A1(n11003), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10935) );
  NAND2_X1 U14002 ( .A1(n11130), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10934) );
  OAI211_X1 U14003 ( .C1(n11155), .C2(n10936), .A(n10935), .B(n10934), .ZN(
        n10937) );
  INV_X1 U14004 ( .A(n10937), .ZN(n10939) );
  NAND2_X1 U14005 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10938) );
  AOI22_X1 U14006 ( .A1(n11129), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11139), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U14007 ( .A1(n11138), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11676), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U14008 ( .A1(n11021), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U14009 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10942) );
  INV_X1 U14010 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11641) );
  INV_X1 U14011 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11870) );
  OAI22_X1 U14012 ( .A1(n11155), .A2(n11641), .B1(n11002), .B2(n11870), .ZN(
        n10947) );
  INV_X1 U14013 ( .A(n10947), .ZN(n10956) );
  AOI22_X1 U14014 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11028), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10955) );
  INV_X1 U14015 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11310) );
  NAND2_X1 U14016 ( .A1(n11003), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10949) );
  NAND2_X1 U14017 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10948) );
  OAI211_X1 U14018 ( .C1(n11031), .C2(n11310), .A(n10949), .B(n10948), .ZN(
        n10950) );
  INV_X1 U14019 ( .A(n10950), .ZN(n10954) );
  INV_X1 U14020 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U14021 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n11130), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U14022 ( .A1(n11676), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10957), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U14023 ( .A1(n11129), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U14024 ( .A1(n11138), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10960) );
  NAND2_X1 U14025 ( .A1(n20285), .A2(n11965), .ZN(n10965) );
  NAND2_X1 U14026 ( .A1(n10967), .A2(n10966), .ZN(n11001) );
  NAND2_X1 U14027 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10969) );
  OAI22_X1 U14028 ( .A1(n11031), .A2(n11905), .B1(n11002), .B2(n11672), .ZN(
        n10974) );
  INV_X1 U14029 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10972) );
  NAND2_X1 U14030 ( .A1(n11003), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10971) );
  NAND2_X1 U14031 ( .A1(n11130), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10970) );
  OAI211_X1 U14032 ( .C1(n11155), .C2(n10972), .A(n10971), .B(n10970), .ZN(
        n10973) );
  OAI22_X1 U14033 ( .A1(n11917), .A2(n11919), .B1(n11845), .B2(n11502), .ZN(
        n10976) );
  INV_X1 U14034 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11915) );
  OAI22_X1 U14035 ( .A1(n11906), .A2(n11915), .B1(n11904), .B2(n11907), .ZN(
        n10975) );
  NOR2_X1 U14036 ( .A1(n10976), .A2(n10975), .ZN(n10983) );
  NAND2_X1 U14037 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10981) );
  NAND2_X1 U14038 ( .A1(n11021), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10980) );
  NAND2_X1 U14039 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10979) );
  NAND2_X1 U14040 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10978) );
  INV_X1 U14041 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11580) );
  INV_X1 U14042 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U14043 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10986) );
  OAI211_X1 U14044 ( .C1(n11155), .C2(n11580), .A(n10987), .B(n10986), .ZN(
        n10988) );
  INV_X1 U14045 ( .A(n10988), .ZN(n10992) );
  AOI22_X1 U14046 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U14047 ( .A1(n11814), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10990) );
  NAND2_X1 U14048 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10989) );
  NAND4_X1 U14049 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n10998) );
  AOI22_X1 U14050 ( .A1(n9659), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U14051 ( .A1(n11138), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10996) );
  INV_X1 U14052 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11588) );
  INV_X1 U14053 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11778) );
  OAI22_X1 U14054 ( .A1(n11917), .A2(n11588), .B1(n11904), .B2(n11778), .ZN(
        n10993) );
  INV_X1 U14055 ( .A(n10993), .ZN(n10995) );
  AOI22_X1 U14056 ( .A1(n11130), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10994) );
  NAND2_X1 U14057 ( .A1(n11050), .A2(n20272), .ZN(n11000) );
  NAND2_X1 U14058 ( .A1(n11040), .A2(n20285), .ZN(n13221) );
  NAND3_X2 U14059 ( .A1(n11001), .A2(n11000), .A3(n10999), .ZN(n11063) );
  NAND2_X1 U14060 ( .A1(n11003), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11005) );
  NAND2_X1 U14061 ( .A1(n11130), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11004) );
  OAI211_X1 U14062 ( .C1(n11155), .C2(n11694), .A(n11005), .B(n11004), .ZN(
        n11006) );
  NAND2_X1 U14063 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11011) );
  NAND2_X1 U14064 ( .A1(n11021), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11010) );
  NAND2_X1 U14065 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11009) );
  NAND2_X1 U14066 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11008) );
  NAND2_X1 U14067 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11014) );
  NAND2_X1 U14068 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11013) );
  OAI211_X1 U14069 ( .C1(n11701), .C2(n10952), .A(n11014), .B(n11013), .ZN(
        n11015) );
  INV_X1 U14070 ( .A(n11015), .ZN(n11016) );
  NAND4_X4 U14071 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n11016), .ZN(
        n20246) );
  AOI22_X1 U14072 ( .A1(n11021), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14073 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11138), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U14074 ( .A1(n11139), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11881), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11024) );
  NAND3_X1 U14075 ( .A1(n11026), .A2(n11025), .A3(n11024), .ZN(n11039) );
  INV_X1 U14076 ( .A(n11155), .ZN(n11027) );
  AOI22_X1 U14077 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11923), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U14078 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11129), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U14079 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11030) );
  NAND2_X1 U14080 ( .A1(n11130), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11029) );
  OAI211_X1 U14081 ( .C1(n11031), .C2(n11731), .A(n11030), .B(n11029), .ZN(
        n11032) );
  INV_X1 U14082 ( .A(n11032), .ZN(n11035) );
  NAND4_X1 U14083 ( .A1(n11037), .A2(n11036), .A3(n11035), .A4(n11034), .ZN(
        n11038) );
  INV_X4 U14084 ( .A(n11067), .ZN(n13352) );
  AND2_X2 U14085 ( .A1(n13226), .A2(n20272), .ZN(n13029) );
  AND2_X4 U14086 ( .A1(n11067), .A2(n20246), .ZN(n14043) );
  INV_X1 U14087 ( .A(n13221), .ZN(n11042) );
  NOR2_X2 U14088 ( .A1(n20246), .A2(n11067), .ZN(n12969) );
  INV_X1 U14089 ( .A(n11965), .ZN(n14305) );
  NAND2_X1 U14090 ( .A1(n12952), .A2(n13352), .ZN(n11044) );
  NAND2_X1 U14091 ( .A1(n9902), .A2(n20246), .ZN(n14012) );
  INV_X1 U14092 ( .A(n13029), .ZN(n11045) );
  NAND2_X1 U14093 ( .A1(n11046), .A2(n13238), .ZN(n11049) );
  NAND2_X1 U14094 ( .A1(n14305), .A2(n20285), .ZN(n11048) );
  NAND2_X1 U14095 ( .A1(n11963), .A2(n13238), .ZN(n11070) );
  NAND2_X1 U14096 ( .A1(n11969), .A2(n14073), .ZN(n13246) );
  NAND2_X1 U14097 ( .A1(n20246), .A2(n20267), .ZN(n11051) );
  NAND2_X1 U14098 ( .A1(n13246), .A2(n11051), .ZN(n12960) );
  NAND2_X1 U14099 ( .A1(n20867), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15953) );
  NAND2_X1 U14100 ( .A1(n15953), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11055) );
  OAI21_X1 U14101 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11057), .ZN(n20596) );
  NAND2_X1 U14102 ( .A1(n15953), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11075) );
  OAI21_X1 U14103 ( .B1(n13040), .B2(n20596), .A(n11075), .ZN(n11058) );
  INV_X1 U14104 ( .A(n11058), .ZN(n11059) );
  INV_X1 U14105 ( .A(n15953), .ZN(n11061) );
  MUX2_X1 U14106 ( .A(n11061), .B(n13040), .S(n20696), .Z(n11062) );
  NAND2_X1 U14107 ( .A1(n11063), .A2(n12969), .ZN(n12959) );
  NOR2_X1 U14108 ( .A1(n11046), .A2(n9902), .ZN(n11065) );
  INV_X1 U14109 ( .A(n12969), .ZN(n13343) );
  NAND2_X1 U14110 ( .A1(n13343), .A2(n12949), .ZN(n12860) );
  OAI22_X1 U14111 ( .A1(n11065), .A2(n12860), .B1(n11064), .B2(n20954), .ZN(
        n11069) );
  NAND2_X1 U14112 ( .A1(n12970), .A2(n11066), .ZN(n13248) );
  NAND2_X1 U14113 ( .A1(n11043), .A2(n20262), .ZN(n13348) );
  NAND4_X1 U14114 ( .A1(n13248), .A2(n16255), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n13348), .ZN(n11068) );
  NOR2_X1 U14115 ( .A1(n11069), .A2(n11068), .ZN(n11072) );
  NAND3_X1 U14116 ( .A1(n11070), .A2(n12972), .A3(n20262), .ZN(n11071) );
  NAND4_X1 U14117 ( .A1(n12959), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n11104) );
  INV_X1 U14118 ( .A(n11074), .ZN(n11077) );
  NAND2_X1 U14119 ( .A1(n11075), .A2(n10901), .ZN(n11076) );
  NAND2_X1 U14120 ( .A1(n11077), .A2(n11076), .ZN(n11078) );
  NAND2_X1 U14121 ( .A1(n11079), .A2(n11080), .ZN(n11212) );
  OAI21_X1 U14122 ( .B1(n11080), .B2(n11079), .A(n11212), .ZN(n13161) );
  INV_X2 U14123 ( .A(n11814), .ZN(n11908) );
  INV_X1 U14124 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11394) );
  OAI22_X1 U14125 ( .A1(n11908), .A2(n11394), .B1(n9643), .B2(n11386), .ZN(
        n11081) );
  INV_X1 U14126 ( .A(n11081), .ZN(n11089) );
  INV_X1 U14127 ( .A(n11028), .ZN(n11910) );
  INV_X2 U14128 ( .A(n11910), .ZN(n11882) );
  AOI22_X1 U14129 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11088) );
  INV_X1 U14130 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11752) );
  NAND2_X1 U14131 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11084) );
  NAND2_X1 U14132 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11083) );
  OAI211_X1 U14133 ( .C1(n11869), .C2(n11752), .A(n11084), .B(n11083), .ZN(
        n11085) );
  INV_X1 U14134 ( .A(n11085), .ZN(n11087) );
  NAND2_X1 U14135 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11086) );
  NAND4_X1 U14136 ( .A1(n11089), .A2(n11088), .A3(n11087), .A4(n11086), .ZN(
        n11101) );
  INV_X2 U14137 ( .A(n11091), .ZN(n11918) );
  AOI22_X1 U14138 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11099) );
  INV_X1 U14139 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11754) );
  INV_X1 U14140 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11092) );
  OAI22_X1 U14141 ( .A1(n11917), .A2(n11754), .B1(n11845), .B2(n11092), .ZN(
        n11093) );
  INV_X1 U14142 ( .A(n11093), .ZN(n11098) );
  AOI22_X1 U14143 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11097) );
  INV_X1 U14144 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11094) );
  INV_X1 U14145 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11753) );
  OAI22_X1 U14146 ( .A1(n11906), .A2(n11094), .B1(n11904), .B2(n11753), .ZN(
        n11095) );
  INV_X1 U14147 ( .A(n11095), .ZN(n11096) );
  NAND4_X1 U14148 ( .A1(n11099), .A2(n11098), .A3(n11097), .A4(n11096), .ZN(
        n11100) );
  NOR2_X1 U14149 ( .A1(n11101), .A2(n11100), .ZN(n13275) );
  NAND2_X1 U14150 ( .A1(n13238), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11126) );
  OR2_X1 U14152 ( .A1(n20246), .A2(n20868), .ZN(n11154) );
  OAI22_X1 U14153 ( .A1(n11994), .A2(n11394), .B1(n13275), .B2(n11154), .ZN(
        n11102) );
  INV_X1 U14154 ( .A(n11104), .ZN(n11105) );
  XNOR2_X1 U14155 ( .A(n11106), .B(n11105), .ZN(n11204) );
  NAND2_X1 U14156 ( .A1(n11204), .A2(n20868), .ZN(n11147) );
  INV_X1 U14157 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11503) );
  OAI22_X1 U14158 ( .A1(n11908), .A2(n11503), .B1(n9643), .B2(n11907), .ZN(
        n11110) );
  NAND2_X1 U14159 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11108) );
  NAND2_X1 U14160 ( .A1(n11130), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11107) );
  OAI211_X1 U14161 ( .C1(n11869), .C2(n11905), .A(n11108), .B(n11107), .ZN(
        n11109) );
  NOR2_X1 U14162 ( .A1(n11110), .A2(n11109), .ZN(n11125) );
  NAND2_X1 U14163 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11115) );
  NAND2_X1 U14164 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11114) );
  NAND2_X1 U14165 ( .A1(n11918), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11113) );
  NAND2_X1 U14166 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11112) );
  INV_X1 U14167 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11916) );
  OAI22_X1 U14168 ( .A1(n11917), .A2(n11672), .B1(n11845), .B2(n11916), .ZN(
        n11117) );
  INV_X1 U14169 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11920) );
  OAI22_X1 U14170 ( .A1(n11906), .A2(n11920), .B1(n11904), .B2(n11502), .ZN(
        n11116) );
  NOR2_X1 U14171 ( .A1(n11117), .A2(n11116), .ZN(n11123) );
  INV_X1 U14172 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11120) );
  NAND2_X1 U14173 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11119) );
  NAND2_X1 U14174 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11118) );
  OAI211_X1 U14175 ( .C1(n11120), .C2(n10952), .A(n11119), .B(n11118), .ZN(
        n11121) );
  INV_X1 U14176 ( .A(n11121), .ZN(n11122) );
  NAND4_X1 U14177 ( .A1(n11125), .A2(n11124), .A3(n11123), .A4(n11122), .ZN(
        n14434) );
  INV_X1 U14178 ( .A(n11126), .ZN(n11180) );
  INV_X1 U14179 ( .A(n14434), .ZN(n11127) );
  NAND2_X1 U14180 ( .A1(n11180), .A2(n11127), .ZN(n11174) );
  OAI22_X1 U14181 ( .A1(n11869), .A2(n11695), .B1(n9643), .B2(n11688), .ZN(
        n11128) );
  INV_X1 U14182 ( .A(n11128), .ZN(n11137) );
  AOI22_X1 U14183 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11884), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11136) );
  INV_X1 U14184 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11699) );
  NAND2_X1 U14185 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14186 ( .A1(n11130), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11131) );
  OAI211_X1 U14187 ( .C1(n11908), .C2(n11699), .A(n11132), .B(n11131), .ZN(
        n11133) );
  INV_X1 U14188 ( .A(n11133), .ZN(n11135) );
  NAND2_X1 U14189 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11134) );
  NAND4_X1 U14190 ( .A1(n11137), .A2(n11136), .A3(n11135), .A4(n11134), .ZN(
        n11145) );
  AOI22_X1 U14191 ( .A1(n11881), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14192 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11926), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U14193 ( .A1(n11918), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11141) );
  AOI22_X1 U14194 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11140) );
  NAND4_X1 U14195 ( .A1(n11143), .A2(n11142), .A3(n11141), .A4(n11140), .ZN(
        n11144) );
  MUX2_X1 U14196 ( .A(n14430), .B(n11174), .S(n13270), .Z(n11146) );
  INV_X1 U14197 ( .A(n13270), .ZN(n11150) );
  INV_X1 U14198 ( .A(n11148), .ZN(n11149) );
  OAI211_X1 U14199 ( .C1(n11150), .C2(n20246), .A(n11149), .B(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n11151) );
  INV_X1 U14200 ( .A(n11151), .ZN(n11152) );
  INV_X1 U14201 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11371) );
  INV_X1 U14202 ( .A(n11154), .ZN(n11172) );
  AOI22_X1 U14203 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11163) );
  INV_X1 U14204 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11718) );
  INV_X1 U14205 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11722) );
  OAI22_X1 U14206 ( .A1(n9643), .A2(n11718), .B1(n11917), .B2(n11722), .ZN(
        n11156) );
  INV_X1 U14207 ( .A(n11156), .ZN(n11162) );
  NAND2_X1 U14208 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11158) );
  NAND2_X1 U14209 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11157) );
  OAI211_X1 U14210 ( .C1(n11908), .C2(n11371), .A(n11158), .B(n11157), .ZN(
        n11159) );
  INV_X1 U14211 ( .A(n11159), .ZN(n11161) );
  NAND2_X1 U14212 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11160) );
  NAND4_X1 U14213 ( .A1(n11163), .A2(n11162), .A3(n11161), .A4(n11160), .ZN(
        n11171) );
  AOI22_X1 U14214 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11169) );
  AOI22_X1 U14215 ( .A1(n11881), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11168) );
  INV_X1 U14216 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11164) );
  INV_X1 U14217 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11729) );
  OAI22_X1 U14218 ( .A1(n11906), .A2(n11164), .B1(n11845), .B2(n11729), .ZN(
        n11165) );
  INV_X1 U14219 ( .A(n11165), .ZN(n11167) );
  AOI22_X1 U14220 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11166) );
  NAND4_X1 U14221 ( .A1(n11169), .A2(n11168), .A3(n11167), .A4(n11166), .ZN(
        n11170) );
  NAND2_X1 U14222 ( .A1(n11172), .A2(n13269), .ZN(n11173) );
  OAI211_X1 U14223 ( .C1(n11994), .C2(n11371), .A(n11174), .B(n11173), .ZN(
        n11183) );
  INV_X1 U14224 ( .A(n11183), .ZN(n11175) );
  INV_X1 U14225 ( .A(n11176), .ZN(n11177) );
  NAND2_X1 U14226 ( .A1(n20301), .A2(n11179), .ZN(n13347) );
  NAND2_X1 U14227 ( .A1(n11180), .A2(n13269), .ZN(n11181) );
  OAI21_X2 U14228 ( .B1(n13347), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11181), 
        .ZN(n11182) );
  INV_X1 U14229 ( .A(n11182), .ZN(n11194) );
  NAND2_X1 U14230 ( .A1(n11195), .A2(n11194), .ZN(n11186) );
  NAND2_X1 U14231 ( .A1(n11186), .A2(n11185), .ZN(n11188) );
  NAND2_X1 U14232 ( .A1(n11188), .A2(n11187), .ZN(n11189) );
  NOR2_X1 U14233 ( .A1(n13221), .A2(n20870), .ZN(n11246) );
  INV_X1 U14234 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n11191) );
  XNOR2_X1 U14235 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13399) );
  AOI21_X1 U14236 ( .B1(n13340), .B2(n13399), .A(n11941), .ZN(n11190) );
  OAI21_X1 U14237 ( .B1(n11936), .B2(n11191), .A(n11190), .ZN(n11192) );
  AOI21_X1 U14238 ( .B1(n11246), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11192), .ZN(n11193) );
  NAND2_X1 U14239 ( .A1(n11941), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11211) );
  NAND2_X1 U14240 ( .A1(n13369), .A2(n11513), .ZN(n11200) );
  INV_X1 U14241 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11197) );
  INV_X1 U14242 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13364) );
  OAI22_X1 U14243 ( .A1(n11936), .A2(n11197), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13364), .ZN(n11198) );
  AOI21_X1 U14244 ( .B1(n11246), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11198), .ZN(n11199) );
  NAND2_X1 U14245 ( .A1(n11200), .A2(n11199), .ZN(n13017) );
  NAND2_X1 U14246 ( .A1(n20328), .A2(n11066), .ZN(n11203) );
  NAND2_X1 U14247 ( .A1(n11203), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13044) );
  INV_X1 U14248 ( .A(n11246), .ZN(n11271) );
  NAND2_X1 U14249 ( .A1(n11942), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11206) );
  NAND2_X1 U14250 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11205) );
  OAI211_X1 U14251 ( .C1(n11271), .C2(n10914), .A(n11206), .B(n11205), .ZN(
        n11207) );
  AOI21_X1 U14252 ( .B1(n20368), .B2(n11513), .A(n11207), .ZN(n11208) );
  OR2_X1 U14253 ( .A1(n13044), .A2(n11208), .ZN(n13045) );
  INV_X1 U14254 ( .A(n11208), .ZN(n13046) );
  OR2_X1 U14255 ( .A1(n13046), .A2(n11935), .ZN(n11209) );
  NAND2_X1 U14256 ( .A1(n13045), .A2(n11209), .ZN(n13016) );
  NAND2_X1 U14257 ( .A1(n13017), .A2(n13016), .ZN(n13385) );
  INV_X1 U14258 ( .A(n13040), .ZN(n11214) );
  NAND2_X1 U14259 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10233), .ZN(
        n20534) );
  NAND2_X1 U14260 ( .A1(n20662), .A2(n20534), .ZN(n11213) );
  NOR3_X1 U14261 ( .A1(n20662), .A2(n20663), .A3(n20592), .ZN(n20807) );
  NAND2_X1 U14262 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20807), .ZN(
        n20857) );
  AOI22_X1 U14263 ( .A1(n11214), .A2(n20542), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15953), .ZN(n11215) );
  INV_X1 U14264 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11791) );
  OAI22_X1 U14265 ( .A1(n11869), .A2(n11791), .B1(n9643), .B2(n11778), .ZN(
        n11218) );
  INV_X1 U14266 ( .A(n11218), .ZN(n11225) );
  AOI22_X1 U14267 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11881), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11224) );
  INV_X1 U14268 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11420) );
  NAND2_X1 U14269 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11220) );
  NAND2_X1 U14270 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11219) );
  OAI211_X1 U14271 ( .C1(n11908), .C2(n11420), .A(n11220), .B(n11219), .ZN(
        n11221) );
  INV_X1 U14272 ( .A(n11221), .ZN(n11223) );
  NAND2_X1 U14273 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11222) );
  NAND4_X1 U14274 ( .A1(n11225), .A2(n11224), .A3(n11223), .A4(n11222), .ZN(
        n11231) );
  AOI22_X1 U14275 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11926), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11229) );
  INV_X2 U14276 ( .A(n11082), .ZN(n11924) );
  AOI22_X1 U14277 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11924), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14278 ( .A1(n11884), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14279 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11226) );
  NAND4_X1 U14280 ( .A1(n11229), .A2(n11228), .A3(n11227), .A4(n11226), .ZN(
        n11230) );
  AOI22_X1 U14281 ( .A1(n11989), .A2(n13499), .B1(n12003), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11232) );
  NAND2_X2 U14282 ( .A1(n11235), .A2(n11234), .ZN(n11277) );
  NAND2_X1 U14283 ( .A1(n11236), .A2(n13370), .ZN(n11237) );
  NAND2_X2 U14284 ( .A1(n11277), .A2(n11237), .ZN(n13371) );
  INV_X1 U14285 ( .A(n13371), .ZN(n11238) );
  NAND2_X1 U14286 ( .A1(n11238), .A2(n11513), .ZN(n11248) );
  INV_X1 U14287 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11244) );
  INV_X1 U14288 ( .A(n11240), .ZN(n11242) );
  INV_X1 U14289 ( .A(n11300), .ZN(n11241) );
  OAI21_X1 U14290 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11242), .A(
        n11241), .ZN(n20138) );
  AOI22_X1 U14291 ( .A1(n13340), .A2(n20138), .B1(n11941), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11243) );
  OAI21_X1 U14292 ( .B1(n11936), .B2(n11244), .A(n11243), .ZN(n11245) );
  AOI21_X1 U14293 ( .B1(n11246), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11245), .ZN(n11247) );
  NAND2_X1 U14294 ( .A1(n13306), .A2(n13305), .ZN(n13304) );
  INV_X1 U14295 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n21084) );
  INV_X1 U14296 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11451) );
  OAI22_X1 U14297 ( .A1(n21084), .A2(n11908), .B1(n9643), .B2(n11451), .ZN(
        n11249) );
  INV_X1 U14298 ( .A(n11249), .ZN(n11257) );
  AOI22_X1 U14299 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11256) );
  INV_X1 U14300 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11252) );
  NAND2_X1 U14301 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11251) );
  NAND2_X1 U14302 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11250) );
  OAI211_X1 U14303 ( .C1(n11869), .C2(n11252), .A(n11251), .B(n11250), .ZN(
        n11253) );
  INV_X1 U14304 ( .A(n11253), .ZN(n11255) );
  NAND2_X1 U14305 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11254) );
  NAND4_X1 U14306 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(
        n11266) );
  AOI22_X1 U14307 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11264) );
  INV_X1 U14308 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11808) );
  INV_X1 U14309 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11453) );
  OAI22_X1 U14310 ( .A1(n11917), .A2(n11808), .B1(n11845), .B2(n11453), .ZN(
        n11258) );
  INV_X1 U14311 ( .A(n11258), .ZN(n11263) );
  AOI22_X1 U14312 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11262) );
  INV_X1 U14313 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11259) );
  INV_X1 U14314 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11809) );
  OAI22_X1 U14315 ( .A1(n11906), .A2(n11259), .B1(n11904), .B2(n11809), .ZN(
        n11260) );
  INV_X1 U14316 ( .A(n11260), .ZN(n11261) );
  NAND4_X1 U14317 ( .A1(n11264), .A2(n11263), .A3(n11262), .A4(n11261), .ZN(
        n11265) );
  NAND2_X1 U14318 ( .A1(n11989), .A2(n13503), .ZN(n11268) );
  NAND2_X1 U14319 ( .A1(n12003), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11267) );
  XNOR2_X1 U14320 ( .A(n11277), .B(n11275), .ZN(n13498) );
  XNOR2_X1 U14321 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n11300), .ZN(
        n14240) );
  INV_X1 U14322 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16258) );
  INV_X1 U14323 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20736) );
  OAI21_X1 U14324 ( .B1(n20736), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20870), .ZN(n11270) );
  NAND2_X1 U14325 ( .A1(n11942), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11269) );
  OAI211_X1 U14326 ( .C1(n11271), .C2(n16258), .A(n11270), .B(n11269), .ZN(
        n11272) );
  OAI21_X1 U14327 ( .B1(n11935), .B2(n14240), .A(n11272), .ZN(n11273) );
  AOI21_X1 U14328 ( .B1(n13498), .B2(n11513), .A(n11274), .ZN(n13423) );
  NOR2_X2 U14329 ( .A1(n11277), .A2(n11276), .ZN(n11297) );
  AOI22_X1 U14330 ( .A1(n11814), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11882), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11285) );
  INV_X1 U14331 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11833) );
  INV_X1 U14332 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11837) );
  OAI22_X1 U14333 ( .A1(n9643), .A2(n11833), .B1(n11917), .B2(n11837), .ZN(
        n11278) );
  INV_X1 U14334 ( .A(n11278), .ZN(n11284) );
  INV_X1 U14335 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11850) );
  NAND2_X1 U14336 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11280) );
  NAND2_X1 U14337 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11279) );
  OAI211_X1 U14338 ( .C1(n11869), .C2(n11850), .A(n11280), .B(n11279), .ZN(
        n11281) );
  INV_X1 U14339 ( .A(n11281), .ZN(n11283) );
  NAND2_X1 U14340 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11282) );
  NAND4_X1 U14341 ( .A1(n11285), .A2(n11284), .A3(n11283), .A4(n11282), .ZN(
        n11293) );
  AOI22_X1 U14342 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11925), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14343 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11290) );
  INV_X1 U14344 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11286) );
  INV_X1 U14345 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11436) );
  OAI22_X1 U14346 ( .A1(n11906), .A2(n11286), .B1(n11904), .B2(n11436), .ZN(
        n11287) );
  INV_X1 U14347 ( .A(n11287), .ZN(n11289) );
  AOI22_X1 U14348 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11288) );
  NAND4_X1 U14349 ( .A1(n11291), .A2(n11290), .A3(n11289), .A4(n11288), .ZN(
        n11292) );
  NAND2_X1 U14350 ( .A1(n11989), .A2(n14412), .ZN(n11295) );
  NAND2_X1 U14351 ( .A1(n12003), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11294) );
  NAND2_X1 U14352 ( .A1(n11295), .A2(n11294), .ZN(n11296) );
  NAND2_X1 U14353 ( .A1(n11297), .A2(n11296), .ZN(n11337) );
  INV_X1 U14354 ( .A(n14403), .ZN(n11299) );
  NAND2_X1 U14355 ( .A1(n11299), .A2(n11513), .ZN(n11306) );
  NOR2_X1 U14356 ( .A1(n11301), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11302) );
  NOR2_X1 U14357 ( .A1(n11328), .A2(n11302), .ZN(n20126) );
  INV_X1 U14358 ( .A(n11941), .ZN(n11554) );
  INV_X1 U14359 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11303) );
  OAI22_X1 U14360 ( .A1(n20126), .A2(n11935), .B1(n11554), .B2(n11303), .ZN(
        n11304) );
  AOI21_X1 U14361 ( .B1(n11942), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11304), .ZN(
        n11305) );
  INV_X1 U14362 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11482) );
  INV_X1 U14363 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11874) );
  OAI22_X1 U14364 ( .A1(n11908), .A2(n11482), .B1(n9643), .B2(n11874), .ZN(
        n11307) );
  INV_X1 U14365 ( .A(n11307), .ZN(n11315) );
  AOI22_X1 U14366 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U14367 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11309) );
  NAND2_X1 U14368 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11308) );
  OAI211_X1 U14369 ( .C1(n11869), .C2(n11310), .A(n11309), .B(n11308), .ZN(
        n11311) );
  INV_X1 U14370 ( .A(n11311), .ZN(n11313) );
  NAND2_X1 U14371 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11312) );
  NAND4_X1 U14372 ( .A1(n11315), .A2(n11314), .A3(n11313), .A4(n11312), .ZN(
        n11325) );
  AOI22_X1 U14373 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11323) );
  INV_X1 U14374 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11316) );
  OAI22_X1 U14375 ( .A1(n11917), .A2(n11870), .B1(n11845), .B2(n11316), .ZN(
        n11317) );
  INV_X1 U14376 ( .A(n11317), .ZN(n11322) );
  AOI22_X1 U14377 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11321) );
  INV_X1 U14378 ( .A(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11318) );
  INV_X1 U14379 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11481) );
  OAI22_X1 U14380 ( .A1(n11906), .A2(n11318), .B1(n11904), .B2(n11481), .ZN(
        n11319) );
  INV_X1 U14381 ( .A(n11319), .ZN(n11320) );
  NAND4_X1 U14382 ( .A1(n11323), .A2(n11322), .A3(n11321), .A4(n11320), .ZN(
        n11324) );
  NAND2_X1 U14383 ( .A1(n11989), .A2(n14419), .ZN(n11327) );
  NAND2_X1 U14384 ( .A1(n12003), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11326) );
  NAND2_X1 U14385 ( .A1(n11337), .A2(n11338), .ZN(n14410) );
  INV_X1 U14386 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11334) );
  INV_X1 U14387 ( .A(n11344), .ZN(n11332) );
  INV_X1 U14388 ( .A(n11328), .ZN(n11330) );
  INV_X1 U14389 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11329) );
  NAND2_X1 U14390 ( .A1(n11330), .A2(n11329), .ZN(n11331) );
  NAND2_X1 U14391 ( .A1(n11332), .A2(n11331), .ZN(n20114) );
  AOI22_X1 U14392 ( .A1(n20114), .A2(n13340), .B1(n11941), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11333) );
  OAI21_X1 U14393 ( .B1(n11936), .B2(n11334), .A(n11333), .ZN(n11335) );
  INV_X1 U14394 ( .A(n11337), .ZN(n11340) );
  NAND2_X1 U14395 ( .A1(n11989), .A2(n14434), .ZN(n11342) );
  NAND2_X1 U14396 ( .A1(n12003), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11341) );
  NAND2_X1 U14397 ( .A1(n11342), .A2(n11341), .ZN(n11343) );
  XNOR2_X2 U14398 ( .A(n14409), .B(n11343), .ZN(n14425) );
  INV_X1 U14399 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11346) );
  OAI21_X1 U14400 ( .B1(n11344), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n11364), .ZN(n20099) );
  AOI22_X1 U14401 ( .A1(n20099), .A2(n13340), .B1(n11941), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11345) );
  OAI21_X1 U14402 ( .B1(n11936), .B2(n11346), .A(n11345), .ZN(n11347) );
  AOI21_X1 U14403 ( .B1(n14425), .B2(n11513), .A(n11347), .ZN(n13540) );
  INV_X1 U14404 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13625) );
  INV_X1 U14405 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11683) );
  OAI22_X1 U14406 ( .A1(n9643), .A2(n11693), .B1(n11845), .B2(n11683), .ZN(
        n11349) );
  INV_X1 U14407 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11696) );
  NOR2_X1 U14408 ( .A1(n10952), .A2(n11696), .ZN(n11348) );
  NOR2_X1 U14409 ( .A1(n11349), .A2(n11348), .ZN(n11353) );
  AOI22_X1 U14410 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11882), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14411 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11924), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11351) );
  NAND2_X1 U14412 ( .A1(n11814), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11350) );
  NAND4_X1 U14413 ( .A1(n11353), .A2(n11352), .A3(n11351), .A4(n11350), .ZN(
        n11359) );
  AOI22_X1 U14414 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14415 ( .A1(n11676), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14416 ( .A1(n11884), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14417 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11354) );
  NAND4_X1 U14418 ( .A1(n11357), .A2(n11356), .A3(n11355), .A4(n11354), .ZN(
        n11358) );
  OR2_X1 U14419 ( .A1(n11359), .A2(n11358), .ZN(n11360) );
  NAND2_X1 U14420 ( .A1(n11513), .A2(n11360), .ZN(n11363) );
  XNOR2_X1 U14421 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11364), .ZN(
        n14634) );
  INV_X1 U14422 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14630) );
  OAI22_X1 U14423 ( .A1(n14634), .A2(n11935), .B1(n11554), .B2(n14630), .ZN(
        n11361) );
  INV_X1 U14424 ( .A(n11361), .ZN(n11362) );
  OAI211_X1 U14425 ( .C1(n13625), .C2(n11936), .A(n11363), .B(n11362), .ZN(
        n13580) );
  AND2_X2 U14426 ( .A1(n13539), .A2(n13580), .ZN(n13578) );
  XOR2_X1 U14427 ( .A(n11383), .B(n11384), .Z(n20081) );
  AOI22_X1 U14428 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14429 ( .A1(n11881), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11925), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14430 ( .A1(n11884), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11926), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14431 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11366) );
  AND4_X1 U14432 ( .A1(n11369), .A2(n11368), .A3(n11367), .A4(n11366), .ZN(
        n11379) );
  AOI22_X1 U14433 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11876), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11378) );
  INV_X1 U14434 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11370) );
  OAI22_X1 U14435 ( .A1(n11869), .A2(n11371), .B1(n9643), .B2(n11370), .ZN(
        n11375) );
  INV_X1 U14436 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11545) );
  NAND2_X1 U14437 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11373) );
  NAND2_X1 U14438 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11372) );
  OAI211_X1 U14439 ( .C1(n11908), .C2(n11545), .A(n11373), .B(n11372), .ZN(
        n11374) );
  NOR2_X1 U14440 ( .A1(n11375), .A2(n11374), .ZN(n11377) );
  NAND2_X1 U14441 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11376) );
  NAND4_X1 U14442 ( .A1(n11379), .A2(n11378), .A3(n11377), .A4(n11376), .ZN(
        n11380) );
  AOI22_X1 U14443 ( .A1(n11513), .A2(n11380), .B1(n11941), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11382) );
  NAND2_X1 U14444 ( .A1(n11942), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11381) );
  OAI211_X1 U14445 ( .C1(n20081), .C2(n11935), .A(n11382), .B(n11381), .ZN(
        n13600) );
  XNOR2_X1 U14446 ( .A(n11406), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14617) );
  INV_X1 U14447 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14392) );
  AOI22_X1 U14448 ( .A1(n11676), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14449 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11926), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11390) );
  INV_X1 U14450 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11385) );
  OAI22_X1 U14451 ( .A1(n11917), .A2(n11386), .B1(n11845), .B2(n11385), .ZN(
        n11387) );
  INV_X1 U14452 ( .A(n11387), .ZN(n11389) );
  AOI22_X1 U14453 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11388) );
  AND4_X1 U14454 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n11400) );
  AOI22_X1 U14455 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11399) );
  OAI22_X1 U14456 ( .A1(n11908), .A2(n11565), .B1(n9643), .B2(n11753), .ZN(
        n11396) );
  NAND2_X1 U14457 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11393) );
  NAND2_X1 U14458 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11392) );
  OAI211_X1 U14459 ( .C1(n11869), .C2(n11394), .A(n11393), .B(n11392), .ZN(
        n11395) );
  NOR2_X1 U14460 ( .A1(n11396), .A2(n11395), .ZN(n11398) );
  NAND2_X1 U14461 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11397) );
  NAND4_X1 U14462 ( .A1(n11400), .A2(n11399), .A3(n11398), .A4(n11397), .ZN(
        n11401) );
  NAND2_X1 U14463 ( .A1(n11513), .A2(n11401), .ZN(n11403) );
  NAND2_X1 U14464 ( .A1(n11941), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11402) );
  OAI211_X1 U14465 ( .C1(n11936), .C2(n14392), .A(n11403), .B(n11402), .ZN(
        n11404) );
  AOI21_X1 U14466 ( .B1(n14617), .B2(n13340), .A(n11404), .ZN(n14222) );
  INV_X1 U14467 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11409) );
  OAI21_X1 U14468 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11407), .A(
        n11429), .ZN(n16120) );
  NAND2_X1 U14469 ( .A1(n16120), .A2(n13340), .ZN(n11408) );
  OAI21_X1 U14470 ( .B1(n11409), .B2(n11554), .A(n11408), .ZN(n11410) );
  AOI21_X1 U14471 ( .B1(n11942), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11410), .ZN(
        n14207) );
  AOI22_X1 U14472 ( .A1(n11884), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14473 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11925), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14474 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11924), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14475 ( .A1(n11881), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11413) );
  AND4_X1 U14476 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n11426) );
  AOI22_X1 U14477 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11880), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11425) );
  INV_X1 U14478 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11417) );
  OAI22_X1 U14479 ( .A1(n11908), .A2(n11588), .B1(n9643), .B2(n11417), .ZN(
        n11422) );
  NAND2_X1 U14480 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11419) );
  NAND2_X1 U14481 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11418) );
  OAI211_X1 U14482 ( .C1(n11869), .C2(n11420), .A(n11419), .B(n11418), .ZN(
        n11421) );
  NOR2_X1 U14483 ( .A1(n11422), .A2(n11421), .ZN(n11424) );
  NAND2_X1 U14484 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11423) );
  NAND4_X1 U14485 ( .A1(n11426), .A2(n11425), .A3(n11424), .A4(n11423), .ZN(
        n11427) );
  NAND2_X1 U14486 ( .A1(n11513), .A2(n11427), .ZN(n14301) );
  INV_X1 U14487 ( .A(n14301), .ZN(n11428) );
  NAND2_X1 U14488 ( .A1(n21148), .A2(n11428), .ZN(n11473) );
  XOR2_X1 U14489 ( .A(n14606), .B(n11474), .Z(n14608) );
  AOI22_X1 U14490 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14491 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11434) );
  INV_X1 U14492 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11430) );
  INV_X1 U14493 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11846) );
  OAI22_X1 U14494 ( .A1(n11906), .A2(n11430), .B1(n11904), .B2(n11846), .ZN(
        n11431) );
  INV_X1 U14495 ( .A(n11431), .ZN(n11433) );
  AOI22_X1 U14496 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11432) );
  AND4_X1 U14497 ( .A1(n11435), .A2(n11434), .A3(n11433), .A4(n11432), .ZN(
        n11445) );
  AOI22_X1 U14498 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11884), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11444) );
  INV_X1 U14499 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11626) );
  OAI22_X1 U14500 ( .A1(n11908), .A2(n11626), .B1(n9643), .B2(n11436), .ZN(
        n11441) );
  INV_X1 U14501 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11439) );
  NAND2_X1 U14502 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11438) );
  NAND2_X1 U14503 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11437) );
  OAI211_X1 U14504 ( .C1(n11869), .C2(n11439), .A(n11438), .B(n11437), .ZN(
        n11440) );
  NOR2_X1 U14505 ( .A1(n11441), .A2(n11440), .ZN(n11443) );
  NAND2_X1 U14506 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11442) );
  NAND4_X1 U14507 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11446) );
  AOI22_X1 U14508 ( .A1(n11513), .A2(n11446), .B1(n11941), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11448) );
  NAND2_X1 U14509 ( .A1(n11942), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11447) );
  OAI211_X1 U14510 ( .C1(n14608), .C2(n11935), .A(n11448), .B(n11447), .ZN(
        n14211) );
  XOR2_X1 U14511 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11449), .Z(
        n16109) );
  AOI22_X1 U14512 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11459) );
  INV_X1 U14513 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11450) );
  OAI22_X1 U14514 ( .A1(n11917), .A2(n11451), .B1(n11845), .B2(n11450), .ZN(
        n11452) );
  INV_X1 U14515 ( .A(n11452), .ZN(n11458) );
  INV_X1 U14516 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11454) );
  OAI22_X1 U14517 ( .A1(n11906), .A2(n11454), .B1(n11849), .B2(n11453), .ZN(
        n11455) );
  INV_X1 U14518 ( .A(n11455), .ZN(n11457) );
  AOI22_X1 U14519 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11456) );
  AND4_X1 U14520 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(
        n11468) );
  AOI22_X1 U14521 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11467) );
  INV_X1 U14522 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11460) );
  OAI22_X1 U14523 ( .A1(n11908), .A2(n11460), .B1(n9643), .B2(n11809), .ZN(
        n11464) );
  NAND2_X1 U14524 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11462) );
  NAND2_X1 U14525 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11461) );
  OAI211_X1 U14526 ( .C1(n11869), .C2(n21084), .A(n11462), .B(n11461), .ZN(
        n11463) );
  NOR2_X1 U14527 ( .A1(n11464), .A2(n11463), .ZN(n11466) );
  NAND2_X1 U14528 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11465) );
  NAND4_X1 U14529 ( .A1(n11468), .A2(n11467), .A3(n11466), .A4(n11465), .ZN(
        n11469) );
  AOI22_X1 U14530 ( .A1(n11513), .A2(n11469), .B1(n11941), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11471) );
  NAND2_X1 U14531 ( .A1(n11942), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11470) );
  OAI211_X1 U14532 ( .C1(n16109), .C2(n11935), .A(n11471), .B(n11470), .ZN(
        n14290) );
  NAND2_X1 U14533 ( .A1(n14211), .A2(n14290), .ZN(n11472) );
  XNOR2_X1 U14534 ( .A(n11497), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14590) );
  NAND2_X1 U14535 ( .A1(n14590), .A2(n13340), .ZN(n11496) );
  INV_X1 U14536 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14385) );
  INV_X1 U14537 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11475) );
  OAI22_X1 U14538 ( .A1(n11906), .A2(n11475), .B1(n11917), .B2(n11874), .ZN(
        n11476) );
  INV_X1 U14539 ( .A(n11476), .ZN(n11480) );
  AOI22_X1 U14540 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14541 ( .A1(n11918), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14542 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11477) );
  AND4_X1 U14543 ( .A1(n11480), .A2(n11479), .A3(n11478), .A4(n11477), .ZN(
        n11490) );
  AOI22_X1 U14544 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11882), .B1(
        n11881), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11489) );
  OAI22_X1 U14545 ( .A1(n11482), .A2(n11869), .B1(n9643), .B2(n11481), .ZN(
        n11486) );
  INV_X1 U14546 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U14547 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11484) );
  NAND2_X1 U14548 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11483) );
  OAI211_X1 U14549 ( .C1(n11908), .C2(n11647), .A(n11484), .B(n11483), .ZN(
        n11485) );
  NOR2_X1 U14550 ( .A1(n11486), .A2(n11485), .ZN(n11488) );
  NAND2_X1 U14551 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11487) );
  NAND4_X1 U14552 ( .A1(n11490), .A2(n11489), .A3(n11488), .A4(n11487), .ZN(
        n11491) );
  NAND2_X1 U14553 ( .A1(n11513), .A2(n11491), .ZN(n11493) );
  NAND2_X1 U14554 ( .A1(n11941), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11492) );
  OAI211_X1 U14555 ( .C1(n11936), .C2(n14385), .A(n11493), .B(n11492), .ZN(
        n11494) );
  INV_X1 U14556 ( .A(n11494), .ZN(n11495) );
  NAND2_X1 U14557 ( .A1(n11496), .A2(n11495), .ZN(n14196) );
  XOR2_X1 U14558 ( .A(n16057), .B(n11517), .Z(n16100) );
  AOI22_X1 U14559 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11926), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14560 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14561 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14562 ( .A1(n11881), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11498) );
  AND4_X1 U14563 ( .A1(n11501), .A2(n11500), .A3(n11499), .A4(n11498), .ZN(
        n11511) );
  AOI22_X1 U14564 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11884), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11510) );
  OAI22_X1 U14565 ( .A1(n11869), .A2(n11503), .B1(n9643), .B2(n11502), .ZN(
        n11507) );
  NAND2_X1 U14566 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11505) );
  NAND2_X1 U14567 ( .A1(n11918), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11504) );
  OAI211_X1 U14568 ( .C1(n11908), .C2(n11919), .A(n11505), .B(n11504), .ZN(
        n11506) );
  NOR2_X1 U14569 ( .A1(n11507), .A2(n11506), .ZN(n11509) );
  NAND2_X1 U14570 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11508) );
  NAND4_X1 U14571 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(
        n11512) );
  AOI22_X1 U14572 ( .A1(n11513), .A2(n11512), .B1(n11941), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11515) );
  NAND2_X1 U14573 ( .A1(n11942), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11514) );
  OAI211_X1 U14574 ( .C1(n16100), .C2(n11935), .A(n11515), .B(n11514), .ZN(
        n11516) );
  INV_X1 U14575 ( .A(n11516), .ZN(n14381) );
  INV_X1 U14576 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14578) );
  XNOR2_X1 U14577 ( .A(n11538), .B(n14578), .ZN(n14582) );
  NAND2_X1 U14578 ( .A1(n14582), .A2(n13340), .ZN(n11537) );
  INV_X1 U14579 ( .A(n12972), .ZN(n14825) );
  NAND2_X1 U14580 ( .A1(n11896), .A2(n11935), .ZN(n11658) );
  AOI22_X1 U14581 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11925), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14582 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11926), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14583 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11520) );
  OAI22_X1 U14584 ( .A1(n11917), .A2(n11693), .B1(n11849), .B2(n11683), .ZN(
        n11518) );
  INV_X1 U14585 ( .A(n11518), .ZN(n11519) );
  AND4_X1 U14586 ( .A1(n11522), .A2(n11521), .A3(n11520), .A4(n11519), .ZN(
        n11532) );
  AOI22_X1 U14587 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11882), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11531) );
  OAI22_X1 U14588 ( .A1(n11908), .A2(n11684), .B1(n11869), .B2(n11523), .ZN(
        n11528) );
  NAND2_X1 U14589 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11526) );
  NAND2_X1 U14590 ( .A1(n11918), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11525) );
  NAND2_X1 U14591 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11524) );
  NAND4_X1 U14592 ( .A1(n11526), .A2(n11525), .A3(n11935), .A4(n11524), .ZN(
        n11527) );
  NOR2_X1 U14593 ( .A1(n11528), .A2(n11527), .ZN(n11530) );
  NAND2_X1 U14594 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11529) );
  NAND4_X1 U14595 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11533) );
  NAND2_X1 U14596 ( .A1(n11658), .A2(n11533), .ZN(n11535) );
  AOI22_X1 U14597 ( .A1(n11942), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20870), .ZN(n11534) );
  NAND2_X1 U14598 ( .A1(n11535), .A2(n11534), .ZN(n11536) );
  XOR2_X1 U14599 ( .A(n16042), .B(n11558), .Z(n16091) );
  AOI22_X1 U14600 ( .A1(n11881), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11926), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11544) );
  INV_X1 U14601 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11539) );
  OAI22_X1 U14602 ( .A1(n11906), .A2(n11539), .B1(n11845), .B2(n11033), .ZN(
        n11540) );
  INV_X1 U14603 ( .A(n11540), .ZN(n11543) );
  AOI22_X1 U14604 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14605 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11541) );
  AND4_X1 U14606 ( .A1(n11544), .A2(n11543), .A3(n11542), .A4(n11541), .ZN(
        n11553) );
  AOI22_X1 U14607 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11884), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11552) );
  OAI22_X1 U14608 ( .A1(n11869), .A2(n11545), .B1(n9643), .B2(n11729), .ZN(
        n11549) );
  NAND2_X1 U14609 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14610 ( .A1(n11918), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11546) );
  OAI211_X1 U14611 ( .C1(n11908), .C2(n11722), .A(n11547), .B(n11546), .ZN(
        n11548) );
  NOR2_X1 U14612 ( .A1(n11549), .A2(n11548), .ZN(n11551) );
  NAND2_X1 U14613 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11550) );
  NAND4_X1 U14614 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11556) );
  INV_X1 U14615 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14370) );
  OAI22_X1 U14616 ( .A1(n11936), .A2(n14370), .B1(n11554), .B2(n16042), .ZN(
        n11555) );
  AOI21_X1 U14617 ( .B1(n11938), .B2(n11556), .A(n11555), .ZN(n11557) );
  OAI21_X1 U14618 ( .B1(n16091), .B2(n11935), .A(n11557), .ZN(n14368) );
  XNOR2_X1 U14619 ( .A(n11578), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16038) );
  AOI22_X1 U14620 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14621 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11924), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11563) );
  INV_X1 U14622 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11559) );
  OAI22_X1 U14623 ( .A1(n11917), .A2(n11753), .B1(n11845), .B2(n11559), .ZN(
        n11560) );
  INV_X1 U14624 ( .A(n11560), .ZN(n11562) );
  AOI22_X1 U14625 ( .A1(n11676), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11561) );
  AND4_X1 U14626 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n11574) );
  AOI22_X1 U14627 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11882), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11573) );
  OAI22_X1 U14628 ( .A1(n11908), .A2(n11754), .B1(n11869), .B2(n11565), .ZN(
        n11570) );
  NAND2_X1 U14629 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11568) );
  NAND2_X1 U14630 ( .A1(n11918), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11567) );
  NAND2_X1 U14631 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11566) );
  NAND4_X1 U14632 ( .A1(n11568), .A2(n11567), .A3(n11935), .A4(n11566), .ZN(
        n11569) );
  NOR2_X1 U14633 ( .A1(n11570), .A2(n11569), .ZN(n11572) );
  NAND2_X1 U14634 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11571) );
  NAND4_X1 U14635 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11576) );
  INV_X1 U14636 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14364) );
  INV_X1 U14637 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14562) );
  OAI22_X1 U14638 ( .A1(n11936), .A2(n14364), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14562), .ZN(n11575) );
  AOI21_X1 U14639 ( .B1(n11658), .B2(n11576), .A(n11575), .ZN(n11577) );
  AOI21_X1 U14640 ( .B1(n16038), .B2(n13340), .A(n11577), .ZN(n14278) );
  OAI21_X1 U14641 ( .B1(n11579), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n11617), .ZN(n16030) );
  OR2_X1 U14642 ( .A1(n16030), .A2(n11935), .ZN(n11600) );
  AOI22_X1 U14643 ( .A1(n11881), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11585) );
  INV_X1 U14644 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11790) );
  OAI22_X1 U14645 ( .A1(n11906), .A2(n11580), .B1(n11845), .B2(n11790), .ZN(
        n11581) );
  INV_X1 U14646 ( .A(n11581), .ZN(n11584) );
  AOI22_X1 U14647 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14648 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11582) );
  AND4_X1 U14649 ( .A1(n11585), .A2(n11584), .A3(n11583), .A4(n11582), .ZN(
        n11594) );
  AOI22_X1 U14650 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11884), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11593) );
  INV_X1 U14651 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11782) );
  OAI22_X1 U14652 ( .A1(n11908), .A2(n11782), .B1(n9643), .B2(n10985), .ZN(
        n11590) );
  NAND2_X1 U14653 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11587) );
  NAND2_X1 U14654 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11586) );
  OAI211_X1 U14655 ( .C1(n11869), .C2(n11588), .A(n11587), .B(n11586), .ZN(
        n11589) );
  NOR2_X1 U14656 ( .A1(n11590), .A2(n11589), .ZN(n11592) );
  NAND2_X1 U14657 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11591) );
  NAND4_X1 U14658 ( .A1(n11594), .A2(n11593), .A3(n11592), .A4(n11591), .ZN(
        n11595) );
  NAND2_X1 U14659 ( .A1(n11938), .A2(n11595), .ZN(n11598) );
  NAND2_X1 U14660 ( .A1(n11942), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U14661 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11596) );
  NAND4_X1 U14662 ( .A1(n11598), .A2(n11935), .A3(n11597), .A4(n11596), .ZN(
        n11599) );
  NAND2_X1 U14663 ( .A1(n11600), .A2(n11599), .ZN(n14272) );
  XNOR2_X1 U14664 ( .A(n11617), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14554) );
  AOI22_X1 U14665 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14666 ( .A1(n11881), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11604) );
  INV_X1 U14667 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11807) );
  OAI22_X1 U14668 ( .A1(n11906), .A2(n11811), .B1(n11845), .B2(n11807), .ZN(
        n11601) );
  INV_X1 U14669 ( .A(n11601), .ZN(n11603) );
  AOI22_X1 U14670 ( .A1(n11884), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11602) );
  AND4_X1 U14671 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11613) );
  AOI22_X1 U14672 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11882), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14673 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11609) );
  NAND2_X1 U14674 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11608) );
  NAND2_X1 U14675 ( .A1(n11814), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11607) );
  AOI21_X1 U14676 ( .B1(n11925), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n13340), .ZN(n11606) );
  AND4_X1 U14677 ( .A1(n11609), .A2(n11608), .A3(n11607), .A4(n11606), .ZN(
        n11611) );
  NAND2_X1 U14678 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11610) );
  NAND4_X1 U14679 ( .A1(n11613), .A2(n11612), .A3(n11611), .A4(n11610), .ZN(
        n11615) );
  INV_X1 U14680 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14357) );
  INV_X1 U14681 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14550) );
  OAI22_X1 U14682 ( .A1(n11936), .A2(n14357), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14550), .ZN(n11614) );
  AOI21_X1 U14683 ( .B1(n11658), .B2(n11615), .A(n11614), .ZN(n11616) );
  AOI21_X1 U14684 ( .B1(n14554), .B2(n13340), .A(n11616), .ZN(n14166) );
  INV_X1 U14685 ( .A(n11618), .ZN(n11620) );
  INV_X1 U14686 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11619) );
  NAND2_X1 U14687 ( .A1(n11620), .A2(n11619), .ZN(n11621) );
  NAND2_X1 U14688 ( .A1(n11663), .A2(n11621), .ZN(n16006) );
  INV_X1 U14689 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14352) );
  AOI22_X1 U14690 ( .A1(n11884), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14691 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11926), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14692 ( .A1(n11918), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11924), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14693 ( .A1(n11881), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11622) );
  AND4_X1 U14694 ( .A1(n11625), .A2(n11624), .A3(n11623), .A4(n11622), .ZN(
        n11635) );
  AOI22_X1 U14695 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11880), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11634) );
  OAI22_X1 U14696 ( .A1(n11155), .A2(n11626), .B1(n9643), .B2(n11846), .ZN(
        n11631) );
  NAND2_X1 U14697 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11629) );
  NAND2_X1 U14698 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11628) );
  OAI211_X1 U14699 ( .C1(n11908), .C2(n11837), .A(n11629), .B(n11628), .ZN(
        n11630) );
  NOR2_X1 U14700 ( .A1(n11631), .A2(n11630), .ZN(n11633) );
  NAND2_X1 U14701 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11632) );
  NAND4_X1 U14702 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11636) );
  NAND2_X1 U14703 ( .A1(n11938), .A2(n11636), .ZN(n11638) );
  OAI21_X1 U14704 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20736), .A(
        n20870), .ZN(n11637) );
  OAI211_X1 U14705 ( .C1(n11936), .C2(n14352), .A(n11638), .B(n11637), .ZN(
        n11639) );
  NAND2_X1 U14706 ( .A1(n11640), .A2(n11639), .ZN(n14262) );
  XNOR2_X1 U14707 ( .A(n11663), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16000) );
  NAND2_X1 U14708 ( .A1(n16000), .A2(n13340), .ZN(n11662) );
  INV_X1 U14709 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15997) );
  AOI22_X1 U14710 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11924), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14711 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14712 ( .A1(n11884), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11644) );
  INV_X1 U14713 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11868) );
  OAI22_X1 U14714 ( .A1(n11906), .A2(n11641), .B1(n11849), .B2(n11868), .ZN(
        n11642) );
  INV_X1 U14715 ( .A(n11642), .ZN(n11643) );
  AND4_X1 U14716 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11656) );
  AOI22_X1 U14717 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11882), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11655) );
  OAI22_X1 U14718 ( .A1(n11647), .A2(n11869), .B1(n11908), .B2(n11870), .ZN(
        n11652) );
  NAND2_X1 U14719 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11650) );
  NAND2_X1 U14720 ( .A1(n11918), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11649) );
  NAND2_X1 U14721 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11648) );
  NAND4_X1 U14722 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11935), .ZN(
        n11651) );
  NOR2_X1 U14723 ( .A1(n11652), .A2(n11651), .ZN(n11654) );
  NAND2_X1 U14724 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11653) );
  NAND4_X1 U14725 ( .A1(n11656), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(
        n11657) );
  NAND2_X1 U14726 ( .A1(n11658), .A2(n11657), .ZN(n11660) );
  NAND2_X1 U14727 ( .A1(n11942), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n11659) );
  OAI211_X1 U14728 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n15997), .A(n11660), 
        .B(n11659), .ZN(n11661) );
  INV_X1 U14729 ( .A(n11665), .ZN(n11667) );
  INV_X1 U14730 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14731 ( .A1(n11667), .A2(n11666), .ZN(n11668) );
  NAND2_X1 U14732 ( .A1(n11746), .A2(n11668), .ZN(n15989) );
  INV_X1 U14733 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14734 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11924), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11671) );
  OAI22_X1 U14735 ( .A1(n11869), .A2(n11919), .B1(n11845), .B2(n11903), .ZN(
        n11669) );
  INV_X1 U14736 ( .A(n11669), .ZN(n11670) );
  OAI211_X1 U14737 ( .C1(n11908), .C2(n11672), .A(n11671), .B(n11670), .ZN(
        n11673) );
  INV_X1 U14738 ( .A(n11673), .ZN(n11675) );
  AOI22_X1 U14739 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11674) );
  OAI211_X1 U14740 ( .C1(n10952), .C2(n11909), .A(n11675), .B(n11674), .ZN(
        n11682) );
  AOI22_X1 U14741 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11882), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14742 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14743 ( .A1(n11676), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14744 ( .A1(n11884), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11677) );
  NAND4_X1 U14745 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11681) );
  NOR2_X1 U14746 ( .A1(n11682), .A2(n11681), .ZN(n11715) );
  OAI22_X1 U14747 ( .A1(n11869), .A2(n11684), .B1(n9643), .B2(n11683), .ZN(
        n11685) );
  INV_X1 U14748 ( .A(n11685), .ZN(n11687) );
  AOI22_X1 U14749 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11686) );
  OAI211_X1 U14750 ( .C1(n11908), .C2(n11688), .A(n11687), .B(n11686), .ZN(
        n11689) );
  INV_X1 U14751 ( .A(n11689), .ZN(n11691) );
  AOI22_X1 U14752 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11690) );
  OAI211_X1 U14753 ( .C1(n10952), .C2(n11692), .A(n11691), .B(n11690), .ZN(
        n11708) );
  OAI22_X1 U14754 ( .A1(n11082), .A2(n11694), .B1(n11810), .B2(n11693), .ZN(
        n11706) );
  OAI22_X1 U14755 ( .A1(n11697), .A2(n11696), .B1(n11906), .B2(n11695), .ZN(
        n11705) );
  INV_X1 U14756 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11698) );
  OAI22_X1 U14757 ( .A1(n11700), .A2(n11699), .B1(n11845), .B2(n11698), .ZN(
        n11704) );
  INV_X1 U14758 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11702) );
  OAI22_X1 U14759 ( .A1(n11917), .A2(n11702), .B1(n11904), .B2(n11701), .ZN(
        n11703) );
  OR4_X1 U14760 ( .A1(n11706), .A2(n11705), .A3(n11704), .A4(n11703), .ZN(
        n11707) );
  NOR2_X1 U14761 ( .A1(n11708), .A2(n11707), .ZN(n11716) );
  XNOR2_X1 U14762 ( .A(n11715), .B(n11716), .ZN(n11712) );
  NAND2_X1 U14763 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11709) );
  NAND2_X1 U14764 ( .A1(n11935), .A2(n11709), .ZN(n11710) );
  AOI21_X1 U14765 ( .B1(n11942), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11710), .ZN(
        n11711) );
  OAI21_X1 U14766 ( .B1(n11896), .B2(n11712), .A(n11711), .ZN(n11713) );
  NAND2_X1 U14767 ( .A1(n11714), .A2(n11713), .ZN(n14342) );
  XNOR2_X1 U14768 ( .A(n11746), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14521) );
  NAND2_X1 U14769 ( .A1(n14521), .A2(n13340), .ZN(n11744) );
  NOR2_X1 U14770 ( .A1(n11716), .A2(n11715), .ZN(n11768) );
  INV_X1 U14771 ( .A(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11717) );
  OAI22_X1 U14772 ( .A1(n11908), .A2(n11718), .B1(n9643), .B2(n11717), .ZN(
        n11719) );
  INV_X1 U14773 ( .A(n11719), .ZN(n11727) );
  AOI22_X1 U14774 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11726) );
  NAND2_X1 U14775 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U14776 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11720) );
  OAI211_X1 U14777 ( .C1(n11869), .C2(n11722), .A(n11721), .B(n11720), .ZN(
        n11723) );
  INV_X1 U14778 ( .A(n11723), .ZN(n11725) );
  NAND2_X1 U14779 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11724) );
  NAND4_X1 U14780 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n11738) );
  AOI22_X1 U14781 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11736) );
  INV_X1 U14782 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11728) );
  OAI22_X1 U14783 ( .A1(n11917), .A2(n11729), .B1(n11845), .B2(n11728), .ZN(
        n11730) );
  INV_X1 U14784 ( .A(n11730), .ZN(n11735) );
  AOI22_X1 U14785 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11734) );
  OAI22_X1 U14786 ( .A1(n11906), .A2(n11731), .B1(n11904), .B2(n11033), .ZN(
        n11732) );
  INV_X1 U14787 ( .A(n11732), .ZN(n11733) );
  NAND4_X1 U14788 ( .A1(n11736), .A2(n11735), .A3(n11734), .A4(n11733), .ZN(
        n11737) );
  OR2_X1 U14789 ( .A1(n11738), .A2(n11737), .ZN(n11767) );
  XNOR2_X1 U14790 ( .A(n11768), .B(n11767), .ZN(n11742) );
  NAND2_X1 U14791 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11739) );
  NAND2_X1 U14792 ( .A1(n11935), .A2(n11739), .ZN(n11740) );
  AOI21_X1 U14793 ( .B1(n11942), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11740), .ZN(
        n11741) );
  OAI21_X1 U14794 ( .B1(n11742), .B2(n11896), .A(n11741), .ZN(n11743) );
  NAND2_X1 U14795 ( .A1(n11744), .A2(n11743), .ZN(n14155) );
  AND2_X2 U14796 ( .A1(n14154), .A2(n11745), .ZN(n14137) );
  INV_X1 U14797 ( .A(n11748), .ZN(n11750) );
  INV_X1 U14798 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11749) );
  NAND2_X1 U14799 ( .A1(n11750), .A2(n11749), .ZN(n11751) );
  NAND2_X1 U14800 ( .A1(n11804), .A2(n11751), .ZN(n14514) );
  INV_X1 U14801 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11760) );
  OAI22_X1 U14802 ( .A1(n11810), .A2(n11753), .B1(n11906), .B2(n11752), .ZN(
        n11757) );
  INV_X1 U14803 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11755) );
  OAI22_X1 U14804 ( .A1(n11910), .A2(n11755), .B1(n11869), .B2(n11754), .ZN(
        n11756) );
  AOI211_X1 U14805 ( .C1(n11814), .C2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n11757), .B(n11756), .ZN(n11759) );
  AOI22_X1 U14806 ( .A1(n11884), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11876), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11758) );
  OAI211_X1 U14807 ( .C1(n10952), .C2(n11760), .A(n11759), .B(n11758), .ZN(
        n11766) );
  AOI22_X1 U14808 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14809 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11924), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U14810 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14811 ( .A1(n11881), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11761) );
  NAND4_X1 U14812 ( .A1(n11764), .A2(n11763), .A3(n11762), .A4(n11761), .ZN(
        n11765) );
  NOR2_X1 U14813 ( .A1(n11766), .A2(n11765), .ZN(n11776) );
  NAND2_X1 U14814 ( .A1(n11768), .A2(n11767), .ZN(n11775) );
  XNOR2_X1 U14815 ( .A(n11776), .B(n11775), .ZN(n11772) );
  NAND2_X1 U14816 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11769) );
  NAND2_X1 U14817 ( .A1(n11935), .A2(n11769), .ZN(n11770) );
  AOI21_X1 U14818 ( .B1(n11942), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11770), .ZN(
        n11771) );
  OAI21_X1 U14819 ( .B1(n11772), .B2(n11896), .A(n11771), .ZN(n11773) );
  XNOR2_X1 U14820 ( .A(n11804), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14510) );
  NOR2_X1 U14821 ( .A1(n11776), .A2(n11775), .ZN(n11825) );
  INV_X1 U14822 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11777) );
  OAI22_X1 U14823 ( .A1(n11908), .A2(n11778), .B1(n9643), .B2(n11777), .ZN(
        n11779) );
  INV_X1 U14824 ( .A(n11779), .ZN(n11788) );
  AOI22_X1 U14825 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11787) );
  NAND2_X1 U14826 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U14827 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11780) );
  OAI211_X1 U14828 ( .C1(n11155), .C2(n11782), .A(n11781), .B(n11780), .ZN(
        n11783) );
  INV_X1 U14829 ( .A(n11783), .ZN(n11786) );
  NAND2_X1 U14830 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11785) );
  NAND4_X1 U14831 ( .A1(n11788), .A2(n11787), .A3(n11786), .A4(n11785), .ZN(
        n11798) );
  AOI22_X1 U14832 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11796) );
  INV_X1 U14833 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n21115) );
  OAI22_X1 U14834 ( .A1(n11917), .A2(n10985), .B1(n11845), .B2(n21115), .ZN(
        n11789) );
  INV_X1 U14835 ( .A(n11789), .ZN(n11795) );
  AOI22_X1 U14836 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11794) );
  OAI22_X1 U14837 ( .A1(n11906), .A2(n11791), .B1(n11904), .B2(n11790), .ZN(
        n11792) );
  INV_X1 U14838 ( .A(n11792), .ZN(n11793) );
  NAND4_X1 U14839 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n11797) );
  OR2_X1 U14840 ( .A1(n11798), .A2(n11797), .ZN(n11824) );
  INV_X1 U14841 ( .A(n11824), .ZN(n11799) );
  XNOR2_X1 U14842 ( .A(n11825), .B(n11799), .ZN(n11802) );
  INV_X1 U14843 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14330) );
  NAND2_X1 U14844 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11800) );
  OAI211_X1 U14845 ( .C1(n11936), .C2(n14330), .A(n11935), .B(n11800), .ZN(
        n11801) );
  AOI21_X1 U14846 ( .B1(n11802), .B2(n11938), .A(n11801), .ZN(n11803) );
  AOI21_X1 U14847 ( .B1(n14510), .B2(n13340), .A(n11803), .ZN(n14125) );
  INV_X1 U14848 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14506) );
  INV_X1 U14849 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14498) );
  NAND2_X1 U14850 ( .A1(n11805), .A2(n14498), .ZN(n11806) );
  INV_X1 U14851 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11817) );
  OAI22_X1 U14852 ( .A1(n11869), .A2(n11808), .B1(n11849), .B2(n11807), .ZN(
        n11813) );
  OAI22_X1 U14853 ( .A1(n11082), .A2(n11811), .B1(n11810), .B2(n11809), .ZN(
        n11812) );
  AOI211_X1 U14854 ( .C1(n11814), .C2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n11813), .B(n11812), .ZN(n11816) );
  AOI22_X1 U14855 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11884), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11815) );
  OAI211_X1 U14856 ( .C1(n10952), .C2(n11817), .A(n11816), .B(n11815), .ZN(
        n11823) );
  AOI22_X1 U14857 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11882), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U14858 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U14859 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11926), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14860 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11818) );
  NAND4_X1 U14861 ( .A1(n11821), .A2(n11820), .A3(n11819), .A4(n11818), .ZN(
        n11822) );
  NOR2_X1 U14862 ( .A1(n11823), .A2(n11822), .ZN(n11831) );
  NAND2_X1 U14863 ( .A1(n11825), .A2(n11824), .ZN(n11830) );
  XOR2_X1 U14864 ( .A(n11831), .B(n11830), .Z(n11828) );
  INV_X1 U14865 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14326) );
  NAND2_X1 U14866 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11826) );
  OAI211_X1 U14867 ( .C1(n11936), .C2(n14326), .A(n11935), .B(n11826), .ZN(
        n11827) );
  AOI21_X1 U14868 ( .B1(n11828), .B2(n11938), .A(n11827), .ZN(n11829) );
  XNOR2_X1 U14869 ( .A(n11863), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14487) );
  NAND2_X1 U14870 ( .A1(n14487), .A2(n13340), .ZN(n11862) );
  NOR2_X1 U14871 ( .A1(n11831), .A2(n11830), .ZN(n11892) );
  INV_X1 U14872 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11832) );
  OAI22_X1 U14873 ( .A1(n11908), .A2(n11833), .B1(n9643), .B2(n11832), .ZN(
        n11834) );
  INV_X1 U14874 ( .A(n11834), .ZN(n11843) );
  AOI22_X1 U14875 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11842) );
  NAND2_X1 U14876 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11836) );
  NAND2_X1 U14877 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11835) );
  OAI211_X1 U14878 ( .C1(n11155), .C2(n11837), .A(n11836), .B(n11835), .ZN(
        n11838) );
  INV_X1 U14879 ( .A(n11838), .ZN(n11841) );
  NAND2_X1 U14880 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11840) );
  NAND4_X1 U14881 ( .A1(n11843), .A2(n11842), .A3(n11841), .A4(n11840), .ZN(
        n11857) );
  AOI22_X1 U14882 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11855) );
  INV_X1 U14883 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11844) );
  OAI22_X1 U14884 ( .A1(n11917), .A2(n11846), .B1(n11845), .B2(n11844), .ZN(
        n11847) );
  INV_X1 U14885 ( .A(n11847), .ZN(n11854) );
  AOI22_X1 U14886 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11853) );
  INV_X1 U14887 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11848) );
  OAI22_X1 U14888 ( .A1(n11906), .A2(n11850), .B1(n11849), .B2(n11848), .ZN(
        n11851) );
  INV_X1 U14889 ( .A(n11851), .ZN(n11852) );
  NAND4_X1 U14890 ( .A1(n11855), .A2(n11854), .A3(n11853), .A4(n11852), .ZN(
        n11856) );
  OR2_X1 U14891 ( .A1(n11857), .A2(n11856), .ZN(n11891) );
  XNOR2_X1 U14892 ( .A(n11892), .B(n11891), .ZN(n11860) );
  INV_X1 U14893 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14489) );
  AOI21_X1 U14894 ( .B1(n14489), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11858) );
  AOI21_X1 U14895 ( .B1(n11942), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11858), .ZN(
        n11859) );
  OAI21_X1 U14896 ( .B1(n11860), .B2(n11896), .A(n11859), .ZN(n11861) );
  NAND2_X1 U14897 ( .A1(n11862), .A2(n11861), .ZN(n14100) );
  NAND2_X1 U14898 ( .A1(n11864), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13336) );
  INV_X1 U14899 ( .A(n11864), .ZN(n11866) );
  INV_X1 U14900 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11865) );
  NAND2_X1 U14901 ( .A1(n11866), .A2(n11865), .ZN(n11867) );
  NAND2_X1 U14902 ( .A1(n13336), .A2(n11867), .ZN(n14475) );
  INV_X1 U14903 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11879) );
  OAI22_X1 U14904 ( .A1(n11870), .A2(n11869), .B1(n9643), .B2(n11868), .ZN(
        n11871) );
  INV_X1 U14905 ( .A(n11871), .ZN(n11873) );
  AOI22_X1 U14906 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11925), .B1(
        n11926), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11872) );
  OAI211_X1 U14907 ( .C1(n11908), .C2(n11874), .A(n11873), .B(n11872), .ZN(
        n11875) );
  INV_X1 U14908 ( .A(n11875), .ZN(n11878) );
  AOI22_X1 U14909 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11877) );
  OAI211_X1 U14910 ( .C1(n10952), .C2(n11879), .A(n11878), .B(n11877), .ZN(
        n11890) );
  AOI22_X1 U14911 ( .A1(n11880), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11918), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U14912 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11881), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U14913 ( .A1(n11884), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14914 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11885) );
  NAND4_X1 U14915 ( .A1(n11888), .A2(n11887), .A3(n11886), .A4(n11885), .ZN(
        n11889) );
  NOR2_X1 U14916 ( .A1(n11890), .A2(n11889), .ZN(n11902) );
  NAND2_X1 U14917 ( .A1(n11892), .A2(n11891), .ZN(n11901) );
  XNOR2_X1 U14918 ( .A(n11902), .B(n11901), .ZN(n11897) );
  NAND2_X1 U14919 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11893) );
  NAND2_X1 U14920 ( .A1(n11935), .A2(n11893), .ZN(n11894) );
  AOI21_X1 U14921 ( .B1(n11942), .B2(P1_EAX_REG_29__SCAN_IN), .A(n11894), .ZN(
        n11895) );
  OAI21_X1 U14922 ( .B1(n11897), .B2(n11896), .A(n11895), .ZN(n11898) );
  INV_X1 U14923 ( .A(n14090), .ZN(n11900) );
  XNOR2_X1 U14924 ( .A(n13336), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14464) );
  NOR2_X1 U14925 ( .A1(n11902), .A2(n11901), .ZN(n11933) );
  OAI22_X1 U14926 ( .A1(n11906), .A2(n11905), .B1(n11904), .B2(n11903), .ZN(
        n11912) );
  OAI22_X1 U14927 ( .A1(n11910), .A2(n11909), .B1(n11908), .B2(n11907), .ZN(
        n11911) );
  AOI211_X1 U14928 ( .C1(n11027), .C2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11912), .B(n11911), .ZN(n11914) );
  AOI22_X1 U14929 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11913) );
  OAI211_X1 U14930 ( .C1(n10952), .C2(n11915), .A(n11914), .B(n11913), .ZN(
        n11931) );
  NOR2_X1 U14931 ( .A1(n11917), .A2(n11916), .ZN(n11922) );
  OAI22_X1 U14932 ( .A1(n11090), .A2(n11920), .B1(n11091), .B2(n11919), .ZN(
        n11921) );
  AOI211_X1 U14933 ( .C1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .C2(n11923), .A(
        n11922), .B(n11921), .ZN(n11929) );
  AOI22_X1 U14934 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11924), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U14935 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11927) );
  NAND3_X1 U14936 ( .A1(n11929), .A2(n11928), .A3(n11927), .ZN(n11930) );
  NOR2_X1 U14937 ( .A1(n11931), .A2(n11930), .ZN(n11932) );
  XNOR2_X1 U14938 ( .A(n11933), .B(n11932), .ZN(n11939) );
  INV_X1 U14939 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14309) );
  NAND2_X1 U14940 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11934) );
  OAI211_X1 U14941 ( .C1(n11936), .C2(n14309), .A(n11935), .B(n11934), .ZN(
        n11937) );
  AOI21_X1 U14942 ( .B1(n11939), .B2(n11938), .A(n11937), .ZN(n11940) );
  NAND2_X1 U14943 ( .A1(n14089), .A2(n14077), .ZN(n11945) );
  AOI22_X1 U14944 ( .A1(n11942), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11941), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11943) );
  INV_X1 U14945 ( .A(n11943), .ZN(n11944) );
  XNOR2_X2 U14946 ( .A(n11945), .B(n11944), .ZN(n14461) );
  XNOR2_X1 U14947 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11961) );
  NAND2_X1 U14948 ( .A1(n11967), .A2(n11961), .ZN(n11948) );
  NAND2_X1 U14949 ( .A1(n20592), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11947) );
  NAND2_X1 U14950 ( .A1(n11948), .A2(n11947), .ZN(n11958) );
  XNOR2_X1 U14951 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11957) );
  NAND2_X1 U14952 ( .A1(n11958), .A2(n11957), .ZN(n11950) );
  NAND2_X1 U14953 ( .A1(n20663), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11949) );
  NAND2_X1 U14954 ( .A1(n11950), .A2(n11949), .ZN(n11960) );
  XNOR2_X1 U14955 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11959) );
  NAND2_X1 U14956 ( .A1(n11960), .A2(n11959), .ZN(n11952) );
  NAND2_X1 U14957 ( .A1(n20662), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11951) );
  NAND2_X1 U14958 ( .A1(n11952), .A2(n11951), .ZN(n11956) );
  NOR2_X1 U14959 ( .A1(n16258), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11953) );
  INV_X1 U14960 ( .A(n11999), .ZN(n12001) );
  XNOR2_X1 U14961 ( .A(n11958), .B(n11957), .ZN(n11991) );
  XNOR2_X1 U14962 ( .A(n11960), .B(n11959), .ZN(n11997) );
  XNOR2_X1 U14963 ( .A(n11967), .B(n11961), .ZN(n11981) );
  NOR4_X1 U14964 ( .A1(n12001), .A2(n11991), .A3(n11997), .A4(n11981), .ZN(
        n11962) );
  NOR2_X1 U14965 ( .A1(n11966), .A2(n11962), .ZN(n12873) );
  NAND2_X1 U14966 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20951) );
  NAND2_X1 U14967 ( .A1(n12873), .A2(n20951), .ZN(n13218) );
  OR2_X1 U14968 ( .A1(n11946), .A2(n13218), .ZN(n12013) );
  NAND2_X1 U14969 ( .A1(n12972), .A2(n11043), .ZN(n11964) );
  AND2_X1 U14970 ( .A1(n13035), .A2(n12969), .ZN(n12962) );
  NAND2_X1 U14971 ( .A1(n11998), .A2(n11966), .ZN(n12011) );
  NAND2_X1 U14972 ( .A1(n11966), .A2(n11989), .ZN(n12009) );
  INV_X1 U14973 ( .A(n11989), .ZN(n11986) );
  INV_X1 U14974 ( .A(n11967), .ZN(n11968) );
  OAI21_X1 U14975 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20696), .A(
        n11968), .ZN(n11970) );
  NOR2_X1 U14976 ( .A1(n11986), .A2(n11970), .ZN(n11974) );
  INV_X1 U14977 ( .A(n11969), .ZN(n12867) );
  INV_X1 U14978 ( .A(n11970), .ZN(n11972) );
  NAND2_X1 U14979 ( .A1(n14305), .A2(n20246), .ZN(n11971) );
  NAND2_X1 U14980 ( .A1(n11971), .A2(n13352), .ZN(n11985) );
  OAI211_X1 U14981 ( .C1(n11043), .C2(n12867), .A(n11972), .B(n11985), .ZN(
        n11973) );
  OAI21_X1 U14982 ( .B1(n11998), .B2(n11974), .A(n11973), .ZN(n11979) );
  INV_X1 U14983 ( .A(n11979), .ZN(n11984) );
  NOR2_X1 U14984 ( .A1(n11965), .A2(n20868), .ZN(n11976) );
  NOR2_X1 U14985 ( .A1(n13352), .A2(n11986), .ZN(n11975) );
  AOI211_X1 U14986 ( .C1(n12003), .C2(n11981), .A(n11976), .B(n11975), .ZN(
        n11980) );
  INV_X1 U14987 ( .A(n11980), .ZN(n11983) );
  INV_X1 U14988 ( .A(n11976), .ZN(n11977) );
  NAND2_X1 U14989 ( .A1(n11977), .A2(n20262), .ZN(n11978) );
  AOI22_X1 U14990 ( .A1(n11981), .A2(n12000), .B1(n11980), .B2(n11979), .ZN(
        n11982) );
  AOI21_X1 U14991 ( .B1(n11984), .B2(n11983), .A(n11982), .ZN(n11993) );
  INV_X1 U14992 ( .A(n11985), .ZN(n11988) );
  NOR2_X1 U14993 ( .A1(n11986), .A2(n11991), .ZN(n11987) );
  AOI211_X1 U14994 ( .C1(n12003), .C2(n11991), .A(n11988), .B(n11987), .ZN(
        n11992) );
  NAND2_X1 U14995 ( .A1(n11989), .A2(n11988), .ZN(n11990) );
  OAI22_X1 U14996 ( .A1(n11993), .A2(n11992), .B1(n11991), .B2(n11990), .ZN(
        n11996) );
  NAND2_X1 U14997 ( .A1(n11994), .A2(n11997), .ZN(n11995) );
  AOI22_X1 U14998 ( .A1(n11998), .A2(n11997), .B1(n11996), .B2(n11995), .ZN(
        n12006) );
  NOR2_X1 U14999 ( .A1(n12003), .A2(n11999), .ZN(n12005) );
  INV_X1 U15000 ( .A(n12000), .ZN(n12002) );
  NAND3_X1 U15001 ( .A1(n12003), .A2(n12002), .A3(n12001), .ZN(n12004) );
  OAI21_X1 U15002 ( .B1(n12006), .B2(n12005), .A(n12004), .ZN(n12007) );
  AOI21_X1 U15003 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20868), .A(
        n12007), .ZN(n12008) );
  NAND2_X1 U15004 ( .A1(n12009), .A2(n12008), .ZN(n12010) );
  NAND2_X1 U15005 ( .A1(n12962), .A2(n13224), .ZN(n12012) );
  INV_X1 U15006 ( .A(n20951), .ZN(n20881) );
  NOR2_X1 U15007 ( .A1(n13231), .A2(n20881), .ZN(n12982) );
  AND2_X1 U15008 ( .A1(n14043), .A2(n12982), .ZN(n12017) );
  NOR2_X1 U15009 ( .A1(n11066), .A2(n20292), .ZN(n12016) );
  AND3_X1 U15010 ( .A1(n12970), .A2(n12016), .A3(n12015), .ZN(n13018) );
  AOI22_X1 U15011 ( .A1(n12014), .A2(n12017), .B1(n13018), .B2(n12969), .ZN(
        n12018) );
  NAND2_X1 U15012 ( .A1(n12987), .A2(n12018), .ZN(n12019) );
  AND2_X1 U15013 ( .A1(n14389), .A2(n9821), .ZN(n12020) );
  NOR2_X1 U15014 ( .A1(n13156), .A2(n13221), .ZN(n12033) );
  NOR4_X1 U15015 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12024) );
  NOR4_X1 U15016 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12023) );
  NOR4_X1 U15017 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12022) );
  NOR4_X1 U15018 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12021) );
  AND4_X1 U15019 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12030) );
  NOR4_X1 U15020 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12028) );
  NOR4_X1 U15021 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12027) );
  NOR4_X1 U15022 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12026) );
  INV_X1 U15023 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n12025) );
  AND4_X1 U15024 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n12029) );
  NAND2_X1 U15025 ( .A1(n12030), .A2(n12029), .ZN(n12031) );
  AOI22_X1 U15026 ( .A1(n14378), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n13156), .ZN(n12032) );
  INV_X1 U15027 ( .A(n12032), .ZN(n12035) );
  NAND2_X1 U15028 ( .A1(n12033), .A2(n20241), .ZN(n14304) );
  INV_X1 U15029 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19420) );
  NOR2_X1 U15030 ( .A1(n12035), .A2(n12034), .ZN(n12036) );
  INV_X2 U15031 ( .A(n12068), .ZN(n12060) );
  INV_X1 U15032 ( .A(n12056), .ZN(n12051) );
  XNOR2_X2 U15033 ( .A(n12051), .B(n12045), .ZN(n12728) );
  INV_X1 U15034 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U15035 ( .A1(n9700), .A2(n12060), .ZN(n12078) );
  INV_X1 U15036 ( .A(n12078), .ZN(n12047) );
  INV_X1 U15037 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12048) );
  NOR2_X1 U15038 ( .A1(n12050), .A2(n12049), .ZN(n12067) );
  NAND2_X1 U15039 ( .A1(n12153), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12066) );
  AND2_X1 U15040 ( .A1(n12051), .A2(n19191), .ZN(n12054) );
  AND2_X1 U15041 ( .A1(n15636), .A2(n12054), .ZN(n12053) );
  AOI22_X1 U15042 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12154), .B1(
        n19429), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12065) );
  INV_X1 U15043 ( .A(n12054), .ZN(n12055) );
  NOR2_X1 U15044 ( .A1(n12941), .A2(n12055), .ZN(n12077) );
  NAND2_X1 U15045 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12059) );
  AND2_X1 U15046 ( .A1(n12056), .A2(n19191), .ZN(n12062) );
  INV_X1 U15047 ( .A(n12062), .ZN(n12057) );
  NAND2_X1 U15048 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12058) );
  AOI22_X1 U15049 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12152), .B1(
        n19487), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12063) );
  OR2_X2 U15050 ( .A1(n12075), .A2(n12072), .ZN(n19700) );
  INV_X1 U15051 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12070) );
  INV_X1 U15052 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12942) );
  NAND2_X1 U15053 ( .A1(n19175), .A2(n15636), .ZN(n12074) );
  INV_X1 U15054 ( .A(n12071), .ZN(n12082) );
  AOI22_X1 U15055 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12140), .B1(
        n9668), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12081) );
  NAND2_X1 U15056 ( .A1(n12145), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12079) );
  INV_X1 U15057 ( .A(n12110), .ZN(n12108) );
  INV_X1 U15058 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12086) );
  INV_X1 U15059 ( .A(n12140), .ZN(n12168) );
  INV_X1 U15060 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12085) );
  OAI22_X1 U15061 ( .A1(n12086), .A2(n12168), .B1(n19700), .B2(n12085), .ZN(
        n12092) );
  INV_X1 U15062 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12090) );
  INV_X1 U15063 ( .A(n9668), .ZN(n12089) );
  INV_X1 U15064 ( .A(n19859), .ZN(n12088) );
  INV_X1 U15065 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12087) );
  OAI22_X1 U15066 ( .A1(n12090), .A2(n12089), .B1(n12088), .B2(n12087), .ZN(
        n12091) );
  NOR2_X1 U15067 ( .A1(n12092), .A2(n12091), .ZN(n12105) );
  INV_X1 U15068 ( .A(n12150), .ZN(n12094) );
  INV_X1 U15069 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12093) );
  INV_X1 U15070 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12725) );
  INV_X1 U15071 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12099) );
  NOR2_X1 U15072 ( .A1(n12101), .A2(n12100), .ZN(n12104) );
  INV_X1 U15073 ( .A(n12135), .ZN(n12102) );
  AOI22_X1 U15074 ( .A1(n12102), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12145), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12103) );
  NAND2_X1 U15075 ( .A1(n10613), .A2(n12115), .ZN(n12117) );
  OAI21_X1 U15076 ( .B1(n12117), .B2(n10598), .A(n12106), .ZN(n12121) );
  NAND2_X1 U15077 ( .A1(n12108), .A2(n12107), .ZN(n12111) );
  NAND2_X1 U15078 ( .A1(n12881), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12880) );
  INV_X1 U15079 ( .A(n12880), .ZN(n12113) );
  NAND2_X1 U15080 ( .A1(n12113), .A2(n12115), .ZN(n12116) );
  NOR2_X1 U15081 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n10613), .ZN(
        n12114) );
  XNOR2_X1 U15082 ( .A(n12115), .B(n12114), .ZN(n12916) );
  NAND2_X1 U15083 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12916), .ZN(
        n12915) );
  NAND2_X1 U15084 ( .A1(n12116), .A2(n12915), .ZN(n12122) );
  XNOR2_X1 U15085 ( .A(n21118), .B(n12122), .ZN(n13736) );
  INV_X1 U15086 ( .A(n12117), .ZN(n12119) );
  NAND3_X1 U15087 ( .A1(n12119), .A2(n10406), .A3(n12118), .ZN(n12120) );
  NAND2_X1 U15088 ( .A1(n12121), .A2(n12120), .ZN(n13734) );
  NAND2_X1 U15089 ( .A1(n13736), .A2(n13734), .ZN(n12124) );
  NAND2_X1 U15090 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12122), .ZN(
        n12123) );
  NAND2_X1 U15091 ( .A1(n12124), .A2(n12123), .ZN(n12125) );
  XNOR2_X1 U15092 ( .A(n12125), .B(n13613), .ZN(n13455) );
  AND2_X1 U15093 ( .A1(n12125), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12126) );
  INV_X1 U15094 ( .A(n12131), .ZN(n12129) );
  XNOR2_X1 U15095 ( .A(n12133), .B(n12132), .ZN(n12130) );
  INV_X1 U15096 ( .A(n12130), .ZN(n12128) );
  NAND2_X1 U15097 ( .A1(n12131), .A2(n12130), .ZN(n13607) );
  INV_X1 U15098 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12137) );
  INV_X1 U15099 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12136) );
  OAI22_X1 U15100 ( .A1(n12137), .A2(n12134), .B1(n12135), .B2(n12136), .ZN(
        n12138) );
  AOI22_X1 U15101 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n12140), .B1(
        n9668), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15102 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19859), .B1(
        n12141), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12148) );
  INV_X1 U15103 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13117) );
  INV_X1 U15104 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12143) );
  OAI22_X1 U15105 ( .A1(n13117), .A2(n12142), .B1(n19700), .B2(n12143), .ZN(
        n12144) );
  INV_X1 U15106 ( .A(n12144), .ZN(n12147) );
  NAND2_X1 U15107 ( .A1(n12145), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12146) );
  AOI22_X1 U15108 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n12150), .B1(
        n12151), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15109 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n12152), .B1(
        n19487), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12157) );
  NAND2_X1 U15110 ( .A1(n12153), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12156) );
  AOI22_X1 U15111 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n12154), .B1(
        n19429), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12155) );
  INV_X1 U15112 ( .A(n12159), .ZN(n12160) );
  NAND2_X1 U15113 ( .A1(n12160), .A2(n10406), .ZN(n12161) );
  NAND2_X1 U15114 ( .A1(n12295), .A2(n13662), .ZN(n13652) );
  INV_X1 U15115 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12166) );
  INV_X1 U15116 ( .A(n12145), .ZN(n12165) );
  INV_X1 U15117 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12164) );
  OAI22_X1 U15118 ( .A1(n12166), .A2(n12165), .B1(n12135), .B2(n12164), .ZN(
        n12167) );
  INV_X1 U15119 ( .A(n12167), .ZN(n12180) );
  INV_X1 U15120 ( .A(n19700), .ZN(n19692) );
  AOI22_X1 U15121 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19692), .B1(
        n9668), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15122 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12151), .B1(
        n12141), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12173) );
  OAI22_X1 U15123 ( .A1(n12169), .A2(n12168), .B1(n12142), .B2(n10698), .ZN(
        n12170) );
  INV_X1 U15124 ( .A(n12170), .ZN(n12172) );
  NAND2_X1 U15125 ( .A1(n12153), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12171) );
  AOI22_X1 U15126 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19859), .B1(
        n12150), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15127 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19487), .B1(
        n19429), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12178) );
  INV_X1 U15128 ( .A(n12134), .ZN(n12175) );
  NAND2_X1 U15129 ( .A1(n12175), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12177) );
  AOI22_X1 U15130 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12152), .B1(
        n12154), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12176) );
  NAND3_X1 U15131 ( .A1(n12180), .A2(n10217), .A3(n10237), .ZN(n12184) );
  INV_X1 U15132 ( .A(n12181), .ZN(n12182) );
  NAND2_X1 U15133 ( .A1(n12182), .A2(n10406), .ZN(n12183) );
  INV_X1 U15134 ( .A(n12190), .ZN(n12185) );
  NAND2_X1 U15135 ( .A1(n12187), .A2(n12190), .ZN(n12188) );
  INV_X1 U15136 ( .A(n12295), .ZN(n12189) );
  NAND2_X1 U15137 ( .A1(n12196), .A2(n13654), .ZN(n12194) );
  NAND2_X1 U15138 ( .A1(n13655), .A2(n12302), .ZN(n12193) );
  INV_X1 U15139 ( .A(n13654), .ZN(n12191) );
  NAND2_X1 U15140 ( .A1(n12191), .A2(n12190), .ZN(n12192) );
  OAI211_X1 U15141 ( .C1(n13655), .C2(n12194), .A(n12193), .B(n12192), .ZN(
        n15600) );
  NAND2_X1 U15142 ( .A1(n15600), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15602) );
  INV_X1 U15143 ( .A(n13655), .ZN(n12195) );
  NAND2_X1 U15144 ( .A1(n12195), .A2(n13654), .ZN(n12197) );
  NAND2_X1 U15145 ( .A1(n12197), .A2(n12196), .ZN(n12198) );
  NAND2_X1 U15146 ( .A1(n12199), .A2(n9942), .ZN(n12201) );
  NAND2_X1 U15147 ( .A1(n12202), .A2(n12201), .ZN(n15298) );
  AND2_X1 U15148 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15549) );
  NAND2_X1 U15149 ( .A1(n15549), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15503) );
  NAND2_X1 U15150 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12203) );
  NOR2_X1 U15151 ( .A1(n15503), .A2(n12203), .ZN(n15508) );
  INV_X1 U15152 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15507) );
  NAND2_X1 U15153 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15450) );
  AND2_X1 U15154 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12486) );
  INV_X1 U15155 ( .A(n15185), .ZN(n12204) );
  NAND2_X1 U15156 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15411) );
  INV_X1 U15157 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15409) );
  INV_X1 U15158 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15365) );
  INV_X1 U15159 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15323) );
  NAND2_X1 U15160 ( .A1(n12508), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12205) );
  OAI21_X1 U15161 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20042), .A(
        n12206), .ZN(n12258) );
  MUX2_X1 U15162 ( .A(n12881), .B(n12258), .S(n12221), .Z(n12274) );
  INV_X1 U15163 ( .A(n12214), .ZN(n12208) );
  OAI21_X1 U15164 ( .B1(n12274), .B2(n12208), .A(n12207), .ZN(n12212) );
  NOR2_X1 U15165 ( .A1(n12210), .A2(n12209), .ZN(n12211) );
  AOI21_X1 U15166 ( .B1(n12212), .B2(n12211), .A(n12235), .ZN(n20047) );
  INV_X1 U15167 ( .A(n12213), .ZN(n12438) );
  AND2_X1 U15168 ( .A1(n10406), .A2(n19378), .ZN(n16415) );
  AND2_X1 U15169 ( .A1(n12438), .A2(n16415), .ZN(n12272) );
  NAND2_X1 U15170 ( .A1(n20047), .A2(n12272), .ZN(n12510) );
  INV_X1 U15171 ( .A(n12258), .ZN(n12218) );
  AND2_X1 U15172 ( .A1(n12214), .A2(n12218), .ZN(n12220) );
  INV_X1 U15173 ( .A(n12216), .ZN(n12217) );
  OAI211_X1 U15174 ( .C1(n10598), .C2(n12218), .A(n12215), .B(n12217), .ZN(
        n12219) );
  OAI21_X1 U15175 ( .B1(n12221), .B2(n12220), .A(n12219), .ZN(n12222) );
  NAND2_X1 U15176 ( .A1(n12229), .A2(n12222), .ZN(n12223) );
  OAI21_X1 U15177 ( .B1(n12257), .B2(n12224), .A(n12223), .ZN(n12228) );
  NAND2_X1 U15178 ( .A1(n19378), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12234) );
  MUX2_X1 U15179 ( .A(n19378), .B(n12234), .S(n12225), .Z(n12226) );
  NAND2_X1 U15180 ( .A1(n12226), .A2(n10598), .ZN(n12227) );
  NAND2_X1 U15181 ( .A1(n12228), .A2(n12227), .ZN(n12232) );
  INV_X1 U15182 ( .A(n12229), .ZN(n12230) );
  AOI21_X1 U15183 ( .B1(n12230), .B2(n10421), .A(n12235), .ZN(n12231) );
  NAND2_X1 U15184 ( .A1(n12232), .A2(n12231), .ZN(n12233) );
  MUX2_X1 U15185 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12233), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12238) );
  NAND2_X1 U15186 ( .A1(n16394), .A2(n10598), .ZN(n19278) );
  AOI21_X1 U15187 ( .B1(n12238), .B2(n12215), .A(n12237), .ZN(n12267) );
  INV_X1 U15188 ( .A(n16385), .ZN(n12239) );
  NOR2_X1 U15189 ( .A1(n16418), .A2(n12239), .ZN(n12251) );
  NOR2_X1 U15190 ( .A1(n12237), .A2(n10598), .ZN(n12461) );
  OAI21_X1 U15191 ( .B1(n12461), .B2(n19378), .A(n19422), .ZN(n12240) );
  NAND2_X1 U15192 ( .A1(n12240), .A2(n10407), .ZN(n12250) );
  INV_X1 U15193 ( .A(n12468), .ZN(n12474) );
  AND2_X1 U15194 ( .A1(n12241), .A2(n12474), .ZN(n12249) );
  NAND2_X1 U15195 ( .A1(n12242), .A2(n12243), .ZN(n12244) );
  NAND2_X1 U15196 ( .A1(n12244), .A2(n19422), .ZN(n12245) );
  NAND2_X1 U15197 ( .A1(n12245), .A2(n16415), .ZN(n12464) );
  NAND2_X1 U15198 ( .A1(n12246), .A2(n10407), .ZN(n12247) );
  NAND2_X1 U15199 ( .A1(n12704), .A2(n12247), .ZN(n12248) );
  NAND4_X1 U15200 ( .A1(n12250), .A2(n12249), .A3(n12464), .A4(n12248), .ZN(
        n12460) );
  AOI21_X1 U15201 ( .B1(n16384), .B2(n12251), .A(n12460), .ZN(n12697) );
  AOI21_X1 U15202 ( .B1(n12252), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12703) );
  NAND2_X1 U15203 ( .A1(n12253), .A2(n12703), .ZN(n12255) );
  INV_X1 U15204 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12254) );
  NAND2_X1 U15205 ( .A1(n12255), .A2(n12254), .ZN(n12256) );
  NAND2_X1 U15206 ( .A1(n12256), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20034) );
  OAI21_X1 U15207 ( .B1(n12258), .B2(n12257), .A(n16384), .ZN(n12259) );
  INV_X1 U15208 ( .A(n12259), .ZN(n12260) );
  NAND2_X1 U15209 ( .A1(n16424), .A2(n12260), .ZN(n12261) );
  NAND2_X1 U15210 ( .A1(n20034), .A2(n12261), .ZN(n20044) );
  NAND3_X1 U15211 ( .A1(n12438), .A2(n10598), .A3(n20044), .ZN(n12265) );
  MUX2_X1 U15212 ( .A(n16418), .B(n10407), .S(n10406), .Z(n12262) );
  NOR2_X1 U15213 ( .A1(n12262), .A2(n19943), .ZN(n12263) );
  NAND2_X1 U15214 ( .A1(n12263), .A2(n16384), .ZN(n12264) );
  NAND3_X1 U15215 ( .A1(n12697), .A2(n12265), .A3(n12264), .ZN(n12266) );
  AOI21_X1 U15216 ( .B1(n19278), .B2(n12267), .A(n12266), .ZN(n12270) );
  INV_X1 U15217 ( .A(n19278), .ZN(n12268) );
  NAND3_X1 U15218 ( .A1(n12268), .A2(n16385), .A3(n10408), .ZN(n12269) );
  NAND3_X1 U15219 ( .A1(n12510), .A2(n12270), .A3(n12269), .ZN(n12271) );
  INV_X1 U15220 ( .A(n12272), .ZN(n20046) );
  OAI21_X1 U15221 ( .B1(n12278), .B2(n12273), .A(n12290), .ZN(n13529) );
  MUX2_X1 U15222 ( .A(n12274), .B(n12693), .S(n9661), .Z(n19193) );
  NOR2_X1 U15223 ( .A1(n19193), .A2(n13721), .ZN(n12913) );
  NAND3_X1 U15224 ( .A1(n9660), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n12275) );
  NAND2_X1 U15225 ( .A1(n12279), .A2(n12275), .ZN(n19173) );
  INV_X1 U15226 ( .A(n19173), .ZN(n12912) );
  NAND2_X1 U15227 ( .A1(n12913), .A2(n12912), .ZN(n12276) );
  NOR2_X1 U15228 ( .A1(n12913), .A2(n12912), .ZN(n12911) );
  AOI21_X1 U15229 ( .B1(n12277), .B2(n12276), .A(n12911), .ZN(n13732) );
  INV_X1 U15230 ( .A(n12278), .ZN(n12282) );
  NAND2_X1 U15231 ( .A1(n12280), .A2(n12279), .ZN(n12281) );
  NAND2_X1 U15232 ( .A1(n12282), .A2(n12281), .ZN(n12283) );
  XNOR2_X1 U15233 ( .A(n12283), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13733) );
  NAND2_X1 U15234 ( .A1(n13732), .A2(n13733), .ZN(n12285) );
  INV_X1 U15235 ( .A(n12283), .ZN(n13571) );
  NAND2_X1 U15236 ( .A1(n13571), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12284) );
  NAND2_X1 U15237 ( .A1(n12285), .A2(n12284), .ZN(n13452) );
  AND2_X1 U15238 ( .A1(n13452), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12286) );
  OR2_X1 U15239 ( .A1(n13452), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12287) );
  INV_X1 U15240 ( .A(n12288), .ZN(n12289) );
  XNOR2_X1 U15241 ( .A(n12290), .B(n12289), .ZN(n19152) );
  XNOR2_X1 U15242 ( .A(n19152), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13611) );
  INV_X1 U15243 ( .A(n13649), .ZN(n12296) );
  NOR2_X1 U15244 ( .A1(n12293), .A2(n12292), .ZN(n12294) );
  OR2_X1 U15245 ( .A1(n12291), .A2(n12294), .ZN(n19142) );
  NAND2_X1 U15246 ( .A1(n12296), .A2(n10238), .ZN(n12299) );
  INV_X1 U15247 ( .A(n13651), .ZN(n12297) );
  NAND2_X1 U15248 ( .A1(n12297), .A2(n13662), .ZN(n12298) );
  NOR2_X1 U15249 ( .A1(n12291), .A2(n12300), .ZN(n12301) );
  OR2_X1 U15250 ( .A1(n12311), .A2(n12301), .ZN(n19131) );
  XNOR2_X1 U15251 ( .A(n12303), .B(n15604), .ZN(n15603) );
  NAND2_X1 U15252 ( .A1(n12306), .A2(n12305), .ZN(n12307) );
  AND2_X1 U15253 ( .A1(n9740), .A2(n12307), .ZN(n12315) );
  AND2_X1 U15254 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12308) );
  NAND2_X1 U15255 ( .A1(n12315), .A2(n12308), .ZN(n16335) );
  INV_X1 U15256 ( .A(n12309), .ZN(n12310) );
  XNOR2_X1 U15257 ( .A(n12311), .B(n12310), .ZN(n19122) );
  NAND2_X1 U15258 ( .A1(n19122), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16333) );
  NAND3_X1 U15259 ( .A1(n12313), .A2(P2_EBX_REG_10__SCAN_IN), .A3(n9661), .ZN(
        n12312) );
  OAI211_X1 U15260 ( .C1(n12313), .C2(P2_EBX_REG_10__SCAN_IN), .A(n12312), .B(
        n12435), .ZN(n19098) );
  OR2_X1 U15261 ( .A1(n19098), .A2(n9942), .ZN(n12314) );
  NAND2_X1 U15262 ( .A1(n12314), .A2(n15546), .ZN(n15290) );
  INV_X1 U15263 ( .A(n12315), .ZN(n13567) );
  OAI21_X1 U15264 ( .B1(n13567), .B2(n9942), .A(n12481), .ZN(n16336) );
  INV_X1 U15265 ( .A(n19122), .ZN(n12316) );
  NAND2_X1 U15266 ( .A1(n12316), .A2(n16374), .ZN(n16332) );
  AND2_X1 U15267 ( .A1(n16336), .A2(n16332), .ZN(n15286) );
  NAND2_X1 U15268 ( .A1(n9660), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12317) );
  XNOR2_X1 U15269 ( .A(n9740), .B(n12317), .ZN(n19112) );
  NAND2_X1 U15270 ( .A1(n19112), .A2(n12433), .ZN(n12318) );
  NAND2_X1 U15271 ( .A1(n12318), .A2(n15591), .ZN(n15594) );
  AND3_X1 U15272 ( .A1(n15290), .A2(n15286), .A3(n15594), .ZN(n12319) );
  INV_X1 U15273 ( .A(n12320), .ZN(n12321) );
  NAND2_X1 U15274 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n12321), .ZN(n12322) );
  NOR2_X1 U15275 ( .A1(n10869), .A2(n12322), .ZN(n12323) );
  NOR2_X1 U15276 ( .A1(n12324), .A2(n12323), .ZN(n19085) );
  AOI21_X1 U15277 ( .B1(n19085), .B2(n12433), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15275) );
  NAND2_X1 U15278 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12325) );
  OR2_X1 U15279 ( .A1(n19098), .A2(n12325), .ZN(n15289) );
  AND2_X1 U15280 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12326) );
  NAND2_X1 U15281 ( .A1(n19112), .A2(n12326), .ZN(n15593) );
  NAND2_X1 U15282 ( .A1(n15289), .A2(n15593), .ZN(n15271) );
  AND2_X1 U15283 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12327) );
  AND2_X1 U15284 ( .A1(n19085), .A2(n12327), .ZN(n15274) );
  NOR2_X1 U15285 ( .A1(n15271), .A2(n15274), .ZN(n12328) );
  NAND2_X1 U15286 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n12330), .ZN(n12331) );
  NOR2_X1 U15287 ( .A1(n10869), .A2(n12331), .ZN(n12332) );
  NOR2_X1 U15288 ( .A1(n12353), .A2(n12332), .ZN(n19074) );
  AND2_X1 U15289 ( .A1(n19074), .A2(n12433), .ZN(n12333) );
  AND2_X1 U15290 ( .A1(n12333), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15262) );
  INV_X1 U15291 ( .A(n12333), .ZN(n12334) );
  NAND2_X1 U15292 ( .A1(n12334), .A2(n15521), .ZN(n15263) );
  AND3_X1 U15293 ( .A1(n12365), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n9660), .ZN(
        n12335) );
  OR2_X1 U15294 ( .A1(n12336), .A2(n12335), .ZN(n18985) );
  OAI21_X1 U15295 ( .B1(n18985), .B2(n9942), .A(n15409), .ZN(n15176) );
  INV_X1 U15296 ( .A(n12337), .ZN(n12338) );
  XNOR2_X1 U15297 ( .A(n12339), .B(n12338), .ZN(n19004) );
  NAND2_X1 U15298 ( .A1(n19004), .A2(n12433), .ZN(n15193) );
  NAND2_X1 U15299 ( .A1(n15193), .A2(n15432), .ZN(n12341) );
  XNOR2_X1 U15300 ( .A(n12344), .B(n9764), .ZN(n19015) );
  NAND2_X1 U15301 ( .A1(n19015), .A2(n12433), .ZN(n12340) );
  INV_X1 U15302 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U15303 ( .A1(n12340), .A2(n15451), .ZN(n15201) );
  NAND2_X1 U15304 ( .A1(n12341), .A2(n15201), .ZN(n15169) );
  OR2_X1 U15305 ( .A1(n12343), .A2(n12342), .ZN(n12345) );
  AND2_X1 U15306 ( .A1(n12345), .A2(n12344), .ZN(n19024) );
  NAND2_X1 U15307 ( .A1(n19024), .A2(n12433), .ZN(n12378) );
  INV_X1 U15308 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15217) );
  NAND2_X1 U15309 ( .A1(n12378), .A2(n15217), .ZN(n15215) );
  NAND2_X1 U15310 ( .A1(n9661), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12347) );
  OAI211_X1 U15311 ( .C1(n12349), .C2(n12347), .A(n12435), .B(n12346), .ZN(
        n14931) );
  OR2_X1 U15312 ( .A1(n14931), .A2(n9942), .ZN(n12348) );
  XNOR2_X1 U15313 ( .A(n12348), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15165) );
  INV_X1 U15314 ( .A(n12349), .ZN(n12351) );
  INV_X1 U15315 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13483) );
  NAND2_X1 U15316 ( .A1(n12357), .A2(n13483), .ZN(n12359) );
  NAND3_X1 U15317 ( .A1(n12359), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n9660), .ZN(
        n12350) );
  NAND2_X1 U15318 ( .A1(n12351), .A2(n12350), .ZN(n19041) );
  OR2_X1 U15319 ( .A1(n19041), .A2(n9942), .ZN(n12352) );
  INV_X1 U15320 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15460) );
  NAND2_X1 U15321 ( .A1(n12352), .A2(n15460), .ZN(n15234) );
  INV_X1 U15322 ( .A(n12357), .ZN(n12355) );
  NAND2_X1 U15323 ( .A1(n10134), .A2(n9765), .ZN(n12354) );
  NAND2_X1 U15324 ( .A1(n12355), .A2(n12354), .ZN(n19066) );
  OR2_X1 U15325 ( .A1(n19066), .A2(n9942), .ZN(n12356) );
  INV_X1 U15326 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15527) );
  NAND2_X1 U15327 ( .A1(n12356), .A2(n15527), .ZN(n15254) );
  AND2_X1 U15328 ( .A1(n15234), .A2(n15254), .ZN(n12361) );
  NAND2_X1 U15329 ( .A1(n9660), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12358) );
  MUX2_X1 U15330 ( .A(n12358), .B(n9660), .S(n12357), .Z(n12360) );
  NAND2_X1 U15331 ( .A1(n19053), .A2(n12433), .ZN(n12373) );
  NAND2_X1 U15332 ( .A1(n12373), .A2(n15507), .ZN(n15241) );
  NAND4_X1 U15333 ( .A1(n15215), .A2(n15165), .A3(n12361), .A4(n15241), .ZN(
        n12362) );
  NOR2_X1 U15334 ( .A1(n15169), .A2(n12362), .ZN(n12367) );
  NAND2_X1 U15335 ( .A1(n9660), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12364) );
  MUX2_X1 U15336 ( .A(n12364), .B(n9661), .S(n12363), .Z(n12366) );
  NAND2_X1 U15337 ( .A1(n12366), .A2(n12365), .ZN(n18993) );
  OR2_X1 U15338 ( .A1(n18993), .A2(n9942), .ZN(n12381) );
  NAND2_X1 U15339 ( .A1(n12381), .A2(n15425), .ZN(n15172) );
  NAND3_X1 U15340 ( .A1(n15176), .A2(n12367), .A3(n15172), .ZN(n12368) );
  INV_X1 U15341 ( .A(n18985), .ZN(n12370) );
  AND2_X1 U15342 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12369) );
  NAND2_X1 U15343 ( .A1(n12370), .A2(n12369), .ZN(n15175) );
  INV_X1 U15344 ( .A(n15193), .ZN(n12372) );
  AND2_X1 U15345 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12371) );
  AND2_X1 U15346 ( .A1(n19015), .A2(n12371), .ZN(n15202) );
  AOI21_X1 U15347 ( .B1(n12372), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15202), .ZN(n15168) );
  INV_X1 U15348 ( .A(n12373), .ZN(n12374) );
  NAND2_X1 U15349 ( .A1(n12374), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15242) );
  NAND2_X1 U15350 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12375) );
  OR2_X1 U15351 ( .A1(n14931), .A2(n12375), .ZN(n15166) );
  NAND2_X1 U15352 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12376) );
  OR2_X1 U15353 ( .A1(n19041), .A2(n12376), .ZN(n15233) );
  NAND2_X1 U15354 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12377) );
  OR2_X1 U15355 ( .A1(n19066), .A2(n12377), .ZN(n15253) );
  AND4_X1 U15356 ( .A1(n15242), .A2(n15166), .A3(n15233), .A4(n15253), .ZN(
        n12380) );
  INV_X1 U15357 ( .A(n12378), .ZN(n12379) );
  NAND2_X1 U15358 ( .A1(n12379), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15167) );
  NAND4_X1 U15359 ( .A1(n15175), .A2(n15168), .A3(n12380), .A4(n15167), .ZN(
        n12382) );
  NOR2_X1 U15360 ( .A1(n12381), .A2(n15425), .ZN(n15174) );
  NOR2_X1 U15361 ( .A1(n12382), .A2(n15174), .ZN(n12383) );
  INV_X1 U15362 ( .A(n12385), .ZN(n12386) );
  NAND2_X1 U15363 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  NAND2_X1 U15364 ( .A1(n12384), .A2(n12388), .ZN(n14911) );
  INV_X1 U15365 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15393) );
  NAND2_X1 U15366 ( .A1(n12389), .A2(n15393), .ZN(n15152) );
  INV_X1 U15367 ( .A(n12389), .ZN(n12390) );
  NAND2_X1 U15368 ( .A1(n12390), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15153) );
  INV_X1 U15369 ( .A(n12391), .ZN(n12392) );
  XNOR2_X1 U15370 ( .A(n12384), .B(n12392), .ZN(n14901) );
  NAND2_X1 U15371 ( .A1(n14901), .A2(n12433), .ZN(n12393) );
  XNOR2_X1 U15372 ( .A(n12393), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15146) );
  NAND2_X1 U15373 ( .A1(n15147), .A2(n15146), .ZN(n15148) );
  OR2_X1 U15374 ( .A1(n12393), .A2(n12491), .ZN(n12394) );
  NAND3_X1 U15375 ( .A1(n12395), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n9661), .ZN(
        n12396) );
  NAND2_X1 U15376 ( .A1(n12396), .A2(n12435), .ZN(n12397) );
  OR2_X1 U15377 ( .A1(n12397), .A2(n12408), .ZN(n16307) );
  NOR2_X1 U15378 ( .A1(n16307), .A2(n9942), .ZN(n12398) );
  INV_X1 U15379 ( .A(n12398), .ZN(n12400) );
  NAND2_X1 U15380 ( .A1(n12400), .A2(n12399), .ZN(n15133) );
  AND2_X1 U15381 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n12412), .ZN(n12402) );
  NAND2_X1 U15382 ( .A1(n12435), .A2(n12403), .ZN(n16291) );
  INV_X1 U15383 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15348) );
  NAND2_X1 U15384 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12404) );
  NAND2_X1 U15385 ( .A1(n12405), .A2(n12421), .ZN(n15113) );
  NAND3_X1 U15386 ( .A1(n9661), .A2(P2_EBX_REG_27__SCAN_IN), .A3(n12406), .ZN(
        n12407) );
  NAND2_X1 U15387 ( .A1(n12415), .A2(n12407), .ZN(n12601) );
  NOR2_X1 U15388 ( .A1(n12408), .A2(n14962), .ZN(n12409) );
  NAND2_X1 U15389 ( .A1(n9660), .A2(n12409), .ZN(n12410) );
  AND2_X1 U15390 ( .A1(n12435), .A2(n12410), .ZN(n12411) );
  NAND2_X1 U15391 ( .A1(n12412), .A2(n12411), .ZN(n14886) );
  NAND2_X1 U15392 ( .A1(n12420), .A2(n15365), .ZN(n15120) );
  AND2_X1 U15393 ( .A1(n12422), .A2(n10214), .ZN(n12427) );
  INV_X1 U15394 ( .A(n12415), .ZN(n12419) );
  INV_X1 U15395 ( .A(n12416), .ZN(n12418) );
  OAI21_X1 U15396 ( .B1(n12419), .B2(n12418), .A(n12417), .ZN(n14864) );
  NAND2_X1 U15397 ( .A1(n15121), .A2(n12421), .ZN(n12574) );
  INV_X1 U15398 ( .A(n12574), .ZN(n12425) );
  INV_X1 U15399 ( .A(n12422), .ZN(n12423) );
  OAI211_X2 U15400 ( .C1(n12427), .C2(n12426), .A(n12425), .B(n12424), .ZN(
        n12542) );
  XNOR2_X1 U15401 ( .A(n12429), .B(n12428), .ZN(n12432) );
  OAI21_X1 U15402 ( .B1(n12432), .B2(n9942), .A(n12539), .ZN(n12540) );
  AOI21_X1 U15403 ( .B1(n12430), .B2(n12433), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12520) );
  INV_X1 U15404 ( .A(n12432), .ZN(n14857) );
  NAND3_X1 U15405 ( .A1(n14857), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12433), .ZN(n12541) );
  OAI21_X1 U15406 ( .B1(n12434), .B2(P2_EBX_REG_30__SCAN_IN), .A(n9660), .ZN(
        n12436) );
  NAND2_X1 U15407 ( .A1(n12436), .A2(n12435), .ZN(n16275) );
  NOR2_X1 U15408 ( .A1(n16275), .A2(n9942), .ZN(n12437) );
  NAND2_X1 U15409 ( .A1(n12438), .A2(n10421), .ZN(n20045) );
  NAND2_X1 U15410 ( .A1(n12546), .A2(n12439), .ZN(n12446) );
  AOI22_X1 U15411 ( .A1(n12440), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12443) );
  NAND2_X1 U15412 ( .A1(n12441), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12442) );
  OAI211_X1 U15413 ( .C1(n10473), .C2(n12444), .A(n12443), .B(n12442), .ZN(
        n12445) );
  INV_X1 U15414 ( .A(n12447), .ZN(n12448) );
  INV_X1 U15415 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15416 ( .A1(n10857), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12449), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12450) );
  OAI21_X1 U15417 ( .B1(n12452), .B2(n12451), .A(n12450), .ZN(n12453) );
  INV_X1 U15418 ( .A(n12453), .ZN(n12454) );
  NAND2_X1 U15419 ( .A1(n12456), .A2(n12457), .ZN(n13061) );
  NAND2_X1 U15420 ( .A1(n10578), .A2(n10598), .ZN(n12458) );
  AND2_X1 U15421 ( .A1(n13061), .A2(n12458), .ZN(n12459) );
  INV_X1 U15422 ( .A(n12460), .ZN(n12462) );
  NAND2_X1 U15423 ( .A1(n12462), .A2(n12461), .ZN(n16393) );
  NAND2_X1 U15424 ( .A1(n12463), .A2(n10598), .ZN(n13711) );
  AOI21_X1 U15425 ( .B1(n13711), .B2(n12464), .A(n10398), .ZN(n12472) );
  AND2_X1 U15426 ( .A1(n10407), .A2(n19378), .ZN(n12470) );
  INV_X1 U15427 ( .A(n12466), .ZN(n14843) );
  OAI21_X1 U15428 ( .B1(n12468), .B2(n12467), .A(n14843), .ZN(n12469) );
  OAI21_X1 U15429 ( .B1(n12465), .B2(n12470), .A(n12469), .ZN(n12471) );
  NOR2_X1 U15430 ( .A1(n12472), .A2(n12471), .ZN(n12473) );
  OAI21_X1 U15431 ( .B1(n12475), .B2(n12474), .A(n12473), .ZN(n13717) );
  NOR2_X1 U15432 ( .A1(n13717), .A2(n12691), .ZN(n12476) );
  OR2_X1 U15433 ( .A1(n12477), .A2(n12476), .ZN(n12478) );
  INV_X1 U15434 ( .A(n19370), .ZN(n15613) );
  NAND3_X1 U15435 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15310) );
  AND2_X1 U15436 ( .A1(n12477), .A2(n19129), .ZN(n19362) );
  INV_X1 U15437 ( .A(n12478), .ZN(n15461) );
  NAND2_X1 U15438 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19371) );
  OR2_X1 U15439 ( .A1(n21118), .A2(n19371), .ZN(n13745) );
  NAND2_X1 U15440 ( .A1(n15461), .A2(n13745), .ZN(n12480) );
  INV_X1 U15441 ( .A(n19362), .ZN(n12479) );
  AND2_X1 U15442 ( .A1(n12480), .A2(n12479), .ZN(n13456) );
  NAND2_X1 U15443 ( .A1(n21118), .A2(n19371), .ZN(n13746) );
  INV_X1 U15444 ( .A(n13746), .ZN(n12498) );
  NOR2_X1 U15445 ( .A1(n13662), .A2(n13656), .ZN(n15605) );
  NAND2_X1 U15446 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15605), .ZN(
        n15610) );
  NOR2_X1 U15447 ( .A1(n12481), .A2(n16374), .ZN(n12499) );
  INV_X1 U15448 ( .A(n12499), .ZN(n16364) );
  OR4_X1 U15449 ( .A1(n12498), .A2(n13613), .A3(n15610), .A4(n16364), .ZN(
        n12482) );
  NAND2_X1 U15450 ( .A1(n19370), .A2(n12482), .ZN(n12483) );
  NAND2_X1 U15451 ( .A1(n13456), .A2(n12483), .ZN(n15580) );
  AND2_X1 U15452 ( .A1(n15508), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12500) );
  INV_X1 U15453 ( .A(n12500), .ZN(n12484) );
  OR2_X1 U15454 ( .A1(n15580), .A2(n12484), .ZN(n12485) );
  NAND2_X1 U15455 ( .A1(n12485), .A2(n15565), .ZN(n15493) );
  INV_X1 U15456 ( .A(n15450), .ZN(n12487) );
  NAND2_X1 U15457 ( .A1(n12487), .A2(n12486), .ZN(n12501) );
  NAND2_X1 U15458 ( .A1(n15565), .A2(n12501), .ZN(n12488) );
  AND2_X1 U15459 ( .A1(n15493), .A2(n12488), .ZN(n15447) );
  NAND2_X1 U15460 ( .A1(n15565), .A2(n15411), .ZN(n12489) );
  AND2_X1 U15461 ( .A1(n15447), .A2(n12489), .ZN(n15410) );
  NAND2_X1 U15462 ( .A1(n19370), .A2(n15409), .ZN(n12490) );
  NAND2_X1 U15463 ( .A1(n15410), .A2(n12490), .ZN(n15398) );
  NOR2_X1 U15464 ( .A1(n12491), .A2(n15393), .ZN(n15370) );
  INV_X1 U15465 ( .A(n15370), .ZN(n15388) );
  NAND2_X1 U15466 ( .A1(n19370), .A2(n15388), .ZN(n12492) );
  NAND2_X1 U15467 ( .A1(n12492), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12493) );
  OR2_X1 U15468 ( .A1(n15398), .A2(n12493), .ZN(n15371) );
  NAND2_X1 U15469 ( .A1(n15371), .A2(n15565), .ZN(n15361) );
  AND2_X1 U15470 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12505) );
  INV_X1 U15471 ( .A(n12505), .ZN(n12494) );
  NAND2_X1 U15472 ( .A1(n15565), .A2(n12494), .ZN(n12495) );
  NAND2_X1 U15473 ( .A1(n15361), .A2(n12495), .ZN(n15338) );
  AOI21_X1 U15474 ( .B1(n15310), .B2(n15565), .A(n15338), .ZN(n15312) );
  OAI21_X1 U15475 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15613), .A(
        n15312), .ZN(n12496) );
  NAND2_X1 U15476 ( .A1(n12496), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12497) );
  INV_X1 U15477 ( .A(n19129), .ZN(n19038) );
  NAND2_X1 U15478 ( .A1(n19038), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12528) );
  OAI211_X1 U15479 ( .C1(n16277), .C2(n16371), .A(n12497), .B(n12528), .ZN(
        n12507) );
  AOI21_X1 U15480 ( .B1(n15458), .B2(n13745), .A(n12498), .ZN(n13458) );
  NAND3_X1 U15481 ( .A1(n13458), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n19370), .ZN(n15617) );
  NAND2_X1 U15482 ( .A1(n15592), .A2(n12500), .ZN(n15497) );
  INV_X1 U15483 ( .A(n15411), .ZN(n12502) );
  NAND2_X1 U15484 ( .A1(n12502), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12503) );
  AND2_X1 U15485 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15370), .ZN(
        n12504) );
  NAND2_X1 U15486 ( .A1(n15366), .A2(n12505), .ZN(n15324) );
  XNOR2_X1 U15487 ( .A(n12538), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15319) );
  INV_X1 U15488 ( .A(n20044), .ZN(n15977) );
  OR2_X1 U15489 ( .A1(n20045), .A2(n15977), .ZN(n12509) );
  NAND2_X1 U15490 ( .A1(n12510), .A2(n12509), .ZN(n12511) );
  NAND2_X1 U15491 ( .A1(n12511), .A2(n19274), .ZN(n18958) );
  NOR2_X2 U15492 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20006) );
  NOR2_X1 U15493 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16422) );
  INV_X1 U15494 ( .A(n16422), .ZN(n12512) );
  NAND2_X1 U15495 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n14846) );
  OAI221_X4 U15496 ( .B1(n12512), .B2(n16421), .C1(n14846), .C2(n16421), .A(
        n19926), .ZN(n19754) );
  INV_X1 U15497 ( .A(n19376), .ZN(n19351) );
  NOR2_X1 U15498 ( .A1(n15315), .A2(n19376), .ZN(n12518) );
  INV_X1 U15499 ( .A(n20008), .ZN(n15625) );
  OR2_X1 U15500 ( .A1(n20006), .A2(n15625), .ZN(n20024) );
  NAND2_X1 U15501 ( .A1(n20024), .A2(n19926), .ZN(n12513) );
  NAND2_X1 U15502 ( .A1(n19926), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12940) );
  NAND2_X1 U15503 ( .A1(n19695), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12514) );
  NAND2_X1 U15504 ( .A1(n12940), .A2(n12514), .ZN(n12927) );
  NAND2_X1 U15505 ( .A1(n19038), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15307) );
  NAND2_X1 U15506 ( .A1(n19349), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12515) );
  OAI211_X1 U15507 ( .C1(n19359), .C2(n12516), .A(n15307), .B(n12515), .ZN(
        n12517) );
  NOR2_X1 U15508 ( .A1(n12518), .A2(n12517), .ZN(n12526) );
  NAND2_X1 U15509 ( .A1(n12519), .A2(n12541), .ZN(n12524) );
  INV_X1 U15510 ( .A(n12520), .ZN(n12522) );
  NAND2_X1 U15511 ( .A1(n12522), .A2(n12521), .ZN(n12523) );
  XNOR2_X1 U15512 ( .A(n12524), .B(n12523), .ZN(n15317) );
  NAND2_X1 U15513 ( .A1(n15317), .A2(n19355), .ZN(n12525) );
  OAI211_X1 U15514 ( .C1(n15319), .C2(n16325), .A(n12526), .B(n12525), .ZN(
        P2_U2984) );
  INV_X1 U15515 ( .A(n16279), .ZN(n12532) );
  NAND2_X1 U15516 ( .A1(n19349), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12527) );
  OAI211_X1 U15517 ( .C1(n19359), .C2(n12529), .A(n12528), .B(n12527), .ZN(
        n12530) );
  INV_X1 U15518 ( .A(n12530), .ZN(n12531) );
  OAI211_X1 U15519 ( .C1(n12536), .C2(n16325), .A(n12535), .B(n12534), .ZN(
        P2_U2983) );
  NAND2_X1 U15520 ( .A1(n12555), .A2(n19352), .ZN(n12554) );
  NAND2_X1 U15521 ( .A1(n12541), .A2(n12540), .ZN(n12543) );
  XOR2_X1 U15522 ( .A(n12543), .B(n12542), .Z(n12564) );
  NOR2_X1 U15523 ( .A1(n12568), .A2(n12544), .ZN(n12545) );
  INV_X1 U15524 ( .A(n14938), .ZN(n12550) );
  NOR2_X1 U15525 ( .A1(n19129), .A2(n19992), .ZN(n12559) );
  AOI21_X1 U15526 ( .B1(n19349), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n12559), .ZN(n12547) );
  OAI21_X1 U15527 ( .B1(n19359), .B2(n12548), .A(n12547), .ZN(n12549) );
  AOI21_X1 U15528 ( .B1(n12550), .B2(n19351), .A(n12549), .ZN(n12551) );
  INV_X1 U15529 ( .A(n12552), .ZN(n12553) );
  NAND2_X1 U15530 ( .A1(n12554), .A2(n12553), .ZN(P2_U2985) );
  NAND2_X1 U15531 ( .A1(n12555), .A2(n16361), .ZN(n12565) );
  NOR2_X1 U15532 ( .A1(n15324), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15342) );
  NOR2_X1 U15533 ( .A1(n15342), .A2(n15338), .ZN(n15330) );
  OAI21_X1 U15534 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15324), .A(
        n15330), .ZN(n12563) );
  AOI21_X1 U15535 ( .B1(n12557), .B2(n14867), .A(n10236), .ZN(n12558) );
  OR4_X1 U15536 ( .A1(n15329), .A2(n15323), .A3(n15324), .A4(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12561) );
  INV_X1 U15537 ( .A(n12559), .ZN(n12560) );
  OAI211_X1 U15538 ( .C1(n15033), .C2(n16371), .A(n12561), .B(n12560), .ZN(
        n12562) );
  OAI21_X1 U15539 ( .B1(n12566), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12537), .ZN(n15320) );
  INV_X1 U15540 ( .A(n12567), .ZN(n12570) );
  INV_X1 U15541 ( .A(n12603), .ZN(n12569) );
  AOI21_X1 U15542 ( .B1(n12570), .B2(n12569), .A(n12568), .ZN(n15327) );
  NAND2_X1 U15543 ( .A1(n19038), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15321) );
  NAND2_X1 U15544 ( .A1(n19349), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12571) );
  OAI211_X1 U15545 ( .C1(n19359), .C2(n12572), .A(n15321), .B(n12571), .ZN(
        n12573) );
  AOI21_X1 U15546 ( .B1(n15327), .B2(n19351), .A(n12573), .ZN(n12581) );
  XOR2_X1 U15547 ( .A(n12575), .B(n12577), .Z(n15103) );
  INV_X1 U15548 ( .A(n12575), .ZN(n12576) );
  OAI22_X1 U15549 ( .A1(n15103), .A2(n15323), .B1(n12577), .B2(n12576), .ZN(
        n12580) );
  XNOR2_X1 U15550 ( .A(n12578), .B(n15329), .ZN(n12579) );
  INV_X1 U15551 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20043) );
  NOR2_X1 U15552 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(n20043), .ZN(n12583) );
  NOR4_X1 U15553 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12582) );
  INV_X1 U15554 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20998) );
  NAND4_X1 U15555 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n12583), .A3(n12582), .A4(
        n20998), .ZN(n12596) );
  NOR2_X1 U15556 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12596), .ZN(n16597)
         );
  INV_X1 U15557 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20947) );
  NOR3_X1 U15558 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20947), .ZN(n12585) );
  NOR4_X1 U15559 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12584) );
  NAND4_X1 U15560 ( .A1(n20241), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12585), .A4(
        n12584), .ZN(U214) );
  NOR4_X1 U15561 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12589) );
  NOR4_X1 U15562 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12588) );
  NOR4_X1 U15563 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12587) );
  NOR4_X1 U15564 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12586) );
  NAND4_X1 U15565 ( .A1(n12589), .A2(n12588), .A3(n12587), .A4(n12586), .ZN(
        n12594) );
  NOR4_X1 U15566 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12592) );
  NOR4_X1 U15567 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12591) );
  NOR4_X1 U15568 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12590) );
  INV_X1 U15569 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19954) );
  NAND4_X1 U15570 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n19954), .ZN(
        n12593) );
  OAI21_X1 U15571 ( .B1(n12594), .B2(n12593), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12595) );
  NOR2_X1 U15572 ( .A1(n19375), .A2(n12596), .ZN(n16512) );
  NAND2_X1 U15573 ( .A1(n16512), .A2(U214), .ZN(U212) );
  INV_X1 U15574 ( .A(n12597), .ZN(n12598) );
  AOI211_X1 U15575 ( .C1(n15107), .C2(n12599), .A(n12598), .B(n19929), .ZN(
        n12612) );
  OAI22_X1 U15576 ( .A1(n15105), .A2(n19097), .B1(n19989), .B2(n19188), .ZN(
        n12611) );
  INV_X1 U15577 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12600) );
  OAI22_X1 U15578 ( .A1(n12601), .A2(n19194), .B1(n12600), .B2(n19156), .ZN(
        n12610) );
  AND2_X1 U15579 ( .A1(n14953), .A2(n12602), .ZN(n12604) );
  OR2_X1 U15580 ( .A1(n12604), .A2(n12603), .ZN(n15340) );
  OR2_X1 U15581 ( .A1(n12606), .A2(n12607), .ZN(n12608) );
  NAND2_X1 U15582 ( .A1(n12605), .A2(n12608), .ZN(n15336) );
  OAI22_X1 U15583 ( .A1(n15340), .A2(n19174), .B1(n15336), .B2(n19154), .ZN(
        n12609) );
  OR4_X1 U15584 ( .A1(n12612), .A2(n12611), .A3(n12610), .A4(n12609), .ZN(
        P2_U2828) );
  INV_X1 U15585 ( .A(n12704), .ZN(n19275) );
  AND2_X1 U15586 ( .A1(n12613), .A2(n19275), .ZN(n19196) );
  INV_X1 U15587 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12614) );
  INV_X1 U15588 ( .A(n12615), .ZN(n18950) );
  OAI211_X1 U15589 ( .C1(n19196), .C2(n12614), .A(n12618), .B(n18950), .ZN(
        P2_U2814) );
  INV_X1 U15590 ( .A(n18952), .ZN(n14848) );
  OAI21_X1 U15591 ( .B1(n12615), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n14848), 
        .ZN(n12616) );
  OAI21_X1 U15592 ( .B1(n14843), .B2(n14848), .A(n12616), .ZN(P2_U3612) );
  INV_X1 U15593 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19324) );
  NAND2_X1 U15594 ( .A1(n10598), .A2(n19924), .ZN(n12617) );
  OR2_X1 U15595 ( .A1(n12618), .A2(n12617), .ZN(n12638) );
  INV_X1 U15596 ( .A(n12638), .ZN(n12672) );
  MUX2_X1 U15597 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n19375), .Z(n19229) );
  NAND2_X1 U15598 ( .A1(n12672), .A2(n19229), .ZN(n12629) );
  INV_X1 U15599 ( .A(n12618), .ZN(n12619) );
  OAI21_X1 U15600 ( .B1(n10406), .B2(n19924), .A(n12619), .ZN(n12634) );
  NAND2_X1 U15601 ( .A1(n12634), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12620) );
  OAI211_X1 U15602 ( .C1(n19324), .C2(n19276), .A(n12629), .B(n12620), .ZN(
        P2_U2977) );
  INV_X1 U15603 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19287) );
  MUX2_X1 U15604 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n19375), .Z(n19224) );
  NAND2_X1 U15605 ( .A1(n12672), .A2(n19224), .ZN(n12627) );
  NAND2_X1 U15606 ( .A1(n12634), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12621) );
  OAI211_X1 U15607 ( .C1(n19287), .C2(n19276), .A(n12627), .B(n12621), .ZN(
        P2_U2964) );
  INV_X1 U15608 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19316) );
  MUX2_X1 U15609 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n19375), .Z(n19219) );
  NAND2_X1 U15610 ( .A1(n12672), .A2(n19219), .ZN(n12631) );
  NAND2_X1 U15611 ( .A1(n12634), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12622) );
  OAI211_X1 U15612 ( .C1(n19316), .C2(n19276), .A(n12631), .B(n12622), .ZN(
        P2_U2981) );
  INV_X1 U15613 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20965) );
  NAND2_X1 U15614 ( .A1(n19375), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12624) );
  INV_X1 U15615 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16551) );
  OR2_X1 U15616 ( .A1(n19375), .A2(n16551), .ZN(n12623) );
  NAND2_X1 U15617 ( .A1(n12624), .A2(n12623), .ZN(n19234) );
  NAND2_X1 U15618 ( .A1(n12672), .A2(n19234), .ZN(n12633) );
  NAND2_X1 U15619 ( .A1(n12634), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12625) );
  OAI211_X1 U15620 ( .C1(n20965), .C2(n19276), .A(n12633), .B(n12625), .ZN(
        P2_U2975) );
  INV_X1 U15621 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19320) );
  NAND2_X1 U15622 ( .A1(n12634), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12626) );
  OAI211_X1 U15623 ( .C1(n19320), .C2(n19276), .A(n12627), .B(n12626), .ZN(
        P2_U2979) );
  INV_X1 U15624 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19291) );
  NAND2_X1 U15625 ( .A1(n12634), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12628) );
  OAI211_X1 U15626 ( .C1(n19291), .C2(n19276), .A(n12629), .B(n12628), .ZN(
        P2_U2962) );
  INV_X1 U15627 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n19283) );
  NAND2_X1 U15628 ( .A1(n12634), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12630) );
  OAI211_X1 U15629 ( .C1(n19283), .C2(n19276), .A(n12631), .B(n12630), .ZN(
        P2_U2966) );
  INV_X1 U15630 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19295) );
  NAND2_X1 U15631 ( .A1(n12634), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12632) );
  OAI211_X1 U15632 ( .C1(n19295), .C2(n19276), .A(n12633), .B(n12632), .ZN(
        P2_U2960) );
  OAI22_X1 U15633 ( .A1(n19375), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19377), .ZN(n19385) );
  INV_X1 U15634 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12635) );
  INV_X1 U15635 ( .A(n12634), .ZN(n12643) );
  INV_X1 U15636 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19312) );
  OAI222_X1 U15637 ( .A1(n12638), .A2(n19385), .B1(n12635), .B2(n12643), .C1(
        n19276), .C2(n19312), .ZN(P2_U2952) );
  INV_X1 U15638 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12637) );
  INV_X1 U15639 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U15640 ( .A1(n19377), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19375), .ZN(n19217) );
  OAI222_X1 U15641 ( .A1(n19276), .A2(n12637), .B1(n12636), .B2(n12643), .C1(
        n12638), .C2(n19217), .ZN(P2_U2982) );
  INV_X1 U15642 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12640) );
  INV_X1 U15643 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12639) );
  OAI222_X1 U15644 ( .A1(n12640), .A2(n19276), .B1(n12639), .B2(n12643), .C1(
        n12638), .C2(n19385), .ZN(P2_U2967) );
  INV_X1 U15645 ( .A(n12643), .ZN(n12678) );
  AOI22_X1 U15646 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12641) );
  AOI22_X1 U15647 ( .A1(n19377), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19375), .ZN(n19412) );
  INV_X1 U15648 ( .A(n19412), .ZN(n15073) );
  NAND2_X1 U15649 ( .A1(n12672), .A2(n15073), .ZN(n12644) );
  NAND2_X1 U15650 ( .A1(n12641), .A2(n12644), .ZN(P2_U2958) );
  AOI22_X1 U15651 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U15652 ( .A1(n19377), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19375), .ZN(n19392) );
  INV_X1 U15653 ( .A(n19392), .ZN(n15097) );
  NAND2_X1 U15654 ( .A1(n12672), .A2(n15097), .ZN(n12664) );
  NAND2_X1 U15655 ( .A1(n12642), .A2(n12664), .ZN(P2_U2968) );
  AOI22_X1 U15656 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n12634), .B1(n12683), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12645) );
  NAND2_X1 U15657 ( .A1(n12645), .A2(n12644), .ZN(P2_U2973) );
  AOI22_X1 U15658 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n12634), .B1(n12683), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12649) );
  INV_X1 U15659 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n12646) );
  OR2_X1 U15660 ( .A1(n19375), .A2(n12646), .ZN(n12648) );
  NAND2_X1 U15661 ( .A1(n19375), .A2(BUF2_REG_7__SCAN_IN), .ZN(n12647) );
  AND2_X1 U15662 ( .A1(n12648), .A2(n12647), .ZN(n19424) );
  INV_X1 U15663 ( .A(n19424), .ZN(n15067) );
  NAND2_X1 U15664 ( .A1(n12672), .A2(n15067), .ZN(n12659) );
  NAND2_X1 U15665 ( .A1(n12649), .A2(n12659), .ZN(P2_U2974) );
  AOI22_X1 U15666 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15667 ( .A1(n19377), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19375), .ZN(n19398) );
  INV_X1 U15668 ( .A(n19398), .ZN(n15087) );
  NAND2_X1 U15669 ( .A1(n12672), .A2(n15087), .ZN(n12681) );
  NAND2_X1 U15670 ( .A1(n12650), .A2(n12681), .ZN(P2_U2955) );
  AOI22_X1 U15671 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12651) );
  INV_X1 U15672 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16556) );
  INV_X1 U15673 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18296) );
  OAI22_X1 U15674 ( .A1(n19375), .A2(n16556), .B1(n18296), .B2(n19377), .ZN(
        n19407) );
  NAND2_X1 U15675 ( .A1(n12672), .A2(n19407), .ZN(n12653) );
  NAND2_X1 U15676 ( .A1(n12651), .A2(n12653), .ZN(P2_U2972) );
  AOI22_X1 U15677 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12652) );
  OAI22_X1 U15678 ( .A1(n19375), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19377), .ZN(n19395) );
  INV_X1 U15679 ( .A(n19395), .ZN(n16317) );
  NAND2_X1 U15680 ( .A1(n12672), .A2(n16317), .ZN(n12684) );
  NAND2_X1 U15681 ( .A1(n12652), .A2(n12684), .ZN(P2_U2969) );
  AOI22_X1 U15682 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U15683 ( .A1(n12654), .A2(n12653), .ZN(P2_U2957) );
  AOI22_X1 U15684 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12658) );
  INV_X1 U15685 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14313) );
  OR2_X1 U15686 ( .A1(n19375), .A2(n14313), .ZN(n12656) );
  NAND2_X1 U15687 ( .A1(n19375), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12655) );
  AND2_X1 U15688 ( .A1(n12656), .A2(n12655), .ZN(n19222) );
  INV_X1 U15689 ( .A(n19222), .ZN(n12657) );
  NAND2_X1 U15690 ( .A1(n12672), .A2(n12657), .ZN(n12679) );
  NAND2_X1 U15691 ( .A1(n12658), .A2(n12679), .ZN(P2_U2980) );
  AOI22_X1 U15692 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12660) );
  NAND2_X1 U15693 ( .A1(n12660), .A2(n12659), .ZN(P2_U2959) );
  AOI22_X1 U15694 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12663) );
  INV_X1 U15695 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13622) );
  OR2_X1 U15696 ( .A1(n19375), .A2(n13622), .ZN(n12662) );
  NAND2_X1 U15697 ( .A1(n19375), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12661) );
  AND2_X1 U15698 ( .A1(n12662), .A2(n12661), .ZN(n19232) );
  INV_X1 U15699 ( .A(n19232), .ZN(n15053) );
  NAND2_X1 U15700 ( .A1(n12672), .A2(n15053), .ZN(n12667) );
  NAND2_X1 U15701 ( .A1(n12663), .A2(n12667), .ZN(P2_U2961) );
  AOI22_X1 U15702 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12665) );
  NAND2_X1 U15703 ( .A1(n12665), .A2(n12664), .ZN(P2_U2953) );
  AOI22_X1 U15704 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12666) );
  OAI22_X1 U15705 ( .A1(n19375), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19377), .ZN(n19402) );
  INV_X1 U15706 ( .A(n19402), .ZN(n16312) );
  NAND2_X1 U15707 ( .A1(n12672), .A2(n16312), .ZN(n12674) );
  NAND2_X1 U15708 ( .A1(n12666), .A2(n12674), .ZN(P2_U2971) );
  AOI22_X1 U15709 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U15710 ( .A1(n12668), .A2(n12667), .ZN(P2_U2976) );
  AOI22_X1 U15711 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12673) );
  INV_X1 U15712 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14324) );
  OR2_X1 U15713 ( .A1(n19375), .A2(n14324), .ZN(n12670) );
  NAND2_X1 U15714 ( .A1(n19375), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12669) );
  AND2_X1 U15715 ( .A1(n12670), .A2(n12669), .ZN(n19227) );
  INV_X1 U15716 ( .A(n19227), .ZN(n12671) );
  NAND2_X1 U15717 ( .A1(n12672), .A2(n12671), .ZN(n12676) );
  NAND2_X1 U15718 ( .A1(n12673), .A2(n12676), .ZN(P2_U2978) );
  AOI22_X1 U15719 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12675) );
  NAND2_X1 U15720 ( .A1(n12675), .A2(n12674), .ZN(P2_U2956) );
  AOI22_X1 U15721 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12677) );
  NAND2_X1 U15722 ( .A1(n12677), .A2(n12676), .ZN(P2_U2963) );
  AOI22_X1 U15723 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12680) );
  NAND2_X1 U15724 ( .A1(n12680), .A2(n12679), .ZN(P2_U2965) );
  AOI22_X1 U15725 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12682) );
  NAND2_X1 U15726 ( .A1(n12682), .A2(n12681), .ZN(P2_U2970) );
  AOI22_X1 U15727 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n12678), .B1(n12683), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U15728 ( .A1(n12685), .A2(n12684), .ZN(P2_U2954) );
  NAND2_X1 U15729 ( .A1(n19411), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15730 ( .A1(n12938), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20006), .B2(n20042), .ZN(n12687) );
  NAND2_X1 U15731 ( .A1(n10598), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12688) );
  AND4_X1 U15732 ( .A1(n10412), .A2(n12688), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19632), .ZN(n12689) );
  INV_X1 U15733 ( .A(n16394), .ZN(n12690) );
  INV_X1 U15734 ( .A(n13061), .ZN(n16390) );
  NAND2_X1 U15735 ( .A1(n12690), .A2(n16390), .ZN(n12698) );
  INV_X1 U15736 ( .A(n12691), .ZN(n13053) );
  NAND2_X1 U15737 ( .A1(n12698), .A2(n13053), .ZN(n12692) );
  MUX2_X1 U15738 ( .A(n15624), .B(n12693), .S(n15004), .Z(n12694) );
  OAI21_X1 U15739 ( .B1(n20037), .B2(n15025), .A(n12694), .ZN(P2_U2887) );
  INV_X1 U15740 ( .A(n16393), .ZN(n12696) );
  AND2_X1 U15741 ( .A1(n12466), .A2(n19924), .ZN(n16386) );
  AND3_X1 U15742 ( .A1(n16384), .A2(n16386), .A3(n10578), .ZN(n12695) );
  AOI21_X1 U15743 ( .B1(n16394), .B2(n12696), .A(n12695), .ZN(n12708) );
  NAND3_X1 U15744 ( .A1(n12708), .A2(n12698), .A3(n12697), .ZN(n12701) );
  NAND2_X1 U15745 ( .A1(n19275), .A2(n16385), .ZN(n12699) );
  NOR2_X1 U15746 ( .A1(n19278), .A2(n12699), .ZN(n12700) );
  INV_X1 U15747 ( .A(n16402), .ZN(n16381) );
  NOR2_X1 U15748 ( .A1(n19926), .A2(n14846), .ZN(n16429) );
  AOI22_X1 U15749 ( .A1(n16429), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n19926), .ZN(n12702) );
  OAI21_X1 U15750 ( .B1(n16381), .B2(n18956), .A(n12702), .ZN(n15644) );
  INV_X1 U15751 ( .A(n15644), .ZN(n13725) );
  OR3_X1 U15752 ( .A1(n12704), .A2(n12703), .A3(n10598), .ZN(n16387) );
  OR3_X1 U15753 ( .A1(n13725), .A2(n20008), .A3(n16387), .ZN(n12705) );
  OAI21_X1 U15754 ( .B1(n16397), .B2(n15644), .A(n12705), .ZN(P2_U3595) );
  INV_X1 U15755 ( .A(n10418), .ZN(n12706) );
  NAND2_X1 U15756 ( .A1(n10224), .A2(n12706), .ZN(n12707) );
  NAND2_X1 U15757 ( .A1(n12708), .A2(n12707), .ZN(n12709) );
  NAND2_X1 U15758 ( .A1(n19239), .A2(n12711), .ZN(n19215) );
  AOI21_X1 U15759 ( .B1(n20037), .B2(n19269), .A(n19265), .ZN(n12721) );
  INV_X1 U15760 ( .A(n12712), .ZN(n12713) );
  XNOR2_X1 U15761 ( .A(n12714), .B(n12713), .ZN(n19184) );
  INV_X1 U15762 ( .A(n19184), .ZN(n12720) );
  NOR3_X1 U15763 ( .A1(n20037), .A2(n19184), .A3(n19216), .ZN(n12715) );
  AOI21_X1 U15764 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n19264), .A(n12715), .ZN(
        n12719) );
  AND2_X1 U15765 ( .A1(n19422), .A2(n19411), .ZN(n12717) );
  INV_X1 U15766 ( .A(n19385), .ZN(n19206) );
  NAND2_X1 U15767 ( .A1(n19241), .A2(n19206), .ZN(n12718) );
  OAI211_X1 U15768 ( .C1(n12721), .C2(n12720), .A(n12719), .B(n12718), .ZN(
        P2_U2919) );
  NAND2_X1 U15769 ( .A1(n12722), .A2(n12873), .ZN(n12864) );
  NOR2_X2 U15770 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20797) );
  NAND2_X1 U15771 ( .A1(n20797), .A2(n20867), .ZN(n20060) );
  INV_X1 U15772 ( .A(n20060), .ZN(n12859) );
  INV_X1 U15773 ( .A(n12857), .ZN(n13088) );
  AOI211_X1 U15774 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n12858), .A(n12859), 
        .B(n13088), .ZN(n12724) );
  INV_X1 U15775 ( .A(n12724), .ZN(P1_U2801) );
  NOR2_X1 U15776 ( .A1(n13008), .A2(n12725), .ZN(n12886) );
  INV_X1 U15777 ( .A(n12940), .ZN(n12727) );
  NAND2_X1 U15778 ( .A1(n12728), .A2(n12727), .ZN(n12730) );
  XNOR2_X1 U15779 ( .A(n20033), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19513) );
  AND2_X1 U15780 ( .A1(n19513), .A2(n20006), .ZN(n19690) );
  AOI21_X1 U15781 ( .B1(n12938), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19690), .ZN(n12729) );
  NAND2_X1 U15782 ( .A1(n12730), .A2(n12729), .ZN(n12731) );
  NAND2_X1 U15783 ( .A1(n12732), .A2(n12731), .ZN(n12733) );
  MUX2_X1 U15784 ( .A(n12734), .B(n19175), .S(n14998), .Z(n12735) );
  OAI21_X1 U15785 ( .B1(n20026), .B2(n15025), .A(n12735), .ZN(P2_U2886) );
  INV_X1 U15786 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17291) );
  NAND2_X1 U15787 ( .A1(n18905), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18775) );
  AOI22_X1 U15788 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12739) );
  INV_X1 U15789 ( .A(n15795), .ZN(n12827) );
  AOI22_X1 U15790 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12738) );
  INV_X1 U15791 ( .A(n12816), .ZN(n15701) );
  INV_X2 U15792 ( .A(n15701), .ZN(n17270) );
  NOR2_X2 U15793 ( .A1(n12740), .A2(n12743), .ZN(n12839) );
  AOI22_X1 U15794 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12737) );
  NOR3_X2 U15795 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18883), .A3(
        n18731), .ZN(n12752) );
  AOI22_X1 U15796 ( .A1(n17264), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12736) );
  NAND4_X1 U15797 ( .A1(n12739), .A2(n12738), .A3(n12737), .A4(n12736), .ZN(
        n12751) );
  AOI22_X1 U15798 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12749) );
  INV_X2 U15799 ( .A(n10212), .ZN(n15834) );
  AOI22_X1 U15800 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9650), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U15801 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U15802 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12746) );
  NAND4_X1 U15803 ( .A1(n12749), .A2(n12748), .A3(n12747), .A4(n12746), .ZN(
        n12750) );
  AOI22_X1 U15804 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U15805 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15806 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12754) );
  BUF_X4 U15807 ( .A(n12752), .Z(n17264) );
  AOI22_X1 U15808 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12753) );
  NAND4_X1 U15809 ( .A1(n12756), .A2(n12755), .A3(n12754), .A4(n12753), .ZN(
        n12762) );
  INV_X2 U15810 ( .A(n9706), .ZN(n17035) );
  AOI22_X1 U15811 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U15812 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U15813 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9645), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U15814 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12757) );
  NAND4_X1 U15815 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12761) );
  OAI22_X1 U15816 ( .A1(n18891), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U15817 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18539), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18901), .ZN(n13691) );
  OAI21_X1 U15818 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18891), .A(
        n12764), .ZN(n12765) );
  OAI22_X1 U15819 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18755), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12765), .ZN(n12771) );
  NOR2_X1 U15820 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18755), .ZN(
        n12766) );
  NAND2_X1 U15821 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12765), .ZN(
        n12770) );
  AOI22_X1 U15822 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12771), .B1(
        n12766), .B2(n12770), .ZN(n12774) );
  AOI21_X1 U15823 ( .B1(n18909), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n13690), .ZN(n15893) );
  AND2_X1 U15824 ( .A1(n13691), .A2(n15893), .ZN(n12773) );
  OAI21_X1 U15825 ( .B1(n12769), .B2(n12768), .A(n12774), .ZN(n12767) );
  INV_X1 U15826 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18721) );
  OAI22_X1 U15827 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18721), .B1(
        n12772), .B2(n12771), .ZN(n13692) );
  AOI211_X1 U15828 ( .C1(n12774), .C2(n12773), .A(n15894), .B(n13692), .ZN(
        n16432) );
  INV_X1 U15829 ( .A(n16432), .ZN(n18717) );
  AOI22_X1 U15830 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U15831 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9645), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12783) );
  INV_X1 U15832 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U15833 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12775) );
  OAI21_X1 U15834 ( .B1(n10230), .B2(n17152), .A(n12775), .ZN(n12781) );
  AOI22_X1 U15835 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U15836 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U15837 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U15838 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12776) );
  NAND4_X1 U15839 ( .A1(n12779), .A2(n12778), .A3(n12777), .A4(n12776), .ZN(
        n12780) );
  AOI22_X1 U15840 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12794) );
  AOI22_X1 U15841 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12793) );
  INV_X1 U15842 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U15843 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12785) );
  OAI21_X1 U15844 ( .B1(n15701), .B2(n17280), .A(n12785), .ZN(n12791) );
  AOI22_X1 U15845 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12789) );
  AOI22_X1 U15846 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U15847 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U15848 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12786) );
  NAND4_X1 U15849 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12790) );
  AOI22_X1 U15850 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U15851 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U15852 ( .A1(n15814), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12795) );
  OAI21_X1 U15853 ( .B1(n12827), .B2(n21083), .A(n12795), .ZN(n12801) );
  AOI22_X1 U15854 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U15855 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12798) );
  AOI22_X1 U15856 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9648), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12797) );
  AOI22_X1 U15857 ( .A1(n17264), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12796) );
  NAND4_X1 U15858 ( .A1(n12799), .A2(n12798), .A3(n12797), .A4(n12796), .ZN(
        n12800) );
  AOI211_X1 U15859 ( .C1(n17247), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n12801), .B(n12800), .ZN(n12802) );
  NAND3_X1 U15860 ( .A1(n12804), .A2(n12803), .A3(n12802), .ZN(n13683) );
  AOI22_X1 U15861 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U15862 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U15863 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U15864 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12805) );
  NAND4_X1 U15865 ( .A1(n12808), .A2(n12807), .A3(n12806), .A4(n12805), .ZN(
        n12814) );
  AOI22_X1 U15866 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U15867 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U15868 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12810) );
  AOI22_X1 U15869 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12809) );
  NAND4_X1 U15870 ( .A1(n12812), .A2(n12811), .A3(n12810), .A4(n12809), .ZN(
        n12813) );
  AOI22_X1 U15871 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U15872 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12824) );
  AOI22_X1 U15873 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12815) );
  OAI21_X1 U15874 ( .B1(n15648), .B2(n20994), .A(n12815), .ZN(n12822) );
  AOI22_X1 U15875 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U15876 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U15877 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U15878 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12817) );
  NAND4_X1 U15879 ( .A1(n12820), .A2(n12819), .A3(n12818), .A4(n12817), .ZN(
        n12821) );
  NOR2_X1 U15880 ( .A1(n18293), .A2(n17317), .ZN(n18726) );
  AOI22_X1 U15881 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U15882 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12835) );
  INV_X1 U15883 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15816) );
  AOI22_X1 U15884 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12826) );
  OAI21_X1 U15885 ( .B1(n9706), .B2(n15816), .A(n12826), .ZN(n12833) );
  AOI22_X1 U15886 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U15887 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9650), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12830) );
  AOI22_X1 U15888 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12829) );
  INV_X2 U15889 ( .A(n12827), .ZN(n17262) );
  AOI22_X1 U15890 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12828) );
  NAND4_X1 U15891 ( .A1(n12831), .A2(n12830), .A3(n12829), .A4(n12828), .ZN(
        n12832) );
  AOI211_X1 U15892 ( .C1(n17247), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n12833), .B(n12832), .ZN(n12834) );
  NAND3_X1 U15893 ( .A1(n12836), .A2(n12835), .A3(n12834), .ZN(n13673) );
  NAND3_X1 U15894 ( .A1(n13686), .A2(n18726), .A3(n13673), .ZN(n15741) );
  NOR2_X1 U15895 ( .A1(n18301), .A2(n13673), .ZN(n13697) );
  NOR2_X1 U15896 ( .A1(n15864), .A2(n13683), .ZN(n18725) );
  NAND2_X1 U15897 ( .A1(n13697), .A2(n18725), .ZN(n13684) );
  NAND2_X1 U15898 ( .A1(n18307), .A2(n18293), .ZN(n12837) );
  NAND2_X1 U15899 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .ZN(n17296) );
  INV_X1 U15900 ( .A(n17296), .ZN(n17301) );
  NAND4_X1 U15901 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n17290), .ZN(n17148) );
  AOI21_X1 U15902 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17278), .A(n17311), .ZN(
        n17259) );
  AOI22_X1 U15903 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U15904 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9645), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U15905 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12839), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12840) );
  OAI21_X1 U15906 ( .B1(n12841), .B2(n17152), .A(n12840), .ZN(n12849) );
  AOI22_X1 U15907 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U15908 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U15909 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U15910 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12844) );
  NAND4_X1 U15911 ( .A1(n12847), .A2(n12846), .A3(n12845), .A4(n12844), .ZN(
        n12848) );
  AOI211_X1 U15912 ( .C1(n9649), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n12849), .B(n12848), .ZN(n12850) );
  NAND3_X1 U15913 ( .A1(n12852), .A2(n12851), .A3(n12850), .ZN(n17425) );
  AOI22_X1 U15914 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17259), .B1(n17311), 
        .B2(n17425), .ZN(n12856) );
  INV_X1 U15915 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n12854) );
  AND2_X1 U15916 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17278), .ZN(n12853) );
  NAND3_X1 U15917 ( .A1(n18307), .A2(n12854), .A3(n12853), .ZN(n12855) );
  NAND2_X1 U15918 ( .A1(n12856), .A2(n12855), .ZN(P3_U2693) );
  NOR2_X1 U15919 ( .A1(n12859), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n12862)
         );
  NAND2_X1 U15920 ( .A1(n20949), .A2(n12860), .ZN(n12861) );
  OAI21_X1 U15921 ( .B1(n20949), .B2(n12862), .A(n12861), .ZN(P1_U3487) );
  INV_X1 U15922 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12879) );
  AND2_X1 U15923 ( .A1(n13231), .A2(n13343), .ZN(n12863) );
  AOI21_X1 U15924 ( .B1(n12864), .B2(n12723), .A(n12863), .ZN(n20056) );
  INV_X2 U15925 ( .A(n14043), .ZN(n13022) );
  NOR2_X1 U15926 ( .A1(n12865), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15973) );
  INV_X1 U15927 ( .A(n15973), .ZN(n13351) );
  NAND3_X1 U15928 ( .A1(n13343), .A2(n13022), .A3(n13351), .ZN(n12866) );
  NAND2_X1 U15929 ( .A1(n12866), .A2(n20951), .ZN(n20952) );
  AND2_X1 U15930 ( .A1(n20056), .A2(n20952), .ZN(n15944) );
  NOR2_X1 U15931 ( .A1(n15944), .A2(n20057), .ZN(n20065) );
  NAND2_X1 U15932 ( .A1(n12867), .A2(n13343), .ZN(n12868) );
  NAND2_X1 U15933 ( .A1(n13035), .A2(n12868), .ZN(n13237) );
  NAND3_X1 U15934 ( .A1(n12869), .A2(n13029), .A3(n20246), .ZN(n12870) );
  NAND2_X1 U15935 ( .A1(n13237), .A2(n12870), .ZN(n12872) );
  NAND2_X1 U15936 ( .A1(n11046), .A2(n20262), .ZN(n13229) );
  NOR2_X1 U15937 ( .A1(n12871), .A2(n13229), .ZN(n13245) );
  MUX2_X1 U15938 ( .A(n12872), .B(n13245), .S(n13224), .Z(n12876) );
  INV_X1 U15939 ( .A(n12722), .ZN(n12874) );
  NOR2_X1 U15940 ( .A1(n12874), .A2(n12873), .ZN(n12875) );
  OAI21_X1 U15941 ( .B1(n12876), .B2(n12875), .A(n20292), .ZN(n15946) );
  INV_X1 U15942 ( .A(n15946), .ZN(n12877) );
  NAND2_X1 U15943 ( .A1(n12877), .A2(n20065), .ZN(n12878) );
  OAI21_X1 U15944 ( .B1(n12879), .B2(n20065), .A(n12878), .ZN(P1_U3484) );
  OAI21_X1 U15945 ( .B1(n12881), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12880), .ZN(n12924) );
  XNOR2_X1 U15946 ( .A(n19193), .B(n13721), .ZN(n12922) );
  OAI22_X1 U15947 ( .A1(n12924), .A2(n19366), .B1(n15597), .B2(n12922), .ZN(
        n12884) );
  AOI22_X1 U15948 ( .A1(n19364), .A2(n19184), .B1(n19362), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12882) );
  NAND2_X1 U15949 ( .A1(n19038), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12923) );
  OAI211_X1 U15950 ( .C1(n15589), .C2(n15624), .A(n12882), .B(n12923), .ZN(
        n12883) );
  AOI211_X1 U15951 ( .C1(n13721), .C2(n19370), .A(n12884), .B(n12883), .ZN(
        n12885) );
  INV_X1 U15952 ( .A(n12885), .ZN(P2_U3046) );
  INV_X1 U15953 ( .A(n20006), .ZN(n19819) );
  NOR2_X1 U15954 ( .A1(n20023), .A2(n20033), .ZN(n19858) );
  INV_X1 U15955 ( .A(n12935), .ZN(n12890) );
  NAND2_X1 U15956 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19722) );
  NAND2_X1 U15957 ( .A1(n19722), .A2(n20023), .ZN(n12889) );
  NAND2_X1 U15958 ( .A1(n12890), .A2(n12889), .ZN(n19514) );
  NOR2_X1 U15959 ( .A1(n19819), .A2(n19514), .ZN(n12891) );
  AOI21_X1 U15960 ( .B1(n12938), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12891), .ZN(n12892) );
  NAND2_X1 U15961 ( .A1(n13924), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12931) );
  INV_X1 U15962 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13574) );
  MUX2_X1 U15963 ( .A(n13574), .B(n15636), .S(n14998), .Z(n12895) );
  OAI21_X1 U15964 ( .B1(n20019), .B2(n15025), .A(n12895), .ZN(P2_U2885) );
  AND2_X1 U15965 ( .A1(n12722), .A2(n20262), .ZN(n14823) );
  NAND2_X1 U15966 ( .A1(n14823), .A2(n15973), .ZN(n12981) );
  NAND2_X1 U15967 ( .A1(n13352), .A2(n15973), .ZN(n12896) );
  NOR2_X1 U15968 ( .A1(n12723), .A2(n12896), .ZN(n15955) );
  INV_X1 U15969 ( .A(n15955), .ZN(n12897) );
  NAND2_X1 U15970 ( .A1(n12981), .A2(n12897), .ZN(n12899) );
  INV_X1 U15971 ( .A(n13036), .ZN(n12898) );
  NAND2_X1 U15972 ( .A1(n20167), .A2(n20246), .ZN(n13145) );
  NOR2_X1 U15973 ( .A1(n20870), .A2(n20867), .ZN(n16262) );
  NAND2_X1 U15974 ( .A1(n20868), .A2(n16262), .ZN(n20165) );
  INV_X2 U15975 ( .A(n20165), .ZN(n20185) );
  NOR2_X4 U15976 ( .A1(n20167), .A2(n20185), .ZN(n20184) );
  AOI22_X1 U15977 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12900) );
  OAI21_X1 U15978 ( .B1(n14330), .B2(n13145), .A(n12900), .ZN(P1_U2910) );
  AOI22_X1 U15979 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12901) );
  OAI21_X1 U15980 ( .B1(n14326), .B2(n13145), .A(n12901), .ZN(P1_U2909) );
  INV_X1 U15981 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U15982 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12902) );
  OAI21_X1 U15983 ( .B1(n12903), .B2(n13145), .A(n12902), .ZN(P1_U2907) );
  INV_X1 U15984 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U15985 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12904) );
  OAI21_X1 U15986 ( .B1(n12905), .B2(n13145), .A(n12904), .ZN(P1_U2912) );
  AOI22_X1 U15987 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12906) );
  OAI21_X1 U15988 ( .B1(n14309), .B2(n13145), .A(n12906), .ZN(P1_U2906) );
  INV_X1 U15989 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U15990 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12907) );
  OAI21_X1 U15991 ( .B1(n12908), .B2(n13145), .A(n12907), .ZN(P1_U2908) );
  INV_X1 U15992 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U15993 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12909) );
  OAI21_X1 U15994 ( .B1(n12910), .B2(n13145), .A(n12909), .ZN(P1_U2911) );
  AOI21_X1 U15995 ( .B1(n12913), .B2(n12912), .A(n12911), .ZN(n12914) );
  XOR2_X1 U15996 ( .A(n12914), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n19360) );
  NOR2_X1 U15997 ( .A1(n19129), .A2(n10428), .ZN(n19363) );
  OAI21_X1 U15998 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12916), .A(
        n12915), .ZN(n19367) );
  NOR2_X1 U15999 ( .A1(n16325), .A2(n19367), .ZN(n12917) );
  AOI211_X1 U16000 ( .C1(n19360), .C2(n19355), .A(n19363), .B(n12917), .ZN(
        n12921) );
  INV_X1 U16001 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12918) );
  MUX2_X1 U16002 ( .A(n19349), .B(n16351), .S(n12918), .Z(n12919) );
  INV_X1 U16003 ( .A(n12919), .ZN(n12920) );
  OAI211_X1 U16004 ( .C1(n19376), .C2(n19175), .A(n12921), .B(n12920), .ZN(
        P2_U3013) );
  INV_X1 U16005 ( .A(n12922), .ZN(n12926) );
  OAI21_X1 U16006 ( .B1(n16325), .B2(n12924), .A(n12923), .ZN(n12925) );
  AOI21_X1 U16007 ( .B1(n19355), .B2(n12926), .A(n12925), .ZN(n12929) );
  OAI21_X1 U16008 ( .B1(n19349), .B2(n12927), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12928) );
  OAI211_X1 U16009 ( .C1(n15624), .C2(n19376), .A(n12929), .B(n12928), .ZN(
        P2_U3014) );
  NAND2_X1 U16010 ( .A1(n12932), .A2(n12931), .ZN(n12933) );
  NAND2_X1 U16011 ( .A1(n12934), .A2(n12933), .ZN(n12997) );
  OAI21_X1 U16012 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12935), .A(
        n20006), .ZN(n12936) );
  NOR2_X1 U16013 ( .A1(n12936), .A2(n19913), .ZN(n12937) );
  AOI21_X1 U16014 ( .B1(n12938), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12937), .ZN(n12939) );
  OAI21_X1 U16015 ( .B1(n12941), .B2(n12940), .A(n12939), .ZN(n12944) );
  NAND2_X1 U16016 ( .A1(n12995), .A2(n12945), .ZN(n12996) );
  INV_X1 U16017 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12946) );
  MUX2_X1 U16018 ( .A(n12946), .B(n12941), .S(n14998), .Z(n12947) );
  OAI21_X1 U16019 ( .B1(n19630), .B2(n15025), .A(n12947), .ZN(P2_U2884) );
  NAND2_X1 U16020 ( .A1(n11066), .A2(n20267), .ZN(n12950) );
  AND2_X1 U16021 ( .A1(n12950), .A2(n20292), .ZN(n12951) );
  OAI211_X1 U16022 ( .C1(n11969), .C2(n20246), .A(n12952), .B(n12951), .ZN(
        n12953) );
  NAND2_X1 U16023 ( .A1(n12953), .A2(n20262), .ZN(n12955) );
  OAI211_X1 U16024 ( .C1(n11963), .C2(n14053), .A(n12955), .B(n12954), .ZN(
        n12956) );
  INV_X1 U16025 ( .A(n12956), .ZN(n12958) );
  AND2_X1 U16026 ( .A1(n13229), .A2(n20246), .ZN(n12957) );
  NAND2_X1 U16027 ( .A1(n11070), .A2(n12957), .ZN(n12984) );
  AND3_X1 U16028 ( .A1(n12959), .A2(n12958), .A3(n12984), .ZN(n13249) );
  NOR2_X1 U16029 ( .A1(n12960), .A2(n14305), .ZN(n12961) );
  NAND3_X1 U16030 ( .A1(n11946), .A2(n13249), .A3(n12961), .ZN(n14824) );
  NAND2_X1 U16031 ( .A1(n20541), .A2(n14824), .ZN(n12978) );
  OR2_X1 U16032 ( .A1(n13245), .A2(n12962), .ZN(n13163) );
  INV_X1 U16033 ( .A(n12963), .ZN(n14829) );
  NAND2_X1 U16034 ( .A1(n14829), .A2(n12964), .ZN(n13164) );
  XNOR2_X1 U16035 ( .A(n13164), .B(n10052), .ZN(n12976) );
  INV_X1 U16036 ( .A(n12965), .ZN(n12968) );
  NAND2_X1 U16037 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12966) );
  NAND2_X1 U16038 ( .A1(n10052), .A2(n12966), .ZN(n12967) );
  NAND3_X1 U16039 ( .A1(n14823), .A2(n12968), .A3(n12967), .ZN(n12974) );
  NAND2_X1 U16040 ( .A1(n12970), .A2(n12969), .ZN(n12971) );
  NOR2_X1 U16041 ( .A1(n12972), .A2(n12971), .ZN(n13167) );
  OAI21_X1 U16042 ( .B1(n13165), .B2(n10052), .A(n10952), .ZN(n12979) );
  NAND2_X1 U16043 ( .A1(n13167), .A2(n12979), .ZN(n12973) );
  NAND2_X1 U16044 ( .A1(n12974), .A2(n12973), .ZN(n12975) );
  AOI21_X1 U16045 ( .B1(n13163), .B2(n12976), .A(n12975), .ZN(n12977) );
  NAND2_X1 U16046 ( .A1(n12978), .A2(n12977), .ZN(n13174) );
  INV_X1 U16047 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20669) );
  AOI22_X1 U16048 ( .A1(n13174), .A2(n16255), .B1(n15956), .B2(n12979), .ZN(
        n12991) );
  INV_X1 U16049 ( .A(n12014), .ZN(n12980) );
  NAND2_X1 U16050 ( .A1(n12981), .A2(n12980), .ZN(n12983) );
  OAI211_X1 U16051 ( .C1(n14043), .C2(n15973), .A(n12983), .B(n12982), .ZN(
        n12989) );
  OR2_X1 U16052 ( .A1(n12722), .A2(n13035), .ZN(n12985) );
  OAI21_X1 U16053 ( .B1(n20267), .B2(n13348), .A(n13234), .ZN(n12986) );
  INV_X1 U16054 ( .A(n12986), .ZN(n12988) );
  NAND2_X1 U16055 ( .A1(n13245), .A2(n13231), .ZN(n13020) );
  NAND2_X1 U16056 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16262), .ZN(n16270) );
  INV_X1 U16057 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20064) );
  OAI22_X1 U16058 ( .A1(n15939), .A2(n20057), .B1(n16270), .B2(n20064), .ZN(
        n16254) );
  AOI21_X1 U16059 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20868), .A(n16254), 
        .ZN(n14833) );
  NAND2_X1 U16060 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14833), .ZN(
        n12990) );
  OAI21_X1 U16061 ( .B1(n12991), .B2(n14833), .A(n12990), .ZN(P1_U3469) );
  AOI22_X1 U16062 ( .A1(n20368), .A2(n14824), .B1(n14825), .B2(n10914), .ZN(
        n15933) );
  OAI21_X1 U16063 ( .B1(n15933), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20867), 
        .ZN(n12992) );
  INV_X1 U16064 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13290) );
  NOR2_X1 U16065 ( .A1(n20867), .A2(n13290), .ZN(n14835) );
  INV_X1 U16066 ( .A(n14835), .ZN(n14832) );
  AOI22_X1 U16067 ( .A1(n12992), .A2(n14832), .B1(n15956), .B2(n10914), .ZN(
        n12994) );
  AOI21_X1 U16068 ( .B1(n14823), .B2(n16255), .A(n14833), .ZN(n12993) );
  OAI22_X1 U16069 ( .A1(n12994), .A2(n14833), .B1(n12993), .B2(n10914), .ZN(
        P1_U3474) );
  INV_X1 U16070 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12998) );
  NOR2_X1 U16071 ( .A1(n13008), .A2(n12998), .ZN(n13001) );
  INV_X1 U16072 ( .A(n13001), .ZN(n13000) );
  NAND2_X1 U16073 ( .A1(n19411), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12999) );
  NAND2_X1 U16074 ( .A1(n13000), .A2(n12999), .ZN(n13002) );
  NAND2_X1 U16075 ( .A1(n13010), .A2(n13001), .ZN(n13146) );
  OAI21_X1 U16076 ( .B1(n13010), .B2(n13002), .A(n13146), .ZN(n19252) );
  INV_X1 U16077 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19155) );
  OR2_X1 U16078 ( .A1(n13004), .A2(n13003), .ZN(n13005) );
  AND2_X1 U16079 ( .A1(n13005), .A2(n13148), .ZN(n19350) );
  INV_X1 U16080 ( .A(n19350), .ZN(n19158) );
  MUX2_X1 U16081 ( .A(n19155), .B(n19158), .S(n14998), .Z(n13006) );
  OAI21_X1 U16082 ( .B1(n19252), .B2(n15025), .A(n13006), .ZN(P2_U2883) );
  AND2_X1 U16083 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13191) );
  NAND4_X1 U16084 ( .A1(n13201), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .A4(n13191), .ZN(n13007) );
  NOR2_X1 U16085 ( .A1(n13008), .A2(n13007), .ZN(n13009) );
  XNOR2_X1 U16086 ( .A(n13127), .B(n13126), .ZN(n13015) );
  NOR2_X1 U16087 ( .A1(n13012), .A2(n13203), .ZN(n13013) );
  NOR2_X1 U16088 ( .A1(n13125), .A2(n13013), .ZN(n16328) );
  INV_X1 U16089 ( .A(n16328), .ZN(n19114) );
  MUX2_X1 U16090 ( .A(n10871), .B(n19114), .S(n14998), .Z(n13014) );
  OAI21_X1 U16091 ( .B1(n13015), .B2(n15025), .A(n13014), .ZN(P2_U2878) );
  OAI21_X1 U16092 ( .B1(n13017), .B2(n13016), .A(n13385), .ZN(n13366) );
  NAND2_X1 U16093 ( .A1(n13018), .A2(n14043), .ZN(n13019) );
  NAND2_X1 U16094 ( .A1(n13020), .A2(n13019), .ZN(n13021) );
  INV_X1 U16095 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13027) );
  MUX2_X1 U16096 ( .A(n14047), .B(n14008), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n13025) );
  INV_X1 U16097 ( .A(n14012), .ZN(n13435) );
  NAND2_X1 U16098 ( .A1(n13435), .A2(n13022), .ZN(n14031) );
  NAND2_X1 U16099 ( .A1(n13022), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13023) );
  AND2_X1 U16100 ( .A1(n14031), .A2(n13023), .ZN(n13024) );
  NAND2_X1 U16101 ( .A1(n13025), .A2(n13024), .ZN(n13295) );
  NAND2_X1 U16102 ( .A1(n14008), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13026) );
  OAI21_X1 U16103 ( .B1(n14073), .B2(P1_EBX_REG_0__SCAN_IN), .A(n13026), .ZN(
        n13115) );
  XNOR2_X1 U16104 ( .A(n13295), .B(n13115), .ZN(n13360) );
  XNOR2_X1 U16105 ( .A(n13360), .B(n13022), .ZN(n13244) );
  OAI222_X1 U16106 ( .A1(n13366), .A2(n16075), .B1(n20161), .B2(n13027), .C1(
        n13244), .C2(n16076), .ZN(P1_U2871) );
  NAND3_X1 U16107 ( .A1(n20868), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16261) );
  INV_X1 U16108 ( .A(n16261), .ZN(n13028) );
  XNOR2_X1 U16109 ( .A(n13270), .B(n13269), .ZN(n13030) );
  OAI211_X1 U16110 ( .C1(n13030), .C2(n20954), .A(n13029), .B(n11965), .ZN(
        n13031) );
  INV_X1 U16111 ( .A(n13031), .ZN(n13032) );
  NAND2_X1 U16112 ( .A1(n11043), .A2(n20272), .ZN(n13276) );
  OAI21_X1 U16113 ( .B1(n20954), .B2(n13270), .A(n13276), .ZN(n13033) );
  INV_X1 U16114 ( .A(n13033), .ZN(n13034) );
  NAND2_X1 U16115 ( .A1(n13048), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13284) );
  XOR2_X1 U16116 ( .A(n13281), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n13217) );
  NAND2_X1 U16117 ( .A1(n13035), .A2(n11969), .ZN(n15947) );
  NAND2_X1 U16118 ( .A1(n13217), .A2(n16141), .ZN(n13043) );
  INV_X1 U16119 ( .A(n20797), .ZN(n20706) );
  NAND2_X1 U16120 ( .A1(n20706), .A2(n13040), .ZN(n20950) );
  NAND2_X1 U16121 ( .A1(n20950), .A2(n20868), .ZN(n13037) );
  NAND2_X1 U16122 ( .A1(n20868), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13039) );
  NAND2_X1 U16123 ( .A1(n20736), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U16124 ( .A1(n13039), .A2(n13038), .ZN(n13049) );
  OR2_X2 U16125 ( .A1(n13040), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20227) );
  INV_X1 U16126 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20939) );
  NOR2_X1 U16127 ( .A1(n20227), .A2(n20939), .ZN(n13254) );
  NOR2_X1 U16128 ( .A1(n16144), .A2(n13364), .ZN(n13041) );
  AOI211_X1 U16129 ( .C1(n16138), .C2(n13364), .A(n13254), .B(n13041), .ZN(
        n13042) );
  OAI211_X1 U16130 ( .C1(n20243), .C2(n13366), .A(n13043), .B(n13042), .ZN(
        P1_U2998) );
  INV_X1 U16131 ( .A(n13044), .ZN(n13047) );
  OAI21_X1 U16132 ( .B1(n13047), .B2(n13046), .A(n13045), .ZN(n13414) );
  OAI21_X1 U16133 ( .B1(n13048), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13284), .ZN(n13268) );
  INV_X2 U16134 ( .A(n20227), .ZN(n16236) );
  NAND2_X1 U16135 ( .A1(n16236), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13261) );
  OAI21_X1 U16136 ( .B1(n16128), .B2(n13049), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13050) );
  OAI211_X1 U16137 ( .C1(n13268), .C2(n20063), .A(n13261), .B(n13050), .ZN(
        n13051) );
  INV_X1 U16138 ( .A(n13051), .ZN(n13052) );
  OAI21_X1 U16139 ( .B1(n20243), .B2(n13414), .A(n13052), .ZN(P1_U2999) );
  INV_X1 U16140 ( .A(n19630), .ZN(n20010) );
  INV_X1 U16141 ( .A(n13717), .ZN(n15635) );
  OR2_X1 U16142 ( .A1(n12941), .A2(n15635), .ZN(n13068) );
  NAND2_X1 U16143 ( .A1(n13054), .A2(n13053), .ZN(n15631) );
  NAND2_X1 U16144 ( .A1(n15631), .A2(n9664), .ZN(n13060) );
  INV_X1 U16145 ( .A(n13056), .ZN(n13057) );
  NAND2_X1 U16146 ( .A1(n13057), .A2(n15646), .ZN(n15630) );
  INV_X1 U16147 ( .A(n12252), .ZN(n13059) );
  NAND2_X1 U16148 ( .A1(n13058), .A2(n13059), .ZN(n15633) );
  NAND3_X1 U16149 ( .A1(n13060), .A2(n15630), .A3(n15633), .ZN(n13065) );
  NAND2_X1 U16150 ( .A1(n16393), .A2(n13061), .ZN(n15640) );
  NAND2_X1 U16151 ( .A1(n15640), .A2(n15630), .ZN(n13063) );
  NAND2_X1 U16152 ( .A1(n13058), .A2(n12252), .ZN(n13062) );
  NAND2_X1 U16153 ( .A1(n13063), .A2(n13062), .ZN(n13064) );
  MUX2_X1 U16154 ( .A(n13065), .B(n13064), .S(n10383), .Z(n13066) );
  NOR2_X1 U16155 ( .A1(n13066), .A2(n10663), .ZN(n13067) );
  NAND2_X1 U16156 ( .A1(n13068), .A2(n13067), .ZN(n16398) );
  AOI22_X1 U16157 ( .A1(n20010), .A2(n16421), .B1(n15625), .B2(n16398), .ZN(
        n13070) );
  NAND2_X1 U16158 ( .A1(n13725), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13069) );
  OAI21_X1 U16159 ( .B1(n13070), .B2(n13725), .A(n13069), .ZN(P2_U3596) );
  NAND2_X1 U16160 ( .A1(n13072), .A2(n13071), .ZN(n13075) );
  INV_X1 U16161 ( .A(n13073), .ZN(n13074) );
  NAND2_X1 U16162 ( .A1(n13075), .A2(n13074), .ZN(n20021) );
  INV_X1 U16163 ( .A(n20021), .ZN(n13086) );
  XNOR2_X1 U16164 ( .A(n20019), .B(n20021), .ZN(n13082) );
  OAI21_X1 U16165 ( .B1(n13076), .B2(n13078), .A(n13077), .ZN(n20031) );
  NOR2_X1 U16166 ( .A1(n20028), .A2(n20031), .ZN(n13079) );
  AOI21_X1 U16167 ( .B1(n20028), .B2(n20031), .A(n13079), .ZN(n19268) );
  NAND2_X1 U16168 ( .A1(n19629), .A2(n19184), .ZN(n19267) );
  NAND2_X1 U16169 ( .A1(n19268), .A2(n19267), .ZN(n19266) );
  INV_X1 U16170 ( .A(n13079), .ZN(n13080) );
  NAND2_X1 U16171 ( .A1(n19266), .A2(n13080), .ZN(n13081) );
  NAND2_X1 U16172 ( .A1(n13082), .A2(n13081), .ZN(n19242) );
  OAI21_X1 U16173 ( .B1(n13082), .B2(n13081), .A(n19242), .ZN(n13083) );
  NAND2_X1 U16174 ( .A1(n13083), .A2(n19269), .ZN(n13085) );
  AOI22_X1 U16175 ( .A1(n19241), .A2(n16317), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19264), .ZN(n13084) );
  OAI211_X1 U16176 ( .C1(n13086), .C2(n19215), .A(n13085), .B(n13084), .ZN(
        P2_U2917) );
  NAND2_X1 U16177 ( .A1(n20954), .A2(n20881), .ZN(n13087) );
  NAND2_X1 U16178 ( .A1(n13110), .A2(n13352), .ZN(n13112) );
  INV_X2 U16179 ( .A(n13112), .ZN(n20217) );
  INV_X2 U16180 ( .A(n13110), .ZN(n20220) );
  AOI22_X1 U16181 ( .A1(n20217), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20220), .ZN(n13092) );
  NOR2_X2 U16182 ( .A1(n20220), .A2(n13352), .ZN(n20205) );
  NAND2_X1 U16183 ( .A1(n20242), .A2(DATAI_4_), .ZN(n13090) );
  NAND2_X1 U16184 ( .A1(n20241), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13089) );
  AND2_X1 U16185 ( .A1(n13090), .A2(n13089), .ZN(n20278) );
  INV_X1 U16186 ( .A(n20278), .ZN(n13091) );
  NAND2_X1 U16187 ( .A1(n20205), .A2(n13091), .ZN(n13320) );
  NAND2_X1 U16188 ( .A1(n13092), .A2(n13320), .ZN(P1_U2956) );
  AOI22_X1 U16189 ( .A1(n20217), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20220), .ZN(n13096) );
  NAND2_X1 U16190 ( .A1(n20242), .A2(DATAI_7_), .ZN(n13094) );
  NAND2_X1 U16191 ( .A1(n20241), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13093) );
  AND2_X1 U16192 ( .A1(n13094), .A2(n13093), .ZN(n20296) );
  INV_X1 U16193 ( .A(n20296), .ZN(n13095) );
  NAND2_X1 U16194 ( .A1(n20205), .A2(n13095), .ZN(n13318) );
  NAND2_X1 U16195 ( .A1(n13096), .A2(n13318), .ZN(P1_U2959) );
  AOI22_X1 U16196 ( .A1(n20217), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20220), .ZN(n13100) );
  NAND2_X1 U16197 ( .A1(n20242), .A2(DATAI_5_), .ZN(n13098) );
  NAND2_X1 U16198 ( .A1(n20241), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13097) );
  AND2_X1 U16199 ( .A1(n13098), .A2(n13097), .ZN(n20282) );
  INV_X1 U16200 ( .A(n20282), .ZN(n13099) );
  NAND2_X1 U16201 ( .A1(n20205), .A2(n13099), .ZN(n13310) );
  NAND2_X1 U16202 ( .A1(n13100), .A2(n13310), .ZN(P1_U2957) );
  AOI22_X1 U16203 ( .A1(n20217), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20220), .ZN(n13104) );
  NAND2_X1 U16204 ( .A1(n20242), .A2(DATAI_3_), .ZN(n13102) );
  NAND2_X1 U16205 ( .A1(n20241), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13101) );
  AND2_X1 U16206 ( .A1(n13102), .A2(n13101), .ZN(n20274) );
  INV_X1 U16207 ( .A(n20274), .ZN(n13103) );
  NAND2_X1 U16208 ( .A1(n20205), .A2(n13103), .ZN(n13308) );
  NAND2_X1 U16209 ( .A1(n13104), .A2(n13308), .ZN(P1_U2955) );
  INV_X1 U16210 ( .A(DATAI_10_), .ZN(n13105) );
  INV_X1 U16211 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16548) );
  MUX2_X1 U16212 ( .A(n13105), .B(n16548), .S(n20241), .Z(n14393) );
  INV_X1 U16213 ( .A(n14393), .ZN(n13106) );
  NAND2_X1 U16214 ( .A1(n20205), .A2(n13106), .ZN(n20211) );
  NAND2_X1 U16215 ( .A1(n20220), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13107) );
  OAI211_X1 U16216 ( .C1(n14330), .C2(n13112), .A(n20211), .B(n13107), .ZN(
        P1_U2947) );
  INV_X1 U16217 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14383) );
  INV_X1 U16218 ( .A(n20205), .ZN(n13111) );
  INV_X1 U16219 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13108) );
  NOR2_X1 U16220 ( .A1(n20242), .A2(n13108), .ZN(n13109) );
  AOI21_X1 U16221 ( .B1(DATAI_15_), .B2(n20242), .A(n13109), .ZN(n14382) );
  INV_X1 U16222 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20163) );
  OAI222_X1 U16223 ( .A1(n13112), .A2(n14383), .B1(n13111), .B2(n14382), .C1(
        n13110), .C2(n20163), .ZN(P1_U2967) );
  OR2_X1 U16224 ( .A1(n14055), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13114) );
  NAND2_X1 U16225 ( .A1(n13115), .A2(n13114), .ZN(n13260) );
  INV_X1 U16226 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13116) );
  OAI222_X1 U16227 ( .A1(n13260), .A2(n16076), .B1(n13116), .B2(n20161), .C1(
        n13414), .C2(n16075), .ZN(P1_U2872) );
  NOR2_X1 U16228 ( .A1(n13146), .A2(n13117), .ZN(n13192) );
  XNOR2_X1 U16229 ( .A(n13192), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13123) );
  INV_X1 U16230 ( .A(n13118), .ZN(n13120) );
  INV_X1 U16231 ( .A(n13119), .ZN(n13195) );
  AOI21_X1 U16232 ( .B1(n13120), .B2(n9762), .A(n13195), .ZN(n19137) );
  NOR2_X1 U16233 ( .A1(n14998), .A2(n19130), .ZN(n13121) );
  AOI21_X1 U16234 ( .B1(n19137), .B2(n14998), .A(n13121), .ZN(n13122) );
  OAI21_X1 U16235 ( .B1(n13123), .B2(n15025), .A(n13122), .ZN(P2_U2881) );
  OAI21_X1 U16236 ( .B1(n13125), .B2(n13124), .A(n13212), .ZN(n19103) );
  OAI211_X1 U16237 ( .C1(n13128), .C2(n13130), .A(n13129), .B(n15012), .ZN(
        n13132) );
  NAND2_X1 U16238 ( .A1(n15015), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13131) );
  OAI211_X1 U16239 ( .C1(n19103), .C2(n15004), .A(n13132), .B(n13131), .ZN(
        P2_U2877) );
  INV_X1 U16240 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13134) );
  AOI22_X1 U16241 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13133) );
  OAI21_X1 U16242 ( .B1(n13134), .B2(n13145), .A(n13133), .ZN(P1_U2913) );
  AOI22_X1 U16243 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13135) );
  OAI21_X1 U16244 ( .B1(n14370), .B2(n13145), .A(n13135), .ZN(P1_U2919) );
  AOI22_X1 U16245 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13136) );
  OAI21_X1 U16246 ( .B1(n14364), .B2(n13145), .A(n13136), .ZN(P1_U2918) );
  INV_X1 U16247 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13138) );
  AOI22_X1 U16248 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13137) );
  OAI21_X1 U16249 ( .B1(n13138), .B2(n13145), .A(n13137), .ZN(P1_U2917) );
  AOI22_X1 U16250 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13139) );
  OAI21_X1 U16251 ( .B1(n14357), .B2(n13145), .A(n13139), .ZN(P1_U2916) );
  INV_X1 U16252 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13141) );
  AOI22_X1 U16253 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13140) );
  OAI21_X1 U16254 ( .B1(n13141), .B2(n13145), .A(n13140), .ZN(P1_U2920) );
  INV_X1 U16255 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13143) );
  AOI22_X1 U16256 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13142) );
  OAI21_X1 U16257 ( .B1(n13143), .B2(n13145), .A(n13142), .ZN(P1_U2914) );
  AOI22_X1 U16258 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13144) );
  OAI21_X1 U16259 ( .B1(n14352), .B2(n13145), .A(n13144), .ZN(P1_U2915) );
  INV_X1 U16260 ( .A(n13146), .ZN(n13147) );
  INV_X1 U16261 ( .A(n13192), .ZN(n13190) );
  OAI211_X1 U16262 ( .C1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .C2(n13147), .A(
        n13190), .B(n15012), .ZN(n13152) );
  NAND2_X1 U16263 ( .A1(n13149), .A2(n13148), .ZN(n13150) );
  AND2_X1 U16264 ( .A1(n13150), .A2(n9762), .ZN(n19148) );
  NAND2_X1 U16265 ( .A1(n14998), .A2(n19148), .ZN(n13151) );
  OAI211_X1 U16266 ( .C1(n14998), .C2(n13153), .A(n13152), .B(n13151), .ZN(
        P2_U2882) );
  INV_X1 U16267 ( .A(n11046), .ZN(n13154) );
  NAND2_X1 U16268 ( .A1(n13154), .A2(n20292), .ZN(n13155) );
  INV_X1 U16269 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20982) );
  NAND2_X1 U16270 ( .A1(n20242), .A2(DATAI_0_), .ZN(n13158) );
  NAND2_X1 U16271 ( .A1(n20241), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13157) );
  AND2_X1 U16272 ( .A1(n13158), .A2(n13157), .ZN(n20254) );
  OAI222_X1 U16273 ( .A1(n14396), .A2(n13414), .B1(n14389), .B2(n20982), .C1(
        n14394), .C2(n20254), .ZN(P1_U2904) );
  NAND2_X1 U16274 ( .A1(n20242), .A2(DATAI_1_), .ZN(n13160) );
  NAND2_X1 U16275 ( .A1(n20241), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13159) );
  AND2_X1 U16276 ( .A1(n13160), .A2(n13159), .ZN(n20264) );
  OAI222_X1 U16277 ( .A1(n14396), .A2(n13366), .B1(n14389), .B2(n11197), .C1(
        n14394), .C2(n20264), .ZN(P1_U2903) );
  NOR2_X1 U16278 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20867), .ZN(n13183) );
  INV_X1 U16279 ( .A(n13162), .ZN(n20252) );
  INV_X1 U16280 ( .A(n13163), .ZN(n13170) );
  INV_X1 U16281 ( .A(n13164), .ZN(n13166) );
  NOR2_X1 U16282 ( .A1(n13166), .A2(n13165), .ZN(n14837) );
  XNOR2_X1 U16283 ( .A(n10051), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13168) );
  AOI22_X1 U16284 ( .A1(n14823), .A2(n13168), .B1(n13167), .B2(n14837), .ZN(
        n13169) );
  OAI21_X1 U16285 ( .B1(n13170), .B2(n14837), .A(n13169), .ZN(n13171) );
  AOI21_X1 U16286 ( .B1(n20252), .B2(n14824), .A(n13171), .ZN(n14840) );
  INV_X1 U16287 ( .A(n14840), .ZN(n13172) );
  INV_X1 U16288 ( .A(n15939), .ZN(n13173) );
  MUX2_X1 U16289 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13172), .S(
        n13173), .Z(n15941) );
  AOI22_X1 U16290 ( .A1(n13183), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15941), .B2(n20867), .ZN(n13176) );
  MUX2_X1 U16291 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13174), .S(
        n13173), .Z(n15932) );
  AOI22_X1 U16292 ( .A1(n13183), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20867), .B2(n15932), .ZN(n13175) );
  NOR2_X1 U16293 ( .A1(n13176), .A2(n13175), .ZN(n15950) );
  INV_X1 U16294 ( .A(n13177), .ZN(n14828) );
  NAND2_X1 U16295 ( .A1(n15950), .A2(n14828), .ZN(n13186) );
  INV_X1 U16296 ( .A(n20406), .ZN(n20666) );
  OR2_X1 U16297 ( .A1(n13178), .A2(n20666), .ZN(n13179) );
  XNOR2_X1 U16298 ( .A(n13179), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14238) );
  INV_X1 U16299 ( .A(n11946), .ZN(n13180) );
  AND2_X1 U16300 ( .A1(n14238), .A2(n13180), .ZN(n16256) );
  OAI21_X1 U16301 ( .B1(n16256), .B2(n15939), .A(n20867), .ZN(n13181) );
  AOI21_X1 U16302 ( .B1(n15939), .B2(n16258), .A(n13181), .ZN(n13182) );
  AOI21_X1 U16303 ( .B1(n13183), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13182), .ZN(n15948) );
  AND3_X1 U16304 ( .A1(n13186), .A2(n15948), .A3(n20064), .ZN(n13185) );
  NOR2_X1 U16305 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20955) );
  AND3_X1 U16306 ( .A1(n13186), .A2(n15948), .A3(n16262), .ZN(n15958) );
  INV_X1 U16307 ( .A(n20368), .ZN(n13410) );
  NAND2_X1 U16308 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20669), .ZN(n13367) );
  INV_X1 U16309 ( .A(n13367), .ZN(n13187) );
  OAI22_X1 U16310 ( .A1(n20328), .A2(n20706), .B1(n13410), .B2(n13187), .ZN(
        n13188) );
  OAI21_X1 U16311 ( .B1(n15958), .B2(n13188), .A(n20239), .ZN(n13189) );
  OAI21_X1 U16312 ( .B1(n20239), .B2(n20696), .A(n13189), .ZN(P1_U3478) );
  NOR2_X1 U16313 ( .A1(n13190), .A2(n10698), .ZN(n13193) );
  NAND2_X1 U16314 ( .A1(n13192), .A2(n13191), .ZN(n13200) );
  OAI211_X1 U16315 ( .C1(n13193), .C2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n15012), .B(n13200), .ZN(n13198) );
  INV_X1 U16316 ( .A(n13194), .ZN(n13204) );
  OAI21_X1 U16317 ( .B1(n13196), .B2(n13195), .A(n13204), .ZN(n19124) );
  INV_X1 U16318 ( .A(n19124), .ZN(n16376) );
  NAND2_X1 U16319 ( .A1(n16376), .A2(n14998), .ZN(n13197) );
  OAI211_X1 U16320 ( .C1(n14998), .C2(n13199), .A(n13198), .B(n13197), .ZN(
        P2_U2880) );
  XOR2_X1 U16321 ( .A(n13201), .B(n13200), .Z(n13207) );
  INV_X1 U16322 ( .A(n13202), .ZN(n13205) );
  AOI21_X1 U16323 ( .B1(n13205), .B2(n13204), .A(n13203), .ZN(n16362) );
  INV_X1 U16324 ( .A(n16362), .ZN(n13562) );
  MUX2_X1 U16325 ( .A(n10870), .B(n13562), .S(n14998), .Z(n13206) );
  OAI21_X1 U16326 ( .B1(n13207), .B2(n15025), .A(n13206), .ZN(P2_U2879) );
  OAI211_X1 U16327 ( .C1(n13209), .C2(n13210), .A(n15012), .B(n13379), .ZN(
        n13215) );
  AND2_X1 U16328 ( .A1(n13212), .A2(n13211), .ZN(n13213) );
  OR2_X1 U16329 ( .A1(n13213), .A2(n9763), .ZN(n15558) );
  INV_X1 U16330 ( .A(n15558), .ZN(n19092) );
  NAND2_X1 U16331 ( .A1(n19092), .A2(n14998), .ZN(n13214) );
  OAI211_X1 U16332 ( .C1(n14998), .C2(n13216), .A(n13215), .B(n13214), .ZN(
        P2_U2876) );
  INV_X1 U16333 ( .A(n13217), .ZN(n13259) );
  NAND2_X1 U16334 ( .A1(n20262), .A2(n13351), .ZN(n13220) );
  INV_X1 U16335 ( .A(n13218), .ZN(n13219) );
  NAND2_X1 U16336 ( .A1(n13220), .A2(n13219), .ZN(n13228) );
  AOI21_X1 U16337 ( .B1(n12014), .B2(n20951), .A(n11043), .ZN(n13223) );
  NOR2_X1 U16338 ( .A1(n20954), .A2(n15973), .ZN(n13222) );
  OAI21_X1 U16339 ( .B1(n13223), .B2(n13222), .A(n13221), .ZN(n13225) );
  NAND2_X1 U16340 ( .A1(n13225), .A2(n13224), .ZN(n13227) );
  MUX2_X1 U16341 ( .A(n13228), .B(n13227), .S(n13226), .Z(n13233) );
  INV_X1 U16342 ( .A(n13229), .ZN(n13230) );
  NAND2_X1 U16343 ( .A1(n13231), .A2(n13230), .ZN(n13232) );
  NAND3_X1 U16344 ( .A1(n13234), .A2(n13233), .A3(n13232), .ZN(n13236) );
  OAI21_X1 U16345 ( .B1(n13238), .B2(n13242), .A(n13237), .ZN(n13239) );
  OR2_X1 U16346 ( .A1(n13240), .A2(n13239), .ZN(n13241) );
  OAI22_X1 U16347 ( .A1(n12723), .A2(n20262), .B1(n11047), .B2(n13242), .ZN(
        n13243) );
  INV_X1 U16348 ( .A(n13244), .ZN(n13255) );
  NAND2_X1 U16349 ( .A1(n13256), .A2(n13245), .ZN(n20229) );
  MUX2_X1 U16350 ( .A(n13246), .B(n13226), .S(n20246), .Z(n13247) );
  NAND3_X1 U16351 ( .A1(n13249), .A2(n13248), .A3(n13247), .ZN(n13250) );
  NAND2_X1 U16352 ( .A1(n13256), .A2(n13250), .ZN(n14788) );
  INV_X1 U16353 ( .A(n14788), .ZN(n13262) );
  NAND2_X1 U16354 ( .A1(n13262), .A2(n13290), .ZN(n13252) );
  INV_X1 U16355 ( .A(n13256), .ZN(n13251) );
  NAND2_X1 U16356 ( .A1(n13251), .A2(n20227), .ZN(n14785) );
  INV_X1 U16357 ( .A(n16171), .ZN(n13291) );
  AOI21_X1 U16358 ( .B1(n16175), .B2(n13290), .A(n13291), .ZN(n13264) );
  INV_X1 U16359 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14822) );
  NOR2_X1 U16360 ( .A1(n13264), .A2(n14822), .ZN(n13253) );
  AOI211_X1 U16361 ( .C1(n16243), .C2(n13255), .A(n13254), .B(n13253), .ZN(
        n13258) );
  NAND2_X1 U16362 ( .A1(n13256), .A2(n14823), .ZN(n14783) );
  OR3_X1 U16363 ( .A1(n14798), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13293), .ZN(n13257) );
  OAI211_X1 U16364 ( .C1(n13259), .C2(n20230), .A(n13258), .B(n13257), .ZN(
        P1_U3030) );
  INV_X1 U16365 ( .A(n13260), .ZN(n13406) );
  INV_X2 U16366 ( .A(n16200), .ZN(n16243) );
  INV_X1 U16367 ( .A(n13261), .ZN(n13266) );
  NOR3_X1 U16368 ( .A1(n16175), .A2(n13262), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13263) );
  AOI21_X1 U16369 ( .B1(n13264), .B2(n14783), .A(n13263), .ZN(n13265) );
  AOI211_X1 U16370 ( .C1(n13406), .C2(n16243), .A(n13266), .B(n13265), .ZN(
        n13267) );
  OAI21_X1 U16371 ( .B1(n13268), .B2(n20230), .A(n13267), .ZN(P1_U3031) );
  NAND2_X1 U16372 ( .A1(n13270), .A2(n13269), .ZN(n13274) );
  NAND2_X1 U16373 ( .A1(n13274), .A2(n13275), .ZN(n13500) );
  INV_X1 U16374 ( .A(n13499), .ZN(n13271) );
  XNOR2_X1 U16375 ( .A(n13500), .B(n13271), .ZN(n13272) );
  INV_X1 U16376 ( .A(n20954), .ZN(n14435) );
  NAND2_X1 U16377 ( .A1(n13272), .A2(n14435), .ZN(n13273) );
  OAI21_X2 U16378 ( .B1(n13371), .B2(n14429), .A(n13273), .ZN(n13494) );
  INV_X1 U16379 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13516) );
  XNOR2_X1 U16380 ( .A(n13494), .B(n13516), .ZN(n13289) );
  OR2_X1 U16381 ( .A1(n13368), .A2(n14429), .ZN(n13280) );
  OAI21_X1 U16382 ( .B1(n13275), .B2(n13274), .A(n13500), .ZN(n13278) );
  INV_X1 U16383 ( .A(n13276), .ZN(n13277) );
  AOI21_X1 U16384 ( .B1(n14435), .B2(n13278), .A(n13277), .ZN(n13279) );
  NAND2_X1 U16385 ( .A1(n13280), .A2(n13279), .ZN(n13396) );
  NAND2_X1 U16386 ( .A1(n13281), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13286) );
  INV_X1 U16387 ( .A(n13282), .ZN(n13283) );
  INV_X1 U16388 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20237) );
  XNOR2_X1 U16389 ( .A(n13287), .B(n20237), .ZN(n13397) );
  NAND2_X1 U16390 ( .A1(n13396), .A2(n13397), .ZN(n13493) );
  NAND2_X1 U16391 ( .A1(n13287), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13491) );
  NAND2_X1 U16392 ( .A1(n13493), .A2(n13491), .ZN(n13288) );
  XNOR2_X1 U16393 ( .A(n13289), .B(n13288), .ZN(n13420) );
  OAI21_X1 U16394 ( .B1(n13290), .B2(n14822), .A(n20237), .ZN(n20224) );
  INV_X1 U16395 ( .A(n16197), .ZN(n16218) );
  NAND2_X1 U16396 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13292) );
  AOI21_X1 U16397 ( .B1(n16218), .B2(n13292), .A(n13291), .ZN(n20236) );
  OAI21_X1 U16398 ( .B1(n20229), .B2(n20224), .A(n20236), .ZN(n13513) );
  INV_X1 U16399 ( .A(n13292), .ZN(n20226) );
  NAND2_X1 U16400 ( .A1(n20226), .A2(n20223), .ZN(n16220) );
  NAND2_X1 U16401 ( .A1(n20229), .A2(n16220), .ZN(n14809) );
  NAND2_X1 U16402 ( .A1(n20224), .A2(n14809), .ZN(n16252) );
  INV_X1 U16403 ( .A(n16252), .ZN(n13294) );
  AOI22_X1 U16404 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13513), .B1(
        n13294), .B2(n13516), .ZN(n13303) );
  INV_X1 U16405 ( .A(n13295), .ZN(n13296) );
  AOI21_X1 U16406 ( .B1(n13360), .B2(n14043), .A(n13296), .ZN(n13389) );
  MUX2_X1 U16407 ( .A(n14047), .B(n14008), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13299) );
  NAND2_X1 U16408 ( .A1(n13022), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13297) );
  AND2_X1 U16409 ( .A1(n14031), .A2(n13297), .ZN(n13298) );
  NAND2_X1 U16410 ( .A1(n13299), .A2(n13298), .ZN(n13388) );
  NAND2_X1 U16411 ( .A1(n13389), .A2(n13388), .ZN(n13387) );
  MUX2_X1 U16412 ( .A(n14048), .B(n14053), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13300) );
  OAI21_X1 U16413 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14055), .A(
        n13300), .ZN(n13301) );
  AOI21_X1 U16414 ( .B1(n13387), .B2(n13301), .A(n10040), .ZN(n20144) );
  AND2_X1 U16415 ( .A1(n16236), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13416) );
  AOI21_X1 U16416 ( .B1(n20144), .B2(n16243), .A(n13416), .ZN(n13302) );
  OAI211_X1 U16417 ( .C1(n20230), .C2(n13420), .A(n13303), .B(n13302), .ZN(
        P1_U3028) );
  OAI21_X1 U16418 ( .B1(n13306), .B2(n13305), .A(n13304), .ZN(n13415) );
  AOI22_X1 U16419 ( .A1(n20144), .A2(n20156), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14296), .ZN(n13307) );
  OAI21_X1 U16420 ( .B1(n13415), .B2(n16075), .A(n13307), .ZN(P1_U2869) );
  AOI22_X1 U16421 ( .A1(n20217), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20220), .ZN(n13309) );
  NAND2_X1 U16422 ( .A1(n13309), .A2(n13308), .ZN(P1_U2940) );
  AOI22_X1 U16423 ( .A1(n20217), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20220), .ZN(n13311) );
  NAND2_X1 U16424 ( .A1(n13311), .A2(n13310), .ZN(P1_U2942) );
  AOI22_X1 U16425 ( .A1(n20217), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20220), .ZN(n13313) );
  INV_X1 U16426 ( .A(n20254), .ZN(n13312) );
  NAND2_X1 U16427 ( .A1(n20205), .A2(n13312), .ZN(n13326) );
  NAND2_X1 U16428 ( .A1(n13313), .A2(n13326), .ZN(P1_U2952) );
  AOI22_X1 U16429 ( .A1(n20217), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20220), .ZN(n13317) );
  NAND2_X1 U16430 ( .A1(n20242), .A2(DATAI_2_), .ZN(n13315) );
  NAND2_X1 U16431 ( .A1(n20241), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13314) );
  AND2_X1 U16432 ( .A1(n13315), .A2(n13314), .ZN(n20269) );
  INV_X1 U16433 ( .A(n20269), .ZN(n13316) );
  NAND2_X1 U16434 ( .A1(n20205), .A2(n13316), .ZN(n13328) );
  NAND2_X1 U16435 ( .A1(n13317), .A2(n13328), .ZN(P1_U2954) );
  AOI22_X1 U16436 ( .A1(n20217), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20220), .ZN(n13319) );
  NAND2_X1 U16437 ( .A1(n13319), .A2(n13318), .ZN(P1_U2944) );
  AOI22_X1 U16438 ( .A1(n20217), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20220), .ZN(n13321) );
  NAND2_X1 U16439 ( .A1(n13321), .A2(n13320), .ZN(P1_U2941) );
  AOI22_X1 U16440 ( .A1(n20217), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20220), .ZN(n13325) );
  NAND2_X1 U16441 ( .A1(n20242), .A2(DATAI_6_), .ZN(n13323) );
  NAND2_X1 U16442 ( .A1(n20241), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13322) );
  AND2_X1 U16443 ( .A1(n13323), .A2(n13322), .ZN(n20287) );
  INV_X1 U16444 ( .A(n20287), .ZN(n13324) );
  NAND2_X1 U16445 ( .A1(n20205), .A2(n13324), .ZN(n13330) );
  NAND2_X1 U16446 ( .A1(n13325), .A2(n13330), .ZN(P1_U2958) );
  AOI22_X1 U16447 ( .A1(n20217), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20220), .ZN(n13327) );
  NAND2_X1 U16448 ( .A1(n13327), .A2(n13326), .ZN(P1_U2937) );
  AOI22_X1 U16449 ( .A1(n20217), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20220), .ZN(n13329) );
  NAND2_X1 U16450 ( .A1(n13329), .A2(n13328), .ZN(P1_U2939) );
  AOI22_X1 U16451 ( .A1(n20217), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20220), .ZN(n13331) );
  NAND2_X1 U16452 ( .A1(n13331), .A2(n13330), .ZN(P1_U2943) );
  AOI22_X1 U16453 ( .A1(n20217), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20220), .ZN(n13333) );
  INV_X1 U16454 ( .A(n20264), .ZN(n13332) );
  NAND2_X1 U16455 ( .A1(n20205), .A2(n13332), .ZN(n13334) );
  NAND2_X1 U16456 ( .A1(n13333), .A2(n13334), .ZN(P1_U2953) );
  AOI22_X1 U16457 ( .A1(n20217), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20220), .ZN(n13335) );
  NAND2_X1 U16458 ( .A1(n13335), .A2(n13334), .ZN(P1_U2938) );
  OAI222_X1 U16459 ( .A1(n14396), .A2(n13415), .B1(n14389), .B2(n11244), .C1(
        n14394), .C2(n20274), .ZN(P1_U2901) );
  INV_X1 U16460 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14466) );
  INV_X1 U16461 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13337) );
  AND2_X1 U16462 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20868), .ZN(n13339) );
  AND2_X1 U16463 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20955), .ZN(n16269) );
  AOI22_X1 U16464 ( .A1(n13340), .A2(n13339), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16269), .ZN(n13341) );
  NAND2_X1 U16465 ( .A1(n20227), .A2(n13341), .ZN(n13342) );
  NAND2_X1 U16466 ( .A1(n14232), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13345) );
  INV_X1 U16467 ( .A(n20949), .ZN(n13349) );
  NOR2_X1 U16468 ( .A1(n13349), .A2(n13343), .ZN(n13344) );
  OR2_X1 U16469 ( .A1(n20119), .A2(n13344), .ZN(n20147) );
  INV_X1 U16470 ( .A(n20147), .ZN(n20132) );
  INV_X1 U16471 ( .A(n13345), .ZN(n13346) );
  NOR2_X1 U16472 ( .A1(n13349), .A2(n13348), .ZN(n20142) );
  INV_X1 U16473 ( .A(n20142), .ZN(n13409) );
  AND2_X1 U16474 ( .A1(n20951), .A2(n20736), .ZN(n15954) );
  INV_X1 U16475 ( .A(n15954), .ZN(n13350) );
  AOI21_X1 U16476 ( .B1(n13352), .B2(n13351), .A(n13350), .ZN(n13356) );
  NAND2_X1 U16477 ( .A1(n20262), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13357) );
  INV_X1 U16478 ( .A(n13357), .ZN(n13353) );
  NOR2_X1 U16479 ( .A1(n13356), .A2(n13353), .ZN(n13354) );
  NAND2_X1 U16480 ( .A1(n14232), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20111) );
  OAI22_X1 U16481 ( .A1(n20111), .A2(n13364), .B1(n14232), .B2(n20939), .ZN(
        n13355) );
  AOI21_X1 U16482 ( .B1(n20143), .B2(P1_EBX_REG_1__SCAN_IN), .A(n13355), .ZN(
        n13362) );
  INV_X1 U16483 ( .A(n20102), .ZN(n20094) );
  NOR2_X1 U16484 ( .A1(n13357), .A2(n15954), .ZN(n13358) );
  AOI22_X1 U16485 ( .A1(n20094), .A2(n20939), .B1(n20145), .B2(n13360), .ZN(
        n13361) );
  OAI211_X1 U16486 ( .C1(n20667), .C2(n13409), .A(n13362), .B(n13361), .ZN(
        n13363) );
  AOI21_X1 U16487 ( .B1(n20140), .B2(n13364), .A(n13363), .ZN(n13365) );
  OAI21_X1 U16488 ( .B1(n20132), .B2(n13366), .A(n13365), .ZN(P1_U2839) );
  INV_X1 U16489 ( .A(n20541), .ZN(n13376) );
  NAND2_X1 U16490 ( .A1(n20239), .A2(n13367), .ZN(n13731) );
  INV_X1 U16491 ( .A(n20239), .ZN(n13728) );
  NOR2_X1 U16492 ( .A1(n13728), .A2(n20706), .ZN(n13727) );
  OR2_X1 U16493 ( .A1(n9665), .A2(n20736), .ZN(n20704) );
  NAND2_X1 U16494 ( .A1(n9665), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20636) );
  OAI22_X1 U16495 ( .A1(n20735), .A2(n20704), .B1(n20502), .B2(n20636), .ZN(
        n13373) );
  INV_X1 U16496 ( .A(n13368), .ZN(n13372) );
  AOI22_X1 U16497 ( .A1(n13373), .A2(n20637), .B1(n13371), .B2(n20736), .ZN(
        n13374) );
  AOI22_X1 U16498 ( .A1(n13727), .A2(n13374), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13728), .ZN(n13375) );
  OAI21_X1 U16499 ( .B1(n13376), .B2(n13731), .A(n13375), .ZN(P1_U3475) );
  OAI21_X1 U16500 ( .B1(n9763), .B2(n13377), .A(n13446), .ZN(n15537) );
  INV_X1 U16501 ( .A(n13380), .ZN(n13378) );
  INV_X1 U16502 ( .A(n13442), .ZN(n13441) );
  OAI211_X1 U16503 ( .C1(n10101), .C2(n13380), .A(n15012), .B(n13441), .ZN(
        n13382) );
  NAND2_X1 U16504 ( .A1(n15015), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13381) );
  OAI211_X1 U16505 ( .C1(n15537), .C2(n15004), .A(n13382), .B(n13381), .ZN(
        P2_U2875) );
  INV_X1 U16506 ( .A(n13383), .ZN(n13384) );
  AOI21_X1 U16507 ( .B1(n13386), .B2(n13385), .A(n13384), .ZN(n13402) );
  NAND2_X1 U16508 ( .A1(n13402), .A2(n20147), .ZN(n13395) );
  OAI21_X1 U16509 ( .B1(n20102), .B2(P1_REIP_REG_1__SCAN_IN), .A(n14232), .ZN(
        n20146) );
  INV_X1 U16510 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13404) );
  INV_X1 U16511 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20892) );
  NOR2_X1 U16512 ( .A1(n20102), .A2(n20939), .ZN(n20150) );
  AOI22_X1 U16513 ( .A1(n20139), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20892), .B2(n20150), .ZN(n13391) );
  OAI21_X1 U16514 ( .B1(n13389), .B2(n13388), .A(n13387), .ZN(n13403) );
  INV_X1 U16515 ( .A(n13403), .ZN(n20234) );
  NAND2_X1 U16516 ( .A1(n20145), .A2(n20234), .ZN(n13390) );
  OAI211_X1 U16517 ( .C1(n20117), .C2(n13404), .A(n13391), .B(n13390), .ZN(
        n13393) );
  NOR2_X1 U16518 ( .A1(n13162), .A2(n13409), .ZN(n13392) );
  AOI211_X1 U16519 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(n20146), .A(n13393), .B(
        n13392), .ZN(n13394) );
  OAI211_X1 U16520 ( .C1(n20098), .C2(n13399), .A(n13395), .B(n13394), .ZN(
        P1_U2838) );
  XNOR2_X1 U16521 ( .A(n13397), .B(n13396), .ZN(n20231) );
  AOI22_X1 U16522 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n16236), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13398) );
  OAI21_X1 U16523 ( .B1(n16135), .B2(n13399), .A(n13398), .ZN(n13400) );
  AOI21_X1 U16524 ( .B1(n13402), .B2(n16140), .A(n13400), .ZN(n13401) );
  OAI21_X1 U16525 ( .B1(n20063), .B2(n20231), .A(n13401), .ZN(P1_U2997) );
  INV_X1 U16526 ( .A(n13402), .ZN(n13405) );
  OAI222_X1 U16527 ( .A1(n13405), .A2(n16075), .B1(n20161), .B2(n13404), .C1(
        n13403), .C2(n16076), .ZN(P1_U2870) );
  OAI222_X1 U16528 ( .A1(n14396), .A2(n13405), .B1(n14389), .B2(n11191), .C1(
        n14394), .C2(n20269), .ZN(P1_U2902) );
  NAND2_X1 U16529 ( .A1(n20098), .A2(n20111), .ZN(n13412) );
  AOI22_X1 U16530 ( .A1(n13406), .A2(n20145), .B1(n20143), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13408) );
  NAND2_X1 U16531 ( .A1(n20102), .A2(n14232), .ZN(n16021) );
  NAND2_X1 U16532 ( .A1(n16021), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13407) );
  OAI211_X1 U16533 ( .C1(n13410), .C2(n13409), .A(n13408), .B(n13407), .ZN(
        n13411) );
  AOI21_X1 U16534 ( .B1(n13412), .B2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n13411), .ZN(n13413) );
  OAI21_X1 U16535 ( .B1(n20132), .B2(n13414), .A(n13413), .ZN(P1_U2840) );
  INV_X1 U16536 ( .A(n13415), .ZN(n20148) );
  AOI21_X1 U16537 ( .B1(n16128), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13416), .ZN(n13417) );
  OAI21_X1 U16538 ( .B1(n16135), .B2(n20138), .A(n13417), .ZN(n13418) );
  AOI21_X1 U16539 ( .B1(n20148), .B2(n16140), .A(n13418), .ZN(n13419) );
  OAI21_X1 U16540 ( .B1(n20063), .B2(n13420), .A(n13419), .ZN(P1_U2996) );
  AOI21_X1 U16541 ( .B1(n13423), .B2(n13304), .A(n13422), .ZN(n13510) );
  INV_X1 U16542 ( .A(n13510), .ZN(n14245) );
  INV_X1 U16543 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14233) );
  NAND2_X1 U16544 ( .A1(n14050), .A2(n14233), .ZN(n13427) );
  INV_X1 U16545 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14399) );
  NAND2_X1 U16546 ( .A1(n14008), .A2(n14399), .ZN(n13425) );
  NAND2_X1 U16547 ( .A1(n14043), .A2(n14233), .ZN(n13424) );
  NAND3_X1 U16548 ( .A1(n13425), .A2(n14053), .A3(n13424), .ZN(n13426) );
  AOI22_X1 U16549 ( .A1(n9767), .A2(n20156), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n14296), .ZN(n13430) );
  OAI21_X1 U16550 ( .B1(n14245), .B2(n16075), .A(n13430), .ZN(P1_U2868) );
  OR2_X1 U16551 ( .A1(n13422), .A2(n13432), .ZN(n13433) );
  NAND2_X1 U16552 ( .A1(n13431), .A2(n13433), .ZN(n20133) );
  INV_X1 U16553 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U16554 ( .A1(n14034), .A2(n13434), .ZN(n13438) );
  INV_X1 U16555 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16246) );
  NAND2_X1 U16556 ( .A1(n14043), .A2(n13434), .ZN(n13436) );
  OAI211_X1 U16557 ( .C1(n14073), .C2(n16246), .A(n13436), .B(n14008), .ZN(
        n13437) );
  OR2_X1 U16558 ( .A1(n16235), .A2(n9774), .ZN(n20129) );
  INV_X1 U16559 ( .A(n20129), .ZN(n16244) );
  AOI22_X1 U16560 ( .A1(n16244), .A2(n20156), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14296), .ZN(n13440) );
  OAI21_X1 U16561 ( .B1(n20133), .B2(n16075), .A(n13440), .ZN(P1_U2867) );
  INV_X1 U16562 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20180) );
  OAI222_X1 U16563 ( .A1(n14245), .A2(n14396), .B1(n20180), .B2(n14389), .C1(
        n14394), .C2(n20278), .ZN(P1_U2900) );
  INV_X1 U16564 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20178) );
  OAI222_X1 U16565 ( .A1(n14396), .A2(n20133), .B1(n14389), .B2(n20178), .C1(
        n14394), .C2(n20282), .ZN(P1_U2899) );
  INV_X1 U16566 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n19065) );
  INV_X1 U16567 ( .A(n13476), .ZN(n13443) );
  OAI211_X1 U16568 ( .C1(n13442), .C2(n13444), .A(n13443), .B(n15012), .ZN(
        n13450) );
  NAND2_X1 U16569 ( .A1(n13446), .A2(n13445), .ZN(n13447) );
  NAND2_X1 U16570 ( .A1(n13479), .A2(n13447), .ZN(n19069) );
  INV_X1 U16571 ( .A(n19069), .ZN(n13448) );
  NAND2_X1 U16572 ( .A1(n13448), .A2(n14998), .ZN(n13449) );
  OAI211_X1 U16573 ( .C1(n14998), .C2(n19065), .A(n13450), .B(n13449), .ZN(
        P2_U2874) );
  XNOR2_X1 U16574 ( .A(n13452), .B(n13613), .ZN(n13453) );
  XNOR2_X1 U16575 ( .A(n13451), .B(n13453), .ZN(n13475) );
  XNOR2_X1 U16576 ( .A(n13454), .B(n13455), .ZN(n13473) );
  OAI21_X1 U16577 ( .B1(n15458), .B2(n13746), .A(n13456), .ZN(n13612) );
  NOR2_X1 U16578 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15613), .ZN(
        n13457) );
  AOI22_X1 U16579 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13612), .B1(
        n13458), .B2(n13457), .ZN(n13464) );
  OAI21_X1 U16580 ( .B1(n13461), .B2(n13460), .A(n13459), .ZN(n20014) );
  INV_X1 U16581 ( .A(n20014), .ZN(n19257) );
  NAND2_X1 U16582 ( .A1(n19038), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13469) );
  INV_X1 U16583 ( .A(n13469), .ZN(n13462) );
  AOI21_X1 U16584 ( .B1(n19364), .B2(n19257), .A(n13462), .ZN(n13463) );
  OAI211_X1 U16585 ( .C1(n12941), .C2(n15589), .A(n13464), .B(n13463), .ZN(
        n13465) );
  AOI21_X1 U16586 ( .B1(n13473), .B2(n16361), .A(n13465), .ZN(n13466) );
  OAI21_X1 U16587 ( .B1(n13475), .B2(n15597), .A(n13466), .ZN(P2_U3043) );
  INV_X1 U16588 ( .A(n13727), .ZN(n13468) );
  XNOR2_X1 U16589 ( .A(n13368), .B(n20636), .ZN(n13467) );
  OAI222_X1 U16590 ( .A1(n13731), .A2(n13162), .B1(n20239), .B2(n20663), .C1(
        n13468), .C2(n13467), .ZN(P1_U3476) );
  OAI21_X1 U16591 ( .B1(n16359), .B2(n13525), .A(n13469), .ZN(n13470) );
  AOI21_X1 U16592 ( .B1(n16351), .B2(n13523), .A(n13470), .ZN(n13471) );
  OAI21_X1 U16593 ( .B1(n12941), .B2(n19376), .A(n13471), .ZN(n13472) );
  AOI21_X1 U16594 ( .B1(n13473), .B2(n19352), .A(n13472), .ZN(n13474) );
  OAI21_X1 U16595 ( .B1(n13475), .B2(n16324), .A(n13474), .ZN(P2_U3011) );
  OAI211_X1 U16596 ( .C1(n13476), .C2(n13477), .A(n13627), .B(n15012), .ZN(
        n13482) );
  INV_X1 U16597 ( .A(n13486), .ZN(n13478) );
  AOI21_X1 U16598 ( .B1(n13480), .B2(n13479), .A(n13478), .ZN(n19058) );
  NAND2_X1 U16599 ( .A1(n19058), .A2(n14998), .ZN(n13481) );
  OAI211_X1 U16600 ( .C1(n14998), .C2(n13483), .A(n13482), .B(n13481), .ZN(
        P2_U2873) );
  XNOR2_X1 U16601 ( .A(n13627), .B(n13626), .ZN(n13490) );
  AND2_X1 U16602 ( .A1(n13486), .A2(n13485), .ZN(n13487) );
  OR2_X1 U16603 ( .A1(n13487), .A2(n13644), .ZN(n15488) );
  NOR2_X1 U16604 ( .A1(n15488), .A2(n15004), .ZN(n13488) );
  AOI21_X1 U16605 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(n15004), .A(n13488), .ZN(
        n13489) );
  OAI21_X1 U16606 ( .B1(n13490), .B2(n15025), .A(n13489), .ZN(P2_U2872) );
  NAND2_X1 U16607 ( .A1(n13494), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13492) );
  NAND3_X1 U16608 ( .A1(n13493), .A2(n13492), .A3(n13491), .ZN(n13497) );
  INV_X1 U16609 ( .A(n13494), .ZN(n13495) );
  NAND2_X1 U16610 ( .A1(n13495), .A2(n13516), .ZN(n13496) );
  NAND2_X1 U16611 ( .A1(n13497), .A2(n13496), .ZN(n14400) );
  INV_X1 U16612 ( .A(n14429), .ZN(n14424) );
  NAND2_X1 U16613 ( .A1(n13498), .A2(n14424), .ZN(n13507) );
  NAND2_X1 U16614 ( .A1(n13500), .A2(n13499), .ZN(n13502) );
  INV_X1 U16615 ( .A(n13503), .ZN(n13501) );
  AOI21_X1 U16616 ( .B1(n13502), .B2(n13501), .A(n20954), .ZN(n13505) );
  INV_X1 U16617 ( .A(n13502), .ZN(n13504) );
  NAND2_X1 U16618 ( .A1(n13504), .A2(n13503), .ZN(n14411) );
  NAND2_X1 U16619 ( .A1(n13505), .A2(n14411), .ZN(n13506) );
  NAND2_X1 U16620 ( .A1(n13507), .A2(n13506), .ZN(n14397) );
  XOR2_X1 U16621 ( .A(n14398), .B(n14397), .Z(n13519) );
  INV_X1 U16622 ( .A(n13519), .ZN(n13512) );
  INV_X1 U16623 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n13590) );
  OR2_X1 U16624 ( .A1(n20227), .A2(n13590), .ZN(n13514) );
  NAND2_X1 U16625 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13508) );
  OAI211_X1 U16626 ( .C1(n16135), .C2(n14240), .A(n13514), .B(n13508), .ZN(
        n13509) );
  AOI21_X1 U16627 ( .B1(n13510), .B2(n16140), .A(n13509), .ZN(n13511) );
  OAI21_X1 U16628 ( .B1(n13512), .B2(n20063), .A(n13511), .ZN(P1_U2995) );
  INV_X1 U16629 ( .A(n9767), .ZN(n14236) );
  NAND2_X1 U16630 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13513), .ZN(
        n13515) );
  OAI211_X1 U16631 ( .C1(n16200), .C2(n14236), .A(n13515), .B(n13514), .ZN(
        n13518) );
  NOR2_X1 U16632 ( .A1(n14399), .A2(n13516), .ZN(n16216) );
  AOI211_X1 U16633 ( .C1(n14399), .C2(n13516), .A(n16216), .B(n16252), .ZN(
        n13517) );
  AOI211_X1 U16634 ( .C1(n16249), .C2(n13519), .A(n13518), .B(n13517), .ZN(
        n13520) );
  INV_X1 U16635 ( .A(n13520), .ZN(P1_U3027) );
  INV_X1 U16636 ( .A(n19196), .ZN(n19159) );
  NAND2_X1 U16637 ( .A1(n19145), .A2(n13521), .ZN(n13522) );
  XNOR2_X1 U16638 ( .A(n13523), .B(n13522), .ZN(n13524) );
  INV_X1 U16639 ( .A(n19929), .ZN(n19178) );
  NAND2_X1 U16640 ( .A1(n13524), .A2(n19178), .ZN(n13533) );
  INV_X1 U16641 ( .A(n12941), .ZN(n13531) );
  OAI22_X1 U16642 ( .A1(n13525), .A2(n19097), .B1(n19154), .B2(n20014), .ZN(
        n13527) );
  NOR2_X1 U16643 ( .A1(n19188), .A2(n10658), .ZN(n13526) );
  AOI211_X1 U16644 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19183), .A(n13527), .B(
        n13526), .ZN(n13528) );
  OAI21_X1 U16645 ( .B1(n13529), .B2(n19194), .A(n13528), .ZN(n13530) );
  AOI21_X1 U16646 ( .B1(n13531), .B2(n19190), .A(n13530), .ZN(n13532) );
  OAI211_X1 U16647 ( .C1(n19159), .C2(n19630), .A(n13533), .B(n13532), .ZN(
        P2_U2852) );
  INV_X1 U16648 ( .A(n13535), .ZN(n13536) );
  AOI21_X1 U16649 ( .B1(n13537), .B2(n13431), .A(n13536), .ZN(n20158) );
  INV_X1 U16650 ( .A(n20158), .ZN(n13538) );
  OAI222_X1 U16651 ( .A1(n14396), .A2(n13538), .B1(n14389), .B2(n11334), .C1(
        n14394), .C2(n20287), .ZN(P1_U2898) );
  AOI21_X1 U16652 ( .B1(n13540), .B2(n13535), .A(n13539), .ZN(n16125) );
  INV_X1 U16653 ( .A(n16125), .ZN(n20105) );
  MUX2_X1 U16654 ( .A(n14048), .B(n14053), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n13541) );
  NAND2_X1 U16655 ( .A1(n13541), .A2(n10225), .ZN(n13550) );
  INV_X1 U16656 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20160) );
  NAND2_X1 U16657 ( .A1(n14050), .A2(n20160), .ZN(n13545) );
  INV_X1 U16658 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16225) );
  NAND2_X1 U16659 ( .A1(n14008), .A2(n16225), .ZN(n13543) );
  NAND2_X1 U16660 ( .A1(n14043), .A2(n20160), .ZN(n13542) );
  NAND3_X1 U16661 ( .A1(n13543), .A2(n14053), .A3(n13542), .ZN(n13544) );
  INV_X1 U16662 ( .A(n16234), .ZN(n13546) );
  NAND2_X1 U16663 ( .A1(n16235), .A2(n13546), .ZN(n13549) );
  NOR2_X1 U16664 ( .A1(n13550), .A2(n16234), .ZN(n13547) );
  INV_X1 U16665 ( .A(n13587), .ZN(n13548) );
  AOI21_X1 U16666 ( .B1(n13550), .B2(n13549), .A(n13548), .ZN(n20108) );
  AOI22_X1 U16667 ( .A1(n20108), .A2(n20156), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14296), .ZN(n13551) );
  OAI21_X1 U16668 ( .B1(n20105), .B2(n16075), .A(n13551), .ZN(P1_U2865) );
  OAI222_X1 U16669 ( .A1(n14396), .A2(n20105), .B1(n14389), .B2(n11346), .C1(
        n14394), .C2(n20296), .ZN(P1_U2897) );
  NOR2_X1 U16670 ( .A1(n19162), .A2(n13552), .ZN(n13553) );
  XNOR2_X1 U16671 ( .A(n13553), .B(n16345), .ZN(n13554) );
  NAND2_X1 U16672 ( .A1(n13554), .A2(n19178), .ZN(n13566) );
  INV_X1 U16673 ( .A(n13555), .ZN(n13559) );
  INV_X1 U16674 ( .A(n15582), .ZN(n13558) );
  AOI21_X1 U16675 ( .B1(n13559), .B2(n13556), .A(n13558), .ZN(n19236) );
  AOI22_X1 U16676 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n19183), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19198), .ZN(n13560) );
  OAI211_X1 U16677 ( .C1(n19188), .C2(n13561), .A(n13560), .B(n19129), .ZN(
        n13564) );
  NOR2_X1 U16678 ( .A1(n13562), .A2(n19174), .ZN(n13563) );
  AOI211_X1 U16679 ( .C1(n19185), .C2(n19236), .A(n13564), .B(n13563), .ZN(
        n13565) );
  OAI211_X1 U16680 ( .C1(n19194), .C2(n13567), .A(n13566), .B(n13565), .ZN(
        P2_U2847) );
  NOR2_X1 U16681 ( .A1(n19162), .A2(n13718), .ZN(n13568) );
  XNOR2_X1 U16682 ( .A(n13568), .B(n13740), .ZN(n13569) );
  NAND2_X1 U16683 ( .A1(n13569), .A2(n19178), .ZN(n13577) );
  NAND2_X1 U16684 ( .A1(n20021), .A2(n19185), .ZN(n13573) );
  INV_X1 U16685 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13737) );
  OAI22_X1 U16686 ( .A1(n13737), .A2(n19097), .B1(n10458), .B2(n19188), .ZN(
        n13570) );
  AOI21_X1 U16687 ( .B1(n19153), .B2(n13571), .A(n13570), .ZN(n13572) );
  OAI211_X1 U16688 ( .C1(n13574), .C2(n19156), .A(n13573), .B(n13572), .ZN(
        n13575) );
  AOI21_X1 U16689 ( .B1(n12060), .B2(n19190), .A(n13575), .ZN(n13576) );
  OAI211_X1 U16690 ( .C1(n20019), .C2(n19159), .A(n13577), .B(n13576), .ZN(
        P2_U2853) );
  INV_X1 U16691 ( .A(n13578), .ZN(n13579) );
  OAI21_X1 U16692 ( .B1(n13539), .B2(n13580), .A(n13579), .ZN(n14631) );
  INV_X1 U16693 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13581) );
  NAND2_X1 U16694 ( .A1(n14050), .A2(n13581), .ZN(n13585) );
  INV_X1 U16695 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16228) );
  NAND2_X1 U16696 ( .A1(n14008), .A2(n16228), .ZN(n13583) );
  NAND2_X1 U16697 ( .A1(n14043), .A2(n13581), .ZN(n13582) );
  NAND3_X1 U16698 ( .A1(n13583), .A2(n14053), .A3(n13582), .ZN(n13584) );
  INV_X1 U16699 ( .A(n13604), .ZN(n13586) );
  AOI21_X1 U16700 ( .B1(n13588), .B2(n13587), .A(n13586), .ZN(n16224) );
  AOI22_X1 U16701 ( .A1(n16224), .A2(n20156), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14296), .ZN(n13589) );
  OAI21_X1 U16702 ( .B1(n14631), .B2(n16075), .A(n13589), .ZN(P1_U2864) );
  INV_X1 U16703 ( .A(n14232), .ZN(n13591) );
  NAND3_X1 U16704 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n14241) );
  NOR2_X1 U16705 ( .A1(n13590), .A2(n14241), .ZN(n20093) );
  INV_X1 U16706 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20898) );
  NAND2_X1 U16707 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20100) );
  NOR2_X1 U16708 ( .A1(n20898), .A2(n20100), .ZN(n13593) );
  NAND3_X1 U16709 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20093), .A3(n13593), 
        .ZN(n20083) );
  NOR2_X1 U16710 ( .A1(n13591), .A2(n20083), .ZN(n14181) );
  INV_X1 U16711 ( .A(n16021), .ZN(n14184) );
  NOR2_X1 U16712 ( .A1(n14181), .A2(n14184), .ZN(n20087) );
  AOI22_X1 U16713 ( .A1(n14634), .A2(n20140), .B1(n20145), .B2(n16224), .ZN(
        n13596) );
  AOI22_X1 U16714 ( .A1(n20143), .A2(P1_EBX_REG_8__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20139), .ZN(n13595) );
  INV_X1 U16715 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13592) );
  NAND4_X1 U16716 ( .A1(n20094), .A2(n20093), .A3(n13593), .A4(n13592), .ZN(
        n13594) );
  NAND4_X1 U16717 ( .A1(n13596), .A2(n13595), .A3(n20227), .A4(n13594), .ZN(
        n13597) );
  AOI21_X1 U16718 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n20087), .A(n13597), .ZN(
        n13598) );
  OAI21_X1 U16719 ( .B1(n14631), .B2(n20104), .A(n13598), .ZN(P1_U2832) );
  OR2_X1 U16720 ( .A1(n13578), .A2(n13600), .ZN(n13601) );
  NAND2_X1 U16721 ( .A1(n13599), .A2(n13601), .ZN(n20086) );
  MUX2_X1 U16722 ( .A(n14048), .B(n14053), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n13602) );
  NAND2_X1 U16723 ( .A1(n13602), .A2(n10227), .ZN(n13603) );
  AND2_X1 U16724 ( .A1(n13604), .A2(n13603), .ZN(n13605) );
  NOR2_X1 U16725 ( .A1(n14224), .A2(n13605), .ZN(n20082) );
  AOI22_X1 U16726 ( .A1(n20082), .A2(n20156), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14296), .ZN(n13606) );
  OAI21_X1 U16727 ( .B1(n20086), .B2(n16075), .A(n13606), .ZN(P1_U2863) );
  NAND2_X1 U16728 ( .A1(n13607), .A2(n13608), .ZN(n13609) );
  XNOR2_X1 U16729 ( .A(n13609), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19353) );
  INV_X1 U16730 ( .A(n19353), .ZN(n13621) );
  XOR2_X1 U16731 ( .A(n13611), .B(n13610), .Z(n19354) );
  AOI21_X1 U16732 ( .B1(n19370), .B2(n13613), .A(n13612), .ZN(n15611) );
  NAND2_X1 U16733 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19348), .ZN(n13614) );
  OAI221_X1 U16734 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15617), .C1(
        n13656), .C2(n15611), .A(n13614), .ZN(n13619) );
  NAND2_X1 U16735 ( .A1(n13615), .A2(n13459), .ZN(n13617) );
  INV_X1 U16736 ( .A(n13658), .ZN(n13616) );
  NAND2_X1 U16737 ( .A1(n13617), .A2(n13616), .ZN(n19250) );
  OAI22_X1 U16738 ( .A1(n19158), .A2(n15589), .B1(n16371), .B2(n19250), .ZN(
        n13618) );
  AOI211_X1 U16739 ( .C1(n19354), .C2(n19361), .A(n13619), .B(n13618), .ZN(
        n13620) );
  OAI21_X1 U16740 ( .B1(n19366), .B2(n13621), .A(n13620), .ZN(P2_U3042) );
  INV_X1 U16741 ( .A(DATAI_9_), .ZN(n13623) );
  MUX2_X1 U16742 ( .A(n13623), .B(n13622), .S(n20241), .Z(n20191) );
  OAI222_X1 U16743 ( .A1(n20086), .A2(n14396), .B1(n20173), .B2(n14389), .C1(
        n14394), .C2(n20191), .ZN(P1_U2895) );
  INV_X1 U16744 ( .A(DATAI_8_), .ZN(n13624) );
  MUX2_X1 U16745 ( .A(n13624), .B(n16551), .S(n20241), .Z(n20188) );
  OAI222_X1 U16746 ( .A1(n14631), .A2(n14396), .B1(n13625), .B2(n14389), .C1(
        n14394), .C2(n20188), .ZN(P1_U2896) );
  AOI22_X1 U16747 ( .A1(n10694), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13631) );
  AOI22_X1 U16748 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10675), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13630) );
  AOI22_X1 U16749 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13629) );
  AOI22_X1 U16750 ( .A1(n10623), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13628) );
  NAND4_X1 U16751 ( .A1(n13631), .A2(n13630), .A3(n13629), .A4(n13628), .ZN(
        n13637) );
  AOI22_X1 U16752 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13834), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13635) );
  AOI22_X1 U16753 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13634) );
  AOI22_X1 U16754 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13633) );
  AOI22_X1 U16755 ( .A1(n13836), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13632) );
  NAND4_X1 U16756 ( .A1(n13635), .A2(n13634), .A3(n13633), .A4(n13632), .ZN(
        n13636) );
  NOR2_X1 U16757 ( .A1(n13637), .A2(n13636), .ZN(n13640) );
  INV_X1 U16758 ( .A(n13640), .ZN(n13638) );
  INV_X1 U16759 ( .A(n13639), .ZN(n13641) );
  AND2_X1 U16760 ( .A1(n13641), .A2(n13640), .ZN(n13642) );
  NOR2_X1 U16761 ( .A1(n13765), .A2(n13642), .ZN(n19211) );
  NAND2_X1 U16762 ( .A1(n19211), .A2(n15012), .ZN(n13647) );
  OR2_X1 U16763 ( .A1(n13644), .A2(n13643), .ZN(n13645) );
  AND2_X1 U16764 ( .A1(n13645), .A2(n15020), .ZN(n15477) );
  NAND2_X1 U16765 ( .A1(n15477), .A2(n14998), .ZN(n13646) );
  OAI211_X1 U16766 ( .C1(n14998), .C2(n13648), .A(n13647), .B(n13646), .ZN(
        P2_U2871) );
  XNOR2_X1 U16767 ( .A(n13649), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13650) );
  XNOR2_X1 U16768 ( .A(n13651), .B(n13650), .ZN(n16353) );
  INV_X1 U16769 ( .A(n16353), .ZN(n13666) );
  NAND2_X1 U16770 ( .A1(n13654), .A2(n13652), .ZN(n13653) );
  AOI22_X1 U16771 ( .A1(n13655), .A2(n13654), .B1(n9795), .B2(n13653), .ZN(
        n16352) );
  AOI211_X1 U16772 ( .C1(n13662), .C2(n13656), .A(n15605), .B(n15617), .ZN(
        n13664) );
  XNOR2_X1 U16773 ( .A(n13658), .B(n13657), .ZN(n19248) );
  OAI22_X1 U16774 ( .A1(n16371), .A2(n19248), .B1(n19129), .B2(n13659), .ZN(
        n13660) );
  AOI21_X1 U16775 ( .B1(n19369), .B2(n19148), .A(n13660), .ZN(n13661) );
  OAI21_X1 U16776 ( .B1(n15611), .B2(n13662), .A(n13661), .ZN(n13663) );
  AOI211_X1 U16777 ( .C1(n16352), .C2(n16361), .A(n13664), .B(n13663), .ZN(
        n13665) );
  OAI21_X1 U16778 ( .B1(n13666), .B2(n15597), .A(n13665), .ZN(P2_U3041) );
  INV_X1 U16779 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17057) );
  AND2_X1 U16780 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n15722) );
  INV_X1 U16781 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16723) );
  INV_X1 U16782 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17075) );
  INV_X1 U16783 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16756) );
  INV_X1 U16784 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17116) );
  NOR4_X1 U16785 ( .A1(n16723), .A2(n17075), .A3(n16756), .A4(n17116), .ZN(
        n13667) );
  NAND4_X1 U16786 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n15722), .A4(n13667), .ZN(n17064) );
  INV_X1 U16787 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17134) );
  INV_X1 U16788 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16813) );
  INV_X1 U16789 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16838) );
  INV_X1 U16790 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17217) );
  NAND2_X1 U16791 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .ZN(n17201) );
  NAND4_X1 U16792 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(P3_EBX_REG_9__SCAN_IN), .ZN(n13668)
         );
  NOR4_X1 U16793 ( .A1(n16838), .A2(n17217), .A3(n17201), .A4(n13668), .ZN(
        n17149) );
  NAND2_X1 U16794 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17150), .ZN(n17133) );
  NAND2_X1 U16795 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17147), .ZN(n17115) );
  NOR3_X1 U16796 ( .A1(n17057), .A2(n17064), .A3(n17115), .ZN(n17054) );
  NAND2_X1 U16797 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17054), .ZN(n13669) );
  NOR2_X1 U16798 ( .A1(n17404), .A2(n13669), .ZN(n13671) );
  INV_X2 U16799 ( .A(n17311), .ZN(n17305) );
  NAND2_X1 U16800 ( .A1(n17305), .A2(n13669), .ZN(n17055) );
  INV_X1 U16801 ( .A(n17055), .ZN(n13670) );
  MUX2_X1 U16802 ( .A(n13671), .B(n13670), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  NOR2_X1 U16803 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18898) );
  INV_X1 U16804 ( .A(n18898), .ZN(n18904) );
  INV_X1 U16805 ( .A(n18293), .ZN(n13672) );
  NAND2_X1 U16806 ( .A1(n18277), .A2(n17404), .ZN(n13685) );
  NAND2_X1 U16807 ( .A1(n13673), .A2(n17317), .ZN(n13677) );
  NOR3_X1 U16808 ( .A1(n18726), .A2(n13697), .A3(n15864), .ZN(n13679) );
  INV_X1 U16809 ( .A(n13673), .ZN(n18297) );
  NOR2_X1 U16810 ( .A1(n18297), .A2(n15864), .ZN(n15899) );
  NOR2_X1 U16811 ( .A1(n18277), .A2(n18929), .ZN(n13674) );
  NAND2_X1 U16812 ( .A1(n17404), .A2(n18744), .ZN(n15983) );
  NAND2_X1 U16813 ( .A1(n13674), .A2(n15983), .ZN(n13701) );
  OAI21_X1 U16814 ( .B1(n13679), .B2(n15899), .A(n13701), .ZN(n13682) );
  NAND2_X1 U16815 ( .A1(n18744), .A2(n18293), .ZN(n13687) );
  NOR2_X1 U16816 ( .A1(n18307), .A2(n18293), .ZN(n13675) );
  NAND2_X1 U16817 ( .A1(n13677), .A2(n13675), .ZN(n13678) );
  INV_X1 U16818 ( .A(n15864), .ZN(n18285) );
  NAND2_X1 U16819 ( .A1(n18277), .A2(n18929), .ZN(n13676) );
  NAND2_X1 U16820 ( .A1(n18285), .A2(n13676), .ZN(n13695) );
  AOI22_X1 U16821 ( .A1(n13687), .A2(n13678), .B1(n13677), .B2(n13695), .ZN(
        n13681) );
  AOI22_X1 U16822 ( .A1(n18277), .A2(n13679), .B1(n18289), .B2(n13685), .ZN(
        n13680) );
  NAND2_X1 U16823 ( .A1(n13681), .A2(n13680), .ZN(n13700) );
  AOI21_X1 U16824 ( .B1(n13683), .B2(n13682), .A(n13700), .ZN(n15744) );
  NAND2_X1 U16825 ( .A1(n13688), .A2(n15744), .ZN(n15747) );
  INV_X1 U16826 ( .A(n15747), .ZN(n18730) );
  NAND2_X1 U16827 ( .A1(n13688), .A2(n15864), .ZN(n13699) );
  OAI21_X1 U16828 ( .B1(n18731), .B2(n18883), .A(n18721), .ZN(n13708) );
  NAND2_X1 U16829 ( .A1(n10213), .A2(n13708), .ZN(n18719) );
  NOR2_X1 U16830 ( .A1(n18904), .A2(n18719), .ZN(n13707) );
  NAND2_X1 U16831 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18794) );
  XOR2_X1 U16832 ( .A(n13691), .B(n13690), .Z(n13693) );
  NOR2_X1 U16833 ( .A1(n9890), .A2(n9891), .ZN(n13703) );
  INV_X1 U16834 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18787) );
  AOI21_X1 U16835 ( .B1(n18807), .B2(n18787), .A(P3_STATE_REG_0__SCAN_IN), 
        .ZN(n18799) );
  NAND2_X1 U16836 ( .A1(n18804), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18940) );
  NOR2_X1 U16837 ( .A1(n18807), .A2(n18940), .ZN(n18795) );
  INV_X2 U16838 ( .A(n18795), .ZN(n18867) );
  NAND2_X1 U16839 ( .A1(n18799), .A2(n18867), .ZN(n16635) );
  INV_X1 U16840 ( .A(n16635), .ZN(n18928) );
  INV_X1 U16841 ( .A(n18744), .ZN(n15984) );
  NOR3_X1 U16842 ( .A1(n13697), .A2(n13696), .A3(n13695), .ZN(n13698) );
  OAI21_X1 U16843 ( .B1(n18293), .B2(n15984), .A(n13698), .ZN(n15865) );
  OAI21_X1 U16844 ( .B1(n15865), .B2(n13700), .A(n13699), .ZN(n13702) );
  NAND2_X1 U16845 ( .A1(n13702), .A2(n13701), .ZN(n15897) );
  AOI21_X1 U16846 ( .B1(n13703), .B2(n17473), .A(n15897), .ZN(n13705) );
  OAI211_X1 U16847 ( .C1(n15741), .C2(n18717), .A(n13705), .B(n15981), .ZN(
        n18752) );
  INV_X1 U16848 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18878) );
  NOR2_X1 U16849 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18878), .ZN(n18276) );
  INV_X1 U16850 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16619) );
  NOR2_X1 U16851 ( .A1(n18905), .A2(n18932), .ZN(n18782) );
  NAND2_X1 U16852 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18782), .ZN(n18876) );
  NOR2_X1 U16853 ( .A1(n16619), .A2(n18876), .ZN(n13706) );
  AOI211_X2 U16854 ( .C1(n18771), .C2(n18752), .A(n18276), .B(n13706), .ZN(
        n18910) );
  MUX2_X1 U16855 ( .A(n13707), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18910), .Z(P3_U3284) );
  NOR2_X1 U16856 ( .A1(n9657), .A2(n13708), .ZN(n18260) );
  INV_X1 U16857 ( .A(n18897), .ZN(n18902) );
  OAI221_X1 U16858 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18905), .C1(n18930), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n18902), .ZN(n18275) );
  OAI221_X1 U16859 ( .B1(n18876), .B2(n18260), .C1(n18876), .C2(n16619), .A(
        n18372), .ZN(n18267) );
  INV_X1 U16860 ( .A(n18267), .ZN(n18262) );
  OAI21_X1 U16861 ( .B1(n18905), .B2(n18930), .A(n18878), .ZN(n16434) );
  INV_X1 U16862 ( .A(n16434), .ZN(n18924) );
  NAND2_X1 U16863 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17897) );
  AOI22_X1 U16864 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .B1(n18924), .B2(n17897), .ZN(n15739) );
  NOR2_X1 U16865 ( .A1(n18262), .A2(n15739), .ZN(n13710) );
  NAND2_X1 U16866 ( .A1(n18930), .A2(n18878), .ZN(n16613) );
  NOR2_X1 U16867 ( .A1(n16613), .A2(n16638), .ZN(n18330) );
  INV_X1 U16868 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18271) );
  NAND2_X1 U16869 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18271), .ZN(n18311) );
  NAND2_X1 U16870 ( .A1(n18311), .A2(n18267), .ZN(n15737) );
  OR2_X1 U16871 ( .A1(n18330), .A2(n15737), .ZN(n13709) );
  MUX2_X1 U16872 ( .A(n13710), .B(n13709), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U16873 ( .A(n13711), .ZN(n13712) );
  NOR2_X1 U16874 ( .A1(n12456), .A2(n13712), .ZN(n15621) );
  XNOR2_X1 U16875 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13715) );
  NAND2_X1 U16876 ( .A1(n13058), .A2(n13713), .ZN(n13714) );
  OAI21_X1 U16877 ( .B1(n15621), .B2(n13715), .A(n13714), .ZN(n13716) );
  AOI21_X1 U16878 ( .B1(n12728), .B2(n13717), .A(n13716), .ZN(n16400) );
  NAND2_X1 U16879 ( .A1(n20028), .A2(n16421), .ZN(n13724) );
  AOI211_X1 U16880 ( .C1(n13720), .C2(n13719), .A(n19162), .B(n13718), .ZN(
        n19179) );
  AOI21_X1 U16881 ( .B1(n19162), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19179), .ZN(n15642) );
  NAND2_X1 U16882 ( .A1(n19145), .A2(n13720), .ZN(n19201) );
  OAI21_X1 U16883 ( .B1(n19145), .B2(n13721), .A(n19201), .ZN(n15628) );
  NAND2_X1 U16884 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15628), .ZN(n15641) );
  INV_X1 U16885 ( .A(n15641), .ZN(n13722) );
  NAND2_X1 U16886 ( .A1(n15642), .A2(n13722), .ZN(n13723) );
  OAI211_X1 U16887 ( .C1(n20008), .C2(n16400), .A(n13724), .B(n13723), .ZN(
        n13726) );
  MUX2_X1 U16888 ( .A(n13726), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n13725), .Z(P2_U3600) );
  OAI211_X1 U16889 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n9665), .A(n13727), 
        .B(n20636), .ZN(n13730) );
  NAND2_X1 U16890 ( .A1(n13728), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13729) );
  OAI211_X1 U16891 ( .C1(n13731), .C2(n20667), .A(n13730), .B(n13729), .ZN(
        P1_U3477) );
  XOR2_X1 U16892 ( .A(n13733), .B(n13732), .Z(n13752) );
  INV_X1 U16893 ( .A(n13734), .ZN(n13735) );
  XNOR2_X1 U16894 ( .A(n13736), .B(n13735), .ZN(n13744) );
  NAND2_X1 U16895 ( .A1(n19038), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13748) );
  OAI21_X1 U16896 ( .B1(n16359), .B2(n13737), .A(n13748), .ZN(n13738) );
  AOI21_X1 U16897 ( .B1(n19352), .B2(n13744), .A(n13738), .ZN(n13739) );
  OAI21_X1 U16898 ( .B1(n13740), .B2(n19359), .A(n13739), .ZN(n13741) );
  AOI21_X1 U16899 ( .B1(n13752), .B2(n19355), .A(n13741), .ZN(n13742) );
  OAI21_X1 U16900 ( .B1(n15636), .B2(n19376), .A(n13742), .ZN(P2_U3012) );
  AOI21_X1 U16901 ( .B1(n13745), .B2(n13746), .A(n15458), .ZN(n13743) );
  INV_X1 U16902 ( .A(n13743), .ZN(n13754) );
  AOI22_X1 U16903 ( .A1(n13744), .A2(n16361), .B1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19362), .ZN(n13750) );
  NAND2_X1 U16904 ( .A1(n20021), .A2(n19364), .ZN(n13749) );
  NAND3_X1 U16905 ( .A1(n15461), .A2(n13746), .A3(n13745), .ZN(n13747) );
  NAND4_X1 U16906 ( .A1(n13750), .A2(n13749), .A3(n13748), .A4(n13747), .ZN(
        n13751) );
  AOI21_X1 U16907 ( .B1(n13752), .B2(n19361), .A(n13751), .ZN(n13753) );
  OAI211_X1 U16908 ( .C1(n15589), .C2(n15636), .A(n13754), .B(n13753), .ZN(
        P2_U3044) );
  AOI22_X1 U16909 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10693), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13758) );
  AOI22_X1 U16910 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13757) );
  AOI22_X1 U16911 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13756) );
  AOI22_X1 U16912 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13755) );
  NAND4_X1 U16913 ( .A1(n13758), .A2(n13757), .A3(n13756), .A4(n13755), .ZN(
        n13764) );
  AOI22_X1 U16914 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n13834), .ZN(n13762) );
  AOI22_X1 U16915 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U16916 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13760) );
  AOI22_X1 U16917 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13759) );
  NAND4_X1 U16918 ( .A1(n13762), .A2(n13761), .A3(n13760), .A4(n13759), .ZN(
        n13763) );
  OR2_X1 U16919 ( .A1(n13764), .A2(n13763), .ZN(n15018) );
  AOI22_X1 U16920 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10693), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13769) );
  AOI22_X1 U16921 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13768) );
  AOI22_X1 U16922 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13767) );
  AOI22_X1 U16923 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13766) );
  NAND4_X1 U16924 ( .A1(n13769), .A2(n13768), .A3(n13767), .A4(n13766), .ZN(
        n13775) );
  AOI22_X1 U16925 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n13834), .ZN(n13773) );
  AOI22_X1 U16926 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13772) );
  AOI22_X1 U16927 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13771) );
  AOI22_X1 U16928 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13770) );
  NAND4_X1 U16929 ( .A1(n13773), .A2(n13772), .A3(n13771), .A4(n13770), .ZN(
        n13774) );
  OR2_X1 U16930 ( .A1(n13775), .A2(n13774), .ZN(n15000) );
  AOI22_X1 U16931 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10693), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13779) );
  AOI22_X1 U16932 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13778) );
  AOI22_X1 U16933 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13777) );
  AOI22_X1 U16934 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13776) );
  NAND4_X1 U16935 ( .A1(n13779), .A2(n13778), .A3(n13777), .A4(n13776), .ZN(
        n13785) );
  AOI22_X1 U16936 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n13834), .ZN(n13783) );
  AOI22_X1 U16937 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13782) );
  AOI22_X1 U16938 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13781) );
  AOI22_X1 U16939 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13780) );
  NAND4_X1 U16940 ( .A1(n13783), .A2(n13782), .A3(n13781), .A4(n13780), .ZN(
        n13784) );
  OR2_X1 U16941 ( .A1(n13785), .A2(n13784), .ZN(n15009) );
  AND2_X1 U16942 ( .A1(n15000), .A2(n15009), .ZN(n13786) );
  AOI22_X1 U16943 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10693), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13790) );
  AOI22_X1 U16944 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13789) );
  AOI22_X1 U16945 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U16946 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13787) );
  NAND4_X1 U16947 ( .A1(n13790), .A2(n13789), .A3(n13788), .A4(n13787), .ZN(
        n13796) );
  AOI22_X1 U16948 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n13834), .ZN(n13794) );
  AOI22_X1 U16949 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13793) );
  AOI22_X1 U16950 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13792) );
  AOI22_X1 U16951 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13791) );
  NAND4_X1 U16952 ( .A1(n13794), .A2(n13793), .A3(n13792), .A4(n13791), .ZN(
        n13795) );
  NOR2_X1 U16953 ( .A1(n13796), .A2(n13795), .ZN(n14990) );
  AOI22_X1 U16954 ( .A1(n10694), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13800) );
  AOI22_X1 U16955 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10675), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13799) );
  AOI22_X1 U16956 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U16957 ( .A1(n10623), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13797) );
  NAND4_X1 U16958 ( .A1(n13800), .A2(n13799), .A3(n13798), .A4(n13797), .ZN(
        n13806) );
  AOI22_X1 U16959 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13834), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13804) );
  AOI22_X1 U16960 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13803) );
  AOI22_X1 U16961 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U16962 ( .A1(n13836), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13801) );
  NAND4_X1 U16963 ( .A1(n13804), .A2(n13803), .A3(n13802), .A4(n13801), .ZN(
        n13805) );
  OR2_X1 U16964 ( .A1(n13806), .A2(n13805), .ZN(n14984) );
  AOI22_X1 U16965 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10693), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U16966 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10675), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13809) );
  AOI22_X1 U16967 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U16968 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13807) );
  NAND4_X1 U16969 ( .A1(n13810), .A2(n13809), .A3(n13808), .A4(n13807), .ZN(
        n13817) );
  AOI22_X1 U16970 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n13834), .ZN(n13815) );
  AOI22_X1 U16971 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13814) );
  AOI22_X1 U16972 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13813) );
  AOI22_X1 U16973 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n13836), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13812) );
  NAND4_X1 U16974 ( .A1(n13815), .A2(n13814), .A3(n13813), .A4(n13812), .ZN(
        n13816) );
  NOR2_X1 U16975 ( .A1(n13817), .A2(n13816), .ZN(n14980) );
  AOI22_X1 U16976 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13819) );
  AOI22_X1 U16977 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13818) );
  AND2_X1 U16978 ( .A1(n13819), .A2(n13818), .ZN(n13822) );
  AOI22_X1 U16979 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13821) );
  AOI22_X1 U16980 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9666), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13820) );
  XNOR2_X1 U16981 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13965) );
  NAND4_X1 U16982 ( .A1(n13822), .A2(n13821), .A3(n13820), .A4(n13965), .ZN(
        n13829) );
  AOI22_X1 U16983 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13824) );
  AOI22_X1 U16984 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13823) );
  AND2_X1 U16985 ( .A1(n13824), .A2(n13823), .ZN(n13827) );
  INV_X1 U16986 ( .A(n13965), .ZN(n13973) );
  AOI22_X1 U16987 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9655), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13826) );
  AOI22_X1 U16988 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13825) );
  NAND4_X1 U16989 ( .A1(n13827), .A2(n13973), .A3(n13826), .A4(n13825), .ZN(
        n13828) );
  AND2_X1 U16990 ( .A1(n13829), .A2(n13828), .ZN(n13865) );
  NAND2_X1 U16991 ( .A1(n13865), .A2(n10598), .ZN(n13846) );
  AOI22_X1 U16992 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10663), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U16993 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10693), .B1(
        n10675), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13832) );
  AOI22_X1 U16994 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10602), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13831) );
  AOI22_X1 U16995 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10623), .B1(
        n10638), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13830) );
  NAND4_X1 U16996 ( .A1(n13833), .A2(n13832), .A3(n13831), .A4(n13830), .ZN(
        n13845) );
  AOI22_X1 U16997 ( .A1(n13835), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n13834), .ZN(n13843) );
  AOI22_X1 U16998 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n13836), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13842) );
  AOI22_X1 U16999 ( .A1(n13811), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13841) );
  AOI22_X1 U17000 ( .A1(n13839), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13840) );
  NAND4_X1 U17001 ( .A1(n13843), .A2(n13842), .A3(n13841), .A4(n13840), .ZN(
        n13844) );
  OR2_X1 U17002 ( .A1(n13845), .A2(n13844), .ZN(n13862) );
  XNOR2_X1 U17003 ( .A(n13846), .B(n13862), .ZN(n13868) );
  NAND2_X1 U17004 ( .A1(n10406), .A2(n13865), .ZN(n14974) );
  AOI22_X1 U17005 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U17006 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13849) );
  AND2_X1 U17007 ( .A1(n13850), .A2(n13849), .ZN(n13853) );
  AOI22_X1 U17008 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13875), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13852) );
  AOI22_X1 U17009 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(n9666), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13851) );
  NAND4_X1 U17010 ( .A1(n13853), .A2(n13852), .A3(n13851), .A4(n13965), .ZN(
        n13861) );
  AOI22_X1 U17011 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13856) );
  AOI22_X1 U17012 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13855) );
  AND2_X1 U17013 ( .A1(n13856), .A2(n13855), .ZN(n13859) );
  AOI22_X1 U17014 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9655), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13858) );
  AOI22_X1 U17015 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13857) );
  NAND4_X1 U17016 ( .A1(n13859), .A2(n13973), .A3(n13858), .A4(n13857), .ZN(
        n13860) );
  NAND2_X1 U17017 ( .A1(n13861), .A2(n13860), .ZN(n13871) );
  NAND2_X1 U17018 ( .A1(n13862), .A2(n13865), .ZN(n13872) );
  XOR2_X1 U17019 ( .A(n13871), .B(n13872), .Z(n13863) );
  NAND2_X1 U17020 ( .A1(n13863), .A2(n13924), .ZN(n14965) );
  INV_X1 U17021 ( .A(n13871), .ZN(n13864) );
  NAND2_X1 U17022 ( .A1(n10406), .A2(n13864), .ZN(n14967) );
  INV_X1 U17023 ( .A(n13865), .ZN(n13866) );
  NOR2_X1 U17024 ( .A1(n14967), .A2(n13866), .ZN(n13867) );
  NAND2_X1 U17025 ( .A1(n13868), .A2(n13867), .ZN(n13869) );
  NOR2_X1 U17026 ( .A1(n13872), .A2(n13871), .ZN(n13886) );
  AOI22_X1 U17027 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13964), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13874) );
  AOI22_X1 U17028 ( .A1(n13972), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13873) );
  AND2_X1 U17029 ( .A1(n13874), .A2(n13873), .ZN(n13878) );
  AOI22_X1 U17030 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13877) );
  AOI22_X1 U17031 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9666), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13876) );
  NAND4_X1 U17032 ( .A1(n13878), .A2(n13877), .A3(n13876), .A4(n13965), .ZN(
        n13885) );
  AOI22_X1 U17033 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13880) );
  AOI22_X1 U17034 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13879) );
  AND2_X1 U17035 ( .A1(n13880), .A2(n13879), .ZN(n13883) );
  AOI22_X1 U17036 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13882) );
  AOI22_X1 U17037 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9666), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13881) );
  NAND4_X1 U17038 ( .A1(n13883), .A2(n13973), .A3(n13882), .A4(n13881), .ZN(
        n13884) );
  AND2_X1 U17039 ( .A1(n13885), .A2(n13884), .ZN(n13887) );
  NAND2_X1 U17040 ( .A1(n13886), .A2(n13887), .ZN(n13909) );
  OAI211_X1 U17041 ( .C1(n13886), .C2(n13887), .A(n13909), .B(n13924), .ZN(
        n13890) );
  INV_X1 U17042 ( .A(n13887), .ZN(n13888) );
  NOR2_X1 U17043 ( .A1(n10598), .A2(n13888), .ZN(n14961) );
  AOI22_X1 U17044 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U17045 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13894) );
  AND2_X1 U17046 ( .A1(n13895), .A2(n13894), .ZN(n13898) );
  AOI22_X1 U17047 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13875), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U17048 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9667), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13896) );
  NAND4_X1 U17049 ( .A1(n13898), .A2(n13897), .A3(n13896), .A4(n13965), .ZN(
        n13905) );
  AOI22_X1 U17050 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17051 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13899) );
  AND2_X1 U17052 ( .A1(n13900), .A2(n13899), .ZN(n13903) );
  AOI22_X1 U17053 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13902) );
  AOI22_X1 U17054 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13901) );
  NAND4_X1 U17055 ( .A1(n13903), .A2(n13973), .A3(n13902), .A4(n13901), .ZN(
        n13904) );
  AND2_X1 U17056 ( .A1(n13905), .A2(n13904), .ZN(n13910) );
  XNOR2_X1 U17057 ( .A(n13909), .B(n13910), .ZN(n13906) );
  NAND2_X1 U17058 ( .A1(n10406), .A2(n13910), .ZN(n14955) );
  NOR2_X2 U17059 ( .A1(n14954), .A2(n13908), .ZN(n13927) );
  INV_X1 U17060 ( .A(n13909), .ZN(n13911) );
  AND2_X1 U17061 ( .A1(n13911), .A2(n13910), .ZN(n13925) );
  AOI22_X1 U17062 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U17063 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13912) );
  AND2_X1 U17064 ( .A1(n13913), .A2(n13912), .ZN(n13916) );
  AOI22_X1 U17065 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9655), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13915) );
  AOI22_X1 U17066 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(n9666), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13914) );
  NAND4_X1 U17067 ( .A1(n13916), .A2(n13915), .A3(n13914), .A4(n13965), .ZN(
        n13923) );
  AOI22_X1 U17068 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13918) );
  AOI22_X1 U17069 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13917) );
  AND2_X1 U17070 ( .A1(n13918), .A2(n13917), .ZN(n13921) );
  AOI22_X1 U17071 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13920) );
  AOI22_X1 U17072 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13919) );
  NAND4_X1 U17073 ( .A1(n13921), .A2(n13973), .A3(n13920), .A4(n13919), .ZN(
        n13922) );
  AND2_X1 U17074 ( .A1(n13923), .A2(n13922), .ZN(n13929) );
  NAND2_X1 U17075 ( .A1(n13925), .A2(n13929), .ZN(n14939) );
  OAI211_X1 U17076 ( .C1(n13925), .C2(n13929), .A(n14939), .B(n13924), .ZN(
        n13926) );
  NAND2_X1 U17077 ( .A1(n10406), .A2(n13929), .ZN(n14946) );
  INV_X1 U17078 ( .A(n13930), .ZN(n13943) );
  AOI22_X1 U17079 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13932) );
  AOI22_X1 U17080 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13931) );
  AND2_X1 U17081 ( .A1(n13932), .A2(n13931), .ZN(n13935) );
  AOI22_X1 U17082 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13934) );
  AOI22_X1 U17083 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n9666), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13933) );
  NAND4_X1 U17084 ( .A1(n13935), .A2(n13934), .A3(n13933), .A4(n13965), .ZN(
        n13942) );
  AOI22_X1 U17085 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13972), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13937) );
  AOI22_X1 U17086 ( .A1(n13964), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13936) );
  AND2_X1 U17087 ( .A1(n13937), .A2(n13936), .ZN(n13940) );
  AOI22_X1 U17088 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U17089 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9666), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13938) );
  NAND4_X1 U17090 ( .A1(n13940), .A2(n13973), .A3(n13939), .A4(n13938), .ZN(
        n13941) );
  AND2_X1 U17091 ( .A1(n13942), .A2(n13941), .ZN(n14940) );
  INV_X1 U17092 ( .A(n14939), .ZN(n13945) );
  AND2_X1 U17093 ( .A1(n10598), .A2(n14940), .ZN(n13944) );
  AND2_X1 U17094 ( .A1(n13945), .A2(n13944), .ZN(n13959) );
  AOI22_X1 U17095 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13947) );
  AOI22_X1 U17096 ( .A1(n13972), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13964), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13946) );
  AND2_X1 U17097 ( .A1(n13947), .A2(n13946), .ZN(n13950) );
  AOI22_X1 U17098 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13949) );
  AOI22_X1 U17099 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9667), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13948) );
  NAND4_X1 U17100 ( .A1(n13950), .A2(n13949), .A3(n13948), .A4(n13965), .ZN(
        n13957) );
  AOI22_X1 U17101 ( .A1(n13854), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13952) );
  AOI22_X1 U17102 ( .A1(n13972), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13964), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13951) );
  AND2_X1 U17103 ( .A1(n13952), .A2(n13951), .ZN(n13955) );
  AOI22_X1 U17104 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13875), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U17105 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9667), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13953) );
  NAND4_X1 U17106 ( .A1(n13955), .A2(n13973), .A3(n13954), .A4(n13953), .ZN(
        n13956) );
  AND2_X1 U17107 ( .A1(n13957), .A2(n13956), .ZN(n13958) );
  NAND2_X1 U17108 ( .A1(n13959), .A2(n13958), .ZN(n13960) );
  OAI21_X1 U17109 ( .B1(n13959), .B2(n13958), .A(n13960), .ZN(n14934) );
  NOR2_X1 U17110 ( .A1(n14935), .A2(n14934), .ZN(n14933) );
  INV_X1 U17111 ( .A(n13960), .ZN(n13961) );
  NOR2_X1 U17112 ( .A1(n14933), .A2(n13961), .ZN(n13981) );
  AOI22_X1 U17113 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9667), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13963) );
  AOI22_X1 U17114 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13875), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13962) );
  NAND2_X1 U17115 ( .A1(n13963), .A2(n13962), .ZN(n13979) );
  AOI22_X1 U17116 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13964), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13967) );
  AOI22_X1 U17117 ( .A1(n13972), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13966) );
  NAND3_X1 U17118 ( .A1(n13967), .A2(n13966), .A3(n13965), .ZN(n13978) );
  AOI22_X1 U17119 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9666), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13970) );
  AOI22_X1 U17120 ( .A1(n13968), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9655), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13969) );
  NAND2_X1 U17121 ( .A1(n13970), .A2(n13969), .ZN(n13977) );
  AOI22_X1 U17122 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13971), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13975) );
  AOI22_X1 U17123 ( .A1(n13972), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13964), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13974) );
  NAND3_X1 U17124 ( .A1(n13975), .A2(n13974), .A3(n13973), .ZN(n13976) );
  OAI22_X1 U17125 ( .A1(n13979), .A2(n13978), .B1(n13977), .B2(n13976), .ZN(
        n13980) );
  XNOR2_X1 U17126 ( .A(n13981), .B(n13980), .ZN(n13990) );
  INV_X1 U17127 ( .A(n19209), .ZN(n15042) );
  INV_X1 U17128 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n13984) );
  AOI22_X1 U17129 ( .A1(n19207), .A2(n19219), .B1(n19264), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n13983) );
  OAI21_X1 U17130 ( .B1(n15042), .B2(n13984), .A(n13983), .ZN(n13986) );
  NOR2_X1 U17131 ( .A1(n15308), .A2(n19215), .ZN(n13985) );
  AOI211_X1 U17132 ( .C1(BUF1_REG_30__SCAN_IN), .C2(n19208), .A(n13986), .B(
        n13985), .ZN(n13987) );
  OAI21_X1 U17133 ( .B1(n13990), .B2(n19216), .A(n13987), .ZN(P2_U2889) );
  NOR2_X1 U17134 ( .A1(n15315), .A2(n15004), .ZN(n13988) );
  AOI21_X1 U17135 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15004), .A(n13988), .ZN(
        n13989) );
  OAI21_X1 U17136 ( .B1(n13990), .B2(n15025), .A(n13989), .ZN(P2_U2857) );
  INV_X1 U17137 ( .A(n14461), .ZN(n14071) );
  NAND2_X1 U17138 ( .A1(n14055), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n13992) );
  NAND2_X1 U17139 ( .A1(n13022), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13991) );
  NAND2_X1 U17140 ( .A1(n13992), .A2(n13991), .ZN(n14074) );
  MUX2_X1 U17141 ( .A(n14047), .B(n14008), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13995) );
  NAND2_X1 U17142 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n13022), .ZN(
        n13993) );
  AND2_X1 U17143 ( .A1(n14031), .A2(n13993), .ZN(n13994) );
  NAND2_X1 U17144 ( .A1(n13995), .A2(n13994), .ZN(n14223) );
  MUX2_X1 U17145 ( .A(n14048), .B(n14053), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13997) );
  INV_X1 U17146 ( .A(n14055), .ZN(n14052) );
  INV_X1 U17147 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16178) );
  NAND2_X1 U17148 ( .A1(n14052), .A2(n16178), .ZN(n13996) );
  MUX2_X1 U17149 ( .A(n14047), .B(n14008), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13998) );
  INV_X1 U17150 ( .A(n13998), .ZN(n14001) );
  NAND2_X1 U17151 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n13022), .ZN(
        n13999) );
  NAND2_X1 U17152 ( .A1(n14031), .A2(n13999), .ZN(n14000) );
  NOR2_X1 U17153 ( .A1(n14001), .A2(n14000), .ZN(n14294) );
  INV_X1 U17154 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16164) );
  INV_X1 U17155 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14286) );
  NAND2_X1 U17156 ( .A1(n14043), .A2(n14286), .ZN(n14002) );
  OAI211_X1 U17157 ( .C1(n14073), .C2(n16164), .A(n14002), .B(n14008), .ZN(
        n14003) );
  OAI21_X1 U17158 ( .B1(n14048), .B2(P1_EBX_REG_13__SCAN_IN), .A(n14003), .ZN(
        n14212) );
  INV_X1 U17159 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14283) );
  NAND2_X1 U17160 ( .A1(n14050), .A2(n14283), .ZN(n14007) );
  INV_X1 U17161 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14440) );
  NAND2_X1 U17162 ( .A1(n14008), .A2(n14440), .ZN(n14005) );
  NAND2_X1 U17163 ( .A1(n14043), .A2(n14283), .ZN(n14004) );
  NAND3_X1 U17164 ( .A1(n14005), .A2(n14053), .A3(n14004), .ZN(n14006) );
  NOR2_X2 U17165 ( .A1(n14213), .A2(n14198), .ZN(n16053) );
  INV_X1 U17166 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n16085) );
  NAND2_X1 U17167 ( .A1(n14034), .A2(n16085), .ZN(n14011) );
  INV_X1 U17168 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16155) );
  NAND2_X1 U17169 ( .A1(n14043), .A2(n16085), .ZN(n14009) );
  OAI211_X1 U17170 ( .C1(n14073), .C2(n16155), .A(n14009), .B(n14008), .ZN(
        n14010) );
  NAND2_X1 U17171 ( .A1(n16053), .A2(n16052), .ZN(n16054) );
  MUX2_X1 U17172 ( .A(n14047), .B(n14012), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n14013) );
  INV_X1 U17173 ( .A(n14013), .ZN(n14016) );
  NAND2_X1 U17174 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n13022), .ZN(
        n14014) );
  NAND2_X1 U17175 ( .A1(n14031), .A2(n14014), .ZN(n14015) );
  NOR2_X1 U17176 ( .A1(n14016), .A2(n14015), .ZN(n14187) );
  MUX2_X1 U17177 ( .A(n14048), .B(n14053), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14018) );
  NAND2_X1 U17178 ( .A1(n14052), .A2(n14446), .ZN(n14017) );
  NAND2_X1 U17179 ( .A1(n14018), .A2(n14017), .ZN(n16046) );
  NOR2_X4 U17180 ( .A1(n16045), .A2(n16046), .ZN(n16044) );
  MUX2_X1 U17181 ( .A(n14047), .B(n14008), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n14021) );
  NAND2_X1 U17182 ( .A1(n13022), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14019) );
  AND2_X1 U17183 ( .A1(n14031), .A2(n14019), .ZN(n14020) );
  NAND2_X1 U17184 ( .A1(n14021), .A2(n14020), .ZN(n14279) );
  INV_X1 U17185 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n16017) );
  NAND2_X1 U17186 ( .A1(n14034), .A2(n16017), .ZN(n14024) );
  INV_X1 U17187 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14538) );
  NAND2_X1 U17188 ( .A1(n14043), .A2(n16017), .ZN(n14022) );
  OAI211_X1 U17189 ( .C1(n14073), .C2(n14538), .A(n14022), .B(n14008), .ZN(
        n14023) );
  INV_X1 U17190 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14172) );
  NAND2_X1 U17191 ( .A1(n14050), .A2(n14172), .ZN(n14028) );
  INV_X1 U17192 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14548) );
  NAND2_X1 U17193 ( .A1(n14008), .A2(n14548), .ZN(n14026) );
  NAND2_X1 U17194 ( .A1(n14043), .A2(n14172), .ZN(n14025) );
  NAND3_X1 U17195 ( .A1(n14026), .A2(n14053), .A3(n14025), .ZN(n14027) );
  AND2_X1 U17196 ( .A1(n14028), .A2(n14027), .ZN(n14171) );
  MUX2_X1 U17197 ( .A(n14048), .B(n14053), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n14029) );
  OAI21_X1 U17198 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14055), .A(
        n14029), .ZN(n14265) );
  MUX2_X1 U17199 ( .A(n14047), .B(n14008), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14033) );
  NAND2_X1 U17200 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n13022), .ZN(
        n14030) );
  AND2_X1 U17201 ( .A1(n14031), .A2(n14030), .ZN(n14032) );
  NAND2_X1 U17202 ( .A1(n14033), .A2(n14032), .ZN(n14260) );
  AND2_X2 U17203 ( .A1(n14268), .A2(n14260), .ZN(n14724) );
  INV_X1 U17204 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n16081) );
  NAND2_X1 U17205 ( .A1(n14034), .A2(n16081), .ZN(n14037) );
  INV_X1 U17206 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14730) );
  NAND2_X1 U17207 ( .A1(n14043), .A2(n16081), .ZN(n14035) );
  OAI211_X1 U17208 ( .C1(n14073), .C2(n14730), .A(n14035), .B(n14008), .ZN(
        n14036) );
  AND2_X1 U17209 ( .A1(n14037), .A2(n14036), .ZN(n14723) );
  MUX2_X1 U17210 ( .A(n14047), .B(n14008), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n14039) );
  NAND2_X1 U17211 ( .A1(n13022), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14038) );
  AND2_X1 U17212 ( .A1(n14039), .A2(n14038), .ZN(n14151) );
  INV_X1 U17213 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14452) );
  INV_X1 U17214 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14040) );
  NAND2_X1 U17215 ( .A1(n14043), .A2(n14040), .ZN(n14041) );
  OAI211_X1 U17216 ( .C1(n14073), .C2(n14452), .A(n14041), .B(n14008), .ZN(
        n14042) );
  OAI21_X1 U17217 ( .B1(n14048), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14042), .ZN(
        n14142) );
  INV_X1 U17218 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14699) );
  NAND2_X1 U17219 ( .A1(n14008), .A2(n14699), .ZN(n14045) );
  INV_X1 U17220 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14253) );
  NAND2_X1 U17221 ( .A1(n14043), .A2(n14253), .ZN(n14044) );
  NAND3_X1 U17222 ( .A1(n14045), .A2(n14053), .A3(n14044), .ZN(n14046) );
  OAI21_X1 U17223 ( .B1(n14047), .B2(P1_EBX_REG_26__SCAN_IN), .A(n14046), .ZN(
        n14131) );
  NAND2_X1 U17224 ( .A1(n14141), .A2(n14131), .ZN(n14133) );
  MUX2_X1 U17225 ( .A(n14048), .B(n14053), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14049) );
  OAI21_X1 U17226 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14055), .A(
        n14049), .ZN(n14120) );
  MUX2_X1 U17227 ( .A(n14050), .B(n13435), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14051) );
  AOI21_X1 U17228 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n13022), .A(
        n14051), .ZN(n14102) );
  NOR2_X1 U17229 ( .A1(n13022), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14054) );
  INV_X1 U17230 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14472) );
  AOI21_X1 U17231 ( .B1(n14052), .B2(n14472), .A(n14054), .ZN(n14072) );
  MUX2_X1 U17232 ( .A(n14054), .B(n14072), .S(n14053), .Z(n14086) );
  AOI22_X1 U17233 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(n14055), .B1(n13022), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14056) );
  XNOR2_X1 U17234 ( .A(n14057), .B(n14056), .ZN(n14655) );
  INV_X1 U17235 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20914) );
  NAND3_X1 U17236 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n14197) );
  NOR2_X1 U17237 ( .A1(n14589), .A2(n14197), .ZN(n14183) );
  NAND4_X1 U17238 ( .A1(n14183), .A2(P1_REIP_REG_15__SCAN_IN), .A3(
        P1_REIP_REG_17__SCAN_IN), .A4(P1_REIP_REG_16__SCAN_IN), .ZN(n16020) );
  NAND2_X1 U17239 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14168) );
  NOR3_X1 U17240 ( .A1(n20083), .A2(n16020), .A3(n14168), .ZN(n14058) );
  NAND4_X1 U17241 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .A4(n14058), .ZN(n14169) );
  NOR2_X1 U17242 ( .A1(n20914), .A2(n14169), .ZN(n15995) );
  NAND2_X1 U17243 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15995), .ZN(n15988) );
  INV_X1 U17244 ( .A(n15988), .ZN(n14059) );
  AND2_X1 U17245 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14059), .ZN(n14156) );
  AND2_X1 U17246 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14060) );
  NAND2_X1 U17247 ( .A1(n14156), .A2(n14060), .ZN(n14112) );
  AND2_X1 U17248 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14103) );
  NAND2_X1 U17249 ( .A1(n14103), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14065) );
  NOR2_X1 U17250 ( .A1(n14112), .A2(n14065), .ZN(n14061) );
  NAND2_X1 U17251 ( .A1(n14232), .A2(n14061), .ZN(n14062) );
  NAND2_X1 U17252 ( .A1(n16021), .A2(n14062), .ZN(n14106) );
  NAND2_X1 U17253 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14063) );
  NAND2_X1 U17254 ( .A1(n16021), .A2(n14063), .ZN(n14064) );
  AND2_X1 U17255 ( .A1(n14106), .A2(n14064), .ZN(n14080) );
  INV_X1 U17256 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14068) );
  AOI22_X1 U17257 ( .A1(n20143), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20139), .ZN(n14067) );
  OR2_X1 U17258 ( .A1(n20102), .A2(n14112), .ZN(n14127) );
  NOR2_X1 U17259 ( .A1(n14127), .A2(n14065), .ZN(n14091) );
  NAND4_X1 U17260 ( .A1(n14091), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_30__SCAN_IN), .A4(n14068), .ZN(n14066) );
  OAI211_X1 U17261 ( .C1(n14080), .C2(n14068), .A(n14067), .B(n14066), .ZN(
        n14069) );
  AOI21_X1 U17262 ( .B1(n14655), .B2(n20145), .A(n14069), .ZN(n14070) );
  OAI21_X1 U17263 ( .B1(n14071), .B2(n20104), .A(n14070), .ZN(P1_U2809) );
  INV_X1 U17264 ( .A(n14078), .ZN(n14468) );
  NAND2_X1 U17265 ( .A1(n14468), .A2(n20119), .ZN(n14084) );
  AOI21_X1 U17266 ( .B1(n14091), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U17267 ( .A1(n20143), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20139), .ZN(n14079) );
  OAI21_X1 U17268 ( .B1(n14081), .B2(n14080), .A(n14079), .ZN(n14082) );
  AOI21_X1 U17269 ( .B1(n20140), .B2(n14464), .A(n14082), .ZN(n14083) );
  OAI211_X1 U17270 ( .C1(n20128), .C2(n14663), .A(n14084), .B(n14083), .ZN(
        P1_U2810) );
  OAI21_X1 U17271 ( .B1(n14101), .B2(n14086), .A(n14085), .ZN(n14667) );
  INV_X1 U17272 ( .A(n14087), .ZN(n14088) );
  NAND2_X1 U17273 ( .A1(n14477), .A2(n20119), .ZN(n14098) );
  INV_X1 U17274 ( .A(n14475), .ZN(n14096) );
  INV_X1 U17275 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14094) );
  NAND2_X1 U17276 ( .A1(n14091), .A2(n14094), .ZN(n14093) );
  AOI22_X1 U17277 ( .A1(n20143), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20139), .ZN(n14092) );
  OAI211_X1 U17278 ( .C1(n14106), .C2(n14094), .A(n14093), .B(n14092), .ZN(
        n14095) );
  AOI21_X1 U17279 ( .B1(n20140), .B2(n14096), .A(n14095), .ZN(n14097) );
  OAI211_X1 U17280 ( .C1(n20128), .C2(n14667), .A(n14098), .B(n14097), .ZN(
        P1_U2811) );
  AOI21_X1 U17281 ( .B1(n14100), .B2(n14099), .A(n14087), .ZN(n14491) );
  INV_X1 U17282 ( .A(n14491), .ZN(n14323) );
  AOI21_X1 U17283 ( .B1(n14102), .B2(n14119), .A(n14101), .ZN(n14684) );
  INV_X1 U17284 ( .A(n14127), .ZN(n14115) );
  AOI21_X1 U17285 ( .B1(n14115), .B2(n14103), .A(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14107) );
  NAND2_X1 U17286 ( .A1(n20140), .A2(n14487), .ZN(n14105) );
  AOI22_X1 U17287 ( .A1(n20143), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20139), .ZN(n14104) );
  OAI211_X1 U17288 ( .C1(n14107), .C2(n14106), .A(n14105), .B(n14104), .ZN(
        n14108) );
  AOI21_X1 U17289 ( .B1(n14684), .B2(n20145), .A(n14108), .ZN(n14109) );
  OAI21_X1 U17290 ( .B1(n14323), .B2(n20104), .A(n14109), .ZN(P1_U2812) );
  INV_X1 U17291 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14128) );
  NOR2_X1 U17292 ( .A1(n14112), .A2(n14128), .ZN(n14113) );
  NAND2_X1 U17293 ( .A1(n14232), .A2(n14113), .ZN(n14114) );
  NAND2_X1 U17294 ( .A1(n16021), .A2(n14114), .ZN(n14126) );
  INV_X1 U17295 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20924) );
  NAND3_X1 U17296 ( .A1(n14115), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n20924), 
        .ZN(n14117) );
  AOI22_X1 U17297 ( .A1(n20143), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20139), .ZN(n14116) );
  OAI211_X1 U17298 ( .C1(n14126), .C2(n20924), .A(n14117), .B(n14116), .ZN(
        n14118) );
  AOI21_X1 U17299 ( .B1(n20140), .B2(n14502), .A(n14118), .ZN(n14122) );
  AOI21_X1 U17300 ( .B1(n14120), .B2(n14133), .A(n10050), .ZN(n14692) );
  NAND2_X1 U17301 ( .A1(n14692), .A2(n20145), .ZN(n14121) );
  OAI211_X1 U17302 ( .C1(n14499), .C2(n20104), .A(n14122), .B(n14121), .ZN(
        P1_U2813) );
  INV_X1 U17303 ( .A(n14110), .ZN(n14124) );
  AOI21_X1 U17304 ( .B1(n14128), .B2(n14127), .A(n14126), .ZN(n14130) );
  OAI22_X1 U17305 ( .A1(n20117), .A2(n14253), .B1(n14506), .B2(n20111), .ZN(
        n14129) );
  AOI211_X1 U17306 ( .C1(n20140), .C2(n14510), .A(n14130), .B(n14129), .ZN(
        n14135) );
  OR2_X1 U17307 ( .A1(n14141), .A2(n14131), .ZN(n14132) );
  AND2_X1 U17308 ( .A1(n14133), .A2(n14132), .ZN(n14701) );
  NAND2_X1 U17309 ( .A1(n14701), .A2(n20145), .ZN(n14134) );
  OAI211_X1 U17310 ( .C1(n14507), .C2(n20104), .A(n14135), .B(n14134), .ZN(
        P1_U2814) );
  INV_X1 U17311 ( .A(n14136), .ZN(n14140) );
  INV_X1 U17313 ( .A(n14138), .ZN(n14139) );
  AOI21_X1 U17314 ( .B1(n14140), .B2(n14139), .A(n14123), .ZN(n14516) );
  INV_X1 U17315 ( .A(n14516), .ZN(n14337) );
  AOI21_X1 U17316 ( .B1(n14142), .B2(n14153), .A(n14141), .ZN(n14709) );
  NOR2_X1 U17317 ( .A1(n20098), .A2(n14514), .ZN(n14149) );
  NAND2_X1 U17318 ( .A1(n14232), .A2(n14156), .ZN(n14143) );
  NAND2_X1 U17319 ( .A1(n16021), .A2(n14143), .ZN(n15987) );
  INV_X1 U17320 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20921) );
  AOI22_X1 U17321 ( .A1(n20143), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20139), .ZN(n14147) );
  INV_X1 U17322 ( .A(n14156), .ZN(n14144) );
  OAI21_X1 U17323 ( .B1(n14144), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14145) );
  OAI211_X1 U17324 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(P1_REIP_REG_24__SCAN_IN), .A(n20094), .B(n14145), .ZN(n14146) );
  OAI211_X1 U17325 ( .C1(n15987), .C2(n20921), .A(n14147), .B(n14146), .ZN(
        n14148) );
  AOI211_X1 U17326 ( .C1(n14709), .C2(n20145), .A(n14149), .B(n14148), .ZN(
        n14150) );
  OAI21_X1 U17327 ( .B1(n14337), .B2(n20104), .A(n14150), .ZN(P1_U2815) );
  NAND2_X1 U17328 ( .A1(n14726), .A2(n14151), .ZN(n14152) );
  NAND2_X1 U17329 ( .A1(n14153), .A2(n14152), .ZN(n14712) );
  INV_X1 U17330 ( .A(n14154), .ZN(n14344) );
  AOI21_X1 U17331 ( .B1(n14155), .B2(n14344), .A(n14138), .ZN(n14525) );
  NAND2_X1 U17332 ( .A1(n14525), .A2(n20119), .ZN(n14163) );
  INV_X1 U17333 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14160) );
  AOI22_X1 U17334 ( .A1(n20143), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20139), .ZN(n14159) );
  NAND2_X1 U17335 ( .A1(n14156), .A2(n14160), .ZN(n14157) );
  OR2_X1 U17336 ( .A1(n20102), .A2(n14157), .ZN(n14158) );
  OAI211_X1 U17337 ( .C1(n15987), .C2(n14160), .A(n14159), .B(n14158), .ZN(
        n14161) );
  AOI21_X1 U17338 ( .B1(n20140), .B2(n14521), .A(n14161), .ZN(n14162) );
  OAI211_X1 U17339 ( .C1(n20128), .C2(n14712), .A(n14163), .B(n14162), .ZN(
        P1_U2816) );
  OAI21_X1 U17340 ( .B1(n14164), .B2(n14166), .A(n14165), .ZN(n14551) );
  INV_X1 U17341 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20084) );
  NOR3_X1 U17342 ( .A1(n20102), .A2(n20083), .A3(n20084), .ZN(n14230) );
  NAND2_X1 U17343 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n14230), .ZN(n16074) );
  NOR3_X1 U17344 ( .A1(n14589), .A2(n14197), .A3(n16074), .ZN(n14179) );
  NAND4_X1 U17345 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_17__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .A4(n14179), .ZN(n16040) );
  INV_X1 U17346 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14167) );
  OAI21_X1 U17347 ( .B1(n14168), .B2(n16040), .A(n14167), .ZN(n14177) );
  INV_X1 U17348 ( .A(n14169), .ZN(n16008) );
  OAI21_X1 U17349 ( .B1(n16008), .B2(n20102), .A(n14232), .ZN(n16012) );
  INV_X1 U17350 ( .A(n14554), .ZN(n14175) );
  INV_X1 U17351 ( .A(n14266), .ZN(n14170) );
  AOI21_X1 U17352 ( .B1(n14171), .B2(n14274), .A(n14170), .ZN(n14768) );
  OAI22_X1 U17353 ( .A1(n20117), .A2(n14172), .B1(n20111), .B2(n14550), .ZN(
        n14173) );
  AOI21_X1 U17354 ( .B1(n14768), .B2(n20145), .A(n14173), .ZN(n14174) );
  OAI21_X1 U17355 ( .B1(n14175), .B2(n20098), .A(n14174), .ZN(n14176) );
  AOI21_X1 U17356 ( .B1(n14177), .B2(n16012), .A(n14176), .ZN(n14178) );
  OAI21_X1 U17357 ( .B1(n14551), .B2(n20104), .A(n14178), .ZN(P1_U2820) );
  INV_X1 U17358 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21094) );
  INV_X1 U17359 ( .A(n14179), .ZN(n14180) );
  NOR2_X1 U17360 ( .A1(n21094), .A2(n14180), .ZN(n16041) );
  INV_X1 U17361 ( .A(n16041), .ZN(n14186) );
  NOR2_X1 U17362 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14180), .ZN(n16059) );
  INV_X1 U17363 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n16199) );
  NOR2_X1 U17364 ( .A1(n16199), .A2(n20084), .ZN(n14182) );
  AOI21_X1 U17365 ( .B1(n14182), .B2(n14181), .A(n14184), .ZN(n16023) );
  INV_X1 U17366 ( .A(n16023), .ZN(n16072) );
  OAI21_X1 U17367 ( .B1(n14184), .B2(n14183), .A(n16072), .ZN(n16051) );
  NOR2_X1 U17368 ( .A1(n16059), .A2(n16051), .ZN(n14185) );
  MUX2_X1 U17369 ( .A(n14186), .B(n14185), .S(P1_REIP_REG_16__SCAN_IN), .Z(
        n14192) );
  NAND2_X1 U17370 ( .A1(n16054), .A2(n14187), .ZN(n14188) );
  NAND2_X1 U17371 ( .A1(n16045), .A2(n14188), .ZN(n14796) );
  AOI22_X1 U17372 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n20143), .B1(n14582), 
        .B2(n20140), .ZN(n14189) );
  OAI21_X1 U17373 ( .B1(n20128), .B2(n14796), .A(n14189), .ZN(n14190) );
  AOI211_X1 U17374 ( .C1(n20139), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n14190), .B(n16236), .ZN(n14191) );
  OAI211_X1 U17375 ( .C1(n14579), .C2(n20104), .A(n14192), .B(n14191), .ZN(
        P1_U2824) );
  OAI21_X1 U17376 ( .B1(n14193), .B2(n14196), .A(n14195), .ZN(n14595) );
  OAI21_X1 U17377 ( .B1(n14197), .B2(n16074), .A(n14589), .ZN(n14202) );
  INV_X1 U17378 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14200) );
  AND2_X1 U17379 ( .A1(n14213), .A2(n14198), .ZN(n14199) );
  OR2_X1 U17380 ( .A1(n14199), .A2(n16053), .ZN(n14816) );
  OAI22_X1 U17381 ( .A1(n14200), .A2(n20111), .B1(n20128), .B2(n14816), .ZN(
        n14201) );
  AOI211_X1 U17382 ( .C1(n16051), .C2(n14202), .A(n16236), .B(n14201), .ZN(
        n14205) );
  INV_X1 U17383 ( .A(n14590), .ZN(n14203) );
  AOI22_X1 U17384 ( .A1(n20140), .A2(n14203), .B1(n20143), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14204) );
  OAI211_X1 U17385 ( .C1(n14595), .C2(n20104), .A(n14205), .B(n14204), .ZN(
        P1_U2826) );
  OAI21_X1 U17386 ( .B1(n21148), .B2(n11411), .A(n14208), .ZN(n14300) );
  OAI21_X1 U17387 ( .B1(n14300), .B2(n14301), .A(n14208), .ZN(n14289) );
  INV_X1 U17388 ( .A(n14193), .ZN(n14210) );
  OAI21_X1 U17389 ( .B1(n14298), .B2(n14294), .A(n14212), .ZN(n14214) );
  AND2_X1 U17390 ( .A1(n14214), .A2(n14213), .ZN(n16165) );
  AOI22_X1 U17391 ( .A1(n16165), .A2(n20145), .B1(n20143), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14215) );
  OAI211_X1 U17392 ( .C1(n20111), .C2(n14606), .A(n14215), .B(n20227), .ZN(
        n14220) );
  NAND2_X1 U17393 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14216) );
  NOR2_X1 U17394 ( .A1(n14216), .A2(n16074), .ZN(n14218) );
  AOI21_X1 U17395 ( .B1(n14216), .B2(n16021), .A(n16023), .ZN(n16062) );
  INV_X1 U17396 ( .A(n16062), .ZN(n14217) );
  MUX2_X1 U17397 ( .A(n14218), .B(n14217), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14219) );
  AOI211_X1 U17398 ( .C1(n14608), .C2(n20140), .A(n14220), .B(n14219), .ZN(
        n14221) );
  OAI21_X1 U17399 ( .B1(n14611), .B2(n20104), .A(n14221), .ZN(P1_U2827) );
  AOI21_X1 U17400 ( .B1(n14222), .B2(n13599), .A(n21148), .ZN(n14619) );
  INV_X1 U17401 ( .A(n14619), .ZN(n14395) );
  NOR2_X1 U17402 ( .A1(n14224), .A2(n14223), .ZN(n14225) );
  OR2_X1 U17403 ( .A1(n9702), .A2(n14225), .ZN(n16201) );
  AOI21_X1 U17404 ( .B1(n20139), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16236), .ZN(n14228) );
  INV_X1 U17405 ( .A(n14617), .ZN(n14226) );
  AOI22_X1 U17406 ( .A1(n20140), .A2(n14226), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n20143), .ZN(n14227) );
  OAI211_X1 U17407 ( .C1(n20128), .C2(n16201), .A(n14228), .B(n14227), .ZN(
        n14229) );
  AOI221_X1 U17408 ( .B1(n16023), .B2(P1_REIP_REG_10__SCAN_IN), .C1(n14230), 
        .C2(n16199), .A(n14229), .ZN(n14231) );
  OAI21_X1 U17409 ( .B1(n14395), .B2(n20104), .A(n14231), .ZN(P1_U2830) );
  OAI21_X1 U17410 ( .B1(n20093), .B2(n20102), .A(n14232), .ZN(n20113) );
  NOR2_X1 U17411 ( .A1(n20117), .A2(n14233), .ZN(n14234) );
  AOI211_X1 U17412 ( .C1(n20139), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16236), .B(n14234), .ZN(n14235) );
  OAI21_X1 U17413 ( .B1(n20128), .B2(n14236), .A(n14235), .ZN(n14237) );
  AOI21_X1 U17414 ( .B1(n20142), .B2(n14238), .A(n14237), .ZN(n14239) );
  OAI21_X1 U17415 ( .B1(n20098), .B2(n14240), .A(n14239), .ZN(n14243) );
  NOR3_X1 U17416 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20102), .A3(n14241), .ZN(
        n14242) );
  AOI211_X1 U17417 ( .C1(P1_REIP_REG_4__SCAN_IN), .C2(n20113), .A(n14243), .B(
        n14242), .ZN(n14244) );
  OAI21_X1 U17418 ( .B1(n20132), .B2(n14245), .A(n14244), .ZN(P1_U2836) );
  INV_X1 U17419 ( .A(n14655), .ZN(n14247) );
  INV_X1 U17420 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14246) );
  OAI22_X1 U17421 ( .A1(n14247), .A2(n16076), .B1(n20161), .B2(n14246), .ZN(
        P1_U2841) );
  INV_X1 U17422 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14248) );
  OAI222_X1 U17423 ( .A1(n16075), .A2(n14078), .B1(n14248), .B2(n20161), .C1(
        n14663), .C2(n16076), .ZN(P1_U2842) );
  INV_X1 U17424 ( .A(n14477), .ZN(n14318) );
  INV_X1 U17425 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14249) );
  OAI222_X1 U17426 ( .A1(n16075), .A2(n14318), .B1(n14249), .B2(n20161), .C1(
        n14667), .C2(n16076), .ZN(P1_U2843) );
  AOI22_X1 U17427 ( .A1(n14684), .A2(n20156), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14296), .ZN(n14250) );
  OAI21_X1 U17428 ( .B1(n14323), .B2(n16075), .A(n14250), .ZN(P1_U2844) );
  AOI22_X1 U17429 ( .A1(n14692), .A2(n20156), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14296), .ZN(n14251) );
  OAI21_X1 U17430 ( .B1(n14499), .B2(n16075), .A(n14251), .ZN(P1_U2845) );
  INV_X1 U17431 ( .A(n14701), .ZN(n14252) );
  AOI22_X1 U17432 ( .A1(n14709), .A2(n20156), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n14296), .ZN(n14254) );
  OAI21_X1 U17433 ( .B1(n14337), .B2(n16075), .A(n14254), .ZN(P1_U2847) );
  INV_X1 U17434 ( .A(n14525), .ZN(n14341) );
  INV_X1 U17435 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14255) );
  OAI222_X1 U17436 ( .A1(n16075), .A2(n14341), .B1(n20161), .B2(n14255), .C1(
        n14712), .C2(n16076), .ZN(P1_U2848) );
  OAI21_X1 U17437 ( .B1(n14256), .B2(n10234), .A(n14258), .ZN(n16002) );
  INV_X1 U17438 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14261) );
  INV_X1 U17439 ( .A(n14724), .ZN(n14259) );
  OAI21_X1 U17440 ( .B1(n14268), .B2(n14260), .A(n14259), .ZN(n16005) );
  OAI222_X1 U17441 ( .A1(n16002), .A2(n16075), .B1(n20161), .B2(n14261), .C1(
        n16005), .C2(n16076), .ZN(P1_U2850) );
  NAND2_X1 U17442 ( .A1(n14165), .A2(n14262), .ZN(n14263) );
  AND2_X1 U17443 ( .A1(n14264), .A2(n14263), .ZN(n16011) );
  INV_X1 U17444 ( .A(n16011), .ZN(n14356) );
  AND2_X1 U17445 ( .A1(n14266), .A2(n14265), .ZN(n14267) );
  NOR2_X1 U17446 ( .A1(n14268), .A2(n14267), .ZN(n16010) );
  AOI22_X1 U17447 ( .A1(n16010), .A2(n20156), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14296), .ZN(n14269) );
  OAI21_X1 U17448 ( .B1(n14356), .B2(n16075), .A(n14269), .ZN(P1_U2851) );
  AOI22_X1 U17449 ( .A1(n14768), .A2(n20156), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n14296), .ZN(n14270) );
  OAI21_X1 U17450 ( .B1(n14551), .B2(n16075), .A(n14270), .ZN(P1_U2852) );
  AND2_X1 U17451 ( .A1(n14271), .A2(n14272), .ZN(n14273) );
  OR2_X1 U17452 ( .A1(n14164), .A2(n14273), .ZN(n14558) );
  OAI21_X1 U17453 ( .B1(n14281), .B2(n14275), .A(n14274), .ZN(n16018) );
  INV_X1 U17454 ( .A(n16018), .ZN(n14776) );
  AOI22_X1 U17455 ( .A1(n14776), .A2(n20156), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14296), .ZN(n14276) );
  OAI21_X1 U17456 ( .B1(n14558), .B2(n16075), .A(n14276), .ZN(P1_U2853) );
  OAI21_X1 U17457 ( .B1(n14277), .B2(n14278), .A(n14271), .ZN(n16035) );
  INV_X1 U17458 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16031) );
  NOR2_X1 U17459 ( .A1(n16044), .A2(n14279), .ZN(n14280) );
  OR2_X1 U17460 ( .A1(n14281), .A2(n14280), .ZN(n16034) );
  OAI222_X1 U17461 ( .A1(n16035), .A2(n16075), .B1(n20161), .B2(n16031), .C1(
        n16034), .C2(n16076), .ZN(P1_U2854) );
  INV_X1 U17462 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14282) );
  OAI222_X1 U17463 ( .A1(n14579), .A2(n16075), .B1(n20161), .B2(n14282), .C1(
        n14796), .C2(n16076), .ZN(P1_U2856) );
  OAI22_X1 U17464 ( .A1(n14816), .A2(n16076), .B1(n14283), .B2(n20161), .ZN(
        n14284) );
  INV_X1 U17465 ( .A(n14284), .ZN(n14285) );
  OAI21_X1 U17466 ( .B1(n14595), .B2(n16075), .A(n14285), .ZN(P1_U2858) );
  NOR2_X1 U17467 ( .A1(n20161), .A2(n14286), .ZN(n14287) );
  AOI21_X1 U17468 ( .B1(n16165), .B2(n20156), .A(n14287), .ZN(n14288) );
  OAI21_X1 U17469 ( .B1(n14611), .B2(n16075), .A(n14288), .ZN(P1_U2859) );
  INV_X1 U17470 ( .A(n14289), .ZN(n14293) );
  INV_X1 U17471 ( .A(n14290), .ZN(n14292) );
  INV_X1 U17472 ( .A(n16108), .ZN(n14388) );
  INV_X1 U17473 ( .A(n14294), .ZN(n14295) );
  XNOR2_X1 U17474 ( .A(n14298), .B(n14295), .ZN(n16182) );
  AOI22_X1 U17475 ( .A1(n16182), .A2(n20156), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14296), .ZN(n14297) );
  OAI21_X1 U17476 ( .B1(n14388), .B2(n16075), .A(n14297), .ZN(P1_U2860) );
  OAI21_X1 U17477 ( .B1(n9702), .B2(n14299), .A(n14298), .ZN(n16067) );
  INV_X1 U17478 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14302) );
  XOR2_X1 U17479 ( .A(n14301), .B(n14300), .Z(n16117) );
  INV_X1 U17480 ( .A(n16117), .ZN(n14391) );
  OAI222_X1 U17481 ( .A1(n16067), .A2(n16076), .B1(n14302), .B2(n20161), .C1(
        n14391), .C2(n16075), .ZN(P1_U2861) );
  INV_X1 U17482 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14303) );
  OAI222_X1 U17483 ( .A1(n16201), .A2(n16076), .B1(n20161), .B2(n14303), .C1(
        n14395), .C2(n16075), .ZN(P1_U2862) );
  AND2_X1 U17484 ( .A1(n14305), .A2(n20292), .ZN(n14306) );
  NAND2_X1 U17485 ( .A1(n14389), .A2(n14306), .ZN(n14375) );
  INV_X1 U17486 ( .A(DATAI_14_), .ZN(n14308) );
  INV_X1 U17487 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14307) );
  MUX2_X1 U17488 ( .A(n14308), .B(n14307), .S(n20241), .Z(n20203) );
  OAI22_X1 U17489 ( .A1(n14375), .A2(n20203), .B1(n14389), .B2(n14309), .ZN(
        n14310) );
  AOI21_X1 U17490 ( .B1(n14377), .B2(BUF1_REG_30__SCAN_IN), .A(n14310), .ZN(
        n14312) );
  NAND2_X1 U17491 ( .A1(n14378), .A2(DATAI_30_), .ZN(n14311) );
  OAI211_X1 U17492 ( .C1(n14078), .C2(n14396), .A(n14312), .B(n14311), .ZN(
        P1_U2874) );
  INV_X1 U17493 ( .A(DATAI_13_), .ZN(n14314) );
  MUX2_X1 U17494 ( .A(n14314), .B(n14313), .S(n20241), .Z(n20200) );
  OAI22_X1 U17495 ( .A1(n14375), .A2(n20200), .B1(n14389), .B2(n12903), .ZN(
        n14315) );
  AOI21_X1 U17496 ( .B1(n14377), .B2(BUF1_REG_29__SCAN_IN), .A(n14315), .ZN(
        n14317) );
  NAND2_X1 U17497 ( .A1(n14378), .A2(DATAI_29_), .ZN(n14316) );
  OAI211_X1 U17498 ( .C1(n14318), .C2(n14396), .A(n14317), .B(n14316), .ZN(
        P1_U2875) );
  INV_X1 U17499 ( .A(DATAI_12_), .ZN(n14319) );
  INV_X1 U17500 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16545) );
  MUX2_X1 U17501 ( .A(n14319), .B(n16545), .S(n20241), .Z(n20197) );
  OAI22_X1 U17502 ( .A1(n14375), .A2(n20197), .B1(n14389), .B2(n12908), .ZN(
        n14320) );
  AOI21_X1 U17503 ( .B1(n14377), .B2(BUF1_REG_28__SCAN_IN), .A(n14320), .ZN(
        n14322) );
  NAND2_X1 U17504 ( .A1(n14378), .A2(DATAI_28_), .ZN(n14321) );
  OAI211_X1 U17505 ( .C1(n14323), .C2(n14396), .A(n14322), .B(n14321), .ZN(
        P1_U2876) );
  INV_X1 U17506 ( .A(DATAI_11_), .ZN(n14325) );
  MUX2_X1 U17507 ( .A(n14325), .B(n14324), .S(n20241), .Z(n20194) );
  OAI22_X1 U17508 ( .A1(n14375), .A2(n20194), .B1(n14389), .B2(n14326), .ZN(
        n14327) );
  AOI21_X1 U17509 ( .B1(n14377), .B2(BUF1_REG_27__SCAN_IN), .A(n14327), .ZN(
        n14329) );
  NAND2_X1 U17510 ( .A1(n14378), .A2(DATAI_27_), .ZN(n14328) );
  OAI211_X1 U17511 ( .C1(n14499), .C2(n14396), .A(n14329), .B(n14328), .ZN(
        P1_U2877) );
  OAI22_X1 U17512 ( .A1(n14375), .A2(n14393), .B1(n14389), .B2(n14330), .ZN(
        n14331) );
  AOI21_X1 U17513 ( .B1(n14377), .B2(BUF1_REG_26__SCAN_IN), .A(n14331), .ZN(
        n14333) );
  NAND2_X1 U17514 ( .A1(n14378), .A2(DATAI_26_), .ZN(n14332) );
  OAI211_X1 U17515 ( .C1(n14507), .C2(n14396), .A(n14333), .B(n14332), .ZN(
        P1_U2878) );
  OAI22_X1 U17516 ( .A1(n14375), .A2(n20191), .B1(n14389), .B2(n12910), .ZN(
        n14334) );
  AOI21_X1 U17517 ( .B1(n14377), .B2(BUF1_REG_25__SCAN_IN), .A(n14334), .ZN(
        n14336) );
  NAND2_X1 U17518 ( .A1(n14378), .A2(DATAI_25_), .ZN(n14335) );
  OAI211_X1 U17519 ( .C1(n14337), .C2(n14396), .A(n14336), .B(n14335), .ZN(
        P1_U2879) );
  OAI22_X1 U17520 ( .A1(n14375), .A2(n20188), .B1(n14389), .B2(n12905), .ZN(
        n14338) );
  AOI21_X1 U17521 ( .B1(n14377), .B2(BUF1_REG_24__SCAN_IN), .A(n14338), .ZN(
        n14340) );
  NAND2_X1 U17522 ( .A1(n14378), .A2(DATAI_24_), .ZN(n14339) );
  OAI211_X1 U17523 ( .C1(n14341), .C2(n14396), .A(n14340), .B(n14339), .ZN(
        P1_U2880) );
  NAND2_X1 U17524 ( .A1(n14258), .A2(n14342), .ZN(n14343) );
  AND2_X1 U17525 ( .A1(n14344), .A2(n14343), .ZN(n16079) );
  INV_X1 U17526 ( .A(n16079), .ZN(n14348) );
  OAI22_X1 U17527 ( .A1(n14375), .A2(n20296), .B1(n14389), .B2(n13134), .ZN(
        n14345) );
  AOI21_X1 U17528 ( .B1(n14377), .B2(BUF1_REG_23__SCAN_IN), .A(n14345), .ZN(
        n14347) );
  NAND2_X1 U17529 ( .A1(n14378), .A2(DATAI_23_), .ZN(n14346) );
  OAI211_X1 U17530 ( .C1(n14348), .C2(n14396), .A(n14347), .B(n14346), .ZN(
        P1_U2881) );
  OAI22_X1 U17531 ( .A1(n14375), .A2(n20287), .B1(n14389), .B2(n13143), .ZN(
        n14349) );
  AOI21_X1 U17532 ( .B1(n14377), .B2(BUF1_REG_22__SCAN_IN), .A(n14349), .ZN(
        n14351) );
  NAND2_X1 U17533 ( .A1(n14378), .A2(DATAI_22_), .ZN(n14350) );
  OAI211_X1 U17534 ( .C1(n16002), .C2(n14396), .A(n14351), .B(n14350), .ZN(
        P1_U2882) );
  OAI22_X1 U17535 ( .A1(n14375), .A2(n20282), .B1(n14389), .B2(n14352), .ZN(
        n14353) );
  AOI21_X1 U17536 ( .B1(n14377), .B2(BUF1_REG_21__SCAN_IN), .A(n14353), .ZN(
        n14355) );
  NAND2_X1 U17537 ( .A1(n14378), .A2(DATAI_21_), .ZN(n14354) );
  OAI211_X1 U17538 ( .C1(n14356), .C2(n14396), .A(n14355), .B(n14354), .ZN(
        P1_U2883) );
  OAI22_X1 U17539 ( .A1(n14375), .A2(n20278), .B1(n14389), .B2(n14357), .ZN(
        n14358) );
  AOI21_X1 U17540 ( .B1(n14377), .B2(BUF1_REG_20__SCAN_IN), .A(n14358), .ZN(
        n14360) );
  NAND2_X1 U17541 ( .A1(n14378), .A2(DATAI_20_), .ZN(n14359) );
  OAI211_X1 U17542 ( .C1(n14551), .C2(n14396), .A(n14360), .B(n14359), .ZN(
        P1_U2884) );
  OAI22_X1 U17543 ( .A1(n14375), .A2(n20274), .B1(n14389), .B2(n13138), .ZN(
        n14361) );
  AOI21_X1 U17544 ( .B1(n14377), .B2(BUF1_REG_19__SCAN_IN), .A(n14361), .ZN(
        n14363) );
  NAND2_X1 U17545 ( .A1(n14378), .A2(DATAI_19_), .ZN(n14362) );
  OAI211_X1 U17546 ( .C1(n14558), .C2(n14396), .A(n14363), .B(n14362), .ZN(
        P1_U2885) );
  OAI22_X1 U17547 ( .A1(n14375), .A2(n20269), .B1(n14389), .B2(n14364), .ZN(
        n14365) );
  AOI21_X1 U17548 ( .B1(n14377), .B2(BUF1_REG_18__SCAN_IN), .A(n14365), .ZN(
        n14367) );
  NAND2_X1 U17549 ( .A1(n14378), .A2(DATAI_18_), .ZN(n14366) );
  OAI211_X1 U17550 ( .C1(n16035), .C2(n14396), .A(n14367), .B(n14366), .ZN(
        P1_U2886) );
  INV_X1 U17551 ( .A(n14368), .ZN(n14369) );
  AOI21_X1 U17552 ( .B1(n14369), .B2(n9672), .A(n14277), .ZN(n16092) );
  INV_X1 U17553 ( .A(n16092), .ZN(n14374) );
  OAI22_X1 U17554 ( .A1(n14375), .A2(n20264), .B1(n14389), .B2(n14370), .ZN(
        n14371) );
  AOI21_X1 U17555 ( .B1(n14377), .B2(BUF1_REG_17__SCAN_IN), .A(n14371), .ZN(
        n14373) );
  NAND2_X1 U17556 ( .A1(n14378), .A2(DATAI_17_), .ZN(n14372) );
  OAI211_X1 U17557 ( .C1(n14374), .C2(n14396), .A(n14373), .B(n14372), .ZN(
        P1_U2887) );
  OAI22_X1 U17558 ( .A1(n14375), .A2(n20254), .B1(n14389), .B2(n13141), .ZN(
        n14376) );
  AOI21_X1 U17559 ( .B1(n14377), .B2(BUF1_REG_16__SCAN_IN), .A(n14376), .ZN(
        n14380) );
  NAND2_X1 U17560 ( .A1(n14378), .A2(DATAI_16_), .ZN(n14379) );
  OAI211_X1 U17561 ( .C1(n14579), .C2(n14396), .A(n14380), .B(n14379), .ZN(
        P1_U2888) );
  AOI21_X1 U17562 ( .B1(n14381), .B2(n14195), .A(n9696), .ZN(n16101) );
  INV_X1 U17563 ( .A(n16101), .ZN(n14384) );
  OAI222_X1 U17564 ( .A1(n14396), .A2(n14384), .B1(n14389), .B2(n14383), .C1(
        n14394), .C2(n14382), .ZN(P1_U2889) );
  OAI222_X1 U17565 ( .A1(n14595), .A2(n14396), .B1(n14385), .B2(n14389), .C1(
        n14394), .C2(n20203), .ZN(P1_U2890) );
  INV_X1 U17566 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14386) );
  OAI222_X1 U17567 ( .A1(n14611), .A2(n14396), .B1(n14386), .B2(n14389), .C1(
        n14394), .C2(n20200), .ZN(P1_U2891) );
  INV_X1 U17568 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14387) );
  OAI222_X1 U17569 ( .A1(n14388), .A2(n14396), .B1(n14387), .B2(n14389), .C1(
        n14394), .C2(n20197), .ZN(P1_U2892) );
  INV_X1 U17570 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14390) );
  OAI222_X1 U17571 ( .A1(n14391), .A2(n14396), .B1(n14390), .B2(n14389), .C1(
        n14394), .C2(n20194), .ZN(P1_U2893) );
  OAI222_X1 U17572 ( .A1(n14396), .A2(n14395), .B1(n14394), .B2(n14393), .C1(
        n14392), .C2(n14389), .ZN(P1_U2894) );
  NAND2_X1 U17573 ( .A1(n14398), .A2(n14397), .ZN(n14402) );
  OR2_X1 U17574 ( .A1(n14400), .A2(n14399), .ZN(n14401) );
  NAND2_X1 U17575 ( .A1(n14402), .A2(n14401), .ZN(n16136) );
  XNOR2_X1 U17576 ( .A(n14411), .B(n14412), .ZN(n14404) );
  NAND2_X1 U17577 ( .A1(n14404), .A2(n14435), .ZN(n14405) );
  XNOR2_X1 U17578 ( .A(n14406), .B(n16246), .ZN(n16137) );
  NAND2_X1 U17579 ( .A1(n16136), .A2(n16137), .ZN(n14408) );
  NAND2_X1 U17580 ( .A1(n14406), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14407) );
  NAND2_X1 U17581 ( .A1(n14408), .A2(n14407), .ZN(n16129) );
  BUF_X1 U17582 ( .A(n14409), .Z(n14432) );
  NAND3_X1 U17583 ( .A1(n14432), .A2(n14410), .A3(n14424), .ZN(n14416) );
  INV_X1 U17584 ( .A(n14411), .ZN(n14413) );
  NAND2_X1 U17585 ( .A1(n14413), .A2(n14412), .ZN(n14421) );
  XNOR2_X1 U17586 ( .A(n14421), .B(n14419), .ZN(n14414) );
  NAND2_X1 U17587 ( .A1(n14414), .A2(n14435), .ZN(n14415) );
  NAND2_X1 U17588 ( .A1(n14416), .A2(n14415), .ZN(n14417) );
  OR2_X1 U17589 ( .A1(n14417), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16131) );
  NAND2_X1 U17590 ( .A1(n16129), .A2(n16131), .ZN(n14418) );
  NAND2_X1 U17591 ( .A1(n14417), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16130) );
  NAND2_X1 U17592 ( .A1(n14418), .A2(n16130), .ZN(n16121) );
  INV_X1 U17593 ( .A(n14419), .ZN(n14420) );
  OR2_X1 U17594 ( .A1(n14421), .A2(n14420), .ZN(n14433) );
  XNOR2_X1 U17595 ( .A(n14433), .B(n14434), .ZN(n14422) );
  AND2_X1 U17596 ( .A1(n14422), .A2(n14435), .ZN(n14423) );
  AOI21_X1 U17597 ( .B1(n14425), .B2(n14424), .A(n14423), .ZN(n16123) );
  INV_X1 U17598 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16122) );
  NAND2_X1 U17599 ( .A1(n16123), .A2(n16122), .ZN(n14426) );
  INV_X1 U17600 ( .A(n16123), .ZN(n14427) );
  NAND2_X1 U17601 ( .A1(n14427), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14428) );
  NOR2_X1 U17602 ( .A1(n14430), .A2(n14429), .ZN(n14431) );
  NAND2_X2 U17603 ( .A1(n14432), .A2(n14431), .ZN(n14449) );
  INV_X1 U17604 ( .A(n14433), .ZN(n14436) );
  NAND3_X1 U17605 ( .A1(n14436), .A2(n14435), .A3(n14434), .ZN(n14437) );
  INV_X1 U17606 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16214) );
  NAND2_X1 U17607 ( .A1(n16112), .A2(n16214), .ZN(n14439) );
  XNOR2_X1 U17608 ( .A(n14449), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14603) );
  INV_X1 U17609 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14737) );
  NAND2_X1 U17610 ( .A1(n16112), .A2(n14737), .ZN(n14602) );
  NAND2_X1 U17611 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14584) );
  OAI21_X1 U17612 ( .B1(n14440), .B2(n14584), .A(n10059), .ZN(n14441) );
  AND2_X1 U17613 ( .A1(n14602), .A2(n14441), .ZN(n14442) );
  NAND2_X1 U17614 ( .A1(n14603), .A2(n14442), .ZN(n14570) );
  XNOR2_X1 U17615 ( .A(n14449), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14575) );
  NAND2_X1 U17616 ( .A1(n16112), .A2(n16155), .ZN(n14443) );
  NAND2_X1 U17617 ( .A1(n14575), .A2(n14443), .ZN(n14573) );
  INV_X1 U17618 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14446) );
  NOR2_X1 U17619 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14597) );
  AND2_X1 U17620 ( .A1(n14597), .A2(n14737), .ZN(n14444) );
  NOR2_X1 U17621 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16097) );
  AND2_X1 U17622 ( .A1(n16097), .A2(n16155), .ZN(n14445) );
  INV_X1 U17623 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14790) );
  NAND2_X1 U17624 ( .A1(n14790), .A2(n14538), .ZN(n14447) );
  NOR2_X2 U17625 ( .A1(n14566), .A2(n14447), .ZN(n14539) );
  NOR2_X1 U17626 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14448) );
  NAND2_X1 U17627 ( .A1(n14539), .A2(n14448), .ZN(n14450) );
  XNOR2_X1 U17628 ( .A(n14449), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14565) );
  NAND2_X1 U17629 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14759) );
  INV_X1 U17630 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14451) );
  NOR2_X1 U17631 ( .A1(n14759), .A2(n14451), .ZN(n14743) );
  AND2_X1 U17632 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14704) );
  AND2_X1 U17633 ( .A1(n14704), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14696) );
  INV_X1 U17634 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14717) );
  NAND3_X1 U17635 ( .A1(n14452), .A2(n14730), .A3(n14717), .ZN(n14481) );
  NAND2_X1 U17636 ( .A1(n9726), .A2(n14601), .ZN(n14453) );
  INV_X1 U17637 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21097) );
  INV_X1 U17638 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14682) );
  NAND2_X1 U17639 ( .A1(n21097), .A2(n14682), .ZN(n14679) );
  NOR2_X1 U17640 ( .A1(n14449), .A2(n14679), .ZN(n14454) );
  AND2_X1 U17641 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U17642 ( .A1(n16112), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14456) );
  XNOR2_X1 U17643 ( .A(n14457), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14657) );
  NAND2_X1 U17644 ( .A1(n16236), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14651) );
  NAND2_X1 U17645 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14458) );
  OAI211_X1 U17646 ( .C1(n14459), .C2(n16135), .A(n14651), .B(n14458), .ZN(
        n14460) );
  OAI21_X1 U17647 ( .B1(n14657), .B2(n20063), .A(n14462), .ZN(P1_U2968) );
  NAND2_X1 U17648 ( .A1(n14464), .A2(n16138), .ZN(n14465) );
  NAND2_X1 U17649 ( .A1(n16236), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14662) );
  OAI211_X1 U17650 ( .C1(n14466), .C2(n16144), .A(n14465), .B(n14662), .ZN(
        n14467) );
  AOI21_X1 U17651 ( .B1(n14468), .B2(n16140), .A(n14467), .ZN(n14469) );
  OAI21_X1 U17652 ( .B1(n14666), .B2(n20063), .A(n14469), .ZN(P1_U2969) );
  MUX2_X1 U17653 ( .A(n10070), .B(n14471), .S(n14470), .Z(n14473) );
  XNOR2_X1 U17654 ( .A(n14473), .B(n14472), .ZN(n14677) );
  NAND2_X1 U17655 ( .A1(n16236), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14671) );
  NAND2_X1 U17656 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14474) );
  OAI211_X1 U17657 ( .C1(n14475), .C2(n16135), .A(n14671), .B(n14474), .ZN(
        n14476) );
  AOI21_X1 U17658 ( .B1(n14477), .B2(n16140), .A(n14476), .ZN(n14478) );
  OAI21_X1 U17659 ( .B1(n14677), .B2(n20063), .A(n14478), .ZN(P1_U2970) );
  AND2_X1 U17660 ( .A1(n14479), .A2(n14601), .ZN(n14512) );
  NOR2_X1 U17661 ( .A1(n14481), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14484) );
  NAND2_X1 U17662 ( .A1(n14485), .A2(n21097), .ZN(n14483) );
  MUX2_X1 U17663 ( .A(n21097), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n16112), .Z(n14482) );
  OAI211_X1 U17664 ( .C1(n14485), .C2(n14484), .A(n14483), .B(n14482), .ZN(
        n14486) );
  XNOR2_X1 U17665 ( .A(n14486), .B(n14682), .ZN(n14686) );
  NAND2_X1 U17666 ( .A1(n14487), .A2(n16138), .ZN(n14488) );
  NAND2_X1 U17667 ( .A1(n16236), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14681) );
  OAI211_X1 U17668 ( .C1(n16144), .C2(n14489), .A(n14488), .B(n14681), .ZN(
        n14490) );
  AOI21_X1 U17669 ( .B1(n14491), .B2(n16140), .A(n14490), .ZN(n14492) );
  OAI21_X1 U17670 ( .B1(n20063), .B2(n14686), .A(n14492), .ZN(P1_U2971) );
  AND2_X1 U17671 ( .A1(n14696), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14640) );
  INV_X1 U17672 ( .A(n14640), .ZN(n14494) );
  NOR2_X1 U17673 ( .A1(n14493), .A2(n14494), .ZN(n14496) );
  MUX2_X1 U17674 ( .A(n14496), .B(n14495), .S(n14601), .Z(n14497) );
  XNOR2_X1 U17675 ( .A(n14497), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14694) );
  NAND2_X1 U17676 ( .A1(n16236), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14689) );
  OAI21_X1 U17677 ( .B1(n16144), .B2(n14498), .A(n14689), .ZN(n14501) );
  NOR2_X1 U17678 ( .A1(n14499), .A2(n20243), .ZN(n14500) );
  OAI21_X1 U17679 ( .B1(n20063), .B2(n14694), .A(n14503), .ZN(P1_U2972) );
  OAI21_X1 U17680 ( .B1(n14505), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14504), .ZN(n14703) );
  NAND2_X1 U17681 ( .A1(n16236), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14698) );
  OAI21_X1 U17682 ( .B1(n16144), .B2(n14506), .A(n14698), .ZN(n14509) );
  NOR2_X1 U17683 ( .A1(n14507), .A2(n20243), .ZN(n14508) );
  OAI21_X1 U17684 ( .B1(n20063), .B2(n14703), .A(n14511), .ZN(P1_U2973) );
  NOR2_X1 U17685 ( .A1(n20227), .A2(n20921), .ZN(n14708) );
  AOI21_X1 U17686 ( .B1(n16128), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14708), .ZN(n14513) );
  OAI21_X1 U17687 ( .B1(n14514), .B2(n16135), .A(n14513), .ZN(n14515) );
  AOI21_X1 U17688 ( .B1(n14516), .B2(n16140), .A(n14515), .ZN(n14517) );
  OAI21_X1 U17689 ( .B1(n20063), .B2(n14711), .A(n14517), .ZN(P1_U2974) );
  NOR2_X1 U17690 ( .A1(n14479), .A2(n14449), .ZN(n14519) );
  MUX2_X1 U17691 ( .A(n16112), .B(n14519), .S(n14518), .Z(n14520) );
  XNOR2_X1 U17692 ( .A(n14520), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14722) );
  INV_X1 U17693 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14523) );
  NAND2_X1 U17694 ( .A1(n14521), .A2(n16138), .ZN(n14522) );
  NAND2_X1 U17695 ( .A1(n16236), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14716) );
  OAI211_X1 U17696 ( .C1(n16144), .C2(n14523), .A(n14522), .B(n14716), .ZN(
        n14524) );
  AOI21_X1 U17697 ( .B1(n14525), .B2(n16140), .A(n14524), .ZN(n14526) );
  OAI21_X1 U17698 ( .B1(n14722), .B2(n20063), .A(n14526), .ZN(P1_U2975) );
  XNOR2_X1 U17699 ( .A(n14449), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14527) );
  XNOR2_X1 U17700 ( .A(n14479), .B(n14527), .ZN(n14735) );
  INV_X1 U17701 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20916) );
  NOR2_X1 U17702 ( .A1(n20227), .A2(n20916), .ZN(n14727) );
  AOI21_X1 U17703 ( .B1(n16128), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14727), .ZN(n14528) );
  OAI21_X1 U17704 ( .B1(n15989), .B2(n16135), .A(n14528), .ZN(n14529) );
  AOI21_X1 U17705 ( .B1(n16079), .B2(n16140), .A(n14529), .ZN(n14530) );
  OAI21_X1 U17706 ( .B1(n14735), .B2(n20063), .A(n14530), .ZN(P1_U2976) );
  NAND2_X1 U17707 ( .A1(n14532), .A2(n14531), .ZN(n14533) );
  XOR2_X1 U17708 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14533), .Z(
        n14751) );
  NAND2_X1 U17709 ( .A1(n16236), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14745) );
  OAI21_X1 U17710 ( .B1(n16144), .B2(n15997), .A(n14745), .ZN(n14535) );
  NOR2_X1 U17711 ( .A1(n16002), .A2(n20243), .ZN(n14534) );
  AOI211_X1 U17712 ( .C1(n16138), .C2(n16000), .A(n14535), .B(n14534), .ZN(
        n14536) );
  OAI21_X1 U17713 ( .B1(n20063), .B2(n14751), .A(n14536), .ZN(P1_U2977) );
  INV_X1 U17714 ( .A(n14537), .ZN(n14780) );
  NOR3_X1 U17715 ( .A1(n14780), .A2(n14601), .A3(n14538), .ZN(n14549) );
  NAND2_X1 U17716 ( .A1(n14539), .A2(n14601), .ZN(n14544) );
  NOR2_X1 U17717 ( .A1(n14544), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14547) );
  AOI21_X1 U17718 ( .B1(n14549), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14547), .ZN(n14540) );
  XOR2_X1 U17719 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n14540), .Z(
        n14757) );
  NOR2_X1 U17720 ( .A1(n20227), .A2(n20914), .ZN(n14753) );
  AOI21_X1 U17721 ( .B1(n16128), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14753), .ZN(n14541) );
  OAI21_X1 U17722 ( .B1(n16006), .B2(n16135), .A(n14541), .ZN(n14542) );
  AOI21_X1 U17723 ( .B1(n16011), .B2(n16140), .A(n14542), .ZN(n14543) );
  OAI21_X1 U17724 ( .B1(n14757), .B2(n20063), .A(n14543), .ZN(P1_U2978) );
  INV_X1 U17725 ( .A(n14544), .ZN(n14545) );
  NOR3_X1 U17726 ( .A1(n14549), .A2(n14545), .A3(n14548), .ZN(n14546) );
  AOI211_X1 U17727 ( .C1(n14549), .C2(n14548), .A(n14547), .B(n14546), .ZN(
        n14770) );
  NAND2_X1 U17728 ( .A1(n16236), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14758) );
  OAI21_X1 U17729 ( .B1(n16144), .B2(n14550), .A(n14758), .ZN(n14553) );
  NOR2_X1 U17730 ( .A1(n14551), .A2(n20243), .ZN(n14552) );
  AOI211_X1 U17731 ( .C1(n16138), .C2(n14554), .A(n14553), .B(n14552), .ZN(
        n14555) );
  OAI21_X1 U17732 ( .B1(n14770), .B2(n20063), .A(n14555), .ZN(P1_U2979) );
  NOR2_X1 U17733 ( .A1(n16112), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14556) );
  MUX2_X1 U17734 ( .A(n14556), .B(n16112), .S(n14537), .Z(n14557) );
  XNOR2_X1 U17735 ( .A(n14557), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14778) );
  INV_X1 U17736 ( .A(n14558), .ZN(n16027) );
  INV_X1 U17737 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n16024) );
  NOR2_X1 U17738 ( .A1(n20227), .A2(n16024), .ZN(n14771) );
  AOI21_X1 U17739 ( .B1(n16128), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n14771), .ZN(n14559) );
  OAI21_X1 U17740 ( .B1(n16030), .B2(n16135), .A(n14559), .ZN(n14560) );
  AOI21_X1 U17741 ( .B1(n16027), .B2(n16140), .A(n14560), .ZN(n14561) );
  OAI21_X1 U17742 ( .B1(n20063), .B2(n14778), .A(n14561), .ZN(P1_U2980) );
  NOR2_X1 U17743 ( .A1(n16144), .A2(n14562), .ZN(n14564) );
  INV_X1 U17744 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14563) );
  NOR2_X1 U17745 ( .A1(n20227), .A2(n14563), .ZN(n14792) );
  AOI211_X1 U17746 ( .C1(n16038), .C2(n16138), .A(n14564), .B(n14792), .ZN(
        n14568) );
  OR2_X1 U17747 ( .A1(n14566), .A2(n14565), .ZN(n14779) );
  NAND3_X1 U17748 ( .A1(n14780), .A2(n16141), .A3(n14779), .ZN(n14567) );
  OAI211_X1 U17749 ( .C1(n16035), .C2(n20243), .A(n14568), .B(n14567), .ZN(
        P1_U2981) );
  AND2_X1 U17750 ( .A1(n14596), .A2(n14569), .ZN(n14586) );
  NOR2_X1 U17751 ( .A1(n14586), .A2(n14570), .ZN(n16095) );
  INV_X1 U17752 ( .A(n14571), .ZN(n14572) );
  NOR2_X1 U17753 ( .A1(n16095), .A2(n14572), .ZN(n14574) );
  NOR2_X1 U17754 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14803) );
  NOR2_X1 U17755 ( .A1(n14574), .A2(n14803), .ZN(n14576) );
  OAI22_X1 U17756 ( .A1(n14576), .A2(n14575), .B1(n14574), .B2(n14573), .ZN(
        n14807) );
  INV_X1 U17757 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14577) );
  OAI22_X1 U17758 ( .A1(n16144), .A2(n14578), .B1(n20227), .B2(n14577), .ZN(
        n14581) );
  NOR2_X1 U17759 ( .A1(n14579), .A2(n20243), .ZN(n14580) );
  AOI211_X1 U17760 ( .C1(n16138), .C2(n14582), .A(n14581), .B(n14580), .ZN(
        n14583) );
  OAI21_X1 U17761 ( .B1(n20063), .B2(n14807), .A(n14583), .ZN(P1_U2983) );
  MUX2_X1 U17762 ( .A(n14440), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .S(
        n16112), .Z(n14588) );
  NAND2_X1 U17763 ( .A1(n16112), .A2(n14584), .ZN(n14599) );
  NAND3_X1 U17764 ( .A1(n14603), .A2(n14602), .A3(n14599), .ZN(n14585) );
  OAI22_X1 U17765 ( .A1(n14586), .A2(n14585), .B1(n16112), .B2(n16164), .ZN(
        n14587) );
  XOR2_X1 U17766 ( .A(n14588), .B(n14587), .Z(n14819) );
  NAND2_X1 U17767 ( .A1(n14819), .A2(n16141), .ZN(n14594) );
  INV_X1 U17768 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14589) );
  OR2_X1 U17769 ( .A1(n20227), .A2(n14589), .ZN(n14815) );
  INV_X1 U17770 ( .A(n14815), .ZN(n14592) );
  NOR2_X1 U17771 ( .A1(n16135), .A2(n14590), .ZN(n14591) );
  AOI211_X1 U17772 ( .C1(n16128), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n14592), .B(n14591), .ZN(n14593) );
  OAI211_X1 U17773 ( .C1(n20243), .C2(n14595), .A(n14594), .B(n14593), .ZN(
        P1_U2985) );
  INV_X1 U17774 ( .A(n14596), .ZN(n16113) );
  INV_X1 U17775 ( .A(n14597), .ZN(n14598) );
  AOI22_X1 U17776 ( .A1(n16113), .A2(n14599), .B1(n10070), .B2(n14598), .ZN(
        n16106) );
  INV_X1 U17777 ( .A(n14602), .ZN(n14600) );
  AOI21_X1 U17778 ( .B1(n14601), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14600), .ZN(n16105) );
  NAND2_X1 U17779 ( .A1(n16106), .A2(n16105), .ZN(n16104) );
  NAND2_X1 U17780 ( .A1(n16104), .A2(n14602), .ZN(n14604) );
  XNOR2_X1 U17781 ( .A(n14604), .B(n14603), .ZN(n16167) );
  NAND2_X1 U17782 ( .A1(n16167), .A2(n16141), .ZN(n14610) );
  INV_X1 U17783 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14606) );
  INV_X1 U17784 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14605) );
  OAI22_X1 U17785 ( .A1(n16144), .A2(n14606), .B1(n20227), .B2(n14605), .ZN(
        n14607) );
  AOI21_X1 U17786 ( .B1(n16138), .B2(n14608), .A(n14607), .ZN(n14609) );
  OAI211_X1 U17787 ( .C1(n20243), .C2(n14611), .A(n14610), .B(n14609), .ZN(
        P1_U2986) );
  NAND2_X1 U17788 ( .A1(n14612), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14614) );
  XNOR2_X1 U17789 ( .A(n16113), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14613) );
  MUX2_X1 U17790 ( .A(n14614), .B(n14613), .S(n16112), .Z(n14615) );
  OR3_X1 U17791 ( .A1(n14612), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n14449), .ZN(n16114) );
  NAND2_X1 U17792 ( .A1(n14615), .A2(n16114), .ZN(n16203) );
  INV_X1 U17793 ( .A(n16203), .ZN(n14621) );
  AOI22_X1 U17794 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n16236), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14616) );
  OAI21_X1 U17795 ( .B1(n16135), .B2(n14617), .A(n14616), .ZN(n14618) );
  AOI21_X1 U17796 ( .B1(n14619), .B2(n16140), .A(n14618), .ZN(n14620) );
  OAI21_X1 U17797 ( .B1(n14621), .B2(n20063), .A(n14620), .ZN(P1_U2989) );
  XNOR2_X1 U17798 ( .A(n14449), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14622) );
  XNOR2_X1 U17799 ( .A(n14623), .B(n14622), .ZN(n16211) );
  NAND2_X1 U17800 ( .A1(n16211), .A2(n16141), .ZN(n14626) );
  NAND2_X1 U17801 ( .A1(n16236), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n16208) );
  OAI21_X1 U17802 ( .B1(n16144), .B2(n11383), .A(n16208), .ZN(n14624) );
  AOI21_X1 U17803 ( .B1(n16138), .B2(n20081), .A(n14624), .ZN(n14625) );
  OAI211_X1 U17804 ( .C1(n20243), .C2(n20086), .A(n14626), .B(n14625), .ZN(
        P1_U2990) );
  XNOR2_X1 U17805 ( .A(n14628), .B(n16228), .ZN(n14629) );
  XNOR2_X1 U17806 ( .A(n14627), .B(n14629), .ZN(n16222) );
  OAI22_X1 U17807 ( .A1(n16144), .A2(n14630), .B1(n20227), .B2(n13592), .ZN(
        n14633) );
  NOR2_X1 U17808 ( .A1(n14631), .A2(n20243), .ZN(n14632) );
  AOI211_X1 U17809 ( .C1(n16138), .C2(n14634), .A(n14633), .B(n14632), .ZN(
        n14635) );
  OAI21_X1 U17810 ( .B1(n20063), .B2(n16222), .A(n14635), .ZN(P1_U2991) );
  NAND2_X1 U17811 ( .A1(n20226), .A2(n16216), .ZN(n16219) );
  NOR2_X1 U17812 ( .A1(n16246), .A2(n16219), .ZN(n16196) );
  NOR3_X1 U17813 ( .A1(n16228), .A2(n16122), .A3(n16225), .ZN(n16195) );
  INV_X1 U17814 ( .A(n16195), .ZN(n14810) );
  INV_X1 U17815 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16207) );
  NOR2_X1 U17816 ( .A1(n16207), .A2(n16214), .ZN(n14811) );
  INV_X1 U17817 ( .A(n14811), .ZN(n16204) );
  NOR2_X1 U17818 ( .A1(n14810), .A2(n16204), .ZN(n14636) );
  NAND2_X1 U17819 ( .A1(n16196), .A2(n14636), .ZN(n16173) );
  NAND3_X1 U17820 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14812) );
  NOR2_X1 U17821 ( .A1(n16173), .A2(n14812), .ZN(n14782) );
  NAND2_X1 U17822 ( .A1(n20223), .A2(n14782), .ZN(n14638) );
  NAND3_X1 U17823 ( .A1(n16216), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n20224), .ZN(n14808) );
  NAND2_X1 U17824 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14636), .ZN(
        n16174) );
  NOR3_X1 U17825 ( .A1(n14737), .A2(n14808), .A3(n16174), .ZN(n14736) );
  NAND3_X1 U17826 ( .A1(n16175), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n14736), .ZN(n14637) );
  NAND2_X1 U17827 ( .A1(n14638), .A2(n14637), .ZN(n14802) );
  NAND2_X1 U17828 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16145) );
  OR3_X1 U17829 ( .A1(n14440), .A2(n14446), .A3(n16145), .ZN(n14789) );
  NOR2_X1 U17830 ( .A1(n14790), .A2(n14789), .ZN(n14641) );
  AND3_X1 U17831 ( .A1(n14641), .A2(n14743), .A3(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14639) );
  NAND3_X1 U17832 ( .A1(n14687), .A2(n14670), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14658) );
  INV_X1 U17833 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14821) );
  NAND2_X1 U17834 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14653) );
  AND2_X1 U17835 ( .A1(n14782), .A2(n14641), .ZN(n14741) );
  AND2_X1 U17836 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14641), .ZN(
        n14740) );
  NAND2_X1 U17837 ( .A1(n14736), .A2(n14740), .ZN(n14642) );
  NAND2_X1 U17838 ( .A1(n16175), .A2(n14642), .ZN(n14643) );
  OAI211_X1 U17839 ( .C1(n16197), .C2(n14741), .A(n16171), .B(n14643), .ZN(
        n14772) );
  OR2_X1 U17840 ( .A1(n14772), .A2(n14759), .ZN(n14645) );
  NAND2_X1 U17841 ( .A1(n14798), .A2(n16171), .ZN(n14644) );
  NAND2_X1 U17842 ( .A1(n14645), .A2(n14644), .ZN(n14744) );
  NAND2_X1 U17843 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14646) );
  NAND2_X1 U17844 ( .A1(n16221), .A2(n14646), .ZN(n14647) );
  NAND2_X1 U17845 ( .A1(n14744), .A2(n14647), .ZN(n14648) );
  AOI21_X1 U17846 ( .B1(n16175), .B2(n14730), .A(n14648), .ZN(n14713) );
  OAI21_X1 U17847 ( .B1(n14696), .B2(n14798), .A(n14713), .ZN(n14695) );
  INV_X1 U17848 ( .A(n14648), .ZN(n14731) );
  NAND2_X1 U17849 ( .A1(n14731), .A2(n14798), .ZN(n14669) );
  OAI21_X1 U17850 ( .B1(n14695), .B2(n14699), .A(n14669), .ZN(n14690) );
  NAND2_X1 U17851 ( .A1(n14690), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14668) );
  INV_X1 U17852 ( .A(n14670), .ZN(n14678) );
  NOR2_X1 U17853 ( .A1(n14668), .A2(n14678), .ZN(n14650) );
  INV_X1 U17854 ( .A(n14669), .ZN(n14649) );
  OAI21_X1 U17855 ( .B1(n14650), .B2(n14649), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14659) );
  NAND3_X1 U17856 ( .A1(n14659), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14669), .ZN(n14652) );
  OAI211_X1 U17857 ( .C1(n14658), .C2(n14653), .A(n14652), .B(n14651), .ZN(
        n14654) );
  AOI21_X1 U17858 ( .B1(n14655), .B2(n16243), .A(n14654), .ZN(n14656) );
  OAI21_X1 U17859 ( .B1(n14657), .B2(n20230), .A(n14656), .ZN(P1_U3000) );
  INV_X1 U17860 ( .A(n14658), .ZN(n14660) );
  OAI21_X1 U17861 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14660), .A(
        n14659), .ZN(n14661) );
  OAI211_X1 U17862 ( .C1(n14663), .C2(n16200), .A(n14662), .B(n14661), .ZN(
        n14664) );
  INV_X1 U17863 ( .A(n14664), .ZN(n14665) );
  OAI21_X1 U17864 ( .B1(n14666), .B2(n20230), .A(n14665), .ZN(P1_U3001) );
  INV_X1 U17865 ( .A(n14667), .ZN(n14675) );
  AOI21_X1 U17866 ( .B1(n14678), .B2(n14669), .A(n14668), .ZN(n14673) );
  AOI21_X1 U17867 ( .B1(n14687), .B2(n14670), .A(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14672) );
  OAI21_X1 U17868 ( .B1(n14673), .B2(n14672), .A(n14671), .ZN(n14674) );
  AOI21_X1 U17869 ( .B1(n14675), .B2(n16243), .A(n14674), .ZN(n14676) );
  OAI21_X1 U17870 ( .B1(n14677), .B2(n20230), .A(n14676), .ZN(P1_U3002) );
  NAND3_X1 U17871 ( .A1(n14687), .A2(n14679), .A3(n14678), .ZN(n14680) );
  OAI211_X1 U17872 ( .C1(n14690), .C2(n14682), .A(n14681), .B(n14680), .ZN(
        n14683) );
  AOI21_X1 U17873 ( .B1(n14684), .B2(n16243), .A(n14683), .ZN(n14685) );
  OAI21_X1 U17874 ( .B1(n14686), .B2(n20230), .A(n14685), .ZN(P1_U3003) );
  NAND2_X1 U17875 ( .A1(n14687), .A2(n21097), .ZN(n14688) );
  OAI211_X1 U17876 ( .C1(n14690), .C2(n21097), .A(n14689), .B(n14688), .ZN(
        n14691) );
  AOI21_X1 U17877 ( .B1(n14692), .B2(n16243), .A(n14691), .ZN(n14693) );
  OAI21_X1 U17878 ( .B1(n14694), .B2(n20230), .A(n14693), .ZN(P1_U3004) );
  INV_X1 U17879 ( .A(n14695), .ZN(n14706) );
  NAND3_X1 U17880 ( .A1(n14728), .A2(n14696), .A3(n14699), .ZN(n14697) );
  OAI211_X1 U17881 ( .C1(n14706), .C2(n14699), .A(n14698), .B(n14697), .ZN(
        n14700) );
  AOI21_X1 U17882 ( .B1(n14701), .B2(n16243), .A(n14700), .ZN(n14702) );
  OAI21_X1 U17883 ( .B1(n14703), .B2(n20230), .A(n14702), .ZN(P1_U3005) );
  AOI21_X1 U17884 ( .B1(n14728), .B2(n14704), .A(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14705) );
  NOR2_X1 U17885 ( .A1(n14706), .A2(n14705), .ZN(n14707) );
  AOI211_X1 U17886 ( .C1(n14709), .C2(n16243), .A(n14708), .B(n14707), .ZN(
        n14710) );
  OAI21_X1 U17887 ( .B1(n14711), .B2(n20230), .A(n14710), .ZN(P1_U3006) );
  INV_X1 U17888 ( .A(n14712), .ZN(n14720) );
  INV_X1 U17889 ( .A(n14713), .ZN(n14714) );
  AOI21_X1 U17890 ( .B1(n20223), .B2(n14730), .A(n14714), .ZN(n14718) );
  NAND3_X1 U17891 ( .A1(n14728), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14717), .ZN(n14715) );
  OAI211_X1 U17892 ( .C1(n14718), .C2(n14717), .A(n14716), .B(n14715), .ZN(
        n14719) );
  AOI21_X1 U17893 ( .B1(n14720), .B2(n16243), .A(n14719), .ZN(n14721) );
  OAI21_X1 U17894 ( .B1(n14722), .B2(n20230), .A(n14721), .ZN(P1_U3007) );
  OR2_X1 U17895 ( .A1(n14724), .A2(n14723), .ZN(n14725) );
  NAND2_X1 U17896 ( .A1(n14726), .A2(n14725), .ZN(n16077) );
  INV_X1 U17897 ( .A(n16077), .ZN(n14733) );
  AOI21_X1 U17898 ( .B1(n14728), .B2(n14730), .A(n14727), .ZN(n14729) );
  OAI21_X1 U17899 ( .B1(n14731), .B2(n14730), .A(n14729), .ZN(n14732) );
  AOI21_X1 U17900 ( .B1(n14733), .B2(n16243), .A(n14732), .ZN(n14734) );
  OAI21_X1 U17901 ( .B1(n14735), .B2(n20230), .A(n14734), .ZN(P1_U3008) );
  INV_X1 U17902 ( .A(n16005), .ZN(n14749) );
  INV_X1 U17903 ( .A(n14783), .ZN(n14760) );
  INV_X1 U17904 ( .A(n14736), .ZN(n14784) );
  NOR2_X1 U17905 ( .A1(n20229), .A2(n14784), .ZN(n14739) );
  NOR3_X1 U17906 ( .A1(n14737), .A2(n16178), .A3(n16173), .ZN(n16162) );
  NAND2_X1 U17907 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16162), .ZN(
        n14781) );
  NOR2_X1 U17908 ( .A1(n14788), .A2(n14781), .ZN(n14738) );
  OR2_X1 U17909 ( .A1(n14739), .A2(n14738), .ZN(n16163) );
  AND2_X1 U17910 ( .A1(n16163), .A2(n14740), .ZN(n14761) );
  AOI21_X1 U17911 ( .B1(n14741), .B2(n14760), .A(n14761), .ZN(n14774) );
  INV_X1 U17912 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14742) );
  NAND2_X1 U17913 ( .A1(n14743), .A2(n14742), .ZN(n14747) );
  NOR3_X1 U17914 ( .A1(n14774), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n14759), .ZN(n14752) );
  INV_X1 U17915 ( .A(n14744), .ZN(n14754) );
  OAI21_X1 U17916 ( .B1(n14752), .B2(n14754), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14746) );
  OAI211_X1 U17917 ( .C1(n14774), .C2(n14747), .A(n14746), .B(n14745), .ZN(
        n14748) );
  AOI21_X1 U17918 ( .B1(n14749), .B2(n16243), .A(n14748), .ZN(n14750) );
  OAI21_X1 U17919 ( .B1(n14751), .B2(n20230), .A(n14750), .ZN(P1_U3009) );
  AOI211_X1 U17920 ( .C1(n14754), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14753), .B(n14752), .ZN(n14756) );
  NAND2_X1 U17921 ( .A1(n16010), .A2(n16243), .ZN(n14755) );
  OAI211_X1 U17922 ( .C1(n14757), .C2(n20230), .A(n14756), .B(n14755), .ZN(
        P1_U3010) );
  INV_X1 U17923 ( .A(n14758), .ZN(n14767) );
  INV_X1 U17924 ( .A(n14772), .ZN(n14765) );
  OAI21_X1 U17925 ( .B1(n14761), .B2(n14760), .A(n14759), .ZN(n14764) );
  INV_X1 U17926 ( .A(n14774), .ZN(n14762) );
  AOI21_X1 U17927 ( .B1(n14762), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14763) );
  AOI21_X1 U17928 ( .B1(n14765), .B2(n14764), .A(n14763), .ZN(n14766) );
  AOI211_X1 U17929 ( .C1(n14768), .C2(n16243), .A(n14767), .B(n14766), .ZN(
        n14769) );
  OAI21_X1 U17930 ( .B1(n14770), .B2(n20230), .A(n14769), .ZN(P1_U3011) );
  AOI21_X1 U17931 ( .B1(n14772), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14771), .ZN(n14773) );
  OAI21_X1 U17932 ( .B1(n14774), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14773), .ZN(n14775) );
  AOI21_X1 U17933 ( .B1(n14776), .B2(n16243), .A(n14775), .ZN(n14777) );
  OAI21_X1 U17934 ( .B1(n14778), .B2(n20230), .A(n14777), .ZN(P1_U3012) );
  NAND3_X1 U17935 ( .A1(n14780), .A2(n16249), .A3(n14779), .ZN(n14795) );
  NOR2_X1 U17936 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14789), .ZN(
        n14793) );
  INV_X1 U17937 ( .A(n14781), .ZN(n14787) );
  NOR2_X1 U17938 ( .A1(n14783), .A2(n14782), .ZN(n16161) );
  AOI21_X1 U17939 ( .B1(n16175), .B2(n14784), .A(n16161), .ZN(n14786) );
  OAI211_X1 U17940 ( .C1(n14788), .C2(n14787), .A(n14786), .B(n14785), .ZN(
        n16166) );
  AOI21_X1 U17941 ( .B1(n16164), .B2(n16163), .A(n16166), .ZN(n14797) );
  INV_X1 U17942 ( .A(n14797), .ZN(n14813) );
  AOI21_X1 U17943 ( .B1(n16221), .B2(n14789), .A(n14813), .ZN(n16146) );
  NOR2_X1 U17944 ( .A1(n16146), .A2(n14790), .ZN(n14791) );
  AOI211_X1 U17945 ( .C1(n14793), .C2(n14802), .A(n14792), .B(n14791), .ZN(
        n14794) );
  OAI211_X1 U17946 ( .C1(n16200), .C2(n16034), .A(n14795), .B(n14794), .ZN(
        P1_U3013) );
  INV_X1 U17947 ( .A(n14796), .ZN(n14801) );
  OAI21_X1 U17948 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14798), .A(
        n14797), .ZN(n16157) );
  NAND2_X1 U17949 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16157), .ZN(
        n14799) );
  OAI21_X1 U17950 ( .B1(n20227), .B2(n14577), .A(n14799), .ZN(n14800) );
  AOI21_X1 U17951 ( .B1(n14801), .B2(n16243), .A(n14800), .ZN(n14806) );
  INV_X1 U17952 ( .A(n16145), .ZN(n14804) );
  NAND2_X1 U17953 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14802), .ZN(
        n16154) );
  OR3_X1 U17954 ( .A1(n14804), .A2(n14803), .A3(n16154), .ZN(n14805) );
  OAI211_X1 U17955 ( .C1(n14807), .C2(n20230), .A(n14806), .B(n14805), .ZN(
        P1_U3015) );
  INV_X1 U17956 ( .A(n14808), .ZN(n16172) );
  NAND2_X1 U17957 ( .A1(n16172), .A2(n14809), .ZN(n16241) );
  NOR2_X1 U17958 ( .A1(n14810), .A2(n16241), .ZN(n16210) );
  NAND2_X1 U17959 ( .A1(n14811), .A2(n16210), .ZN(n16194) );
  NOR2_X1 U17960 ( .A1(n14812), .A2(n16194), .ZN(n14814) );
  MUX2_X1 U17961 ( .A(n14814), .B(n14813), .S(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n14818) );
  OAI21_X1 U17962 ( .B1(n14816), .B2(n16200), .A(n14815), .ZN(n14817) );
  AOI211_X1 U17963 ( .C1(n14819), .C2(n16249), .A(n14818), .B(n14817), .ZN(
        n14820) );
  INV_X1 U17964 ( .A(n14820), .ZN(P1_U3017) );
  AOI22_X1 U17965 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14822), .B2(n14821), .ZN(
        n14836) );
  INV_X1 U17966 ( .A(n14823), .ZN(n15934) );
  INV_X1 U17967 ( .A(n20667), .ZN(n20739) );
  NAND2_X1 U17968 ( .A1(n20739), .A2(n14824), .ZN(n14827) );
  NAND3_X1 U17969 ( .A1(n14825), .A2(n14828), .A3(n14829), .ZN(n14826) );
  OAI211_X1 U17970 ( .C1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n15934), .A(
        n14827), .B(n14826), .ZN(n15935) );
  NAND2_X1 U17971 ( .A1(n15935), .A2(n16255), .ZN(n14831) );
  NAND3_X1 U17972 ( .A1(n14829), .A2(n15956), .A3(n14828), .ZN(n14830) );
  OAI211_X1 U17973 ( .C1(n14836), .C2(n14832), .A(n14831), .B(n14830), .ZN(
        n14834) );
  INV_X1 U17974 ( .A(n14833), .ZN(n16259) );
  MUX2_X1 U17975 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14834), .S(
        n16259), .Z(P1_U3473) );
  INV_X1 U17976 ( .A(n16255), .ZN(n14839) );
  AOI22_X1 U17977 ( .A1(n14837), .A2(n15956), .B1(n14836), .B2(n14835), .ZN(
        n14838) );
  OAI21_X1 U17978 ( .B1(n14840), .B2(n14839), .A(n14838), .ZN(n14841) );
  MUX2_X1 U17979 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14841), .S(
        n16259), .Z(P1_U3472) );
  OAI21_X1 U17980 ( .B1(n12215), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19938), 
        .ZN(n14842) );
  NAND3_X1 U17981 ( .A1(n14843), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14842), 
        .ZN(n14845) );
  OAI22_X1 U17982 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16422), .B1(n19943), 
        .B2(n20035), .ZN(n14844) );
  NAND2_X1 U17983 ( .A1(n14845), .A2(n14844), .ZN(n14850) );
  NOR2_X1 U17984 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14846), .ZN(n19325) );
  INV_X1 U17985 ( .A(n19325), .ZN(n19280) );
  OAI21_X1 U17986 ( .B1(n16419), .B2(n20035), .A(n19632), .ZN(n14847) );
  OAI211_X1 U17987 ( .C1(n19943), .C2(n19280), .A(n14848), .B(n14847), .ZN(
        n14849) );
  MUX2_X1 U17988 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n14850), .S(n14849), 
        .Z(P2_U3610) );
  AOI211_X1 U17989 ( .C1(n14851), .C2(n14852), .A(n9752), .B(n19929), .ZN(
        n14853) );
  INV_X1 U17990 ( .A(n14853), .ZN(n14859) );
  AOI22_X1 U17991 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19198), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19170), .ZN(n14855) );
  NAND2_X1 U17992 ( .A1(n19183), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14854) );
  OAI211_X1 U17993 ( .C1(n15033), .C2(n19154), .A(n14855), .B(n14854), .ZN(
        n14856) );
  AOI21_X1 U17994 ( .B1(n19153), .B2(n14857), .A(n14856), .ZN(n14858) );
  OAI211_X1 U17995 ( .C1(n14938), .C2(n19174), .A(n14859), .B(n14858), .ZN(
        P2_U2826) );
  INV_X1 U17996 ( .A(n15327), .ZN(n14942) );
  AOI211_X1 U17997 ( .C1(n14862), .C2(n14861), .A(n14860), .B(n19929), .ZN(
        n14863) );
  INV_X1 U17998 ( .A(n14863), .ZN(n14873) );
  INV_X1 U17999 ( .A(n14864), .ZN(n14871) );
  NAND2_X1 U18000 ( .A1(n12605), .A2(n14865), .ZN(n14866) );
  NAND2_X1 U18001 ( .A1(n14867), .A2(n14866), .ZN(n15322) );
  NAND2_X1 U18002 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19183), .ZN(n14869) );
  AOI22_X1 U18003 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19198), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19170), .ZN(n14868) );
  OAI211_X1 U18004 ( .C1(n15322), .C2(n19154), .A(n14869), .B(n14868), .ZN(
        n14870) );
  AOI21_X1 U18005 ( .B1(n14871), .B2(n19153), .A(n14870), .ZN(n14872) );
  OAI211_X1 U18006 ( .C1(n19174), .C2(n14942), .A(n14873), .B(n14872), .ZN(
        P2_U2827) );
  AOI211_X1 U18007 ( .C1(n9688), .C2(n15128), .A(n19929), .B(n14874), .ZN(
        n14875) );
  INV_X1 U18008 ( .A(n14875), .ZN(n14885) );
  AND2_X1 U18009 ( .A1(n15062), .A2(n14876), .ZN(n14877) );
  NOR2_X1 U18010 ( .A1(n15048), .A2(n14877), .ZN(n15358) );
  AOI22_X1 U18011 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19198), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19170), .ZN(n14878) );
  OAI21_X1 U18012 ( .B1(n19156), .B2(n14962), .A(n14878), .ZN(n14883) );
  NAND2_X1 U18013 ( .A1(n14879), .A2(n14880), .ZN(n14881) );
  NAND2_X1 U18014 ( .A1(n14951), .A2(n14881), .ZN(n15362) );
  NOR2_X1 U18015 ( .A1(n15362), .A2(n19174), .ZN(n14882) );
  AOI211_X1 U18016 ( .C1(n19185), .C2(n15358), .A(n14883), .B(n14882), .ZN(
        n14884) );
  OAI211_X1 U18017 ( .C1(n19194), .C2(n14886), .A(n14885), .B(n14884), .ZN(
        P2_U2830) );
  NOR2_X1 U18018 ( .A1(n14904), .A2(n14887), .ZN(n14888) );
  OR2_X1 U18019 ( .A1(n14969), .A2(n14888), .ZN(n15142) );
  NAND2_X1 U18020 ( .A1(n14909), .A2(n14890), .ZN(n14891) );
  NAND2_X1 U18021 ( .A1(n9718), .A2(n14891), .ZN(n15383) );
  INV_X1 U18022 ( .A(n15383), .ZN(n14895) );
  AOI22_X1 U18023 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19198), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19170), .ZN(n14892) );
  OAI21_X1 U18024 ( .B1(n19156), .B2(n14893), .A(n14892), .ZN(n14894) );
  AOI21_X1 U18025 ( .B1(n14895), .B2(n19185), .A(n14894), .ZN(n14896) );
  OAI21_X1 U18026 ( .B1(n15142), .B2(n19174), .A(n14896), .ZN(n14900) );
  AOI211_X1 U18027 ( .C1(n14898), .C2(n15143), .A(n19929), .B(n14897), .ZN(
        n14899) );
  AOI211_X1 U18028 ( .C1(n19153), .C2(n14901), .A(n14900), .B(n14899), .ZN(
        n14902) );
  INV_X1 U18029 ( .A(n14902), .ZN(P2_U2832) );
  AND2_X1 U18030 ( .A1(n9694), .A2(n14903), .ZN(n14905) );
  OR2_X1 U18031 ( .A1(n14905), .A2(n14904), .ZN(n15401) );
  OR2_X1 U18032 ( .A1(n14907), .A2(n14906), .ZN(n14908) );
  NAND2_X1 U18033 ( .A1(n14909), .A2(n14908), .ZN(n15395) );
  AOI22_X1 U18034 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19198), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19170), .ZN(n14914) );
  INV_X1 U18035 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n14910) );
  OAI22_X1 U18036 ( .A1(n14911), .A2(n19194), .B1(n19156), .B2(n14910), .ZN(
        n14912) );
  INV_X1 U18037 ( .A(n14912), .ZN(n14913) );
  OAI211_X1 U18038 ( .C1(n15395), .C2(n19154), .A(n14914), .B(n14913), .ZN(
        n14918) );
  AOI211_X1 U18039 ( .C1(n14916), .C2(n9768), .A(n14915), .B(n19929), .ZN(
        n14917) );
  NOR2_X1 U18040 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  OAI21_X1 U18041 ( .B1(n15401), .B2(n19174), .A(n14919), .ZN(P2_U2833) );
  NAND2_X1 U18042 ( .A1(n14920), .A2(n14921), .ZN(n14922) );
  AND2_X1 U18043 ( .A1(n15094), .A2(n14922), .ZN(n19210) );
  NAND2_X1 U18044 ( .A1(n19185), .A2(n19210), .ZN(n14928) );
  NOR2_X1 U18045 ( .A1(n19162), .A2(n14923), .ZN(n19047) );
  XNOR2_X1 U18046 ( .A(n19047), .B(n15226), .ZN(n14926) );
  AOI22_X1 U18047 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19198), .B1(
        P2_EBX_REG_16__SCAN_IN), .B2(n19183), .ZN(n14924) );
  INV_X1 U18048 ( .A(n14924), .ZN(n14925) );
  AOI211_X1 U18049 ( .C1(n19178), .C2(n14926), .A(n14925), .B(n19038), .ZN(
        n14927) );
  OAI211_X1 U18050 ( .C1(n19188), .C2(n19970), .A(n14928), .B(n14927), .ZN(
        n14929) );
  AOI21_X1 U18051 ( .B1(n15477), .B2(n19190), .A(n14929), .ZN(n14930) );
  OAI21_X1 U18052 ( .B1(n14931), .B2(n19194), .A(n14930), .ZN(P2_U2839) );
  NAND2_X1 U18053 ( .A1(n16279), .A2(n14998), .ZN(n14932) );
  OAI21_X1 U18054 ( .B1(n14998), .B2(n16273), .A(n14932), .ZN(P2_U2856) );
  INV_X1 U18055 ( .A(n14933), .ZN(n15027) );
  NAND2_X1 U18056 ( .A1(n14935), .A2(n14934), .ZN(n15026) );
  NAND3_X1 U18057 ( .A1(n15027), .A2(n15012), .A3(n15026), .ZN(n14937) );
  NAND2_X1 U18058 ( .A1(n15015), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14936) );
  OAI211_X1 U18059 ( .C1(n15004), .C2(n14938), .A(n14937), .B(n14936), .ZN(
        P2_U2858) );
  NAND2_X1 U18060 ( .A1(n13930), .A2(n14939), .ZN(n14941) );
  XNOR2_X1 U18061 ( .A(n14941), .B(n14940), .ZN(n15039) );
  NOR2_X1 U18062 ( .A1(n14942), .A2(n15004), .ZN(n14943) );
  AOI21_X1 U18063 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15004), .A(n14943), .ZN(
        n14944) );
  OAI21_X1 U18064 ( .B1(n15039), .B2(n15025), .A(n14944), .ZN(P2_U2859) );
  NAND2_X1 U18065 ( .A1(n15040), .A2(n15012), .ZN(n14949) );
  NAND2_X1 U18066 ( .A1(n15015), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14948) );
  OAI211_X1 U18067 ( .C1(n15340), .C2(n15004), .A(n14949), .B(n14948), .ZN(
        P2_U2860) );
  NAND2_X1 U18068 ( .A1(n14951), .A2(n14950), .ZN(n14952) );
  NAND2_X1 U18069 ( .A1(n14953), .A2(n14952), .ZN(n16294) );
  AOI21_X1 U18070 ( .B1(n14956), .B2(n14955), .A(n14954), .ZN(n15046) );
  NAND2_X1 U18071 ( .A1(n15046), .A2(n15012), .ZN(n14958) );
  NAND2_X1 U18072 ( .A1(n15015), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14957) );
  OAI211_X1 U18073 ( .C1(n16294), .C2(n15004), .A(n14958), .B(n14957), .ZN(
        P2_U2861) );
  OAI21_X1 U18074 ( .B1(n14959), .B2(n14961), .A(n14960), .ZN(n15058) );
  MUX2_X1 U18075 ( .A(n15362), .B(n14962), .S(n15015), .Z(n14963) );
  OAI21_X1 U18076 ( .B1(n15058), .B2(n15025), .A(n14963), .ZN(P2_U2862) );
  AOI21_X1 U18077 ( .B1(n14964), .B2(n14965), .A(n9679), .ZN(n14966) );
  XOR2_X1 U18078 ( .A(n14967), .B(n14966), .Z(n15059) );
  OR2_X1 U18079 ( .A1(n14969), .A2(n14968), .ZN(n14970) );
  NAND2_X1 U18080 ( .A1(n14879), .A2(n14970), .ZN(n16301) );
  NOR2_X1 U18081 ( .A1(n16301), .A2(n15004), .ZN(n14971) );
  AOI21_X1 U18082 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15004), .A(n14971), .ZN(
        n14972) );
  OAI21_X1 U18083 ( .B1(n15059), .B2(n15025), .A(n14972), .ZN(P2_U2863) );
  AOI21_X1 U18084 ( .B1(n14975), .B2(n14974), .A(n14973), .ZN(n15071) );
  NAND2_X1 U18085 ( .A1(n15071), .A2(n15012), .ZN(n14977) );
  NAND2_X1 U18086 ( .A1(n15015), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14976) );
  OAI211_X1 U18087 ( .C1(n15142), .C2(n15004), .A(n14977), .B(n14976), .ZN(
        P2_U2864) );
  AOI21_X1 U18088 ( .B1(n14980), .B2(n14978), .A(n14979), .ZN(n15077) );
  NAND2_X1 U18089 ( .A1(n15077), .A2(n15012), .ZN(n14982) );
  NAND2_X1 U18090 ( .A1(n15015), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14981) );
  OAI211_X1 U18091 ( .C1(n15401), .C2(n15004), .A(n14982), .B(n14981), .ZN(
        P2_U2865) );
  OAI21_X1 U18092 ( .B1(n14983), .B2(n14984), .A(n14978), .ZN(n15083) );
  NAND2_X1 U18093 ( .A1(n15015), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14988) );
  NAND2_X1 U18094 ( .A1(n9742), .A2(n14985), .ZN(n14986) );
  NAND2_X1 U18095 ( .A1(n9694), .A2(n14986), .ZN(n18979) );
  OR2_X1 U18096 ( .A1(n18979), .A2(n15004), .ZN(n14987) );
  OAI211_X1 U18097 ( .C1(n15083), .C2(n15025), .A(n14988), .B(n14987), .ZN(
        P2_U2866) );
  AND2_X1 U18098 ( .A1(n14989), .A2(n14990), .ZN(n14991) );
  NOR2_X1 U18099 ( .A1(n14983), .A2(n14991), .ZN(n16313) );
  NAND2_X1 U18100 ( .A1(n16313), .A2(n15012), .ZN(n14996) );
  OR2_X1 U18101 ( .A1(n14992), .A2(n14993), .ZN(n14994) );
  AND2_X1 U18102 ( .A1(n9742), .A2(n14994), .ZN(n18996) );
  NAND2_X1 U18103 ( .A1(n18996), .A2(n14998), .ZN(n14995) );
  OAI211_X1 U18104 ( .C1(n14998), .C2(n14997), .A(n14996), .B(n14995), .ZN(
        P2_U2867) );
  AND2_X1 U18105 ( .A1(n14999), .A2(n15009), .ZN(n15010) );
  OAI21_X1 U18106 ( .B1(n15010), .B2(n15000), .A(n14989), .ZN(n15092) );
  NOR2_X1 U18107 ( .A1(n15008), .A2(n15001), .ZN(n15002) );
  OR2_X1 U18108 ( .A1(n14992), .A2(n15002), .ZN(n19008) );
  NOR2_X1 U18109 ( .A1(n19008), .A2(n15004), .ZN(n15003) );
  AOI21_X1 U18110 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15004), .A(n15003), .ZN(
        n15005) );
  OAI21_X1 U18111 ( .B1(n15092), .B2(n15025), .A(n15005), .ZN(P2_U2868) );
  AND2_X1 U18112 ( .A1(n15022), .A2(n15006), .ZN(n15007) );
  NOR2_X1 U18113 ( .A1(n15008), .A2(n15007), .ZN(n19019) );
  INV_X1 U18114 ( .A(n19019), .ZN(n15016) );
  INV_X1 U18115 ( .A(n15009), .ZN(n15011) );
  INV_X1 U18116 ( .A(n14999), .ZN(n15017) );
  AOI21_X1 U18117 ( .B1(n15011), .B2(n15017), .A(n15010), .ZN(n16319) );
  NAND2_X1 U18118 ( .A1(n16319), .A2(n15012), .ZN(n15014) );
  NAND2_X1 U18119 ( .A1(n15015), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15013) );
  OAI211_X1 U18120 ( .C1(n15016), .C2(n15015), .A(n15014), .B(n15013), .ZN(
        P2_U2869) );
  OAI21_X1 U18121 ( .B1(n13765), .B2(n15018), .A(n15017), .ZN(n15102) );
  NAND2_X1 U18122 ( .A1(n15020), .A2(n15019), .ZN(n15021) );
  NAND2_X1 U18123 ( .A1(n15022), .A2(n15021), .ZN(n15467) );
  NOR2_X1 U18124 ( .A1(n15467), .A2(n15004), .ZN(n15023) );
  AOI21_X1 U18125 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15004), .A(n15023), .ZN(
        n15024) );
  OAI21_X1 U18126 ( .B1(n15102), .B2(n15025), .A(n15024), .ZN(P2_U2870) );
  NAND3_X1 U18127 ( .A1(n15027), .A2(n19269), .A3(n15026), .ZN(n15032) );
  INV_X1 U18128 ( .A(n19207), .ZN(n15041) );
  INV_X1 U18129 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19285) );
  OAI22_X1 U18130 ( .A1(n15041), .A2(n19222), .B1(n19239), .B2(n19285), .ZN(
        n15030) );
  INV_X1 U18131 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n15028) );
  NOR2_X1 U18132 ( .A1(n15042), .A2(n15028), .ZN(n15029) );
  AOI211_X1 U18133 ( .C1(BUF1_REG_29__SCAN_IN), .C2(n19208), .A(n15030), .B(
        n15029), .ZN(n15031) );
  OAI211_X1 U18134 ( .C1(n19215), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        P2_U2890) );
  INV_X1 U18135 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n15035) );
  AOI22_X1 U18136 ( .A1(n19207), .A2(n19224), .B1(n19264), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15034) );
  OAI21_X1 U18137 ( .B1(n15042), .B2(n15035), .A(n15034), .ZN(n15037) );
  NOR2_X1 U18138 ( .A1(n15322), .A2(n19215), .ZN(n15036) );
  AOI211_X1 U18139 ( .C1(n19208), .C2(BUF1_REG_28__SCAN_IN), .A(n15037), .B(
        n15036), .ZN(n15038) );
  OAI21_X1 U18140 ( .B1(n15039), .B2(n19216), .A(n15038), .ZN(P2_U2891) );
  INV_X1 U18141 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19289) );
  OAI22_X1 U18142 ( .A1(n15041), .A2(n19227), .B1(n19239), .B2(n19289), .ZN(
        n15044) );
  NOR2_X1 U18143 ( .A1(n15042), .A2(n17338), .ZN(n15043) );
  AOI211_X1 U18144 ( .C1(BUF1_REG_27__SCAN_IN), .C2(n19208), .A(n15044), .B(
        n15043), .ZN(n15045) );
  NAND2_X1 U18145 ( .A1(n15046), .A2(n19269), .ZN(n15052) );
  AOI22_X1 U18146 ( .A1(n19207), .A2(n19229), .B1(n19264), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15051) );
  AOI21_X1 U18147 ( .B1(n10173), .B2(n10174), .A(n12606), .ZN(n16297) );
  AOI22_X1 U18148 ( .A1(n16297), .A2(n19265), .B1(n19208), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15050) );
  NAND2_X1 U18149 ( .A1(n19209), .A2(BUF2_REG_26__SCAN_IN), .ZN(n15049) );
  NAND4_X1 U18150 ( .A1(n15052), .A2(n15051), .A3(n15050), .A4(n15049), .ZN(
        P2_U2893) );
  INV_X1 U18151 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19293) );
  NAND2_X1 U18152 ( .A1(n19207), .A2(n15053), .ZN(n15054) );
  OAI21_X1 U18153 ( .B1(n19239), .B2(n19293), .A(n15054), .ZN(n15055) );
  AOI21_X1 U18154 ( .B1(n15358), .B2(n19265), .A(n15055), .ZN(n15057) );
  AOI22_X1 U18155 ( .A1(n19208), .A2(BUF1_REG_25__SCAN_IN), .B1(n19209), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15056) );
  OAI211_X1 U18156 ( .C1(n15058), .C2(n19216), .A(n15057), .B(n15056), .ZN(
        P2_U2894) );
  OR2_X1 U18157 ( .A1(n15059), .A2(n19216), .ZN(n15066) );
  AOI22_X1 U18158 ( .A1(n19207), .A2(n19234), .B1(n19264), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n15065) );
  AOI22_X1 U18159 ( .A1(n19208), .A2(BUF1_REG_24__SCAN_IN), .B1(n19209), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15064) );
  NAND2_X1 U18160 ( .A1(n9718), .A2(n15060), .ZN(n15061) );
  AND2_X1 U18161 ( .A1(n15062), .A2(n15061), .ZN(n16299) );
  NAND2_X1 U18162 ( .A1(n16299), .A2(n19265), .ZN(n15063) );
  NAND4_X1 U18163 ( .A1(n15066), .A2(n15065), .A3(n15064), .A4(n15063), .ZN(
        P2_U2895) );
  AOI22_X1 U18164 ( .A1(n19208), .A2(BUF1_REG_23__SCAN_IN), .B1(n19209), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U18165 ( .A1(n19207), .A2(n15067), .B1(n19264), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15068) );
  OAI211_X1 U18166 ( .C1(n15383), .C2(n19215), .A(n15069), .B(n15068), .ZN(
        n15070) );
  AOI21_X1 U18167 ( .B1(n15071), .B2(n19269), .A(n15070), .ZN(n15072) );
  INV_X1 U18168 ( .A(n15072), .ZN(P2_U2896) );
  AOI22_X1 U18169 ( .A1(n19208), .A2(BUF1_REG_22__SCAN_IN), .B1(n19209), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n15075) );
  AOI22_X1 U18170 ( .A1(n19207), .A2(n15073), .B1(n19264), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15074) );
  OAI211_X1 U18171 ( .C1(n19215), .C2(n15395), .A(n15075), .B(n15074), .ZN(
        n15076) );
  AOI21_X1 U18172 ( .B1(n15077), .B2(n19269), .A(n15076), .ZN(n15078) );
  INV_X1 U18173 ( .A(n15078), .ZN(P2_U2897) );
  XNOR2_X1 U18174 ( .A(n15422), .B(n9776), .ZN(n15407) );
  INV_X1 U18175 ( .A(n15407), .ZN(n18978) );
  AOI22_X1 U18176 ( .A1(n19208), .A2(BUF1_REG_21__SCAN_IN), .B1(n19209), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15080) );
  AOI22_X1 U18177 ( .A1(n19207), .A2(n19407), .B1(n19264), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15079) );
  OAI211_X1 U18178 ( .C1(n18978), .C2(n19215), .A(n15080), .B(n15079), .ZN(
        n15081) );
  INV_X1 U18179 ( .A(n15081), .ZN(n15082) );
  OAI21_X1 U18180 ( .B1(n15083), .B2(n19216), .A(n15082), .ZN(P2_U2898) );
  OR2_X1 U18181 ( .A1(n15445), .A2(n15085), .ZN(n15086) );
  NAND2_X1 U18182 ( .A1(n15084), .A2(n15086), .ZN(n19007) );
  AOI22_X1 U18183 ( .A1(n19208), .A2(BUF1_REG_19__SCAN_IN), .B1(n19209), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n15089) );
  AOI22_X1 U18184 ( .A1(n19207), .A2(n15087), .B1(n19264), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15088) );
  OAI211_X1 U18185 ( .C1(n19215), .C2(n19007), .A(n15089), .B(n15088), .ZN(
        n15090) );
  INV_X1 U18186 ( .A(n15090), .ZN(n15091) );
  OAI21_X1 U18187 ( .B1(n15092), .B2(n19216), .A(n15091), .ZN(P2_U2900) );
  AND2_X1 U18188 ( .A1(n15094), .A2(n15093), .ZN(n15096) );
  OR2_X1 U18189 ( .A1(n15096), .A2(n15095), .ZN(n19035) );
  AOI22_X1 U18190 ( .A1(n19208), .A2(BUF1_REG_17__SCAN_IN), .B1(n19209), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n15099) );
  AOI22_X1 U18191 ( .A1(n19207), .A2(n15097), .B1(n19264), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15098) );
  OAI211_X1 U18192 ( .C1(n19215), .C2(n19035), .A(n15099), .B(n15098), .ZN(
        n15100) );
  INV_X1 U18193 ( .A(n15100), .ZN(n15101) );
  OAI21_X1 U18194 ( .B1(n15102), .B2(n19216), .A(n15101), .ZN(P2_U2902) );
  XNOR2_X1 U18195 ( .A(n15103), .B(n15323), .ZN(n15345) );
  AOI21_X1 U18196 ( .B1(n15323), .B2(n15104), .A(n12566), .ZN(n15343) );
  NAND2_X1 U18197 ( .A1(n19038), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15335) );
  OAI21_X1 U18198 ( .B1(n16359), .B2(n15105), .A(n15335), .ZN(n15106) );
  AOI21_X1 U18199 ( .B1(n16351), .B2(n15107), .A(n15106), .ZN(n15108) );
  OAI21_X1 U18200 ( .B1(n15340), .B2(n19376), .A(n15108), .ZN(n15109) );
  AOI21_X1 U18201 ( .B1(n15343), .B2(n19352), .A(n15109), .ZN(n15110) );
  OAI21_X1 U18202 ( .B1(n15345), .B2(n16324), .A(n15110), .ZN(P2_U2987) );
  OAI21_X1 U18203 ( .B1(n15111), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15104), .ZN(n15355) );
  INV_X1 U18204 ( .A(n15120), .ZN(n15112) );
  OAI21_X1 U18205 ( .B1(n15123), .B2(n15112), .A(n15121), .ZN(n15114) );
  XNOR2_X1 U18206 ( .A(n15114), .B(n15113), .ZN(n15352) );
  NOR2_X1 U18207 ( .A1(n16294), .A2(n19376), .ZN(n15118) );
  NAND2_X1 U18208 ( .A1(n19038), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15347) );
  NAND2_X1 U18209 ( .A1(n19349), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15115) );
  OAI211_X1 U18210 ( .C1(n19359), .C2(n15116), .A(n15347), .B(n15115), .ZN(
        n15117) );
  AOI211_X1 U18211 ( .C1(n15352), .C2(n19355), .A(n15118), .B(n15117), .ZN(
        n15119) );
  OAI21_X1 U18212 ( .B1(n15355), .B2(n16325), .A(n15119), .ZN(P2_U2988) );
  NAND2_X1 U18213 ( .A1(n15121), .A2(n15120), .ZN(n15122) );
  XNOR2_X1 U18214 ( .A(n15123), .B(n15122), .ZN(n15369) );
  INV_X1 U18215 ( .A(n15111), .ZN(n15357) );
  NAND2_X1 U18216 ( .A1(n15124), .A2(n15365), .ZN(n15356) );
  NAND3_X1 U18217 ( .A1(n15357), .A2(n19352), .A3(n15356), .ZN(n15130) );
  NAND2_X1 U18218 ( .A1(n19038), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15360) );
  OAI21_X1 U18219 ( .B1(n16359), .B2(n15125), .A(n15360), .ZN(n15127) );
  NOR2_X1 U18220 ( .A1(n15362), .A2(n19376), .ZN(n15126) );
  AOI211_X1 U18221 ( .C1(n16351), .C2(n15128), .A(n15127), .B(n15126), .ZN(
        n15129) );
  OAI211_X1 U18222 ( .C1(n16324), .C2(n15369), .A(n15130), .B(n15129), .ZN(
        P2_U2989) );
  INV_X1 U18223 ( .A(n15131), .ZN(n15132) );
  OAI21_X1 U18224 ( .B1(n15132), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15124), .ZN(n15379) );
  NAND2_X1 U18225 ( .A1(n9748), .A2(n15133), .ZN(n15134) );
  XNOR2_X1 U18226 ( .A(n15135), .B(n15134), .ZN(n15377) );
  NOR2_X1 U18227 ( .A1(n19129), .A2(n19983), .ZN(n15373) );
  NOR2_X1 U18228 ( .A1(n19359), .A2(n15136), .ZN(n15137) );
  AOI211_X1 U18229 ( .C1(n19349), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15373), .B(n15137), .ZN(n15138) );
  OAI21_X1 U18230 ( .B1(n16301), .B2(n19376), .A(n15138), .ZN(n15139) );
  AOI21_X1 U18231 ( .B1(n15377), .B2(n19355), .A(n15139), .ZN(n15140) );
  OAI21_X1 U18232 ( .B1(n15379), .B2(n16325), .A(n15140), .ZN(P2_U2990) );
  OAI21_X1 U18233 ( .B1(n15141), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15131), .ZN(n15380) );
  INV_X1 U18234 ( .A(n15142), .ZN(n15385) );
  NAND2_X1 U18235 ( .A1(n16351), .A2(n15143), .ZN(n15144) );
  NAND2_X1 U18236 ( .A1(n19038), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15381) );
  OAI211_X1 U18237 ( .C1(n16359), .C2(n15145), .A(n15144), .B(n15381), .ZN(
        n15150) );
  NOR2_X1 U18238 ( .A1(n15147), .A2(n15146), .ZN(n15386) );
  INV_X1 U18239 ( .A(n15148), .ZN(n15387) );
  NOR3_X1 U18240 ( .A1(n15386), .A2(n15387), .A3(n16324), .ZN(n15149) );
  AOI211_X1 U18241 ( .C1(n19351), .C2(n15385), .A(n15150), .B(n15149), .ZN(
        n15151) );
  OAI21_X1 U18242 ( .B1(n15380), .B2(n16325), .A(n15151), .ZN(P2_U2991) );
  OAI21_X1 U18243 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n9670), .A(
        n10199), .ZN(n15405) );
  NAND2_X1 U18244 ( .A1(n15153), .A2(n15152), .ZN(n15154) );
  XNOR2_X1 U18245 ( .A(n15155), .B(n15154), .ZN(n15403) );
  NOR2_X1 U18246 ( .A1(n19129), .A2(n19979), .ZN(n15397) );
  NOR2_X1 U18247 ( .A1(n19359), .A2(n15156), .ZN(n15157) );
  AOI211_X1 U18248 ( .C1(n19349), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15397), .B(n15157), .ZN(n15158) );
  OAI21_X1 U18249 ( .B1(n15401), .B2(n19376), .A(n15158), .ZN(n15159) );
  AOI21_X1 U18250 ( .B1(n15403), .B2(n19355), .A(n15159), .ZN(n15160) );
  OAI21_X1 U18251 ( .B1(n15405), .B2(n16325), .A(n15160), .ZN(P2_U2992) );
  INV_X1 U18252 ( .A(n15161), .ZN(n15256) );
  INV_X1 U18253 ( .A(n15253), .ZN(n15162) );
  INV_X1 U18254 ( .A(n15241), .ZN(n15163) );
  INV_X1 U18255 ( .A(n15233), .ZN(n15164) );
  INV_X1 U18256 ( .A(n15165), .ZN(n15223) );
  NAND3_X1 U18257 ( .A1(n15214), .A2(n15215), .A3(n15167), .ZN(n15213) );
  INV_X1 U18258 ( .A(n15168), .ZN(n15171) );
  INV_X1 U18259 ( .A(n15169), .ZN(n15170) );
  INV_X1 U18260 ( .A(n15174), .ZN(n15173) );
  NOR2_X1 U18261 ( .A1(n15187), .A2(n15174), .ZN(n15178) );
  NAND2_X1 U18262 ( .A1(n15176), .A2(n15175), .ZN(n15177) );
  XNOR2_X1 U18263 ( .A(n15178), .B(n15177), .ZN(n15418) );
  AOI21_X1 U18265 ( .B1(n15409), .B2(n15180), .A(n9670), .ZN(n15415) );
  AND2_X1 U18266 ( .A1(n19038), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15406) );
  AOI21_X1 U18267 ( .B1(n19349), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15406), .ZN(n15182) );
  NAND2_X1 U18268 ( .A1(n16351), .A2(n18983), .ZN(n15181) );
  OAI211_X1 U18269 ( .C1(n18979), .C2(n19376), .A(n15182), .B(n15181), .ZN(
        n15183) );
  AOI21_X1 U18270 ( .B1(n15415), .B2(n19352), .A(n15183), .ZN(n15184) );
  OAI21_X1 U18271 ( .B1(n15418), .B2(n16324), .A(n15184), .ZN(P2_U2993) );
  OAI21_X1 U18272 ( .B1(n15185), .B2(n15432), .A(n15425), .ZN(n15186) );
  NAND2_X1 U18273 ( .A1(n15186), .A2(n15180), .ZN(n15431) );
  NAND2_X1 U18274 ( .A1(n15419), .A2(n19355), .ZN(n15192) );
  NOR2_X1 U18275 ( .A1(n19129), .A2(n15188), .ZN(n15423) );
  AOI21_X1 U18276 ( .B1(n19349), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15423), .ZN(n15189) );
  OAI21_X1 U18277 ( .B1(n19359), .B2(n18991), .A(n15189), .ZN(n15190) );
  AOI21_X1 U18278 ( .B1(n18996), .B2(n19351), .A(n15190), .ZN(n15191) );
  OAI211_X1 U18279 ( .C1(n16325), .C2(n15431), .A(n15192), .B(n15191), .ZN(
        P2_U2994) );
  OAI21_X1 U18280 ( .B1(n15212), .B2(n15202), .A(n15201), .ZN(n15195) );
  XNOR2_X1 U18281 ( .A(n15193), .B(n15432), .ZN(n15194) );
  XNOR2_X1 U18282 ( .A(n15195), .B(n15194), .ZN(n15442) );
  XNOR2_X1 U18283 ( .A(n15185), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15440) );
  NAND2_X1 U18284 ( .A1(n19038), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15433) );
  OAI21_X1 U18285 ( .B1(n16359), .B2(n15196), .A(n15433), .ZN(n15197) );
  AOI21_X1 U18286 ( .B1(n16351), .B2(n19003), .A(n15197), .ZN(n15198) );
  OAI21_X1 U18287 ( .B1(n19008), .B2(n19376), .A(n15198), .ZN(n15199) );
  AOI21_X1 U18288 ( .B1(n15440), .B2(n19352), .A(n15199), .ZN(n15200) );
  OAI21_X1 U18289 ( .B1(n15442), .B2(n16324), .A(n15200), .ZN(P2_U2995) );
  INV_X1 U18290 ( .A(n15201), .ZN(n15203) );
  NOR2_X1 U18291 ( .A1(n15203), .A2(n15202), .ZN(n15204) );
  XNOR2_X1 U18292 ( .A(n15212), .B(n15204), .ZN(n15457) );
  NAND2_X1 U18293 ( .A1(n19038), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15446) );
  NAND2_X1 U18294 ( .A1(n19349), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15205) );
  OAI211_X1 U18295 ( .C1(n19359), .C2(n19014), .A(n15446), .B(n15205), .ZN(
        n15210) );
  NAND2_X1 U18296 ( .A1(n15206), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15207) );
  NAND2_X1 U18297 ( .A1(n15207), .A2(n15451), .ZN(n15208) );
  NAND2_X1 U18298 ( .A1(n15208), .A2(n15185), .ZN(n15454) );
  NOR2_X1 U18299 ( .A1(n15454), .A2(n16325), .ZN(n15209) );
  AOI211_X1 U18300 ( .C1(n19351), .C2(n19019), .A(n15210), .B(n15209), .ZN(
        n15211) );
  OAI21_X1 U18301 ( .B1(n15457), .B2(n16324), .A(n15211), .ZN(P2_U2996) );
  INV_X1 U18302 ( .A(n15212), .ZN(n15216) );
  AOI22_X1 U18303 ( .A1(n15216), .A2(n15215), .B1(n15214), .B2(n15213), .ZN(
        n15465) );
  XNOR2_X1 U18304 ( .A(n15206), .B(n15217), .ZN(n15221) );
  NAND2_X1 U18305 ( .A1(n19038), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15468) );
  OAI21_X1 U18306 ( .B1(n16359), .B2(n10239), .A(n15468), .ZN(n15218) );
  AOI21_X1 U18307 ( .B1(n16351), .B2(n19028), .A(n15218), .ZN(n15219) );
  OAI21_X1 U18308 ( .B1(n15467), .B2(n19376), .A(n15219), .ZN(n15220) );
  AOI21_X1 U18309 ( .B1(n15221), .B2(n19352), .A(n15220), .ZN(n15222) );
  OAI21_X1 U18310 ( .B1(n15465), .B2(n16324), .A(n15222), .ZN(P2_U2997) );
  XNOR2_X1 U18311 ( .A(n15224), .B(n15223), .ZN(n15487) );
  NOR2_X1 U18312 ( .A1(n19129), .A2(n19970), .ZN(n15480) );
  AOI21_X1 U18313 ( .B1(n19349), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15480), .ZN(n15225) );
  OAI21_X1 U18314 ( .B1(n19359), .B2(n15226), .A(n15225), .ZN(n15231) );
  INV_X1 U18315 ( .A(n15227), .ZN(n15228) );
  AOI21_X1 U18316 ( .B1(n15228), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15229) );
  NOR3_X1 U18317 ( .A1(n15229), .A2(n15206), .A3(n16325), .ZN(n15230) );
  AOI211_X1 U18318 ( .C1(n19351), .C2(n15477), .A(n15231), .B(n15230), .ZN(
        n15232) );
  OAI21_X1 U18319 ( .B1(n16324), .B2(n15487), .A(n15232), .ZN(P2_U2998) );
  XNOR2_X1 U18320 ( .A(n15227), .B(n15460), .ZN(n15501) );
  NAND2_X1 U18321 ( .A1(n15234), .A2(n15233), .ZN(n15235) );
  XNOR2_X1 U18322 ( .A(n15236), .B(n15235), .ZN(n15499) );
  NAND2_X1 U18323 ( .A1(n19038), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15491) );
  OAI21_X1 U18324 ( .B1(n16359), .B2(n19036), .A(n15491), .ZN(n15237) );
  AOI21_X1 U18325 ( .B1(n16351), .B2(n19044), .A(n15237), .ZN(n15238) );
  OAI21_X1 U18326 ( .B1(n15488), .B2(n19376), .A(n15238), .ZN(n15239) );
  AOI21_X1 U18327 ( .B1(n15499), .B2(n19355), .A(n15239), .ZN(n15240) );
  OAI21_X1 U18328 ( .B1(n16325), .B2(n15501), .A(n15240), .ZN(P2_U2999) );
  NAND2_X1 U18329 ( .A1(n15242), .A2(n15241), .ZN(n15243) );
  XNOR2_X1 U18330 ( .A(n15244), .B(n15243), .ZN(n15518) );
  NAND2_X1 U18331 ( .A1(n15245), .A2(n15507), .ZN(n15246) );
  AND2_X1 U18332 ( .A1(n15227), .A2(n15246), .ZN(n15516) );
  NAND2_X1 U18333 ( .A1(n19058), .A2(n19351), .ZN(n15248) );
  AOI22_X1 U18334 ( .A1(n19349), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19038), .ZN(n15247) );
  OAI211_X1 U18335 ( .C1(n19359), .C2(n19051), .A(n15248), .B(n15247), .ZN(
        n15249) );
  AOI21_X1 U18336 ( .B1(n15516), .B2(n19352), .A(n15249), .ZN(n15250) );
  OAI21_X1 U18337 ( .B1(n15518), .B2(n16324), .A(n15250), .ZN(P2_U3000) );
  NAND2_X1 U18338 ( .A1(n15285), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15270) );
  OAI21_X1 U18339 ( .B1(n15270), .B2(n15521), .A(n15527), .ZN(n15252) );
  NAND2_X1 U18340 ( .A1(n15252), .A2(n15245), .ZN(n15532) );
  NAND2_X1 U18341 ( .A1(n15254), .A2(n15253), .ZN(n15255) );
  XNOR2_X1 U18342 ( .A(n15256), .B(n15255), .ZN(n15530) );
  NAND2_X1 U18343 ( .A1(n19038), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15520) );
  OAI21_X1 U18344 ( .B1(n16359), .B2(n15257), .A(n15520), .ZN(n15258) );
  AOI21_X1 U18345 ( .B1(n16351), .B2(n19064), .A(n15258), .ZN(n15259) );
  OAI21_X1 U18346 ( .B1(n19376), .B2(n19069), .A(n15259), .ZN(n15260) );
  AOI21_X1 U18347 ( .B1(n15530), .B2(n19355), .A(n15260), .ZN(n15261) );
  OAI21_X1 U18348 ( .B1(n15532), .B2(n16325), .A(n15261), .ZN(P2_U3001) );
  XNOR2_X1 U18349 ( .A(n15270), .B(n15521), .ZN(n15545) );
  INV_X1 U18350 ( .A(n15262), .ZN(n15264) );
  NAND2_X1 U18351 ( .A1(n15264), .A2(n15263), .ZN(n15265) );
  NOR2_X1 U18352 ( .A1(n19129), .A2(n19964), .ZN(n15538) );
  NOR2_X1 U18353 ( .A1(n19359), .A2(n19079), .ZN(n15266) );
  AOI211_X1 U18354 ( .C1(n19349), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15538), .B(n15266), .ZN(n15267) );
  OAI21_X1 U18355 ( .B1(n19376), .B2(n15537), .A(n15267), .ZN(n15268) );
  AOI21_X1 U18356 ( .B1(n15543), .B2(n19355), .A(n15268), .ZN(n15269) );
  OAI21_X1 U18357 ( .B1(n15545), .B2(n16325), .A(n15269), .ZN(P2_U3002) );
  OAI21_X1 U18358 ( .B1(n15285), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15270), .ZN(n15564) );
  INV_X1 U18359 ( .A(n15271), .ZN(n15272) );
  NAND2_X1 U18360 ( .A1(n15273), .A2(n15272), .ZN(n15277) );
  NOR2_X1 U18361 ( .A1(n15275), .A2(n15274), .ZN(n15276) );
  XNOR2_X1 U18362 ( .A(n15277), .B(n15276), .ZN(n15559) );
  INV_X1 U18363 ( .A(n15559), .ZN(n15282) );
  NOR2_X1 U18364 ( .A1(n19129), .A2(n15278), .ZN(n15554) );
  NOR2_X1 U18365 ( .A1(n16359), .A2(n19087), .ZN(n15279) );
  AOI211_X1 U18366 ( .C1(n19090), .C2(n16351), .A(n15554), .B(n15279), .ZN(
        n15280) );
  OAI21_X1 U18367 ( .B1(n19376), .B2(n15558), .A(n15280), .ZN(n15281) );
  AOI21_X1 U18368 ( .B1(n15282), .B2(n19355), .A(n15281), .ZN(n15283) );
  OAI21_X1 U18369 ( .B1(n15564), .B2(n16325), .A(n15283), .ZN(P2_U3003) );
  AOI21_X1 U18370 ( .B1(n15251), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15284) );
  NAND2_X1 U18371 ( .A1(n15287), .A2(n15286), .ZN(n15596) );
  INV_X1 U18372 ( .A(n15594), .ZN(n15288) );
  OAI21_X1 U18373 ( .B1(n15596), .B2(n15288), .A(n15593), .ZN(n15292) );
  NAND2_X1 U18374 ( .A1(n15290), .A2(n15289), .ZN(n15291) );
  XNOR2_X1 U18375 ( .A(n15292), .B(n15291), .ZN(n15577) );
  NOR2_X1 U18376 ( .A1(n19129), .A2(n19961), .ZN(n15570) );
  NOR2_X1 U18377 ( .A1(n19359), .A2(n19102), .ZN(n15293) );
  AOI211_X1 U18378 ( .C1(n19349), .C2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15570), .B(n15293), .ZN(n15294) );
  OAI21_X1 U18379 ( .B1(n19376), .B2(n19103), .A(n15294), .ZN(n15295) );
  AOI21_X1 U18380 ( .B1(n15577), .B2(n19355), .A(n15295), .ZN(n15296) );
  OAI21_X1 U18381 ( .B1(n15579), .B2(n16325), .A(n15296), .ZN(P2_U3004) );
  XNOR2_X1 U18382 ( .A(n15298), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15299) );
  XNOR2_X1 U18383 ( .A(n15297), .B(n15299), .ZN(n16380) );
  NAND2_X1 U18384 ( .A1(n16333), .A2(n16332), .ZN(n15301) );
  XOR2_X1 U18385 ( .A(n15301), .B(n15300), .Z(n16377) );
  OAI22_X1 U18386 ( .A1(n16359), .A2(n15302), .B1(n20984), .B2(n19129), .ZN(
        n15303) );
  AOI21_X1 U18387 ( .B1(n16351), .B2(n19120), .A(n15303), .ZN(n15304) );
  OAI21_X1 U18388 ( .B1(n19376), .B2(n19124), .A(n15304), .ZN(n15305) );
  AOI21_X1 U18389 ( .B1(n16377), .B2(n19355), .A(n15305), .ZN(n15306) );
  OAI21_X1 U18390 ( .B1(n16380), .B2(n16325), .A(n15306), .ZN(P2_U3007) );
  OAI21_X1 U18391 ( .B1(n15308), .B2(n16371), .A(n15307), .ZN(n15309) );
  INV_X1 U18392 ( .A(n15309), .ZN(n15311) );
  INV_X1 U18393 ( .A(n15313), .ZN(n15314) );
  OAI21_X1 U18394 ( .B1(n15315), .B2(n15589), .A(n15314), .ZN(n15316) );
  OAI21_X1 U18395 ( .B1(n15319), .B2(n19366), .A(n15318), .ZN(P2_U3016) );
  INV_X1 U18396 ( .A(n15320), .ZN(n15332) );
  OAI21_X1 U18397 ( .B1(n15322), .B2(n16371), .A(n15321), .ZN(n15326) );
  NOR3_X1 U18398 ( .A1(n15324), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15323), .ZN(n15325) );
  AOI211_X1 U18399 ( .C1(n15327), .C2(n19369), .A(n15326), .B(n15325), .ZN(
        n15328) );
  OAI21_X1 U18400 ( .B1(n15330), .B2(n15329), .A(n15328), .ZN(n15331) );
  OAI21_X1 U18401 ( .B1(n15334), .B2(n15597), .A(n15333), .ZN(P2_U3018) );
  OAI21_X1 U18402 ( .B1(n15336), .B2(n16371), .A(n15335), .ZN(n15337) );
  AOI21_X1 U18403 ( .B1(n15338), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15337), .ZN(n15339) );
  OAI21_X1 U18404 ( .B1(n15340), .B2(n15589), .A(n15339), .ZN(n15341) );
  AOI211_X1 U18405 ( .C1(n15343), .C2(n16361), .A(n15342), .B(n15341), .ZN(
        n15344) );
  OAI21_X1 U18406 ( .B1(n15345), .B2(n15597), .A(n15344), .ZN(P2_U3019) );
  XNOR2_X1 U18407 ( .A(n15348), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15351) );
  NAND2_X1 U18408 ( .A1(n16297), .A2(n19364), .ZN(n15346) );
  OAI211_X1 U18409 ( .C1(n15361), .C2(n15348), .A(n15347), .B(n15346), .ZN(
        n15350) );
  NOR2_X1 U18410 ( .A1(n16294), .A2(n15589), .ZN(n15349) );
  AOI211_X1 U18411 ( .C1(n15351), .C2(n15366), .A(n15350), .B(n15349), .ZN(
        n15354) );
  NAND2_X1 U18412 ( .A1(n15352), .A2(n19361), .ZN(n15353) );
  OAI211_X1 U18413 ( .C1(n15355), .C2(n19366), .A(n15354), .B(n15353), .ZN(
        P2_U3020) );
  NAND3_X1 U18414 ( .A1(n15357), .A2(n16361), .A3(n15356), .ZN(n15368) );
  NAND2_X1 U18415 ( .A1(n15358), .A2(n19364), .ZN(n15359) );
  OAI211_X1 U18416 ( .C1(n15361), .C2(n15365), .A(n15360), .B(n15359), .ZN(
        n15364) );
  NOR2_X1 U18417 ( .A1(n15362), .A2(n15589), .ZN(n15363) );
  AOI211_X1 U18418 ( .C1(n15366), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        n15367) );
  OAI211_X1 U18419 ( .C1(n15369), .C2(n15597), .A(n15368), .B(n15367), .ZN(
        P2_U3021) );
  AND2_X1 U18420 ( .A1(n15394), .A2(n15370), .ZN(n15372) );
  OAI21_X1 U18421 ( .B1(n15372), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15371), .ZN(n15375) );
  AOI21_X1 U18422 ( .B1(n16299), .B2(n19364), .A(n15373), .ZN(n15374) );
  OAI211_X1 U18423 ( .C1(n16301), .C2(n15589), .A(n15375), .B(n15374), .ZN(
        n15376) );
  AOI21_X1 U18424 ( .B1(n15377), .B2(n19361), .A(n15376), .ZN(n15378) );
  OAI21_X1 U18425 ( .B1(n15379), .B2(n19366), .A(n15378), .ZN(P2_U3022) );
  OR2_X1 U18426 ( .A1(n15380), .A2(n19366), .ZN(n15392) );
  NAND2_X1 U18427 ( .A1(n15398), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15382) );
  OAI211_X1 U18428 ( .C1(n16371), .C2(n15383), .A(n15382), .B(n15381), .ZN(
        n15384) );
  AOI21_X1 U18429 ( .B1(n15385), .B2(n19369), .A(n15384), .ZN(n15391) );
  OR3_X1 U18430 ( .A1(n15387), .A2(n15386), .A3(n15597), .ZN(n15390) );
  OAI211_X1 U18431 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15394), .B(n15388), .ZN(
        n15389) );
  NAND4_X1 U18432 ( .A1(n15392), .A2(n15391), .A3(n15390), .A4(n15389), .ZN(
        P2_U3023) );
  NAND2_X1 U18433 ( .A1(n15394), .A2(n15393), .ZN(n15400) );
  NOR2_X1 U18434 ( .A1(n15395), .A2(n16371), .ZN(n15396) );
  AOI211_X1 U18435 ( .C1(n15398), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15397), .B(n15396), .ZN(n15399) );
  OAI211_X1 U18436 ( .C1(n15401), .C2(n15589), .A(n15400), .B(n15399), .ZN(
        n15402) );
  AOI21_X1 U18437 ( .B1(n15403), .B2(n19361), .A(n15402), .ZN(n15404) );
  OAI21_X1 U18438 ( .B1(n15405), .B2(n19366), .A(n15404), .ZN(P2_U3024) );
  INV_X1 U18439 ( .A(n18979), .ZN(n15414) );
  AOI21_X1 U18440 ( .B1(n19364), .B2(n15407), .A(n15406), .ZN(n15408) );
  OAI21_X1 U18441 ( .B1(n15410), .B2(n15409), .A(n15408), .ZN(n15413) );
  NOR3_X1 U18442 ( .A1(n15438), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15411), .ZN(n15412) );
  AOI211_X1 U18443 ( .C1(n15414), .C2(n19369), .A(n15413), .B(n15412), .ZN(
        n15417) );
  NAND2_X1 U18444 ( .A1(n15415), .A2(n16361), .ZN(n15416) );
  OAI211_X1 U18445 ( .C1(n15418), .C2(n15597), .A(n15417), .B(n15416), .ZN(
        P2_U3025) );
  NAND2_X1 U18446 ( .A1(n15419), .A2(n19361), .ZN(n15430) );
  NAND2_X1 U18447 ( .A1(n15084), .A2(n15420), .ZN(n15421) );
  AND2_X1 U18448 ( .A1(n15422), .A2(n15421), .ZN(n18995) );
  AOI21_X1 U18449 ( .B1(n19364), .B2(n18995), .A(n15423), .ZN(n15424) );
  OAI21_X1 U18450 ( .B1(n15447), .B2(n15425), .A(n15424), .ZN(n15428) );
  XNOR2_X1 U18451 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15426) );
  NOR2_X1 U18452 ( .A1(n15438), .A2(n15426), .ZN(n15427) );
  AOI211_X1 U18453 ( .C1(n18996), .C2(n19369), .A(n15428), .B(n15427), .ZN(
        n15429) );
  OAI211_X1 U18454 ( .C1(n15431), .C2(n19366), .A(n15430), .B(n15429), .ZN(
        P2_U3026) );
  INV_X1 U18455 ( .A(n19008), .ZN(n15436) );
  NOR2_X1 U18456 ( .A1(n15447), .A2(n15432), .ZN(n15435) );
  OAI21_X1 U18457 ( .B1(n16371), .B2(n19007), .A(n15433), .ZN(n15434) );
  AOI211_X1 U18458 ( .C1(n15436), .C2(n19369), .A(n15435), .B(n15434), .ZN(
        n15437) );
  OAI21_X1 U18459 ( .B1(n15438), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15437), .ZN(n15439) );
  AOI21_X1 U18460 ( .B1(n15440), .B2(n16361), .A(n15439), .ZN(n15441) );
  OAI21_X1 U18461 ( .B1(n15442), .B2(n15597), .A(n15441), .ZN(P2_U3027) );
  NOR2_X1 U18462 ( .A1(n15095), .A2(n15443), .ZN(n15444) );
  OR2_X1 U18463 ( .A1(n15445), .A2(n15444), .ZN(n16318) );
  OAI21_X1 U18464 ( .B1(n16371), .B2(n16318), .A(n15446), .ZN(n15449) );
  NOR2_X1 U18465 ( .A1(n15447), .A2(n15451), .ZN(n15448) );
  AOI211_X1 U18466 ( .C1(n19019), .C2(n19369), .A(n15449), .B(n15448), .ZN(
        n15453) );
  NOR2_X1 U18467 ( .A1(n15497), .A2(n15450), .ZN(n15466) );
  NAND3_X1 U18468 ( .A1(n15466), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15451), .ZN(n15452) );
  OAI211_X1 U18469 ( .C1(n15454), .C2(n19366), .A(n15453), .B(n15452), .ZN(
        n15455) );
  INV_X1 U18470 ( .A(n15455), .ZN(n15456) );
  OAI21_X1 U18471 ( .B1(n15457), .B2(n15597), .A(n15456), .ZN(P2_U3028) );
  AND2_X1 U18472 ( .A1(n19366), .A2(n15458), .ZN(n15459) );
  OR2_X1 U18473 ( .A1(n15206), .A2(n15459), .ZN(n15464) );
  NAND2_X1 U18474 ( .A1(n15461), .A2(n15460), .ZN(n15462) );
  AND2_X1 U18475 ( .A1(n15493), .A2(n15462), .ZN(n15463) );
  AND2_X1 U18476 ( .A1(n15464), .A2(n15463), .ZN(n15476) );
  OAI21_X1 U18477 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15613), .A(
        n15476), .ZN(n15474) );
  NOR2_X1 U18478 ( .A1(n15465), .A2(n15597), .ZN(n15473) );
  AOI21_X1 U18479 ( .B1(n15206), .B2(n16361), .A(n15466), .ZN(n15471) );
  INV_X1 U18480 ( .A(n15467), .ZN(n19030) );
  OAI21_X1 U18481 ( .B1(n16371), .B2(n19035), .A(n15468), .ZN(n15469) );
  AOI21_X1 U18482 ( .B1(n19030), .B2(n19369), .A(n15469), .ZN(n15470) );
  OAI21_X1 U18483 ( .B1(n15471), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15470), .ZN(n15472) );
  AOI211_X1 U18484 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n15474), .A(
        n15473), .B(n15472), .ZN(n15475) );
  INV_X1 U18485 ( .A(n15475), .ZN(P2_U3029) );
  INV_X1 U18486 ( .A(n15476), .ZN(n15485) );
  INV_X1 U18487 ( .A(n15477), .ZN(n15483) );
  OAI21_X1 U18488 ( .B1(n15227), .B2(n19366), .A(n15497), .ZN(n15479) );
  NAND3_X1 U18489 ( .A1(n15479), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n15478), .ZN(n15482) );
  AOI21_X1 U18490 ( .B1(n19364), .B2(n19210), .A(n15480), .ZN(n15481) );
  OAI211_X1 U18491 ( .C1(n15483), .C2(n15589), .A(n15482), .B(n15481), .ZN(
        n15484) );
  AOI21_X1 U18492 ( .B1(n15485), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15484), .ZN(n15486) );
  OAI21_X1 U18493 ( .B1(n15487), .B2(n15597), .A(n15486), .ZN(P2_U3030) );
  INV_X1 U18494 ( .A(n15488), .ZN(n19045) );
  OR2_X1 U18495 ( .A1(n9749), .A2(n15489), .ZN(n15490) );
  NAND2_X1 U18496 ( .A1(n14920), .A2(n15490), .ZN(n19218) );
  OAI21_X1 U18497 ( .B1(n16371), .B2(n19218), .A(n15491), .ZN(n15492) );
  AOI21_X1 U18498 ( .B1(n19045), .B2(n19369), .A(n15492), .ZN(n15496) );
  INV_X1 U18499 ( .A(n15493), .ZN(n15494) );
  NAND2_X1 U18500 ( .A1(n15494), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15495) );
  OAI211_X1 U18501 ( .C1(n15497), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15496), .B(n15495), .ZN(n15498) );
  AOI21_X1 U18502 ( .B1(n15499), .B2(n19361), .A(n15498), .ZN(n15500) );
  OAI21_X1 U18503 ( .B1(n19366), .B2(n15501), .A(n15500), .ZN(P2_U3031) );
  INV_X1 U18504 ( .A(n15503), .ZN(n15502) );
  NAND2_X1 U18505 ( .A1(n15592), .A2(n15502), .ZN(n15505) );
  NOR2_X1 U18506 ( .A1(n15505), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15542) );
  AND2_X1 U18507 ( .A1(n19370), .A2(n15503), .ZN(n15504) );
  OR2_X1 U18508 ( .A1(n15580), .A2(n15504), .ZN(n15536) );
  NOR2_X1 U18509 ( .A1(n15542), .A2(n15536), .ZN(n15528) );
  OR2_X1 U18510 ( .A1(n15505), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15522) );
  NAND2_X1 U18511 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19348), .ZN(n15506) );
  OAI221_X1 U18512 ( .B1(n15507), .B2(n15528), .C1(n15507), .C2(n15522), .A(
        n15506), .ZN(n15515) );
  NAND3_X1 U18513 ( .A1(n15592), .A2(n15508), .A3(n15507), .ZN(n15513) );
  NOR2_X1 U18514 ( .A1(n15510), .A2(n15509), .ZN(n15511) );
  OR2_X1 U18515 ( .A1(n9749), .A2(n15511), .ZN(n19221) );
  INV_X1 U18516 ( .A(n19221), .ZN(n19057) );
  AOI22_X1 U18517 ( .A1(n19058), .A2(n19369), .B1(n19364), .B2(n19057), .ZN(
        n15512) );
  NAND2_X1 U18518 ( .A1(n15513), .A2(n15512), .ZN(n15514) );
  AOI211_X1 U18519 ( .C1(n15516), .C2(n16361), .A(n15515), .B(n15514), .ZN(
        n15517) );
  OAI21_X1 U18520 ( .B1(n15597), .B2(n15518), .A(n15517), .ZN(P2_U3032) );
  XNOR2_X1 U18521 ( .A(n15533), .B(n15519), .ZN(n19223) );
  INV_X1 U18522 ( .A(n19223), .ZN(n15525) );
  OAI21_X1 U18523 ( .B1(n19069), .B2(n15589), .A(n15520), .ZN(n15524) );
  NOR2_X1 U18524 ( .A1(n15522), .A2(n15521), .ZN(n15523) );
  AOI211_X1 U18525 ( .C1(n19364), .C2(n15525), .A(n15524), .B(n15523), .ZN(
        n15526) );
  OAI21_X1 U18526 ( .B1(n15528), .B2(n15527), .A(n15526), .ZN(n15529) );
  AOI21_X1 U18527 ( .B1(n15530), .B2(n19361), .A(n15529), .ZN(n15531) );
  OAI21_X1 U18528 ( .B1(n15532), .B2(n19366), .A(n15531), .ZN(P2_U3033) );
  INV_X1 U18529 ( .A(n15533), .ZN(n15534) );
  OAI21_X1 U18530 ( .B1(n15550), .B2(n15535), .A(n15534), .ZN(n19226) );
  NAND2_X1 U18531 ( .A1(n15536), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15540) );
  INV_X1 U18532 ( .A(n15537), .ZN(n19081) );
  AOI21_X1 U18533 ( .B1(n19081), .B2(n19369), .A(n15538), .ZN(n15539) );
  OAI211_X1 U18534 ( .C1(n16371), .C2(n19226), .A(n15540), .B(n15539), .ZN(
        n15541) );
  AOI211_X1 U18535 ( .C1(n15543), .C2(n19361), .A(n15542), .B(n15541), .ZN(
        n15544) );
  OAI21_X1 U18536 ( .B1(n15545), .B2(n19366), .A(n15544), .ZN(P2_U3034) );
  INV_X1 U18537 ( .A(n15565), .ZN(n15547) );
  NOR2_X1 U18538 ( .A1(n15580), .A2(n15591), .ZN(n15575) );
  NAND3_X1 U18539 ( .A1(n15592), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n15546), .ZN(n15573) );
  OAI21_X1 U18540 ( .B1(n15547), .B2(n15575), .A(n15573), .ZN(n15562) );
  INV_X1 U18541 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15548) );
  NAND3_X1 U18542 ( .A1(n15592), .A2(n15549), .A3(n15548), .ZN(n15557) );
  INV_X1 U18543 ( .A(n15550), .ZN(n15553) );
  NAND2_X1 U18544 ( .A1(n15568), .A2(n15551), .ZN(n15552) );
  NAND2_X1 U18545 ( .A1(n15553), .A2(n15552), .ZN(n19228) );
  INV_X1 U18546 ( .A(n19228), .ZN(n15555) );
  AOI21_X1 U18547 ( .B1(n19364), .B2(n15555), .A(n15554), .ZN(n15556) );
  OAI211_X1 U18548 ( .C1(n15558), .C2(n15589), .A(n15557), .B(n15556), .ZN(
        n15561) );
  NOR2_X1 U18549 ( .A1(n15559), .A2(n15597), .ZN(n15560) );
  AOI211_X1 U18550 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15562), .A(
        n15561), .B(n15560), .ZN(n15563) );
  OAI21_X1 U18551 ( .B1(n15564), .B2(n19366), .A(n15563), .ZN(P2_U3035) );
  NAND2_X1 U18552 ( .A1(n15565), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15574) );
  INV_X1 U18553 ( .A(n19103), .ZN(n15571) );
  NAND2_X1 U18554 ( .A1(n15584), .A2(n15566), .ZN(n15567) );
  NAND2_X1 U18555 ( .A1(n15568), .A2(n15567), .ZN(n19231) );
  NOR2_X1 U18556 ( .A1(n16371), .A2(n19231), .ZN(n15569) );
  AOI211_X1 U18557 ( .C1(n15571), .C2(n19369), .A(n15570), .B(n15569), .ZN(
        n15572) );
  OAI211_X1 U18558 ( .C1(n15575), .C2(n15574), .A(n15573), .B(n15572), .ZN(
        n15576) );
  AOI21_X1 U18559 ( .B1(n15577), .B2(n19361), .A(n15576), .ZN(n15578) );
  OAI21_X1 U18560 ( .B1(n15579), .B2(n19366), .A(n15578), .ZN(P2_U3036) );
  XNOR2_X1 U18561 ( .A(n15251), .B(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16326) );
  NAND2_X1 U18562 ( .A1(n15580), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15588) );
  NAND2_X1 U18563 ( .A1(n15582), .A2(n15581), .ZN(n15583) );
  NAND2_X1 U18564 ( .A1(n15584), .A2(n15583), .ZN(n19233) );
  INV_X1 U18565 ( .A(n19233), .ZN(n15586) );
  NOR2_X1 U18566 ( .A1(n10748), .A2(n19129), .ZN(n15585) );
  AOI21_X1 U18567 ( .B1(n19364), .B2(n15586), .A(n15585), .ZN(n15587) );
  OAI211_X1 U18568 ( .C1(n15589), .C2(n19114), .A(n15588), .B(n15587), .ZN(
        n15590) );
  AOI21_X1 U18569 ( .B1(n15592), .B2(n15591), .A(n15590), .ZN(n15599) );
  NAND2_X1 U18570 ( .A1(n15594), .A2(n15593), .ZN(n15595) );
  XNOR2_X1 U18571 ( .A(n15596), .B(n15595), .ZN(n16323) );
  OR2_X1 U18572 ( .A1(n16323), .A2(n15597), .ZN(n15598) );
  OAI211_X1 U18573 ( .C1(n16326), .C2(n19366), .A(n15599), .B(n15598), .ZN(
        P2_U3037) );
  OAI21_X1 U18574 ( .B1(n15601), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15602), .ZN(n16346) );
  XOR2_X1 U18575 ( .A(n9750), .B(n15603), .Z(n16348) );
  NAND2_X1 U18576 ( .A1(n15605), .A2(n15604), .ZN(n15616) );
  NOR2_X1 U18577 ( .A1(n10493), .A2(n19129), .ZN(n15609) );
  XOR2_X1 U18578 ( .A(n15607), .B(n15606), .Z(n19240) );
  NOR2_X1 U18579 ( .A1(n16371), .A2(n19240), .ZN(n15608) );
  AOI211_X1 U18580 ( .C1(n19137), .C2(n19369), .A(n15609), .B(n15608), .ZN(
        n15615) );
  INV_X1 U18581 ( .A(n15610), .ZN(n15612) );
  OAI21_X1 U18582 ( .B1(n15613), .B2(n15612), .A(n15611), .ZN(n16373) );
  NAND2_X1 U18583 ( .A1(n16373), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15614) );
  OAI211_X1 U18584 ( .C1(n15617), .C2(n15616), .A(n15615), .B(n15614), .ZN(
        n15618) );
  AOI21_X1 U18585 ( .B1(n16348), .B2(n19361), .A(n15618), .ZN(n15619) );
  OAI21_X1 U18586 ( .B1(n19366), .B2(n16346), .A(n15619), .ZN(P2_U3040) );
  INV_X1 U18587 ( .A(n12726), .ZN(n15626) );
  INV_X1 U18588 ( .A(n13058), .ZN(n15622) );
  MUX2_X1 U18589 ( .A(n15622), .B(n15621), .S(n15620), .Z(n15623) );
  OAI21_X1 U18590 ( .B1(n15624), .B2(n15635), .A(n15623), .ZN(n16404) );
  AOI22_X1 U18591 ( .A1(n15626), .A2(n16421), .B1(n16404), .B2(n15625), .ZN(
        n15627) );
  OAI21_X1 U18592 ( .B1(n15628), .B2(n16424), .A(n15627), .ZN(n15629) );
  MUX2_X1 U18593 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15629), .S(
        n15644), .Z(P2_U3601) );
  INV_X1 U18594 ( .A(n20019), .ZN(n19243) );
  NAND2_X1 U18595 ( .A1(n9664), .A2(n15630), .ZN(n15639) );
  INV_X1 U18596 ( .A(n15631), .ZN(n15634) );
  OAI22_X1 U18597 ( .A1(n15634), .A2(n15639), .B1(n15632), .B2(n15633), .ZN(
        n15638) );
  NOR2_X1 U18598 ( .A1(n15636), .A2(n15635), .ZN(n15637) );
  AOI211_X1 U18599 ( .C1(n15640), .C2(n15639), .A(n15638), .B(n15637), .ZN(
        n16382) );
  OAI22_X1 U18600 ( .A1(n16382), .A2(n20008), .B1(n15642), .B2(n15641), .ZN(
        n15643) );
  AOI21_X1 U18601 ( .B1(n16421), .B2(n19243), .A(n15643), .ZN(n15645) );
  MUX2_X1 U18602 ( .A(n9640), .B(n15645), .S(n15644), .Z(n15647) );
  INV_X1 U18603 ( .A(n15647), .ZN(P2_U3599) );
  AOI22_X1 U18604 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15652) );
  AOI22_X1 U18605 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15651) );
  AOI22_X1 U18606 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9648), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15650) );
  AOI22_X1 U18607 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15649) );
  NAND4_X1 U18608 ( .A1(n15652), .A2(n15651), .A3(n15650), .A4(n15649), .ZN(
        n15658) );
  AOI22_X1 U18609 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9645), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U18610 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15655) );
  AOI22_X1 U18611 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15654) );
  AOI22_X1 U18612 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15653) );
  NAND4_X1 U18613 ( .A1(n15656), .A2(n15655), .A3(n15654), .A4(n15653), .ZN(
        n15657) );
  NOR2_X1 U18614 ( .A1(n15658), .A2(n15657), .ZN(n17066) );
  AOI22_X1 U18615 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15662) );
  AOI22_X1 U18616 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9657), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15661) );
  AOI22_X1 U18617 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15660) );
  AOI22_X1 U18618 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15659) );
  NAND4_X1 U18619 ( .A1(n15662), .A2(n15661), .A3(n15660), .A4(n15659), .ZN(
        n15668) );
  AOI22_X1 U18620 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15666) );
  AOI22_X1 U18621 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15665) );
  AOI22_X1 U18622 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15664) );
  AOI22_X1 U18623 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15663) );
  NAND4_X1 U18624 ( .A1(n15666), .A2(n15665), .A3(n15664), .A4(n15663), .ZN(
        n15667) );
  NOR2_X1 U18625 ( .A1(n15668), .A2(n15667), .ZN(n17077) );
  AOI22_X1 U18626 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9649), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15673) );
  AOI22_X1 U18627 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15672) );
  AOI22_X1 U18628 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15671) );
  AOI22_X1 U18629 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15670) );
  NAND4_X1 U18630 ( .A1(n15673), .A2(n15672), .A3(n15671), .A4(n15670), .ZN(
        n15679) );
  AOI22_X1 U18631 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15677) );
  AOI22_X1 U18632 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15676) );
  AOI22_X1 U18633 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15675) );
  AOI22_X1 U18634 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15674) );
  NAND4_X1 U18635 ( .A1(n15677), .A2(n15676), .A3(n15675), .A4(n15674), .ZN(
        n15678) );
  NOR2_X1 U18636 ( .A1(n15679), .A2(n15678), .ZN(n17088) );
  AOI22_X1 U18637 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15683) );
  AOI22_X1 U18638 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15682) );
  AOI22_X1 U18639 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15681) );
  AOI22_X1 U18640 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15680) );
  NAND4_X1 U18641 ( .A1(n15683), .A2(n15682), .A3(n15681), .A4(n15680), .ZN(
        n15689) );
  AOI22_X1 U18642 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15687) );
  AOI22_X1 U18643 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9644), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15686) );
  AOI22_X1 U18644 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15685) );
  AOI22_X1 U18645 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15684) );
  NAND4_X1 U18646 ( .A1(n15687), .A2(n15686), .A3(n15685), .A4(n15684), .ZN(
        n15688) );
  NOR2_X1 U18647 ( .A1(n15689), .A2(n15688), .ZN(n17089) );
  NOR2_X1 U18648 ( .A1(n17088), .A2(n17089), .ZN(n17087) );
  AOI22_X1 U18649 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n9642), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15699) );
  AOI22_X1 U18650 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9645), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15698) );
  INV_X1 U18651 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17306) );
  AOI22_X1 U18652 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9650), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15690) );
  OAI21_X1 U18653 ( .B1(n9706), .B2(n17306), .A(n15690), .ZN(n15696) );
  AOI22_X1 U18654 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17269), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17252), .ZN(n15694) );
  AOI22_X1 U18655 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9648), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15693) );
  AOI22_X1 U18656 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17270), .ZN(n15692) );
  AOI22_X1 U18657 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15691) );
  NAND4_X1 U18658 ( .A1(n15694), .A2(n15693), .A3(n15692), .A4(n15691), .ZN(
        n15695) );
  AOI211_X1 U18659 ( .C1(n15834), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n15696), .B(n15695), .ZN(n15697) );
  NAND3_X1 U18660 ( .A1(n15699), .A2(n15698), .A3(n15697), .ZN(n17083) );
  NAND2_X1 U18661 ( .A1(n17087), .A2(n17083), .ZN(n17082) );
  NOR2_X1 U18662 ( .A1(n17077), .A2(n17082), .ZN(n17076) );
  AOI22_X1 U18663 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15710) );
  AOI22_X1 U18664 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15709) );
  AOI22_X1 U18665 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15700) );
  OAI21_X1 U18666 ( .B1(n15701), .B2(n21083), .A(n15700), .ZN(n15707) );
  AOI22_X1 U18667 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15705) );
  AOI22_X1 U18668 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15704) );
  AOI22_X1 U18669 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15703) );
  AOI22_X1 U18670 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15702) );
  NAND4_X1 U18671 ( .A1(n15705), .A2(n15704), .A3(n15703), .A4(n15702), .ZN(
        n15706) );
  AOI211_X1 U18672 ( .C1(n9649), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n15707), .B(n15706), .ZN(n15708) );
  NAND3_X1 U18673 ( .A1(n15710), .A2(n15709), .A3(n15708), .ZN(n17072) );
  NAND2_X1 U18674 ( .A1(n17076), .A2(n17072), .ZN(n17071) );
  NOR2_X1 U18675 ( .A1(n17066), .A2(n17071), .ZN(n17065) );
  AOI22_X1 U18676 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9650), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15720) );
  AOI22_X1 U18677 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15719) );
  AOI22_X1 U18678 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15711) );
  OAI21_X1 U18679 ( .B1(n15648), .B2(n15816), .A(n15711), .ZN(n15717) );
  AOI22_X1 U18680 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15715) );
  AOI22_X1 U18681 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15714) );
  AOI22_X1 U18682 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15713) );
  AOI22_X1 U18683 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15712) );
  NAND4_X1 U18684 ( .A1(n15715), .A2(n15714), .A3(n15713), .A4(n15712), .ZN(
        n15716) );
  AOI211_X1 U18685 ( .C1(n9657), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n15717), .B(n15716), .ZN(n15718) );
  NAND3_X1 U18686 ( .A1(n15720), .A2(n15719), .A3(n15718), .ZN(n15721) );
  NAND2_X1 U18687 ( .A1(n17065), .A2(n15721), .ZN(n17059) );
  OAI21_X1 U18688 ( .B1(n17065), .B2(n15721), .A(n17059), .ZN(n17333) );
  NAND2_X1 U18689 ( .A1(n18307), .A2(n17314), .ZN(n17308) );
  INV_X1 U18690 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16783) );
  NAND2_X1 U18691 ( .A1(n18307), .A2(n17147), .ZN(n17129) );
  NAND2_X1 U18692 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17117), .ZN(n17104) );
  NAND2_X1 U18693 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17086), .ZN(n17081) );
  NAND2_X1 U18694 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17080), .ZN(n17070) );
  NAND2_X1 U18695 ( .A1(n17305), .A2(n17070), .ZN(n17068) );
  OAI21_X1 U18696 ( .B1(n15722), .B2(n17308), .A(n17068), .ZN(n17061) );
  INV_X1 U18697 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17069) );
  NOR3_X1 U18698 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17069), .A3(n17070), .ZN(
        n15723) );
  AOI21_X1 U18699 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17061), .A(n15723), .ZN(
        n15724) );
  OAI21_X1 U18700 ( .B1(n17333), .B2(n17305), .A(n15724), .ZN(P3_U2675) );
  AOI22_X1 U18701 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15728) );
  AOI22_X1 U18702 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15727) );
  AOI22_X1 U18703 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9657), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15726) );
  AOI22_X1 U18704 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15725) );
  NAND4_X1 U18705 ( .A1(n15728), .A2(n15727), .A3(n15726), .A4(n15725), .ZN(
        n15734) );
  AOI22_X1 U18706 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15732) );
  AOI22_X1 U18707 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15731) );
  AOI22_X1 U18708 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15730) );
  AOI22_X1 U18709 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15729) );
  NAND4_X1 U18710 ( .A1(n15732), .A2(n15731), .A3(n15730), .A4(n15729), .ZN(
        n15733) );
  NOR2_X1 U18711 ( .A1(n15734), .A2(n15733), .ZN(n17410) );
  NAND2_X1 U18712 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17245), .ZN(n17244) );
  NOR2_X1 U18713 ( .A1(n17404), .A2(n17244), .ZN(n17232) );
  AOI21_X1 U18714 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17232), .A(n17311), .ZN(
        n17231) );
  AND2_X1 U18715 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17232), .ZN(n15735) );
  INV_X1 U18716 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17215) );
  AOI22_X1 U18717 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17231), .B1(n15735), 
        .B2(n17215), .ZN(n15736) );
  OAI21_X1 U18718 ( .B1(n17410), .B2(n17305), .A(n15736), .ZN(P3_U2690) );
  NAND2_X1 U18719 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18490) );
  INV_X1 U18720 ( .A(n17897), .ZN(n18783) );
  NOR2_X1 U18721 ( .A1(n16434), .A2(n18783), .ZN(n15738) );
  AOI221_X1 U18722 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18490), .C1(n15738), 
        .C2(n18490), .A(n15737), .ZN(n18266) );
  NOR2_X1 U18723 ( .A1(n15739), .A2(n18539), .ZN(n15740) );
  OAI21_X1 U18724 ( .B1(n15740), .B2(n18330), .A(n18267), .ZN(n18264) );
  AOI22_X1 U18725 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18266), .B1(
        n18264), .B2(n18263), .ZN(P3_U2865) );
  INV_X1 U18726 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21110) );
  INV_X1 U18727 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18073) );
  INV_X1 U18728 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18056) );
  NOR2_X1 U18729 ( .A1(n18073), .A2(n18056), .ZN(n18047) );
  INV_X1 U18730 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17714) );
  INV_X1 U18731 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18021) );
  NAND2_X1 U18732 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17680) );
  NOR3_X1 U18733 ( .A1(n17714), .A2(n18021), .A3(n17680), .ZN(n15916) );
  AND2_X1 U18734 ( .A1(n18047), .A2(n15916), .ZN(n18004) );
  NAND2_X1 U18735 ( .A1(n18004), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17944) );
  INV_X1 U18736 ( .A(n17944), .ZN(n15926) );
  INV_X1 U18737 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18106) );
  INV_X1 U18738 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18149) );
  INV_X1 U18739 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18145) );
  NOR2_X1 U18740 ( .A1(n18149), .A2(n18145), .ZN(n18131) );
  NAND2_X1 U18741 ( .A1(n18131), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18134) );
  INV_X1 U18742 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17805) );
  NOR2_X1 U18743 ( .A1(n18134), .A2(n17805), .ZN(n18094) );
  NAND2_X1 U18744 ( .A1(n18094), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17773) );
  NOR2_X1 U18745 ( .A1(n18106), .A2(n17773), .ZN(n18067) );
  NAND2_X1 U18746 ( .A1(n18067), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17736) );
  INV_X1 U18747 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18192) );
  INV_X1 U18748 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18209) );
  INV_X1 U18749 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18212) );
  NOR3_X1 U18750 ( .A1(n18192), .A2(n18209), .A3(n18212), .ZN(n18187) );
  AOI21_X1 U18751 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18229) );
  INV_X1 U18752 ( .A(n18229), .ZN(n15742) );
  NAND2_X1 U18753 ( .A1(n18187), .A2(n15742), .ZN(n18159) );
  NAND3_X1 U18754 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15748) );
  NOR2_X1 U18755 ( .A1(n18159), .A2(n15748), .ZN(n18063) );
  NAND2_X1 U18756 ( .A1(n18043), .A2(n18063), .ZN(n18045) );
  NAND2_X1 U18757 ( .A1(n18929), .A2(n15743), .ZN(n15745) );
  OAI21_X1 U18758 ( .B1(n15746), .B2(n15745), .A(n15744), .ZN(n18724) );
  AOI21_X2 U18759 ( .B1(n18725), .B2(n18729), .A(n18724), .ZN(n18745) );
  AOI21_X1 U18760 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18065), .A(
        n18749), .ZN(n18225) );
  NAND3_X1 U18761 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18187), .ZN(n18158) );
  NOR2_X1 U18762 ( .A1(n15748), .A2(n18158), .ZN(n18093) );
  NAND2_X1 U18763 ( .A1(n18043), .A2(n18093), .ZN(n15925) );
  OAI22_X1 U18764 ( .A1(n18742), .A2(n18045), .B1(n18225), .B2(n15925), .ZN(
        n16496) );
  NAND2_X1 U18765 ( .A1(n15926), .A2(n16496), .ZN(n17967) );
  INV_X1 U18766 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17961) );
  NAND3_X1 U18767 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17614) );
  NOR2_X1 U18768 ( .A1(n17961), .A2(n17614), .ZN(n16459) );
  NAND2_X1 U18769 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16459), .ZN(
        n15749) );
  NOR3_X1 U18770 ( .A1(n21110), .A2(n17967), .A3(n15749), .ZN(n16482) );
  INV_X1 U18771 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17948) );
  AOI22_X1 U18772 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15753) );
  AOI22_X1 U18773 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15752) );
  AOI22_X1 U18774 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15751) );
  AOI22_X1 U18775 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15750) );
  NAND4_X1 U18776 ( .A1(n15753), .A2(n15752), .A3(n15751), .A4(n15750), .ZN(
        n15759) );
  AOI22_X1 U18777 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9649), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15757) );
  AOI22_X1 U18778 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15756) );
  AOI22_X1 U18779 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15755) );
  AOI22_X1 U18780 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15754) );
  NAND4_X1 U18781 ( .A1(n15757), .A2(n15756), .A3(n15755), .A4(n15754), .ZN(
        n15758) );
  AOI22_X1 U18782 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15763) );
  AOI22_X1 U18783 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15762) );
  AOI22_X1 U18784 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15761) );
  AOI22_X1 U18785 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15760) );
  NAND4_X1 U18786 ( .A1(n15763), .A2(n15762), .A3(n15761), .A4(n15760), .ZN(
        n15770) );
  AOI22_X1 U18787 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15768) );
  AOI22_X1 U18788 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15767) );
  AOI22_X1 U18789 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15766) );
  AOI22_X1 U18790 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9657), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15765) );
  NAND4_X1 U18791 ( .A1(n15768), .A2(n15767), .A3(n15766), .A4(n15765), .ZN(
        n15769) );
  AOI22_X1 U18792 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15774) );
  AOI22_X1 U18793 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15773) );
  AOI22_X1 U18794 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15772) );
  AOI22_X1 U18795 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15771) );
  NAND4_X1 U18796 ( .A1(n15774), .A2(n15773), .A3(n15772), .A4(n15771), .ZN(
        n15780) );
  AOI22_X1 U18797 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15778) );
  AOI22_X1 U18798 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15777) );
  AOI22_X1 U18799 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15776) );
  AOI22_X1 U18800 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15775) );
  NAND4_X1 U18801 ( .A1(n15778), .A2(n15777), .A3(n15776), .A4(n15775), .ZN(
        n15779) );
  AOI22_X1 U18802 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15791) );
  AOI22_X1 U18803 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15790) );
  INV_X1 U18804 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15782) );
  AOI22_X1 U18805 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15781) );
  OAI21_X1 U18806 ( .B1(n15827), .B2(n15782), .A(n15781), .ZN(n15788) );
  AOI22_X1 U18807 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15786) );
  AOI22_X1 U18808 ( .A1(n15669), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15785) );
  AOI22_X1 U18809 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15784) );
  AOI22_X1 U18810 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15783) );
  NAND4_X1 U18811 ( .A1(n15786), .A2(n15785), .A3(n15784), .A4(n15783), .ZN(
        n15787) );
  AOI211_X1 U18812 ( .C1(n9645), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n15788), .B(n15787), .ZN(n15789) );
  AOI22_X1 U18813 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9649), .B1(n9644), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15794) );
  AOI22_X1 U18814 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17263), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n15814), .ZN(n15793) );
  AOI22_X1 U18815 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n15795), .ZN(n15800) );
  AOI22_X1 U18816 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n15796), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n15804), .ZN(n15799) );
  AOI22_X1 U18817 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n9648), .ZN(n15798) );
  AOI22_X1 U18818 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17270), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17264), .ZN(n15797) );
  AOI22_X1 U18819 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17035), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17269), .ZN(n15801) );
  NAND2_X1 U18820 ( .A1(n17459), .A2(n15840), .ZN(n15839) );
  AOI22_X1 U18821 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15813) );
  AOI22_X1 U18822 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15812) );
  AOI22_X1 U18823 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15802) );
  OAI21_X1 U18824 ( .B1(n15803), .B2(n21083), .A(n15802), .ZN(n15810) );
  AOI22_X1 U18825 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15808) );
  AOI22_X1 U18826 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15807) );
  AOI22_X1 U18827 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15806) );
  AOI22_X1 U18828 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15805) );
  NAND4_X1 U18829 ( .A1(n15808), .A2(n15807), .A3(n15806), .A4(n15805), .ZN(
        n15809) );
  AOI211_X1 U18830 ( .C1(n9650), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n15810), .B(n15809), .ZN(n15811) );
  NAND3_X1 U18831 ( .A1(n15813), .A2(n15812), .A3(n15811), .ZN(n15869) );
  NAND2_X1 U18832 ( .A1(n15839), .A2(n15869), .ZN(n15848) );
  NOR2_X1 U18833 ( .A1(n17450), .A2(n15848), .ZN(n15838) );
  AOI22_X1 U18834 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15825) );
  AOI22_X1 U18835 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15824) );
  AOI22_X1 U18836 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15815) );
  OAI21_X1 U18837 ( .B1(n10212), .B2(n15816), .A(n15815), .ZN(n15822) );
  AOI22_X1 U18838 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9644), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15820) );
  AOI22_X1 U18839 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15819) );
  AOI22_X1 U18840 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15818) );
  AOI22_X1 U18841 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15817) );
  NAND4_X1 U18842 ( .A1(n15820), .A2(n15819), .A3(n15818), .A4(n15817), .ZN(
        n15821) );
  AOI211_X1 U18843 ( .C1(n17035), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n15822), .B(n15821), .ZN(n15823) );
  NAND3_X1 U18844 ( .A1(n15825), .A2(n15824), .A3(n15823), .ZN(n15867) );
  NAND2_X1 U18845 ( .A1(n15838), .A2(n15867), .ZN(n15852) );
  NOR2_X1 U18846 ( .A1(n17444), .A2(n15852), .ZN(n15856) );
  AOI22_X1 U18847 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15837) );
  AOI22_X1 U18848 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15836) );
  AOI22_X1 U18849 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15826) );
  OAI21_X1 U18850 ( .B1(n15827), .B2(n17280), .A(n15826), .ZN(n15833) );
  AOI22_X1 U18851 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15831) );
  AOI22_X1 U18852 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9645), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15830) );
  AOI22_X1 U18853 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15829) );
  AOI22_X1 U18854 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15828) );
  NAND4_X1 U18855 ( .A1(n15831), .A2(n15830), .A3(n15829), .A4(n15828), .ZN(
        n15832) );
  AOI211_X1 U18856 ( .C1(n15834), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n15833), .B(n15832), .ZN(n15835) );
  NAND2_X1 U18857 ( .A1(n15856), .A2(n16498), .ZN(n15857) );
  XOR2_X1 U18858 ( .A(n15838), .B(n15867), .Z(n15850) );
  XNOR2_X1 U18859 ( .A(n15839), .B(n15869), .ZN(n15845) );
  NOR2_X1 U18860 ( .A1(n15845), .A2(n18212), .ZN(n15846) );
  INV_X1 U18861 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18222) );
  NOR2_X1 U18862 ( .A1(n15843), .A2(n18222), .ZN(n15844) );
  INV_X1 U18863 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18886) );
  NOR2_X1 U18864 ( .A1(n15870), .A2(n18886), .ZN(n15842) );
  NAND3_X1 U18865 ( .A1(n17937), .A2(n15870), .A3(n18886), .ZN(n15841) );
  OAI221_X1 U18866 ( .B1(n15842), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n17937), .C2(n15870), .A(n15841), .ZN(n17919) );
  NOR2_X1 U18867 ( .A1(n17919), .A2(n17918), .ZN(n17917) );
  NOR2_X1 U18868 ( .A1(n15844), .A2(n17917), .ZN(n17908) );
  XOR2_X1 U18869 ( .A(n15845), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n17907) );
  NOR2_X1 U18870 ( .A1(n17908), .A2(n17907), .ZN(n17906) );
  NOR2_X1 U18871 ( .A1(n15847), .A2(n18209), .ZN(n15849) );
  XNOR2_X1 U18872 ( .A(n15848), .B(n17450), .ZN(n17895) );
  XOR2_X1 U18873 ( .A(n18192), .B(n15850), .Z(n17885) );
  XNOR2_X1 U18874 ( .A(n15852), .B(n17444), .ZN(n15854) );
  NOR2_X1 U18875 ( .A1(n15853), .A2(n15854), .ZN(n15855) );
  INV_X1 U18876 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18186) );
  INV_X1 U18877 ( .A(n16498), .ZN(n17441) );
  XOR2_X1 U18878 ( .A(n15856), .B(n17441), .Z(n15859) );
  NAND2_X1 U18879 ( .A1(n15858), .A2(n15859), .ZN(n17864) );
  NAND2_X1 U18880 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17864), .ZN(
        n15861) );
  NOR2_X1 U18881 ( .A1(n15857), .A2(n15861), .ZN(n15863) );
  INV_X1 U18882 ( .A(n15857), .ZN(n15862) );
  OR2_X1 U18883 ( .A1(n15859), .A2(n15858), .ZN(n17865) );
  OAI21_X1 U18884 ( .B1(n15862), .B2(n15861), .A(n17865), .ZN(n15860) );
  INV_X1 U18885 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18162) );
  INV_X1 U18886 ( .A(n18067), .ZN(n18082) );
  INV_X1 U18887 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17987) );
  NOR2_X1 U18888 ( .A1(n17987), .A2(n17944), .ZN(n15912) );
  INV_X1 U18889 ( .A(n15912), .ZN(n17641) );
  NAND3_X1 U18890 ( .A1(n17951), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16502) );
  NOR2_X1 U18891 ( .A1(n18281), .A2(n15864), .ZN(n15896) );
  NAND2_X1 U18892 ( .A1(n15896), .A2(n17317), .ZN(n15901) );
  NAND2_X1 U18893 ( .A1(n16499), .A2(n17441), .ZN(n18166) );
  INV_X1 U18894 ( .A(n15867), .ZN(n17447) );
  INV_X1 U18895 ( .A(n17450), .ZN(n15879) );
  NAND2_X1 U18896 ( .A1(n15878), .A2(n15879), .ZN(n15866) );
  OAI21_X1 U18897 ( .B1(n16498), .B2(n16495), .A(n17849), .ZN(n15890) );
  INV_X1 U18898 ( .A(n15890), .ZN(n15889) );
  XNOR2_X1 U18899 ( .A(n15867), .B(n15866), .ZN(n15882) );
  XNOR2_X1 U18900 ( .A(n15869), .B(n15868), .ZN(n15874) );
  OR2_X1 U18901 ( .A1(n18222), .A2(n15872), .ZN(n15873) );
  NAND2_X1 U18902 ( .A1(n15870), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15871) );
  XNOR2_X1 U18903 ( .A(n15872), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17922) );
  NAND2_X1 U18904 ( .A1(n17921), .A2(n17922), .ZN(n17920) );
  NAND2_X1 U18905 ( .A1(n15874), .A2(n15876), .ZN(n15877) );
  XOR2_X1 U18906 ( .A(n15879), .B(n15878), .Z(n15880) );
  XOR2_X1 U18907 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15880), .Z(
        n17900) );
  NAND2_X1 U18908 ( .A1(n17899), .A2(n17900), .ZN(n17898) );
  NAND2_X1 U18909 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15880), .ZN(
        n15881) );
  NAND2_X1 U18910 ( .A1(n15882), .A2(n15884), .ZN(n15885) );
  XOR2_X1 U18911 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15887), .Z(
        n17872) );
  NAND2_X1 U18912 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15887), .ZN(
        n15888) );
  NAND2_X1 U18913 ( .A1(n17870), .A2(n15888), .ZN(n15891) );
  NAND2_X1 U18914 ( .A1(n15889), .A2(n15891), .ZN(n15892) );
  XNOR2_X1 U18915 ( .A(n15891), .B(n15890), .ZN(n17859) );
  NAND2_X1 U18916 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17859), .ZN(
        n17858) );
  NAND2_X1 U18917 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17981), .ZN(
        n17631) );
  NOR2_X1 U18918 ( .A1(n17948), .A2(n17631), .ZN(n17630) );
  NAND2_X1 U18919 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17630), .ZN(
        n15923) );
  INV_X1 U18920 ( .A(n15923), .ZN(n17950) );
  NAND3_X1 U18921 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n17950), .ZN(n16501) );
  OAI22_X1 U18922 ( .A1(n17985), .A2(n16502), .B1(n18166), .B2(n16501), .ZN(
        n15904) );
  AOI21_X1 U18923 ( .B1(n15894), .B2(n15893), .A(n9891), .ZN(n18714) );
  INV_X1 U18924 ( .A(n18714), .ZN(n15902) );
  OAI21_X1 U18925 ( .B1(n18285), .B2(n18929), .A(n16635), .ZN(n15895) );
  OAI21_X1 U18926 ( .B1(n15896), .B2(n15895), .A(n18794), .ZN(n16616) );
  NOR3_X1 U18927 ( .A1(n15899), .A2(n9891), .A3(n16616), .ZN(n15898) );
  AOI211_X1 U18928 ( .C1(n15899), .C2(n16432), .A(n15898), .B(n15897), .ZN(
        n15900) );
  OAI21_X1 U18929 ( .B1(n15902), .B2(n15901), .A(n15900), .ZN(n15903) );
  OAI21_X1 U18930 ( .B1(n16482), .B2(n15904), .A(n18248), .ZN(n15972) );
  NOR2_X1 U18931 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18904), .ZN(n18946) );
  INV_X2 U18932 ( .A(n18236), .ZN(n18252) );
  INV_X1 U18933 ( .A(n16499), .ZN(n18713) );
  INV_X1 U18934 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16472) );
  NOR4_X1 U18935 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15906) );
  INV_X1 U18936 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18081) );
  NAND4_X1 U18937 ( .A1(n15906), .A2(n18106), .A3(n17805), .A4(n18081), .ZN(
        n15907) );
  AOI21_X1 U18938 ( .B1(n15910), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15909), .ZN(n17732) );
  NAND2_X1 U18939 ( .A1(n15911), .A2(n15910), .ZN(n17737) );
  NAND2_X1 U18940 ( .A1(n17737), .A2(n15912), .ZN(n15914) );
  INV_X1 U18941 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18035) );
  NAND2_X1 U18942 ( .A1(n17721), .A2(n18035), .ZN(n15913) );
  NOR2_X1 U18943 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15913), .ZN(
        n17673) );
  NAND2_X1 U18944 ( .A1(n17673), .A2(n18021), .ZN(n17666) );
  NAND2_X1 U18945 ( .A1(n15914), .A2(n10226), .ZN(n15915) );
  NAND2_X1 U18946 ( .A1(n18047), .A2(n17737), .ZN(n17671) );
  NOR2_X1 U18947 ( .A1(n17619), .A2(n17849), .ZN(n15918) );
  NAND2_X1 U18948 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17954) );
  AND2_X1 U18949 ( .A1(n17833), .A2(n17954), .ZN(n15917) );
  AOI22_X1 U18950 ( .A1(n17833), .A2(n21110), .B1(n15964), .B2(n9851), .ZN(
        n15921) );
  XNOR2_X1 U18951 ( .A(n16472), .B(n15921), .ZN(n16475) );
  AOI22_X1 U18952 ( .A1(n18252), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18070), 
        .B2(n16475), .ZN(n15931) );
  INV_X1 U18953 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17945) );
  NOR3_X1 U18954 ( .A1(n21110), .A2(n17945), .A3(n16472), .ZN(n16461) );
  INV_X1 U18955 ( .A(n16461), .ZN(n15924) );
  NOR2_X1 U18956 ( .A1(n15922), .A2(n15924), .ZN(n16470) );
  NOR2_X1 U18957 ( .A1(n17985), .A2(n18242), .ZN(n18241) );
  INV_X1 U18958 ( .A(n18241), .ZN(n18258) );
  NOR2_X1 U18959 ( .A1(n15924), .A2(n15923), .ZN(n16449) );
  OR2_X1 U18960 ( .A1(n16449), .A2(n16498), .ZN(n16471) );
  INV_X1 U18961 ( .A(n18196), .ZN(n18256) );
  OAI22_X1 U18962 ( .A1(n16470), .A2(n18258), .B1(n16471), .B2(n18256), .ZN(
        n15968) );
  NAND2_X1 U18963 ( .A1(n18236), .A2(n18242), .ZN(n18211) );
  INV_X1 U18964 ( .A(n15925), .ZN(n18044) );
  NAND2_X1 U18965 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18044), .ZN(
        n18064) );
  NAND3_X1 U18966 ( .A1(n15926), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16459), .ZN(n16497) );
  NOR2_X1 U18967 ( .A1(n18064), .A2(n16497), .ZN(n15928) );
  OAI21_X1 U18968 ( .B1(n17944), .B2(n18045), .A(n18718), .ZN(n17989) );
  INV_X1 U18969 ( .A(n16459), .ZN(n17946) );
  NAND2_X1 U18970 ( .A1(n15926), .A2(n18044), .ZN(n17947) );
  AOI222_X1 U18971 ( .A1(n18749), .A2(n17946), .B1(n18749), .B2(n17947), .C1(
        n17946), .C2(n18718), .ZN(n15927) );
  OAI211_X1 U18972 ( .C1(n18745), .C2(n15928), .A(n17989), .B(n15927), .ZN(
        n15966) );
  AOI211_X1 U18973 ( .C1(n18140), .C2(n17945), .A(n18244), .B(n15966), .ZN(
        n16504) );
  INV_X1 U18974 ( .A(n18006), .ZN(n18161) );
  NAND2_X1 U18975 ( .A1(n18161), .A2(n18248), .ZN(n18237) );
  OAI22_X1 U18976 ( .A1(n18151), .A2(n16504), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18237), .ZN(n15929) );
  OAI21_X1 U18977 ( .B1(n15968), .B2(n15929), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15930) );
  OAI211_X1 U18978 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15972), .A(
        n15931), .B(n15930), .ZN(P3_U2833) );
  INV_X1 U18979 ( .A(n15932), .ZN(n15943) );
  OAI211_X1 U18980 ( .C1(n10914), .C2(n15934), .A(n15933), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15936) );
  OAI21_X1 U18981 ( .B1(n15936), .B2(n20592), .A(n15935), .ZN(n15938) );
  NAND2_X1 U18982 ( .A1(n15936), .A2(n20592), .ZN(n15937) );
  OAI21_X1 U18983 ( .B1(n15939), .B2(n15938), .A(n15937), .ZN(n15940) );
  AOI222_X1 U18984 ( .A1(n15941), .A2(n20663), .B1(n15941), .B2(n15940), .C1(
        n20663), .C2(n15940), .ZN(n15942) );
  AOI222_X1 U18985 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15943), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15942), .C1(n15943), 
        .C2(n15942), .ZN(n15951) );
  OAI21_X1 U18986 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15944), .ZN(n15945) );
  NAND4_X1 U18987 ( .A1(n15948), .A2(n15947), .A3(n15946), .A4(n15945), .ZN(
        n15949) );
  AOI211_X1 U18988 ( .C1(n15951), .C2(n20240), .A(n15950), .B(n15949), .ZN(
        n15963) );
  NAND3_X1 U18989 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20881), .A3(n20868), 
        .ZN(n15952) );
  AOI22_X1 U18990 ( .A1(n15955), .A2(n15954), .B1(n15953), .B2(n15952), .ZN(
        n16263) );
  OAI221_X1 U18991 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15963), 
        .A(n16263), .ZN(n16271) );
  AND2_X1 U18992 ( .A1(n20955), .A2(n15956), .ZN(n15957) );
  NOR2_X1 U18993 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15957), .ZN(n15961) );
  AOI211_X1 U18994 ( .C1(n20881), .C2(n20870), .A(n15958), .B(n16269), .ZN(
        n15959) );
  NAND2_X1 U18995 ( .A1(n16271), .A2(n15959), .ZN(n15960) );
  AOI22_X1 U18996 ( .A1(n16271), .A2(n15961), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15960), .ZN(n15962) );
  OAI21_X1 U18997 ( .B1(n15963), .B2(n20057), .A(n15962), .ZN(P1_U3161) );
  INV_X1 U18998 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16460) );
  NAND2_X1 U18999 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16460), .ZN(
        n15971) );
  OAI21_X1 U19000 ( .B1(n15965), .B2(n16460), .A(n16445), .ZN(n16457) );
  AOI22_X1 U19001 ( .A1(n18252), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n18070), 
        .B2(n16457), .ZN(n15970) );
  AOI21_X1 U19002 ( .B1(n18248), .B2(n15966), .A(n18244), .ZN(n15967) );
  OAI21_X1 U19003 ( .B1(n16461), .B2(n18237), .A(n15967), .ZN(n16491) );
  OAI21_X1 U19004 ( .B1(n16491), .B2(n15968), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15969) );
  OAI211_X1 U19005 ( .C1(n15972), .C2(n15971), .A(n15970), .B(n15969), .ZN(
        P3_U2832) );
  INV_X1 U19006 ( .A(HOLD), .ZN(n20873) );
  INV_X1 U19007 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20889) );
  NAND2_X1 U19008 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20889), .ZN(n20878) );
  AOI21_X1 U19009 ( .B1(n20881), .B2(P1_STATE_REG_1__SCAN_IN), .A(n15973), 
        .ZN(n15975) );
  OAI211_X1 U19010 ( .C1(n20889), .C2(n20873), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n15974) );
  OAI211_X1 U19011 ( .C1(n20873), .C2(n20878), .A(n15975), .B(n15974), .ZN(
        P1_U3195) );
  AND2_X1 U19012 ( .A1(n20184), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19013 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15976) );
  NOR3_X1 U19014 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19926), .A3(n19924), 
        .ZN(n16414) );
  NOR4_X1 U19015 ( .A1(n15976), .A2(n16422), .A3(n16429), .A4(n16414), .ZN(
        P2_U3178) );
  AOI221_X1 U19016 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16429), .C1(n15977), .C2(
        n16429), .A(n19868), .ZN(n20040) );
  INV_X1 U19017 ( .A(n20040), .ZN(n20041) );
  NOR2_X1 U19018 ( .A1(n15978), .A2(n20041), .ZN(P2_U3047) );
  NAND3_X1 U19019 ( .A1(n18277), .A2(n18281), .A3(n15979), .ZN(n15980) );
  NAND2_X1 U19020 ( .A1(n18307), .A2(n17316), .ZN(n17467) );
  INV_X1 U19021 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17543) );
  INV_X1 U19022 ( .A(n17316), .ZN(n15982) );
  AOI22_X1 U19023 ( .A1(n17466), .A2(BUF2_REG_0__SCAN_IN), .B1(n17465), .B2(
        n15985), .ZN(n15986) );
  OAI221_X1 U19024 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17467), .C1(n17543), 
        .C2(n17316), .A(n15986), .ZN(P3_U2735) );
  AOI221_X1 U19025 ( .B1(n20102), .B2(n20916), .C1(n15988), .C2(n20916), .A(
        n15987), .ZN(n15991) );
  OAI22_X1 U19026 ( .A1(n20098), .A2(n15989), .B1(n16081), .B2(n20117), .ZN(
        n15990) );
  AOI211_X1 U19027 ( .C1(n20139), .C2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15991), .B(n15990), .ZN(n15994) );
  NOR2_X1 U19028 ( .A1(n16077), .A2(n20128), .ZN(n15992) );
  AOI21_X1 U19029 ( .B1(n16079), .B2(n20119), .A(n15992), .ZN(n15993) );
  NAND2_X1 U19030 ( .A1(n15994), .A2(n15993), .ZN(P1_U2817) );
  NOR2_X1 U19031 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n20102), .ZN(n16007) );
  INV_X1 U19032 ( .A(n15995), .ZN(n15996) );
  NOR3_X1 U19033 ( .A1(n20102), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n15996), 
        .ZN(n15999) );
  OAI22_X1 U19034 ( .A1(n20117), .A2(n14261), .B1(n15997), .B2(n20111), .ZN(
        n15998) );
  AOI211_X1 U19035 ( .C1(n20140), .C2(n16000), .A(n15999), .B(n15998), .ZN(
        n16001) );
  OAI21_X1 U19036 ( .B1(n16002), .B2(n20104), .A(n16001), .ZN(n16003) );
  AOI221_X1 U19037 ( .B1(n16012), .B2(P1_REIP_REG_22__SCAN_IN), .C1(n16007), 
        .C2(P1_REIP_REG_22__SCAN_IN), .A(n16003), .ZN(n16004) );
  OAI21_X1 U19038 ( .B1(n20128), .B2(n16005), .A(n16004), .ZN(P1_U2818) );
  INV_X1 U19039 ( .A(n16006), .ZN(n16009) );
  AOI22_X1 U19040 ( .A1(n16009), .A2(n20140), .B1(n16008), .B2(n16007), .ZN(
        n16016) );
  AOI22_X1 U19041 ( .A1(n20143), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20139), .ZN(n16015) );
  AOI22_X1 U19042 ( .A1(n16011), .A2(n20119), .B1(n20145), .B2(n16010), .ZN(
        n16014) );
  NAND2_X1 U19043 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n16012), .ZN(n16013) );
  NAND4_X1 U19044 ( .A1(n16016), .A2(n16015), .A3(n16014), .A4(n16013), .ZN(
        P1_U2819) );
  OAI22_X1 U19045 ( .A1(n16018), .A2(n20128), .B1(n16017), .B2(n20117), .ZN(
        n16019) );
  AOI211_X1 U19046 ( .C1(n20139), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16236), .B(n16019), .ZN(n16029) );
  XNOR2_X1 U19047 ( .A(P1_REIP_REG_19__SCAN_IN), .B(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n16025) );
  AND2_X1 U19048 ( .A1(n16021), .A2(n16020), .ZN(n16022) );
  NOR2_X1 U19049 ( .A1(n16023), .A2(n16022), .ZN(n16050) );
  OAI22_X1 U19050 ( .A1(n16040), .A2(n16025), .B1(n16050), .B2(n16024), .ZN(
        n16026) );
  AOI21_X1 U19051 ( .B1(n16027), .B2(n20119), .A(n16026), .ZN(n16028) );
  OAI211_X1 U19052 ( .C1(n16030), .C2(n20098), .A(n16029), .B(n16028), .ZN(
        P1_U2821) );
  OAI22_X1 U19053 ( .A1(n16050), .A2(n14563), .B1(n16031), .B2(n20117), .ZN(
        n16032) );
  AOI211_X1 U19054 ( .C1(n20139), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16032), .B(n16236), .ZN(n16033) );
  INV_X1 U19055 ( .A(n16033), .ZN(n16037) );
  OAI22_X1 U19056 ( .A1(n16035), .A2(n20104), .B1(n20128), .B2(n16034), .ZN(
        n16036) );
  AOI211_X1 U19057 ( .C1(n16038), .C2(n20140), .A(n16037), .B(n16036), .ZN(
        n16039) );
  OAI21_X1 U19058 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n16040), .A(n16039), 
        .ZN(P1_U2822) );
  AOI21_X1 U19059 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n16041), .A(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16049) );
  INV_X1 U19060 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n16083) );
  OAI22_X1 U19061 ( .A1(n20117), .A2(n16083), .B1(n16042), .B2(n20111), .ZN(
        n16043) );
  AOI211_X1 U19062 ( .C1(n20140), .C2(n16091), .A(n16236), .B(n16043), .ZN(
        n16048) );
  AOI21_X1 U19063 ( .B1(n16046), .B2(n16045), .A(n16044), .ZN(n16147) );
  AOI22_X1 U19064 ( .A1(n16092), .A2(n20119), .B1(n20145), .B2(n16147), .ZN(
        n16047) );
  OAI211_X1 U19065 ( .C1(n16050), .C2(n16049), .A(n16048), .B(n16047), .ZN(
        P1_U2823) );
  AOI22_X1 U19066 ( .A1(n16101), .A2(n20119), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n16051), .ZN(n16061) );
  OR2_X1 U19067 ( .A1(n16053), .A2(n16052), .ZN(n16055) );
  AND2_X1 U19068 ( .A1(n16055), .A2(n16054), .ZN(n16153) );
  AOI22_X1 U19069 ( .A1(n16153), .A2(n20145), .B1(n20143), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n16056) );
  OAI211_X1 U19070 ( .C1(n20111), .C2(n16057), .A(n16056), .B(n20227), .ZN(
        n16058) );
  AOI211_X1 U19071 ( .C1(n20140), .C2(n16100), .A(n16059), .B(n16058), .ZN(
        n16060) );
  NAND2_X1 U19072 ( .A1(n16061), .A2(n16060), .ZN(P1_U2825) );
  AOI22_X1 U19073 ( .A1(n16109), .A2(n20140), .B1(n20145), .B2(n16182), .ZN(
        n16066) );
  AOI22_X1 U19074 ( .A1(n20143), .A2(P1_EBX_REG_12__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20139), .ZN(n16065) );
  INV_X1 U19075 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n16073) );
  INV_X1 U19076 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n16184) );
  AOI221_X1 U19077 ( .B1(n16073), .B2(n16184), .C1(n16074), .C2(n16184), .A(
        n16062), .ZN(n16063) );
  AOI21_X1 U19078 ( .B1(n16108), .B2(n20119), .A(n16063), .ZN(n16064) );
  NAND4_X1 U19079 ( .A1(n16066), .A2(n16065), .A3(n16064), .A4(n20227), .ZN(
        P1_U2828) );
  AOI21_X1 U19080 ( .B1(n20139), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16236), .ZN(n16069) );
  INV_X1 U19081 ( .A(n16067), .ZN(n16189) );
  AOI22_X1 U19082 ( .A1(n16189), .A2(n20145), .B1(n20143), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n16068) );
  OAI211_X1 U19083 ( .C1(n16120), .C2(n20098), .A(n16069), .B(n16068), .ZN(
        n16070) );
  AOI21_X1 U19084 ( .B1(n20119), .B2(n16117), .A(n16070), .ZN(n16071) );
  OAI221_X1 U19085 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16074), .C1(n16073), 
        .C2(n16072), .A(n16071), .ZN(P1_U2829) );
  INV_X1 U19086 ( .A(n16075), .ZN(n20157) );
  NOR2_X1 U19087 ( .A1(n16077), .A2(n16076), .ZN(n16078) );
  AOI21_X1 U19088 ( .B1(n16079), .B2(n20157), .A(n16078), .ZN(n16080) );
  OAI21_X1 U19089 ( .B1(n20161), .B2(n16081), .A(n16080), .ZN(P1_U2849) );
  AOI22_X1 U19090 ( .A1(n16092), .A2(n20157), .B1(n20156), .B2(n16147), .ZN(
        n16082) );
  OAI21_X1 U19091 ( .B1(n20161), .B2(n16083), .A(n16082), .ZN(P1_U2855) );
  AOI22_X1 U19092 ( .A1(n16101), .A2(n20157), .B1(n20156), .B2(n16153), .ZN(
        n16084) );
  OAI21_X1 U19093 ( .B1(n20161), .B2(n16085), .A(n16084), .ZN(P1_U2857) );
  NAND2_X1 U19094 ( .A1(n16087), .A2(n16086), .ZN(n16088) );
  NOR2_X1 U19095 ( .A1(n16088), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16089) );
  MUX2_X1 U19096 ( .A(n16089), .B(n16088), .S(n16112), .Z(n16090) );
  XNOR2_X1 U19097 ( .A(n16090), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16152) );
  AOI22_X1 U19098 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16236), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16094) );
  AOI22_X1 U19099 ( .A1(n16092), .A2(n16140), .B1(n16091), .B2(n16138), .ZN(
        n16093) );
  OAI211_X1 U19100 ( .C1(n16152), .C2(n20063), .A(n16094), .B(n16093), .ZN(
        P1_U2982) );
  INV_X1 U19101 ( .A(n16095), .ZN(n16096) );
  OAI21_X1 U19102 ( .B1(n16097), .B2(n16112), .A(n16096), .ZN(n16099) );
  XNOR2_X1 U19103 ( .A(n14449), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16098) );
  XNOR2_X1 U19104 ( .A(n16099), .B(n16098), .ZN(n16160) );
  AOI22_X1 U19105 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16236), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16103) );
  AOI22_X1 U19106 ( .A1(n16101), .A2(n16140), .B1(n16100), .B2(n16138), .ZN(
        n16102) );
  OAI211_X1 U19107 ( .C1(n16160), .C2(n20063), .A(n16103), .B(n16102), .ZN(
        P1_U2984) );
  OAI21_X1 U19108 ( .B1(n16106), .B2(n16105), .A(n16104), .ZN(n16107) );
  INV_X1 U19109 ( .A(n16107), .ZN(n16188) );
  AOI22_X1 U19110 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16236), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16111) );
  AOI22_X1 U19111 ( .A1(n16138), .A2(n16109), .B1(n16140), .B2(n16108), .ZN(
        n16110) );
  OAI211_X1 U19112 ( .C1(n16188), .C2(n20063), .A(n16111), .B(n16110), .ZN(
        P1_U2987) );
  AOI22_X1 U19113 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16236), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16119) );
  NAND3_X1 U19114 ( .A1(n16113), .A2(n16112), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16115) );
  NAND2_X1 U19115 ( .A1(n16115), .A2(n16114), .ZN(n16116) );
  XOR2_X1 U19116 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16116), .Z(
        n16190) );
  AOI22_X1 U19117 ( .A1(n16141), .A2(n16190), .B1(n16140), .B2(n16117), .ZN(
        n16118) );
  OAI211_X1 U19118 ( .C1(n16135), .C2(n16120), .A(n16119), .B(n16118), .ZN(
        P1_U2988) );
  AOI22_X1 U19119 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16236), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16127) );
  XNOR2_X1 U19120 ( .A(n16123), .B(n16122), .ZN(n16124) );
  XNOR2_X1 U19121 ( .A(n16121), .B(n16124), .ZN(n16230) );
  AOI22_X1 U19122 ( .A1(n16230), .A2(n16141), .B1(n16125), .B2(n16140), .ZN(
        n16126) );
  OAI211_X1 U19123 ( .C1(n16135), .C2(n20099), .A(n16127), .B(n16126), .ZN(
        P1_U2992) );
  AOI22_X1 U19124 ( .A1(n16128), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16236), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16134) );
  NAND2_X1 U19125 ( .A1(n16131), .A2(n16130), .ZN(n16132) );
  XNOR2_X1 U19126 ( .A(n16129), .B(n16132), .ZN(n16238) );
  AOI22_X1 U19127 ( .A1(n16141), .A2(n16238), .B1(n20158), .B2(n16140), .ZN(
        n16133) );
  OAI211_X1 U19128 ( .C1(n16135), .C2(n20114), .A(n16134), .B(n16133), .ZN(
        P1_U2993) );
  XOR2_X1 U19129 ( .A(n16136), .B(n16137), .Z(n16250) );
  INV_X1 U19130 ( .A(n20133), .ZN(n16139) );
  AOI222_X1 U19131 ( .A1(n16250), .A2(n16141), .B1(n16140), .B2(n16139), .C1(
        n20126), .C2(n16138), .ZN(n16143) );
  INV_X1 U19132 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20896) );
  NOR2_X1 U19133 ( .A1(n20227), .A2(n20896), .ZN(n16242) );
  INV_X1 U19134 ( .A(n16242), .ZN(n16142) );
  OAI211_X1 U19135 ( .C1(n11303), .C2(n16144), .A(n16143), .B(n16142), .ZN(
        P1_U2994) );
  OAI21_X1 U19136 ( .B1(n16145), .B2(n16154), .A(n14446), .ZN(n16149) );
  INV_X1 U19137 ( .A(n16146), .ZN(n16148) );
  AOI22_X1 U19138 ( .A1(n16149), .A2(n16148), .B1(n16243), .B2(n16147), .ZN(
        n16151) );
  NAND2_X1 U19139 ( .A1(n16236), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16150) );
  OAI211_X1 U19140 ( .C1(n16152), .C2(n20230), .A(n16151), .B(n16150), .ZN(
        P1_U3014) );
  AOI22_X1 U19141 ( .A1(n16153), .A2(n16243), .B1(n16236), .B2(
        P1_REIP_REG_15__SCAN_IN), .ZN(n16159) );
  INV_X1 U19142 ( .A(n16154), .ZN(n16156) );
  AOI22_X1 U19143 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16157), .B1(
        n16156), .B2(n16155), .ZN(n16158) );
  OAI211_X1 U19144 ( .C1(n16160), .C2(n20230), .A(n16159), .B(n16158), .ZN(
        P1_U3016) );
  AOI22_X1 U19145 ( .A1(n16236), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n16162), 
        .B2(n16161), .ZN(n16170) );
  AOI22_X1 U19146 ( .A1(n16165), .A2(n16243), .B1(n16164), .B2(n16163), .ZN(
        n16169) );
  AOI22_X1 U19147 ( .A1(n16167), .A2(n16249), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16166), .ZN(n16168) );
  NAND3_X1 U19148 ( .A1(n16170), .A2(n16169), .A3(n16168), .ZN(P1_U3018) );
  NOR2_X1 U19149 ( .A1(n16178), .A2(n16194), .ZN(n16181) );
  OAI21_X1 U19150 ( .B1(n20229), .B2(n16172), .A(n16171), .ZN(n16217) );
  INV_X1 U19151 ( .A(n16217), .ZN(n16177) );
  AOI22_X1 U19152 ( .A1(n16175), .A2(n16174), .B1(n16218), .B2(n16173), .ZN(
        n16176) );
  NAND2_X1 U19153 ( .A1(n16177), .A2(n16176), .ZN(n16191) );
  AOI21_X1 U19154 ( .B1(n20223), .B2(n16178), .A(n16191), .ZN(n16179) );
  INV_X1 U19155 ( .A(n16179), .ZN(n16180) );
  MUX2_X1 U19156 ( .A(n16181), .B(n16180), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n16186) );
  NAND2_X1 U19157 ( .A1(n16182), .A2(n16243), .ZN(n16183) );
  OAI21_X1 U19158 ( .B1(n16184), .B2(n20227), .A(n16183), .ZN(n16185) );
  NOR2_X1 U19159 ( .A1(n16186), .A2(n16185), .ZN(n16187) );
  OAI21_X1 U19160 ( .B1(n16188), .B2(n20230), .A(n16187), .ZN(P1_U3019) );
  AOI22_X1 U19161 ( .A1(n16189), .A2(n16243), .B1(n16236), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16193) );
  AOI22_X1 U19162 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16191), .B1(
        n16249), .B2(n16190), .ZN(n16192) );
  OAI211_X1 U19163 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16194), .A(
        n16193), .B(n16192), .ZN(P1_U3020) );
  OAI21_X1 U19164 ( .B1(n16197), .B2(n16196), .A(n16195), .ZN(n16198) );
  AOI21_X1 U19165 ( .B1(n16221), .B2(n16198), .A(n16217), .ZN(n16215) );
  OAI22_X1 U19166 ( .A1(n16201), .A2(n16200), .B1(n16199), .B2(n20227), .ZN(
        n16202) );
  AOI21_X1 U19167 ( .B1(n16249), .B2(n16203), .A(n16202), .ZN(n16206) );
  OAI211_X1 U19168 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n16210), .B(n16204), .ZN(n16205) );
  OAI211_X1 U19169 ( .C1(n16215), .C2(n16207), .A(n16206), .B(n16205), .ZN(
        P1_U3021) );
  INV_X1 U19170 ( .A(n16208), .ZN(n16209) );
  AOI21_X1 U19171 ( .B1(n20082), .B2(n16243), .A(n16209), .ZN(n16213) );
  AOI22_X1 U19172 ( .A1(n16211), .A2(n16249), .B1(n16210), .B2(n16214), .ZN(
        n16212) );
  OAI211_X1 U19173 ( .C1(n16215), .C2(n16214), .A(n16213), .B(n16212), .ZN(
        P1_U3022) );
  NAND2_X1 U19174 ( .A1(n16216), .A2(n16246), .ZN(n16253) );
  AOI21_X1 U19175 ( .B1(n16219), .B2(n16218), .A(n16217), .ZN(n16247) );
  OAI21_X1 U19176 ( .B1(n16220), .B2(n16253), .A(n16247), .ZN(n16237) );
  AOI21_X1 U19177 ( .B1(n16225), .B2(n16221), .A(n16237), .ZN(n16233) );
  INV_X1 U19178 ( .A(n16222), .ZN(n16223) );
  AOI222_X1 U19179 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n16236), .B1(n16243), 
        .B2(n16224), .C1(n16249), .C2(n16223), .ZN(n16227) );
  NOR2_X1 U19180 ( .A1(n16225), .A2(n16241), .ZN(n16229) );
  OAI221_X1 U19181 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16228), .C2(n16122), .A(
        n16229), .ZN(n16226) );
  OAI211_X1 U19182 ( .C1(n16233), .C2(n16228), .A(n16227), .B(n16226), .ZN(
        P1_U3023) );
  AOI22_X1 U19183 ( .A1(n20108), .A2(n16243), .B1(n16236), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16232) );
  AOI22_X1 U19184 ( .A1(n16230), .A2(n16249), .B1(n16122), .B2(n16229), .ZN(
        n16231) );
  OAI211_X1 U19185 ( .C1(n16233), .C2(n16122), .A(n16232), .B(n16231), .ZN(
        P1_U3024) );
  XNOR2_X1 U19186 ( .A(n16235), .B(n16234), .ZN(n20155) );
  AOI22_X1 U19187 ( .A1(n20155), .A2(n16243), .B1(n16236), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16240) );
  AOI22_X1 U19188 ( .A1(n16238), .A2(n16249), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16237), .ZN(n16239) );
  OAI211_X1 U19189 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16241), .A(
        n16240), .B(n16239), .ZN(P1_U3025) );
  AOI21_X1 U19190 ( .B1(n16244), .B2(n16243), .A(n16242), .ZN(n16245) );
  OAI21_X1 U19191 ( .B1(n16247), .B2(n16246), .A(n16245), .ZN(n16248) );
  AOI21_X1 U19192 ( .B1(n16250), .B2(n16249), .A(n16248), .ZN(n16251) );
  OAI21_X1 U19193 ( .B1(n16253), .B2(n16252), .A(n16251), .ZN(P1_U3026) );
  NAND3_X1 U19194 ( .A1(n16256), .A2(n16255), .A3(n16254), .ZN(n16257) );
  OAI21_X1 U19195 ( .B1(n16259), .B2(n16258), .A(n16257), .ZN(P1_U3468) );
  NAND4_X1 U19196 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20870), .A4(n20951), .ZN(n16260) );
  AND2_X1 U19197 ( .A1(n16261), .A2(n16260), .ZN(n20869) );
  INV_X1 U19198 ( .A(n16262), .ZN(n16264) );
  AOI21_X1 U19199 ( .B1(n20869), .B2(n16264), .A(n16263), .ZN(n16268) );
  NOR2_X1 U19200 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20951), .ZN(n16265) );
  NOR2_X1 U19201 ( .A1(n20868), .A2(n16265), .ZN(n16266) );
  AOI21_X1 U19202 ( .B1(n16266), .B2(n16271), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n16267) );
  NOR3_X1 U19203 ( .A1(n16269), .A2(n16268), .A3(n16267), .ZN(P1_U3162) );
  OAI221_X1 U19204 ( .B1(n20669), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20669), 
        .C2(n16271), .A(n16270), .ZN(P1_U3466) );
  OAI22_X1 U19205 ( .A1(n16273), .A2(n16272), .B1(n12451), .B2(n19188), .ZN(
        n16274) );
  INV_X1 U19206 ( .A(n16274), .ZN(n16285) );
  OAI22_X1 U19207 ( .A1(n16275), .A2(n19194), .B1(n19097), .B2(n21100), .ZN(
        n16276) );
  INV_X1 U19208 ( .A(n16276), .ZN(n16284) );
  NOR2_X1 U19209 ( .A1(n16277), .A2(n19154), .ZN(n16278) );
  AOI21_X1 U19210 ( .B1(n16279), .B2(n19190), .A(n16278), .ZN(n16283) );
  NAND2_X1 U19211 ( .A1(n16281), .A2(n16280), .ZN(n16282) );
  NAND4_X1 U19212 ( .A1(n16285), .A2(n16284), .A3(n16283), .A4(n16282), .ZN(
        P2_U2824) );
  AOI211_X1 U19213 ( .C1(n16288), .C2(n16286), .A(n16287), .B(n19929), .ZN(
        n16296) );
  AOI22_X1 U19214 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19198), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19170), .ZN(n16290) );
  NAND2_X1 U19215 ( .A1(n19183), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16289) );
  OAI211_X1 U19216 ( .C1(n16291), .C2(n19194), .A(n16290), .B(n16289), .ZN(
        n16292) );
  INV_X1 U19217 ( .A(n16292), .ZN(n16293) );
  OAI21_X1 U19218 ( .B1(n16294), .B2(n19174), .A(n16293), .ZN(n16295) );
  AOI211_X1 U19219 ( .C1(n19185), .C2(n16297), .A(n16296), .B(n16295), .ZN(
        n16298) );
  INV_X1 U19220 ( .A(n16298), .ZN(P2_U2829) );
  INV_X1 U19221 ( .A(n16299), .ZN(n16300) );
  OAI22_X1 U19222 ( .A1(n16301), .A2(n19174), .B1(n16300), .B2(n19154), .ZN(
        n16302) );
  INV_X1 U19223 ( .A(n16302), .ZN(n16311) );
  AOI211_X1 U19224 ( .C1(n16305), .C2(n16303), .A(n16304), .B(n19929), .ZN(
        n16309) );
  AOI22_X1 U19225 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19183), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19170), .ZN(n16306) );
  OAI21_X1 U19226 ( .B1(n16307), .B2(n19194), .A(n16306), .ZN(n16308) );
  AOI211_X1 U19227 ( .C1(n19198), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16309), .B(n16308), .ZN(n16310) );
  NAND2_X1 U19228 ( .A1(n16311), .A2(n16310), .ZN(P2_U2831) );
  AOI22_X1 U19229 ( .A1(n19207), .A2(n16312), .B1(n19264), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16316) );
  AOI22_X1 U19230 ( .A1(n19209), .A2(BUF2_REG_20__SCAN_IN), .B1(n19208), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16315) );
  AOI22_X1 U19231 ( .A1(n16313), .A2(n19269), .B1(n19265), .B2(n18995), .ZN(
        n16314) );
  NAND3_X1 U19232 ( .A1(n16316), .A2(n16315), .A3(n16314), .ZN(P2_U2899) );
  AOI22_X1 U19233 ( .A1(n19207), .A2(n16317), .B1(n19264), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16322) );
  AOI22_X1 U19234 ( .A1(n19209), .A2(BUF2_REG_18__SCAN_IN), .B1(n19208), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16321) );
  INV_X1 U19235 ( .A(n16318), .ZN(n19018) );
  AOI22_X1 U19236 ( .A1(n16319), .A2(n19269), .B1(n19265), .B2(n19018), .ZN(
        n16320) );
  NAND3_X1 U19237 ( .A1(n16322), .A2(n16321), .A3(n16320), .ZN(P2_U2901) );
  AOI22_X1 U19238 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19348), .B1(n16351), 
        .B2(n19110), .ZN(n16330) );
  OAI22_X1 U19239 ( .A1(n16326), .A2(n16325), .B1(n16324), .B2(n16323), .ZN(
        n16327) );
  AOI21_X1 U19240 ( .B1(n19351), .B2(n16328), .A(n16327), .ZN(n16329) );
  OAI211_X1 U19241 ( .C1(n16359), .C2(n16331), .A(n16330), .B(n16329), .ZN(
        P2_U3005) );
  AOI22_X1 U19242 ( .A1(n19349), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19348), .ZN(n16344) );
  INV_X1 U19243 ( .A(n16332), .ZN(n16334) );
  OAI21_X1 U19244 ( .B1(n15300), .B2(n16334), .A(n16333), .ZN(n16338) );
  NAND2_X1 U19245 ( .A1(n16336), .A2(n16335), .ZN(n16337) );
  XNOR2_X1 U19246 ( .A(n16338), .B(n16337), .ZN(n16363) );
  OAI21_X1 U19247 ( .B1(n16339), .B2(n16341), .A(n16340), .ZN(n16342) );
  INV_X1 U19248 ( .A(n16342), .ZN(n16360) );
  AOI222_X1 U19249 ( .A1(n16363), .A2(n19355), .B1(n19351), .B2(n16362), .C1(
        n19352), .C2(n16360), .ZN(n16343) );
  OAI211_X1 U19250 ( .C1(n19359), .C2(n16345), .A(n16344), .B(n16343), .ZN(
        P2_U3006) );
  AOI22_X1 U19251 ( .A1(n19349), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19348), .ZN(n16350) );
  INV_X1 U19252 ( .A(n16346), .ZN(n16347) );
  AOI222_X1 U19253 ( .A1(n16348), .A2(n19355), .B1(n19351), .B2(n19137), .C1(
        n19352), .C2(n16347), .ZN(n16349) );
  OAI211_X1 U19254 ( .C1(n19359), .C2(n19135), .A(n16350), .B(n16349), .ZN(
        P2_U3008) );
  AOI22_X1 U19255 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19348), .B1(n16351), 
        .B2(n19147), .ZN(n16357) );
  AOI22_X1 U19256 ( .A1(n16353), .A2(n19355), .B1(n19352), .B2(n16352), .ZN(
        n16354) );
  INV_X1 U19257 ( .A(n16354), .ZN(n16355) );
  AOI21_X1 U19258 ( .B1(n19351), .B2(n19148), .A(n16355), .ZN(n16356) );
  OAI211_X1 U19259 ( .C1(n16359), .C2(n16358), .A(n16357), .B(n16356), .ZN(
        P2_U3009) );
  AOI22_X1 U19260 ( .A1(n16373), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19364), .B2(n19236), .ZN(n16368) );
  AOI222_X1 U19261 ( .A1(n16363), .A2(n19361), .B1(n19369), .B2(n16362), .C1(
        n16361), .C2(n16360), .ZN(n16367) );
  NAND2_X1 U19262 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19348), .ZN(n16366) );
  OAI211_X1 U19263 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16375), .B(n16364), .ZN(n16365) );
  NAND4_X1 U19264 ( .A1(n16368), .A2(n16367), .A3(n16366), .A4(n16365), .ZN(
        P2_U3038) );
  OAI21_X1 U19265 ( .B1(n16370), .B2(n16369), .A(n13556), .ZN(n19238) );
  OAI22_X1 U19266 ( .A1(n16371), .A2(n19238), .B1(n20984), .B2(n19129), .ZN(
        n16372) );
  AOI221_X1 U19267 ( .B1(n16375), .B2(n16374), .C1(n16373), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16372), .ZN(n16379) );
  AOI22_X1 U19268 ( .A1(n16377), .A2(n19361), .B1(n19369), .B2(n16376), .ZN(
        n16378) );
  OAI211_X1 U19269 ( .C1(n19366), .C2(n16380), .A(n16379), .B(n16378), .ZN(
        P2_U3039) );
  MUX2_X1 U19270 ( .A(n16398), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16381), .Z(n16412) );
  INV_X1 U19271 ( .A(n16382), .ZN(n16383) );
  MUX2_X1 U19272 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16383), .S(
        n16402), .Z(n16411) );
  INV_X1 U19273 ( .A(n16384), .ZN(n16389) );
  NOR4_X1 U19274 ( .A1(n16389), .A2(n10092), .A3(n16386), .A4(n16385), .ZN(
        n18957) );
  OAI21_X1 U19275 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18957), .ZN(n16388) );
  OAI211_X1 U19276 ( .C1(n12215), .C2(n12213), .A(n16388), .B(n16387), .ZN(
        n16395) );
  NAND2_X1 U19277 ( .A1(n16389), .A2(n10578), .ZN(n16392) );
  NAND2_X1 U19278 ( .A1(n16394), .A2(n16390), .ZN(n16391) );
  OAI211_X1 U19279 ( .C1(n16394), .C2(n16393), .A(n16392), .B(n16391), .ZN(
        n20048) );
  NOR2_X1 U19280 ( .A1(n16395), .A2(n20048), .ZN(n16396) );
  OAI21_X1 U19281 ( .B1(n16397), .B2(n16402), .A(n16396), .ZN(n16410) );
  INV_X1 U19282 ( .A(n16398), .ZN(n16401) );
  OAI21_X1 U19283 ( .B1(n20042), .B2(n16404), .A(n20033), .ZN(n16399) );
  AOI22_X1 U19284 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16401), .B1(
        n16400), .B2(n16399), .ZN(n16403) );
  OAI211_X1 U19285 ( .C1(n19722), .C2(n16404), .A(n16403), .B(n16402), .ZN(
        n16405) );
  INV_X1 U19286 ( .A(n16405), .ZN(n16406) );
  OAI211_X1 U19287 ( .C1(n20023), .C2(n16406), .A(n16411), .B(n10561), .ZN(
        n16408) );
  AOI22_X1 U19288 ( .A1(n16412), .A2(n10561), .B1(n20023), .B2(n16406), .ZN(
        n16407) );
  AOI21_X1 U19289 ( .B1(n16408), .B2(n16407), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16409) );
  AOI211_X1 U19290 ( .C1(n16412), .C2(n16411), .A(n16410), .B(n16409), .ZN(
        n16428) );
  AOI211_X1 U19291 ( .C1(n16429), .C2(n20044), .A(n16414), .B(n16413), .ZN(
        n16427) );
  INV_X1 U19292 ( .A(n16415), .ZN(n16416) );
  NOR3_X1 U19293 ( .A1(n16418), .A2(n16417), .A3(n16416), .ZN(n16420) );
  NOR3_X1 U19294 ( .A1(n16420), .A2(n16419), .A3(n20035), .ZN(n16423) );
  AOI22_X1 U19295 ( .A1(n19943), .A2(n16423), .B1(n16422), .B2(n16421), .ZN(
        n16425) );
  OAI221_X1 U19296 ( .B1(n19926), .B2(n16428), .C1(n19926), .C2(n16424), .A(
        n16423), .ZN(n19925) );
  NAND2_X1 U19297 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19925), .ZN(n16430) );
  OAI21_X1 U19298 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16425), .A(n16430), 
        .ZN(n16426) );
  OAI211_X1 U19299 ( .C1(n16428), .C2(n18956), .A(n16427), .B(n16426), .ZN(
        P2_U3176) );
  AOI21_X1 U19300 ( .B1(n16430), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16429), 
        .ZN(n16431) );
  INV_X1 U19301 ( .A(n16431), .ZN(P2_U3593) );
  INV_X1 U19302 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18887) );
  NAND2_X1 U19303 ( .A1(n16470), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16433) );
  XNOR2_X1 U19304 ( .A(n18887), .B(n16433), .ZN(n16485) );
  NAND3_X1 U19305 ( .A1(n17939), .A2(n16638), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n17787) );
  NAND2_X1 U19306 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17784) );
  INV_X1 U19307 ( .A(n17784), .ZN(n16839) );
  NAND2_X1 U19308 ( .A1(n16839), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17742) );
  NAND2_X1 U19309 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17743) );
  NAND2_X1 U19310 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17706) );
  INV_X1 U19311 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17687) );
  INV_X1 U19312 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17676) );
  INV_X1 U19313 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17662) );
  NOR2_X1 U19314 ( .A1(n17676), .A2(n17662), .ZN(n17658) );
  INV_X1 U19315 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17622) );
  NAND2_X1 U19316 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17624) );
  NAND2_X1 U19317 ( .A1(n17609), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17589) );
  NAND2_X1 U19318 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17590) );
  NAND2_X1 U19319 ( .A1(n16469), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16439) );
  INV_X1 U19320 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17933) );
  NAND2_X1 U19321 ( .A1(n16452), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16437) );
  INV_X1 U19322 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16664) );
  XNOR2_X2 U19323 ( .A(n16437), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16641) );
  INV_X1 U19324 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18864) );
  NOR2_X1 U19325 ( .A1(n18864), .A2(n18236), .ZN(n16488) );
  INV_X1 U19326 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16455) );
  NOR2_X1 U19327 ( .A1(n18930), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n17782) );
  OAI21_X1 U19328 ( .B1(n17933), .B2(n17648), .A(n18373), .ZN(n17741) );
  INV_X1 U19329 ( .A(n17741), .ZN(n17705) );
  NOR2_X1 U19330 ( .A1(n17705), .A2(n16439), .ZN(n16440) );
  INV_X1 U19331 ( .A(n16440), .ZN(n16454) );
  NOR2_X1 U19332 ( .A1(n16455), .A2(n16454), .ZN(n16442) );
  NOR2_X1 U19333 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17648), .ZN(
        n16477) );
  NAND2_X1 U19334 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n10229), .ZN(
        n16647) );
  NAND2_X1 U19335 ( .A1(n17621), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16651) );
  INV_X1 U19336 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17639) );
  NOR2_X1 U19337 ( .A1(n16651), .A2(n17639), .ZN(n16653) );
  NAND2_X1 U19338 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16653), .ZN(
        n17578) );
  INV_X1 U19339 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16717) );
  NOR2_X1 U19340 ( .A1(n17578), .A2(n16717), .ZN(n16657) );
  INV_X1 U19341 ( .A(n16657), .ZN(n16438) );
  NOR2_X1 U19342 ( .A1(n16438), .A2(n17590), .ZN(n16642) );
  INV_X1 U19343 ( .A(n17782), .ZN(n17938) );
  INV_X2 U19344 ( .A(n18373), .ZN(n18655) );
  NAND2_X1 U19345 ( .A1(n18655), .A2(n16439), .ZN(n16466) );
  OAI211_X1 U19346 ( .C1(n16642), .C2(n17938), .A(n17939), .B(n16466), .ZN(
        n16467) );
  AOI211_X1 U19347 ( .C1(n16440), .C2(n16455), .A(n16477), .B(n16467), .ZN(
        n16453) );
  INV_X1 U19348 ( .A(n16453), .ZN(n16441) );
  MUX2_X1 U19349 ( .A(n16442), .B(n16441), .S(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n16443) );
  AOI211_X1 U19350 ( .C1(n17799), .C2(n16641), .A(n16488), .B(n16443), .ZN(
        n16451) );
  NOR2_X1 U19351 ( .A1(n18887), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16489) );
  INV_X1 U19352 ( .A(n16489), .ZN(n16448) );
  OAI21_X1 U19353 ( .B1(n17833), .B2(n9729), .A(n16444), .ZN(n16447) );
  NAND2_X1 U19354 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18887), .ZN(
        n16484) );
  INV_X1 U19355 ( .A(n16484), .ZN(n16446) );
  NAND2_X1 U19356 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16449), .ZN(
        n16450) );
  XOR2_X1 U19357 ( .A(n18887), .B(n16450), .Z(n16487) );
  NAND2_X1 U19358 ( .A1(n17441), .A2(n17883), .ZN(n17850) );
  INV_X1 U19359 ( .A(n17850), .ZN(n17774) );
  INV_X1 U19360 ( .A(n16452), .ZN(n16476) );
  AOI22_X1 U19361 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16452), .B1(
        n16476), .B2(n16455), .ZN(n16667) );
  AOI21_X1 U19362 ( .B1(n16455), .B2(n16454), .A(n16453), .ZN(n16456) );
  AOI21_X1 U19363 ( .B1(n16667), .B2(n17799), .A(n16456), .ZN(n16465) );
  INV_X1 U19364 ( .A(n17883), .ZN(n17942) );
  OAI22_X1 U19365 ( .A1(n16470), .A2(n17943), .B1(n17942), .B2(n16471), .ZN(
        n16458) );
  AOI22_X1 U19366 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16458), .B1(
        n17748), .B2(n16457), .ZN(n16464) );
  NAND2_X1 U19367 ( .A1(n18252), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16463) );
  NOR2_X1 U19368 ( .A1(n17944), .A2(n17751), .ZN(n17656) );
  AND2_X1 U19369 ( .A1(n16459), .A2(n17656), .ZN(n17604) );
  NAND3_X1 U19370 ( .A1(n16461), .A2(n17604), .A3(n16460), .ZN(n16462) );
  NAND4_X1 U19371 ( .A1(n16465), .A2(n16464), .A3(n16463), .A4(n16462), .ZN(
        P3_U2800) );
  INV_X1 U19372 ( .A(n16466), .ZN(n16468) );
  AOI22_X1 U19373 ( .A1(n16469), .A2(n16468), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16467), .ZN(n16481) );
  AOI211_X1 U19374 ( .C1(n16472), .C2(n16502), .A(n16470), .B(n17943), .ZN(
        n16474) );
  AOI211_X1 U19375 ( .C1(n16472), .C2(n16501), .A(n17942), .B(n16471), .ZN(
        n16473) );
  AOI211_X1 U19376 ( .C1(n16475), .C2(n17748), .A(n16474), .B(n16473), .ZN(
        n16480) );
  NAND2_X1 U19377 ( .A1(n18252), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16479) );
  OAI21_X1 U19378 ( .B1(n16642), .B2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16476), .ZN(n16677) );
  INV_X1 U19379 ( .A(n16677), .ZN(n16679) );
  OAI21_X1 U19380 ( .B1(n16477), .B2(n17799), .A(n16679), .ZN(n16478) );
  NAND4_X1 U19381 ( .A1(n16481), .A2(n16480), .A3(n16479), .A4(n16478), .ZN(
        P3_U2801) );
  NAND2_X1 U19382 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16482), .ZN(
        n16483) );
  OAI22_X1 U19383 ( .A1(n17985), .A2(n16485), .B1(n16484), .B2(n16483), .ZN(
        n16486) );
  AOI21_X1 U19384 ( .B1(n16487), .B2(n18126), .A(n16486), .ZN(n16494) );
  INV_X1 U19385 ( .A(n18237), .ZN(n18203) );
  AOI21_X1 U19386 ( .B1(n16489), .B2(n18203), .A(n16488), .ZN(n16493) );
  OAI211_X1 U19387 ( .C1(n16494), .C2(n18242), .A(n16493), .B(n16492), .ZN(
        P3_U2831) );
  AOI22_X1 U19388 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17849), .B1(
        n17833), .B2(n21110), .ZN(n17585) );
  AOI21_X1 U19389 ( .B1(n17833), .B2(n17597), .A(n17595), .ZN(n17584) );
  NOR2_X1 U19390 ( .A1(n17585), .A2(n17584), .ZN(n17583) );
  OAI211_X1 U19391 ( .C1(n17595), .C2(n16495), .A(n21110), .B(n18070), .ZN(
        n16509) );
  OAI22_X1 U19392 ( .A1(n18127), .A2(n17985), .B1(n18125), .B2(n18166), .ZN(
        n18041) );
  AOI21_X1 U19393 ( .B1(n18043), .B2(n18041), .A(n16496), .ZN(n18010) );
  NOR2_X1 U19394 ( .A1(n18010), .A2(n18242), .ZN(n18016) );
  NOR2_X1 U19395 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16497), .ZN(
        n17588) );
  AOI22_X1 U19396 ( .A1(n18252), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n18016), 
        .B2(n17588), .ZN(n16508) );
  NAND2_X1 U19397 ( .A1(n16499), .A2(n16498), .ZN(n18099) );
  NOR3_X1 U19398 ( .A1(n16500), .A2(n17583), .A3(n18099), .ZN(n16506) );
  AOI22_X1 U19399 ( .A1(n18716), .A2(n16502), .B1(n18126), .B2(n16501), .ZN(
        n16503) );
  NAND2_X1 U19400 ( .A1(n16504), .A2(n16503), .ZN(n16505) );
  OAI211_X1 U19401 ( .C1(n16506), .C2(n16505), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18236), .ZN(n16507) );
  OAI211_X1 U19402 ( .C1(n17583), .C2(n16509), .A(n16508), .B(n16507), .ZN(
        P3_U2834) );
  NOR3_X1 U19403 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16511) );
  NOR4_X1 U19404 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16510) );
  INV_X2 U19405 ( .A(n16603), .ZN(U215) );
  NAND4_X1 U19406 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16511), .A3(n16510), .A4(
        U215), .ZN(U213) );
  INV_X1 U19407 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16605) );
  INV_X2 U19408 ( .A(U214), .ZN(n16566) );
  INV_X1 U19409 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n21081) );
  OAI222_X1 U19410 ( .A1(U212), .A2(n16605), .B1(n16568), .B2(n19420), .C1(
        U214), .C2(n21081), .ZN(U216) );
  INV_X1 U19411 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16514) );
  INV_X2 U19412 ( .A(U212), .ZN(n16565) );
  AOI22_X1 U19413 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16565), .ZN(n16513) );
  OAI21_X1 U19414 ( .B1(n16514), .B2(n16568), .A(n16513), .ZN(U217) );
  INV_X1 U19415 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16516) );
  AOI22_X1 U19416 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16565), .ZN(n16515) );
  OAI21_X1 U19417 ( .B1(n16516), .B2(n16568), .A(n16515), .ZN(U218) );
  INV_X1 U19418 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n21131) );
  AOI22_X1 U19419 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16565), .ZN(n16517) );
  OAI21_X1 U19420 ( .B1(n21131), .B2(n16568), .A(n16517), .ZN(U219) );
  INV_X1 U19421 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16519) );
  AOI22_X1 U19422 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16565), .ZN(n16518) );
  OAI21_X1 U19423 ( .B1(n16519), .B2(n16568), .A(n16518), .ZN(U220) );
  INV_X1 U19424 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16521) );
  AOI22_X1 U19425 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16565), .ZN(n16520) );
  OAI21_X1 U19426 ( .B1(n16521), .B2(n16568), .A(n16520), .ZN(U221) );
  INV_X1 U19427 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16523) );
  AOI22_X1 U19428 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16565), .ZN(n16522) );
  OAI21_X1 U19429 ( .B1(n16523), .B2(n16568), .A(n16522), .ZN(U222) );
  INV_X1 U19430 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16525) );
  AOI22_X1 U19431 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16565), .ZN(n16524) );
  OAI21_X1 U19432 ( .B1(n16525), .B2(n16568), .A(n16524), .ZN(U223) );
  INV_X1 U19433 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16527) );
  AOI22_X1 U19434 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16565), .ZN(n16526) );
  OAI21_X1 U19435 ( .B1(n16527), .B2(n16568), .A(n16526), .ZN(U224) );
  INV_X1 U19436 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16529) );
  AOI22_X1 U19437 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16565), .ZN(n16528) );
  OAI21_X1 U19438 ( .B1(n16529), .B2(n16568), .A(n16528), .ZN(U225) );
  INV_X1 U19439 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19406) );
  AOI22_X1 U19440 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16565), .ZN(n16530) );
  OAI21_X1 U19441 ( .B1(n19406), .B2(n16568), .A(n16530), .ZN(U226) );
  INV_X1 U19442 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16532) );
  AOI22_X1 U19443 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16565), .ZN(n16531) );
  OAI21_X1 U19444 ( .B1(n16532), .B2(n16568), .A(n16531), .ZN(U227) );
  INV_X1 U19445 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16534) );
  AOI22_X1 U19446 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16565), .ZN(n16533) );
  OAI21_X1 U19447 ( .B1(n16534), .B2(n16568), .A(n16533), .ZN(U228) );
  INV_X1 U19448 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16536) );
  AOI22_X1 U19449 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16565), .ZN(n16535) );
  OAI21_X1 U19450 ( .B1(n16536), .B2(n16568), .A(n16535), .ZN(U229) );
  INV_X1 U19451 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16538) );
  AOI22_X1 U19452 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16565), .ZN(n16537) );
  OAI21_X1 U19453 ( .B1(n16538), .B2(n16568), .A(n16537), .ZN(U230) );
  INV_X1 U19454 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16540) );
  AOI22_X1 U19455 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16565), .ZN(n16539) );
  OAI21_X1 U19456 ( .B1(n16540), .B2(n16568), .A(n16539), .ZN(U231) );
  AOI22_X1 U19457 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16565), .ZN(n16541) );
  OAI21_X1 U19458 ( .B1(n13108), .B2(n16568), .A(n16541), .ZN(U232) );
  AOI22_X1 U19459 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16565), .ZN(n16542) );
  OAI21_X1 U19460 ( .B1(n14307), .B2(n16568), .A(n16542), .ZN(U233) );
  AOI22_X1 U19461 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16565), .ZN(n16543) );
  OAI21_X1 U19462 ( .B1(n14313), .B2(n16568), .A(n16543), .ZN(U234) );
  AOI22_X1 U19463 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16565), .ZN(n16544) );
  OAI21_X1 U19464 ( .B1(n16545), .B2(n16568), .A(n16544), .ZN(U235) );
  AOI22_X1 U19465 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16565), .ZN(n16546) );
  OAI21_X1 U19466 ( .B1(n14324), .B2(n16568), .A(n16546), .ZN(U236) );
  AOI22_X1 U19467 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16565), .ZN(n16547) );
  OAI21_X1 U19468 ( .B1(n16548), .B2(n16568), .A(n16547), .ZN(U237) );
  AOI22_X1 U19469 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16565), .ZN(n16549) );
  OAI21_X1 U19470 ( .B1(n13622), .B2(n16568), .A(n16549), .ZN(U238) );
  AOI22_X1 U19471 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16565), .ZN(n16550) );
  OAI21_X1 U19472 ( .B1(n16551), .B2(n16568), .A(n16550), .ZN(U239) );
  AOI22_X1 U19473 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16565), .ZN(n16552) );
  OAI21_X1 U19474 ( .B1(n12646), .B2(n16568), .A(n16552), .ZN(U240) );
  INV_X1 U19475 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16554) );
  AOI22_X1 U19476 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16565), .ZN(n16553) );
  OAI21_X1 U19477 ( .B1(n16554), .B2(n16568), .A(n16553), .ZN(U241) );
  AOI22_X1 U19478 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16565), .ZN(n16555) );
  OAI21_X1 U19479 ( .B1(n16556), .B2(n16568), .A(n16555), .ZN(U242) );
  INV_X1 U19480 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16558) );
  AOI22_X1 U19481 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16565), .ZN(n16557) );
  OAI21_X1 U19482 ( .B1(n16558), .B2(n16568), .A(n16557), .ZN(U243) );
  INV_X1 U19483 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16560) );
  AOI22_X1 U19484 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16565), .ZN(n16559) );
  OAI21_X1 U19485 ( .B1(n16560), .B2(n16568), .A(n16559), .ZN(U244) );
  INV_X1 U19486 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16562) );
  AOI22_X1 U19487 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16565), .ZN(n16561) );
  OAI21_X1 U19488 ( .B1(n16562), .B2(n16568), .A(n16561), .ZN(U245) );
  INV_X1 U19489 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16564) );
  AOI22_X1 U19490 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16565), .ZN(n16563) );
  OAI21_X1 U19491 ( .B1(n16564), .B2(n16568), .A(n16563), .ZN(U246) );
  INV_X1 U19492 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16569) );
  AOI22_X1 U19493 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16566), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16565), .ZN(n16567) );
  OAI21_X1 U19494 ( .B1(n16569), .B2(n16568), .A(n16567), .ZN(U247) );
  OAI22_X1 U19495 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16603), .ZN(n16570) );
  INV_X1 U19496 ( .A(n16570), .ZN(U251) );
  OAI22_X1 U19497 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16603), .ZN(n16571) );
  INV_X1 U19498 ( .A(n16571), .ZN(U252) );
  OAI22_X1 U19499 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16603), .ZN(n16572) );
  INV_X1 U19500 ( .A(n16572), .ZN(U253) );
  OAI22_X1 U19501 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16603), .ZN(n16573) );
  INV_X1 U19502 ( .A(n16573), .ZN(U254) );
  OAI22_X1 U19503 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16603), .ZN(n16574) );
  INV_X1 U19504 ( .A(n16574), .ZN(U255) );
  OAI22_X1 U19505 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16603), .ZN(n16575) );
  INV_X1 U19506 ( .A(n16575), .ZN(U256) );
  OAI22_X1 U19507 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16603), .ZN(n16576) );
  INV_X1 U19508 ( .A(n16576), .ZN(U257) );
  OAI22_X1 U19509 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16603), .ZN(n16577) );
  INV_X1 U19510 ( .A(n16577), .ZN(U258) );
  OAI22_X1 U19511 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16603), .ZN(n16578) );
  INV_X1 U19512 ( .A(n16578), .ZN(U259) );
  OAI22_X1 U19513 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16597), .ZN(n16579) );
  INV_X1 U19514 ( .A(n16579), .ZN(U260) );
  OAI22_X1 U19515 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16597), .ZN(n16580) );
  INV_X1 U19516 ( .A(n16580), .ZN(U261) );
  OAI22_X1 U19517 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16603), .ZN(n16581) );
  INV_X1 U19518 ( .A(n16581), .ZN(U262) );
  OAI22_X1 U19519 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16603), .ZN(n16582) );
  INV_X1 U19520 ( .A(n16582), .ZN(U263) );
  OAI22_X1 U19521 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16603), .ZN(n16583) );
  INV_X1 U19522 ( .A(n16583), .ZN(U264) );
  OAI22_X1 U19523 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16603), .ZN(n16584) );
  INV_X1 U19524 ( .A(n16584), .ZN(U265) );
  OAI22_X1 U19525 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16597), .ZN(n16585) );
  INV_X1 U19526 ( .A(n16585), .ZN(U266) );
  OAI22_X1 U19527 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16597), .ZN(n16586) );
  INV_X1 U19528 ( .A(n16586), .ZN(U267) );
  OAI22_X1 U19529 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16597), .ZN(n16587) );
  INV_X1 U19530 ( .A(n16587), .ZN(U268) );
  OAI22_X1 U19531 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16597), .ZN(n16588) );
  INV_X1 U19532 ( .A(n16588), .ZN(U269) );
  OAI22_X1 U19533 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16597), .ZN(n16589) );
  INV_X1 U19534 ( .A(n16589), .ZN(U270) );
  OAI22_X1 U19535 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16597), .ZN(n16590) );
  INV_X1 U19536 ( .A(n16590), .ZN(U271) );
  OAI22_X1 U19537 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16603), .ZN(n16591) );
  INV_X1 U19538 ( .A(n16591), .ZN(U272) );
  OAI22_X1 U19539 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16603), .ZN(n16592) );
  INV_X1 U19540 ( .A(n16592), .ZN(U273) );
  OAI22_X1 U19541 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16597), .ZN(n16593) );
  INV_X1 U19542 ( .A(n16593), .ZN(U274) );
  OAI22_X1 U19543 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16603), .ZN(n16594) );
  INV_X1 U19544 ( .A(n16594), .ZN(U275) );
  OAI22_X1 U19545 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16603), .ZN(n16595) );
  INV_X1 U19546 ( .A(n16595), .ZN(U276) );
  OAI22_X1 U19547 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16603), .ZN(n16596) );
  INV_X1 U19548 ( .A(n16596), .ZN(U277) );
  OAI22_X1 U19549 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16597), .ZN(n16598) );
  INV_X1 U19550 ( .A(n16598), .ZN(U278) );
  OAI22_X1 U19551 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16603), .ZN(n16599) );
  INV_X1 U19552 ( .A(n16599), .ZN(U279) );
  OAI22_X1 U19553 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16603), .ZN(n16600) );
  INV_X1 U19554 ( .A(n16600), .ZN(U280) );
  OAI22_X1 U19555 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16603), .ZN(n16602) );
  INV_X1 U19556 ( .A(n16602), .ZN(U281) );
  INV_X1 U19557 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19418) );
  AOI22_X1 U19558 ( .A1(n16603), .A2(n16605), .B1(n19418), .B2(U215), .ZN(U282) );
  INV_X1 U19559 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16604) );
  AOI222_X1 U19560 ( .A1(n21081), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16605), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16604), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16606) );
  INV_X2 U19561 ( .A(n16608), .ZN(n16607) );
  INV_X1 U19562 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18824) );
  INV_X1 U19563 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19962) );
  AOI22_X1 U19564 ( .A1(n16607), .A2(n18824), .B1(n19962), .B2(n16608), .ZN(
        U347) );
  INV_X1 U19565 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18822) );
  INV_X1 U19566 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19960) );
  AOI22_X1 U19567 ( .A1(n16607), .A2(n18822), .B1(n19960), .B2(n16608), .ZN(
        U348) );
  INV_X1 U19568 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n21129) );
  INV_X1 U19569 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19959) );
  AOI22_X1 U19570 ( .A1(n16607), .A2(n21129), .B1(n19959), .B2(n16608), .ZN(
        U349) );
  INV_X1 U19571 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18819) );
  INV_X1 U19572 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19958) );
  AOI22_X1 U19573 ( .A1(n16607), .A2(n18819), .B1(n19958), .B2(n16608), .ZN(
        U350) );
  INV_X1 U19574 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18817) );
  INV_X1 U19575 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19957) );
  AOI22_X1 U19576 ( .A1(n16607), .A2(n18817), .B1(n19957), .B2(n16608), .ZN(
        U351) );
  INV_X1 U19577 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18814) );
  INV_X1 U19578 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19956) );
  AOI22_X1 U19579 ( .A1(n16607), .A2(n18814), .B1(n19956), .B2(n16608), .ZN(
        U352) );
  INV_X1 U19580 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18813) );
  INV_X1 U19581 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19955) );
  AOI22_X1 U19582 ( .A1(n16607), .A2(n18813), .B1(n19955), .B2(n16608), .ZN(
        U353) );
  INV_X1 U19583 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18811) );
  AOI22_X1 U19584 ( .A1(n16607), .A2(n18811), .B1(n19954), .B2(n16608), .ZN(
        U354) );
  INV_X1 U19585 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18865) );
  INV_X1 U19586 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19996) );
  AOI22_X1 U19587 ( .A1(n16607), .A2(n18865), .B1(n19996), .B2(n16608), .ZN(
        U355) );
  INV_X1 U19588 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18863) );
  INV_X1 U19589 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19993) );
  AOI22_X1 U19590 ( .A1(n16607), .A2(n18863), .B1(n19993), .B2(n16608), .ZN(
        U356) );
  INV_X1 U19591 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18860) );
  INV_X1 U19592 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19991) );
  AOI22_X1 U19593 ( .A1(n16607), .A2(n18860), .B1(n19991), .B2(n16608), .ZN(
        U357) );
  INV_X1 U19594 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18859) );
  INV_X1 U19595 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19988) );
  AOI22_X1 U19596 ( .A1(n16607), .A2(n18859), .B1(n19988), .B2(n16608), .ZN(
        U358) );
  INV_X1 U19597 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18857) );
  INV_X1 U19598 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19987) );
  AOI22_X1 U19599 ( .A1(n16607), .A2(n18857), .B1(n19987), .B2(n16608), .ZN(
        U359) );
  INV_X1 U19600 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18854) );
  INV_X1 U19601 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19986) );
  AOI22_X1 U19602 ( .A1(n16607), .A2(n18854), .B1(n19986), .B2(n16608), .ZN(
        U360) );
  INV_X1 U19603 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18852) );
  INV_X1 U19604 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19984) );
  AOI22_X1 U19605 ( .A1(n16607), .A2(n18852), .B1(n19984), .B2(n16608), .ZN(
        U361) );
  INV_X1 U19606 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18850) );
  INV_X1 U19607 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19982) );
  AOI22_X1 U19608 ( .A1(n16607), .A2(n18850), .B1(n19982), .B2(n16608), .ZN(
        U362) );
  INV_X1 U19609 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18848) );
  INV_X1 U19610 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19980) );
  AOI22_X1 U19611 ( .A1(n16607), .A2(n18848), .B1(n19980), .B2(n16608), .ZN(
        U363) );
  INV_X1 U19612 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18846) );
  INV_X1 U19613 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19978) );
  AOI22_X1 U19614 ( .A1(n16607), .A2(n18846), .B1(n19978), .B2(n16608), .ZN(
        U364) );
  INV_X1 U19615 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18810) );
  INV_X1 U19616 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19953) );
  AOI22_X1 U19617 ( .A1(n16607), .A2(n18810), .B1(n19953), .B2(n16608), .ZN(
        U365) );
  INV_X1 U19618 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18843) );
  INV_X1 U19619 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19977) );
  AOI22_X1 U19620 ( .A1(n16607), .A2(n18843), .B1(n19977), .B2(n16608), .ZN(
        U366) );
  INV_X1 U19621 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18842) );
  INV_X1 U19622 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19976) );
  AOI22_X1 U19623 ( .A1(n16607), .A2(n18842), .B1(n19976), .B2(n16608), .ZN(
        U367) );
  INV_X1 U19624 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18840) );
  INV_X1 U19625 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19974) );
  AOI22_X1 U19626 ( .A1(n16607), .A2(n18840), .B1(n19974), .B2(n16608), .ZN(
        U368) );
  INV_X1 U19627 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18837) );
  INV_X1 U19628 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19973) );
  AOI22_X1 U19629 ( .A1(n16607), .A2(n18837), .B1(n19973), .B2(n16608), .ZN(
        U369) );
  INV_X1 U19630 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18836) );
  INV_X1 U19631 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19971) );
  AOI22_X1 U19632 ( .A1(n16607), .A2(n18836), .B1(n19971), .B2(n16608), .ZN(
        U370) );
  INV_X1 U19633 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18834) );
  INV_X1 U19634 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19969) );
  AOI22_X1 U19635 ( .A1(n16607), .A2(n18834), .B1(n19969), .B2(n16608), .ZN(
        U371) );
  INV_X1 U19636 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18832) );
  INV_X1 U19637 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19968) );
  AOI22_X1 U19638 ( .A1(n16607), .A2(n18832), .B1(n19968), .B2(n16608), .ZN(
        U372) );
  INV_X1 U19639 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18830) );
  INV_X1 U19640 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19967) );
  AOI22_X1 U19641 ( .A1(n16607), .A2(n18830), .B1(n19967), .B2(n16608), .ZN(
        U373) );
  INV_X1 U19642 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18828) );
  INV_X1 U19643 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19965) );
  AOI22_X1 U19644 ( .A1(n16607), .A2(n18828), .B1(n19965), .B2(n16608), .ZN(
        U374) );
  INV_X1 U19645 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18826) );
  INV_X1 U19646 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19963) );
  AOI22_X1 U19647 ( .A1(n16607), .A2(n18826), .B1(n19963), .B2(n16608), .ZN(
        U375) );
  INV_X1 U19648 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18808) );
  INV_X1 U19649 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19952) );
  AOI22_X1 U19650 ( .A1(n16607), .A2(n18808), .B1(n19952), .B2(n16608), .ZN(
        U376) );
  NOR2_X1 U19651 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18804), .ZN(n18793) );
  NAND2_X1 U19652 ( .A1(n18787), .A2(n18804), .ZN(n18792) );
  INV_X1 U19653 ( .A(n18792), .ZN(n16609) );
  AOI21_X1 U19654 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18793), .A(n16609), 
        .ZN(n18786) );
  INV_X1 U19655 ( .A(n18786), .ZN(n18874) );
  AOI21_X1 U19656 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18874), .ZN(n16610) );
  INV_X1 U19657 ( .A(n16610), .ZN(P3_U2633) );
  NAND2_X1 U19658 ( .A1(n18712), .A2(n16617), .ZN(n16611) );
  OAI21_X1 U19659 ( .B1(n18925), .B2(n16611), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16612) );
  OAI21_X1 U19660 ( .B1(n16613), .B2(n18775), .A(n16612), .ZN(P3_U2634) );
  AOI21_X1 U19661 ( .B1(n18807), .B2(n18804), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16614) );
  AOI22_X1 U19662 ( .A1(n18939), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16614), 
        .B2(n18940), .ZN(P3_U2635) );
  NOR2_X1 U19663 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n16615) );
  OAI21_X1 U19664 ( .B1(n16615), .B2(BS16), .A(n18874), .ZN(n18873) );
  OAI21_X1 U19665 ( .B1(n18874), .B2(n16638), .A(n18873), .ZN(P3_U2636) );
  AND3_X1 U19666 ( .A1(n18712), .A2(n16617), .A3(n16616), .ZN(n18723) );
  NOR2_X1 U19667 ( .A1(n18723), .A2(n18925), .ZN(n18920) );
  OAI21_X1 U19668 ( .B1(n18920), .B2(n16619), .A(n16618), .ZN(P3_U2637) );
  NOR4_X1 U19669 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16623) );
  NOR4_X1 U19670 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16622) );
  NOR4_X1 U19671 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16621) );
  NOR4_X1 U19672 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16620) );
  NAND4_X1 U19673 ( .A1(n16623), .A2(n16622), .A3(n16621), .A4(n16620), .ZN(
        n16629) );
  NOR4_X1 U19674 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16627) );
  AOI211_X1 U19675 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_21__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16626) );
  NOR4_X1 U19676 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16625) );
  NOR4_X1 U19677 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16624) );
  NAND4_X1 U19678 ( .A1(n16627), .A2(n16626), .A3(n16625), .A4(n16624), .ZN(
        n16628) );
  NOR2_X1 U19679 ( .A1(n16629), .A2(n16628), .ZN(n18915) );
  INV_X1 U19680 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16631) );
  NOR3_X1 U19681 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16632) );
  OAI21_X1 U19682 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16632), .A(n18915), .ZN(
        n16630) );
  OAI21_X1 U19683 ( .B1(n18915), .B2(n16631), .A(n16630), .ZN(P3_U2638) );
  INV_X1 U19684 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18911) );
  INV_X1 U19685 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21132) );
  AOI21_X1 U19686 ( .B1(n18911), .B2(n21132), .A(n16632), .ZN(n16634) );
  INV_X1 U19687 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16633) );
  INV_X1 U19688 ( .A(n18915), .ZN(n18917) );
  AOI22_X1 U19689 ( .A1(n18915), .A2(n16634), .B1(n16633), .B2(n18917), .ZN(
        P3_U2639) );
  NAND4_X1 U19690 ( .A1(n18930), .A2(n18932), .A3(n16638), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18781) );
  INV_X1 U19691 ( .A(n18781), .ZN(n17006) );
  INV_X1 U19692 ( .A(n18616), .ZN(n18776) );
  NOR2_X1 U19693 ( .A1(n18775), .A2(n18776), .ZN(n18769) );
  AOI211_X1 U19694 ( .C1(n16635), .C2(n18281), .A(n9890), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18766) );
  INV_X1 U19695 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18861) );
  INV_X1 U19696 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18858) );
  NOR2_X1 U19697 ( .A1(n18861), .A2(n18858), .ZN(n16636) );
  INV_X1 U19698 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18856) );
  INV_X1 U19699 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18851) );
  INV_X1 U19700 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18838) );
  INV_X1 U19701 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18833) );
  INV_X1 U19702 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18827) );
  INV_X1 U19703 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18809) );
  NOR2_X1 U19704 ( .A1(n18911), .A2(n18809), .ZN(n16996) );
  AND2_X1 U19705 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n16996), .ZN(n16926) );
  NAND3_X1 U19706 ( .A1(n16926), .A2(P3_REIP_REG_5__SCAN_IN), .A3(
        P3_REIP_REG_4__SCAN_IN), .ZN(n16874) );
  NAND3_X1 U19707 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n16875) );
  NOR2_X1 U19708 ( .A1(n16874), .A2(n16875), .ZN(n16889) );
  NAND4_X1 U19709 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16889), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16862) );
  NOR2_X1 U19710 ( .A1(n18827), .A2(n16862), .ZN(n16851) );
  NAND3_X1 U19711 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16851), .ZN(n16841) );
  NOR2_X1 U19712 ( .A1(n18833), .A2(n16841), .ZN(n16815) );
  NAND2_X1 U19713 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n16815), .ZN(n16803) );
  NOR2_X1 U19714 ( .A1(n18838), .A2(n16803), .ZN(n16751) );
  NAND3_X1 U19715 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n16752) );
  NAND2_X1 U19716 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16760) );
  NOR2_X1 U19717 ( .A1(n16752), .A2(n16760), .ZN(n16740) );
  NAND3_X1 U19718 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16751), .A3(n16740), 
        .ZN(n16718) );
  NOR2_X1 U19719 ( .A1(n18851), .A2(n16718), .ZN(n16724) );
  NAND2_X1 U19720 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16724), .ZN(n16703) );
  NOR2_X1 U19721 ( .A1(n18856), .A2(n16703), .ZN(n16658) );
  NOR2_X1 U19722 ( .A1(n16658), .A2(n17018), .ZN(n16704) );
  NOR2_X1 U19723 ( .A1(n16999), .A2(n16704), .ZN(n16706) );
  OAI221_X1 U19724 ( .B1(n17018), .B2(P3_REIP_REG_29__SCAN_IN), .C1(n17018), 
        .C2(n16636), .A(n16706), .ZN(n16674) );
  INV_X1 U19725 ( .A(n16640), .ZN(n16637) );
  AOI211_X4 U19726 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18929), .A(n18766), .B(
        n16637), .ZN(n17026) );
  AOI22_X1 U19727 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n16674), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n17026), .ZN(n16663) );
  NAND2_X1 U19728 ( .A1(n16638), .A2(n18794), .ZN(n16639) );
  NOR3_X1 U19729 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16998) );
  INV_X1 U19730 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16991) );
  NAND2_X1 U19731 ( .A1(n16998), .A2(n16991), .ZN(n16990) );
  NOR2_X1 U19732 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16990), .ZN(n16964) );
  INV_X1 U19733 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17283) );
  NAND2_X1 U19734 ( .A1(n16964), .A2(n17283), .ZN(n16960) );
  INV_X1 U19735 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16939) );
  NAND2_X1 U19736 ( .A1(n16942), .A2(n16939), .ZN(n16936) );
  INV_X1 U19737 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16912) );
  NAND2_X1 U19738 ( .A1(n16903), .A2(n16912), .ZN(n16887) );
  INV_X1 U19739 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16883) );
  NAND2_X1 U19740 ( .A1(n16886), .A2(n16883), .ZN(n16882) );
  NAND2_X1 U19741 ( .A1(n16869), .A2(n17215), .ZN(n16852) );
  NAND2_X1 U19742 ( .A1(n16840), .A2(n16838), .ZN(n16831) );
  NAND2_X1 U19743 ( .A1(n16816), .A2(n16813), .ZN(n16806) );
  NAND2_X1 U19744 ( .A1(n16794), .A2(n17134), .ZN(n16787) );
  NAND2_X1 U19745 ( .A1(n16775), .A2(n17116), .ZN(n16769) );
  INV_X1 U19746 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16747) );
  NAND2_X1 U19747 ( .A1(n16755), .A2(n16747), .ZN(n16746) );
  NOR2_X1 U19748 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16746), .ZN(n16731) );
  NAND2_X1 U19749 ( .A1(n16731), .A2(n16723), .ZN(n16722) );
  NOR2_X1 U19750 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16722), .ZN(n16707) );
  NAND2_X1 U19751 ( .A1(n16707), .A2(n17069), .ZN(n16699) );
  NOR2_X1 U19752 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16699), .ZN(n16685) );
  NAND2_X1 U19753 ( .A1(n16685), .A2(n17057), .ZN(n16665) );
  NOR2_X1 U19754 ( .A1(n16997), .A2(n16665), .ZN(n16668) );
  INV_X1 U19755 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16661) );
  INV_X1 U19756 ( .A(n17006), .ZN(n17016) );
  INV_X1 U19757 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n21125) );
  NAND2_X1 U19758 ( .A1(n16657), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16656) );
  AOI21_X1 U19759 ( .B1(n21125), .B2(n16656), .A(n16642), .ZN(n17581) );
  NAND2_X1 U19760 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17686), .ZN(
        n17660) );
  INV_X1 U19761 ( .A(n16647), .ZN(n16648) );
  AOI21_X1 U19762 ( .B1(n17687), .B2(n17660), .A(n16648), .ZN(n17690) );
  NOR2_X1 U19763 ( .A1(n17933), .A2(n17728), .ZN(n16643) );
  INV_X1 U19764 ( .A(n16643), .ZN(n16818) );
  NOR2_X1 U19765 ( .A1(n17727), .A2(n16818), .ZN(n17701) );
  XOR2_X1 U19766 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B(n17701), .Z(
        n17720) );
  INV_X1 U19767 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16980) );
  AOI21_X1 U19768 ( .B1(n17727), .B2(n16818), .A(n17701), .ZN(n17730) );
  NOR2_X1 U19769 ( .A1(n17720), .A2(n16798), .ZN(n16797) );
  NOR2_X1 U19770 ( .A1(n16797), .A2(n16979), .ZN(n16786) );
  INV_X1 U19771 ( .A(n16786), .ZN(n16646) );
  INV_X1 U19772 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17709) );
  NAND2_X1 U19773 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17701), .ZN(
        n16644) );
  AOI22_X1 U19774 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17686), .B1(
        n17709), .B2(n16644), .ZN(n17703) );
  INV_X1 U19775 ( .A(n17703), .ZN(n16645) );
  NAND2_X1 U19776 ( .A1(n16646), .A2(n16645), .ZN(n16784) );
  NOR2_X1 U19777 ( .A1(n16773), .A2(n16979), .ZN(n16765) );
  AOI22_X1 U19778 ( .A1(n16648), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n17676), .B2(n16647), .ZN(n17679) );
  NAND2_X1 U19779 ( .A1(n16648), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16649) );
  AOI21_X1 U19780 ( .B1(n17662), .B2(n16649), .A(n17621), .ZN(n17665) );
  NOR2_X1 U19781 ( .A1(n16753), .A2(n16979), .ZN(n16742) );
  OAI21_X1 U19782 ( .B1(n17621), .B2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16651), .ZN(n16650) );
  INV_X1 U19783 ( .A(n16650), .ZN(n17649) );
  NOR2_X1 U19784 ( .A1(n16742), .A2(n17649), .ZN(n16741) );
  OR2_X1 U19785 ( .A1(n16741), .A2(n16979), .ZN(n16732) );
  AOI21_X1 U19786 ( .B1(n16651), .B2(n17639), .A(n16653), .ZN(n17636) );
  NAND2_X1 U19787 ( .A1(n16732), .A2(n16652), .ZN(n16733) );
  OAI21_X1 U19788 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16653), .A(
        n17578), .ZN(n16654) );
  INV_X1 U19789 ( .A(n16654), .ZN(n17627) );
  NOR2_X1 U19790 ( .A1(n16720), .A2(n17627), .ZN(n16719) );
  OR2_X1 U19791 ( .A1(n16719), .A2(n16979), .ZN(n16708) );
  AOI21_X1 U19792 ( .B1(n17578), .B2(n16717), .A(n16657), .ZN(n17613) );
  INV_X1 U19793 ( .A(n17613), .ZN(n16655) );
  NAND2_X1 U19794 ( .A1(n16708), .A2(n16655), .ZN(n16709) );
  OAI21_X1 U19795 ( .B1(n16657), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16656), .ZN(n17599) );
  INV_X1 U19796 ( .A(n17599), .ZN(n16695) );
  NOR2_X1 U19797 ( .A1(n16693), .A2(n16979), .ZN(n16687) );
  OR2_X1 U19798 ( .A1(n16686), .A2(n16979), .ZN(n16676) );
  NOR4_X1 U19799 ( .A1(n16667), .A2(n16979), .A3(n17016), .A4(n16666), .ZN(
        n16660) );
  INV_X1 U19800 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18866) );
  NAND2_X1 U19801 ( .A1(n16983), .A2(n16658), .ZN(n16692) );
  NOR3_X1 U19802 ( .A1(n18861), .A2(n18858), .A3(n16692), .ZN(n16675) );
  NAND2_X1 U19803 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16675), .ZN(n16671) );
  AOI221_X1 U19804 ( .B1(P3_REIP_REG_31__SCAN_IN), .B2(P3_REIP_REG_30__SCAN_IN), .C1(n18864), .C2(n18866), .A(n16671), .ZN(n16659) );
  AOI211_X1 U19805 ( .C1(n16668), .C2(n16661), .A(n16660), .B(n16659), .ZN(
        n16662) );
  OAI211_X1 U19806 ( .C1(n16664), .C2(n17014), .A(n16663), .B(n16662), .ZN(
        P3_U2640) );
  AOI22_X1 U19807 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16940), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n16674), .ZN(n16670) );
  NAND2_X1 U19808 ( .A1(n17025), .A2(n16665), .ZN(n16682) );
  OAI211_X1 U19809 ( .C1(P3_REIP_REG_30__SCAN_IN), .C2(n16671), .A(n16670), 
        .B(n16669), .ZN(P3_U2641) );
  NOR2_X1 U19810 ( .A1(n16685), .A2(n17057), .ZN(n16683) );
  INV_X1 U19811 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18862) );
  INV_X1 U19812 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16672) );
  OAI22_X1 U19813 ( .A1(n16672), .A2(n17014), .B1(n17017), .B2(n17057), .ZN(
        n16673) );
  AOI221_X1 U19814 ( .B1(n16675), .B2(n18862), .C1(n16674), .C2(
        P3_REIP_REG_29__SCAN_IN), .A(n16673), .ZN(n16681) );
  INV_X1 U19815 ( .A(n16676), .ZN(n16678) );
  OAI221_X1 U19816 ( .B1(n16679), .B2(n16678), .C1(n16677), .C2(n16676), .A(
        n17006), .ZN(n16680) );
  OAI211_X1 U19817 ( .C1(n16683), .C2(n16682), .A(n16681), .B(n16680), .ZN(
        P3_U2642) );
  NOR3_X1 U19818 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18858), .A3(n16692), 
        .ZN(n16684) );
  AOI21_X1 U19819 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17026), .A(n16684), .ZN(
        n16691) );
  OAI21_X1 U19820 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16692), .A(n16706), 
        .ZN(n16698) );
  AOI211_X1 U19821 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16699), .A(n16685), .B(
        n16997), .ZN(n16689) );
  AOI211_X1 U19822 ( .C1(n17581), .C2(n16687), .A(n16686), .B(n17016), .ZN(
        n16688) );
  AOI211_X1 U19823 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16698), .A(n16689), 
        .B(n16688), .ZN(n16690) );
  OAI211_X1 U19824 ( .C1(n21125), .C2(n17014), .A(n16691), .B(n16690), .ZN(
        P3_U2643) );
  AOI22_X1 U19825 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16940), .B1(
        n17026), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16702) );
  INV_X1 U19826 ( .A(n16692), .ZN(n16697) );
  AOI211_X1 U19827 ( .C1(n16695), .C2(n16694), .A(n16693), .B(n17016), .ZN(
        n16696) );
  AOI221_X1 U19828 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16698), .C1(n16697), 
        .C2(n16698), .A(n16696), .ZN(n16701) );
  OAI211_X1 U19829 ( .C1(n16707), .C2(n17069), .A(n17025), .B(n16699), .ZN(
        n16700) );
  NAND3_X1 U19830 ( .A1(n16702), .A2(n16701), .A3(n16700), .ZN(P3_U2644) );
  INV_X1 U19831 ( .A(n16703), .ZN(n16705) );
  AOI22_X1 U19832 ( .A1(n17026), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16705), 
        .B2(n16704), .ZN(n16716) );
  INV_X1 U19833 ( .A(n16706), .ZN(n16714) );
  AOI211_X1 U19834 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16722), .A(n16707), .B(
        n16997), .ZN(n16713) );
  INV_X1 U19835 ( .A(n16708), .ZN(n16711) );
  INV_X1 U19836 ( .A(n16709), .ZN(n16710) );
  AOI211_X1 U19837 ( .C1(n17613), .C2(n16711), .A(n16710), .B(n17016), .ZN(
        n16712) );
  AOI211_X1 U19838 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16714), .A(n16713), 
        .B(n16712), .ZN(n16715) );
  OAI211_X1 U19839 ( .C1(n16717), .C2(n17014), .A(n16716), .B(n16715), .ZN(
        P3_U2645) );
  AOI22_X1 U19840 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16940), .B1(
        n17026), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16728) );
  NOR2_X1 U19841 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17018), .ZN(n16729) );
  INV_X1 U19842 ( .A(n16718), .ZN(n16730) );
  OAI21_X1 U19843 ( .B1(n16730), .B2(n17018), .A(n17027), .ZN(n16745) );
  AOI211_X1 U19844 ( .C1(n17627), .C2(n16720), .A(n16719), .B(n17016), .ZN(
        n16721) );
  AOI221_X1 U19845 ( .B1(n16729), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n16745), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n16721), .ZN(n16727) );
  OAI211_X1 U19846 ( .C1(n16731), .C2(n16723), .A(n17025), .B(n16722), .ZN(
        n16726) );
  INV_X1 U19847 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18853) );
  NAND3_X1 U19848 ( .A1(n16983), .A2(n16724), .A3(n18853), .ZN(n16725) );
  NAND4_X1 U19849 ( .A1(n16728), .A2(n16727), .A3(n16726), .A4(n16725), .ZN(
        P3_U2646) );
  AOI22_X1 U19850 ( .A1(n17026), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16730), 
        .B2(n16729), .ZN(n16739) );
  AOI211_X1 U19851 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16746), .A(n16731), .B(
        n16997), .ZN(n16737) );
  INV_X1 U19852 ( .A(n16732), .ZN(n16735) );
  INV_X1 U19853 ( .A(n16733), .ZN(n16734) );
  AOI211_X1 U19854 ( .C1(n17636), .C2(n16735), .A(n16734), .B(n17016), .ZN(
        n16736) );
  AOI211_X1 U19855 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16745), .A(n16737), 
        .B(n16736), .ZN(n16738) );
  OAI211_X1 U19856 ( .C1(n17639), .C2(n17014), .A(n16739), .B(n16738), .ZN(
        P3_U2647) );
  NAND2_X1 U19857 ( .A1(n16740), .A2(n16800), .ZN(n16750) );
  AOI211_X1 U19858 ( .C1(n17649), .C2(n16742), .A(n16741), .B(n17016), .ZN(
        n16744) );
  OAI22_X1 U19859 ( .A1(n17622), .A2(n17014), .B1(n17017), .B2(n16747), .ZN(
        n16743) );
  AOI211_X1 U19860 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16745), .A(n16744), 
        .B(n16743), .ZN(n16749) );
  OAI211_X1 U19861 ( .C1(n16755), .C2(n16747), .A(n17025), .B(n16746), .ZN(
        n16748) );
  OAI211_X1 U19862 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16750), .A(n16749), 
        .B(n16748), .ZN(P3_U2648) );
  INV_X1 U19863 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18847) );
  NAND2_X1 U19864 ( .A1(n16751), .A2(n17027), .ZN(n16796) );
  NAND2_X1 U19865 ( .A1(n17027), .A2(n17018), .ZN(n17024) );
  OAI21_X1 U19866 ( .B1(n16752), .B2(n16796), .A(n17024), .ZN(n16778) );
  AOI211_X1 U19867 ( .C1(n17665), .C2(n16754), .A(n16753), .B(n17016), .ZN(
        n16759) );
  AOI211_X1 U19868 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16769), .A(n16755), .B(
        n16997), .ZN(n16758) );
  OAI22_X1 U19869 ( .A1(n17662), .A2(n17014), .B1(n17017), .B2(n16756), .ZN(
        n16757) );
  NOR3_X1 U19870 ( .A1(n16759), .A2(n16758), .A3(n16757), .ZN(n16762) );
  INV_X1 U19871 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18844) );
  NAND3_X1 U19872 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n16800), .ZN(n16779) );
  NOR2_X1 U19873 ( .A1(n18844), .A2(n16779), .ZN(n16767) );
  OAI211_X1 U19874 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16767), .B(n16760), .ZN(n16761) );
  OAI211_X1 U19875 ( .C1(n18847), .C2(n16778), .A(n16762), .B(n16761), .ZN(
        P3_U2649) );
  AOI22_X1 U19876 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16940), .B1(
        n17026), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16772) );
  INV_X1 U19877 ( .A(n16778), .ZN(n16768) );
  INV_X1 U19878 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18845) );
  INV_X1 U19879 ( .A(n16763), .ZN(n16764) );
  AOI211_X1 U19880 ( .C1(n17679), .C2(n16765), .A(n16764), .B(n17016), .ZN(
        n16766) );
  AOI221_X1 U19881 ( .B1(n16768), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n16767), 
        .C2(n18845), .A(n16766), .ZN(n16771) );
  OAI211_X1 U19882 ( .C1(n16775), .C2(n17116), .A(n17025), .B(n16769), .ZN(
        n16770) );
  NAND3_X1 U19883 ( .A1(n16772), .A2(n16771), .A3(n16770), .ZN(P3_U2650) );
  AOI211_X1 U19884 ( .C1(n17690), .C2(n16774), .A(n16773), .B(n17016), .ZN(
        n16777) );
  AOI211_X1 U19885 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16787), .A(n16775), .B(
        n16997), .ZN(n16776) );
  AOI211_X1 U19886 ( .C1(n16940), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16777), .B(n16776), .ZN(n16782) );
  AOI21_X1 U19887 ( .B1(n18844), .B2(n16779), .A(n16778), .ZN(n16780) );
  INV_X1 U19888 ( .A(n16780), .ZN(n16781) );
  OAI211_X1 U19889 ( .C1(n16783), .C2(n17017), .A(n16782), .B(n16781), .ZN(
        P3_U2651) );
  NAND2_X1 U19890 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16800), .ZN(n16793) );
  INV_X1 U19891 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18841) );
  INV_X1 U19892 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18839) );
  AOI22_X1 U19893 ( .A1(n16800), .A2(n18839), .B1(n17024), .B2(n16796), .ZN(
        n16792) );
  INV_X1 U19894 ( .A(n16784), .ZN(n16785) );
  AOI211_X1 U19895 ( .C1(n17703), .C2(n16786), .A(n16785), .B(n17016), .ZN(
        n16790) );
  OAI211_X1 U19896 ( .C1(n16794), .C2(n17134), .A(n17025), .B(n16787), .ZN(
        n16788) );
  OAI211_X1 U19897 ( .C1(n17017), .C2(n17134), .A(n18236), .B(n16788), .ZN(
        n16789) );
  AOI211_X1 U19898 ( .C1(n16940), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16790), .B(n16789), .ZN(n16791) );
  OAI221_X1 U19899 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(n16793), .C1(n18841), 
        .C2(n16792), .A(n16791), .ZN(P3_U2652) );
  INV_X1 U19900 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17717) );
  AOI211_X1 U19901 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16806), .A(n16794), .B(
        n16997), .ZN(n16795) );
  AOI211_X1 U19902 ( .C1(n17026), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18252), .B(
        n16795), .ZN(n16802) );
  AND2_X1 U19903 ( .A1(n17024), .A2(n16796), .ZN(n16811) );
  AOI211_X1 U19904 ( .C1(n17720), .C2(n16798), .A(n16797), .B(n17016), .ZN(
        n16799) );
  AOI221_X1 U19905 ( .B1(n16811), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n16800), 
        .C2(n18839), .A(n16799), .ZN(n16801) );
  OAI211_X1 U19906 ( .C1(n17717), .C2(n17014), .A(n16802), .B(n16801), .ZN(
        P3_U2653) );
  OAI21_X1 U19907 ( .B1(n17018), .B2(n16803), .A(n18838), .ZN(n16810) );
  AOI211_X1 U19908 ( .C1(n17730), .C2(n16805), .A(n16804), .B(n17016), .ZN(
        n16809) );
  OAI211_X1 U19909 ( .C1(n16816), .C2(n16813), .A(n17025), .B(n16806), .ZN(
        n16807) );
  OAI21_X1 U19910 ( .B1(n17014), .B2(n17727), .A(n16807), .ZN(n16808) );
  AOI211_X1 U19911 ( .C1(n16811), .C2(n16810), .A(n16809), .B(n16808), .ZN(
        n16812) );
  OAI211_X1 U19912 ( .C1(n17017), .C2(n16813), .A(n16812), .B(n18236), .ZN(
        P3_U2654) );
  NOR2_X1 U19913 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n17018), .ZN(n16814) );
  AOI22_X1 U19914 ( .A1(n17026), .A2(P3_EBX_REG_16__SCAN_IN), .B1(n16815), 
        .B2(n16814), .ZN(n16824) );
  AOI211_X1 U19915 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16831), .A(n16816), .B(
        n16997), .ZN(n16817) );
  AOI211_X1 U19916 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n16940), .A(
        n18252), .B(n16817), .ZN(n16823) );
  INV_X1 U19917 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17762) );
  INV_X1 U19918 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17768) );
  INV_X1 U19919 ( .A(n16919), .ZN(n17844) );
  NAND2_X1 U19920 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17844), .ZN(
        n16950) );
  NOR2_X1 U19921 ( .A1(n17828), .A2(n16950), .ZN(n16876) );
  NAND2_X1 U19922 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16876), .ZN(
        n17781) );
  OR2_X1 U19923 ( .A1(n17784), .A2(n17781), .ZN(n16849) );
  NOR2_X1 U19924 ( .A1(n17768), .A2(n16849), .ZN(n17740) );
  INV_X1 U19925 ( .A(n17740), .ZN(n16826) );
  NOR2_X1 U19926 ( .A1(n17762), .A2(n16826), .ZN(n16825) );
  OAI21_X1 U19927 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16825), .A(
        n16818), .ZN(n17746) );
  NOR2_X1 U19928 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17933), .ZN(
        n17007) );
  NAND3_X1 U19929 ( .A1(n9779), .A2(n16819), .A3(n17007), .ZN(n16828) );
  OAI21_X1 U19930 ( .B1(n17762), .B2(n16828), .A(n16641), .ZN(n16827) );
  AOI21_X1 U19931 ( .B1(n17746), .B2(n16827), .A(n17016), .ZN(n16820) );
  OAI21_X1 U19932 ( .B1(n17746), .B2(n16827), .A(n16820), .ZN(n16822) );
  AOI21_X1 U19933 ( .B1(n16841), .B2(n16983), .A(n16999), .ZN(n16834) );
  INV_X1 U19934 ( .A(n16834), .ZN(n16845) );
  NOR3_X1 U19935 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n17018), .A3(n16841), 
        .ZN(n16836) );
  OAI21_X1 U19936 ( .B1(n16845), .B2(n16836), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n16821) );
  NAND4_X1 U19937 ( .A1(n16824), .A2(n16823), .A3(n16822), .A4(n16821), .ZN(
        P3_U2655) );
  AOI21_X1 U19938 ( .B1(n17762), .B2(n16826), .A(n16825), .ZN(n17752) );
  INV_X1 U19939 ( .A(n16827), .ZN(n16830) );
  NAND2_X1 U19940 ( .A1(n16979), .A2(n17006), .ZN(n17010) );
  INV_X1 U19941 ( .A(n17010), .ZN(n16902) );
  AOI21_X1 U19942 ( .B1(n17752), .B2(n16828), .A(n17016), .ZN(n16829) );
  OAI22_X1 U19943 ( .A1(n17752), .A2(n16830), .B1(n16902), .B2(n16829), .ZN(
        n16833) );
  OAI211_X1 U19944 ( .C1(n16840), .C2(n16838), .A(n17025), .B(n16831), .ZN(
        n16832) );
  OAI211_X1 U19945 ( .C1(n16834), .C2(n18833), .A(n16833), .B(n16832), .ZN(
        n16835) );
  AOI211_X1 U19946 ( .C1(n16940), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16836), .B(n16835), .ZN(n16837) );
  OAI211_X1 U19947 ( .C1(n17017), .C2(n16838), .A(n16837), .B(n18236), .ZN(
        P3_U2656) );
  AOI21_X1 U19948 ( .B1(n17768), .B2(n16849), .A(n17740), .ZN(n17770) );
  AOI21_X1 U19949 ( .B1(n9779), .B2(n17007), .A(n16979), .ZN(n16868) );
  INV_X1 U19950 ( .A(n16868), .ZN(n16866) );
  OAI21_X1 U19951 ( .B1(n16979), .B2(n16839), .A(n16866), .ZN(n16858) );
  XNOR2_X1 U19952 ( .A(n17770), .B(n16858), .ZN(n16848) );
  AOI22_X1 U19953 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16940), .B1(
        n17026), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16847) );
  AOI211_X1 U19954 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16852), .A(n16840), .B(
        n16997), .ZN(n16844) );
  INV_X1 U19955 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18829) );
  NAND3_X1 U19956 ( .A1(n16841), .A2(n16851), .A3(n16983), .ZN(n16842) );
  OAI21_X1 U19957 ( .B1(n18829), .B2(n16842), .A(n18236), .ZN(n16843) );
  AOI211_X1 U19958 ( .C1(n16845), .C2(P3_REIP_REG_14__SCAN_IN), .A(n16844), 
        .B(n16843), .ZN(n16846) );
  OAI211_X1 U19959 ( .C1(n17016), .C2(n16848), .A(n16847), .B(n16846), .ZN(
        P3_U2657) );
  INV_X1 U19960 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16865) );
  NOR2_X1 U19961 ( .A1(n16865), .A2(n17781), .ZN(n16864) );
  OAI21_X1 U19962 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16864), .A(
        n16849), .ZN(n17786) );
  OAI21_X1 U19963 ( .B1(n16979), .B2(n16980), .A(n17006), .ZN(n16944) );
  INV_X1 U19964 ( .A(n16944), .ZN(n17021) );
  OAI21_X1 U19965 ( .B1(n16864), .B2(n16979), .A(n17021), .ZN(n16861) );
  AOI21_X1 U19966 ( .B1(n16983), .B2(n16862), .A(n16999), .ZN(n16879) );
  OAI21_X1 U19967 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17018), .A(n16879), 
        .ZN(n16857) );
  INV_X1 U19968 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16850) );
  OAI22_X1 U19969 ( .A1(n16850), .A2(n17014), .B1(n17017), .B2(n17215), .ZN(
        n16856) );
  NAND2_X1 U19970 ( .A1(n16983), .A2(n16851), .ZN(n16854) );
  OAI211_X1 U19971 ( .C1(n16869), .C2(n17215), .A(n17025), .B(n16852), .ZN(
        n16853) );
  OAI211_X1 U19972 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16854), .A(n18236), 
        .B(n16853), .ZN(n16855) );
  AOI211_X1 U19973 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16857), .A(n16856), 
        .B(n16855), .ZN(n16860) );
  NAND3_X1 U19974 ( .A1(n17006), .A2(n17786), .A3(n16858), .ZN(n16859) );
  OAI211_X1 U19975 ( .C1(n17786), .C2(n16861), .A(n16860), .B(n16859), .ZN(
        P3_U2658) );
  NOR3_X1 U19976 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17018), .A3(n16862), 
        .ZN(n16863) );
  AOI211_X1 U19977 ( .C1(n17026), .C2(P3_EBX_REG_12__SCAN_IN), .A(n18252), .B(
        n16863), .ZN(n16873) );
  AOI21_X1 U19978 ( .B1(n16865), .B2(n17781), .A(n16864), .ZN(n17798) );
  INV_X1 U19979 ( .A(n17798), .ZN(n16867) );
  AOI221_X1 U19980 ( .B1(n17798), .B2(n16868), .C1(n16867), .C2(n16866), .A(
        n17016), .ZN(n16871) );
  AOI211_X1 U19981 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16882), .A(n16869), .B(
        n16997), .ZN(n16870) );
  AOI211_X1 U19982 ( .C1(n16940), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16871), .B(n16870), .ZN(n16872) );
  OAI211_X1 U19983 ( .C1(n16879), .C2(n18827), .A(n16873), .B(n16872), .ZN(
        P3_U2659) );
  INV_X1 U19984 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18823) );
  INV_X1 U19985 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18821) );
  NOR2_X1 U19986 ( .A1(n18823), .A2(n18821), .ZN(n16895) );
  NOR2_X1 U19987 ( .A1(n17018), .A2(n16874), .ZN(n16932) );
  INV_X1 U19988 ( .A(n16932), .ZN(n16941) );
  NOR2_X1 U19989 ( .A1(n16875), .A2(n16941), .ZN(n16909) );
  AOI21_X1 U19990 ( .B1(n16895), .B2(n16909), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16880) );
  OAI21_X1 U19991 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16876), .A(
        n17781), .ZN(n17819) );
  INV_X1 U19992 ( .A(n16876), .ZN(n16890) );
  OAI21_X1 U19993 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16890), .A(
        n16641), .ZN(n16877) );
  XNOR2_X1 U19994 ( .A(n17819), .B(n16877), .ZN(n16878) );
  OAI22_X1 U19995 ( .A1(n16880), .A2(n16879), .B1(n17016), .B2(n16878), .ZN(
        n16881) );
  AOI211_X1 U19996 ( .C1(n17026), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18252), .B(
        n16881), .ZN(n16885) );
  OAI211_X1 U19997 ( .C1(n16886), .C2(n16883), .A(n17025), .B(n16882), .ZN(
        n16884) );
  OAI211_X1 U19998 ( .C1(n17014), .C2(n17808), .A(n16885), .B(n16884), .ZN(
        P3_U2660) );
  INV_X1 U19999 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17820) );
  AOI211_X1 U20000 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16887), .A(n16886), .B(
        n16997), .ZN(n16888) );
  AOI211_X1 U20001 ( .C1(n17026), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18252), .B(
        n16888), .ZN(n16899) );
  OAI21_X1 U20002 ( .B1(n16889), .B2(n17018), .A(n17027), .ZN(n16921) );
  INV_X1 U20003 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16901) );
  INV_X1 U20004 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17862) );
  NOR2_X1 U20005 ( .A1(n17862), .A2(n16950), .ZN(n16928) );
  NAND2_X1 U20006 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16928), .ZN(
        n16917) );
  NOR2_X1 U20007 ( .A1(n16901), .A2(n16917), .ZN(n16891) );
  OAI21_X1 U20008 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16891), .A(
        n16890), .ZN(n17831) );
  INV_X1 U20009 ( .A(n17831), .ZN(n16893) );
  NOR2_X1 U20010 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16917), .ZN(
        n16906) );
  AOI21_X1 U20011 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16906), .A(
        n16979), .ZN(n16905) );
  INV_X1 U20012 ( .A(n16905), .ZN(n16892) );
  AOI221_X1 U20013 ( .B1(n16893), .B2(n16905), .C1(n17831), .C2(n16892), .A(
        n17016), .ZN(n16897) );
  INV_X1 U20014 ( .A(n16909), .ZN(n16894) );
  AOI211_X1 U20015 ( .C1(n18823), .C2(n18821), .A(n16895), .B(n16894), .ZN(
        n16896) );
  AOI211_X1 U20016 ( .C1(n16921), .C2(P3_REIP_REG_10__SCAN_IN), .A(n16897), 
        .B(n16896), .ZN(n16898) );
  OAI211_X1 U20017 ( .C1(n17820), .C2(n17014), .A(n16899), .B(n16898), .ZN(
        P3_U2661) );
  AOI21_X1 U20018 ( .B1(n17025), .B2(n16903), .A(n17026), .ZN(n16913) );
  INV_X1 U20019 ( .A(n16917), .ZN(n16900) );
  OAI22_X1 U20020 ( .A1(n16901), .A2(n16900), .B1(n16917), .B2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16904) );
  AOI22_X1 U20021 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16940), .B1(
        n16904), .B2(n16902), .ZN(n16911) );
  OR2_X1 U20022 ( .A1(n16997), .A2(n16903), .ZN(n16915) );
  INV_X1 U20023 ( .A(n16904), .ZN(n17839) );
  OAI211_X1 U20024 ( .C1(n16906), .C2(n17839), .A(n17006), .B(n16905), .ZN(
        n16907) );
  OAI211_X1 U20025 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16915), .A(n18236), .B(
        n16907), .ZN(n16908) );
  AOI221_X1 U20026 ( .B1(n16921), .B2(P3_REIP_REG_9__SCAN_IN), .C1(n16909), 
        .C2(n18821), .A(n16908), .ZN(n16910) );
  OAI211_X1 U20027 ( .C1(n16913), .C2(n16912), .A(n16911), .B(n16910), .ZN(
        P3_U2662) );
  INV_X1 U20028 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18818) );
  INV_X1 U20029 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18816) );
  NOR4_X1 U20030 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18818), .A3(n18816), .A4(
        n16941), .ZN(n16914) );
  AOI21_X1 U20031 ( .B1(n16940), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16914), .ZN(n16925) );
  AOI21_X1 U20032 ( .B1(n16936), .B2(P3_EBX_REG_8__SCAN_IN), .A(n16915), .ZN(
        n16916) );
  AOI21_X1 U20033 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17026), .A(n16916), .ZN(
        n16924) );
  OAI21_X1 U20034 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16928), .A(
        n16917), .ZN(n16918) );
  INV_X1 U20035 ( .A(n16918), .ZN(n17845) );
  NOR2_X1 U20036 ( .A1(n16919), .A2(n17862), .ZN(n17854) );
  AOI21_X1 U20037 ( .B1(n17854), .B2(n17007), .A(n16979), .ZN(n16920) );
  XOR2_X1 U20038 ( .A(n17845), .B(n16920), .Z(n16922) );
  AOI22_X1 U20039 ( .A1(n17006), .A2(n16922), .B1(P3_REIP_REG_8__SCAN_IN), 
        .B2(n16921), .ZN(n16923) );
  NAND4_X1 U20040 ( .A1(n16925), .A2(n16924), .A3(n16923), .A4(n18236), .ZN(
        P3_U2663) );
  NAND2_X1 U20041 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n16927) );
  NAND2_X1 U20042 ( .A1(n16926), .A2(n17027), .ZN(n16963) );
  OAI21_X1 U20043 ( .B1(n16927), .B2(n16963), .A(n17024), .ZN(n16957) );
  OAI21_X1 U20044 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16941), .A(n16957), .ZN(
        n16948) );
  AOI21_X1 U20045 ( .B1(n17862), .B2(n16950), .A(n16928), .ZN(n17867) );
  OAI21_X1 U20046 ( .B1(n16950), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16641), .ZN(n16929) );
  INV_X1 U20047 ( .A(n16929), .ZN(n16931) );
  OAI21_X1 U20048 ( .B1(n17867), .B2(n16931), .A(n17006), .ZN(n16930) );
  AOI21_X1 U20049 ( .B1(n17867), .B2(n16931), .A(n16930), .ZN(n16935) );
  NAND3_X1 U20050 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16932), .A3(n18818), 
        .ZN(n16933) );
  OAI211_X1 U20051 ( .C1(n17862), .C2(n17014), .A(n18236), .B(n16933), .ZN(
        n16934) );
  AOI211_X1 U20052 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n16948), .A(n16935), .B(
        n16934), .ZN(n16938) );
  OAI211_X1 U20053 ( .C1(n16942), .C2(n16939), .A(n17025), .B(n16936), .ZN(
        n16937) );
  OAI211_X1 U20054 ( .C1(n16939), .C2(n17017), .A(n16938), .B(n16937), .ZN(
        P3_U2664) );
  AOI22_X1 U20055 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16940), .B1(
        n17026), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n16953) );
  NAND2_X1 U20056 ( .A1(n18816), .A2(n16941), .ZN(n16947) );
  AOI211_X1 U20057 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16960), .A(n16942), .B(
        n16997), .ZN(n16946) );
  NAND2_X1 U20058 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17878), .ZN(
        n16955) );
  INV_X1 U20059 ( .A(n16955), .ZN(n16943) );
  OAI21_X1 U20060 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16943), .A(
        n16950), .ZN(n17881) );
  AOI211_X1 U20061 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16641), .A(
        n17881), .B(n16944), .ZN(n16945) );
  AOI211_X1 U20062 ( .C1(n16948), .C2(n16947), .A(n16946), .B(n16945), .ZN(
        n16952) );
  NOR2_X1 U20063 ( .A1(n16979), .A2(n17016), .ZN(n16949) );
  OAI211_X1 U20064 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n16950), .A(
        n16949), .B(n17881), .ZN(n16951) );
  NAND4_X1 U20065 ( .A1(n16953), .A2(n16952), .A3(n18236), .A4(n16951), .ZN(
        P3_U2665) );
  INV_X1 U20066 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18812) );
  NAND3_X1 U20067 ( .A1(n16983), .A2(P3_REIP_REG_3__SCAN_IN), .A3(n16996), 
        .ZN(n16978) );
  INV_X1 U20068 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18815) );
  OAI21_X1 U20069 ( .B1(n18812), .B2(n16978), .A(n18815), .ZN(n16954) );
  INV_X1 U20070 ( .A(n16954), .ZN(n16958) );
  NOR2_X1 U20071 ( .A1(n17933), .A2(n17888), .ZN(n16967) );
  OAI21_X1 U20072 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16967), .A(
        n16955), .ZN(n17893) );
  AOI21_X1 U20073 ( .B1(n16980), .B2(n16967), .A(n16979), .ZN(n16970) );
  XOR2_X1 U20074 ( .A(n17893), .B(n16970), .Z(n16956) );
  OAI22_X1 U20075 ( .A1(n16958), .A2(n16957), .B1(n17016), .B2(n16956), .ZN(
        n16959) );
  AOI211_X1 U20076 ( .C1(n17026), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18252), .B(
        n16959), .ZN(n16962) );
  OAI211_X1 U20077 ( .C1(n16964), .C2(n17283), .A(n17025), .B(n16960), .ZN(
        n16961) );
  OAI211_X1 U20078 ( .C1(n17014), .C2(n17887), .A(n16962), .B(n16961), .ZN(
        P3_U2666) );
  NAND2_X1 U20079 ( .A1(n17024), .A2(n16963), .ZN(n16984) );
  AOI211_X1 U20080 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16990), .A(n16964), .B(
        n16997), .ZN(n16976) );
  NOR2_X1 U20081 ( .A1(n9888), .A2(n18944), .ZN(n18947) );
  AOI221_X1 U20082 ( .B1(n18947), .B2(n17247), .C1(n18947), .C2(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n18252), .ZN(n16965) );
  INV_X1 U20083 ( .A(n16965), .ZN(n16975) );
  INV_X1 U20084 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16969) );
  NAND2_X1 U20085 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16966), .ZN(
        n16981) );
  AOI21_X1 U20086 ( .B1(n16969), .B2(n16981), .A(n16967), .ZN(n16968) );
  INV_X1 U20087 ( .A(n16968), .ZN(n17901) );
  OAI22_X1 U20088 ( .A1(n16969), .A2(n17014), .B1(n17901), .B2(n17010), .ZN(
        n16974) );
  NAND2_X1 U20089 ( .A1(n16966), .A2(n16969), .ZN(n17905) );
  INV_X1 U20090 ( .A(n17905), .ZN(n16971) );
  AOI22_X1 U20091 ( .A1(n17007), .A2(n16971), .B1(n16970), .B2(n17901), .ZN(
        n16972) );
  OAI22_X1 U20092 ( .A1(n16972), .A2(n17016), .B1(n17017), .B2(n17291), .ZN(
        n16973) );
  NOR4_X1 U20093 ( .A1(n16976), .A2(n16975), .A3(n16974), .A4(n16973), .ZN(
        n16977) );
  OAI221_X1 U20094 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16978), .C1(n18812), 
        .C2(n16984), .A(n16977), .ZN(P3_U2667) );
  NAND2_X1 U20095 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16995) );
  INV_X1 U20096 ( .A(n16995), .ZN(n16982) );
  AOI21_X1 U20097 ( .B1(n16982), .B2(n16980), .A(n16979), .ZN(n17005) );
  OAI21_X1 U20098 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16982), .A(
        n16981), .ZN(n17916) );
  XNOR2_X1 U20099 ( .A(n17005), .B(n17916), .ZN(n16989) );
  INV_X1 U20100 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n21123) );
  NAND2_X1 U20101 ( .A1(n16983), .A2(n16996), .ZN(n16985) );
  AOI21_X1 U20102 ( .B1(n21123), .B2(n16985), .A(n16984), .ZN(n16988) );
  NOR2_X1 U20103 ( .A1(n18909), .A2(n18731), .ZN(n18728) );
  OAI21_X1 U20104 ( .B1(n18728), .B2(n18883), .A(n10230), .ZN(n18881) );
  AOI22_X1 U20105 ( .A1(n18881), .A2(n18947), .B1(n17026), .B2(
        P3_EBX_REG_3__SCAN_IN), .ZN(n16986) );
  INV_X1 U20106 ( .A(n16986), .ZN(n16987) );
  AOI211_X1 U20107 ( .C1(n16989), .C2(n17006), .A(n16988), .B(n16987), .ZN(
        n16993) );
  OAI211_X1 U20108 ( .C1(n16998), .C2(n16991), .A(n17025), .B(n16990), .ZN(
        n16992) );
  OAI211_X1 U20109 ( .C1(n17014), .C2(n16994), .A(n16993), .B(n16992), .ZN(
        P3_U2668) );
  OAI21_X1 U20110 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16995), .ZN(n17923) );
  AOI211_X1 U20111 ( .C1(n18911), .C2(n18809), .A(n16996), .B(n17018), .ZN(
        n17004) );
  INV_X1 U20112 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17307) );
  INV_X1 U20113 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17313) );
  NAND2_X1 U20114 ( .A1(n17307), .A2(n17313), .ZN(n17011) );
  AOI211_X1 U20115 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17011), .A(n16998), .B(
        n16997), .ZN(n17003) );
  INV_X1 U20116 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17297) );
  OAI22_X1 U20117 ( .A1(n17927), .A2(n17014), .B1(n17017), .B2(n17297), .ZN(
        n17002) );
  AOI21_X1 U20118 ( .B1(n18891), .B2(n18739), .A(n18728), .ZN(n18888) );
  AOI22_X1 U20119 ( .A1(n16999), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18888), 
        .B2(n18947), .ZN(n17000) );
  INV_X1 U20120 ( .A(n17000), .ZN(n17001) );
  NOR4_X1 U20121 ( .A1(n17004), .A2(n17003), .A3(n17002), .A4(n17001), .ZN(
        n17009) );
  OAI211_X1 U20122 ( .C1(n17007), .C2(n17923), .A(n17006), .B(n17005), .ZN(
        n17008) );
  OAI211_X1 U20123 ( .C1(n17010), .C2(n17923), .A(n17009), .B(n17008), .ZN(
        P3_U2669) );
  NAND2_X1 U20124 ( .A1(n17011), .A2(n17296), .ZN(n17309) );
  INV_X1 U20125 ( .A(n17309), .ZN(n17013) );
  AND2_X1 U20126 ( .A1(n18739), .A2(n17012), .ZN(n18896) );
  AOI22_X1 U20127 ( .A1(n17025), .A2(n17013), .B1(n18896), .B2(n18947), .ZN(
        n17023) );
  NAND2_X1 U20128 ( .A1(n16641), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17015) );
  OAI21_X1 U20129 ( .B1(n17016), .B2(n17015), .A(n17014), .ZN(n17020) );
  OAI22_X1 U20130 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17018), .B1(n17017), 
        .B2(n17307), .ZN(n17019) );
  AOI221_X1 U20131 ( .B1(n17021), .B2(n17933), .C1(n17020), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17019), .ZN(n17022) );
  OAI211_X1 U20132 ( .C1(n17027), .C2(n18911), .A(n17023), .B(n17022), .ZN(
        P3_U2670) );
  AOI22_X1 U20133 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17024), .B1(n18947), 
        .B2(n18909), .ZN(n17030) );
  OAI21_X1 U20134 ( .B1(n17026), .B2(n17025), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17029) );
  NAND3_X1 U20135 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18904), .A3(
        n17027), .ZN(n17028) );
  NAND3_X1 U20136 ( .A1(n17030), .A2(n17029), .A3(n17028), .ZN(P3_U2671) );
  AOI22_X1 U20137 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20138 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20139 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U20140 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17031) );
  NAND4_X1 U20141 ( .A1(n17034), .A2(n17033), .A3(n17032), .A4(n17031), .ZN(
        n17041) );
  AOI22_X1 U20142 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20143 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20144 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20145 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17036) );
  NAND4_X1 U20146 ( .A1(n17039), .A2(n17038), .A3(n17037), .A4(n17036), .ZN(
        n17040) );
  NOR2_X1 U20147 ( .A1(n17041), .A2(n17040), .ZN(n17060) );
  NOR2_X1 U20148 ( .A1(n17060), .A2(n17059), .ZN(n17058) );
  AOI22_X1 U20149 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20150 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20151 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20152 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17042) );
  NAND4_X1 U20153 ( .A1(n17045), .A2(n17044), .A3(n17043), .A4(n17042), .ZN(
        n17052) );
  AOI22_X1 U20154 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17050) );
  AOI22_X1 U20155 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20156 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9649), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20157 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17047) );
  NAND4_X1 U20158 ( .A1(n17050), .A2(n17049), .A3(n17048), .A4(n17047), .ZN(
        n17051) );
  NOR2_X1 U20159 ( .A1(n17052), .A2(n17051), .ZN(n17053) );
  XOR2_X1 U20160 ( .A(n17058), .B(n17053), .Z(n17324) );
  NOR2_X1 U20161 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17054), .ZN(n17056) );
  OAI22_X1 U20162 ( .A1(n17324), .A2(n17305), .B1(n17056), .B2(n17055), .ZN(
        P3_U2673) );
  NAND2_X1 U20163 ( .A1(n17117), .A2(n17057), .ZN(n17063) );
  AOI21_X1 U20164 ( .B1(n17060), .B2(n17059), .A(n17058), .ZN(n17325) );
  AOI22_X1 U20165 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17061), .B1(n17325), 
        .B2(n17311), .ZN(n17062) );
  OAI21_X1 U20166 ( .B1(n17064), .B2(n17063), .A(n17062), .ZN(P3_U2674) );
  AOI21_X1 U20167 ( .B1(n17066), .B2(n17071), .A(n17065), .ZN(n17334) );
  NAND2_X1 U20168 ( .A1(n17334), .A2(n17311), .ZN(n17067) );
  OAI221_X1 U20169 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17070), .C1(n17069), 
        .C2(n17068), .A(n17067), .ZN(P3_U2676) );
  INV_X1 U20170 ( .A(n17070), .ZN(n17074) );
  AOI21_X1 U20171 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17305), .A(n17080), .ZN(
        n17073) );
  OAI21_X1 U20172 ( .B1(n17076), .B2(n17072), .A(n17071), .ZN(n17343) );
  OAI22_X1 U20173 ( .A1(n17074), .A2(n17073), .B1(n17305), .B2(n17343), .ZN(
        P3_U2677) );
  NOR2_X1 U20174 ( .A1(n17075), .A2(n17081), .ZN(n17085) );
  AOI21_X1 U20175 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17305), .A(n17085), .ZN(
        n17079) );
  AOI21_X1 U20176 ( .B1(n17077), .B2(n17082), .A(n17076), .ZN(n17344) );
  INV_X1 U20177 ( .A(n17344), .ZN(n17078) );
  OAI22_X1 U20178 ( .A1(n17080), .A2(n17079), .B1(n17305), .B2(n17078), .ZN(
        P3_U2678) );
  INV_X1 U20179 ( .A(n17081), .ZN(n17092) );
  AOI21_X1 U20180 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17305), .A(n17092), .ZN(
        n17084) );
  OAI21_X1 U20181 ( .B1(n17087), .B2(n17083), .A(n17082), .ZN(n17353) );
  OAI22_X1 U20182 ( .A1(n17085), .A2(n17084), .B1(n17305), .B2(n17353), .ZN(
        P3_U2679) );
  AOI21_X1 U20183 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17305), .A(n17086), .ZN(
        n17091) );
  AOI21_X1 U20184 ( .B1(n17089), .B2(n17088), .A(n17087), .ZN(n17354) );
  INV_X1 U20185 ( .A(n17354), .ZN(n17090) );
  OAI22_X1 U20186 ( .A1(n17092), .A2(n17091), .B1(n17305), .B2(n17090), .ZN(
        P3_U2680) );
  AOI22_X1 U20187 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20188 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U20189 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U20190 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17093) );
  NAND4_X1 U20191 ( .A1(n17096), .A2(n17095), .A3(n17094), .A4(n17093), .ZN(
        n17102) );
  AOI22_X1 U20192 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9650), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20193 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20194 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20195 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17097) );
  NAND4_X1 U20196 ( .A1(n17100), .A2(n17099), .A3(n17098), .A4(n17097), .ZN(
        n17101) );
  NOR2_X1 U20197 ( .A1(n17102), .A2(n17101), .ZN(n17362) );
  NAND3_X1 U20198 ( .A1(n17104), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17305), 
        .ZN(n17103) );
  OAI221_X1 U20199 ( .B1(n17104), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17305), 
        .C2(n17362), .A(n17103), .ZN(P3_U2681) );
  AOI22_X1 U20200 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17108) );
  AOI22_X1 U20201 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17107) );
  AOI22_X1 U20202 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20203 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17105) );
  NAND4_X1 U20204 ( .A1(n17108), .A2(n17107), .A3(n17106), .A4(n17105), .ZN(
        n17114) );
  AOI22_X1 U20205 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20206 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20207 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20208 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17109) );
  NAND4_X1 U20209 ( .A1(n17112), .A2(n17111), .A3(n17110), .A4(n17109), .ZN(
        n17113) );
  NOR2_X1 U20210 ( .A1(n17114), .A2(n17113), .ZN(n17368) );
  AND2_X1 U20211 ( .A1(n17305), .A2(n17115), .ZN(n17130) );
  AOI22_X1 U20212 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17130), .B1(n17117), 
        .B2(n17116), .ZN(n17118) );
  OAI21_X1 U20213 ( .B1(n17368), .B2(n17305), .A(n17118), .ZN(P3_U2682) );
  AOI22_X1 U20214 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9645), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20215 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17121) );
  AOI22_X1 U20216 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12816), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U20217 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17119) );
  NAND4_X1 U20218 ( .A1(n17122), .A2(n17121), .A3(n17120), .A4(n17119), .ZN(
        n17128) );
  AOI22_X1 U20219 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20220 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17125) );
  AOI22_X1 U20221 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U20222 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9657), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17123) );
  NAND4_X1 U20223 ( .A1(n17126), .A2(n17125), .A3(n17124), .A4(n17123), .ZN(
        n17127) );
  NOR2_X1 U20224 ( .A1(n17128), .A2(n17127), .ZN(n17376) );
  INV_X1 U20225 ( .A(n17129), .ZN(n17131) );
  OAI21_X1 U20226 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17131), .A(n17130), .ZN(
        n17132) );
  OAI21_X1 U20227 ( .B1(n17376), .B2(n17305), .A(n17132), .ZN(P3_U2683) );
  AOI21_X1 U20228 ( .B1(n17134), .B2(n17133), .A(n17311), .ZN(n17135) );
  INV_X1 U20229 ( .A(n17135), .ZN(n17146) );
  AOI22_X1 U20230 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U20231 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20232 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20233 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17136) );
  NAND4_X1 U20234 ( .A1(n17139), .A2(n17138), .A3(n17137), .A4(n17136), .ZN(
        n17145) );
  AOI22_X1 U20235 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20236 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20237 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20238 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17140) );
  NAND4_X1 U20239 ( .A1(n17143), .A2(n17142), .A3(n17141), .A4(n17140), .ZN(
        n17144) );
  NOR2_X1 U20240 ( .A1(n17145), .A2(n17144), .ZN(n17380) );
  OAI22_X1 U20241 ( .A1(n17147), .A2(n17146), .B1(n17380), .B2(n17305), .ZN(
        P3_U2684) );
  NOR2_X1 U20242 ( .A1(n17404), .A2(n17148), .ZN(n17261) );
  NAND4_X1 U20243 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n17149), .A4(n17261), .ZN(n17163) );
  NOR2_X1 U20244 ( .A1(n17311), .A2(n17150), .ZN(n17175) );
  AOI22_X1 U20245 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9648), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20246 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20247 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17151) );
  OAI21_X1 U20248 ( .B1(n12827), .B2(n17152), .A(n17151), .ZN(n17158) );
  AOI22_X1 U20249 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17156) );
  AOI22_X1 U20250 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12839), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20251 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20252 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12752), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17153) );
  NAND4_X1 U20253 ( .A1(n17156), .A2(n17155), .A3(n17154), .A4(n17153), .ZN(
        n17157) );
  AOI211_X1 U20254 ( .C1(n17247), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17158), .B(n17157), .ZN(n17159) );
  NAND3_X1 U20255 ( .A1(n17161), .A2(n17160), .A3(n17159), .ZN(n17381) );
  AOI22_X1 U20256 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17175), .B1(n17311), 
        .B2(n17381), .ZN(n17162) );
  OAI21_X1 U20257 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17163), .A(n17162), .ZN(
        P3_U2685) );
  AOI22_X1 U20258 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17190), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17167) );
  AOI22_X1 U20259 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9648), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20260 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17270), .ZN(n17165) );
  AOI22_X1 U20261 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17252), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12752), .ZN(n17164) );
  NAND4_X1 U20262 ( .A1(n17167), .A2(n17166), .A3(n17165), .A4(n17164), .ZN(
        n17173) );
  AOI22_X1 U20263 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17171) );
  AOI22_X1 U20264 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n15814), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17170) );
  AOI22_X1 U20265 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n12839), .ZN(n17169) );
  AOI22_X1 U20266 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n9645), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17168) );
  NAND4_X1 U20267 ( .A1(n17171), .A2(n17170), .A3(n17169), .A4(n17168), .ZN(
        n17172) );
  NOR2_X1 U20268 ( .A1(n17173), .A2(n17172), .ZN(n17392) );
  INV_X1 U20269 ( .A(n17174), .ZN(n17176) );
  OAI21_X1 U20270 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17176), .A(n17175), .ZN(
        n17177) );
  OAI21_X1 U20271 ( .B1(n17392), .B2(n17305), .A(n17177), .ZN(P3_U2686) );
  INV_X1 U20272 ( .A(n17232), .ZN(n17178) );
  NOR2_X1 U20273 ( .A1(n17201), .A2(n17178), .ZN(n17218) );
  NAND3_X1 U20274 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17218), .ZN(n17202) );
  AOI22_X1 U20275 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17182) );
  AOI22_X1 U20276 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U20277 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20278 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12752), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17179) );
  NAND4_X1 U20279 ( .A1(n17182), .A2(n17181), .A3(n17180), .A4(n17179), .ZN(
        n17188) );
  AOI22_X1 U20280 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12816), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17186) );
  AOI22_X1 U20281 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12839), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20282 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20283 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17183) );
  NAND4_X1 U20284 ( .A1(n17186), .A2(n17185), .A3(n17184), .A4(n17183), .ZN(
        n17187) );
  NOR2_X1 U20285 ( .A1(n17188), .A2(n17187), .ZN(n17398) );
  NAND3_X1 U20286 ( .A1(n17202), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17305), 
        .ZN(n17189) );
  OAI221_X1 U20287 ( .B1(n17202), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n17305), 
        .C2(n17398), .A(n17189), .ZN(P3_U2687) );
  AOI22_X1 U20288 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20289 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12816), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20290 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12752), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20291 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17191) );
  NAND4_X1 U20292 ( .A1(n17194), .A2(n17193), .A3(n17192), .A4(n17191), .ZN(
        n17200) );
  AOI22_X1 U20293 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12839), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U20294 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9644), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20295 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U20296 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17195) );
  NAND4_X1 U20297 ( .A1(n17198), .A2(n17197), .A3(n17196), .A4(n17195), .ZN(
        n17199) );
  NOR2_X1 U20298 ( .A1(n17200), .A2(n17199), .ZN(n17402) );
  NOR3_X1 U20299 ( .A1(n17217), .A2(n17201), .A3(n17244), .ZN(n17203) );
  OAI211_X1 U20300 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17203), .A(n17202), .B(
        n17305), .ZN(n17204) );
  OAI21_X1 U20301 ( .B1(n17402), .B2(n17305), .A(n17204), .ZN(P3_U2688) );
  AOI22_X1 U20302 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20303 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17207) );
  AOI22_X1 U20304 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12839), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U20305 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12752), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17205) );
  NAND4_X1 U20306 ( .A1(n17208), .A2(n17207), .A3(n17206), .A4(n17205), .ZN(
        n17214) );
  AOI22_X1 U20307 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20308 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20309 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9648), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20310 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17209) );
  NAND4_X1 U20311 ( .A1(n17212), .A2(n17211), .A3(n17210), .A4(n17209), .ZN(
        n17213) );
  NOR2_X1 U20312 ( .A1(n17214), .A2(n17213), .ZN(n17406) );
  INV_X1 U20313 ( .A(n17308), .ZN(n17310) );
  AOI21_X1 U20314 ( .B1(n17215), .B2(n17310), .A(n17231), .ZN(n17216) );
  INV_X1 U20315 ( .A(n17216), .ZN(n17219) );
  AOI22_X1 U20316 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17219), .B1(n17218), 
        .B2(n17217), .ZN(n17220) );
  OAI21_X1 U20317 ( .B1(n17406), .B2(n17305), .A(n17220), .ZN(P3_U2689) );
  AOI22_X1 U20318 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20319 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20320 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20321 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12752), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17221) );
  NAND4_X1 U20322 ( .A1(n17224), .A2(n17223), .A3(n17222), .A4(n17221), .ZN(
        n17230) );
  AOI22_X1 U20323 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20324 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12839), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20325 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9644), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20326 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17225) );
  NAND4_X1 U20327 ( .A1(n17228), .A2(n17227), .A3(n17226), .A4(n17225), .ZN(
        n17229) );
  NOR2_X1 U20328 ( .A1(n17230), .A2(n17229), .ZN(n17415) );
  OAI21_X1 U20329 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17232), .A(n17231), .ZN(
        n17233) );
  OAI21_X1 U20330 ( .B1(n17415), .B2(n17305), .A(n17233), .ZN(P3_U2691) );
  AOI22_X1 U20331 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20332 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20333 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U20334 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12752), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17234) );
  NAND4_X1 U20335 ( .A1(n17237), .A2(n17236), .A3(n17235), .A4(n17234), .ZN(
        n17243) );
  AOI22_X1 U20336 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9650), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20337 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17263), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U20338 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U20339 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12839), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17238) );
  NAND4_X1 U20340 ( .A1(n17241), .A2(n17240), .A3(n17239), .A4(n17238), .ZN(
        n17242) );
  NOR2_X1 U20341 ( .A1(n17243), .A2(n17242), .ZN(n17419) );
  OAI21_X1 U20342 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17245), .A(n17244), .ZN(
        n17246) );
  AOI22_X1 U20343 ( .A1(n17311), .A2(n17419), .B1(n17246), .B2(n17305), .ZN(
        P3_U2692) );
  AOI22_X1 U20344 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17247), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U20345 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17263), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U20346 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12838), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17249) );
  AOI22_X1 U20347 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12752), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17248) );
  NAND4_X1 U20348 ( .A1(n17251), .A2(n17250), .A3(n17249), .A4(n17248), .ZN(
        n17258) );
  AOI22_X1 U20349 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17262), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U20350 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n12839), .ZN(n17255) );
  AOI22_X1 U20351 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n9645), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9648), .ZN(n17254) );
  AOI22_X1 U20352 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9642), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17252), .ZN(n17253) );
  NAND4_X1 U20353 ( .A1(n17256), .A2(n17255), .A3(n17254), .A4(n17253), .ZN(
        n17257) );
  NOR2_X1 U20354 ( .A1(n17258), .A2(n17257), .ZN(n17430) );
  OAI21_X1 U20355 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17278), .A(n17259), .ZN(
        n17260) );
  OAI21_X1 U20356 ( .B1(n17430), .B2(n17305), .A(n17260), .ZN(P3_U2694) );
  OAI21_X1 U20357 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17261), .A(n17305), .ZN(
        n17277) );
  AOI22_X1 U20358 ( .A1(n15834), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U20359 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17267) );
  AOI22_X1 U20360 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15804), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17266) );
  AOI22_X1 U20361 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17264), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17265) );
  NAND4_X1 U20362 ( .A1(n17268), .A2(n17267), .A3(n17266), .A4(n17265), .ZN(
        n17276) );
  AOI22_X1 U20363 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15814), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U20364 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9645), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U20365 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17272) );
  AOI22_X1 U20366 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9649), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17271) );
  NAND4_X1 U20367 ( .A1(n17274), .A2(n17273), .A3(n17272), .A4(n17271), .ZN(
        n17275) );
  NOR2_X1 U20368 ( .A1(n17276), .A2(n17275), .ZN(n17438) );
  OAI22_X1 U20369 ( .A1(n17278), .A2(n17277), .B1(n17438), .B2(n17305), .ZN(
        P3_U2695) );
  NAND2_X1 U20370 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n17279) );
  NOR4_X1 U20371 ( .A1(n17404), .A2(n17291), .A3(n17295), .A4(n17279), .ZN(
        n17286) );
  AOI21_X1 U20372 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17305), .A(n17286), .ZN(
        n17281) );
  OAI22_X1 U20373 ( .A1(n17282), .A2(n17281), .B1(n17280), .B2(n17305), .ZN(
        P3_U2696) );
  NOR4_X1 U20374 ( .A1(n17404), .A2(n17283), .A3(n17291), .A4(n17295), .ZN(
        n17289) );
  AOI21_X1 U20375 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17305), .A(n17289), .ZN(
        n17285) );
  INV_X1 U20376 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17284) );
  OAI22_X1 U20377 ( .A1(n17286), .A2(n17285), .B1(n17284), .B2(n17305), .ZN(
        P3_U2697) );
  OAI21_X1 U20378 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17290), .A(n17305), .ZN(
        n17288) );
  INV_X1 U20379 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17287) );
  OAI22_X1 U20380 ( .A1(n17289), .A2(n17288), .B1(n17287), .B2(n17305), .ZN(
        P3_U2698) );
  INV_X1 U20381 ( .A(n17290), .ZN(n17293) );
  AOI21_X1 U20382 ( .B1(n17291), .B2(n17295), .A(n17311), .ZN(n17292) );
  AOI22_X1 U20383 ( .A1(n17293), .A2(n17292), .B1(
        P3_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n17311), .ZN(n17294) );
  INV_X1 U20384 ( .A(n17294), .ZN(P3_U2699) );
  INV_X1 U20385 ( .A(n17295), .ZN(n17300) );
  NOR3_X1 U20386 ( .A1(n17297), .A2(n17296), .A3(n17308), .ZN(n17304) );
  AOI21_X1 U20387 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17305), .A(n17304), .ZN(
        n17299) );
  INV_X1 U20388 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17298) );
  OAI22_X1 U20389 ( .A1(n17300), .A2(n17299), .B1(n17298), .B2(n17305), .ZN(
        P3_U2700) );
  AOI22_X1 U20390 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17305), .B1(n17301), .B2(
        n17310), .ZN(n17303) );
  INV_X1 U20391 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17302) );
  OAI22_X1 U20392 ( .A1(n17304), .A2(n17303), .B1(n17302), .B2(n17305), .ZN(
        P3_U2701) );
  OAI222_X1 U20393 ( .A1(n17309), .A2(n17308), .B1(n17307), .B2(n17314), .C1(
        n17306), .C2(n17305), .ZN(P3_U2702) );
  AOI22_X1 U20394 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17311), .B1(
        n17310), .B2(n17313), .ZN(n17312) );
  OAI21_X1 U20395 ( .B1(n17314), .B2(n17313), .A(n17312), .ZN(P3_U2703) );
  INV_X1 U20396 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17537) );
  INV_X1 U20397 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17533) );
  INV_X1 U20398 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17577) );
  INV_X1 U20399 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21109) );
  NAND3_X1 U20400 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .ZN(n17440) );
  INV_X1 U20401 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17547) );
  AND4_X1 U20402 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17315)
         );
  NAND2_X1 U20403 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .ZN(n17360) );
  NAND2_X1 U20404 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17350), .ZN(n17349) );
  NAND2_X1 U20405 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17329), .ZN(n17326) );
  NAND2_X1 U20406 ( .A1(n17321), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17320) );
  NAND2_X1 U20407 ( .A1(n17317), .A2(n17435), .ZN(n17367) );
  OAI22_X1 U20408 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17467), .B1(n17435), 
        .B2(n17321), .ZN(n17318) );
  AOI22_X1 U20409 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17393), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17318), .ZN(n17319) );
  OAI21_X1 U20410 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17320), .A(n17319), .ZN(
        P3_U2704) );
  NAND2_X1 U20411 ( .A1(n18297), .A2(n17435), .ZN(n17387) );
  AOI22_X1 U20412 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17394), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17393), .ZN(n17323) );
  OAI211_X1 U20413 ( .C1(n17321), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17458), .B(
        n17320), .ZN(n17322) );
  OAI211_X1 U20414 ( .C1(n17324), .C2(n17460), .A(n17323), .B(n17322), .ZN(
        P3_U2705) );
  AOI22_X1 U20415 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17394), .B1(n17465), .B2(
        n17325), .ZN(n17328) );
  OAI211_X1 U20416 ( .C1(n17329), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17458), .B(
        n17326), .ZN(n17327) );
  OAI211_X1 U20417 ( .C1(n17367), .C2(n15028), .A(n17328), .B(n17327), .ZN(
        P3_U2706) );
  AOI22_X1 U20418 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17394), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17393), .ZN(n17332) );
  AOI211_X1 U20419 ( .C1(n17537), .C2(n17335), .A(n17329), .B(n17435), .ZN(
        n17330) );
  INV_X1 U20420 ( .A(n17330), .ZN(n17331) );
  OAI211_X1 U20421 ( .C1(n17333), .C2(n17460), .A(n17332), .B(n17331), .ZN(
        P3_U2707) );
  INV_X1 U20422 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20423 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17394), .B1(n17465), .B2(
        n17334), .ZN(n17337) );
  OAI211_X1 U20424 ( .C1(n17339), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17458), .B(
        n17335), .ZN(n17336) );
  OAI211_X1 U20425 ( .C1(n17367), .C2(n17338), .A(n17337), .B(n17336), .ZN(
        P3_U2708) );
  AOI22_X1 U20426 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17394), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17393), .ZN(n17342) );
  AOI211_X1 U20427 ( .C1(n17533), .C2(n17345), .A(n17339), .B(n17435), .ZN(
        n17340) );
  INV_X1 U20428 ( .A(n17340), .ZN(n17341) );
  OAI211_X1 U20429 ( .C1(n17343), .C2(n17460), .A(n17342), .B(n17341), .ZN(
        P3_U2709) );
  INV_X1 U20430 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18280) );
  AOI22_X1 U20431 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17394), .B1(n17465), .B2(
        n17344), .ZN(n17348) );
  OAI211_X1 U20432 ( .C1(n17346), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17458), .B(
        n17345), .ZN(n17347) );
  OAI211_X1 U20433 ( .C1(n17367), .C2(n18280), .A(n17348), .B(n17347), .ZN(
        P3_U2710) );
  AOI22_X1 U20434 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17394), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17393), .ZN(n17352) );
  OAI211_X1 U20435 ( .C1(n17350), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17458), .B(
        n17349), .ZN(n17351) );
  OAI211_X1 U20436 ( .C1(n17353), .C2(n17460), .A(n17352), .B(n17351), .ZN(
        P3_U2711) );
  INV_X1 U20437 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U20438 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17394), .B1(n17465), .B2(
        n17354), .ZN(n17358) );
  OAI211_X1 U20439 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17356), .A(n17458), .B(
        n17355), .ZN(n17357) );
  OAI211_X1 U20440 ( .C1(n17367), .C2(n17359), .A(n17358), .B(n17357), .ZN(
        P3_U2712) );
  INV_X1 U20441 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18300) );
  INV_X1 U20442 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17518) );
  INV_X1 U20443 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17516) );
  INV_X1 U20444 ( .A(n17384), .ZN(n17388) );
  NAND2_X1 U20445 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17382), .ZN(n17377) );
  NAND2_X1 U20446 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17373), .ZN(n17372) );
  NAND2_X1 U20447 ( .A1(n17458), .A2(n17372), .ZN(n17371) );
  OAI21_X1 U20448 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17467), .A(n17371), .ZN(
        n17365) );
  NOR3_X1 U20449 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17360), .A3(n17377), .ZN(
        n17364) );
  INV_X1 U20450 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n17361) );
  OAI22_X1 U20451 ( .A1(n17362), .A2(n17460), .B1(n17361), .B2(n17367), .ZN(
        n17363) );
  AOI211_X1 U20452 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17365), .A(n17364), .B(
        n17363), .ZN(n17366) );
  OAI21_X1 U20453 ( .B1(n18300), .B2(n17387), .A(n17366), .ZN(P3_U2713) );
  INV_X1 U20454 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17523) );
  INV_X1 U20455 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19405) );
  OAI22_X1 U20456 ( .A1(n17368), .A2(n17460), .B1(n19405), .B2(n17367), .ZN(
        n17369) );
  AOI21_X1 U20457 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17394), .A(n17369), .ZN(
        n17370) );
  OAI221_X1 U20458 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17372), .C1(n17523), 
        .C2(n17371), .A(n17370), .ZN(P3_U2714) );
  AOI22_X1 U20459 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17394), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17393), .ZN(n17375) );
  OAI211_X1 U20460 ( .C1(n17373), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17458), .B(
        n17372), .ZN(n17374) );
  OAI211_X1 U20461 ( .C1(n17376), .C2(n17460), .A(n17375), .B(n17374), .ZN(
        P3_U2715) );
  AOI22_X1 U20462 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17394), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17393), .ZN(n17379) );
  OAI211_X1 U20463 ( .C1(n17382), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17458), .B(
        n17377), .ZN(n17378) );
  OAI211_X1 U20464 ( .C1(n17380), .C2(n17460), .A(n17379), .B(n17378), .ZN(
        P3_U2716) );
  INV_X1 U20465 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18284) );
  AOI22_X1 U20466 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17393), .B1(n17465), .B2(
        n17381), .ZN(n17386) );
  INV_X1 U20467 ( .A(n17382), .ZN(n17383) );
  OAI211_X1 U20468 ( .C1(n17384), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17458), .B(
        n17383), .ZN(n17385) );
  OAI211_X1 U20469 ( .C1(n17387), .C2(n18284), .A(n17386), .B(n17385), .ZN(
        P3_U2717) );
  AOI22_X1 U20470 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17394), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17393), .ZN(n17391) );
  INV_X1 U20471 ( .A(n17395), .ZN(n17389) );
  OAI211_X1 U20472 ( .C1(n17389), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17458), .B(
        n17388), .ZN(n17390) );
  OAI211_X1 U20473 ( .C1(n17392), .C2(n17460), .A(n17391), .B(n17390), .ZN(
        P3_U2718) );
  AOI22_X1 U20474 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17394), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17393), .ZN(n17397) );
  OAI211_X1 U20475 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17399), .A(n17458), .B(
        n17395), .ZN(n17396) );
  OAI211_X1 U20476 ( .C1(n17398), .C2(n17460), .A(n17397), .B(n17396), .ZN(
        P3_U2719) );
  AOI211_X1 U20477 ( .C1(n17577), .C2(n17403), .A(n17435), .B(n17399), .ZN(
        n17400) );
  AOI21_X1 U20478 ( .B1(n17466), .B2(BUF2_REG_15__SCAN_IN), .A(n17400), .ZN(
        n17401) );
  OAI21_X1 U20479 ( .B1(n17402), .B2(n17460), .A(n17401), .ZN(P3_U2720) );
  INV_X1 U20480 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n17409) );
  INV_X1 U20481 ( .A(n17403), .ZN(n17408) );
  NAND2_X1 U20482 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .ZN(n17405) );
  INV_X1 U20483 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17561) );
  NOR3_X1 U20484 ( .A1(n17404), .A2(n21109), .A3(n17439), .ZN(n17429) );
  NAND2_X1 U20485 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17429), .ZN(n17428) );
  NOR2_X1 U20486 ( .A1(n17561), .A2(n17428), .ZN(n17423) );
  NAND2_X1 U20487 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17423), .ZN(n17414) );
  NOR2_X1 U20488 ( .A1(n17405), .A2(n17414), .ZN(n17412) );
  AOI21_X1 U20489 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17458), .A(n17412), .ZN(
        n17407) );
  OAI222_X1 U20490 ( .A1(n17463), .A2(n17409), .B1(n17408), .B2(n17407), .C1(
        n17460), .C2(n17406), .ZN(P3_U2721) );
  INV_X1 U20491 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17413) );
  INV_X1 U20492 ( .A(n17414), .ZN(n17421) );
  AOI22_X1 U20493 ( .A1(n17421), .A2(P3_EAX_REG_12__SCAN_IN), .B1(
        P3_EAX_REG_13__SCAN_IN), .B2(n17458), .ZN(n17411) );
  OAI222_X1 U20494 ( .A1(n17463), .A2(n17413), .B1(n17412), .B2(n17411), .C1(
        n17460), .C2(n17410), .ZN(P3_U2722) );
  INV_X1 U20495 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17418) );
  INV_X1 U20496 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17567) );
  NOR2_X1 U20497 ( .A1(n17567), .A2(n17414), .ZN(n17417) );
  AOI21_X1 U20498 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17458), .A(n17421), .ZN(
        n17416) );
  OAI222_X1 U20499 ( .A1(n17463), .A2(n17418), .B1(n17417), .B2(n17416), .C1(
        n17460), .C2(n17415), .ZN(P3_U2723) );
  INV_X1 U20500 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17422) );
  AOI21_X1 U20501 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17458), .A(n17423), .ZN(
        n17420) );
  OAI222_X1 U20502 ( .A1(n17463), .A2(n17422), .B1(n17421), .B2(n17420), .C1(
        n17460), .C2(n17419), .ZN(P3_U2724) );
  INV_X1 U20503 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17427) );
  AOI211_X1 U20504 ( .C1(n17561), .C2(n17428), .A(n17435), .B(n17423), .ZN(
        n17424) );
  AOI21_X1 U20505 ( .B1(n17465), .B2(n17425), .A(n17424), .ZN(n17426) );
  OAI21_X1 U20506 ( .B1(n17427), .B2(n17463), .A(n17426), .ZN(P3_U2725) );
  INV_X1 U20507 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17433) );
  INV_X1 U20508 ( .A(n17428), .ZN(n17432) );
  AOI21_X1 U20509 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17458), .A(n17429), .ZN(
        n17431) );
  OAI222_X1 U20510 ( .A1(n17463), .A2(n17433), .B1(n17432), .B2(n17431), .C1(
        n17460), .C2(n17430), .ZN(P3_U2726) );
  AOI211_X1 U20511 ( .C1(n21109), .C2(n17439), .A(n17435), .B(n17434), .ZN(
        n17436) );
  AOI21_X1 U20512 ( .B1(n17466), .B2(BUF2_REG_8__SCAN_IN), .A(n17436), .ZN(
        n17437) );
  OAI21_X1 U20513 ( .B1(n17438), .B2(n17460), .A(n17437), .ZN(P3_U2727) );
  INV_X1 U20514 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18304) );
  INV_X1 U20515 ( .A(n17439), .ZN(n17443) );
  INV_X1 U20516 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17545) );
  NOR3_X1 U20517 ( .A1(n17545), .A2(n17543), .A3(n17467), .ZN(n17457) );
  NAND2_X1 U20518 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17457), .ZN(n17453) );
  NOR2_X1 U20519 ( .A1(n17440), .A2(n17453), .ZN(n17449) );
  AOI22_X1 U20520 ( .A1(n17449), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17458), .ZN(n17442) );
  OAI222_X1 U20521 ( .A1(n17463), .A2(n18304), .B1(n17443), .B2(n17442), .C1(
        n17460), .C2(n17441), .ZN(P3_U2728) );
  AND2_X1 U20522 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17449), .ZN(n17446) );
  AOI21_X1 U20523 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17458), .A(n17449), .ZN(
        n17445) );
  OAI222_X1 U20524 ( .A1(n18300), .A2(n17463), .B1(n17446), .B2(n17445), .C1(
        n17460), .C2(n17444), .ZN(P3_U2729) );
  INV_X1 U20525 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17549) );
  NOR2_X1 U20526 ( .A1(n17549), .A2(n17453), .ZN(n17456) );
  AOI22_X1 U20527 ( .A1(n17456), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n17458), .ZN(n17448) );
  OAI222_X1 U20528 ( .A1(n18296), .A2(n17463), .B1(n17449), .B2(n17448), .C1(
        n17460), .C2(n17447), .ZN(P3_U2730) );
  INV_X1 U20529 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18292) );
  AND2_X1 U20530 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17456), .ZN(n17452) );
  AOI21_X1 U20531 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17458), .A(n17456), .ZN(
        n17451) );
  OAI222_X1 U20532 ( .A1(n18292), .A2(n17463), .B1(n17452), .B2(n17451), .C1(
        n17460), .C2(n17450), .ZN(P3_U2731) );
  INV_X1 U20533 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18288) );
  INV_X1 U20534 ( .A(n17453), .ZN(n17462) );
  AOI21_X1 U20535 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17458), .A(n17462), .ZN(
        n17455) );
  OAI222_X1 U20536 ( .A1(n18288), .A2(n17463), .B1(n17456), .B2(n17455), .C1(
        n17460), .C2(n17454), .ZN(P3_U2732) );
  AOI21_X1 U20537 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17458), .A(n17457), .ZN(
        n17461) );
  OAI222_X1 U20538 ( .A1(n18284), .A2(n17463), .B1(n17462), .B2(n17461), .C1(
        n17460), .C2(n17459), .ZN(P3_U2733) );
  AOI22_X1 U20539 ( .A1(n17466), .A2(BUF2_REG_1__SCAN_IN), .B1(n17465), .B2(
        n17464), .ZN(n17472) );
  NOR2_X1 U20540 ( .A1(n17543), .A2(n17467), .ZN(n17470) );
  NOR2_X1 U20541 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17467), .ZN(n17469) );
  OAI22_X1 U20542 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17470), .B1(n17469), .B2(
        n17468), .ZN(n17471) );
  NAND2_X1 U20543 ( .A1(n17472), .A2(n17471), .ZN(P3_U2734) );
  OR2_X1 U20544 ( .A1(n18905), .A2(n17938), .ZN(n18927) );
  NOR2_X4 U20545 ( .A1(n17507), .A2(n17491), .ZN(n17502) );
  AND2_X1 U20546 ( .A1(n17502), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20547 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17541) );
  AOI22_X1 U20548 ( .A1(n17507), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17474) );
  OAI21_X1 U20549 ( .B1(n17541), .B2(n17489), .A(n17474), .ZN(P3_U2737) );
  INV_X1 U20550 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U20551 ( .A1(n17507), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17475) );
  OAI21_X1 U20552 ( .B1(n17539), .B2(n17489), .A(n17475), .ZN(P3_U2738) );
  AOI22_X1 U20553 ( .A1(n17507), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17476) );
  OAI21_X1 U20554 ( .B1(n17537), .B2(n17489), .A(n17476), .ZN(P3_U2739) );
  INV_X1 U20555 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17535) );
  AOI22_X1 U20556 ( .A1(n17507), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17477) );
  OAI21_X1 U20557 ( .B1(n17535), .B2(n17489), .A(n17477), .ZN(P3_U2740) );
  AOI22_X1 U20558 ( .A1(n17507), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17478) );
  OAI21_X1 U20559 ( .B1(n17533), .B2(n17489), .A(n17478), .ZN(P3_U2741) );
  INV_X1 U20560 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17531) );
  AOI22_X1 U20561 ( .A1(n17507), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17479) );
  OAI21_X1 U20562 ( .B1(n17531), .B2(n17489), .A(n17479), .ZN(P3_U2742) );
  INV_X1 U20563 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17529) );
  INV_X2 U20564 ( .A(n18927), .ZN(n17507) );
  AOI22_X1 U20565 ( .A1(n17507), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17480) );
  OAI21_X1 U20566 ( .B1(n17529), .B2(n17489), .A(n17480), .ZN(P3_U2743) );
  INV_X1 U20567 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17527) );
  AOI22_X1 U20568 ( .A1(n17507), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17481) );
  OAI21_X1 U20569 ( .B1(n17527), .B2(n17489), .A(n17481), .ZN(P3_U2744) );
  INV_X1 U20570 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17525) );
  AOI22_X1 U20571 ( .A1(n17507), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17482) );
  OAI21_X1 U20572 ( .B1(n17525), .B2(n17489), .A(n17482), .ZN(P3_U2745) );
  AOI22_X1 U20573 ( .A1(n17507), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17483) );
  OAI21_X1 U20574 ( .B1(n17523), .B2(n17489), .A(n17483), .ZN(P3_U2746) );
  INV_X1 U20575 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20986) );
  AOI22_X1 U20576 ( .A1(n17507), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17484) );
  OAI21_X1 U20577 ( .B1(n20986), .B2(n17489), .A(n17484), .ZN(P3_U2747) );
  INV_X1 U20578 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17520) );
  AOI22_X1 U20579 ( .A1(n17507), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17485) );
  OAI21_X1 U20580 ( .B1(n17520), .B2(n17489), .A(n17485), .ZN(P3_U2748) );
  AOI22_X1 U20581 ( .A1(n17507), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17486) );
  OAI21_X1 U20582 ( .B1(n17518), .B2(n17489), .A(n17486), .ZN(P3_U2749) );
  AOI22_X1 U20583 ( .A1(n17507), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17487) );
  OAI21_X1 U20584 ( .B1(n17516), .B2(n17489), .A(n17487), .ZN(P3_U2750) );
  INV_X1 U20585 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U20586 ( .A1(n17507), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17488) );
  OAI21_X1 U20587 ( .B1(n17514), .B2(n17489), .A(n17488), .ZN(P3_U2751) );
  AOI22_X1 U20588 ( .A1(n17507), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17490) );
  OAI21_X1 U20589 ( .B1(n17577), .B2(n17509), .A(n17490), .ZN(P3_U2752) );
  INV_X1 U20590 ( .A(P3_LWORD_REG_14__SCAN_IN), .ZN(n17572) );
  AOI22_X1 U20591 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17491), .B1(n17502), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17492) );
  OAI21_X1 U20592 ( .B1(n18927), .B2(n17572), .A(n17492), .ZN(P3_U2753) );
  INV_X1 U20593 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17569) );
  AOI22_X1 U20594 ( .A1(n17507), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17493) );
  OAI21_X1 U20595 ( .B1(n17569), .B2(n17509), .A(n17493), .ZN(P3_U2754) );
  AOI22_X1 U20596 ( .A1(n17507), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17494) );
  OAI21_X1 U20597 ( .B1(n17567), .B2(n17509), .A(n17494), .ZN(P3_U2755) );
  INV_X1 U20598 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17563) );
  AOI22_X1 U20599 ( .A1(n17507), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17495) );
  OAI21_X1 U20600 ( .B1(n17563), .B2(n17509), .A(n17495), .ZN(P3_U2756) );
  AOI22_X1 U20601 ( .A1(n17507), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17496) );
  OAI21_X1 U20602 ( .B1(n17561), .B2(n17509), .A(n17496), .ZN(P3_U2757) );
  INV_X1 U20603 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17559) );
  AOI22_X1 U20604 ( .A1(n17507), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17497) );
  OAI21_X1 U20605 ( .B1(n17559), .B2(n17509), .A(n17497), .ZN(P3_U2758) );
  AOI22_X1 U20606 ( .A1(n17507), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17498) );
  OAI21_X1 U20607 ( .B1(n21109), .B2(n17509), .A(n17498), .ZN(P3_U2759) );
  INV_X1 U20608 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17556) );
  AOI22_X1 U20609 ( .A1(n17507), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17499) );
  OAI21_X1 U20610 ( .B1(n17556), .B2(n17509), .A(n17499), .ZN(P3_U2760) );
  INV_X1 U20611 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U20612 ( .A1(n17507), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17500) );
  OAI21_X1 U20613 ( .B1(n17554), .B2(n17509), .A(n17500), .ZN(P3_U2761) );
  INV_X1 U20614 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n21096) );
  AOI22_X1 U20615 ( .A1(n17507), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17501) );
  OAI21_X1 U20616 ( .B1(n21096), .B2(n17509), .A(n17501), .ZN(P3_U2762) );
  INV_X1 U20617 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17551) );
  AOI22_X1 U20618 ( .A1(n17507), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17503) );
  OAI21_X1 U20619 ( .B1(n17551), .B2(n17509), .A(n17503), .ZN(P3_U2763) );
  AOI22_X1 U20620 ( .A1(n17507), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17504) );
  OAI21_X1 U20621 ( .B1(n17549), .B2(n17509), .A(n17504), .ZN(P3_U2764) );
  AOI22_X1 U20622 ( .A1(n17507), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17505) );
  OAI21_X1 U20623 ( .B1(n17547), .B2(n17509), .A(n17505), .ZN(P3_U2765) );
  AOI22_X1 U20624 ( .A1(n17507), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17506) );
  OAI21_X1 U20625 ( .B1(n17545), .B2(n17509), .A(n17506), .ZN(P3_U2766) );
  AOI22_X1 U20626 ( .A1(n17507), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17502), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17508) );
  OAI21_X1 U20627 ( .B1(n17543), .B2(n17509), .A(n17508), .ZN(P3_U2767) );
  NOR2_X1 U20628 ( .A1(n18929), .A2(n17510), .ZN(n18765) );
  AND2_X1 U20629 ( .A1(n17511), .A2(n18765), .ZN(n17570) );
  OAI211_X1 U20630 ( .C1(n18281), .C2(n18794), .A(n17512), .B(n17511), .ZN(
        n17574) );
  AOI22_X1 U20631 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17575), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17564), .ZN(n17513) );
  OAI21_X1 U20632 ( .B1(n17514), .B2(n9646), .A(n17513), .ZN(P3_U2768) );
  AOI22_X1 U20633 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17575), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17564), .ZN(n17515) );
  OAI21_X1 U20634 ( .B1(n17516), .B2(n9646), .A(n17515), .ZN(P3_U2769) );
  AOI22_X1 U20635 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17575), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17564), .ZN(n17517) );
  OAI21_X1 U20636 ( .B1(n17518), .B2(n9646), .A(n17517), .ZN(P3_U2770) );
  AOI22_X1 U20637 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17564), .ZN(n17519) );
  OAI21_X1 U20638 ( .B1(n17520), .B2(n9646), .A(n17519), .ZN(P3_U2771) );
  AOI22_X1 U20639 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17564), .ZN(n17521) );
  OAI21_X1 U20640 ( .B1(n20986), .B2(n9646), .A(n17521), .ZN(P3_U2772) );
  AOI22_X1 U20641 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17564), .ZN(n17522) );
  OAI21_X1 U20642 ( .B1(n17523), .B2(n9646), .A(n17522), .ZN(P3_U2773) );
  AOI22_X1 U20643 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17564), .ZN(n17524) );
  OAI21_X1 U20644 ( .B1(n17525), .B2(n9646), .A(n17524), .ZN(P3_U2774) );
  AOI22_X1 U20645 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17564), .ZN(n17526) );
  OAI21_X1 U20646 ( .B1(n17527), .B2(n9646), .A(n17526), .ZN(P3_U2775) );
  AOI22_X1 U20647 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17564), .ZN(n17528) );
  OAI21_X1 U20648 ( .B1(n17529), .B2(n9646), .A(n17528), .ZN(P3_U2776) );
  AOI22_X1 U20649 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17564), .ZN(n17530) );
  OAI21_X1 U20650 ( .B1(n17531), .B2(n9646), .A(n17530), .ZN(P3_U2777) );
  AOI22_X1 U20651 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17564), .ZN(n17532) );
  OAI21_X1 U20652 ( .B1(n17533), .B2(n9646), .A(n17532), .ZN(P3_U2778) );
  AOI22_X1 U20653 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17574), .ZN(n17534) );
  OAI21_X1 U20654 ( .B1(n17535), .B2(n9646), .A(n17534), .ZN(P3_U2779) );
  AOI22_X1 U20655 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17575), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17574), .ZN(n17536) );
  OAI21_X1 U20656 ( .B1(n17537), .B2(n9646), .A(n17536), .ZN(P3_U2780) );
  AOI22_X1 U20657 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17575), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17574), .ZN(n17538) );
  OAI21_X1 U20658 ( .B1(n17539), .B2(n9646), .A(n17538), .ZN(P3_U2781) );
  AOI22_X1 U20659 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17575), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17574), .ZN(n17540) );
  OAI21_X1 U20660 ( .B1(n17541), .B2(n9646), .A(n17540), .ZN(P3_U2782) );
  AOI22_X1 U20661 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17574), .ZN(n17542) );
  OAI21_X1 U20662 ( .B1(n17543), .B2(n9646), .A(n17542), .ZN(P3_U2783) );
  AOI22_X1 U20663 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17574), .ZN(n17544) );
  OAI21_X1 U20664 ( .B1(n17545), .B2(n9646), .A(n17544), .ZN(P3_U2784) );
  AOI22_X1 U20665 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17574), .ZN(n17546) );
  OAI21_X1 U20666 ( .B1(n17547), .B2(n9646), .A(n17546), .ZN(P3_U2785) );
  AOI22_X1 U20667 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17574), .ZN(n17548) );
  OAI21_X1 U20668 ( .B1(n17549), .B2(n9646), .A(n17548), .ZN(P3_U2786) );
  AOI22_X1 U20669 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17564), .ZN(n17550) );
  OAI21_X1 U20670 ( .B1(n17551), .B2(n9646), .A(n17550), .ZN(P3_U2787) );
  AOI22_X1 U20671 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17564), .ZN(n17552) );
  OAI21_X1 U20672 ( .B1(n21096), .B2(n9646), .A(n17552), .ZN(P3_U2788) );
  AOI22_X1 U20673 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17564), .ZN(n17553) );
  OAI21_X1 U20674 ( .B1(n17554), .B2(n9646), .A(n17553), .ZN(P3_U2789) );
  AOI22_X1 U20675 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17564), .ZN(n17555) );
  OAI21_X1 U20676 ( .B1(n17556), .B2(n9646), .A(n17555), .ZN(P3_U2790) );
  AOI22_X1 U20677 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17564), .ZN(n17557) );
  OAI21_X1 U20678 ( .B1(n21109), .B2(n9646), .A(n17557), .ZN(P3_U2791) );
  AOI22_X1 U20679 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17564), .ZN(n17558) );
  OAI21_X1 U20680 ( .B1(n17559), .B2(n9646), .A(n17558), .ZN(P3_U2792) );
  AOI22_X1 U20681 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17565), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17564), .ZN(n17560) );
  OAI21_X1 U20682 ( .B1(n17561), .B2(n9646), .A(n17560), .ZN(P3_U2793) );
  AOI22_X1 U20683 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17564), .ZN(n17562) );
  OAI21_X1 U20684 ( .B1(n17563), .B2(n9646), .A(n17562), .ZN(P3_U2794) );
  AOI22_X1 U20685 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17565), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17564), .ZN(n17566) );
  OAI21_X1 U20686 ( .B1(n17567), .B2(n9646), .A(n17566), .ZN(P3_U2795) );
  AOI22_X1 U20687 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17574), .ZN(n17568) );
  OAI21_X1 U20688 ( .B1(n17569), .B2(n9646), .A(n17568), .ZN(P3_U2796) );
  AOI22_X1 U20689 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17575), .B1(
        P3_EAX_REG_14__SCAN_IN), .B2(n17570), .ZN(n17571) );
  OAI21_X1 U20690 ( .B1(n17573), .B2(n17572), .A(n17571), .ZN(P3_U2797) );
  AOI22_X1 U20691 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17575), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17574), .ZN(n17576) );
  OAI21_X1 U20692 ( .B1(n17577), .B2(n9646), .A(n17576), .ZN(P3_U2798) );
  INV_X1 U20693 ( .A(n17578), .ZN(n17579) );
  OAI21_X1 U20694 ( .B1(n17579), .B2(n17938), .A(n17939), .ZN(n17580) );
  AOI21_X1 U20695 ( .B1(n18783), .B2(n17589), .A(n17580), .ZN(n17611) );
  OAI21_X1 U20696 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17648), .A(
        n17611), .ZN(n17601) );
  AOI22_X1 U20697 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17601), .B1(
        n17799), .B2(n17581), .ZN(n17594) );
  INV_X1 U20698 ( .A(n17751), .ZN(n17642) );
  NOR2_X1 U20699 ( .A1(n17932), .A2(n17774), .ZN(n17696) );
  OAI22_X1 U20700 ( .A1(n17951), .A2(n17943), .B1(n17950), .B2(n17850), .ZN(
        n17615) );
  NOR2_X1 U20701 ( .A1(n17945), .A2(n17615), .ZN(n17582) );
  NOR3_X1 U20702 ( .A1(n17696), .A2(n17582), .A3(n21110), .ZN(n17587) );
  AOI211_X1 U20703 ( .C1(n17585), .C2(n17584), .A(n17583), .B(n17851), .ZN(
        n17586) );
  AOI211_X1 U20704 ( .C1(n17588), .C2(n17642), .A(n17587), .B(n17586), .ZN(
        n17593) );
  NAND2_X1 U20705 ( .A1(n18252), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17592) );
  NOR2_X1 U20706 ( .A1(n17705), .A2(n17589), .ZN(n17603) );
  OAI211_X1 U20707 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17603), .B(n17590), .ZN(n17591) );
  NAND4_X1 U20708 ( .A1(n17594), .A2(n17593), .A3(n17592), .A4(n17591), .ZN(
        P3_U2802) );
  INV_X1 U20709 ( .A(n17595), .ZN(n17596) );
  NAND2_X1 U20710 ( .A1(n17597), .A2(n17596), .ZN(n17598) );
  XOR2_X1 U20711 ( .A(n17598), .B(n17849), .Z(n17959) );
  INV_X1 U20712 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17602) );
  OAI22_X1 U20713 ( .A1(n18236), .A2(n18858), .B1(n17787), .B2(n17599), .ZN(
        n17600) );
  AOI221_X1 U20714 ( .B1(n17603), .B2(n17602), .C1(n17601), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17600), .ZN(n17606) );
  AOI22_X1 U20715 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17615), .B1(
        n17604), .B2(n17945), .ZN(n17605) );
  OAI211_X1 U20716 ( .C1(n17959), .C2(n17851), .A(n17606), .B(n17605), .ZN(
        P3_U2803) );
  AOI21_X1 U20717 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17608), .A(
        n17607), .ZN(n17966) );
  AOI21_X1 U20718 ( .B1(n18655), .B2(n17609), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17610) );
  OAI22_X1 U20719 ( .A1(n17611), .A2(n17610), .B1(n18236), .B2(n18856), .ZN(
        n17612) );
  AOI221_X1 U20720 ( .B1(n17799), .B2(n17613), .C1(n17689), .C2(n17613), .A(
        n17612), .ZN(n17617) );
  NOR2_X1 U20721 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17614), .ZN(
        n17965) );
  AOI22_X1 U20722 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17615), .B1(
        n17656), .B2(n17965), .ZN(n17616) );
  OAI211_X1 U20723 ( .C1(n17966), .C2(n17851), .A(n17617), .B(n17616), .ZN(
        P3_U2804) );
  OAI21_X1 U20724 ( .B1(n17849), .B2(n17619), .A(n17618), .ZN(n17620) );
  XOR2_X1 U20725 ( .A(n17620), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17978) );
  NAND2_X1 U20726 ( .A1(n18655), .A2(n17623), .ZN(n17653) );
  OAI211_X1 U20727 ( .C1(n17621), .C2(n17938), .A(n17939), .B(n17653), .ZN(
        n17650) );
  AOI21_X1 U20728 ( .B1(n17689), .B2(n17622), .A(n17650), .ZN(n17637) );
  INV_X1 U20729 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21128) );
  NOR2_X1 U20730 ( .A1(n17705), .A2(n17623), .ZN(n17640) );
  OAI211_X1 U20731 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17640), .B(n17624), .ZN(n17625) );
  NAND2_X1 U20732 ( .A1(n18151), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17976) );
  OAI211_X1 U20733 ( .C1(n17637), .C2(n21128), .A(n17625), .B(n17976), .ZN(
        n17626) );
  AOI21_X1 U20734 ( .B1(n17799), .B2(n17627), .A(n17626), .ZN(n17633) );
  AOI21_X1 U20735 ( .B1(n17948), .B2(n17629), .A(n17628), .ZN(n17972) );
  AOI21_X1 U20736 ( .B1(n17948), .B2(n17631), .A(n17630), .ZN(n17968) );
  AOI22_X1 U20737 ( .A1(n17932), .A2(n17972), .B1(n17774), .B2(n17968), .ZN(
        n17632) );
  OAI211_X1 U20738 ( .C1(n17851), .C2(n17978), .A(n17633), .B(n17632), .ZN(
        P3_U2805) );
  AOI21_X1 U20739 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17635), .A(
        n17634), .ZN(n17993) );
  NOR2_X1 U20740 ( .A1(n18236), .A2(n18851), .ZN(n17979) );
  OAI22_X1 U20741 ( .A1(n17637), .A2(n17639), .B1(n17787), .B2(n16652), .ZN(
        n17638) );
  AOI211_X1 U20742 ( .C1(n17640), .C2(n17639), .A(n17979), .B(n17638), .ZN(
        n17644) );
  OAI22_X1 U20743 ( .A1(n17986), .A2(n17943), .B1(n17981), .B2(n17850), .ZN(
        n17655) );
  NOR2_X1 U20744 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17641), .ZN(
        n17980) );
  AOI22_X1 U20745 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17655), .B1(
        n17642), .B2(n17980), .ZN(n17643) );
  OAI211_X1 U20746 ( .C1(n17993), .C2(n17851), .A(n17644), .B(n17643), .ZN(
        P3_U2806) );
  AOI22_X1 U20747 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17849), .B1(
        n17645), .B2(n17666), .ZN(n17646) );
  NAND2_X1 U20748 ( .A1(n17684), .A2(n17646), .ZN(n17647) );
  XOR2_X1 U20749 ( .A(n17647), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n17998) );
  NAND2_X1 U20750 ( .A1(n17787), .A2(n17648), .ZN(n17725) );
  AOI22_X1 U20751 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17650), .B1(
        n17649), .B2(n17725), .ZN(n17651) );
  NAND2_X1 U20752 ( .A1(n18151), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17997) );
  OAI211_X1 U20753 ( .C1(n17653), .C2(n17652), .A(n17651), .B(n17997), .ZN(
        n17654) );
  AOI221_X1 U20754 ( .B1(n17656), .B2(n17987), .C1(n17655), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17654), .ZN(n17657) );
  OAI21_X1 U20755 ( .B1(n17851), .B2(n17998), .A(n17657), .ZN(P3_U2807) );
  INV_X1 U20756 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18015) );
  NAND2_X1 U20757 ( .A1(n18004), .A2(n18015), .ZN(n18009) );
  NAND2_X1 U20758 ( .A1(n10229), .A2(n17741), .ZN(n17677) );
  AOI211_X1 U20759 ( .C1(n17676), .C2(n17662), .A(n17658), .B(n17677), .ZN(
        n17664) );
  INV_X1 U20760 ( .A(n10229), .ZN(n17659) );
  AOI22_X1 U20761 ( .A1(n17782), .A2(n17660), .B1(n18783), .B2(n17659), .ZN(
        n17661) );
  NAND2_X1 U20762 ( .A1(n17661), .A2(n17939), .ZN(n17695) );
  AOI21_X1 U20763 ( .B1(n17689), .B2(n17687), .A(n17695), .ZN(n17675) );
  NAND2_X1 U20764 ( .A1(n18151), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18013) );
  OAI21_X1 U20765 ( .B1(n17675), .B2(n17662), .A(n18013), .ZN(n17663) );
  AOI211_X1 U20766 ( .C1(n17665), .C2(n17799), .A(n17664), .B(n17663), .ZN(
        n17670) );
  AOI22_X1 U20767 ( .A1(n9653), .A2(n18075), .B1(n17774), .B2(n18077), .ZN(
        n17750) );
  OAI21_X1 U20768 ( .B1(n18004), .B2(n17696), .A(n17750), .ZN(n17681) );
  INV_X1 U20769 ( .A(n17666), .ZN(n17667) );
  OAI221_X1 U20770 ( .B1(n17667), .B2(n18004), .C1(n17667), .C2(n17737), .A(
        n17684), .ZN(n17668) );
  XOR2_X1 U20771 ( .A(n18015), .B(n17668), .Z(n18011) );
  AOI22_X1 U20772 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17681), .B1(
        n17748), .B2(n18011), .ZN(n17669) );
  OAI211_X1 U20773 ( .C1(n17751), .C2(n18009), .A(n17670), .B(n17669), .ZN(
        P3_U2808) );
  INV_X1 U20774 ( .A(n17680), .ZN(n18003) );
  NOR3_X1 U20775 ( .A1(n17714), .A2(n17849), .A3(n17671), .ZN(n17699) );
  AOI22_X1 U20776 ( .A1(n18003), .A2(n17699), .B1(n9840), .B2(n17673), .ZN(
        n17674) );
  XOR2_X1 U20777 ( .A(n17674), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n18027) );
  NAND2_X1 U20778 ( .A1(n18252), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18025) );
  OAI221_X1 U20779 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17677), .C1(
        n17676), .C2(n17675), .A(n18025), .ZN(n17678) );
  AOI21_X1 U20780 ( .B1(n17799), .B2(n17679), .A(n17678), .ZN(n17683) );
  NOR2_X1 U20781 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17680), .ZN(
        n18024) );
  NAND2_X1 U20782 ( .A1(n18047), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18017) );
  NOR2_X1 U20783 ( .A1(n17751), .A2(n18017), .ZN(n17712) );
  AOI22_X1 U20784 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17681), .B1(
        n18024), .B2(n17712), .ZN(n17682) );
  OAI211_X1 U20785 ( .C1(n18027), .C2(n17851), .A(n17683), .B(n17682), .ZN(
        P3_U2809) );
  OAI221_X1 U20786 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17721), 
        .C1(n18035), .C2(n17699), .A(n17684), .ZN(n17685) );
  XOR2_X1 U20787 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17685), .Z(
        n18034) );
  INV_X1 U20788 ( .A(n17686), .ZN(n17688) );
  OAI21_X1 U20789 ( .B1(n17688), .B2(n18373), .A(n17687), .ZN(n17694) );
  INV_X1 U20790 ( .A(n17690), .ZN(n17691) );
  AOI21_X1 U20791 ( .B1(n17787), .B2(n17648), .A(n17691), .ZN(n17693) );
  NOR2_X1 U20792 ( .A1(n18236), .A2(n18844), .ZN(n17692) );
  AOI211_X1 U20793 ( .C1(n17695), .C2(n17694), .A(n17693), .B(n17692), .ZN(
        n17698) );
  NOR2_X1 U20794 ( .A1(n18035), .A2(n18017), .ZN(n18030) );
  OAI21_X1 U20795 ( .B1(n17696), .B2(n18030), .A(n17750), .ZN(n17711) );
  NOR2_X1 U20796 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18035), .ZN(
        n18028) );
  AOI22_X1 U20797 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17711), .B1(
        n17712), .B2(n18028), .ZN(n17697) );
  OAI211_X1 U20798 ( .C1(n17851), .C2(n18034), .A(n17698), .B(n17697), .ZN(
        P3_U2810) );
  AOI21_X1 U20799 ( .B1(n9840), .B2(n17721), .A(n17699), .ZN(n17700) );
  XOR2_X1 U20800 ( .A(n17700), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n18040) );
  INV_X1 U20801 ( .A(n17939), .ZN(n17912) );
  AOI21_X1 U20802 ( .B1(n17704), .B2(n18783), .A(n17912), .ZN(n17726) );
  OAI21_X1 U20803 ( .B1(n17938), .B2(n17701), .A(n17726), .ZN(n17702) );
  INV_X1 U20804 ( .A(n17702), .ZN(n17716) );
  AOI22_X1 U20805 ( .A1(n18252), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n17799), 
        .B2(n17703), .ZN(n17708) );
  NOR2_X1 U20806 ( .A1(n17705), .A2(n17704), .ZN(n17715) );
  OAI211_X1 U20807 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17715), .B(n17706), .ZN(n17707) );
  OAI211_X1 U20808 ( .C1(n17716), .C2(n17709), .A(n17708), .B(n17707), .ZN(
        n17710) );
  AOI221_X1 U20809 ( .B1(n17712), .B2(n18035), .C1(n17711), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17710), .ZN(n17713) );
  OAI21_X1 U20810 ( .B1(n18040), .B2(n17851), .A(n17713), .ZN(P3_U2811) );
  NAND2_X1 U20811 ( .A1(n18047), .A2(n17714), .ZN(n18055) );
  INV_X1 U20812 ( .A(n17715), .ZN(n17718) );
  NAND2_X1 U20813 ( .A1(n18252), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18053) );
  OAI221_X1 U20814 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17718), .C1(
        n17717), .C2(n17716), .A(n18053), .ZN(n17719) );
  AOI21_X1 U20815 ( .B1(n17799), .B2(n17720), .A(n17719), .ZN(n17724) );
  OAI21_X1 U20816 ( .B1(n18047), .B2(n17751), .A(n17750), .ZN(n17733) );
  AOI21_X1 U20817 ( .B1(n17833), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17721), .ZN(n17722) );
  XOR2_X1 U20818 ( .A(n17722), .B(n9840), .Z(n18051) );
  AOI22_X1 U20819 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17733), .B1(
        n17748), .B2(n18051), .ZN(n17723) );
  OAI211_X1 U20820 ( .C1(n17751), .C2(n18055), .A(n17724), .B(n17723), .ZN(
        P3_U2812) );
  NAND2_X1 U20821 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18056), .ZN(
        n18062) );
  INV_X1 U20822 ( .A(n17725), .ZN(n17924) );
  AOI221_X1 U20823 ( .B1(n17728), .B2(n17727), .C1(n18373), .C2(n17727), .A(
        n17726), .ZN(n17729) );
  NOR2_X1 U20824 ( .A1(n18236), .A2(n18838), .ZN(n18059) );
  AOI211_X1 U20825 ( .C1(n17730), .C2(n17725), .A(n17729), .B(n18059), .ZN(
        n17735) );
  OAI21_X1 U20826 ( .B1(n17732), .B2(n18056), .A(n17731), .ZN(n18060) );
  AOI22_X1 U20827 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17733), .B1(
        n17748), .B2(n18060), .ZN(n17734) );
  OAI211_X1 U20828 ( .C1(n17751), .C2(n18062), .A(n17735), .B(n17734), .ZN(
        P3_U2813) );
  INV_X1 U20829 ( .A(n18125), .ZN(n17813) );
  NAND2_X1 U20830 ( .A1(n17833), .A2(n17813), .ZN(n17832) );
  OAI22_X1 U20831 ( .A1(n17833), .A2(n17737), .B1(n17832), .B2(n17736), .ZN(
        n17738) );
  XOR2_X1 U20832 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17738), .Z(
        n18069) );
  AOI21_X1 U20833 ( .B1(n18783), .B2(n17739), .A(n17912), .ZN(n17767) );
  OAI21_X1 U20834 ( .B1(n17740), .B2(n17938), .A(n17767), .ZN(n17753) );
  AOI22_X1 U20835 ( .A1(n18252), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17753), .ZN(n17745) );
  NAND2_X1 U20836 ( .A1(n9779), .A2(n17741), .ZN(n17802) );
  NOR2_X1 U20837 ( .A1(n17742), .A2(n17802), .ZN(n17763) );
  OAI211_X1 U20838 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17763), .B(n17743), .ZN(n17744) );
  OAI211_X1 U20839 ( .C1(n17787), .C2(n17746), .A(n17745), .B(n17744), .ZN(
        n17747) );
  AOI21_X1 U20840 ( .B1(n17748), .B2(n18069), .A(n17747), .ZN(n17749) );
  OAI221_X1 U20841 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17751), 
        .C1(n18073), .C2(n17750), .A(n17749), .ZN(P3_U2814) );
  NOR2_X1 U20842 ( .A1(n17771), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18089) );
  NAND2_X1 U20843 ( .A1(n17932), .A2(n18075), .ZN(n17765) );
  AOI22_X1 U20844 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17753), .B1(
        n17799), .B2(n17752), .ZN(n17754) );
  NAND2_X1 U20845 ( .A1(n18252), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18086) );
  NAND2_X1 U20846 ( .A1(n17754), .A2(n18086), .ZN(n17761) );
  NOR2_X1 U20847 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17772), .ZN(
        n18080) );
  NAND2_X1 U20848 ( .A1(n17774), .A2(n18077), .ZN(n17759) );
  INV_X1 U20849 ( .A(n18134), .ZN(n18117) );
  NAND3_X1 U20850 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18117), .A3(
        n17755), .ZN(n17757) );
  INV_X1 U20851 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17779) );
  NOR4_X1 U20852 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n17833), .A4(n15905), .ZN(
        n17811) );
  INV_X1 U20853 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17815) );
  NAND2_X1 U20854 ( .A1(n17811), .A2(n17815), .ZN(n17795) );
  AOI22_X1 U20855 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17833), .B1(
        n18106), .B2(n17805), .ZN(n17756) );
  AOI221_X1 U20856 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17757), 
        .C1(n17779), .C2(n17795), .A(n17756), .ZN(n17758) );
  XOR2_X1 U20857 ( .A(n18081), .B(n17758), .Z(n18078) );
  OAI22_X1 U20858 ( .A1(n18080), .A2(n17759), .B1(n17851), .B2(n18078), .ZN(
        n17760) );
  AOI211_X1 U20859 ( .C1(n17763), .C2(n17762), .A(n17761), .B(n17760), .ZN(
        n17764) );
  OAI21_X1 U20860 ( .B1(n18089), .B2(n17765), .A(n17764), .ZN(P3_U2815) );
  INV_X1 U20861 ( .A(n17773), .ZN(n18095) );
  NOR2_X1 U20862 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17795), .ZN(
        n17777) );
  AOI22_X1 U20863 ( .A1(n17822), .A2(n18095), .B1(n17777), .B2(n17779), .ZN(
        n17766) );
  XOR2_X1 U20864 ( .A(n17766), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18100) );
  INV_X1 U20865 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18831) );
  NOR2_X1 U20866 ( .A1(n18236), .A2(n18831), .ZN(n18103) );
  NAND2_X1 U20867 ( .A1(n9779), .A2(n18655), .ZN(n17810) );
  AOI221_X1 U20868 ( .B1(n17784), .B2(n17768), .C1(n17810), .C2(n17768), .A(
        n17767), .ZN(n17769) );
  AOI211_X1 U20869 ( .C1(n17770), .C2(n17725), .A(n18103), .B(n17769), .ZN(
        n17776) );
  INV_X1 U20870 ( .A(n18094), .ZN(n17791) );
  NOR2_X1 U20871 ( .A1(n17791), .A2(n18127), .ZN(n17790) );
  INV_X1 U20872 ( .A(n17790), .ZN(n18111) );
  AOI221_X1 U20873 ( .B1(n17779), .B2(n18106), .C1(n18111), .C2(n18106), .A(
        n17771), .ZN(n18101) );
  AOI221_X1 U20874 ( .B1(n17773), .B2(n18106), .C1(n18125), .C2(n18106), .A(
        n17772), .ZN(n18091) );
  AOI22_X1 U20875 ( .A1(n9653), .A2(n18101), .B1(n17774), .B2(n18091), .ZN(
        n17775) );
  OAI211_X1 U20876 ( .C1(n18100), .C2(n17851), .A(n17776), .B(n17775), .ZN(
        P3_U2816) );
  NAND3_X1 U20877 ( .A1(n18131), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n17822), .ZN(n17794) );
  INV_X1 U20878 ( .A(n17777), .ZN(n17778) );
  OAI21_X1 U20879 ( .B1(n17805), .B2(n17794), .A(n17778), .ZN(n17780) );
  XOR2_X1 U20880 ( .A(n17780), .B(n17779), .Z(n18116) );
  AOI21_X1 U20881 ( .B1(n17782), .B2(n17781), .A(n17912), .ZN(n17783) );
  OAI21_X1 U20882 ( .B1(n9779), .B2(n17897), .A(n17783), .ZN(n17800) );
  NOR2_X1 U20883 ( .A1(n18236), .A2(n18829), .ZN(n17789) );
  OAI21_X1 U20884 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17784), .ZN(n17785) );
  OAI22_X1 U20885 ( .A1(n17787), .A2(n17786), .B1(n17802), .B2(n17785), .ZN(
        n17788) );
  AOI211_X1 U20886 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17800), .A(
        n17789), .B(n17788), .ZN(n17793) );
  NOR2_X1 U20887 ( .A1(n17791), .A2(n18125), .ZN(n18108) );
  OAI22_X1 U20888 ( .A1(n17790), .A2(n17943), .B1(n18108), .B2(n17850), .ZN(
        n17804) );
  NOR2_X1 U20889 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17791), .ZN(
        n18107) );
  AOI22_X1 U20890 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17804), .B1(
        n18107), .B2(n17841), .ZN(n17792) );
  OAI211_X1 U20891 ( .C1(n18116), .C2(n17851), .A(n17793), .B(n17792), .ZN(
        P3_U2817) );
  NAND2_X1 U20892 ( .A1(n17795), .A2(n17794), .ZN(n17796) );
  XOR2_X1 U20893 ( .A(n17805), .B(n17796), .Z(n18123) );
  INV_X1 U20894 ( .A(n17841), .ZN(n17797) );
  NOR2_X1 U20895 ( .A1(n17797), .A2(n18134), .ZN(n17806) );
  AOI22_X1 U20896 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17800), .B1(
        n17799), .B2(n17798), .ZN(n17801) );
  NAND2_X1 U20897 ( .A1(n18151), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18121) );
  OAI211_X1 U20898 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17802), .A(
        n17801), .B(n18121), .ZN(n17803) );
  AOI221_X1 U20899 ( .B1(n17806), .B2(n17805), .C1(n17804), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17803), .ZN(n17807) );
  OAI21_X1 U20900 ( .B1(n18123), .B2(n17851), .A(n17807), .ZN(P3_U2818) );
  NAND2_X1 U20901 ( .A1(n17939), .A2(n17897), .ZN(n17934) );
  NAND3_X1 U20902 ( .A1(n17878), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18655), .ZN(n17860) );
  OAI22_X1 U20903 ( .A1(n17877), .A2(n17808), .B1(n17828), .B2(n17860), .ZN(
        n17809) );
  AOI22_X1 U20904 ( .A1(n18252), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17810), 
        .B2(n17809), .ZN(n17818) );
  INV_X1 U20905 ( .A(n18131), .ZN(n17814) );
  NOR2_X1 U20906 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17814), .ZN(
        n18124) );
  AOI21_X1 U20907 ( .B1(n17822), .B2(n18131), .A(n17811), .ZN(n17812) );
  XOR2_X1 U20908 ( .A(n17812), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18139) );
  OAI22_X1 U20909 ( .A1(n17813), .A2(n17850), .B1(n17943), .B2(n9813), .ZN(
        n17842) );
  AOI21_X1 U20910 ( .B1(n17814), .B2(n17841), .A(n17842), .ZN(n17825) );
  OAI22_X1 U20911 ( .A1(n18139), .A2(n17851), .B1(n17825), .B2(n17815), .ZN(
        n17816) );
  AOI21_X1 U20912 ( .B1(n18124), .B2(n17841), .A(n17816), .ZN(n17817) );
  OAI211_X1 U20913 ( .C1(n17924), .C2(n17819), .A(n17818), .B(n17817), .ZN(
        P3_U2819) );
  NAND2_X1 U20914 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17853) );
  NOR2_X1 U20915 ( .A1(n17853), .A2(n17860), .ZN(n17836) );
  NAND2_X1 U20916 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17836), .ZN(
        n17835) );
  OAI21_X1 U20917 ( .B1(n17877), .B2(n17820), .A(n17835), .ZN(n17827) );
  NOR3_X1 U20918 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17833), .A3(
        n15905), .ZN(n17821) );
  AOI21_X1 U20919 ( .B1(n17822), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17821), .ZN(n17823) );
  XNOR2_X1 U20920 ( .A(n18145), .B(n17823), .ZN(n18148) );
  AOI21_X1 U20921 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17841), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17824) );
  OAI22_X1 U20922 ( .A1(n18148), .A2(n17851), .B1(n17825), .B2(n17824), .ZN(
        n17826) );
  AOI221_X1 U20923 ( .B1(n17828), .B2(n17827), .C1(n17860), .C2(n17827), .A(
        n17826), .ZN(n17830) );
  NAND2_X1 U20924 ( .A1(n18252), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17829) );
  OAI211_X1 U20925 ( .C1(n17924), .C2(n17831), .A(n17830), .B(n17829), .ZN(
        P3_U2820) );
  OAI21_X1 U20926 ( .B1(n15905), .B2(n17833), .A(n17832), .ZN(n17834) );
  XOR2_X1 U20927 ( .A(n17834), .B(n18149), .Z(n18157) );
  OAI211_X1 U20928 ( .C1(n17836), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17934), .B(n17835), .ZN(n17838) );
  NAND2_X1 U20929 ( .A1(n18252), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17837) );
  OAI211_X1 U20930 ( .C1(n17924), .C2(n17839), .A(n17838), .B(n17837), .ZN(
        n17840) );
  AOI221_X1 U20931 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17842), .C1(
        n18149), .C2(n17841), .A(n17840), .ZN(n17843) );
  OAI21_X1 U20932 ( .B1(n18157), .B2(n17851), .A(n17843), .ZN(P3_U2821) );
  OAI21_X1 U20933 ( .B1(n17844), .B2(n17897), .A(n17939), .ZN(n17861) );
  AOI22_X1 U20934 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17861), .B1(
        n17845), .B2(n17725), .ZN(n17857) );
  AOI21_X1 U20935 ( .B1(n17847), .B2(n18162), .A(n17846), .ZN(n18164) );
  AOI21_X1 U20936 ( .B1(n17849), .B2(n18167), .A(n17848), .ZN(n18173) );
  OAI22_X1 U20937 ( .A1(n18173), .A2(n17851), .B1(n17850), .B2(n18167), .ZN(
        n17852) );
  AOI21_X1 U20938 ( .B1(n17932), .B2(n18164), .A(n17852), .ZN(n17856) );
  NAND2_X1 U20939 ( .A1(n18252), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18170) );
  OAI211_X1 U20940 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17854), .A(
        n18655), .B(n17853), .ZN(n17855) );
  NAND4_X1 U20941 ( .A1(n17857), .A2(n17856), .A3(n18170), .A4(n17855), .ZN(
        P3_U2822) );
  OAI21_X1 U20942 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17859), .A(
        n17858), .ZN(n18182) );
  INV_X1 U20943 ( .A(n17860), .ZN(n17863) );
  NOR2_X1 U20944 ( .A1(n18236), .A2(n18818), .ZN(n18174) );
  AOI221_X1 U20945 ( .B1(n17863), .B2(n17862), .C1(n17861), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18174), .ZN(n17869) );
  NAND2_X1 U20946 ( .A1(n17865), .A2(n17864), .ZN(n17866) );
  INV_X1 U20947 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18177) );
  XOR2_X1 U20948 ( .A(n17866), .B(n18177), .Z(n18178) );
  AOI22_X1 U20949 ( .A1(n17932), .A2(n18178), .B1(n17867), .B2(n17725), .ZN(
        n17868) );
  OAI211_X1 U20950 ( .C1(n17942), .C2(n18182), .A(n17869), .B(n17868), .ZN(
        P3_U2823) );
  NAND2_X1 U20951 ( .A1(n17878), .A2(n18655), .ZN(n17873) );
  OAI21_X1 U20952 ( .B1(n17872), .B2(n17871), .A(n17870), .ZN(n18190) );
  OAI22_X1 U20953 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17873), .B1(
        n17942), .B2(n18190), .ZN(n17874) );
  AOI21_X1 U20954 ( .B1(n18252), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17874), .ZN(
        n17880) );
  AOI21_X1 U20955 ( .B1(n17876), .B2(n18186), .A(n17875), .ZN(n18185) );
  AOI21_X1 U20956 ( .B1(n18655), .B2(n17878), .A(n17877), .ZN(n17890) );
  AOI22_X1 U20957 ( .A1(n9653), .A2(n18185), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17890), .ZN(n17879) );
  OAI211_X1 U20958 ( .C1(n17924), .C2(n17881), .A(n17880), .B(n17879), .ZN(
        P3_U2824) );
  XOR2_X1 U20959 ( .A(n17882), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18195) );
  AOI22_X1 U20960 ( .A1(n17883), .A2(n18195), .B1(n18151), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17892) );
  AOI21_X1 U20961 ( .B1(n17886), .B2(n17885), .A(n17884), .ZN(n18194) );
  OAI21_X1 U20962 ( .B1(n17912), .B2(n17888), .A(n17887), .ZN(n17889) );
  AOI22_X1 U20963 ( .A1(n17932), .A2(n18194), .B1(n17890), .B2(n17889), .ZN(
        n17891) );
  OAI211_X1 U20964 ( .C1(n17924), .C2(n17893), .A(n17892), .B(n17891), .ZN(
        P3_U2825) );
  AOI21_X1 U20965 ( .B1(n17896), .B2(n17895), .A(n17894), .ZN(n18206) );
  AOI22_X1 U20966 ( .A1(n9653), .A2(n18206), .B1(n18151), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n17904) );
  OAI21_X1 U20967 ( .B1(n16966), .B2(n17897), .A(n17939), .ZN(n17913) );
  OAI21_X1 U20968 ( .B1(n17900), .B2(n17899), .A(n17898), .ZN(n18204) );
  OAI22_X1 U20969 ( .A1(n17924), .A2(n17901), .B1(n17942), .B2(n18204), .ZN(
        n17902) );
  AOI21_X1 U20970 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17913), .A(
        n17902), .ZN(n17903) );
  OAI211_X1 U20971 ( .C1(n18373), .C2(n17905), .A(n17904), .B(n17903), .ZN(
        P3_U2826) );
  AOI21_X1 U20972 ( .B1(n17908), .B2(n17907), .A(n17906), .ZN(n18214) );
  OAI21_X1 U20973 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17910), .A(
        n17909), .ZN(n18219) );
  OAI22_X1 U20974 ( .A1(n17942), .A2(n18219), .B1(n18236), .B2(n21123), .ZN(
        n17911) );
  AOI21_X1 U20975 ( .B1(n9653), .B2(n18214), .A(n17911), .ZN(n17915) );
  NOR2_X1 U20976 ( .A1(n17912), .A2(n17927), .ZN(n17928) );
  OAI21_X1 U20977 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17928), .A(
        n17913), .ZN(n17914) );
  OAI211_X1 U20978 ( .C1(n17924), .C2(n17916), .A(n17915), .B(n17914), .ZN(
        P3_U2827) );
  AOI21_X1 U20979 ( .B1(n17919), .B2(n17918), .A(n17917), .ZN(n18228) );
  NOR2_X1 U20980 ( .A1(n18236), .A2(n18809), .ZN(n18233) );
  OAI21_X1 U20981 ( .B1(n17922), .B2(n17921), .A(n17920), .ZN(n18235) );
  OAI22_X1 U20982 ( .A1(n17924), .A2(n17923), .B1(n17942), .B2(n18235), .ZN(
        n17925) );
  AOI211_X1 U20983 ( .C1(n17932), .C2(n18228), .A(n18233), .B(n17925), .ZN(
        n17926) );
  OAI221_X1 U20984 ( .B1(n17928), .B2(n17927), .C1(n17928), .C2(n18373), .A(
        n17926), .ZN(P3_U2828) );
  OAI21_X1 U20985 ( .B1(n17930), .B2(n9674), .A(n17929), .ZN(n18247) );
  NAND2_X1 U20986 ( .A1(n18886), .A2(n17937), .ZN(n17931) );
  XNOR2_X1 U20987 ( .A(n17931), .B(n17930), .ZN(n18240) );
  AOI22_X1 U20988 ( .A1(n9653), .A2(n18240), .B1(n18151), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17936) );
  AOI22_X1 U20989 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17934), .B1(
        n17725), .B2(n17933), .ZN(n17935) );
  OAI211_X1 U20990 ( .C1(n17942), .C2(n18247), .A(n17936), .B(n17935), .ZN(
        P3_U2829) );
  AOI21_X1 U20991 ( .B1(n17937), .B2(n18886), .A(n9674), .ZN(n18259) );
  INV_X1 U20992 ( .A(n18259), .ZN(n18257) );
  NAND3_X1 U20993 ( .A1(n18905), .A2(n17939), .A3(n17938), .ZN(n17940) );
  AOI22_X1 U20994 ( .A1(n18252), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17940), .ZN(n17941) );
  OAI221_X1 U20995 ( .B1(n18259), .B2(n17943), .C1(n18257), .C2(n17942), .A(
        n17941), .ZN(P3_U2830) );
  NOR2_X1 U20996 ( .A1(n17944), .A2(n18010), .ZN(n17995) );
  INV_X1 U20997 ( .A(n17995), .ZN(n17960) );
  AOI221_X1 U20998 ( .B1(n17946), .B2(n17945), .C1(n17960), .C2(n17945), .A(
        n18242), .ZN(n17956) );
  NOR2_X1 U20999 ( .A1(n18065), .A2(n18718), .ZN(n18243) );
  INV_X1 U21000 ( .A(n18243), .ZN(n17953) );
  AND2_X1 U21001 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17970) );
  NAND2_X1 U21002 ( .A1(n18065), .A2(n18886), .ZN(n18201) );
  INV_X1 U21003 ( .A(n18201), .ZN(n18221) );
  NOR2_X1 U21004 ( .A1(n18749), .A2(n18065), .ZN(n18050) );
  INV_X1 U21005 ( .A(n18050), .ZN(n18220) );
  OAI21_X1 U21006 ( .B1(n18221), .B2(n17947), .A(n18220), .ZN(n17983) );
  OAI211_X1 U21007 ( .C1(n18006), .C2(n17970), .A(n17989), .B(n17983), .ZN(
        n17971) );
  AOI21_X1 U21008 ( .B1(n18749), .B2(n17948), .A(n18126), .ZN(n17949) );
  OAI22_X1 U21009 ( .A1(n17951), .A2(n17985), .B1(n17950), .B2(n17949), .ZN(
        n17952) );
  OAI211_X1 U21010 ( .C1(n18249), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17962), .ZN(n17955) );
  AOI22_X1 U21011 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18244), .B1(
        n17956), .B2(n17955), .ZN(n17958) );
  NAND2_X1 U21012 ( .A1(n18252), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17957) );
  OAI211_X1 U21013 ( .C1(n17959), .C2(n18172), .A(n17958), .B(n17957), .ZN(
        P3_U2835) );
  NOR2_X1 U21014 ( .A1(n18242), .A2(n17960), .ZN(n17964) );
  NOR2_X1 U21015 ( .A1(n18236), .A2(n18856), .ZN(n17963) );
  NOR2_X1 U21016 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17967), .ZN(
        n17969) );
  AOI22_X1 U21017 ( .A1(n17970), .A2(n17969), .B1(n18126), .B2(n17968), .ZN(
        n17974) );
  AOI22_X1 U21018 ( .A1(n18716), .A2(n17972), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17971), .ZN(n17973) );
  AOI21_X1 U21019 ( .B1(n17974), .B2(n17973), .A(n18242), .ZN(n17975) );
  AOI21_X1 U21020 ( .B1(n18244), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17975), .ZN(n17977) );
  OAI211_X1 U21021 ( .C1(n17978), .C2(n18172), .A(n17977), .B(n17976), .ZN(
        P3_U2837) );
  AOI21_X1 U21022 ( .B1(n17980), .B2(n18016), .A(n17979), .ZN(n17992) );
  OAI21_X1 U21023 ( .B1(n18166), .B2(n17981), .A(n18211), .ZN(n17982) );
  INV_X1 U21024 ( .A(n17982), .ZN(n17984) );
  OAI211_X1 U21025 ( .C1(n17986), .C2(n17985), .A(n17984), .B(n17983), .ZN(
        n17990) );
  NOR2_X1 U21026 ( .A1(n17987), .A2(n17990), .ZN(n17988) );
  AOI21_X1 U21027 ( .B1(n17989), .B2(n17988), .A(n18252), .ZN(n17994) );
  OAI211_X1 U21028 ( .C1(n18161), .C2(n17990), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17994), .ZN(n17991) );
  OAI211_X1 U21029 ( .C1(n17993), .C2(n18172), .A(n17992), .B(n17991), .ZN(
        P3_U2838) );
  OAI221_X1 U21030 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17995), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18211), .A(n17994), .ZN(
        n17996) );
  OAI211_X1 U21031 ( .C1(n17998), .C2(n18172), .A(n17997), .B(n17996), .ZN(
        P3_U2839) );
  OAI21_X1 U21032 ( .B1(n18064), .B2(n18017), .A(n18065), .ZN(n18002) );
  OAI21_X1 U21033 ( .B1(n18045), .B2(n18017), .A(n18718), .ZN(n18001) );
  AOI21_X1 U21034 ( .B1(n18044), .B2(n18030), .A(n18249), .ZN(n17999) );
  INV_X1 U21035 ( .A(n17999), .ZN(n18000) );
  NAND3_X1 U21036 ( .A1(n18002), .A2(n18001), .A3(n18000), .ZN(n18020) );
  AOI22_X1 U21037 ( .A1(n18716), .A2(n18075), .B1(n18126), .B2(n18077), .ZN(
        n18019) );
  NOR2_X1 U21038 ( .A1(n18716), .A2(n18126), .ZN(n18130) );
  OAI222_X1 U21039 ( .A1(n18004), .A2(n18130), .B1(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n18249), .C1(n18243), .C2(
        n18003), .ZN(n18005) );
  INV_X1 U21040 ( .A(n18005), .ZN(n18022) );
  OAI211_X1 U21041 ( .C1(n18006), .C2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n18019), .B(n18022), .ZN(n18007) );
  OAI21_X1 U21042 ( .B1(n18020), .B2(n18007), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18008) );
  OAI21_X1 U21043 ( .B1(n18010), .B2(n18009), .A(n18008), .ZN(n18012) );
  AOI22_X1 U21044 ( .A1(n18248), .A2(n18012), .B1(n18070), .B2(n18011), .ZN(
        n18014) );
  OAI211_X1 U21045 ( .C1(n18211), .C2(n18015), .A(n18014), .B(n18013), .ZN(
        P3_U2840) );
  INV_X1 U21046 ( .A(n18016), .ZN(n18018) );
  NOR2_X1 U21047 ( .A1(n18018), .A2(n18017), .ZN(n18036) );
  NAND2_X1 U21048 ( .A1(n18248), .A2(n18019), .ZN(n18068) );
  NOR2_X1 U21049 ( .A1(n18068), .A2(n18020), .ZN(n18029) );
  AOI211_X1 U21050 ( .C1(n18029), .C2(n18022), .A(n18252), .B(n18021), .ZN(
        n18023) );
  AOI21_X1 U21051 ( .B1(n18036), .B2(n18024), .A(n18023), .ZN(n18026) );
  OAI211_X1 U21052 ( .C1(n18027), .C2(n18172), .A(n18026), .B(n18025), .ZN(
        P3_U2841) );
  AOI22_X1 U21053 ( .A1(n18252), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18036), 
        .B2(n18028), .ZN(n18033) );
  AOI221_X1 U21054 ( .B1(n18030), .B2(n18029), .C1(n18130), .C2(n18029), .A(
        n18252), .ZN(n18037) );
  NOR3_X1 U21055 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18243), .A3(
        n18930), .ZN(n18031) );
  OAI21_X1 U21056 ( .B1(n18037), .B2(n18031), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18032) );
  OAI211_X1 U21057 ( .C1(n18172), .C2(n18034), .A(n18033), .B(n18032), .ZN(
        P3_U2842) );
  AOI22_X1 U21058 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18037), .B1(
        n18036), .B2(n18035), .ZN(n18039) );
  NAND2_X1 U21059 ( .A1(n18252), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18038) );
  OAI211_X1 U21060 ( .C1(n18040), .C2(n18172), .A(n18039), .B(n18038), .ZN(
        P3_U2843) );
  INV_X1 U21061 ( .A(n18041), .ZN(n18042) );
  NAND2_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18200) );
  OAI22_X1 U21063 ( .A1(n18229), .A2(n18742), .B1(n18225), .B2(n18200), .ZN(
        n18216) );
  NAND2_X1 U21064 ( .A1(n18187), .A2(n18216), .ZN(n18176) );
  NOR3_X1 U21065 ( .A1(n18177), .A2(n18186), .A3(n18176), .ZN(n18163) );
  NAND2_X1 U21066 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18163), .ZN(
        n18090) );
  NAND2_X1 U21067 ( .A1(n18043), .A2(n18150), .ZN(n18074) );
  NAND3_X1 U21068 ( .A1(n18044), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18201), .ZN(n18049) );
  NAND2_X1 U21069 ( .A1(n18718), .A2(n18045), .ZN(n18046) );
  AOI22_X1 U21070 ( .A1(n18047), .A2(n18046), .B1(n18130), .B2(n18742), .ZN(
        n18048) );
  AOI211_X1 U21071 ( .C1(n18220), .C2(n18049), .A(n18048), .B(n18068), .ZN(
        n18057) );
  AOI221_X1 U21072 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18057), 
        .C1(n18050), .C2(n18057), .A(n18252), .ZN(n18052) );
  AOI22_X1 U21073 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18052), .B1(
        n18070), .B2(n18051), .ZN(n18054) );
  OAI211_X1 U21074 ( .C1(n18055), .C2(n18074), .A(n18054), .B(n18053), .ZN(
        P3_U2844) );
  NOR3_X1 U21075 ( .A1(n18252), .A2(n18057), .A3(n18056), .ZN(n18058) );
  AOI211_X1 U21076 ( .C1(n18070), .C2(n18060), .A(n18059), .B(n18058), .ZN(
        n18061) );
  OAI21_X1 U21077 ( .B1(n18074), .B2(n18062), .A(n18061), .ZN(P3_U2845) );
  INV_X1 U21078 ( .A(n18140), .ZN(n18112) );
  NOR2_X1 U21079 ( .A1(n18063), .A2(n18742), .ZN(n18133) );
  NOR2_X1 U21080 ( .A1(n18249), .A2(n18093), .ZN(n18141) );
  NOR2_X1 U21081 ( .A1(n18133), .A2(n18141), .ZN(n18152) );
  OAI21_X1 U21082 ( .B1(n18081), .B2(n18065), .A(n18064), .ZN(n18066) );
  OAI211_X1 U21083 ( .C1(n18112), .C2(n18067), .A(n18152), .B(n18066), .ZN(
        n18084) );
  OAI221_X1 U21084 ( .B1(n18068), .B2(n18161), .C1(n18068), .C2(n18084), .A(
        n18236), .ZN(n18072) );
  AOI22_X1 U21085 ( .A1(n18252), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18070), 
        .B2(n18069), .ZN(n18071) );
  OAI221_X1 U21086 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18074), 
        .C1(n18073), .C2(n18072), .A(n18071), .ZN(P3_U2846) );
  AND2_X1 U21087 ( .A1(n18075), .A2(n18716), .ZN(n18076) );
  AOI22_X1 U21088 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18244), .B1(
        n18248), .B2(n18076), .ZN(n18088) );
  NAND2_X1 U21089 ( .A1(n18126), .A2(n18077), .ZN(n18079) );
  OAI22_X1 U21090 ( .A1(n18080), .A2(n18079), .B1(n18099), .B2(n18078), .ZN(
        n18085) );
  OAI21_X1 U21091 ( .B1(n18082), .B2(n18090), .A(n18081), .ZN(n18083) );
  OAI221_X1 U21092 ( .B1(n18085), .B2(n18084), .C1(n18085), .C2(n18083), .A(
        n18248), .ZN(n18087) );
  OAI211_X1 U21093 ( .C1(n18089), .C2(n18088), .A(n18087), .B(n18086), .ZN(
        P3_U2847) );
  NOR2_X1 U21094 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18090), .ZN(
        n18092) );
  AOI22_X1 U21095 ( .A1(n18095), .A2(n18092), .B1(n18126), .B2(n18091), .ZN(
        n18098) );
  AND2_X1 U21096 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18093), .ZN(
        n18129) );
  OAI221_X1 U21097 ( .B1(n18745), .B2(n18094), .C1(n18745), .C2(n18129), .A(
        n18152), .ZN(n18110) );
  OAI22_X1 U21098 ( .A1(n18112), .A2(n18095), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18243), .ZN(n18096) );
  OAI21_X1 U21099 ( .B1(n18110), .B2(n18096), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18097) );
  OAI211_X1 U21100 ( .C1(n18100), .C2(n18099), .A(n18098), .B(n18097), .ZN(
        n18102) );
  AOI22_X1 U21101 ( .A1(n18248), .A2(n18102), .B1(n18241), .B2(n18101), .ZN(
        n18105) );
  INV_X1 U21102 ( .A(n18103), .ZN(n18104) );
  OAI211_X1 U21103 ( .C1(n18211), .C2(n18106), .A(n18105), .B(n18104), .ZN(
        P3_U2848) );
  AOI22_X1 U21104 ( .A1(n18252), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18150), 
        .B2(n18107), .ZN(n18115) );
  OAI22_X1 U21105 ( .A1(n18112), .A2(n18117), .B1(n18108), .B2(n18166), .ZN(
        n18109) );
  AOI211_X1 U21106 ( .C1(n18716), .C2(n18111), .A(n18110), .B(n18109), .ZN(
        n18119) );
  OAI211_X1 U21107 ( .C1(n18112), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18248), .B(n18119), .ZN(n18113) );
  NAND3_X1 U21108 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18236), .A3(
        n18113), .ZN(n18114) );
  OAI211_X1 U21109 ( .C1(n18116), .C2(n18172), .A(n18115), .B(n18114), .ZN(
        P3_U2849) );
  AOI22_X1 U21110 ( .A1(n18117), .A2(n18150), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18248), .ZN(n18118) );
  AOI21_X1 U21111 ( .B1(n18119), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18118), .ZN(n18120) );
  AOI21_X1 U21112 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18244), .A(
        n18120), .ZN(n18122) );
  OAI211_X1 U21113 ( .C1(n18123), .C2(n18172), .A(n18122), .B(n18121), .ZN(
        P3_U2850) );
  AOI22_X1 U21114 ( .A1(n18252), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18150), 
        .B2(n18124), .ZN(n18138) );
  AOI22_X1 U21115 ( .A1(n18716), .A2(n18127), .B1(n18126), .B2(n18125), .ZN(
        n18128) );
  OAI211_X1 U21116 ( .C1(n18745), .C2(n18129), .A(n18248), .B(n18128), .ZN(
        n18153) );
  OAI22_X1 U21117 ( .A1(n18745), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n18131), .B2(n18130), .ZN(n18132) );
  NOR3_X1 U21118 ( .A1(n18133), .A2(n18153), .A3(n18132), .ZN(n18143) );
  NAND2_X1 U21119 ( .A1(n18140), .A2(n18134), .ZN(n18135) );
  OAI211_X1 U21120 ( .C1(n18745), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18143), .B(n18135), .ZN(n18136) );
  OAI211_X1 U21121 ( .C1(n18141), .C2(n18136), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18236), .ZN(n18137) );
  OAI211_X1 U21122 ( .C1(n18139), .C2(n18172), .A(n18138), .B(n18137), .ZN(
        P3_U2851) );
  OAI21_X1 U21123 ( .B1(n18141), .B2(n18149), .A(n18140), .ZN(n18142) );
  AOI21_X1 U21124 ( .B1(n18143), .B2(n18142), .A(n18151), .ZN(n18144) );
  AOI22_X1 U21125 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18144), .B1(
        n18151), .B2(P3_REIP_REG_10__SCAN_IN), .ZN(n18147) );
  NAND3_X1 U21126 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18150), .A3(
        n18145), .ZN(n18146) );
  OAI211_X1 U21127 ( .C1(n18148), .C2(n18172), .A(n18147), .B(n18146), .ZN(
        P3_U2852) );
  AOI22_X1 U21128 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18151), .B1(n18150), 
        .B2(n18149), .ZN(n18156) );
  INV_X1 U21129 ( .A(n18152), .ZN(n18154) );
  OAI211_X1 U21130 ( .C1(n18154), .C2(n18153), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18236), .ZN(n18155) );
  OAI211_X1 U21131 ( .C1(n18157), .C2(n18172), .A(n18156), .B(n18155), .ZN(
        P3_U2853) );
  AOI22_X1 U21132 ( .A1(n18718), .A2(n18159), .B1(n18220), .B2(n18158), .ZN(
        n18160) );
  NAND2_X1 U21133 ( .A1(n18160), .A2(n18201), .ZN(n18183) );
  AOI211_X1 U21134 ( .C1(n18161), .C2(n18186), .A(n18177), .B(n18183), .ZN(
        n18175) );
  OAI21_X1 U21135 ( .B1(n18175), .B2(n18237), .A(n18211), .ZN(n18169) );
  AOI22_X1 U21136 ( .A1(n18716), .A2(n18164), .B1(n18163), .B2(n18162), .ZN(
        n18165) );
  OAI21_X1 U21137 ( .B1(n18167), .B2(n18166), .A(n18165), .ZN(n18168) );
  AOI22_X1 U21138 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18169), .B1(
        n18248), .B2(n18168), .ZN(n18171) );
  OAI211_X1 U21139 ( .C1(n18173), .C2(n18172), .A(n18171), .B(n18170), .ZN(
        P3_U2854) );
  AOI21_X1 U21140 ( .B1(n18244), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18174), .ZN(n18181) );
  AOI221_X1 U21141 ( .B1(n18186), .B2(n18177), .C1(n18176), .C2(n18177), .A(
        n18175), .ZN(n18179) );
  AOI22_X1 U21142 ( .A1(n18248), .A2(n18179), .B1(n18241), .B2(n18178), .ZN(
        n18180) );
  OAI211_X1 U21143 ( .C1(n18256), .C2(n18182), .A(n18181), .B(n18180), .ZN(
        P3_U2855) );
  OAI21_X1 U21144 ( .B1(n18242), .B2(n18183), .A(n18236), .ZN(n18191) );
  OAI22_X1 U21145 ( .A1(n18186), .A2(n18191), .B1(n18236), .B2(n18816), .ZN(
        n18184) );
  AOI21_X1 U21146 ( .B1(n18241), .B2(n18185), .A(n18184), .ZN(n18189) );
  NAND4_X1 U21147 ( .A1(n18248), .A2(n18187), .A3(n18186), .A4(n18216), .ZN(
        n18188) );
  OAI211_X1 U21148 ( .C1(n18190), .C2(n18256), .A(n18189), .B(n18188), .ZN(
        P3_U2856) );
  NAND4_X1 U21149 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18248), .A4(n18216), .ZN(
        n18199) );
  OAI22_X1 U21150 ( .A1(n18192), .A2(n18191), .B1(n18236), .B2(n18815), .ZN(
        n18193) );
  INV_X1 U21151 ( .A(n18193), .ZN(n18198) );
  AOI22_X1 U21152 ( .A1(n18196), .A2(n18195), .B1(n18241), .B2(n18194), .ZN(
        n18197) );
  OAI211_X1 U21153 ( .C1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n18199), .A(
        n18198), .B(n18197), .ZN(P3_U2857) );
  NAND3_X1 U21154 ( .A1(n18248), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18216), .ZN(n18210) );
  AOI22_X1 U21155 ( .A1(n18718), .A2(n18229), .B1(n18220), .B2(n18200), .ZN(
        n18202) );
  NAND3_X1 U21156 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18202), .A3(
        n18201), .ZN(n18215) );
  AOI21_X1 U21157 ( .B1(n18203), .B2(n18215), .A(n18244), .ZN(n18208) );
  OAI22_X1 U21158 ( .A1(n18236), .A2(n18812), .B1(n18256), .B2(n18204), .ZN(
        n18205) );
  AOI21_X1 U21159 ( .B1(n18241), .B2(n18206), .A(n18205), .ZN(n18207) );
  OAI221_X1 U21160 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18210), .C1(
        n18209), .C2(n18208), .A(n18207), .ZN(P3_U2858) );
  OAI22_X1 U21161 ( .A1(n18212), .A2(n18211), .B1(n18236), .B2(n21123), .ZN(
        n18213) );
  AOI21_X1 U21162 ( .B1(n18241), .B2(n18214), .A(n18213), .ZN(n18218) );
  OAI211_X1 U21163 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18216), .A(
        n18248), .B(n18215), .ZN(n18217) );
  OAI211_X1 U21164 ( .C1(n18219), .C2(n18256), .A(n18218), .B(n18217), .ZN(
        P3_U2859) );
  OAI21_X1 U21165 ( .B1(n18221), .B2(n9850), .A(n18220), .ZN(n18224) );
  NAND2_X1 U21166 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18223) );
  AOI221_X1 U21167 ( .B1(n18742), .B2(n18224), .C1(n18223), .C2(n18224), .A(
        n18222), .ZN(n18227) );
  NOR3_X1 U21168 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n9850), .A3(
        n18225), .ZN(n18226) );
  AOI211_X1 U21169 ( .C1(n18228), .C2(n18716), .A(n18227), .B(n18226), .ZN(
        n18231) );
  NAND2_X1 U21170 ( .A1(n18718), .A2(n18229), .ZN(n18230) );
  AOI21_X1 U21171 ( .B1(n18231), .B2(n18230), .A(n18242), .ZN(n18232) );
  AOI211_X1 U21172 ( .C1(n18244), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18233), .B(n18232), .ZN(n18234) );
  OAI21_X1 U21173 ( .B1(n18256), .B2(n18235), .A(n18234), .ZN(P3_U2860) );
  NOR2_X1 U21174 ( .A1(n18236), .A2(n18911), .ZN(n18239) );
  AOI211_X1 U21175 ( .C1(n18249), .C2(n18886), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18237), .ZN(n18238) );
  AOI211_X1 U21176 ( .C1(n18241), .C2(n18240), .A(n18239), .B(n18238), .ZN(
        n18246) );
  NOR3_X1 U21177 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18243), .A3(
        n18242), .ZN(n18251) );
  OAI21_X1 U21178 ( .B1(n18244), .B2(n18251), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18245) );
  OAI211_X1 U21179 ( .C1(n18247), .C2(n18256), .A(n18246), .B(n18245), .ZN(
        P3_U2861) );
  AOI21_X1 U21180 ( .B1(n18249), .B2(n18248), .A(n18886), .ZN(n18250) );
  NOR2_X1 U21181 ( .A1(n18251), .A2(n18250), .ZN(n18254) );
  INV_X1 U21182 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18253) );
  MUX2_X1 U21183 ( .A(n18254), .B(n18253), .S(n18252), .Z(n18255) );
  OAI221_X1 U21184 ( .B1(n18259), .B2(n18258), .C1(n18257), .C2(n18256), .A(
        n18255), .ZN(P3_U2862) );
  OAI211_X1 U21185 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18260), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18773)
         );
  OAI21_X1 U21186 ( .B1(n18262), .B2(n18924), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18261) );
  OAI221_X1 U21187 ( .B1(n18262), .B2(n18773), .C1(n18262), .C2(n18311), .A(
        n18261), .ZN(P3_U2863) );
  INV_X1 U21188 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18757) );
  NOR2_X1 U21189 ( .A1(n18263), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18443) );
  INV_X1 U21190 ( .A(n18443), .ZN(n18396) );
  NOR2_X1 U21191 ( .A1(n18757), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18540) );
  NAND2_X1 U21192 ( .A1(n18330), .A2(n18540), .ZN(n18562) );
  AND2_X1 U21193 ( .A1(n18396), .A2(n18562), .ZN(n18265) );
  OAI22_X1 U21194 ( .A1(n18266), .A2(n18757), .B1(n18265), .B2(n18264), .ZN(
        P3_U2866) );
  NOR2_X1 U21195 ( .A1(n18755), .A2(n18267), .ZN(P3_U2867) );
  NAND2_X1 U21196 ( .A1(n18655), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18469) );
  NAND2_X1 U21197 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18272) );
  INV_X1 U21198 ( .A(n18272), .ZN(n18270) );
  NOR2_X1 U21199 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18539), .ZN(
        n18514) );
  NAND2_X1 U21200 ( .A1(n18270), .A2(n18514), .ZN(n18624) );
  NOR2_X1 U21201 ( .A1(n18272), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18654) );
  NAND2_X1 U21202 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18654), .ZN(
        n18709) );
  INV_X1 U21203 ( .A(n18709), .ZN(n18687) );
  INV_X1 U21204 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18268) );
  NOR2_X2 U21205 ( .A1(n18268), .A2(n18373), .ZN(n18656) );
  INV_X1 U21206 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18269) );
  NOR2_X2 U21207 ( .A1(n18372), .A2(n18269), .ZN(n18650) );
  NAND2_X1 U21208 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18537) );
  INV_X1 U21209 ( .A(n18537), .ZN(n18750) );
  NAND2_X1 U21210 ( .A1(n18750), .A2(n18270), .ZN(n18660) );
  NOR2_X1 U21211 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18751) );
  NOR2_X1 U21212 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18351) );
  NAND2_X1 U21213 ( .A1(n18751), .A2(n18351), .ZN(n18371) );
  NAND2_X1 U21214 ( .A1(n18660), .A2(n18371), .ZN(n18273) );
  INV_X1 U21215 ( .A(n18273), .ZN(n18331) );
  NOR2_X1 U21216 ( .A1(n18616), .A2(n18331), .ZN(n18305) );
  AOI22_X1 U21217 ( .A1(n18687), .A2(n18656), .B1(n18650), .B2(n18305), .ZN(
        n18279) );
  NOR2_X1 U21218 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18271), .ZN(
        n18488) );
  NOR2_X1 U21219 ( .A1(n18514), .A2(n18488), .ZN(n18563) );
  NOR2_X1 U21220 ( .A1(n18563), .A2(n18272), .ZN(n18615) );
  AOI21_X1 U21221 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18372), .ZN(n18274) );
  AOI22_X1 U21222 ( .A1(n18655), .A2(n18615), .B1(n18274), .B2(n18273), .ZN(
        n18308) );
  INV_X1 U21223 ( .A(n18371), .ZN(n18364) );
  NAND2_X1 U21224 ( .A1(n18276), .A2(n18275), .ZN(n18306) );
  NOR2_X1 U21225 ( .A1(n18277), .A2(n18306), .ZN(n18466) );
  AOI22_X1 U21226 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18308), .B1(
        n18364), .B2(n18466), .ZN(n18278) );
  OAI211_X1 U21227 ( .C1(n18469), .C2(n18624), .A(n18279), .B(n18278), .ZN(
        P3_U2868) );
  NOR2_X1 U21228 ( .A1(n18280), .A2(n18373), .ZN(n18591) );
  INV_X1 U21229 ( .A(n18591), .ZN(n18666) );
  INV_X1 U21230 ( .A(n18624), .ZN(n18644) );
  AND2_X1 U21231 ( .A1(n18655), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18662) );
  AND2_X1 U21232 ( .A1(n18621), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18661) );
  AOI22_X1 U21233 ( .A1(n18644), .A2(n18662), .B1(n18305), .B2(n18661), .ZN(
        n18283) );
  NOR2_X1 U21234 ( .A1(n18281), .A2(n18306), .ZN(n18663) );
  AOI22_X1 U21235 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18308), .B1(
        n18364), .B2(n18663), .ZN(n18282) );
  OAI211_X1 U21236 ( .C1(n18709), .C2(n18666), .A(n18283), .B(n18282), .ZN(
        P3_U2869) );
  NAND2_X1 U21237 ( .A1(n18655), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18631) );
  NAND2_X1 U21238 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18655), .ZN(n18672) );
  INV_X1 U21239 ( .A(n18672), .ZN(n18628) );
  NOR2_X2 U21240 ( .A1(n18372), .A2(n18284), .ZN(n18667) );
  AOI22_X1 U21241 ( .A1(n18687), .A2(n18628), .B1(n18305), .B2(n18667), .ZN(
        n18287) );
  AOI22_X1 U21242 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18308), .B1(
        n18364), .B2(n18669), .ZN(n18286) );
  OAI211_X1 U21243 ( .C1(n18624), .C2(n18631), .A(n18287), .B(n18286), .ZN(
        P3_U2870) );
  NAND2_X1 U21244 ( .A1(n18655), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18600) );
  NAND2_X1 U21245 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18655), .ZN(n18678) );
  INV_X1 U21246 ( .A(n18678), .ZN(n18597) );
  NOR2_X2 U21247 ( .A1(n18372), .A2(n18288), .ZN(n18673) );
  AOI22_X1 U21248 ( .A1(n18687), .A2(n18597), .B1(n18305), .B2(n18673), .ZN(
        n18291) );
  NOR2_X1 U21249 ( .A1(n18289), .A2(n18306), .ZN(n18675) );
  AOI22_X1 U21250 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18308), .B1(
        n18364), .B2(n18675), .ZN(n18290) );
  OAI211_X1 U21251 ( .C1(n18624), .C2(n18600), .A(n18291), .B(n18290), .ZN(
        P3_U2871) );
  NAND2_X1 U21252 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18655), .ZN(n18684) );
  NAND2_X1 U21253 ( .A1(n18655), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18576) );
  INV_X1 U21254 ( .A(n18576), .ZN(n18680) );
  NOR2_X2 U21255 ( .A1(n18372), .A2(n18292), .ZN(n18679) );
  AOI22_X1 U21256 ( .A1(n18644), .A2(n18680), .B1(n18305), .B2(n18679), .ZN(
        n18295) );
  NOR2_X2 U21257 ( .A1(n18293), .A2(n18306), .ZN(n18681) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18308), .B1(
        n18364), .B2(n18681), .ZN(n18294) );
  OAI211_X1 U21259 ( .C1(n18709), .C2(n18684), .A(n18295), .B(n18294), .ZN(
        P3_U2872) );
  NOR2_X1 U21260 ( .A1(n18373), .A2(n19405), .ZN(n18686) );
  INV_X1 U21261 ( .A(n18686), .ZN(n18606) );
  NAND2_X1 U21262 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18655), .ZN(n18692) );
  INV_X1 U21263 ( .A(n18692), .ZN(n18603) );
  NOR2_X2 U21264 ( .A1(n18372), .A2(n18296), .ZN(n18685) );
  AOI22_X1 U21265 ( .A1(n18687), .A2(n18603), .B1(n18305), .B2(n18685), .ZN(
        n18299) );
  NOR2_X2 U21266 ( .A1(n18297), .A2(n18306), .ZN(n18688) );
  AOI22_X1 U21267 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18308), .B1(
        n18364), .B2(n18688), .ZN(n18298) );
  OAI211_X1 U21268 ( .C1(n18624), .C2(n18606), .A(n18299), .B(n18298), .ZN(
        P3_U2873) );
  NAND2_X1 U21269 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18655), .ZN(n18641) );
  NAND2_X1 U21270 ( .A1(n18655), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18698) );
  INV_X1 U21271 ( .A(n18698), .ZN(n18638) );
  NOR2_X2 U21272 ( .A1(n18372), .A2(n18300), .ZN(n18693) );
  AOI22_X1 U21273 ( .A1(n18644), .A2(n18638), .B1(n18305), .B2(n18693), .ZN(
        n18303) );
  NOR2_X2 U21274 ( .A1(n18301), .A2(n18306), .ZN(n18695) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18308), .B1(
        n18364), .B2(n18695), .ZN(n18302) );
  OAI211_X1 U21276 ( .C1(n18709), .C2(n18641), .A(n18303), .B(n18302), .ZN(
        P3_U2874) );
  NOR2_X1 U21277 ( .A1(n18373), .A2(n19418), .ZN(n18702) );
  INV_X1 U21278 ( .A(n18702), .ZN(n18649) );
  NAND2_X1 U21279 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18655), .ZN(n18708) );
  INV_X1 U21280 ( .A(n18708), .ZN(n18643) );
  NOR2_X2 U21281 ( .A1(n18304), .A2(n18372), .ZN(n18700) );
  AOI22_X1 U21282 ( .A1(n18644), .A2(n18643), .B1(n18305), .B2(n18700), .ZN(
        n18310) );
  NOR2_X2 U21283 ( .A1(n18307), .A2(n18306), .ZN(n18703) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18308), .B1(
        n18364), .B2(n18703), .ZN(n18309) );
  OAI211_X1 U21285 ( .C1(n18709), .C2(n18649), .A(n18310), .B(n18309), .ZN(
        P3_U2875) );
  INV_X1 U21286 ( .A(n18466), .ZN(n18659) );
  NAND2_X1 U21287 ( .A1(n18488), .A2(n18351), .ZN(n18386) );
  INV_X1 U21288 ( .A(n18660), .ZN(n18704) );
  INV_X1 U21289 ( .A(n18469), .ZN(n18651) );
  INV_X1 U21290 ( .A(n18351), .ZN(n18397) );
  NAND2_X1 U21291 ( .A1(n18539), .A2(n18776), .ZN(n18489) );
  NOR2_X1 U21292 ( .A1(n18397), .A2(n18489), .ZN(n18326) );
  AOI22_X1 U21293 ( .A1(n18704), .A2(n18651), .B1(n18650), .B2(n18326), .ZN(
        n18313) );
  NOR2_X1 U21294 ( .A1(n18757), .A2(n18490), .ZN(n18652) );
  NAND2_X1 U21295 ( .A1(n18621), .A2(n18311), .ZN(n18491) );
  NOR2_X1 U21296 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18491), .ZN(
        n18398) );
  AOI22_X1 U21297 ( .A1(n18655), .A2(n18652), .B1(n18351), .B2(n18398), .ZN(
        n18327) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18327), .B1(
        n18644), .B2(n18656), .ZN(n18312) );
  OAI211_X1 U21299 ( .C1(n18659), .C2(n18386), .A(n18313), .B(n18312), .ZN(
        P3_U2876) );
  INV_X1 U21300 ( .A(n18663), .ZN(n18594) );
  AOI22_X1 U21301 ( .A1(n18644), .A2(n18591), .B1(n18661), .B2(n18326), .ZN(
        n18315) );
  AOI22_X1 U21302 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18327), .B1(
        n18704), .B2(n18662), .ZN(n18314) );
  OAI211_X1 U21303 ( .C1(n18594), .C2(n18386), .A(n18315), .B(n18314), .ZN(
        P3_U2877) );
  AOI22_X1 U21304 ( .A1(n18644), .A2(n18628), .B1(n18667), .B2(n18326), .ZN(
        n18317) );
  INV_X1 U21305 ( .A(n18386), .ZN(n18392) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18327), .B1(
        n18669), .B2(n18392), .ZN(n18316) );
  OAI211_X1 U21307 ( .C1(n18660), .C2(n18631), .A(n18317), .B(n18316), .ZN(
        P3_U2878) );
  INV_X1 U21308 ( .A(n18600), .ZN(n18674) );
  AOI22_X1 U21309 ( .A1(n18704), .A2(n18674), .B1(n18673), .B2(n18326), .ZN(
        n18319) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18327), .B1(
        n18675), .B2(n18392), .ZN(n18318) );
  OAI211_X1 U21311 ( .C1(n18624), .C2(n18678), .A(n18319), .B(n18318), .ZN(
        P3_U2879) );
  INV_X1 U21312 ( .A(n18684), .ZN(n18573) );
  AOI22_X1 U21313 ( .A1(n18644), .A2(n18573), .B1(n18679), .B2(n18326), .ZN(
        n18321) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18327), .B1(
        n18681), .B2(n18392), .ZN(n18320) );
  OAI211_X1 U21315 ( .C1(n18660), .C2(n18576), .A(n18321), .B(n18320), .ZN(
        P3_U2880) );
  AOI22_X1 U21316 ( .A1(n18644), .A2(n18603), .B1(n18685), .B2(n18326), .ZN(
        n18323) );
  AOI22_X1 U21317 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18327), .B1(
        n18688), .B2(n18392), .ZN(n18322) );
  OAI211_X1 U21318 ( .C1(n18660), .C2(n18606), .A(n18323), .B(n18322), .ZN(
        P3_U2881) );
  AOI22_X1 U21319 ( .A1(n18704), .A2(n18638), .B1(n18693), .B2(n18326), .ZN(
        n18325) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18327), .B1(
        n18695), .B2(n18392), .ZN(n18324) );
  OAI211_X1 U21321 ( .C1(n18624), .C2(n18641), .A(n18325), .B(n18324), .ZN(
        P3_U2882) );
  AOI22_X1 U21322 ( .A1(n18704), .A2(n18643), .B1(n18700), .B2(n18326), .ZN(
        n18329) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18327), .B1(
        n18703), .B2(n18392), .ZN(n18328) );
  OAI211_X1 U21324 ( .C1(n18624), .C2(n18649), .A(n18329), .B(n18328), .ZN(
        P3_U2883) );
  NAND2_X1 U21325 ( .A1(n18514), .A2(n18351), .ZN(n18414) );
  AOI21_X1 U21326 ( .B1(n18386), .B2(n18414), .A(n18616), .ZN(n18347) );
  AOI22_X1 U21327 ( .A1(n18704), .A2(n18656), .B1(n18650), .B2(n18347), .ZN(
        n18334) );
  INV_X1 U21328 ( .A(n18414), .ZN(n18416) );
  INV_X1 U21329 ( .A(n18330), .ZN(n18618) );
  AOI221_X1 U21330 ( .B1(n18331), .B2(n18386), .C1(n18618), .C2(n18386), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18332) );
  OAI21_X1 U21331 ( .B1(n18416), .B2(n18332), .A(n18621), .ZN(n18348) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18348), .B1(
        n18364), .B2(n18651), .ZN(n18333) );
  OAI211_X1 U21333 ( .C1(n18659), .C2(n18414), .A(n18334), .B(n18333), .ZN(
        P3_U2884) );
  AOI22_X1 U21334 ( .A1(n18704), .A2(n18591), .B1(n18661), .B2(n18347), .ZN(
        n18336) );
  AOI22_X1 U21335 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18348), .B1(
        n18364), .B2(n18662), .ZN(n18335) );
  OAI211_X1 U21336 ( .C1(n18594), .C2(n18414), .A(n18336), .B(n18335), .ZN(
        P3_U2885) );
  AOI22_X1 U21337 ( .A1(n18704), .A2(n18628), .B1(n18667), .B2(n18347), .ZN(
        n18338) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18348), .B1(
        n18669), .B2(n18416), .ZN(n18337) );
  OAI211_X1 U21339 ( .C1(n18371), .C2(n18631), .A(n18338), .B(n18337), .ZN(
        P3_U2886) );
  AOI22_X1 U21340 ( .A1(n18364), .A2(n18674), .B1(n18673), .B2(n18347), .ZN(
        n18340) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18348), .B1(
        n18675), .B2(n18416), .ZN(n18339) );
  OAI211_X1 U21342 ( .C1(n18660), .C2(n18678), .A(n18340), .B(n18339), .ZN(
        P3_U2887) );
  AOI22_X1 U21343 ( .A1(n18364), .A2(n18680), .B1(n18679), .B2(n18347), .ZN(
        n18342) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18348), .B1(
        n18681), .B2(n18416), .ZN(n18341) );
  OAI211_X1 U21345 ( .C1(n18660), .C2(n18684), .A(n18342), .B(n18341), .ZN(
        P3_U2888) );
  AOI22_X1 U21346 ( .A1(n18364), .A2(n18686), .B1(n18685), .B2(n18347), .ZN(
        n18344) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18348), .B1(
        n18688), .B2(n18416), .ZN(n18343) );
  OAI211_X1 U21348 ( .C1(n18660), .C2(n18692), .A(n18344), .B(n18343), .ZN(
        P3_U2889) );
  INV_X1 U21349 ( .A(n18641), .ZN(n18694) );
  AOI22_X1 U21350 ( .A1(n18704), .A2(n18694), .B1(n18693), .B2(n18347), .ZN(
        n18346) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18348), .B1(
        n18695), .B2(n18416), .ZN(n18345) );
  OAI211_X1 U21352 ( .C1(n18371), .C2(n18698), .A(n18346), .B(n18345), .ZN(
        P3_U2890) );
  AOI22_X1 U21353 ( .A1(n18364), .A2(n18643), .B1(n18700), .B2(n18347), .ZN(
        n18350) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18348), .B1(
        n18703), .B2(n18416), .ZN(n18349) );
  OAI211_X1 U21355 ( .C1(n18660), .C2(n18649), .A(n18350), .B(n18349), .ZN(
        P3_U2891) );
  AOI22_X1 U21356 ( .A1(n18364), .A2(n18656), .B1(n18650), .B2(n18367), .ZN(
        n18353) );
  AOI21_X1 U21357 ( .B1(n18539), .B2(n18618), .A(n18491), .ZN(n18442) );
  NAND2_X1 U21358 ( .A1(n18351), .A2(n18442), .ZN(n18368) );
  NAND2_X1 U21359 ( .A1(n18750), .A2(n18351), .ZN(n18441) );
  INV_X1 U21360 ( .A(n18441), .ZN(n18428) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18368), .B1(
        n18466), .B2(n18428), .ZN(n18352) );
  OAI211_X1 U21362 ( .C1(n18469), .C2(n18386), .A(n18353), .B(n18352), .ZN(
        P3_U2892) );
  AOI22_X1 U21363 ( .A1(n18662), .A2(n18392), .B1(n18661), .B2(n18367), .ZN(
        n18355) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18368), .B1(
        n18663), .B2(n18428), .ZN(n18354) );
  OAI211_X1 U21365 ( .C1(n18371), .C2(n18666), .A(n18355), .B(n18354), .ZN(
        P3_U2893) );
  AOI22_X1 U21366 ( .A1(n18364), .A2(n18628), .B1(n18667), .B2(n18367), .ZN(
        n18357) );
  AOI22_X1 U21367 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18368), .B1(
        n18669), .B2(n18428), .ZN(n18356) );
  OAI211_X1 U21368 ( .C1(n18631), .C2(n18386), .A(n18357), .B(n18356), .ZN(
        P3_U2894) );
  AOI22_X1 U21369 ( .A1(n18674), .A2(n18392), .B1(n18673), .B2(n18367), .ZN(
        n18359) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18368), .B1(
        n18675), .B2(n18428), .ZN(n18358) );
  OAI211_X1 U21371 ( .C1(n18371), .C2(n18678), .A(n18359), .B(n18358), .ZN(
        P3_U2895) );
  AOI22_X1 U21372 ( .A1(n18680), .A2(n18392), .B1(n18679), .B2(n18367), .ZN(
        n18361) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18368), .B1(
        n18681), .B2(n18428), .ZN(n18360) );
  OAI211_X1 U21374 ( .C1(n18371), .C2(n18684), .A(n18361), .B(n18360), .ZN(
        P3_U2896) );
  AOI22_X1 U21375 ( .A1(n18686), .A2(n18392), .B1(n18685), .B2(n18367), .ZN(
        n18363) );
  AOI22_X1 U21376 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18368), .B1(
        n18688), .B2(n18428), .ZN(n18362) );
  OAI211_X1 U21377 ( .C1(n18371), .C2(n18692), .A(n18363), .B(n18362), .ZN(
        P3_U2897) );
  AOI22_X1 U21378 ( .A1(n18364), .A2(n18694), .B1(n18693), .B2(n18367), .ZN(
        n18366) );
  AOI22_X1 U21379 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18368), .B1(
        n18695), .B2(n18428), .ZN(n18365) );
  OAI211_X1 U21380 ( .C1(n18698), .C2(n18386), .A(n18366), .B(n18365), .ZN(
        P3_U2898) );
  AOI22_X1 U21381 ( .A1(n18643), .A2(n18392), .B1(n18700), .B2(n18367), .ZN(
        n18370) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18368), .B1(
        n18703), .B2(n18428), .ZN(n18369) );
  OAI211_X1 U21383 ( .C1(n18371), .C2(n18649), .A(n18370), .B(n18369), .ZN(
        P3_U2899) );
  NAND2_X1 U21384 ( .A1(n18751), .A2(n18443), .ZN(n18463) );
  NOR2_X1 U21385 ( .A1(n18428), .A2(n18456), .ZN(n18420) );
  NOR2_X1 U21386 ( .A1(n18616), .A2(n18420), .ZN(n18391) );
  AOI22_X1 U21387 ( .A1(n18656), .A2(n18392), .B1(n18650), .B2(n18391), .ZN(
        n18377) );
  NOR2_X1 U21388 ( .A1(n18392), .A2(n18416), .ZN(n18374) );
  OAI22_X1 U21389 ( .A1(n18374), .A2(n18373), .B1(n18420), .B2(n18372), .ZN(
        n18375) );
  OAI21_X1 U21390 ( .B1(n18456), .B2(n18878), .A(n18375), .ZN(n18393) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18393), .B1(
        n18466), .B2(n18456), .ZN(n18376) );
  OAI211_X1 U21392 ( .C1(n18469), .C2(n18414), .A(n18377), .B(n18376), .ZN(
        P3_U2900) );
  AOI22_X1 U21393 ( .A1(n18662), .A2(n18416), .B1(n18661), .B2(n18391), .ZN(
        n18379) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18393), .B1(
        n18663), .B2(n18456), .ZN(n18378) );
  OAI211_X1 U21395 ( .C1(n18666), .C2(n18386), .A(n18379), .B(n18378), .ZN(
        P3_U2901) );
  INV_X1 U21396 ( .A(n18631), .ZN(n18668) );
  AOI22_X1 U21397 ( .A1(n18668), .A2(n18416), .B1(n18667), .B2(n18391), .ZN(
        n18381) );
  AOI22_X1 U21398 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18393), .B1(
        n18669), .B2(n18456), .ZN(n18380) );
  OAI211_X1 U21399 ( .C1(n18672), .C2(n18386), .A(n18381), .B(n18380), .ZN(
        P3_U2902) );
  AOI22_X1 U21400 ( .A1(n18674), .A2(n18416), .B1(n18673), .B2(n18391), .ZN(
        n18383) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18393), .B1(
        n18675), .B2(n18456), .ZN(n18382) );
  OAI211_X1 U21402 ( .C1(n18678), .C2(n18386), .A(n18383), .B(n18382), .ZN(
        P3_U2903) );
  AOI22_X1 U21403 ( .A1(n18680), .A2(n18416), .B1(n18679), .B2(n18391), .ZN(
        n18385) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18393), .B1(
        n18681), .B2(n18456), .ZN(n18384) );
  OAI211_X1 U21405 ( .C1(n18684), .C2(n18386), .A(n18385), .B(n18384), .ZN(
        P3_U2904) );
  AOI22_X1 U21406 ( .A1(n18603), .A2(n18392), .B1(n18685), .B2(n18391), .ZN(
        n18388) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18393), .B1(
        n18688), .B2(n18456), .ZN(n18387) );
  OAI211_X1 U21408 ( .C1(n18606), .C2(n18414), .A(n18388), .B(n18387), .ZN(
        P3_U2905) );
  AOI22_X1 U21409 ( .A1(n18694), .A2(n18392), .B1(n18693), .B2(n18391), .ZN(
        n18390) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18393), .B1(
        n18695), .B2(n18456), .ZN(n18389) );
  OAI211_X1 U21411 ( .C1(n18698), .C2(n18414), .A(n18390), .B(n18389), .ZN(
        P3_U2906) );
  AOI22_X1 U21412 ( .A1(n18702), .A2(n18392), .B1(n18700), .B2(n18391), .ZN(
        n18395) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18393), .B1(
        n18703), .B2(n18456), .ZN(n18394) );
  OAI211_X1 U21414 ( .C1(n18708), .C2(n18414), .A(n18395), .B(n18394), .ZN(
        P3_U2907) );
  NAND2_X1 U21415 ( .A1(n18488), .A2(n18443), .ZN(n18482) );
  NOR2_X1 U21416 ( .A1(n18489), .A2(n18396), .ZN(n18415) );
  AOI22_X1 U21417 ( .A1(n18656), .A2(n18416), .B1(n18650), .B2(n18415), .ZN(
        n18401) );
  NOR2_X1 U21418 ( .A1(n18539), .A2(n18397), .ZN(n18399) );
  AOI22_X1 U21419 ( .A1(n18655), .A2(n18399), .B1(n18398), .B2(n18443), .ZN(
        n18417) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18417), .B1(
        n18651), .B2(n18428), .ZN(n18400) );
  OAI211_X1 U21421 ( .C1(n18659), .C2(n18482), .A(n18401), .B(n18400), .ZN(
        P3_U2908) );
  AOI22_X1 U21422 ( .A1(n18591), .A2(n18416), .B1(n18661), .B2(n18415), .ZN(
        n18403) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18417), .B1(
        n18662), .B2(n18428), .ZN(n18402) );
  OAI211_X1 U21424 ( .C1(n18594), .C2(n18482), .A(n18403), .B(n18402), .ZN(
        P3_U2909) );
  INV_X1 U21425 ( .A(n18669), .ZN(n18548) );
  AOI22_X1 U21426 ( .A1(n18628), .A2(n18416), .B1(n18667), .B2(n18415), .ZN(
        n18405) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18417), .B1(
        n18668), .B2(n18428), .ZN(n18404) );
  OAI211_X1 U21428 ( .C1(n18548), .C2(n18482), .A(n18405), .B(n18404), .ZN(
        P3_U2910) );
  INV_X1 U21429 ( .A(n18675), .ZN(n18551) );
  AOI22_X1 U21430 ( .A1(n18597), .A2(n18416), .B1(n18673), .B2(n18415), .ZN(
        n18407) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18417), .B1(
        n18674), .B2(n18428), .ZN(n18406) );
  OAI211_X1 U21432 ( .C1(n18551), .C2(n18482), .A(n18407), .B(n18406), .ZN(
        P3_U2911) );
  AOI22_X1 U21433 ( .A1(n18680), .A2(n18428), .B1(n18679), .B2(n18415), .ZN(
        n18409) );
  INV_X1 U21434 ( .A(n18482), .ZN(n18484) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18417), .B1(
        n18681), .B2(n18484), .ZN(n18408) );
  OAI211_X1 U21436 ( .C1(n18684), .C2(n18414), .A(n18409), .B(n18408), .ZN(
        P3_U2912) );
  AOI22_X1 U21437 ( .A1(n18603), .A2(n18416), .B1(n18685), .B2(n18415), .ZN(
        n18411) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18417), .B1(
        n18688), .B2(n18484), .ZN(n18410) );
  OAI211_X1 U21439 ( .C1(n18606), .C2(n18441), .A(n18411), .B(n18410), .ZN(
        P3_U2913) );
  AOI22_X1 U21440 ( .A1(n18638), .A2(n18428), .B1(n18693), .B2(n18415), .ZN(
        n18413) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18417), .B1(
        n18695), .B2(n18484), .ZN(n18412) );
  OAI211_X1 U21442 ( .C1(n18641), .C2(n18414), .A(n18413), .B(n18412), .ZN(
        P3_U2914) );
  AOI22_X1 U21443 ( .A1(n18702), .A2(n18416), .B1(n18700), .B2(n18415), .ZN(
        n18419) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18417), .B1(
        n18703), .B2(n18484), .ZN(n18418) );
  OAI211_X1 U21445 ( .C1(n18708), .C2(n18441), .A(n18419), .B(n18418), .ZN(
        P3_U2915) );
  NAND2_X1 U21446 ( .A1(n18514), .A2(n18443), .ZN(n18513) );
  INV_X1 U21447 ( .A(n18513), .ZN(n18506) );
  NOR2_X1 U21448 ( .A1(n18484), .A2(n18506), .ZN(n18464) );
  OAI21_X1 U21449 ( .B1(n18420), .B2(n18618), .A(n18464), .ZN(n18421) );
  OAI211_X1 U21450 ( .C1(n18506), .C2(n18878), .A(n18621), .B(n18421), .ZN(
        n18438) );
  NOR2_X1 U21451 ( .A1(n18616), .A2(n18464), .ZN(n18437) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18438), .B1(
        n18650), .B2(n18437), .ZN(n18423) );
  AOI22_X1 U21453 ( .A1(n18651), .A2(n18456), .B1(n18656), .B2(n18428), .ZN(
        n18422) );
  OAI211_X1 U21454 ( .C1(n18659), .C2(n18513), .A(n18423), .B(n18422), .ZN(
        P3_U2916) );
  AOI22_X1 U21455 ( .A1(n18591), .A2(n18428), .B1(n18661), .B2(n18437), .ZN(
        n18425) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18438), .B1(
        n18662), .B2(n18456), .ZN(n18424) );
  OAI211_X1 U21457 ( .C1(n18594), .C2(n18513), .A(n18425), .B(n18424), .ZN(
        P3_U2917) );
  AOI22_X1 U21458 ( .A1(n18628), .A2(n18428), .B1(n18667), .B2(n18437), .ZN(
        n18427) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18438), .B1(
        n18668), .B2(n18456), .ZN(n18426) );
  OAI211_X1 U21460 ( .C1(n18548), .C2(n18513), .A(n18427), .B(n18426), .ZN(
        P3_U2918) );
  AOI22_X1 U21461 ( .A1(n18597), .A2(n18428), .B1(n18673), .B2(n18437), .ZN(
        n18430) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18438), .B1(
        n18674), .B2(n18456), .ZN(n18429) );
  OAI211_X1 U21463 ( .C1(n18551), .C2(n18513), .A(n18430), .B(n18429), .ZN(
        P3_U2919) );
  AOI22_X1 U21464 ( .A1(n18680), .A2(n18456), .B1(n18679), .B2(n18437), .ZN(
        n18432) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18438), .B1(
        n18681), .B2(n18506), .ZN(n18431) );
  OAI211_X1 U21466 ( .C1(n18684), .C2(n18441), .A(n18432), .B(n18431), .ZN(
        P3_U2920) );
  AOI22_X1 U21467 ( .A1(n18686), .A2(n18456), .B1(n18685), .B2(n18437), .ZN(
        n18434) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18438), .B1(
        n18688), .B2(n18506), .ZN(n18433) );
  OAI211_X1 U21469 ( .C1(n18692), .C2(n18441), .A(n18434), .B(n18433), .ZN(
        P3_U2921) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18438), .B1(
        n18693), .B2(n18437), .ZN(n18436) );
  AOI22_X1 U21471 ( .A1(n18695), .A2(n18506), .B1(n18638), .B2(n18456), .ZN(
        n18435) );
  OAI211_X1 U21472 ( .C1(n18641), .C2(n18441), .A(n18436), .B(n18435), .ZN(
        P3_U2922) );
  AOI22_X1 U21473 ( .A1(n18643), .A2(n18456), .B1(n18700), .B2(n18437), .ZN(
        n18440) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18438), .B1(
        n18703), .B2(n18506), .ZN(n18439) );
  OAI211_X1 U21475 ( .C1(n18649), .C2(n18441), .A(n18440), .B(n18439), .ZN(
        P3_U2923) );
  AOI22_X1 U21476 ( .A1(n18656), .A2(n18456), .B1(n18650), .B2(n18459), .ZN(
        n18445) );
  NAND2_X1 U21477 ( .A1(n18442), .A2(n18443), .ZN(n18460) );
  NAND2_X1 U21478 ( .A1(n18750), .A2(n18443), .ZN(n18536) );
  INV_X1 U21479 ( .A(n18536), .ZN(n18517) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18460), .B1(
        n18466), .B2(n18517), .ZN(n18444) );
  OAI211_X1 U21481 ( .C1(n18469), .C2(n18482), .A(n18445), .B(n18444), .ZN(
        P3_U2924) );
  AOI22_X1 U21482 ( .A1(n18591), .A2(n18456), .B1(n18661), .B2(n18459), .ZN(
        n18447) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18460), .B1(
        n18662), .B2(n18484), .ZN(n18446) );
  OAI211_X1 U21484 ( .C1(n18594), .C2(n18536), .A(n18447), .B(n18446), .ZN(
        P3_U2925) );
  AOI22_X1 U21485 ( .A1(n18628), .A2(n18456), .B1(n18667), .B2(n18459), .ZN(
        n18449) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18460), .B1(
        n18669), .B2(n18517), .ZN(n18448) );
  OAI211_X1 U21487 ( .C1(n18631), .C2(n18482), .A(n18449), .B(n18448), .ZN(
        P3_U2926) );
  AOI22_X1 U21488 ( .A1(n18674), .A2(n18484), .B1(n18673), .B2(n18459), .ZN(
        n18451) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18460), .B1(
        n18597), .B2(n18456), .ZN(n18450) );
  OAI211_X1 U21490 ( .C1(n18551), .C2(n18536), .A(n18451), .B(n18450), .ZN(
        P3_U2927) );
  AOI22_X1 U21491 ( .A1(n18680), .A2(n18484), .B1(n18679), .B2(n18459), .ZN(
        n18453) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18460), .B1(
        n18681), .B2(n18517), .ZN(n18452) );
  OAI211_X1 U21493 ( .C1(n18684), .C2(n18463), .A(n18453), .B(n18452), .ZN(
        P3_U2928) );
  AOI22_X1 U21494 ( .A1(n18686), .A2(n18484), .B1(n18685), .B2(n18459), .ZN(
        n18455) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18460), .B1(
        n18688), .B2(n18517), .ZN(n18454) );
  OAI211_X1 U21496 ( .C1(n18692), .C2(n18463), .A(n18455), .B(n18454), .ZN(
        P3_U2929) );
  AOI22_X1 U21497 ( .A1(n18694), .A2(n18456), .B1(n18693), .B2(n18459), .ZN(
        n18458) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18460), .B1(
        n18695), .B2(n18517), .ZN(n18457) );
  OAI211_X1 U21499 ( .C1(n18698), .C2(n18482), .A(n18458), .B(n18457), .ZN(
        P3_U2930) );
  AOI22_X1 U21500 ( .A1(n18643), .A2(n18484), .B1(n18700), .B2(n18459), .ZN(
        n18462) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18460), .B1(
        n18703), .B2(n18517), .ZN(n18461) );
  OAI211_X1 U21502 ( .C1(n18649), .C2(n18463), .A(n18462), .B(n18461), .ZN(
        P3_U2931) );
  NOR2_X1 U21503 ( .A1(n18517), .A2(n18541), .ZN(n18515) );
  OAI21_X1 U21504 ( .B1(n18464), .B2(n18618), .A(n18515), .ZN(n18465) );
  OAI211_X1 U21505 ( .C1(n18541), .C2(n18878), .A(n18621), .B(n18465), .ZN(
        n18485) );
  NOR2_X1 U21506 ( .A1(n18616), .A2(n18515), .ZN(n18483) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18485), .B1(
        n18650), .B2(n18483), .ZN(n18468) );
  AOI22_X1 U21508 ( .A1(n18466), .A2(n18541), .B1(n18656), .B2(n18484), .ZN(
        n18467) );
  OAI211_X1 U21509 ( .C1(n18469), .C2(n18513), .A(n18468), .B(n18467), .ZN(
        P3_U2932) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18485), .B1(
        n18661), .B2(n18483), .ZN(n18471) );
  AOI22_X1 U21511 ( .A1(n18663), .A2(n18541), .B1(n18662), .B2(n18506), .ZN(
        n18470) );
  OAI211_X1 U21512 ( .C1(n18666), .C2(n18482), .A(n18471), .B(n18470), .ZN(
        P3_U2933) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18485), .B1(
        n18667), .B2(n18483), .ZN(n18473) );
  AOI22_X1 U21514 ( .A1(n18669), .A2(n18541), .B1(n18628), .B2(n18484), .ZN(
        n18472) );
  OAI211_X1 U21515 ( .C1(n18631), .C2(n18513), .A(n18473), .B(n18472), .ZN(
        P3_U2934) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18485), .B1(
        n18673), .B2(n18483), .ZN(n18475) );
  AOI22_X1 U21517 ( .A1(n18674), .A2(n18506), .B1(n18675), .B2(n18541), .ZN(
        n18474) );
  OAI211_X1 U21518 ( .C1(n18678), .C2(n18482), .A(n18475), .B(n18474), .ZN(
        P3_U2935) );
  AOI22_X1 U21519 ( .A1(n18573), .A2(n18484), .B1(n18679), .B2(n18483), .ZN(
        n18477) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18485), .B1(
        n18681), .B2(n18541), .ZN(n18476) );
  OAI211_X1 U21521 ( .C1(n18576), .C2(n18513), .A(n18477), .B(n18476), .ZN(
        P3_U2936) );
  AOI22_X1 U21522 ( .A1(n18686), .A2(n18506), .B1(n18685), .B2(n18483), .ZN(
        n18479) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18485), .B1(
        n18688), .B2(n18541), .ZN(n18478) );
  OAI211_X1 U21524 ( .C1(n18692), .C2(n18482), .A(n18479), .B(n18478), .ZN(
        P3_U2937) );
  AOI22_X1 U21525 ( .A1(n18638), .A2(n18506), .B1(n18693), .B2(n18483), .ZN(
        n18481) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18485), .B1(
        n18695), .B2(n18541), .ZN(n18480) );
  OAI211_X1 U21527 ( .C1(n18641), .C2(n18482), .A(n18481), .B(n18480), .ZN(
        P3_U2938) );
  AOI22_X1 U21528 ( .A1(n18702), .A2(n18484), .B1(n18700), .B2(n18483), .ZN(
        n18487) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18485), .B1(
        n18703), .B2(n18541), .ZN(n18486) );
  OAI211_X1 U21530 ( .C1(n18708), .C2(n18513), .A(n18487), .B(n18486), .ZN(
        P3_U2939) );
  NAND2_X1 U21531 ( .A1(n18488), .A2(n18540), .ZN(n18581) );
  INV_X1 U21532 ( .A(n18540), .ZN(n18538) );
  NOR2_X1 U21533 ( .A1(n18489), .A2(n18538), .ZN(n18509) );
  AOI22_X1 U21534 ( .A1(n18656), .A2(n18506), .B1(n18650), .B2(n18509), .ZN(
        n18495) );
  NOR2_X1 U21535 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18490), .ZN(
        n18493) );
  INV_X1 U21536 ( .A(n18491), .ZN(n18653) );
  NOR2_X1 U21537 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18538), .ZN(
        n18492) );
  AOI22_X1 U21538 ( .A1(n18655), .A2(n18493), .B1(n18653), .B2(n18492), .ZN(
        n18510) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18510), .B1(
        n18651), .B2(n18517), .ZN(n18494) );
  OAI211_X1 U21540 ( .C1(n18659), .C2(n18581), .A(n18495), .B(n18494), .ZN(
        P3_U2940) );
  AOI22_X1 U21541 ( .A1(n18591), .A2(n18506), .B1(n18661), .B2(n18509), .ZN(
        n18497) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18510), .B1(
        n18662), .B2(n18517), .ZN(n18496) );
  OAI211_X1 U21543 ( .C1(n18594), .C2(n18581), .A(n18497), .B(n18496), .ZN(
        P3_U2941) );
  AOI22_X1 U21544 ( .A1(n18668), .A2(n18517), .B1(n18667), .B2(n18509), .ZN(
        n18499) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18510), .B1(
        n18628), .B2(n18506), .ZN(n18498) );
  OAI211_X1 U21546 ( .C1(n18548), .C2(n18581), .A(n18499), .B(n18498), .ZN(
        P3_U2942) );
  AOI22_X1 U21547 ( .A1(n18674), .A2(n18517), .B1(n18673), .B2(n18509), .ZN(
        n18501) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18510), .B1(
        n18597), .B2(n18506), .ZN(n18500) );
  OAI211_X1 U21549 ( .C1(n18551), .C2(n18581), .A(n18501), .B(n18500), .ZN(
        P3_U2943) );
  AOI22_X1 U21550 ( .A1(n18680), .A2(n18517), .B1(n18679), .B2(n18509), .ZN(
        n18503) );
  INV_X1 U21551 ( .A(n18581), .ZN(n18583) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18510), .B1(
        n18681), .B2(n18583), .ZN(n18502) );
  OAI211_X1 U21553 ( .C1(n18684), .C2(n18513), .A(n18503), .B(n18502), .ZN(
        P3_U2944) );
  AOI22_X1 U21554 ( .A1(n18603), .A2(n18506), .B1(n18685), .B2(n18509), .ZN(
        n18505) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18510), .B1(
        n18688), .B2(n18583), .ZN(n18504) );
  OAI211_X1 U21556 ( .C1(n18606), .C2(n18536), .A(n18505), .B(n18504), .ZN(
        P3_U2945) );
  AOI22_X1 U21557 ( .A1(n18694), .A2(n18506), .B1(n18693), .B2(n18509), .ZN(
        n18508) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18510), .B1(
        n18695), .B2(n18583), .ZN(n18507) );
  OAI211_X1 U21559 ( .C1(n18698), .C2(n18536), .A(n18508), .B(n18507), .ZN(
        P3_U2946) );
  AOI22_X1 U21560 ( .A1(n18643), .A2(n18517), .B1(n18700), .B2(n18509), .ZN(
        n18512) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18510), .B1(
        n18703), .B2(n18583), .ZN(n18511) );
  OAI211_X1 U21562 ( .C1(n18649), .C2(n18513), .A(n18512), .B(n18511), .ZN(
        P3_U2947) );
  NAND2_X1 U21563 ( .A1(n18514), .A2(n18540), .ZN(n18609) );
  AOI21_X1 U21564 ( .B1(n18581), .B2(n18609), .A(n18616), .ZN(n18532) );
  AOI22_X1 U21565 ( .A1(n18651), .A2(n18541), .B1(n18650), .B2(n18532), .ZN(
        n18519) );
  INV_X1 U21566 ( .A(n18609), .ZN(n18611) );
  OAI211_X1 U21567 ( .C1(n18515), .C2(n18618), .A(n18581), .B(n18609), .ZN(
        n18516) );
  OAI211_X1 U21568 ( .C1(n18611), .C2(n18878), .A(n18621), .B(n18516), .ZN(
        n18533) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18533), .B1(
        n18656), .B2(n18517), .ZN(n18518) );
  OAI211_X1 U21570 ( .C1(n18659), .C2(n18609), .A(n18519), .B(n18518), .ZN(
        P3_U2948) );
  AOI22_X1 U21571 ( .A1(n18662), .A2(n18541), .B1(n18661), .B2(n18532), .ZN(
        n18521) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18533), .B1(
        n18663), .B2(n18611), .ZN(n18520) );
  OAI211_X1 U21573 ( .C1(n18666), .C2(n18536), .A(n18521), .B(n18520), .ZN(
        P3_U2949) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18533), .B1(
        n18667), .B2(n18532), .ZN(n18523) );
  AOI22_X1 U21575 ( .A1(n18668), .A2(n18541), .B1(n18669), .B2(n18611), .ZN(
        n18522) );
  OAI211_X1 U21576 ( .C1(n18672), .C2(n18536), .A(n18523), .B(n18522), .ZN(
        P3_U2950) );
  AOI22_X1 U21577 ( .A1(n18674), .A2(n18541), .B1(n18673), .B2(n18532), .ZN(
        n18525) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18533), .B1(
        n18675), .B2(n18611), .ZN(n18524) );
  OAI211_X1 U21579 ( .C1(n18678), .C2(n18536), .A(n18525), .B(n18524), .ZN(
        P3_U2951) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18533), .B1(
        n18679), .B2(n18532), .ZN(n18527) );
  AOI22_X1 U21581 ( .A1(n18681), .A2(n18611), .B1(n18680), .B2(n18541), .ZN(
        n18526) );
  OAI211_X1 U21582 ( .C1(n18684), .C2(n18536), .A(n18527), .B(n18526), .ZN(
        P3_U2952) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18533), .B1(
        n18685), .B2(n18532), .ZN(n18529) );
  AOI22_X1 U21584 ( .A1(n18686), .A2(n18541), .B1(n18688), .B2(n18611), .ZN(
        n18528) );
  OAI211_X1 U21585 ( .C1(n18692), .C2(n18536), .A(n18529), .B(n18528), .ZN(
        P3_U2953) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18533), .B1(
        n18693), .B2(n18532), .ZN(n18531) );
  AOI22_X1 U21587 ( .A1(n18695), .A2(n18611), .B1(n18638), .B2(n18541), .ZN(
        n18530) );
  OAI211_X1 U21588 ( .C1(n18641), .C2(n18536), .A(n18531), .B(n18530), .ZN(
        P3_U2954) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18533), .B1(
        n18700), .B2(n18532), .ZN(n18535) );
  AOI22_X1 U21590 ( .A1(n18703), .A2(n18611), .B1(n18643), .B2(n18541), .ZN(
        n18534) );
  OAI211_X1 U21591 ( .C1(n18649), .C2(n18536), .A(n18535), .B(n18534), .ZN(
        P3_U2955) );
  NOR2_X2 U21592 ( .A1(n18537), .A2(n18538), .ZN(n18627) );
  INV_X1 U21593 ( .A(n18627), .ZN(n18648) );
  NOR2_X1 U21594 ( .A1(n18539), .A2(n18538), .ZN(n18588) );
  AND2_X1 U21595 ( .A1(n18776), .A2(n18588), .ZN(n18558) );
  AOI22_X1 U21596 ( .A1(n18651), .A2(n18583), .B1(n18650), .B2(n18558), .ZN(
        n18543) );
  OAI211_X1 U21597 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18655), .A(
        n18653), .B(n18540), .ZN(n18559) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18559), .B1(
        n18656), .B2(n18541), .ZN(n18542) );
  OAI211_X1 U21599 ( .C1(n18659), .C2(n18648), .A(n18543), .B(n18542), .ZN(
        P3_U2956) );
  AOI22_X1 U21600 ( .A1(n18591), .A2(n18541), .B1(n18661), .B2(n18558), .ZN(
        n18545) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18559), .B1(
        n18662), .B2(n18583), .ZN(n18544) );
  OAI211_X1 U21602 ( .C1(n18594), .C2(n18648), .A(n18545), .B(n18544), .ZN(
        P3_U2957) );
  AOI22_X1 U21603 ( .A1(n18628), .A2(n18541), .B1(n18667), .B2(n18558), .ZN(
        n18547) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18559), .B1(
        n18668), .B2(n18583), .ZN(n18546) );
  OAI211_X1 U21605 ( .C1(n18548), .C2(n18648), .A(n18547), .B(n18546), .ZN(
        P3_U2958) );
  AOI22_X1 U21606 ( .A1(n18597), .A2(n18541), .B1(n18673), .B2(n18558), .ZN(
        n18550) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18559), .B1(
        n18674), .B2(n18583), .ZN(n18549) );
  OAI211_X1 U21608 ( .C1(n18551), .C2(n18648), .A(n18550), .B(n18549), .ZN(
        P3_U2959) );
  AOI22_X1 U21609 ( .A1(n18573), .A2(n18541), .B1(n18679), .B2(n18558), .ZN(
        n18553) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18559), .B1(
        n18681), .B2(n18627), .ZN(n18552) );
  OAI211_X1 U21611 ( .C1(n18576), .C2(n18581), .A(n18553), .B(n18552), .ZN(
        P3_U2960) );
  AOI22_X1 U21612 ( .A1(n18603), .A2(n18541), .B1(n18685), .B2(n18558), .ZN(
        n18555) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18559), .B1(
        n18688), .B2(n18627), .ZN(n18554) );
  OAI211_X1 U21614 ( .C1(n18606), .C2(n18581), .A(n18555), .B(n18554), .ZN(
        P3_U2961) );
  AOI22_X1 U21615 ( .A1(n18694), .A2(n18541), .B1(n18693), .B2(n18558), .ZN(
        n18557) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18559), .B1(
        n18695), .B2(n18627), .ZN(n18556) );
  OAI211_X1 U21617 ( .C1(n18698), .C2(n18581), .A(n18557), .B(n18556), .ZN(
        P3_U2962) );
  AOI22_X1 U21618 ( .A1(n18702), .A2(n18541), .B1(n18700), .B2(n18558), .ZN(
        n18561) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18559), .B1(
        n18703), .B2(n18627), .ZN(n18560) );
  OAI211_X1 U21620 ( .C1(n18708), .C2(n18581), .A(n18561), .B(n18560), .ZN(
        P3_U2963) );
  INV_X1 U21621 ( .A(n18654), .ZN(n18587) );
  NOR2_X2 U21622 ( .A1(n18587), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18701) );
  INV_X1 U21623 ( .A(n18701), .ZN(n18691) );
  AOI21_X1 U21624 ( .B1(n18648), .B2(n18691), .A(n18616), .ZN(n18582) );
  AOI22_X1 U21625 ( .A1(n18651), .A2(n18611), .B1(n18650), .B2(n18582), .ZN(
        n18566) );
  AOI221_X1 U21626 ( .B1(n18563), .B2(n18648), .C1(n18562), .C2(n18648), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18564) );
  OAI21_X1 U21627 ( .B1(n18701), .B2(n18564), .A(n18621), .ZN(n18584) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18584), .B1(
        n18656), .B2(n18583), .ZN(n18565) );
  OAI211_X1 U21629 ( .C1(n18659), .C2(n18691), .A(n18566), .B(n18565), .ZN(
        P3_U2964) );
  AOI22_X1 U21630 ( .A1(n18662), .A2(n18611), .B1(n18661), .B2(n18582), .ZN(
        n18568) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18584), .B1(
        n18663), .B2(n18701), .ZN(n18567) );
  OAI211_X1 U21632 ( .C1(n18666), .C2(n18581), .A(n18568), .B(n18567), .ZN(
        P3_U2965) );
  AOI22_X1 U21633 ( .A1(n18628), .A2(n18583), .B1(n18667), .B2(n18582), .ZN(
        n18570) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18584), .B1(
        n18669), .B2(n18701), .ZN(n18569) );
  OAI211_X1 U21635 ( .C1(n18631), .C2(n18609), .A(n18570), .B(n18569), .ZN(
        P3_U2966) );
  AOI22_X1 U21636 ( .A1(n18674), .A2(n18611), .B1(n18673), .B2(n18582), .ZN(
        n18572) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18584), .B1(
        n18675), .B2(n18701), .ZN(n18571) );
  OAI211_X1 U21638 ( .C1(n18678), .C2(n18581), .A(n18572), .B(n18571), .ZN(
        P3_U2967) );
  AOI22_X1 U21639 ( .A1(n18573), .A2(n18583), .B1(n18679), .B2(n18582), .ZN(
        n18575) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18584), .B1(
        n18681), .B2(n18701), .ZN(n18574) );
  OAI211_X1 U21641 ( .C1(n18576), .C2(n18609), .A(n18575), .B(n18574), .ZN(
        P3_U2968) );
  AOI22_X1 U21642 ( .A1(n18686), .A2(n18611), .B1(n18685), .B2(n18582), .ZN(
        n18578) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18584), .B1(
        n18688), .B2(n18701), .ZN(n18577) );
  OAI211_X1 U21644 ( .C1(n18692), .C2(n18581), .A(n18578), .B(n18577), .ZN(
        P3_U2969) );
  AOI22_X1 U21645 ( .A1(n18638), .A2(n18611), .B1(n18693), .B2(n18582), .ZN(
        n18580) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18584), .B1(
        n18695), .B2(n18701), .ZN(n18579) );
  OAI211_X1 U21647 ( .C1(n18641), .C2(n18581), .A(n18580), .B(n18579), .ZN(
        P3_U2970) );
  AOI22_X1 U21648 ( .A1(n18702), .A2(n18583), .B1(n18700), .B2(n18582), .ZN(
        n18586) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18584), .B1(
        n18703), .B2(n18701), .ZN(n18585) );
  OAI211_X1 U21650 ( .C1(n18708), .C2(n18609), .A(n18586), .B(n18585), .ZN(
        P3_U2971) );
  NOR2_X1 U21651 ( .A1(n18616), .A2(n18587), .ZN(n18610) );
  AOI22_X1 U21652 ( .A1(n18651), .A2(n18627), .B1(n18650), .B2(n18610), .ZN(
        n18590) );
  AOI22_X1 U21653 ( .A1(n18655), .A2(n18588), .B1(n18654), .B2(n18653), .ZN(
        n18612) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18612), .B1(
        n18656), .B2(n18611), .ZN(n18589) );
  OAI211_X1 U21655 ( .C1(n18659), .C2(n18709), .A(n18590), .B(n18589), .ZN(
        P3_U2972) );
  AOI22_X1 U21656 ( .A1(n18591), .A2(n18611), .B1(n18661), .B2(n18610), .ZN(
        n18593) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18612), .B1(
        n18662), .B2(n18627), .ZN(n18592) );
  OAI211_X1 U21658 ( .C1(n18709), .C2(n18594), .A(n18593), .B(n18592), .ZN(
        P3_U2973) );
  AOI22_X1 U21659 ( .A1(n18668), .A2(n18627), .B1(n18667), .B2(n18610), .ZN(
        n18596) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18612), .B1(
        n18687), .B2(n18669), .ZN(n18595) );
  OAI211_X1 U21661 ( .C1(n18672), .C2(n18609), .A(n18596), .B(n18595), .ZN(
        P3_U2974) );
  AOI22_X1 U21662 ( .A1(n18597), .A2(n18611), .B1(n18673), .B2(n18610), .ZN(
        n18599) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18612), .B1(
        n18687), .B2(n18675), .ZN(n18598) );
  OAI211_X1 U21664 ( .C1(n18600), .C2(n18648), .A(n18599), .B(n18598), .ZN(
        P3_U2975) );
  AOI22_X1 U21665 ( .A1(n18680), .A2(n18627), .B1(n18679), .B2(n18610), .ZN(
        n18602) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18612), .B1(
        n18687), .B2(n18681), .ZN(n18601) );
  OAI211_X1 U21667 ( .C1(n18684), .C2(n18609), .A(n18602), .B(n18601), .ZN(
        P3_U2976) );
  AOI22_X1 U21668 ( .A1(n18603), .A2(n18611), .B1(n18685), .B2(n18610), .ZN(
        n18605) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18612), .B1(
        n18687), .B2(n18688), .ZN(n18604) );
  OAI211_X1 U21670 ( .C1(n18606), .C2(n18648), .A(n18605), .B(n18604), .ZN(
        P3_U2977) );
  AOI22_X1 U21671 ( .A1(n18638), .A2(n18627), .B1(n18693), .B2(n18610), .ZN(
        n18608) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18612), .B1(
        n18687), .B2(n18695), .ZN(n18607) );
  OAI211_X1 U21673 ( .C1(n18641), .C2(n18609), .A(n18608), .B(n18607), .ZN(
        P3_U2978) );
  AOI22_X1 U21674 ( .A1(n18702), .A2(n18611), .B1(n18700), .B2(n18610), .ZN(
        n18614) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18612), .B1(
        n18687), .B2(n18703), .ZN(n18613) );
  OAI211_X1 U21676 ( .C1(n18708), .C2(n18648), .A(n18614), .B(n18613), .ZN(
        P3_U2979) );
  INV_X1 U21677 ( .A(n18615), .ZN(n18617) );
  NOR2_X1 U21678 ( .A1(n18616), .A2(n18617), .ZN(n18642) );
  AOI22_X1 U21679 ( .A1(n18651), .A2(n18701), .B1(n18650), .B2(n18642), .ZN(
        n18623) );
  NOR2_X1 U21680 ( .A1(n18627), .A2(n18701), .ZN(n18619) );
  OAI21_X1 U21681 ( .B1(n18619), .B2(n18618), .A(n18617), .ZN(n18620) );
  OAI211_X1 U21682 ( .C1(n18644), .C2(n18878), .A(n18621), .B(n18620), .ZN(
        n18645) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18645), .B1(
        n18656), .B2(n18627), .ZN(n18622) );
  OAI211_X1 U21684 ( .C1(n18624), .C2(n18659), .A(n18623), .B(n18622), .ZN(
        P3_U2980) );
  AOI22_X1 U21685 ( .A1(n18662), .A2(n18701), .B1(n18661), .B2(n18642), .ZN(
        n18626) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18645), .B1(
        n18644), .B2(n18663), .ZN(n18625) );
  OAI211_X1 U21687 ( .C1(n18666), .C2(n18648), .A(n18626), .B(n18625), .ZN(
        P3_U2981) );
  AOI22_X1 U21688 ( .A1(n18628), .A2(n18627), .B1(n18667), .B2(n18642), .ZN(
        n18630) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18645), .B1(
        n18644), .B2(n18669), .ZN(n18629) );
  OAI211_X1 U21690 ( .C1(n18631), .C2(n18691), .A(n18630), .B(n18629), .ZN(
        P3_U2982) );
  AOI22_X1 U21691 ( .A1(n18674), .A2(n18701), .B1(n18673), .B2(n18642), .ZN(
        n18633) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18645), .B1(
        n18644), .B2(n18675), .ZN(n18632) );
  OAI211_X1 U21693 ( .C1(n18678), .C2(n18648), .A(n18633), .B(n18632), .ZN(
        P3_U2983) );
  AOI22_X1 U21694 ( .A1(n18680), .A2(n18701), .B1(n18679), .B2(n18642), .ZN(
        n18635) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18645), .B1(
        n18644), .B2(n18681), .ZN(n18634) );
  OAI211_X1 U21696 ( .C1(n18684), .C2(n18648), .A(n18635), .B(n18634), .ZN(
        P3_U2984) );
  AOI22_X1 U21697 ( .A1(n18686), .A2(n18701), .B1(n18685), .B2(n18642), .ZN(
        n18637) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18645), .B1(
        n18644), .B2(n18688), .ZN(n18636) );
  OAI211_X1 U21699 ( .C1(n18692), .C2(n18648), .A(n18637), .B(n18636), .ZN(
        P3_U2985) );
  AOI22_X1 U21700 ( .A1(n18638), .A2(n18701), .B1(n18693), .B2(n18642), .ZN(
        n18640) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18645), .B1(
        n18644), .B2(n18695), .ZN(n18639) );
  OAI211_X1 U21702 ( .C1(n18641), .C2(n18648), .A(n18640), .B(n18639), .ZN(
        P3_U2986) );
  AOI22_X1 U21703 ( .A1(n18643), .A2(n18701), .B1(n18700), .B2(n18642), .ZN(
        n18647) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18645), .B1(
        n18644), .B2(n18703), .ZN(n18646) );
  OAI211_X1 U21705 ( .C1(n18649), .C2(n18648), .A(n18647), .B(n18646), .ZN(
        P3_U2987) );
  AND2_X1 U21706 ( .A1(n18776), .A2(n18652), .ZN(n18699) );
  AOI22_X1 U21707 ( .A1(n18651), .A2(n18687), .B1(n18650), .B2(n18699), .ZN(
        n18658) );
  AOI22_X1 U21708 ( .A1(n18655), .A2(n18654), .B1(n18653), .B2(n18652), .ZN(
        n18705) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18705), .B1(
        n18656), .B2(n18701), .ZN(n18657) );
  OAI211_X1 U21710 ( .C1(n18660), .C2(n18659), .A(n18658), .B(n18657), .ZN(
        P3_U2988) );
  AOI22_X1 U21711 ( .A1(n18687), .A2(n18662), .B1(n18661), .B2(n18699), .ZN(
        n18665) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18705), .B1(
        n18704), .B2(n18663), .ZN(n18664) );
  OAI211_X1 U21713 ( .C1(n18666), .C2(n18691), .A(n18665), .B(n18664), .ZN(
        P3_U2989) );
  AOI22_X1 U21714 ( .A1(n18687), .A2(n18668), .B1(n18667), .B2(n18699), .ZN(
        n18671) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18705), .B1(
        n18704), .B2(n18669), .ZN(n18670) );
  OAI211_X1 U21716 ( .C1(n18672), .C2(n18691), .A(n18671), .B(n18670), .ZN(
        P3_U2990) );
  AOI22_X1 U21717 ( .A1(n18687), .A2(n18674), .B1(n18673), .B2(n18699), .ZN(
        n18677) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18705), .B1(
        n18704), .B2(n18675), .ZN(n18676) );
  OAI211_X1 U21719 ( .C1(n18678), .C2(n18691), .A(n18677), .B(n18676), .ZN(
        P3_U2991) );
  AOI22_X1 U21720 ( .A1(n18687), .A2(n18680), .B1(n18679), .B2(n18699), .ZN(
        n18683) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18705), .B1(
        n18704), .B2(n18681), .ZN(n18682) );
  OAI211_X1 U21722 ( .C1(n18684), .C2(n18691), .A(n18683), .B(n18682), .ZN(
        P3_U2992) );
  AOI22_X1 U21723 ( .A1(n18687), .A2(n18686), .B1(n18685), .B2(n18699), .ZN(
        n18690) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18705), .B1(
        n18704), .B2(n18688), .ZN(n18689) );
  OAI211_X1 U21725 ( .C1(n18692), .C2(n18691), .A(n18690), .B(n18689), .ZN(
        P3_U2993) );
  AOI22_X1 U21726 ( .A1(n18694), .A2(n18701), .B1(n18693), .B2(n18699), .ZN(
        n18697) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18705), .B1(
        n18704), .B2(n18695), .ZN(n18696) );
  OAI211_X1 U21728 ( .C1(n18709), .C2(n18698), .A(n18697), .B(n18696), .ZN(
        P3_U2994) );
  AOI22_X1 U21729 ( .A1(n18702), .A2(n18701), .B1(n18700), .B2(n18699), .ZN(
        n18707) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18705), .B1(
        n18704), .B2(n18703), .ZN(n18706) );
  OAI211_X1 U21731 ( .C1(n18709), .C2(n18708), .A(n18707), .B(n18706), .ZN(
        P3_U2995) );
  NOR2_X1 U21732 ( .A1(n10213), .A2(n18710), .ZN(n18711) );
  OAI22_X1 U21733 ( .A1(n18714), .A2(n18713), .B1(n18712), .B2(n18711), .ZN(
        n18715) );
  AOI221_X1 U21734 ( .B1(n18718), .B2(n18717), .C1(n18716), .C2(n18717), .A(
        n18715), .ZN(n18922) );
  OAI211_X1 U21735 ( .C1(n18721), .C2(n18752), .A(n18720), .B(n18719), .ZN(
        n18722) );
  AOI221_X1 U21736 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n18723), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n18723), .A(n18722), .ZN(n18764) );
  INV_X1 U21737 ( .A(n18752), .ZN(n18743) );
  AOI21_X1 U21738 ( .B1(n18726), .B2(n18725), .A(n18724), .ZN(n18737) );
  AOI22_X1 U21739 ( .A1(n18891), .A2(n18739), .B1(n18731), .B2(n18749), .ZN(
        n18727) );
  OAI21_X1 U21740 ( .B1(n18737), .B2(n18728), .A(n18727), .ZN(n18882) );
  NOR2_X1 U21741 ( .A1(n18743), .A2(n18882), .ZN(n18734) );
  AND2_X1 U21742 ( .A1(n18891), .A2(n18739), .ZN(n18732) );
  OAI21_X1 U21743 ( .B1(n18745), .B2(n18909), .A(n18729), .ZN(n18736) );
  NOR2_X1 U21744 ( .A1(n18730), .A2(n18736), .ZN(n18746) );
  OAI22_X1 U21745 ( .A1(n18732), .A2(n18742), .B1(n18746), .B2(n18731), .ZN(
        n18879) );
  NAND2_X1 U21746 ( .A1(n18883), .A2(n18879), .ZN(n18733) );
  OAI22_X1 U21747 ( .A1(n18734), .A2(n18883), .B1(n18743), .B2(n18733), .ZN(
        n18759) );
  NAND2_X1 U21748 ( .A1(n18901), .A2(n18891), .ZN(n18735) );
  OAI221_X1 U21749 ( .B1(n18901), .B2(n18891), .C1(n10213), .C2(n18736), .A(
        n18735), .ZN(n18741) );
  INV_X1 U21750 ( .A(n18737), .ZN(n18738) );
  NAND3_X1 U21751 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18739), .A3(
        n18738), .ZN(n18740) );
  OAI211_X1 U21752 ( .C1(n18888), .C2(n18742), .A(n18741), .B(n18740), .ZN(
        n18889) );
  AOI22_X1 U21753 ( .A1(n18743), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18889), .B2(n18752), .ZN(n18758) );
  NAND2_X1 U21754 ( .A1(n18745), .A2(n18744), .ZN(n18748) );
  INV_X1 U21755 ( .A(n18746), .ZN(n18747) );
  AOI22_X1 U21756 ( .A1(n18896), .A2(n18748), .B1(n18901), .B2(n18747), .ZN(
        n18892) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18749), .B1(
        n18748), .B2(n18909), .ZN(n18903) );
  AOI222_X1 U21758 ( .A1(n18892), .A2(n18903), .B1(n18892), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n18903), .C2(n18750), .ZN(
        n18753) );
  AOI21_X1 U21759 ( .B1(n18753), .B2(n18752), .A(n18751), .ZN(n18754) );
  AOI222_X1 U21760 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18758), 
        .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18754), .C1(n18758), 
        .C2(n18754), .ZN(n18756) );
  OAI211_X1 U21761 ( .C1(n18759), .C2(n18757), .A(n18756), .B(n18755), .ZN(
        n18763) );
  NOR2_X1 U21762 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18761) );
  INV_X1 U21763 ( .A(n18758), .ZN(n18760) );
  OAI21_X1 U21764 ( .B1(n18761), .B2(n18760), .A(n18759), .ZN(n18762) );
  NAND4_X1 U21765 ( .A1(n18922), .A2(n18764), .A3(n18763), .A4(n18762), .ZN(
        n18770) );
  AOI211_X1 U21766 ( .C1(n18766), .C2(n18765), .A(n18925), .B(n18770), .ZN(
        n18875) );
  NOR2_X1 U21767 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18794), .ZN(n18774) );
  NOR2_X1 U21768 ( .A1(n18875), .A2(n18774), .ZN(n18777) );
  NOR2_X1 U21769 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18935) );
  NAND2_X1 U21770 ( .A1(n9890), .A2(n17507), .ZN(n18780) );
  INV_X1 U21771 ( .A(n18780), .ZN(n18767) );
  AOI211_X1 U21772 ( .C1(n18897), .C2(n18935), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18767), .ZN(n18768) );
  AOI211_X1 U21773 ( .C1(n18771), .C2(n18770), .A(n18769), .B(n18768), .ZN(
        n18772) );
  OAI221_X1 U21774 ( .B1(n18932), .B2(n18777), .C1(n18932), .C2(n18773), .A(
        n18772), .ZN(P3_U2996) );
  NAND2_X1 U21775 ( .A1(n18774), .A2(n18782), .ZN(n18785) );
  INV_X1 U21776 ( .A(n18775), .ZN(n18778) );
  NAND3_X1 U21777 ( .A1(n18778), .A2(n18777), .A3(n18776), .ZN(n18779) );
  NAND4_X1 U21778 ( .A1(n18781), .A2(n18780), .A3(n18785), .A4(n18779), .ZN(
        P3_U2997) );
  OR3_X1 U21779 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18783), .A3(n18782), 
        .ZN(n18784) );
  AND3_X1 U21780 ( .A1(n18785), .A2(n18876), .A3(n18784), .ZN(P3_U2998) );
  AND2_X1 U21781 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(
        P3_U2999) );
  AND2_X1 U21782 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(
        P3_U3000) );
  AND2_X1 U21783 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(
        P3_U3001) );
  AND2_X1 U21784 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_28__SCAN_IN), .ZN(
        P3_U3002) );
  AND2_X1 U21785 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(
        P3_U3003) );
  AND2_X1 U21786 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(
        P3_U3004) );
  AND2_X1 U21787 ( .A1(n18786), .A2(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(
        P3_U3005) );
  AND2_X1 U21788 ( .A1(n18786), .A2(P3_DATAWIDTH_REG_24__SCAN_IN), .ZN(
        P3_U3006) );
  AND2_X1 U21789 ( .A1(n18786), .A2(P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(
        P3_U3007) );
  AND2_X1 U21790 ( .A1(n18786), .A2(P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(
        P3_U3008) );
  AND2_X1 U21791 ( .A1(n18786), .A2(P3_DATAWIDTH_REG_20__SCAN_IN), .ZN(
        P3_U3010) );
  AND2_X1 U21792 ( .A1(n18786), .A2(P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(
        P3_U3011) );
  AND2_X1 U21793 ( .A1(n18786), .A2(P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(
        P3_U3012) );
  AND2_X1 U21794 ( .A1(n18786), .A2(P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(
        P3_U3013) );
  AND2_X1 U21795 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(
        P3_U3014) );
  AND2_X1 U21796 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(
        P3_U3015) );
  AND2_X1 U21797 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(
        P3_U3016) );
  AND2_X1 U21798 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(
        P3_U3017) );
  AND2_X1 U21799 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(
        P3_U3018) );
  AND2_X1 U21800 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(
        P3_U3019) );
  AND2_X1 U21801 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(
        P3_U3020) );
  AND2_X1 U21802 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(P3_U3021) );
  AND2_X1 U21803 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(P3_U3022) );
  AND2_X1 U21804 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(P3_U3023) );
  AND2_X1 U21805 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(P3_U3024) );
  AND2_X1 U21806 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(P3_U3025) );
  AND2_X1 U21807 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(P3_U3026) );
  AND2_X1 U21808 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(P3_U3027) );
  AND2_X1 U21809 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(P3_U3028) );
  NOR2_X1 U21810 ( .A1(n18787), .A2(n20873), .ZN(n18791) );
  NOR2_X1 U21811 ( .A1(n18807), .A2(n20873), .ZN(n18802) );
  INV_X1 U21812 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18937) );
  NOR3_X1 U21813 ( .A1(n18791), .A2(n18802), .A3(n18937), .ZN(n18790) );
  INV_X1 U21814 ( .A(NA), .ZN(n20883) );
  NAND2_X1 U21815 ( .A1(n9890), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18800) );
  INV_X1 U21816 ( .A(n18800), .ZN(n18798) );
  OAI21_X1 U21817 ( .B1(n18798), .B2(n18804), .A(n18807), .ZN(n18788) );
  OAI21_X1 U21818 ( .B1(n18792), .B2(n20883), .A(n18788), .ZN(n18805) );
  INV_X1 U21819 ( .A(n18805), .ZN(n18789) );
  OAI21_X1 U21820 ( .B1(n18939), .B2(n18790), .A(n18789), .ZN(P3_U3029) );
  AOI211_X1 U21821 ( .C1(n18791), .C2(n18807), .A(n18798), .B(n18799), .ZN(
        n18797) );
  OAI211_X1 U21822 ( .C1(n18793), .C2(n20873), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .B(n18792), .ZN(n18796) );
  AOI22_X1 U21823 ( .A1(n18797), .A2(n18796), .B1(n18795), .B2(n18794), .ZN(
        P3_U3030) );
  NOR2_X1 U21824 ( .A1(n18799), .A2(n18798), .ZN(n18806) );
  OAI22_X1 U21825 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18800), .ZN(n18801) );
  OAI22_X1 U21826 ( .A1(n18802), .A2(n18801), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18803) );
  OAI22_X1 U21827 ( .A1(n18806), .A2(n18805), .B1(n18804), .B2(n18803), .ZN(
        P3_U3031) );
  OAI222_X1 U21828 ( .A1(n18911), .A2(n18867), .B1(n18808), .B2(n18939), .C1(
        n18809), .C2(n18855), .ZN(P3_U3032) );
  OAI222_X1 U21829 ( .A1(n18855), .A2(n21123), .B1(n18810), .B2(n18939), .C1(
        n18809), .C2(n18867), .ZN(P3_U3033) );
  OAI222_X1 U21830 ( .A1(n21123), .A2(n18867), .B1(n18811), .B2(n18939), .C1(
        n18812), .C2(n18855), .ZN(P3_U3034) );
  OAI222_X1 U21831 ( .A1(n18855), .A2(n18815), .B1(n18813), .B2(n18939), .C1(
        n18812), .C2(n18867), .ZN(P3_U3035) );
  OAI222_X1 U21832 ( .A1(n18815), .A2(n18867), .B1(n18814), .B2(n18939), .C1(
        n18816), .C2(n18855), .ZN(P3_U3036) );
  OAI222_X1 U21833 ( .A1(n18855), .A2(n18818), .B1(n18817), .B2(n18939), .C1(
        n18816), .C2(n18867), .ZN(P3_U3037) );
  INV_X1 U21834 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18820) );
  OAI222_X1 U21835 ( .A1(n18855), .A2(n18820), .B1(n18819), .B2(n18939), .C1(
        n18818), .C2(n18867), .ZN(P3_U3038) );
  OAI222_X1 U21836 ( .A1(n18820), .A2(n18867), .B1(n21129), .B2(n18939), .C1(
        n18821), .C2(n18855), .ZN(P3_U3039) );
  OAI222_X1 U21837 ( .A1(n18855), .A2(n18823), .B1(n18822), .B2(n18939), .C1(
        n18821), .C2(n18867), .ZN(P3_U3040) );
  INV_X1 U21838 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18825) );
  OAI222_X1 U21839 ( .A1(n18855), .A2(n18825), .B1(n18824), .B2(n18939), .C1(
        n18823), .C2(n18867), .ZN(P3_U3041) );
  OAI222_X1 U21840 ( .A1(n18855), .A2(n18827), .B1(n18826), .B2(n18939), .C1(
        n18825), .C2(n18867), .ZN(P3_U3042) );
  OAI222_X1 U21841 ( .A1(n18855), .A2(n18829), .B1(n18828), .B2(n18939), .C1(
        n18827), .C2(n18867), .ZN(P3_U3043) );
  OAI222_X1 U21842 ( .A1(n18855), .A2(n18831), .B1(n18830), .B2(n18939), .C1(
        n18829), .C2(n18867), .ZN(P3_U3044) );
  OAI222_X1 U21843 ( .A1(n18855), .A2(n18833), .B1(n18832), .B2(n18939), .C1(
        n18831), .C2(n18867), .ZN(P3_U3045) );
  INV_X1 U21844 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18835) );
  OAI222_X1 U21845 ( .A1(n18855), .A2(n18835), .B1(n18834), .B2(n18939), .C1(
        n18833), .C2(n18867), .ZN(P3_U3046) );
  OAI222_X1 U21846 ( .A1(n18855), .A2(n18838), .B1(n18836), .B2(n18939), .C1(
        n18835), .C2(n18867), .ZN(P3_U3047) );
  OAI222_X1 U21847 ( .A1(n18838), .A2(n18867), .B1(n18837), .B2(n18939), .C1(
        n18839), .C2(n18855), .ZN(P3_U3048) );
  OAI222_X1 U21848 ( .A1(n18855), .A2(n18841), .B1(n18840), .B2(n18939), .C1(
        n18839), .C2(n18867), .ZN(P3_U3049) );
  OAI222_X1 U21849 ( .A1(n18855), .A2(n18844), .B1(n18842), .B2(n18939), .C1(
        n18841), .C2(n18867), .ZN(P3_U3050) );
  OAI222_X1 U21850 ( .A1(n18844), .A2(n18867), .B1(n18843), .B2(n18939), .C1(
        n18845), .C2(n18855), .ZN(P3_U3051) );
  OAI222_X1 U21851 ( .A1(n18855), .A2(n18847), .B1(n18846), .B2(n18939), .C1(
        n18845), .C2(n18867), .ZN(P3_U3052) );
  INV_X1 U21852 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18849) );
  OAI222_X1 U21853 ( .A1(n18855), .A2(n18849), .B1(n18848), .B2(n18939), .C1(
        n18847), .C2(n18867), .ZN(P3_U3053) );
  OAI222_X1 U21854 ( .A1(n18855), .A2(n18851), .B1(n18850), .B2(n18939), .C1(
        n18849), .C2(n18867), .ZN(P3_U3054) );
  OAI222_X1 U21855 ( .A1(n18855), .A2(n18853), .B1(n18852), .B2(n18939), .C1(
        n18851), .C2(n18867), .ZN(P3_U3055) );
  OAI222_X1 U21856 ( .A1(n18855), .A2(n18856), .B1(n18854), .B2(n18939), .C1(
        n18853), .C2(n18867), .ZN(P3_U3056) );
  OAI222_X1 U21857 ( .A1(n18855), .A2(n18858), .B1(n18857), .B2(n18939), .C1(
        n18856), .C2(n18867), .ZN(P3_U3057) );
  OAI222_X1 U21858 ( .A1(n18855), .A2(n18861), .B1(n18859), .B2(n18939), .C1(
        n18858), .C2(n18867), .ZN(P3_U3058) );
  OAI222_X1 U21859 ( .A1(n18861), .A2(n18867), .B1(n18860), .B2(n18939), .C1(
        n18862), .C2(n18855), .ZN(P3_U3059) );
  OAI222_X1 U21860 ( .A1(n18855), .A2(n18866), .B1(n18863), .B2(n18939), .C1(
        n18862), .C2(n18867), .ZN(P3_U3060) );
  OAI222_X1 U21861 ( .A1(n18867), .A2(n18866), .B1(n18865), .B2(n18939), .C1(
        n18864), .C2(n18855), .ZN(P3_U3061) );
  OAI22_X1 U21862 ( .A1(n18940), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18939), .ZN(n18868) );
  INV_X1 U21863 ( .A(n18868), .ZN(P3_U3274) );
  OAI22_X1 U21864 ( .A1(n18940), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18939), .ZN(n18869) );
  INV_X1 U21865 ( .A(n18869), .ZN(P3_U3275) );
  OAI22_X1 U21866 ( .A1(n18940), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18939), .ZN(n18870) );
  INV_X1 U21867 ( .A(n18870), .ZN(P3_U3276) );
  OAI22_X1 U21868 ( .A1(n18940), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18939), .ZN(n18871) );
  INV_X1 U21869 ( .A(n18871), .ZN(P3_U3277) );
  OAI21_X1 U21870 ( .B1(n18874), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18873), 
        .ZN(n18872) );
  INV_X1 U21871 ( .A(n18872), .ZN(P3_U3280) );
  OAI21_X1 U21872 ( .B1(n21132), .B2(n18874), .A(n18873), .ZN(P3_U3281) );
  INV_X1 U21873 ( .A(n18875), .ZN(n18877) );
  OAI221_X1 U21874 ( .B1(n18878), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18878), 
        .C2(n18877), .A(n18876), .ZN(P3_U3282) );
  NOR2_X1 U21875 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18904), .ZN(
        n18880) );
  AOI22_X1 U21876 ( .A1(n18897), .A2(n18881), .B1(n18880), .B2(n18879), .ZN(
        n18885) );
  AOI21_X1 U21877 ( .B1(n18898), .B2(n18882), .A(n18910), .ZN(n18884) );
  OAI22_X1 U21878 ( .A1(n18910), .A2(n18885), .B1(n18884), .B2(n18883), .ZN(
        P3_U3285) );
  NOR2_X1 U21879 ( .A1(n18905), .A2(n18886), .ZN(n18894) );
  OAI22_X1 U21880 ( .A1(n18887), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n9850), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18893) );
  AOI222_X1 U21881 ( .A1(n18889), .A2(n18898), .B1(n18894), .B2(n18893), .C1(
        n18897), .C2(n18888), .ZN(n18890) );
  INV_X1 U21882 ( .A(n18910), .ZN(n18907) );
  AOI22_X1 U21883 ( .A1(n18910), .A2(n18891), .B1(n18890), .B2(n18907), .ZN(
        P3_U3288) );
  INV_X1 U21884 ( .A(n18892), .ZN(n18899) );
  INV_X1 U21885 ( .A(n18893), .ZN(n18895) );
  AOI222_X1 U21886 ( .A1(n18899), .A2(n18898), .B1(n18897), .B2(n18896), .C1(
        n18895), .C2(n18894), .ZN(n18900) );
  AOI22_X1 U21887 ( .A1(n18910), .A2(n18901), .B1(n18900), .B2(n18907), .ZN(
        P3_U3289) );
  OAI222_X1 U21888 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18905), .B1(
        n18904), .B2(n18903), .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(
        n18902), .ZN(n18906) );
  INV_X1 U21889 ( .A(n18906), .ZN(n18908) );
  AOI22_X1 U21890 ( .A1(n18910), .A2(n18909), .B1(n18908), .B2(n18907), .ZN(
        P3_U3290) );
  AOI21_X1 U21891 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18912) );
  AOI22_X1 U21892 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18912), .B2(n18911), .ZN(n18914) );
  INV_X1 U21893 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18913) );
  AOI22_X1 U21894 ( .A1(n18915), .A2(n18914), .B1(n18913), .B2(n18917), .ZN(
        P3_U3292) );
  INV_X1 U21895 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18918) );
  NOR2_X1 U21896 ( .A1(n18917), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18916) );
  AOI22_X1 U21897 ( .A1(n18918), .A2(n18917), .B1(n18253), .B2(n18916), .ZN(
        P3_U3293) );
  INV_X1 U21898 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18919) );
  AOI22_X1 U21899 ( .A1(n18939), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18919), 
        .B2(n18940), .ZN(P3_U3294) );
  INV_X1 U21900 ( .A(n18920), .ZN(n18923) );
  NAND2_X1 U21901 ( .A1(n18923), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18921) );
  OAI21_X1 U21902 ( .B1(n18923), .B2(n18922), .A(n18921), .ZN(P3_U3295) );
  AOI21_X1 U21903 ( .B1(n18925), .B2(n18924), .A(n18945), .ZN(n18926) );
  OAI21_X1 U21904 ( .B1(n9890), .B2(n18927), .A(n18926), .ZN(n18938) );
  OAI21_X1 U21905 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18929), .A(n18928), 
        .ZN(n18931) );
  AOI211_X1 U21906 ( .C1(n18943), .C2(n18931), .A(n9890), .B(n18930), .ZN(
        n18933) );
  NOR2_X1 U21907 ( .A1(n18933), .A2(n18932), .ZN(n18934) );
  OAI21_X1 U21908 ( .B1(n18935), .B2(n18934), .A(n18938), .ZN(n18936) );
  OAI21_X1 U21909 ( .B1(n18938), .B2(n18937), .A(n18936), .ZN(P3_U3296) );
  OAI22_X1 U21910 ( .A1(n18940), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18939), .ZN(n18941) );
  INV_X1 U21911 ( .A(n18941), .ZN(P3_U3297) );
  OAI21_X1 U21912 ( .B1(n18946), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n18944), 
        .ZN(n18942) );
  OAI21_X1 U21913 ( .B1(n18944), .B2(n18943), .A(n18942), .ZN(P3_U3298) );
  NOR3_X1 U21914 ( .A1(P3_MEMORYFETCH_REG_SCAN_IN), .A2(n18946), .A3(n18945), 
        .ZN(n18948) );
  NOR2_X1 U21915 ( .A1(n18948), .A2(n18947), .ZN(P3_U3299) );
  INV_X1 U21916 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19951) );
  NAND2_X1 U21917 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19951), .ZN(n19941) );
  INV_X1 U21918 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18953) );
  AOI22_X1 U21919 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19941), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n18953), .ZN(n20004) );
  AOI21_X1 U21920 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20004), .ZN(n18949) );
  INV_X1 U21921 ( .A(n18949), .ZN(P2_U2815) );
  INV_X1 U21922 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18951) );
  OAI22_X1 U21923 ( .A1(n18952), .A2(n18951), .B1(n19926), .B2(n18950), .ZN(
        P2_U2816) );
  NAND2_X1 U21924 ( .A1(n18953), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20052) );
  INV_X2 U21925 ( .A(n20052), .ZN(n19995) );
  INV_X1 U21926 ( .A(n18955), .ZN(n19946) );
  NAND2_X1 U21927 ( .A1(n19946), .A2(n20052), .ZN(n19937) );
  AOI21_X1 U21928 ( .B1(n18953), .B2(n19937), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18954) );
  AOI21_X1 U21929 ( .B1(n19995), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n18954), 
        .ZN(P2_U2817) );
  OAI21_X1 U21930 ( .B1(n18955), .B2(BS16), .A(n20004), .ZN(n20002) );
  OAI21_X1 U21931 ( .B1(n20004), .B2(n19695), .A(n20002), .ZN(P2_U2818) );
  NOR2_X1 U21932 ( .A1(n18957), .A2(n18956), .ZN(n20050) );
  OAI21_X1 U21933 ( .B1(n20050), .B2(n12254), .A(n18958), .ZN(P2_U2819) );
  NOR4_X1 U21934 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18968) );
  NOR4_X1 U21935 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18967) );
  NOR4_X1 U21936 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18959) );
  INV_X1 U21937 ( .A(P2_DATAWIDTH_REG_20__SCAN_IN), .ZN(n19933) );
  INV_X1 U21938 ( .A(P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20975) );
  NAND3_X1 U21939 ( .A1(n18959), .A2(n19933), .A3(n20975), .ZN(n18965) );
  NOR4_X1 U21940 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18963) );
  NOR4_X1 U21941 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18962) );
  NOR4_X1 U21942 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18961) );
  NOR4_X1 U21943 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18960) );
  NAND4_X1 U21944 ( .A1(n18963), .A2(n18962), .A3(n18961), .A4(n18960), .ZN(
        n18964) );
  AOI211_X1 U21945 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n18965), .B(n18964), .ZN(n18966) );
  NAND3_X1 U21946 ( .A1(n18968), .A2(n18967), .A3(n18966), .ZN(n18975) );
  NOR2_X1 U21947 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18975), .ZN(n18970) );
  INV_X1 U21948 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20000) );
  AOI22_X1 U21949 ( .A1(n18970), .A2(n10440), .B1(n18975), .B2(n20000), .ZN(
        P2_U2820) );
  OR3_X1 U21950 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18974) );
  INV_X1 U21951 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18969) );
  AOI22_X1 U21952 ( .A1(n18970), .A2(n18974), .B1(n18975), .B2(n18969), .ZN(
        P2_U2821) );
  INV_X1 U21953 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20003) );
  NAND2_X1 U21954 ( .A1(n18970), .A2(n20003), .ZN(n18973) );
  INV_X1 U21955 ( .A(n18975), .ZN(n18977) );
  OAI21_X1 U21956 ( .B1(n10428), .B2(n10440), .A(n18977), .ZN(n18971) );
  OAI21_X1 U21957 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18977), .A(n18971), 
        .ZN(n18972) );
  OAI221_X1 U21958 ( .B1(n18973), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18973), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18972), .ZN(P2_U2822) );
  INV_X1 U21959 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18976) );
  OAI221_X1 U21960 ( .B1(n18977), .B2(n18976), .C1(n18975), .C2(n18974), .A(
        n18973), .ZN(P2_U2823) );
  OAI22_X1 U21961 ( .A1(n18979), .A2(n19174), .B1(n18978), .B2(n19154), .ZN(
        n18980) );
  INV_X1 U21962 ( .A(n18980), .ZN(n18989) );
  AOI211_X1 U21963 ( .C1(n18983), .C2(n18982), .A(n18981), .B(n19929), .ZN(
        n18987) );
  AOI22_X1 U21964 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n19183), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19170), .ZN(n18984) );
  OAI21_X1 U21965 ( .B1(n18985), .B2(n19194), .A(n18984), .ZN(n18986) );
  AOI211_X1 U21966 ( .C1(n19198), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n18987), .B(n18986), .ZN(n18988) );
  NAND2_X1 U21967 ( .A1(n18989), .A2(n18988), .ZN(P2_U2834) );
  OAI21_X1 U21968 ( .B1(n18991), .B2(n18990), .A(n19178), .ZN(n18999) );
  AOI22_X1 U21969 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19198), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19170), .ZN(n18992) );
  OAI21_X1 U21970 ( .B1(n18993), .B2(n19194), .A(n18992), .ZN(n18994) );
  AOI21_X1 U21971 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n19183), .A(n18994), .ZN(
        n18998) );
  AOI22_X1 U21972 ( .A1(n18996), .A2(n19190), .B1(n18995), .B2(n19185), .ZN(
        n18997) );
  OAI211_X1 U21973 ( .C1(n19000), .C2(n18999), .A(n18998), .B(n18997), .ZN(
        P2_U2835) );
  NAND2_X1 U21974 ( .A1(n19145), .A2(n19001), .ZN(n19002) );
  XOR2_X1 U21975 ( .A(n19003), .B(n19002), .Z(n19012) );
  AOI22_X1 U21976 ( .A1(n19004), .A2(n19153), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n19183), .ZN(n19005) );
  OAI211_X1 U21977 ( .C1(n19975), .C2(n19188), .A(n19005), .B(n19129), .ZN(
        n19006) );
  AOI21_X1 U21978 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19198), .A(
        n19006), .ZN(n19011) );
  OAI22_X1 U21979 ( .A1(n19008), .A2(n19174), .B1(n19007), .B2(n19154), .ZN(
        n19009) );
  INV_X1 U21980 ( .A(n19009), .ZN(n19010) );
  OAI211_X1 U21981 ( .C1(n19929), .C2(n19012), .A(n19011), .B(n19010), .ZN(
        P2_U2836) );
  NOR2_X1 U21982 ( .A1(n19162), .A2(n19013), .ZN(n19032) );
  XOR2_X1 U21983 ( .A(n19032), .B(n19014), .Z(n19022) );
  AOI22_X1 U21984 ( .A1(n19015), .A2(n19153), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19183), .ZN(n19016) );
  OAI211_X1 U21985 ( .C1(n10834), .C2(n19188), .A(n19016), .B(n19129), .ZN(
        n19017) );
  AOI21_X1 U21986 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19198), .A(
        n19017), .ZN(n19021) );
  AOI22_X1 U21987 ( .A1(n19019), .A2(n19190), .B1(n19018), .B2(n19185), .ZN(
        n19020) );
  OAI211_X1 U21988 ( .C1(n19929), .C2(n19022), .A(n19021), .B(n19020), .ZN(
        P2_U2837) );
  NAND2_X1 U21989 ( .A1(n19162), .A2(n19178), .ZN(n19182) );
  INV_X1 U21990 ( .A(n19028), .ZN(n19026) );
  OAI22_X1 U21991 ( .A1(n10239), .A2(n19097), .B1(n19972), .B2(n19188), .ZN(
        n19023) );
  AOI211_X1 U21992 ( .C1(n19024), .C2(n19153), .A(n19038), .B(n19023), .ZN(
        n19025) );
  OAI21_X1 U21993 ( .B1(n19182), .B2(n19026), .A(n19025), .ZN(n19027) );
  AOI21_X1 U21994 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n19183), .A(n19027), .ZN(
        n19034) );
  AOI21_X1 U21995 ( .B1(n19029), .B2(n19028), .A(n19929), .ZN(n19031) );
  AOI22_X1 U21996 ( .A1(n19032), .A2(n19031), .B1(n19030), .B2(n19190), .ZN(
        n19033) );
  OAI211_X1 U21997 ( .C1(n19035), .C2(n19154), .A(n19034), .B(n19033), .ZN(
        P2_U2838) );
  INV_X1 U21998 ( .A(n19182), .ZN(n19197) );
  NAND2_X1 U21999 ( .A1(n19197), .A2(n19044), .ZN(n19040) );
  OAI22_X1 U22000 ( .A1(n19036), .A2(n19097), .B1(n21116), .B2(n19188), .ZN(
        n19037) );
  NOR2_X1 U22001 ( .A1(n19038), .A2(n19037), .ZN(n19039) );
  OAI211_X1 U22002 ( .C1(n19194), .C2(n19041), .A(n19040), .B(n19039), .ZN(
        n19042) );
  AOI21_X1 U22003 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(n19183), .A(n19042), .ZN(
        n19049) );
  AOI21_X1 U22004 ( .B1(n19044), .B2(n19043), .A(n19929), .ZN(n19046) );
  AOI22_X1 U22005 ( .A1(n19047), .A2(n19046), .B1(n19045), .B2(n19190), .ZN(
        n19048) );
  OAI211_X1 U22006 ( .C1(n19218), .C2(n19154), .A(n19049), .B(n19048), .ZN(
        P2_U2840) );
  NOR2_X1 U22007 ( .A1(n19162), .A2(n19050), .ZN(n19052) );
  XOR2_X1 U22008 ( .A(n19052), .B(n19051), .Z(n19061) );
  INV_X1 U22009 ( .A(n19053), .ZN(n19055) );
  AOI22_X1 U22010 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19198), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19183), .ZN(n19054) );
  OAI21_X1 U22011 ( .B1(n19055), .B2(n19194), .A(n19054), .ZN(n19056) );
  AOI211_X1 U22012 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19170), .A(n19348), 
        .B(n19056), .ZN(n19060) );
  AOI22_X1 U22013 ( .A1(n19058), .A2(n19190), .B1(n19185), .B2(n19057), .ZN(
        n19059) );
  OAI211_X1 U22014 ( .C1(n19929), .C2(n19061), .A(n19060), .B(n19059), .ZN(
        P2_U2841) );
  NAND2_X1 U22015 ( .A1(n19145), .A2(n19062), .ZN(n19063) );
  XOR2_X1 U22016 ( .A(n19064), .B(n19063), .Z(n19073) );
  OAI21_X1 U22017 ( .B1(n19966), .B2(n19188), .A(n19129), .ZN(n19068) );
  OAI22_X1 U22018 ( .A1(n19066), .A2(n19194), .B1(n19156), .B2(n19065), .ZN(
        n19067) );
  AOI211_X1 U22019 ( .C1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n19198), .A(
        n19068), .B(n19067), .ZN(n19072) );
  OAI22_X1 U22020 ( .A1(n19069), .A2(n19174), .B1(n19223), .B2(n19154), .ZN(
        n19070) );
  INV_X1 U22021 ( .A(n19070), .ZN(n19071) );
  OAI211_X1 U22022 ( .C1(n19929), .C2(n19073), .A(n19072), .B(n19071), .ZN(
        P2_U2842) );
  INV_X1 U22023 ( .A(n19074), .ZN(n19076) );
  AOI22_X1 U22024 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19198), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n19183), .ZN(n19075) );
  OAI21_X1 U22025 ( .B1(n19076), .B2(n19194), .A(n19075), .ZN(n19077) );
  AOI211_X1 U22026 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19170), .A(n19348), 
        .B(n19077), .ZN(n19084) );
  NOR2_X1 U22027 ( .A1(n19162), .A2(n19078), .ZN(n19080) );
  XNOR2_X1 U22028 ( .A(n19080), .B(n19079), .ZN(n19082) );
  AOI22_X1 U22029 ( .A1(n19082), .A2(n19178), .B1(n19190), .B2(n19081), .ZN(
        n19083) );
  OAI211_X1 U22030 ( .C1(n19226), .C2(n19154), .A(n19084), .B(n19083), .ZN(
        P2_U2843) );
  AOI22_X1 U22031 ( .A1(n19085), .A2(n19153), .B1(P2_EBX_REG_11__SCAN_IN), 
        .B2(n19183), .ZN(n19086) );
  OAI21_X1 U22032 ( .B1(n19087), .B2(n19097), .A(n19086), .ZN(n19088) );
  AOI211_X1 U22033 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19170), .A(n19038), 
        .B(n19088), .ZN(n19095) );
  NAND2_X1 U22034 ( .A1(n19145), .A2(n19089), .ZN(n19091) );
  XNOR2_X1 U22035 ( .A(n19091), .B(n19090), .ZN(n19093) );
  AOI22_X1 U22036 ( .A1(n19093), .A2(n19178), .B1(n19190), .B2(n19092), .ZN(
        n19094) );
  OAI211_X1 U22037 ( .C1(n19228), .C2(n19154), .A(n19095), .B(n19094), .ZN(
        P2_U2844) );
  INV_X1 U22038 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19108) );
  INV_X1 U22039 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n19096) );
  OAI22_X1 U22040 ( .A1(n19098), .A2(n19194), .B1(n19097), .B2(n19096), .ZN(
        n19099) );
  AOI211_X1 U22041 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19170), .A(n19348), 
        .B(n19099), .ZN(n19107) );
  NOR2_X1 U22042 ( .A1(n19162), .A2(n19100), .ZN(n19101) );
  XNOR2_X1 U22043 ( .A(n19102), .B(n19101), .ZN(n19105) );
  OAI22_X1 U22044 ( .A1(n19103), .A2(n19174), .B1(n19154), .B2(n19231), .ZN(
        n19104) );
  AOI21_X1 U22045 ( .B1(n19105), .B2(n19178), .A(n19104), .ZN(n19106) );
  OAI211_X1 U22046 ( .C1(n19156), .C2(n19108), .A(n19107), .B(n19106), .ZN(
        P2_U2845) );
  NAND2_X1 U22047 ( .A1(n19145), .A2(n19109), .ZN(n19111) );
  XOR2_X1 U22048 ( .A(n19111), .B(n19110), .Z(n19118) );
  AOI22_X1 U22049 ( .A1(n19112), .A2(n19153), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19183), .ZN(n19113) );
  OAI211_X1 U22050 ( .C1(n10748), .C2(n19188), .A(n19113), .B(n19129), .ZN(
        n19116) );
  OAI22_X1 U22051 ( .A1(n19114), .A2(n19174), .B1(n19154), .B2(n19233), .ZN(
        n19115) );
  AOI211_X1 U22052 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19198), .A(
        n19116), .B(n19115), .ZN(n19117) );
  OAI21_X1 U22053 ( .B1(n19118), .B2(n19929), .A(n19117), .ZN(P2_U2846) );
  NAND2_X1 U22054 ( .A1(n19145), .A2(n19119), .ZN(n19121) );
  XOR2_X1 U22055 ( .A(n19121), .B(n19120), .Z(n19128) );
  AOI22_X1 U22056 ( .A1(n19122), .A2(n19153), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19183), .ZN(n19123) );
  OAI211_X1 U22057 ( .C1(n20984), .C2(n19188), .A(n19123), .B(n19129), .ZN(
        n19126) );
  OAI22_X1 U22058 ( .A1(n19124), .A2(n19174), .B1(n19238), .B2(n19154), .ZN(
        n19125) );
  AOI211_X1 U22059 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19198), .A(
        n19126), .B(n19125), .ZN(n19127) );
  OAI21_X1 U22060 ( .B1(n19128), .B2(n19929), .A(n19127), .ZN(P2_U2848) );
  OAI21_X1 U22061 ( .B1(n10493), .B2(n19188), .A(n19129), .ZN(n19133) );
  OAI22_X1 U22062 ( .A1(n19131), .A2(n19194), .B1(n19156), .B2(n19130), .ZN(
        n19132) );
  AOI211_X1 U22063 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19198), .A(
        n19133), .B(n19132), .ZN(n19140) );
  NOR2_X1 U22064 ( .A1(n19162), .A2(n19134), .ZN(n19136) );
  XNOR2_X1 U22065 ( .A(n19136), .B(n19135), .ZN(n19138) );
  AOI22_X1 U22066 ( .A1(n19138), .A2(n19178), .B1(n19190), .B2(n19137), .ZN(
        n19139) );
  OAI211_X1 U22067 ( .C1(n19154), .C2(n19240), .A(n19140), .B(n19139), .ZN(
        P2_U2849) );
  AOI22_X1 U22068 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19198), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19183), .ZN(n19141) );
  OAI21_X1 U22069 ( .B1(n19194), .B2(n19142), .A(n19141), .ZN(n19143) );
  AOI211_X1 U22070 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19170), .A(n19348), .B(
        n19143), .ZN(n19151) );
  NAND2_X1 U22071 ( .A1(n19145), .A2(n19144), .ZN(n19146) );
  XNOR2_X1 U22072 ( .A(n19147), .B(n19146), .ZN(n19149) );
  AOI22_X1 U22073 ( .A1(n19149), .A2(n19178), .B1(n19190), .B2(n19148), .ZN(
        n19150) );
  OAI211_X1 U22074 ( .C1(n19154), .C2(n19248), .A(n19151), .B(n19150), .ZN(
        P2_U2850) );
  AOI22_X1 U22075 ( .A1(n19153), .A2(n19152), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19198), .ZN(n19169) );
  OAI22_X1 U22076 ( .A1(n19156), .A2(n19155), .B1(n19154), .B2(n19250), .ZN(
        n19157) );
  AOI211_X1 U22077 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19170), .A(n19348), .B(
        n19157), .ZN(n19168) );
  OAI22_X1 U22078 ( .A1(n19252), .A2(n19159), .B1(n19174), .B2(n19158), .ZN(
        n19160) );
  INV_X1 U22079 ( .A(n19160), .ZN(n19167) );
  INV_X1 U22080 ( .A(n19358), .ZN(n19165) );
  NOR2_X1 U22081 ( .A1(n19162), .A2(n19161), .ZN(n19164) );
  AOI21_X1 U22082 ( .B1(n19165), .B2(n19164), .A(n19929), .ZN(n19163) );
  OAI21_X1 U22083 ( .B1(n19165), .B2(n19164), .A(n19163), .ZN(n19166) );
  NAND4_X1 U22084 ( .A1(n19169), .A2(n19168), .A3(n19167), .A4(n19166), .ZN(
        P2_U2851) );
  AOI22_X1 U22085 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19198), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19170), .ZN(n19172) );
  NAND2_X1 U22086 ( .A1(n19183), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n19171) );
  OAI211_X1 U22087 ( .C1(n19194), .C2(n19173), .A(n19172), .B(n19171), .ZN(
        n19177) );
  NOR2_X1 U22088 ( .A1(n19175), .A2(n19174), .ZN(n19176) );
  AOI211_X1 U22089 ( .C1(n19185), .C2(n20031), .A(n19177), .B(n19176), .ZN(
        n19181) );
  AOI22_X1 U22090 ( .A1(n19179), .A2(n19178), .B1(n19196), .B2(n20028), .ZN(
        n19180) );
  OAI211_X1 U22091 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19182), .A(
        n19181), .B(n19180), .ZN(P2_U2854) );
  NAND2_X1 U22092 ( .A1(n19183), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n19187) );
  NAND2_X1 U22093 ( .A1(n19185), .A2(n19184), .ZN(n19186) );
  OAI211_X1 U22094 ( .C1(n10440), .C2(n19188), .A(n19187), .B(n19186), .ZN(
        n19189) );
  AOI21_X1 U22095 ( .B1(n19191), .B2(n19190), .A(n19189), .ZN(n19192) );
  OAI21_X1 U22096 ( .B1(n19194), .B2(n19193), .A(n19192), .ZN(n19195) );
  AOI21_X1 U22097 ( .B1(n19629), .B2(n19196), .A(n19195), .ZN(n19200) );
  OAI21_X1 U22098 ( .B1(n19198), .B2(n19197), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19199) );
  OAI211_X1 U22099 ( .C1(n19201), .C2(n19929), .A(n19200), .B(n19199), .ZN(
        P2_U2855) );
  OR2_X1 U22100 ( .A1(n16277), .A2(n19215), .ZN(n19203) );
  NAND2_X1 U22101 ( .A1(n19209), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19202) );
  AND2_X1 U22102 ( .A1(n19203), .A2(n19202), .ZN(n19205) );
  AOI22_X1 U22103 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19264), .B1(n19208), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19204) );
  NAND2_X1 U22104 ( .A1(n19205), .A2(n19204), .ZN(P2_U2888) );
  AOI22_X1 U22105 ( .A1(n19207), .A2(n19206), .B1(n19264), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19214) );
  AOI22_X1 U22106 ( .A1(n19209), .A2(BUF2_REG_16__SCAN_IN), .B1(n19208), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19213) );
  AOI22_X1 U22107 ( .A1(n19211), .A2(n19269), .B1(n19265), .B2(n19210), .ZN(
        n19212) );
  NAND3_X1 U22108 ( .A1(n19214), .A2(n19213), .A3(n19212), .ZN(P2_U2903) );
  AND2_X1 U22109 ( .A1(n19216), .A2(n19215), .ZN(n19249) );
  OAI222_X1 U22110 ( .A1(n19218), .A2(n19249), .B1(n12637), .B2(n19239), .C1(
        n19217), .C2(n19273), .ZN(P2_U2904) );
  AOI22_X1 U22111 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19264), .B1(n19219), 
        .B2(n19241), .ZN(n19220) );
  OAI21_X1 U22112 ( .B1(n19249), .B2(n19221), .A(n19220), .ZN(P2_U2905) );
  INV_X1 U22113 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19318) );
  OAI222_X1 U22114 ( .A1(n19223), .A2(n19249), .B1(n19318), .B2(n19239), .C1(
        n19273), .C2(n19222), .ZN(P2_U2906) );
  AOI22_X1 U22115 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19264), .B1(n19224), 
        .B2(n19241), .ZN(n19225) );
  OAI21_X1 U22116 ( .B1(n19249), .B2(n19226), .A(n19225), .ZN(P2_U2907) );
  INV_X1 U22117 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19322) );
  OAI222_X1 U22118 ( .A1(n19228), .A2(n19249), .B1(n19322), .B2(n19239), .C1(
        n19273), .C2(n19227), .ZN(P2_U2908) );
  AOI22_X1 U22119 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19264), .B1(n19229), 
        .B2(n19241), .ZN(n19230) );
  OAI21_X1 U22120 ( .B1(n19249), .B2(n19231), .A(n19230), .ZN(P2_U2909) );
  INV_X1 U22121 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19327) );
  OAI222_X1 U22122 ( .A1(n19233), .A2(n19249), .B1(n19327), .B2(n19239), .C1(
        n19273), .C2(n19232), .ZN(P2_U2910) );
  INV_X1 U22123 ( .A(n19249), .ZN(n19235) );
  AOI22_X1 U22124 ( .A1(n19236), .A2(n19235), .B1(n19234), .B2(n19241), .ZN(
        n19237) );
  OAI21_X1 U22125 ( .B1(n19239), .B2(n20965), .A(n19237), .ZN(P2_U2911) );
  OAI222_X1 U22126 ( .A1(n19238), .A2(n19249), .B1(n19330), .B2(n19239), .C1(
        n19273), .C2(n19424), .ZN(P2_U2912) );
  OAI222_X1 U22127 ( .A1(n19240), .A2(n19249), .B1(n19333), .B2(n19239), .C1(
        n19273), .C2(n19412), .ZN(P2_U2913) );
  AOI22_X1 U22128 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19264), .B1(n19407), .B2(
        n19241), .ZN(n19247) );
  OAI21_X1 U22129 ( .B1(n20021), .B2(n19243), .A(n19242), .ZN(n19259) );
  XNOR2_X1 U22130 ( .A(n19630), .B(n19257), .ZN(n19260) );
  NAND2_X1 U22131 ( .A1(n19259), .A2(n19260), .ZN(n19258) );
  OAI21_X1 U22132 ( .B1(n20010), .B2(n19257), .A(n19258), .ZN(n19244) );
  NAND2_X1 U22133 ( .A1(n19244), .A2(n19250), .ZN(n19253) );
  INV_X1 U22134 ( .A(n19252), .ZN(n19245) );
  NAND3_X1 U22135 ( .A1(n19253), .A2(n19245), .A3(n19269), .ZN(n19246) );
  OAI211_X1 U22136 ( .C1(n19249), .C2(n19248), .A(n19247), .B(n19246), .ZN(
        P2_U2914) );
  INV_X1 U22137 ( .A(n19250), .ZN(n19251) );
  AOI22_X1 U22138 ( .A1(n19265), .A2(n19251), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19264), .ZN(n19256) );
  XNOR2_X1 U22139 ( .A(n19253), .B(n19252), .ZN(n19254) );
  NAND2_X1 U22140 ( .A1(n19254), .A2(n19269), .ZN(n19255) );
  OAI211_X1 U22141 ( .C1(n19402), .C2(n19273), .A(n19256), .B(n19255), .ZN(
        P2_U2915) );
  AOI22_X1 U22142 ( .A1(n19265), .A2(n19257), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19264), .ZN(n19263) );
  OAI21_X1 U22143 ( .B1(n19260), .B2(n19259), .A(n19258), .ZN(n19261) );
  NAND2_X1 U22144 ( .A1(n19261), .A2(n19269), .ZN(n19262) );
  OAI211_X1 U22145 ( .C1(n19398), .C2(n19273), .A(n19263), .B(n19262), .ZN(
        P2_U2916) );
  AOI22_X1 U22146 ( .A1(n19265), .A2(n20031), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19264), .ZN(n19272) );
  OAI21_X1 U22147 ( .B1(n19268), .B2(n19267), .A(n19266), .ZN(n19270) );
  NAND2_X1 U22148 ( .A1(n19270), .A2(n19269), .ZN(n19271) );
  OAI211_X1 U22149 ( .C1(n19392), .C2(n19273), .A(n19272), .B(n19271), .ZN(
        P2_U2918) );
  NAND2_X1 U22150 ( .A1(n19275), .A2(n19274), .ZN(n19277) );
  OAI21_X1 U22151 ( .B1(n19278), .B2(n19277), .A(n19276), .ZN(n19279) );
  AND2_X1 U22152 ( .A1(n19279), .A2(n19938), .ZN(n19313) );
  AND2_X1 U22153 ( .A1(n19331), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NAND2_X1 U22154 ( .A1(n19313), .A2(n19281), .ZN(n19311) );
  AOI22_X1 U22155 ( .A1(n19345), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n19282) );
  OAI21_X1 U22156 ( .B1(n19283), .B2(n19311), .A(n19282), .ZN(P2_U2921) );
  AOI22_X1 U22157 ( .A1(n19345), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19284) );
  OAI21_X1 U22158 ( .B1(n19285), .B2(n19311), .A(n19284), .ZN(P2_U2922) );
  AOI22_X1 U22159 ( .A1(n19345), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19331), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19286) );
  OAI21_X1 U22160 ( .B1(n19287), .B2(n19311), .A(n19286), .ZN(P2_U2923) );
  AOI22_X1 U22161 ( .A1(n19345), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19331), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19288) );
  OAI21_X1 U22162 ( .B1(n19289), .B2(n19311), .A(n19288), .ZN(P2_U2924) );
  AOI22_X1 U22163 ( .A1(n19345), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19331), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19290) );
  OAI21_X1 U22164 ( .B1(n19291), .B2(n19311), .A(n19290), .ZN(P2_U2925) );
  AOI22_X1 U22165 ( .A1(n19345), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19331), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19292) );
  OAI21_X1 U22166 ( .B1(n19293), .B2(n19311), .A(n19292), .ZN(P2_U2926) );
  AOI22_X1 U22167 ( .A1(n19345), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19331), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19294) );
  OAI21_X1 U22168 ( .B1(n19295), .B2(n19311), .A(n19294), .ZN(P2_U2927) );
  INV_X1 U22169 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19297) );
  AOI22_X1 U22170 ( .A1(n19345), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19296) );
  OAI21_X1 U22171 ( .B1(n19297), .B2(n19311), .A(n19296), .ZN(P2_U2928) );
  INV_X1 U22172 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19299) );
  AOI22_X1 U22173 ( .A1(n19345), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19298) );
  OAI21_X1 U22174 ( .B1(n19299), .B2(n19311), .A(n19298), .ZN(P2_U2929) );
  INV_X1 U22175 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19301) );
  AOI22_X1 U22176 ( .A1(n19345), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19300) );
  OAI21_X1 U22177 ( .B1(n19301), .B2(n19311), .A(n19300), .ZN(P2_U2930) );
  INV_X1 U22178 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19303) );
  AOI22_X1 U22179 ( .A1(n19345), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19302) );
  OAI21_X1 U22180 ( .B1(n19303), .B2(n19311), .A(n19302), .ZN(P2_U2931) );
  INV_X1 U22181 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19305) );
  AOI22_X1 U22182 ( .A1(n19345), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19304) );
  OAI21_X1 U22183 ( .B1(n19305), .B2(n19311), .A(n19304), .ZN(P2_U2932) );
  INV_X1 U22184 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19307) );
  AOI22_X1 U22185 ( .A1(n19325), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19306) );
  OAI21_X1 U22186 ( .B1(n19307), .B2(n19311), .A(n19306), .ZN(P2_U2933) );
  INV_X1 U22187 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19309) );
  AOI22_X1 U22188 ( .A1(n19325), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19308) );
  OAI21_X1 U22189 ( .B1(n19309), .B2(n19311), .A(n19308), .ZN(P2_U2934) );
  AOI22_X1 U22190 ( .A1(n19325), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19310) );
  OAI21_X1 U22191 ( .B1(n19312), .B2(n19311), .A(n19310), .ZN(P2_U2935) );
  AOI22_X1 U22192 ( .A1(n19325), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19314) );
  OAI21_X1 U22193 ( .B1(n12637), .B2(n19347), .A(n19314), .ZN(P2_U2936) );
  AOI22_X1 U22194 ( .A1(n19325), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19315) );
  OAI21_X1 U22195 ( .B1(n19316), .B2(n19347), .A(n19315), .ZN(P2_U2937) );
  AOI22_X1 U22196 ( .A1(n19325), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19317) );
  OAI21_X1 U22197 ( .B1(n19318), .B2(n19347), .A(n19317), .ZN(P2_U2938) );
  AOI22_X1 U22198 ( .A1(n19325), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19319) );
  OAI21_X1 U22199 ( .B1(n19320), .B2(n19347), .A(n19319), .ZN(P2_U2939) );
  AOI22_X1 U22200 ( .A1(n19325), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19321) );
  OAI21_X1 U22201 ( .B1(n19322), .B2(n19347), .A(n19321), .ZN(P2_U2940) );
  AOI22_X1 U22202 ( .A1(n19325), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19331), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19323) );
  OAI21_X1 U22203 ( .B1(n19324), .B2(n19347), .A(n19323), .ZN(P2_U2941) );
  AOI22_X1 U22204 ( .A1(n19325), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19331), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19326) );
  OAI21_X1 U22205 ( .B1(n19327), .B2(n19347), .A(n19326), .ZN(P2_U2942) );
  AOI22_X1 U22206 ( .A1(n19345), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19331), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19328) );
  OAI21_X1 U22207 ( .B1(n20965), .B2(n19347), .A(n19328), .ZN(P2_U2943) );
  AOI22_X1 U22208 ( .A1(n19345), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19331), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19329) );
  OAI21_X1 U22209 ( .B1(n19330), .B2(n19347), .A(n19329), .ZN(P2_U2944) );
  AOI22_X1 U22210 ( .A1(n19345), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19331), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19332) );
  OAI21_X1 U22211 ( .B1(n19333), .B2(n19347), .A(n19332), .ZN(P2_U2945) );
  INV_X1 U22212 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19335) );
  AOI22_X1 U22213 ( .A1(n19345), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19334) );
  OAI21_X1 U22214 ( .B1(n19335), .B2(n19347), .A(n19334), .ZN(P2_U2946) );
  INV_X1 U22215 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19337) );
  AOI22_X1 U22216 ( .A1(n19345), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19336) );
  OAI21_X1 U22217 ( .B1(n19337), .B2(n19347), .A(n19336), .ZN(P2_U2947) );
  INV_X1 U22218 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19339) );
  AOI22_X1 U22219 ( .A1(n19345), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19338) );
  OAI21_X1 U22220 ( .B1(n19339), .B2(n19347), .A(n19338), .ZN(P2_U2948) );
  INV_X1 U22221 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19341) );
  AOI22_X1 U22222 ( .A1(n19345), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19340) );
  OAI21_X1 U22223 ( .B1(n19341), .B2(n19347), .A(n19340), .ZN(P2_U2949) );
  INV_X1 U22224 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19343) );
  AOI22_X1 U22225 ( .A1(n19345), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19342) );
  OAI21_X1 U22226 ( .B1(n19343), .B2(n19347), .A(n19342), .ZN(P2_U2950) );
  AOI22_X1 U22227 ( .A1(n19345), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19344), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19346) );
  OAI21_X1 U22228 ( .B1(n12640), .B2(n19347), .A(n19346), .ZN(P2_U2951) );
  AOI22_X1 U22229 ( .A1(n19349), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19348), .ZN(n19357) );
  AOI222_X1 U22230 ( .A1(n19355), .A2(n19354), .B1(n19353), .B2(n19352), .C1(
        n19351), .C2(n19350), .ZN(n19356) );
  OAI211_X1 U22231 ( .C1(n19359), .C2(n19358), .A(n19357), .B(n19356), .ZN(
        P2_U3010) );
  AOI22_X1 U22232 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19362), .B1(
        n19361), .B2(n19360), .ZN(n19374) );
  AOI21_X1 U22233 ( .B1(n19364), .B2(n20031), .A(n19363), .ZN(n19365) );
  OAI21_X1 U22234 ( .B1(n19367), .B2(n19366), .A(n19365), .ZN(n19368) );
  AOI21_X1 U22235 ( .B1(n12728), .B2(n19369), .A(n19368), .ZN(n19373) );
  OAI211_X1 U22236 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n19371), .B(n19370), .ZN(n19372) );
  NAND3_X1 U22237 ( .A1(n19374), .A2(n19373), .A3(n19372), .ZN(P2_U3045) );
  AOI22_X1 U22238 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19415), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19416), .ZN(n19761) );
  AOI22_X1 U22239 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19415), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19416), .ZN(n19873) );
  INV_X1 U22240 ( .A(n19873), .ZN(n19758) );
  AND2_X1 U22241 ( .A1(n19378), .A2(n19421), .ZN(n19861) );
  NAND2_X1 U22242 ( .A1(n10561), .A2(n20023), .ZN(n19481) );
  INV_X1 U22243 ( .A(n19481), .ZN(n19482) );
  NAND2_X1 U22244 ( .A1(n19482), .A2(n20033), .ZN(n19430) );
  NOR2_X1 U22245 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19430), .ZN(
        n19423) );
  AOI22_X1 U22246 ( .A1(n19758), .A2(n19917), .B1(n19861), .B2(n19423), .ZN(
        n19391) );
  INV_X1 U22247 ( .A(n19454), .ZN(n19379) );
  OAI21_X1 U22248 ( .B1(n19917), .B2(n19379), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19380) );
  NAND2_X1 U22249 ( .A1(n19380), .A2(n20006), .ZN(n19389) );
  NOR2_X1 U22250 ( .A1(n19913), .A2(n19423), .ZN(n19388) );
  INV_X1 U22251 ( .A(n19388), .ZN(n19384) );
  INV_X1 U22252 ( .A(n12142), .ZN(n19386) );
  INV_X1 U22253 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19632) );
  OAI21_X1 U22254 ( .B1(n19386), .B2(n20035), .A(n19632), .ZN(n19382) );
  INV_X1 U22255 ( .A(n19423), .ZN(n19381) );
  AOI21_X1 U22256 ( .B1(n19382), .B2(n19381), .A(n19754), .ZN(n19383) );
  NOR2_X2 U22257 ( .A1(n19385), .A2(n19754), .ZN(n19862) );
  OAI21_X1 U22258 ( .B1(n19386), .B2(n19423), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19387) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19426), .B1(
        n19862), .B2(n19425), .ZN(n19390) );
  OAI211_X1 U22260 ( .C1(n19761), .C2(n19454), .A(n19391), .B(n19390), .ZN(
        P2_U3048) );
  AOI22_X1 U22261 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19415), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19416), .ZN(n19832) );
  AOI22_X1 U22262 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19415), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19416), .ZN(n19879) );
  AOI22_X1 U22263 ( .A1(n19829), .A2(n19917), .B1(n19874), .B2(n19423), .ZN(
        n19394) );
  NOR2_X2 U22264 ( .A1(n19392), .A2(n19754), .ZN(n19875) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19426), .B1(
        n19875), .B2(n19425), .ZN(n19393) );
  OAI211_X1 U22266 ( .C1(n19832), .C2(n19454), .A(n19394), .B(n19393), .ZN(
        P2_U3049) );
  AOI22_X1 U22267 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19415), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19416), .ZN(n19836) );
  AOI22_X1 U22268 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19415), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19416), .ZN(n19885) );
  INV_X1 U22269 ( .A(n19885), .ZN(n19833) );
  NOR2_X2 U22270 ( .A1(n10407), .A2(n19401), .ZN(n19880) );
  AOI22_X1 U22271 ( .A1(n19833), .A2(n19917), .B1(n19880), .B2(n19423), .ZN(
        n19397) );
  NOR2_X2 U22272 ( .A1(n19395), .A2(n19754), .ZN(n19881) );
  AOI22_X1 U22273 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19426), .B1(
        n19881), .B2(n19425), .ZN(n19396) );
  OAI211_X1 U22274 ( .C1(n19836), .C2(n19454), .A(n19397), .B(n19396), .ZN(
        P2_U3050) );
  AOI22_X1 U22275 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19415), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19416), .ZN(n19840) );
  AOI22_X1 U22276 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19415), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19416), .ZN(n19891) );
  AND2_X1 U22277 ( .A1(n10397), .A2(n19421), .ZN(n19886) );
  AOI22_X1 U22278 ( .A1(n19837), .A2(n19917), .B1(n19886), .B2(n19423), .ZN(
        n19400) );
  NOR2_X2 U22279 ( .A1(n19398), .A2(n19754), .ZN(n19887) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19426), .B1(
        n19887), .B2(n19425), .ZN(n19399) );
  OAI211_X1 U22281 ( .C1(n19840), .C2(n19454), .A(n19400), .B(n19399), .ZN(
        P2_U3051) );
  AOI22_X1 U22282 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19415), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19416), .ZN(n19897) );
  AOI22_X1 U22283 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19416), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19415), .ZN(n19844) );
  INV_X1 U22284 ( .A(n19844), .ZN(n19894) );
  NOR2_X2 U22285 ( .A1(n12237), .A2(n19401), .ZN(n19892) );
  AOI22_X1 U22286 ( .A1(n19894), .A2(n19917), .B1(n19892), .B2(n19423), .ZN(
        n19404) );
  NOR2_X2 U22287 ( .A1(n19402), .A2(n19754), .ZN(n19893) );
  AOI22_X1 U22288 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19426), .B1(
        n19893), .B2(n19425), .ZN(n19403) );
  OAI211_X1 U22289 ( .C1(n19897), .C2(n19454), .A(n19404), .B(n19403), .ZN(
        P2_U3052) );
  INV_X1 U22290 ( .A(n19415), .ZN(n19419) );
  INV_X1 U22291 ( .A(n19416), .ZN(n19417) );
  AOI22_X1 U22292 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19416), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19415), .ZN(n19803) );
  AOI22_X1 U22293 ( .A1(n19900), .A2(n19917), .B1(n19898), .B2(n19423), .ZN(
        n19410) );
  INV_X1 U22294 ( .A(n19407), .ZN(n19408) );
  NOR2_X2 U22295 ( .A1(n19408), .A2(n19754), .ZN(n19899) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19426), .B1(
        n19899), .B2(n19425), .ZN(n19409) );
  OAI211_X1 U22297 ( .C1(n19905), .C2(n19454), .A(n19410), .B(n19409), .ZN(
        P2_U3053) );
  AOI22_X1 U22298 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19415), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19416), .ZN(n19808) );
  AOI22_X1 U22299 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19416), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19415), .ZN(n19911) );
  INV_X1 U22300 ( .A(n19911), .ZN(n19804) );
  AND2_X1 U22301 ( .A1(n19411), .A2(n19421), .ZN(n19906) );
  AOI22_X1 U22302 ( .A1(n19804), .A2(n19917), .B1(n19906), .B2(n19423), .ZN(
        n19414) );
  NOR2_X2 U22303 ( .A1(n19412), .A2(n19754), .ZN(n19907) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19426), .B1(
        n19907), .B2(n19425), .ZN(n19413) );
  OAI211_X1 U22305 ( .C1(n19808), .C2(n19454), .A(n19414), .B(n19413), .ZN(
        P2_U3054) );
  AOI22_X1 U22306 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19416), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19415), .ZN(n19857) );
  AND2_X1 U22307 ( .A1(n19422), .A2(n19421), .ZN(n19912) );
  AOI22_X1 U22308 ( .A1(n19852), .A2(n19917), .B1(n19912), .B2(n19423), .ZN(
        n19428) );
  NOR2_X2 U22309 ( .A1(n19754), .A2(n19424), .ZN(n19914) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19426), .B1(
        n19914), .B2(n19425), .ZN(n19427) );
  OAI211_X1 U22311 ( .C1(n19857), .C2(n19454), .A(n19428), .B(n19427), .ZN(
        P2_U3055) );
  NAND2_X1 U22312 ( .A1(n20033), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19661) );
  NOR2_X1 U22313 ( .A1(n19661), .A2(n19481), .ZN(n19449) );
  NOR3_X1 U22314 ( .A1(n19429), .A2(n19449), .A3(n20035), .ZN(n19431) );
  AOI211_X2 U22315 ( .C1(n19430), .C2(n20035), .A(n19602), .B(n19431), .ZN(
        n19450) );
  AOI22_X1 U22316 ( .A1(n19450), .A2(n19862), .B1(n19861), .B2(n19449), .ZN(
        n19436) );
  AND2_X1 U22317 ( .A1(n19630), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19604) );
  INV_X1 U22318 ( .A(n19604), .ZN(n19544) );
  OAI21_X1 U22319 ( .B1(n19544), .B2(n19662), .A(n19430), .ZN(n19434) );
  INV_X1 U22320 ( .A(n19449), .ZN(n19432) );
  AOI211_X1 U22321 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19432), .A(n19754), 
        .B(n19431), .ZN(n19433) );
  NAND2_X1 U22322 ( .A1(n19434), .A2(n19433), .ZN(n19451) );
  NOR2_X2 U22323 ( .A1(n19662), .A2(n19608), .ZN(n19477) );
  INV_X1 U22324 ( .A(n19761), .ZN(n19870) );
  AOI22_X1 U22325 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19451), .B1(
        n19477), .B2(n19870), .ZN(n19435) );
  OAI211_X1 U22326 ( .C1(n19873), .C2(n19454), .A(n19436), .B(n19435), .ZN(
        P2_U3056) );
  AOI22_X1 U22327 ( .A1(n19450), .A2(n19875), .B1(n19874), .B2(n19449), .ZN(
        n19438) );
  INV_X1 U22328 ( .A(n19832), .ZN(n19876) );
  AOI22_X1 U22329 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19451), .B1(
        n19477), .B2(n19876), .ZN(n19437) );
  OAI211_X1 U22330 ( .C1(n19879), .C2(n19454), .A(n19438), .B(n19437), .ZN(
        P2_U3057) );
  AOI22_X1 U22331 ( .A1(n19450), .A2(n19881), .B1(n19880), .B2(n19449), .ZN(
        n19440) );
  INV_X1 U22332 ( .A(n19836), .ZN(n19882) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19451), .B1(
        n19477), .B2(n19882), .ZN(n19439) );
  OAI211_X1 U22334 ( .C1(n19885), .C2(n19454), .A(n19440), .B(n19439), .ZN(
        P2_U3058) );
  AOI22_X1 U22335 ( .A1(n19450), .A2(n19887), .B1(n19886), .B2(n19449), .ZN(
        n19442) );
  INV_X1 U22336 ( .A(n19840), .ZN(n19888) );
  AOI22_X1 U22337 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19451), .B1(
        n19477), .B2(n19888), .ZN(n19441) );
  OAI211_X1 U22338 ( .C1(n19891), .C2(n19454), .A(n19442), .B(n19441), .ZN(
        P2_U3059) );
  AOI22_X1 U22339 ( .A1(n19450), .A2(n19893), .B1(n19892), .B2(n19449), .ZN(
        n19444) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19451), .B1(
        n19477), .B2(n19841), .ZN(n19443) );
  OAI211_X1 U22341 ( .C1(n19844), .C2(n19454), .A(n19444), .B(n19443), .ZN(
        P2_U3060) );
  AOI22_X1 U22342 ( .A1(n19450), .A2(n19899), .B1(n19898), .B2(n19449), .ZN(
        n19446) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19451), .B1(
        n19477), .B2(n19800), .ZN(n19445) );
  OAI211_X1 U22344 ( .C1(n19803), .C2(n19454), .A(n19446), .B(n19445), .ZN(
        P2_U3061) );
  AOI22_X1 U22345 ( .A1(n19450), .A2(n19907), .B1(n19906), .B2(n19449), .ZN(
        n19448) );
  INV_X1 U22346 ( .A(n19808), .ZN(n19908) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19451), .B1(
        n19477), .B2(n19908), .ZN(n19447) );
  OAI211_X1 U22348 ( .C1(n19911), .C2(n19454), .A(n19448), .B(n19447), .ZN(
        P2_U3062) );
  AOI22_X1 U22349 ( .A1(n19450), .A2(n19914), .B1(n19912), .B2(n19449), .ZN(
        n19453) );
  INV_X1 U22350 ( .A(n19857), .ZN(n19916) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19451), .B1(
        n19477), .B2(n19916), .ZN(n19452) );
  OAI211_X1 U22352 ( .C1(n19922), .C2(n19454), .A(n19453), .B(n19452), .ZN(
        P2_U3063) );
  NOR2_X1 U22353 ( .A1(n20033), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19691) );
  NAND2_X1 U22354 ( .A1(n19691), .A2(n19482), .ZN(n19456) );
  AND2_X1 U22355 ( .A1(n12168), .A2(n19456), .ZN(n19455) );
  NAND2_X1 U22356 ( .A1(n19513), .A2(n19482), .ZN(n19458) );
  OAI22_X1 U22357 ( .A1(n19455), .A2(n20035), .B1(n19819), .B2(n19458), .ZN(
        n19476) );
  INV_X1 U22358 ( .A(n19456), .ZN(n19475) );
  AOI22_X1 U22359 ( .A1(n19476), .A2(n19862), .B1(n19861), .B2(n19475), .ZN(
        n19462) );
  AOI21_X1 U22360 ( .B1(n12168), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19460) );
  OAI21_X1 U22361 ( .B1(n19507), .B2(n19477), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19457) );
  NAND2_X1 U22362 ( .A1(n19458), .A2(n19457), .ZN(n19459) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19478), .B1(
        n19477), .B2(n19758), .ZN(n19461) );
  OAI211_X1 U22364 ( .C1(n19761), .C2(n19503), .A(n19462), .B(n19461), .ZN(
        P2_U3064) );
  AOI22_X1 U22365 ( .A1(n19476), .A2(n19875), .B1(n19874), .B2(n19475), .ZN(
        n19464) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19478), .B1(
        n19477), .B2(n19829), .ZN(n19463) );
  OAI211_X1 U22367 ( .C1(n19832), .C2(n19503), .A(n19464), .B(n19463), .ZN(
        P2_U3065) );
  AOI22_X1 U22368 ( .A1(n19476), .A2(n19881), .B1(n19880), .B2(n19475), .ZN(
        n19466) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19478), .B1(
        n19477), .B2(n19833), .ZN(n19465) );
  OAI211_X1 U22370 ( .C1(n19836), .C2(n19503), .A(n19466), .B(n19465), .ZN(
        P2_U3066) );
  AOI22_X1 U22371 ( .A1(n19476), .A2(n19887), .B1(n19886), .B2(n19475), .ZN(
        n19468) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19478), .B1(
        n19477), .B2(n19837), .ZN(n19467) );
  OAI211_X1 U22373 ( .C1(n19840), .C2(n19503), .A(n19468), .B(n19467), .ZN(
        P2_U3067) );
  AOI22_X1 U22374 ( .A1(n19476), .A2(n19893), .B1(n19892), .B2(n19475), .ZN(
        n19470) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19478), .B1(
        n19477), .B2(n19894), .ZN(n19469) );
  OAI211_X1 U22376 ( .C1(n19897), .C2(n19503), .A(n19470), .B(n19469), .ZN(
        P2_U3068) );
  AOI22_X1 U22377 ( .A1(n19476), .A2(n19899), .B1(n19898), .B2(n19475), .ZN(
        n19472) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19478), .B1(
        n19477), .B2(n19900), .ZN(n19471) );
  OAI211_X1 U22379 ( .C1(n19905), .C2(n19503), .A(n19472), .B(n19471), .ZN(
        P2_U3069) );
  AOI22_X1 U22380 ( .A1(n19476), .A2(n19907), .B1(n19906), .B2(n19475), .ZN(
        n19474) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19478), .B1(
        n19477), .B2(n19804), .ZN(n19473) );
  OAI211_X1 U22382 ( .C1(n19808), .C2(n19503), .A(n19474), .B(n19473), .ZN(
        P2_U3070) );
  AOI22_X1 U22383 ( .A1(n19476), .A2(n19914), .B1(n19912), .B2(n19475), .ZN(
        n19480) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19478), .B1(
        n19477), .B2(n19852), .ZN(n19479) );
  OAI211_X1 U22385 ( .C1(n19857), .C2(n19503), .A(n19480), .B(n19479), .ZN(
        P2_U3071) );
  NOR2_X2 U22386 ( .A1(n19608), .A2(n20007), .ZN(n19540) );
  NOR2_X1 U22387 ( .A1(n19722), .A2(n19481), .ZN(n19506) );
  AOI22_X1 U22388 ( .A1(n19870), .A2(n19540), .B1(n19506), .B2(n19861), .ZN(
        n19492) );
  OAI21_X1 U22389 ( .B1(n19544), .B2(n20007), .A(n20006), .ZN(n19490) );
  NAND2_X1 U22390 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19482), .ZN(
        n19489) );
  INV_X1 U22391 ( .A(n19489), .ZN(n19486) );
  NAND2_X1 U22392 ( .A1(n19487), .A2(n19632), .ZN(n19484) );
  INV_X1 U22393 ( .A(n19506), .ZN(n19483) );
  NAND3_X1 U22394 ( .A1(n19484), .A2(n19819), .A3(n19483), .ZN(n19485) );
  OAI211_X1 U22395 ( .C1(n19490), .C2(n19486), .A(n19868), .B(n19485), .ZN(
        n19509) );
  OAI21_X1 U22396 ( .B1(n19487), .B2(n19506), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19488) );
  OAI21_X1 U22397 ( .B1(n19490), .B2(n19489), .A(n19488), .ZN(n19508) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19509), .B1(
        n19862), .B2(n19508), .ZN(n19491) );
  OAI211_X1 U22399 ( .C1(n19873), .C2(n19503), .A(n19492), .B(n19491), .ZN(
        P2_U3072) );
  INV_X1 U22400 ( .A(n19540), .ZN(n19517) );
  AOI22_X1 U22401 ( .A1(n19829), .A2(n19507), .B1(n19506), .B2(n19874), .ZN(
        n19494) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19509), .B1(
        n19875), .B2(n19508), .ZN(n19493) );
  OAI211_X1 U22403 ( .C1(n19832), .C2(n19517), .A(n19494), .B(n19493), .ZN(
        P2_U3073) );
  AOI22_X1 U22404 ( .A1(n19882), .A2(n19540), .B1(n19506), .B2(n19880), .ZN(
        n19496) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19509), .B1(
        n19881), .B2(n19508), .ZN(n19495) );
  OAI211_X1 U22406 ( .C1(n19885), .C2(n19503), .A(n19496), .B(n19495), .ZN(
        P2_U3074) );
  AOI22_X1 U22407 ( .A1(n19888), .A2(n19540), .B1(n19506), .B2(n19886), .ZN(
        n19498) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19509), .B1(
        n19887), .B2(n19508), .ZN(n19497) );
  OAI211_X1 U22409 ( .C1(n19891), .C2(n19503), .A(n19498), .B(n19497), .ZN(
        P2_U3075) );
  AOI22_X1 U22410 ( .A1(n19841), .A2(n19540), .B1(n19506), .B2(n19892), .ZN(
        n19500) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19509), .B1(
        n19893), .B2(n19508), .ZN(n19499) );
  OAI211_X1 U22412 ( .C1(n19844), .C2(n19503), .A(n19500), .B(n19499), .ZN(
        P2_U3076) );
  AOI22_X1 U22413 ( .A1(n19800), .A2(n19540), .B1(n19506), .B2(n19898), .ZN(
        n19502) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19509), .B1(
        n19899), .B2(n19508), .ZN(n19501) );
  OAI211_X1 U22415 ( .C1(n19803), .C2(n19503), .A(n19502), .B(n19501), .ZN(
        P2_U3077) );
  AOI22_X1 U22416 ( .A1(n19804), .A2(n19507), .B1(n19506), .B2(n19906), .ZN(
        n19505) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19509), .B1(
        n19907), .B2(n19508), .ZN(n19504) );
  OAI211_X1 U22418 ( .C1(n19808), .C2(n19517), .A(n19505), .B(n19504), .ZN(
        P2_U3078) );
  AOI22_X1 U22419 ( .A1(n19852), .A2(n19507), .B1(n19506), .B2(n19912), .ZN(
        n19511) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19509), .B1(
        n19914), .B2(n19508), .ZN(n19510) );
  OAI211_X1 U22421 ( .C1(n19857), .C2(n19517), .A(n19511), .B(n19510), .ZN(
        P2_U3079) );
  NOR3_X1 U22422 ( .A1(n20023), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19548) );
  NAND2_X1 U22423 ( .A1(n20042), .A2(n19548), .ZN(n19518) );
  AND2_X1 U22424 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19518), .ZN(n19512) );
  NAND2_X1 U22425 ( .A1(n12134), .A2(n19512), .ZN(n19520) );
  NOR2_X1 U22426 ( .A1(n19514), .A2(n19513), .ZN(n19750) );
  NAND2_X1 U22427 ( .A1(n19750), .A2(n10561), .ZN(n19516) );
  AOI21_X1 U22428 ( .B1(n19516), .B2(n20035), .A(n19602), .ZN(n19515) );
  INV_X1 U22429 ( .A(n19518), .ZN(n19538) );
  AOI22_X1 U22430 ( .A1(n19539), .A2(n19862), .B1(n19861), .B2(n19538), .ZN(
        n19525) );
  INV_X1 U22431 ( .A(n19516), .ZN(n19523) );
  AOI21_X1 U22432 ( .B1(n19517), .B2(n19571), .A(n19695), .ZN(n19522) );
  NAND2_X1 U22433 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19518), .ZN(n19519) );
  AND3_X1 U22434 ( .A1(n19520), .A2(n19868), .A3(n19519), .ZN(n19521) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19758), .ZN(n19524) );
  OAI211_X1 U22436 ( .C1(n19761), .C2(n19571), .A(n19525), .B(n19524), .ZN(
        P2_U3080) );
  AOI22_X1 U22437 ( .A1(n19539), .A2(n19875), .B1(n19874), .B2(n19538), .ZN(
        n19527) );
  AOI22_X1 U22438 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19829), .ZN(n19526) );
  OAI211_X1 U22439 ( .C1(n19832), .C2(n19571), .A(n19527), .B(n19526), .ZN(
        P2_U3081) );
  AOI22_X1 U22440 ( .A1(n19539), .A2(n19881), .B1(n19880), .B2(n19538), .ZN(
        n19529) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19833), .ZN(n19528) );
  OAI211_X1 U22442 ( .C1(n19836), .C2(n19571), .A(n19529), .B(n19528), .ZN(
        P2_U3082) );
  AOI22_X1 U22443 ( .A1(n19539), .A2(n19887), .B1(n19886), .B2(n19538), .ZN(
        n19531) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19837), .ZN(n19530) );
  OAI211_X1 U22445 ( .C1(n19840), .C2(n19571), .A(n19531), .B(n19530), .ZN(
        P2_U3083) );
  AOI22_X1 U22446 ( .A1(n19539), .A2(n19893), .B1(n19892), .B2(n19538), .ZN(
        n19533) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19894), .ZN(n19532) );
  OAI211_X1 U22448 ( .C1(n19897), .C2(n19571), .A(n19533), .B(n19532), .ZN(
        P2_U3084) );
  AOI22_X1 U22449 ( .A1(n19539), .A2(n19899), .B1(n19898), .B2(n19538), .ZN(
        n19535) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19900), .ZN(n19534) );
  OAI211_X1 U22451 ( .C1(n19905), .C2(n19571), .A(n19535), .B(n19534), .ZN(
        P2_U3085) );
  AOI22_X1 U22452 ( .A1(n19539), .A2(n19907), .B1(n19906), .B2(n19538), .ZN(
        n19537) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19804), .ZN(n19536) );
  OAI211_X1 U22454 ( .C1(n19808), .C2(n19571), .A(n19537), .B(n19536), .ZN(
        P2_U3086) );
  AOI22_X1 U22455 ( .A1(n19539), .A2(n19914), .B1(n19912), .B2(n19538), .ZN(
        n19543) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19852), .ZN(n19542) );
  OAI211_X1 U22457 ( .C1(n19857), .C2(n19571), .A(n19543), .B(n19542), .ZN(
        P2_U3087) );
  INV_X1 U22458 ( .A(n19548), .ZN(n19550) );
  NOR2_X1 U22459 ( .A1(n20042), .A2(n19550), .ZN(n19576) );
  AOI22_X1 U22460 ( .A1(n19870), .A2(n19590), .B1(n9784), .B2(n19861), .ZN(
        n19553) );
  OAI21_X1 U22461 ( .B1(n19544), .B2(n19788), .A(n20006), .ZN(n19551) );
  NAND2_X1 U22462 ( .A1(n12154), .A2(n19632), .ZN(n19546) );
  INV_X1 U22463 ( .A(n19576), .ZN(n19545) );
  NAND3_X1 U22464 ( .A1(n19546), .A2(n19819), .A3(n19545), .ZN(n19547) );
  OAI211_X1 U22465 ( .C1(n19551), .C2(n19548), .A(n19868), .B(n19547), .ZN(
        n19568) );
  OAI21_X1 U22466 ( .B1(n12154), .B2(n19576), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19549) );
  OAI21_X1 U22467 ( .B1(n19551), .B2(n19550), .A(n19549), .ZN(n19567) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19568), .B1(
        n19862), .B2(n19567), .ZN(n19552) );
  OAI211_X1 U22469 ( .C1(n19873), .C2(n19571), .A(n19553), .B(n19552), .ZN(
        P2_U3088) );
  AOI22_X1 U22470 ( .A1(n19829), .A2(n19558), .B1(n19874), .B2(n9784), .ZN(
        n19555) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19568), .B1(
        n19875), .B2(n19567), .ZN(n19554) );
  OAI211_X1 U22472 ( .C1(n19832), .C2(n19600), .A(n19555), .B(n19554), .ZN(
        P2_U3089) );
  AOI22_X1 U22473 ( .A1(n19833), .A2(n19558), .B1(n9784), .B2(n19880), .ZN(
        n19557) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19568), .B1(
        n19881), .B2(n19567), .ZN(n19556) );
  OAI211_X1 U22475 ( .C1(n19836), .C2(n19600), .A(n19557), .B(n19556), .ZN(
        P2_U3090) );
  AOI22_X1 U22476 ( .A1(n19837), .A2(n19558), .B1(n9784), .B2(n19886), .ZN(
        n19560) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19568), .B1(
        n19887), .B2(n19567), .ZN(n19559) );
  OAI211_X1 U22478 ( .C1(n19840), .C2(n19600), .A(n19560), .B(n19559), .ZN(
        P2_U3091) );
  AOI22_X1 U22479 ( .A1(n19841), .A2(n19590), .B1(n9784), .B2(n19892), .ZN(
        n19562) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19568), .B1(
        n19893), .B2(n19567), .ZN(n19561) );
  OAI211_X1 U22481 ( .C1(n19844), .C2(n19571), .A(n19562), .B(n19561), .ZN(
        P2_U3092) );
  AOI22_X1 U22482 ( .A1(n19800), .A2(n19590), .B1(n9784), .B2(n19898), .ZN(
        n19564) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19568), .B1(
        n19899), .B2(n19567), .ZN(n19563) );
  OAI211_X1 U22484 ( .C1(n19803), .C2(n19571), .A(n19564), .B(n19563), .ZN(
        P2_U3093) );
  AOI22_X1 U22485 ( .A1(n19908), .A2(n19590), .B1(n9784), .B2(n19906), .ZN(
        n19566) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19568), .B1(
        n19907), .B2(n19567), .ZN(n19565) );
  OAI211_X1 U22487 ( .C1(n19911), .C2(n19571), .A(n19566), .B(n19565), .ZN(
        P2_U3094) );
  AOI22_X1 U22488 ( .A1(n19916), .A2(n19590), .B1(n9784), .B2(n19912), .ZN(
        n19570) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19568), .B1(
        n19914), .B2(n19567), .ZN(n19569) );
  OAI211_X1 U22490 ( .C1(n19922), .C2(n19571), .A(n19570), .B(n19569), .ZN(
        P2_U3095) );
  NAND2_X1 U22491 ( .A1(n10561), .A2(n19858), .ZN(n19603) );
  NOR2_X1 U22492 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19603), .ZN(
        n19595) );
  OR3_X1 U22493 ( .A1(n12145), .A2(n19595), .A3(n20035), .ZN(n19577) );
  NOR2_X1 U22494 ( .A1(n19576), .A2(n19595), .ZN(n19573) );
  OAI21_X1 U22495 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19573), .A(n20035), 
        .ZN(n19574) );
  AND2_X1 U22496 ( .A1(n19577), .A2(n19574), .ZN(n19596) );
  AOI22_X1 U22497 ( .A1(n19596), .A2(n19862), .B1(n19861), .B2(n19595), .ZN(
        n19581) );
  AOI21_X1 U22498 ( .B1(n19600), .B2(n19621), .A(n19695), .ZN(n19575) );
  AOI221_X1 U22499 ( .B1(n19632), .B2(n19576), .C1(n19632), .C2(n19575), .A(
        n19595), .ZN(n19579) );
  INV_X1 U22500 ( .A(n19577), .ZN(n19578) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19597), .B1(
        n19590), .B2(n19758), .ZN(n19580) );
  OAI211_X1 U22502 ( .C1(n19761), .C2(n19621), .A(n19581), .B(n19580), .ZN(
        P2_U3096) );
  AOI22_X1 U22503 ( .A1(n19596), .A2(n19875), .B1(n19874), .B2(n19595), .ZN(
        n19583) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19597), .B1(
        n19590), .B2(n19829), .ZN(n19582) );
  OAI211_X1 U22505 ( .C1(n19832), .C2(n19621), .A(n19583), .B(n19582), .ZN(
        P2_U3097) );
  AOI22_X1 U22506 ( .A1(n19596), .A2(n19881), .B1(n19880), .B2(n19595), .ZN(
        n19585) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19597), .B1(
        n19625), .B2(n19882), .ZN(n19584) );
  OAI211_X1 U22508 ( .C1(n19885), .C2(n19600), .A(n19585), .B(n19584), .ZN(
        P2_U3098) );
  AOI22_X1 U22509 ( .A1(n19596), .A2(n19887), .B1(n19886), .B2(n19595), .ZN(
        n19587) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19597), .B1(
        n19625), .B2(n19888), .ZN(n19586) );
  OAI211_X1 U22511 ( .C1(n19891), .C2(n19600), .A(n19587), .B(n19586), .ZN(
        P2_U3099) );
  AOI22_X1 U22512 ( .A1(n19596), .A2(n19893), .B1(n19892), .B2(n19595), .ZN(
        n19589) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19597), .B1(
        n19625), .B2(n19841), .ZN(n19588) );
  OAI211_X1 U22514 ( .C1(n19844), .C2(n19600), .A(n19589), .B(n19588), .ZN(
        P2_U3100) );
  AOI22_X1 U22515 ( .A1(n19596), .A2(n19899), .B1(n19898), .B2(n19595), .ZN(
        n19592) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19597), .B1(
        n19590), .B2(n19900), .ZN(n19591) );
  OAI211_X1 U22517 ( .C1(n19905), .C2(n19621), .A(n19592), .B(n19591), .ZN(
        P2_U3101) );
  AOI22_X1 U22518 ( .A1(n19596), .A2(n19907), .B1(n19906), .B2(n19595), .ZN(
        n19594) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19597), .B1(
        n19625), .B2(n19908), .ZN(n19593) );
  OAI211_X1 U22520 ( .C1(n19911), .C2(n19600), .A(n19594), .B(n19593), .ZN(
        P2_U3102) );
  AOI22_X1 U22521 ( .A1(n19596), .A2(n19914), .B1(n19912), .B2(n19595), .ZN(
        n19599) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19597), .B1(
        n19625), .B2(n19916), .ZN(n19598) );
  OAI211_X1 U22523 ( .C1(n19922), .C2(n19600), .A(n19599), .B(n19598), .ZN(
        P2_U3103) );
  NOR2_X1 U22524 ( .A1(n20042), .A2(n19603), .ZN(n19637) );
  INV_X1 U22525 ( .A(n19637), .ZN(n19634) );
  NAND2_X1 U22526 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19634), .ZN(n19601) );
  NOR2_X1 U22527 ( .A1(n12152), .A2(n19601), .ZN(n19605) );
  AOI211_X2 U22528 ( .C1(n19603), .C2(n20035), .A(n19602), .B(n19605), .ZN(
        n19624) );
  AOI22_X1 U22529 ( .A1(n19624), .A2(n19862), .B1(n19861), .B2(n19637), .ZN(
        n19610) );
  INV_X1 U22530 ( .A(n19603), .ZN(n19607) );
  INV_X1 U22531 ( .A(n19814), .ZN(n19863) );
  AND2_X1 U22532 ( .A1(n19604), .A2(n19863), .ZN(n20005) );
  AOI211_X1 U22533 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19634), .A(n19754), 
        .B(n19605), .ZN(n19606) );
  OAI21_X1 U22534 ( .B1(n19607), .B2(n20005), .A(n19606), .ZN(n19626) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19870), .ZN(n19609) );
  OAI211_X1 U22536 ( .C1(n19873), .C2(n19621), .A(n19610), .B(n19609), .ZN(
        P2_U3104) );
  AOI22_X1 U22537 ( .A1(n19624), .A2(n19875), .B1(n19874), .B2(n19637), .ZN(
        n19612) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19876), .ZN(n19611) );
  OAI211_X1 U22539 ( .C1(n19879), .C2(n19621), .A(n19612), .B(n19611), .ZN(
        P2_U3105) );
  AOI22_X1 U22540 ( .A1(n19624), .A2(n19881), .B1(n19880), .B2(n19637), .ZN(
        n19614) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19882), .ZN(n19613) );
  OAI211_X1 U22542 ( .C1(n19885), .C2(n19621), .A(n19614), .B(n19613), .ZN(
        P2_U3106) );
  AOI22_X1 U22543 ( .A1(n19624), .A2(n19887), .B1(n19886), .B2(n19637), .ZN(
        n19616) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19888), .ZN(n19615) );
  OAI211_X1 U22545 ( .C1(n19891), .C2(n19621), .A(n19616), .B(n19615), .ZN(
        P2_U3107) );
  AOI22_X1 U22546 ( .A1(n19624), .A2(n19893), .B1(n19892), .B2(n19637), .ZN(
        n19618) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19841), .ZN(n19617) );
  OAI211_X1 U22548 ( .C1(n19844), .C2(n19621), .A(n19618), .B(n19617), .ZN(
        P2_U3108) );
  AOI22_X1 U22549 ( .A1(n19624), .A2(n19899), .B1(n19898), .B2(n19637), .ZN(
        n19620) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19800), .ZN(n19619) );
  OAI211_X1 U22551 ( .C1(n19803), .C2(n19621), .A(n19620), .B(n19619), .ZN(
        P2_U3109) );
  AOI22_X1 U22552 ( .A1(n19624), .A2(n19907), .B1(n19906), .B2(n19637), .ZN(
        n19623) );
  AOI22_X1 U22553 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19626), .B1(
        n19625), .B2(n19804), .ZN(n19622) );
  OAI211_X1 U22554 ( .C1(n19808), .C2(n19660), .A(n19623), .B(n19622), .ZN(
        P2_U3110) );
  AOI22_X1 U22555 ( .A1(n19624), .A2(n19914), .B1(n19912), .B2(n19637), .ZN(
        n19628) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19626), .B1(
        n19625), .B2(n19852), .ZN(n19627) );
  OAI211_X1 U22557 ( .C1(n19857), .C2(n19660), .A(n19628), .B(n19627), .ZN(
        P2_U3111) );
  NAND2_X1 U22558 ( .A1(n20023), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19726) );
  NOR2_X1 U22559 ( .A1(n19726), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19666) );
  INV_X1 U22560 ( .A(n19666), .ZN(n19668) );
  NOR2_X1 U22561 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19668), .ZN(
        n19655) );
  AOI22_X1 U22562 ( .A1(n19758), .A2(n19650), .B1(n19861), .B2(n19655), .ZN(
        n19641) );
  AOI21_X1 U22563 ( .B1(n19660), .B2(n19684), .A(n19695), .ZN(n19631) );
  NOR2_X1 U22564 ( .A1(n19631), .A2(n19819), .ZN(n19636) );
  OAI21_X1 U22565 ( .B1(n9668), .B2(n20035), .A(n19632), .ZN(n19633) );
  AOI21_X1 U22566 ( .B1(n19636), .B2(n19634), .A(n19633), .ZN(n19635) );
  OAI21_X1 U22567 ( .B1(n19655), .B2(n19637), .A(n19636), .ZN(n19639) );
  OAI21_X1 U22568 ( .B1(n9668), .B2(n19655), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19638) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19657), .B1(
        n19862), .B2(n19656), .ZN(n19640) );
  OAI211_X1 U22570 ( .C1(n19761), .C2(n19684), .A(n19641), .B(n19640), .ZN(
        P2_U3112) );
  AOI22_X1 U22571 ( .A1(n19829), .A2(n19650), .B1(n19874), .B2(n19655), .ZN(
        n19643) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19875), .ZN(n19642) );
  OAI211_X1 U22573 ( .C1(n19832), .C2(n19684), .A(n19643), .B(n19642), .ZN(
        P2_U3113) );
  AOI22_X1 U22574 ( .A1(n19833), .A2(n19650), .B1(n19880), .B2(n19655), .ZN(
        n19645) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19881), .ZN(n19644) );
  OAI211_X1 U22576 ( .C1(n19836), .C2(n19684), .A(n19645), .B(n19644), .ZN(
        P2_U3114) );
  AOI22_X1 U22577 ( .A1(n19837), .A2(n19650), .B1(n19886), .B2(n19655), .ZN(
        n19647) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19887), .ZN(n19646) );
  OAI211_X1 U22579 ( .C1(n19840), .C2(n19684), .A(n19647), .B(n19646), .ZN(
        P2_U3115) );
  AOI22_X1 U22580 ( .A1(n19841), .A2(n19685), .B1(n19892), .B2(n19655), .ZN(
        n19649) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19893), .ZN(n19648) );
  OAI211_X1 U22582 ( .C1(n19844), .C2(n19660), .A(n19649), .B(n19648), .ZN(
        P2_U3116) );
  AOI22_X1 U22583 ( .A1(n19900), .A2(n19650), .B1(n19898), .B2(n19655), .ZN(
        n19652) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19899), .ZN(n19651) );
  OAI211_X1 U22585 ( .C1(n19905), .C2(n19684), .A(n19652), .B(n19651), .ZN(
        P2_U3117) );
  AOI22_X1 U22586 ( .A1(n19908), .A2(n19685), .B1(n19906), .B2(n19655), .ZN(
        n19654) );
  AOI22_X1 U22587 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19907), .ZN(n19653) );
  OAI211_X1 U22588 ( .C1(n19911), .C2(n19660), .A(n19654), .B(n19653), .ZN(
        P2_U3118) );
  AOI22_X1 U22589 ( .A1(n19916), .A2(n19685), .B1(n19912), .B2(n19655), .ZN(
        n19659) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19914), .ZN(n19658) );
  OAI211_X1 U22591 ( .C1(n19922), .C2(n19660), .A(n19659), .B(n19658), .ZN(
        P2_U3119) );
  NOR2_X1 U22592 ( .A1(n19661), .A2(n19726), .ZN(n19697) );
  AOI22_X1 U22593 ( .A1(n19758), .A2(n19685), .B1(n19861), .B2(n19697), .ZN(
        n19671) );
  NAND2_X1 U22594 ( .A1(n20010), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19782) );
  OAI21_X1 U22595 ( .B1(n19782), .B2(n19662), .A(n20006), .ZN(n19669) );
  OAI21_X1 U22596 ( .B1(n12151), .B2(n20035), .A(n19632), .ZN(n19664) );
  INV_X1 U22597 ( .A(n19697), .ZN(n19663) );
  AOI21_X1 U22598 ( .B1(n19664), .B2(n19663), .A(n19754), .ZN(n19665) );
  OAI21_X1 U22599 ( .B1(n19669), .B2(n19666), .A(n19665), .ZN(n19687) );
  OAI21_X1 U22600 ( .B1(n12151), .B2(n19697), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19667) );
  OAI21_X1 U22601 ( .B1(n19669), .B2(n19668), .A(n19667), .ZN(n19686) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19687), .B1(
        n19862), .B2(n19686), .ZN(n19670) );
  OAI211_X1 U22603 ( .C1(n19761), .C2(n19696), .A(n19671), .B(n19670), .ZN(
        P2_U3120) );
  AOI22_X1 U22604 ( .A1(n19876), .A2(n19718), .B1(n19874), .B2(n19697), .ZN(
        n19673) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19687), .B1(
        n19875), .B2(n19686), .ZN(n19672) );
  OAI211_X1 U22606 ( .C1(n19879), .C2(n19684), .A(n19673), .B(n19672), .ZN(
        P2_U3121) );
  AOI22_X1 U22607 ( .A1(n19882), .A2(n19718), .B1(n19880), .B2(n19697), .ZN(
        n19675) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19687), .B1(
        n19881), .B2(n19686), .ZN(n19674) );
  OAI211_X1 U22609 ( .C1(n19885), .C2(n19684), .A(n19675), .B(n19674), .ZN(
        P2_U3122) );
  AOI22_X1 U22610 ( .A1(n19888), .A2(n19718), .B1(n19886), .B2(n19697), .ZN(
        n19677) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19687), .B1(
        n19887), .B2(n19686), .ZN(n19676) );
  OAI211_X1 U22612 ( .C1(n19891), .C2(n19684), .A(n19677), .B(n19676), .ZN(
        P2_U3123) );
  AOI22_X1 U22613 ( .A1(n19841), .A2(n19718), .B1(n19892), .B2(n19697), .ZN(
        n19679) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19687), .B1(
        n19893), .B2(n19686), .ZN(n19678) );
  OAI211_X1 U22615 ( .C1(n19844), .C2(n19684), .A(n19679), .B(n19678), .ZN(
        P2_U3124) );
  AOI22_X1 U22616 ( .A1(n19900), .A2(n19685), .B1(n19898), .B2(n19697), .ZN(
        n19681) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19687), .B1(
        n19899), .B2(n19686), .ZN(n19680) );
  OAI211_X1 U22618 ( .C1(n19905), .C2(n19696), .A(n19681), .B(n19680), .ZN(
        P2_U3125) );
  AOI22_X1 U22619 ( .A1(n19908), .A2(n19718), .B1(n19906), .B2(n19697), .ZN(
        n19683) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19687), .B1(
        n19907), .B2(n19686), .ZN(n19682) );
  OAI211_X1 U22621 ( .C1(n19911), .C2(n19684), .A(n19683), .B(n19682), .ZN(
        P2_U3126) );
  AOI22_X1 U22622 ( .A1(n19852), .A2(n19685), .B1(n19912), .B2(n19697), .ZN(
        n19689) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19687), .B1(
        n19914), .B2(n19686), .ZN(n19688) );
  OAI211_X1 U22624 ( .C1(n19857), .C2(n19696), .A(n19689), .B(n19688), .ZN(
        P2_U3127) );
  INV_X1 U22625 ( .A(n19690), .ZN(n19694) );
  INV_X1 U22626 ( .A(n19726), .ZN(n19723) );
  AND2_X1 U22627 ( .A1(n19691), .A2(n19723), .ZN(n19716) );
  OAI21_X1 U22628 ( .B1(n19692), .B2(n19716), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19693) );
  OAI21_X1 U22629 ( .B1(n19726), .B2(n19694), .A(n19693), .ZN(n19717) );
  AOI22_X1 U22630 ( .A1(n19717), .A2(n19862), .B1(n19861), .B2(n19716), .ZN(
        n19703) );
  AOI21_X1 U22631 ( .B1(n19749), .B2(n19696), .A(n19695), .ZN(n19698) );
  NOR2_X1 U22632 ( .A1(n19698), .A2(n19697), .ZN(n19699) );
  AOI211_X1 U22633 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19700), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19699), .ZN(n19701) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19719), .B1(
        n19718), .B2(n19758), .ZN(n19702) );
  OAI211_X1 U22635 ( .C1(n19761), .C2(n19749), .A(n19703), .B(n19702), .ZN(
        P2_U3128) );
  AOI22_X1 U22636 ( .A1(n19717), .A2(n19875), .B1(n19874), .B2(n19716), .ZN(
        n19705) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19719), .B1(
        n19718), .B2(n19829), .ZN(n19704) );
  OAI211_X1 U22638 ( .C1(n19832), .C2(n19749), .A(n19705), .B(n19704), .ZN(
        P2_U3129) );
  AOI22_X1 U22639 ( .A1(n19717), .A2(n19881), .B1(n19880), .B2(n19716), .ZN(
        n19707) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19719), .B1(
        n19718), .B2(n19833), .ZN(n19706) );
  OAI211_X1 U22641 ( .C1(n19836), .C2(n19749), .A(n19707), .B(n19706), .ZN(
        P2_U3130) );
  AOI22_X1 U22642 ( .A1(n19717), .A2(n19887), .B1(n19886), .B2(n19716), .ZN(
        n19709) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19719), .B1(
        n19718), .B2(n19837), .ZN(n19708) );
  OAI211_X1 U22644 ( .C1(n19840), .C2(n19749), .A(n19709), .B(n19708), .ZN(
        P2_U3131) );
  AOI22_X1 U22645 ( .A1(n19717), .A2(n19893), .B1(n19892), .B2(n19716), .ZN(
        n19711) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19719), .B1(
        n19718), .B2(n19894), .ZN(n19710) );
  OAI211_X1 U22647 ( .C1(n19897), .C2(n19749), .A(n19711), .B(n19710), .ZN(
        P2_U3132) );
  AOI22_X1 U22648 ( .A1(n19717), .A2(n19899), .B1(n19898), .B2(n19716), .ZN(
        n19713) );
  AOI22_X1 U22649 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19719), .B1(
        n19718), .B2(n19900), .ZN(n19712) );
  OAI211_X1 U22650 ( .C1(n19905), .C2(n19749), .A(n19713), .B(n19712), .ZN(
        P2_U3133) );
  AOI22_X1 U22651 ( .A1(n19717), .A2(n19907), .B1(n19906), .B2(n19716), .ZN(
        n19715) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19719), .B1(
        n19718), .B2(n19804), .ZN(n19714) );
  OAI211_X1 U22653 ( .C1(n19808), .C2(n19749), .A(n19715), .B(n19714), .ZN(
        P2_U3134) );
  AOI22_X1 U22654 ( .A1(n19717), .A2(n19914), .B1(n19912), .B2(n19716), .ZN(
        n19721) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19719), .B1(
        n19718), .B2(n19852), .ZN(n19720) );
  OAI211_X1 U22656 ( .C1(n19857), .C2(n19749), .A(n19721), .B(n19720), .ZN(
        P2_U3135) );
  NOR2_X1 U22657 ( .A1(n19722), .A2(n19726), .ZN(n19744) );
  NAND2_X1 U22658 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19723), .ZN(
        n19724) );
  OAI21_X1 U22659 ( .B1(n19724), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20035), 
        .ZN(n19725) );
  AOI22_X1 U22660 ( .A1(n19745), .A2(n19862), .B1(n19861), .B2(n19744), .ZN(
        n19731) );
  NOR3_X1 U22661 ( .A1(n19782), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n20007), 
        .ZN(n19729) );
  AOI211_X1 U22662 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20042), .A(n20033), 
        .B(n19726), .ZN(n19728) );
  OAI211_X1 U22663 ( .C1(n19729), .C2(n19728), .A(n19868), .B(n19727), .ZN(
        n19746) );
  NOR2_X2 U22664 ( .A1(n19789), .A2(n20007), .ZN(n19776) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19746), .B1(
        n19776), .B2(n19870), .ZN(n19730) );
  OAI211_X1 U22666 ( .C1(n19873), .C2(n19749), .A(n19731), .B(n19730), .ZN(
        P2_U3136) );
  AOI22_X1 U22667 ( .A1(n19745), .A2(n19875), .B1(n19874), .B2(n19744), .ZN(
        n19733) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19746), .B1(
        n19776), .B2(n19876), .ZN(n19732) );
  OAI211_X1 U22669 ( .C1(n19879), .C2(n19749), .A(n19733), .B(n19732), .ZN(
        P2_U3137) );
  AOI22_X1 U22670 ( .A1(n19745), .A2(n19881), .B1(n19880), .B2(n19744), .ZN(
        n19735) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19746), .B1(
        n19776), .B2(n19882), .ZN(n19734) );
  OAI211_X1 U22672 ( .C1(n19885), .C2(n19749), .A(n19735), .B(n19734), .ZN(
        P2_U3138) );
  AOI22_X1 U22673 ( .A1(n19745), .A2(n19887), .B1(n19886), .B2(n19744), .ZN(
        n19737) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19746), .B1(
        n19776), .B2(n19888), .ZN(n19736) );
  OAI211_X1 U22675 ( .C1(n19891), .C2(n19749), .A(n19737), .B(n19736), .ZN(
        P2_U3139) );
  AOI22_X1 U22676 ( .A1(n19745), .A2(n19893), .B1(n19892), .B2(n19744), .ZN(
        n19739) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19746), .B1(
        n19776), .B2(n19841), .ZN(n19738) );
  OAI211_X1 U22678 ( .C1(n19844), .C2(n19749), .A(n19739), .B(n19738), .ZN(
        P2_U3140) );
  AOI22_X1 U22679 ( .A1(n19745), .A2(n19899), .B1(n19898), .B2(n19744), .ZN(
        n19741) );
  AOI22_X1 U22680 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19746), .B1(
        n19776), .B2(n19800), .ZN(n19740) );
  OAI211_X1 U22681 ( .C1(n19803), .C2(n19749), .A(n19741), .B(n19740), .ZN(
        P2_U3141) );
  AOI22_X1 U22682 ( .A1(n19745), .A2(n19907), .B1(n19906), .B2(n19744), .ZN(
        n19743) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19746), .B1(
        n19776), .B2(n19908), .ZN(n19742) );
  OAI211_X1 U22684 ( .C1(n19911), .C2(n19749), .A(n19743), .B(n19742), .ZN(
        P2_U3142) );
  AOI22_X1 U22685 ( .A1(n19745), .A2(n19914), .B1(n19912), .B2(n19744), .ZN(
        n19748) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19746), .B1(
        n19776), .B2(n19916), .ZN(n19747) );
  OAI211_X1 U22687 ( .C1(n19922), .C2(n19749), .A(n19748), .B(n19747), .ZN(
        P2_U3143) );
  NAND3_X1 U22688 ( .A1(n20033), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19785) );
  NOR2_X1 U22689 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19785), .ZN(
        n19774) );
  NOR3_X1 U22690 ( .A1(n12102), .A2(n19774), .A3(n20035), .ZN(n19753) );
  NAND2_X1 U22691 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19750), .ZN(
        n19755) );
  INV_X1 U22692 ( .A(n19755), .ZN(n19751) );
  AOI21_X1 U22693 ( .B1(n19751), .B2(n19632), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19752) );
  AOI22_X1 U22694 ( .A1(n19775), .A2(n19862), .B1(n19861), .B2(n19774), .ZN(
        n19760) );
  OAI21_X1 U22695 ( .B1(n19805), .B2(n19776), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19756) );
  AOI211_X1 U22696 ( .C1(n19756), .C2(n19755), .A(n19754), .B(n19753), .ZN(
        n19757) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19758), .ZN(n19759) );
  OAI211_X1 U22698 ( .C1(n19761), .C2(n19813), .A(n19760), .B(n19759), .ZN(
        P2_U3144) );
  AOI22_X1 U22699 ( .A1(n19775), .A2(n19875), .B1(n19874), .B2(n19774), .ZN(
        n19763) );
  AOI22_X1 U22700 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19829), .ZN(n19762) );
  OAI211_X1 U22701 ( .C1(n19832), .C2(n19813), .A(n19763), .B(n19762), .ZN(
        P2_U3145) );
  AOI22_X1 U22702 ( .A1(n19775), .A2(n19881), .B1(n19880), .B2(n19774), .ZN(
        n19765) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19833), .ZN(n19764) );
  OAI211_X1 U22704 ( .C1(n19836), .C2(n19813), .A(n19765), .B(n19764), .ZN(
        P2_U3146) );
  AOI22_X1 U22705 ( .A1(n19775), .A2(n19887), .B1(n19886), .B2(n19774), .ZN(
        n19767) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19837), .ZN(n19766) );
  OAI211_X1 U22707 ( .C1(n19840), .C2(n19813), .A(n19767), .B(n19766), .ZN(
        P2_U3147) );
  AOI22_X1 U22708 ( .A1(n19775), .A2(n19893), .B1(n19892), .B2(n19774), .ZN(
        n19769) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19894), .ZN(n19768) );
  OAI211_X1 U22710 ( .C1(n19897), .C2(n19813), .A(n19769), .B(n19768), .ZN(
        P2_U3148) );
  AOI22_X1 U22711 ( .A1(n19775), .A2(n19899), .B1(n19898), .B2(n19774), .ZN(
        n19771) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19900), .ZN(n19770) );
  OAI211_X1 U22713 ( .C1(n19905), .C2(n19813), .A(n19771), .B(n19770), .ZN(
        P2_U3149) );
  AOI22_X1 U22714 ( .A1(n19775), .A2(n19907), .B1(n19906), .B2(n19774), .ZN(
        n19773) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19804), .ZN(n19772) );
  OAI211_X1 U22716 ( .C1(n19808), .C2(n19813), .A(n19773), .B(n19772), .ZN(
        P2_U3150) );
  AOI22_X1 U22717 ( .A1(n19775), .A2(n19914), .B1(n19912), .B2(n19774), .ZN(
        n19779) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19852), .ZN(n19778) );
  OAI211_X1 U22719 ( .C1(n19857), .C2(n19813), .A(n19779), .B(n19778), .ZN(
        P2_U3151) );
  NOR2_X1 U22720 ( .A1(n20042), .A2(n19785), .ZN(n19818) );
  NOR3_X1 U22721 ( .A1(n12141), .A2(n19818), .A3(n20035), .ZN(n19784) );
  INV_X1 U22722 ( .A(n19785), .ZN(n19780) );
  AOI21_X1 U22723 ( .B1(n19632), .B2(n19780), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19781) );
  NOR2_X1 U22724 ( .A1(n19784), .A2(n19781), .ZN(n19809) );
  AOI22_X1 U22725 ( .A1(n19809), .A2(n19862), .B1(n19861), .B2(n19818), .ZN(
        n19791) );
  INV_X1 U22726 ( .A(n19782), .ZN(n19864) );
  INV_X1 U22727 ( .A(n19788), .ZN(n19783) );
  NAND2_X1 U22728 ( .A1(n19864), .A2(n19783), .ZN(n19786) );
  AOI21_X1 U22729 ( .B1(n19786), .B2(n19785), .A(n19784), .ZN(n19787) );
  OAI211_X1 U22730 ( .C1(n19818), .C2(n19632), .A(n19787), .B(n19868), .ZN(
        n19810) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19810), .B1(
        n19851), .B2(n19870), .ZN(n19790) );
  OAI211_X1 U22732 ( .C1(n19873), .C2(n19813), .A(n19791), .B(n19790), .ZN(
        P2_U3152) );
  AOI22_X1 U22733 ( .A1(n19809), .A2(n19875), .B1(n19874), .B2(n19818), .ZN(
        n19793) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19810), .B1(
        n19851), .B2(n19876), .ZN(n19792) );
  OAI211_X1 U22735 ( .C1(n19879), .C2(n19813), .A(n19793), .B(n19792), .ZN(
        P2_U3153) );
  AOI22_X1 U22736 ( .A1(n19809), .A2(n19881), .B1(n19880), .B2(n19818), .ZN(
        n19795) );
  AOI22_X1 U22737 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19810), .B1(
        n19851), .B2(n19882), .ZN(n19794) );
  OAI211_X1 U22738 ( .C1(n19885), .C2(n19813), .A(n19795), .B(n19794), .ZN(
        P2_U3154) );
  AOI22_X1 U22739 ( .A1(n19809), .A2(n19887), .B1(n19886), .B2(n19818), .ZN(
        n19797) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19810), .B1(
        n19805), .B2(n19837), .ZN(n19796) );
  OAI211_X1 U22741 ( .C1(n19840), .C2(n19849), .A(n19797), .B(n19796), .ZN(
        P2_U3155) );
  AOI22_X1 U22742 ( .A1(n19809), .A2(n19893), .B1(n19892), .B2(n19818), .ZN(
        n19799) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19810), .B1(
        n19805), .B2(n19894), .ZN(n19798) );
  OAI211_X1 U22744 ( .C1(n19897), .C2(n19849), .A(n19799), .B(n19798), .ZN(
        P2_U3156) );
  AOI22_X1 U22745 ( .A1(n19809), .A2(n19899), .B1(n19898), .B2(n19818), .ZN(
        n19802) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19810), .B1(
        n19851), .B2(n19800), .ZN(n19801) );
  OAI211_X1 U22747 ( .C1(n19803), .C2(n19813), .A(n19802), .B(n19801), .ZN(
        P2_U3157) );
  AOI22_X1 U22748 ( .A1(n19809), .A2(n19907), .B1(n19906), .B2(n19818), .ZN(
        n19807) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19810), .B1(
        n19805), .B2(n19804), .ZN(n19806) );
  OAI211_X1 U22750 ( .C1(n19808), .C2(n19849), .A(n19807), .B(n19806), .ZN(
        P2_U3158) );
  AOI22_X1 U22751 ( .A1(n19809), .A2(n19914), .B1(n19912), .B2(n19818), .ZN(
        n19812) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19810), .B1(
        n19851), .B2(n19916), .ZN(n19811) );
  OAI211_X1 U22753 ( .C1(n19922), .C2(n19813), .A(n19812), .B(n19811), .ZN(
        P2_U3159) );
  INV_X1 U22754 ( .A(n19858), .ZN(n19816) );
  NOR3_X2 U22755 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10561), .A3(
        n19816), .ZN(n19850) );
  AOI22_X1 U22756 ( .A1(n19870), .A2(n19901), .B1(n19861), .B2(n19850), .ZN(
        n19828) );
  OAI21_X1 U22757 ( .B1(n19901), .B2(n19851), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19817) );
  NAND2_X1 U22758 ( .A1(n19817), .A2(n20006), .ZN(n19826) );
  NOR2_X1 U22759 ( .A1(n19850), .A2(n19818), .ZN(n19825) );
  INV_X1 U22760 ( .A(n19825), .ZN(n19823) );
  INV_X1 U22761 ( .A(n12153), .ZN(n19821) );
  INV_X1 U22762 ( .A(n19850), .ZN(n19820) );
  OAI211_X1 U22763 ( .C1(n19821), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19820), 
        .B(n19819), .ZN(n19822) );
  OAI211_X1 U22764 ( .C1(n19826), .C2(n19823), .A(n19868), .B(n19822), .ZN(
        n19854) );
  OAI21_X1 U22765 ( .B1(n12153), .B2(n19850), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19824) );
  AOI22_X1 U22766 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19854), .B1(
        n19862), .B2(n19853), .ZN(n19827) );
  OAI211_X1 U22767 ( .C1(n19873), .C2(n19849), .A(n19828), .B(n19827), .ZN(
        P2_U3160) );
  AOI22_X1 U22768 ( .A1(n19829), .A2(n19851), .B1(n19874), .B2(n19850), .ZN(
        n19831) );
  AOI22_X1 U22769 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19854), .B1(
        n19875), .B2(n19853), .ZN(n19830) );
  OAI211_X1 U22770 ( .C1(n19832), .C2(n19921), .A(n19831), .B(n19830), .ZN(
        P2_U3161) );
  AOI22_X1 U22771 ( .A1(n19833), .A2(n19851), .B1(n19880), .B2(n19850), .ZN(
        n19835) );
  AOI22_X1 U22772 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19854), .B1(
        n19881), .B2(n19853), .ZN(n19834) );
  OAI211_X1 U22773 ( .C1(n19836), .C2(n19921), .A(n19835), .B(n19834), .ZN(
        P2_U3162) );
  AOI22_X1 U22774 ( .A1(n19837), .A2(n19851), .B1(n19886), .B2(n19850), .ZN(
        n19839) );
  AOI22_X1 U22775 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19854), .B1(
        n19887), .B2(n19853), .ZN(n19838) );
  OAI211_X1 U22776 ( .C1(n19840), .C2(n19921), .A(n19839), .B(n19838), .ZN(
        P2_U3163) );
  AOI22_X1 U22777 ( .A1(n19841), .A2(n19901), .B1(n19892), .B2(n19850), .ZN(
        n19843) );
  AOI22_X1 U22778 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19854), .B1(
        n19893), .B2(n19853), .ZN(n19842) );
  OAI211_X1 U22779 ( .C1(n19844), .C2(n19849), .A(n19843), .B(n19842), .ZN(
        P2_U3164) );
  AOI22_X1 U22780 ( .A1(n19900), .A2(n19851), .B1(n19898), .B2(n19850), .ZN(
        n19846) );
  AOI22_X1 U22781 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19854), .B1(
        n19899), .B2(n19853), .ZN(n19845) );
  OAI211_X1 U22782 ( .C1(n19905), .C2(n19921), .A(n19846), .B(n19845), .ZN(
        P2_U3165) );
  AOI22_X1 U22783 ( .A1(n19908), .A2(n19901), .B1(n19906), .B2(n19850), .ZN(
        n19848) );
  AOI22_X1 U22784 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19854), .B1(
        n19907), .B2(n19853), .ZN(n19847) );
  OAI211_X1 U22785 ( .C1(n19911), .C2(n19849), .A(n19848), .B(n19847), .ZN(
        P2_U3166) );
  AOI22_X1 U22786 ( .A1(n19852), .A2(n19851), .B1(n19912), .B2(n19850), .ZN(
        n19856) );
  AOI22_X1 U22787 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19854), .B1(
        n19914), .B2(n19853), .ZN(n19855) );
  OAI211_X1 U22788 ( .C1(n19857), .C2(n19921), .A(n19856), .B(n19855), .ZN(
        P2_U3167) );
  NAND2_X1 U22789 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19858), .ZN(
        n19866) );
  OR2_X1 U22790 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19866), .ZN(n19860) );
  NOR3_X1 U22791 ( .A1(n19859), .A2(n19913), .A3(n20035), .ZN(n19865) );
  AOI21_X1 U22792 ( .B1(n20035), .B2(n19860), .A(n19865), .ZN(n19915) );
  AOI22_X1 U22793 ( .A1(n19915), .A2(n19862), .B1(n19913), .B2(n19861), .ZN(
        n19872) );
  NAND2_X1 U22794 ( .A1(n19864), .A2(n19863), .ZN(n19867) );
  AOI21_X1 U22795 ( .B1(n19867), .B2(n19866), .A(n19865), .ZN(n19869) );
  OAI211_X1 U22796 ( .C1(n19913), .C2(n19632), .A(n19869), .B(n19868), .ZN(
        n19918) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19918), .B1(
        n19917), .B2(n19870), .ZN(n19871) );
  OAI211_X1 U22798 ( .C1(n19873), .C2(n19921), .A(n19872), .B(n19871), .ZN(
        P2_U3168) );
  AOI22_X1 U22799 ( .A1(n19915), .A2(n19875), .B1(n19913), .B2(n19874), .ZN(
        n19878) );
  AOI22_X1 U22800 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19918), .B1(
        n19917), .B2(n19876), .ZN(n19877) );
  OAI211_X1 U22801 ( .C1(n19879), .C2(n19921), .A(n19878), .B(n19877), .ZN(
        P2_U3169) );
  AOI22_X1 U22802 ( .A1(n19915), .A2(n19881), .B1(n19913), .B2(n19880), .ZN(
        n19884) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19918), .B1(
        n19917), .B2(n19882), .ZN(n19883) );
  OAI211_X1 U22804 ( .C1(n19885), .C2(n19921), .A(n19884), .B(n19883), .ZN(
        P2_U3170) );
  AOI22_X1 U22805 ( .A1(n19915), .A2(n19887), .B1(n19913), .B2(n19886), .ZN(
        n19890) );
  AOI22_X1 U22806 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19918), .B1(
        n19917), .B2(n19888), .ZN(n19889) );
  OAI211_X1 U22807 ( .C1(n19891), .C2(n19921), .A(n19890), .B(n19889), .ZN(
        P2_U3171) );
  INV_X1 U22808 ( .A(n19917), .ZN(n19904) );
  AOI22_X1 U22809 ( .A1(n19915), .A2(n19893), .B1(n19913), .B2(n19892), .ZN(
        n19896) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19918), .B1(
        n19901), .B2(n19894), .ZN(n19895) );
  OAI211_X1 U22811 ( .C1(n19897), .C2(n19904), .A(n19896), .B(n19895), .ZN(
        P2_U3172) );
  AOI22_X1 U22812 ( .A1(n19915), .A2(n19899), .B1(n19913), .B2(n19898), .ZN(
        n19903) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19918), .B1(
        n19901), .B2(n19900), .ZN(n19902) );
  OAI211_X1 U22814 ( .C1(n19905), .C2(n19904), .A(n19903), .B(n19902), .ZN(
        P2_U3173) );
  AOI22_X1 U22815 ( .A1(n19915), .A2(n19907), .B1(n19913), .B2(n19906), .ZN(
        n19910) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19918), .B1(
        n19917), .B2(n19908), .ZN(n19909) );
  OAI211_X1 U22817 ( .C1(n19911), .C2(n19921), .A(n19910), .B(n19909), .ZN(
        P2_U3174) );
  AOI22_X1 U22818 ( .A1(n19915), .A2(n19914), .B1(n19913), .B2(n19912), .ZN(
        n19920) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19918), .B1(
        n19917), .B2(n19916), .ZN(n19919) );
  OAI211_X1 U22820 ( .C1(n19922), .C2(n19921), .A(n19920), .B(n19919), .ZN(
        P2_U3175) );
  OAI211_X1 U22821 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19924), .A(n19925), 
        .B(n19923), .ZN(n19931) );
  INV_X1 U22822 ( .A(n19925), .ZN(n19928) );
  NOR2_X1 U22823 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19926), .ZN(n19927) );
  OAI211_X1 U22824 ( .C1(n19928), .C2(n19927), .A(n19943), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19930) );
  OAI211_X1 U22825 ( .C1(n19932), .C2(n19931), .A(n19930), .B(n19929), .ZN(
        P2_U3177) );
  INV_X1 U22826 ( .A(n20004), .ZN(n19934) );
  AND2_X1 U22827 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19934), .ZN(
        P2_U3179) );
  AND2_X1 U22828 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19934), .ZN(
        P2_U3180) );
  AND2_X1 U22829 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19934), .ZN(
        P2_U3181) );
  AND2_X1 U22830 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19934), .ZN(
        P2_U3182) );
  AND2_X1 U22831 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19934), .ZN(
        P2_U3183) );
  AND2_X1 U22832 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19934), .ZN(
        P2_U3184) );
  AND2_X1 U22833 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19934), .ZN(
        P2_U3185) );
  AND2_X1 U22834 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19934), .ZN(
        P2_U3186) );
  AND2_X1 U22835 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19934), .ZN(
        P2_U3187) );
  AND2_X1 U22836 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19934), .ZN(
        P2_U3188) );
  AND2_X1 U22837 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19934), .ZN(
        P2_U3189) );
  NOR2_X1 U22838 ( .A1(n19933), .A2(n20004), .ZN(P2_U3190) );
  AND2_X1 U22839 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19934), .ZN(
        P2_U3191) );
  AND2_X1 U22840 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19934), .ZN(
        P2_U3192) );
  AND2_X1 U22841 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19934), .ZN(
        P2_U3193) );
  AND2_X1 U22842 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19934), .ZN(
        P2_U3194) );
  AND2_X1 U22843 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19934), .ZN(
        P2_U3195) );
  AND2_X1 U22844 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19934), .ZN(
        P2_U3196) );
  AND2_X1 U22845 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19934), .ZN(
        P2_U3197) );
  AND2_X1 U22846 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19934), .ZN(
        P2_U3198) );
  AND2_X1 U22847 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19934), .ZN(
        P2_U3199) );
  AND2_X1 U22848 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19934), .ZN(
        P2_U3200) );
  AND2_X1 U22849 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19934), .ZN(P2_U3201) );
  AND2_X1 U22850 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19934), .ZN(P2_U3202) );
  NOR2_X1 U22851 ( .A1(n20975), .A2(n20004), .ZN(P2_U3203) );
  AND2_X1 U22852 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19934), .ZN(P2_U3204) );
  AND2_X1 U22853 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19934), .ZN(P2_U3205) );
  AND2_X1 U22854 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19934), .ZN(P2_U3206) );
  AND2_X1 U22855 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19934), .ZN(P2_U3207) );
  AND2_X1 U22856 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19934), .ZN(P2_U3208) );
  NAND2_X1 U22857 ( .A1(n19943), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19945) );
  NAND3_X1 U22858 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19945), .ZN(n19935) );
  NOR3_X1 U22859 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20883), .ZN(n19950) );
  AOI21_X1 U22860 ( .B1(n19951), .B2(n19935), .A(n19950), .ZN(n19936) );
  OAI221_X1 U22861 ( .B1(n19937), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n19937), .C2(n20873), .A(n19936), .ZN(P2_U3209) );
  AOI21_X1 U22862 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20873), .A(n19951), 
        .ZN(n19942) );
  NOR2_X1 U22863 ( .A1(n18953), .A2(n19942), .ZN(n19939) );
  AOI21_X1 U22864 ( .B1(n19939), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .A(n19938), .ZN(n19940) );
  OAI211_X1 U22865 ( .C1(n20873), .C2(n19941), .A(n19940), .B(n19945), .ZN(
        P2_U3210) );
  AND2_X1 U22866 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19944) );
  AOI21_X1 U22867 ( .B1(n19944), .B2(n19943), .A(n19942), .ZN(n19949) );
  OAI22_X1 U22868 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19946), .B1(NA), 
        .B2(n19945), .ZN(n19947) );
  OAI211_X1 U22869 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19947), .ZN(n19948) );
  OAI21_X1 U22870 ( .B1(n19950), .B2(n19949), .A(n19948), .ZN(P2_U3211) );
  OAI222_X1 U22871 ( .A1(n19997), .A2(n10458), .B1(n19952), .B2(n19995), .C1(
        n10428), .C2(n19994), .ZN(P2_U3212) );
  OAI222_X1 U22872 ( .A1(n19997), .A2(n10658), .B1(n19953), .B2(n19995), .C1(
        n10458), .C2(n19994), .ZN(P2_U3213) );
  OAI222_X1 U22873 ( .A1(n19997), .A2(n10674), .B1(n19954), .B2(n19995), .C1(
        n10658), .C2(n19994), .ZN(P2_U3214) );
  OAI222_X1 U22874 ( .A1(n19997), .A2(n13659), .B1(n19955), .B2(n19995), .C1(
        n10674), .C2(n19994), .ZN(P2_U3215) );
  OAI222_X1 U22875 ( .A1(n19997), .A2(n10493), .B1(n19956), .B2(n19995), .C1(
        n13659), .C2(n19994), .ZN(P2_U3216) );
  OAI222_X1 U22876 ( .A1(n19997), .A2(n20984), .B1(n19957), .B2(n19995), .C1(
        n10493), .C2(n19994), .ZN(P2_U3217) );
  OAI222_X1 U22877 ( .A1(n19997), .A2(n13561), .B1(n19958), .B2(n19995), .C1(
        n20984), .C2(n19994), .ZN(P2_U3218) );
  OAI222_X1 U22878 ( .A1(n19997), .A2(n10748), .B1(n19959), .B2(n19995), .C1(
        n13561), .C2(n19994), .ZN(P2_U3219) );
  OAI222_X1 U22879 ( .A1(n19997), .A2(n19961), .B1(n19960), .B2(n19995), .C1(
        n10748), .C2(n19994), .ZN(P2_U3220) );
  OAI222_X1 U22880 ( .A1(n19997), .A2(n15278), .B1(n19962), .B2(n19995), .C1(
        n19961), .C2(n19994), .ZN(P2_U3221) );
  OAI222_X1 U22881 ( .A1(n19997), .A2(n19964), .B1(n19963), .B2(n19995), .C1(
        n15278), .C2(n19994), .ZN(P2_U3222) );
  OAI222_X1 U22882 ( .A1(n19997), .A2(n19966), .B1(n19965), .B2(n19995), .C1(
        n19964), .C2(n19994), .ZN(P2_U3223) );
  OAI222_X1 U22883 ( .A1(n19997), .A2(n10814), .B1(n19967), .B2(n19995), .C1(
        n19966), .C2(n19994), .ZN(P2_U3224) );
  OAI222_X1 U22884 ( .A1(n19997), .A2(n21116), .B1(n19968), .B2(n19995), .C1(
        n10814), .C2(n19994), .ZN(P2_U3225) );
  OAI222_X1 U22885 ( .A1(n19997), .A2(n19970), .B1(n19969), .B2(n19995), .C1(
        n21116), .C2(n19994), .ZN(P2_U3226) );
  OAI222_X1 U22886 ( .A1(n19997), .A2(n19972), .B1(n19971), .B2(n19995), .C1(
        n19970), .C2(n19994), .ZN(P2_U3227) );
  OAI222_X1 U22887 ( .A1(n19997), .A2(n10834), .B1(n19973), .B2(n19995), .C1(
        n19972), .C2(n19994), .ZN(P2_U3228) );
  OAI222_X1 U22888 ( .A1(n19997), .A2(n19975), .B1(n19974), .B2(n19995), .C1(
        n10834), .C2(n19994), .ZN(P2_U3229) );
  OAI222_X1 U22889 ( .A1(n19997), .A2(n15188), .B1(n19976), .B2(n19995), .C1(
        n19975), .C2(n19994), .ZN(P2_U3230) );
  OAI222_X1 U22890 ( .A1(n19997), .A2(n10533), .B1(n19977), .B2(n19995), .C1(
        n15188), .C2(n19994), .ZN(P2_U3231) );
  OAI222_X1 U22891 ( .A1(n19997), .A2(n19979), .B1(n19978), .B2(n19995), .C1(
        n10533), .C2(n19994), .ZN(P2_U3232) );
  OAI222_X1 U22892 ( .A1(n19997), .A2(n19981), .B1(n19980), .B2(n19995), .C1(
        n19979), .C2(n19994), .ZN(P2_U3233) );
  OAI222_X1 U22893 ( .A1(n19997), .A2(n19983), .B1(n19982), .B2(n19995), .C1(
        n19981), .C2(n19994), .ZN(P2_U3234) );
  OAI222_X1 U22894 ( .A1(n19997), .A2(n19985), .B1(n19984), .B2(n19995), .C1(
        n19983), .C2(n19994), .ZN(P2_U3235) );
  OAI222_X1 U22895 ( .A1(n19997), .A2(n10850), .B1(n19986), .B2(n19995), .C1(
        n19985), .C2(n19994), .ZN(P2_U3236) );
  OAI222_X1 U22896 ( .A1(n19997), .A2(n19989), .B1(n19987), .B2(n19995), .C1(
        n10850), .C2(n19994), .ZN(P2_U3237) );
  OAI222_X1 U22897 ( .A1(n19994), .A2(n19989), .B1(n19988), .B2(n19995), .C1(
        n19990), .C2(n19997), .ZN(P2_U3238) );
  OAI222_X1 U22898 ( .A1(n19997), .A2(n19992), .B1(n19991), .B2(n19995), .C1(
        n19990), .C2(n19994), .ZN(P2_U3239) );
  OAI222_X1 U22899 ( .A1(n19997), .A2(n10859), .B1(n19993), .B2(n19995), .C1(
        n19992), .C2(n19994), .ZN(P2_U3240) );
  OAI222_X1 U22900 ( .A1(n19997), .A2(n12451), .B1(n19996), .B2(n19995), .C1(
        n10859), .C2(n19994), .ZN(P2_U3241) );
  OAI22_X1 U22901 ( .A1(n20052), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19995), .ZN(n19998) );
  INV_X1 U22902 ( .A(n19998), .ZN(P2_U3585) );
  MUX2_X1 U22903 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20052), .Z(P2_U3586) );
  OAI22_X1 U22904 ( .A1(n20052), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19995), .ZN(n19999) );
  INV_X1 U22905 ( .A(n19999), .ZN(P2_U3587) );
  AOI22_X1 U22906 ( .A1(n19995), .A2(n20000), .B1(n20998), .B2(n20052), .ZN(
        P2_U3588) );
  OAI21_X1 U22907 ( .B1(n20004), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20002), 
        .ZN(n20001) );
  INV_X1 U22908 ( .A(n20001), .ZN(P2_U3591) );
  OAI21_X1 U22909 ( .B1(n20004), .B2(n20003), .A(n20002), .ZN(P2_U3592) );
  NAND2_X1 U22910 ( .A1(n20005), .A2(n20006), .ZN(n20013) );
  NAND2_X1 U22911 ( .A1(n20006), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20029) );
  OR2_X1 U22912 ( .A1(n20007), .A2(n20029), .ZN(n20017) );
  NAND3_X1 U22913 ( .A1(n20028), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20008), 
        .ZN(n20009) );
  NAND2_X1 U22914 ( .A1(n20009), .A2(n20024), .ZN(n20018) );
  NAND2_X1 U22915 ( .A1(n20017), .A2(n20018), .ZN(n20011) );
  NAND2_X1 U22916 ( .A1(n20011), .A2(n20010), .ZN(n20012) );
  OAI211_X1 U22917 ( .C1(n20014), .C2(n19632), .A(n20013), .B(n20012), .ZN(
        n20015) );
  INV_X1 U22918 ( .A(n20015), .ZN(n20016) );
  AOI22_X1 U22919 ( .A1(n20040), .A2(n10561), .B1(n20016), .B2(n20041), .ZN(
        P2_U3602) );
  OAI21_X1 U22920 ( .B1(n20019), .B2(n20018), .A(n20017), .ZN(n20020) );
  AOI21_X1 U22921 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20021), .A(n20020), 
        .ZN(n20022) );
  AOI22_X1 U22922 ( .A1(n20040), .A2(n20023), .B1(n20022), .B2(n20041), .ZN(
        P2_U3603) );
  INV_X1 U22923 ( .A(n20024), .ZN(n20036) );
  AND2_X1 U22924 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20025) );
  OR3_X1 U22925 ( .A1(n20026), .A2(n20036), .A3(n20025), .ZN(n20027) );
  OAI21_X1 U22926 ( .B1(n20029), .B2(n20028), .A(n20027), .ZN(n20030) );
  AOI21_X1 U22927 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20031), .A(n20030), 
        .ZN(n20032) );
  AOI22_X1 U22928 ( .A1(n20040), .A2(n20033), .B1(n20032), .B2(n20041), .ZN(
        P2_U3604) );
  OAI22_X1 U22929 ( .A1(n20037), .A2(n20036), .B1(n20035), .B2(n20034), .ZN(
        n20038) );
  AOI21_X1 U22930 ( .B1(n20042), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20038), 
        .ZN(n20039) );
  OAI22_X1 U22931 ( .A1(n20042), .A2(n20041), .B1(n20040), .B2(n20039), .ZN(
        P2_U3605) );
  AOI22_X1 U22932 ( .A1(n19995), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20043), 
        .B2(n20052), .ZN(P2_U3608) );
  OAI22_X1 U22933 ( .A1(n20047), .A2(n20046), .B1(n20045), .B2(n20044), .ZN(
        n20049) );
  OR2_X1 U22934 ( .A1(n20049), .A2(n20048), .ZN(n20051) );
  MUX2_X1 U22935 ( .A(P2_MORE_REG_SCAN_IN), .B(n20051), .S(n20050), .Z(
        P2_U3609) );
  OAI22_X1 U22936 ( .A1(n20052), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19995), .ZN(n20053) );
  INV_X1 U22937 ( .A(n20053), .ZN(P2_U3611) );
  AND2_X1 U22938 ( .A1(n20878), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n20055) );
  INV_X1 U22939 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20054) );
  INV_X1 U22940 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20884) );
  NAND2_X1 U22941 ( .A1(n20884), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20932) );
  AOI21_X1 U22942 ( .B1(n20055), .B2(n20054), .A(n20948), .ZN(P1_U2802) );
  INV_X1 U22943 ( .A(n20056), .ZN(n20058) );
  OAI21_X1 U22944 ( .B1(n20058), .B2(n20057), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20059) );
  OAI21_X1 U22945 ( .B1(n20060), .B2(n20868), .A(n20059), .ZN(P1_U2803) );
  NAND2_X1 U22946 ( .A1(n20889), .A2(n20884), .ZN(n20877) );
  INV_X1 U22947 ( .A(n20877), .ZN(n20062) );
  OAI21_X1 U22948 ( .B1(n20062), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20960), .ZN(
        n20061) );
  OAI21_X1 U22949 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20960), .A(n20061), 
        .ZN(P1_U2804) );
  AOI21_X1 U22950 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20878), .A(n20948), 
        .ZN(n20938) );
  OAI21_X1 U22951 ( .B1(BS16), .B2(n20062), .A(n20938), .ZN(n20936) );
  OAI21_X1 U22952 ( .B1(n20938), .B2(n20736), .A(n20936), .ZN(P1_U2805) );
  OAI21_X1 U22953 ( .B1(n20065), .B2(n20064), .A(n20063), .ZN(P1_U2806) );
  NOR4_X1 U22954 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20069) );
  NOR4_X1 U22955 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20068) );
  NOR4_X1 U22956 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20067) );
  NOR4_X1 U22957 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20066) );
  NAND4_X1 U22958 ( .A1(n20069), .A2(n20068), .A3(n20067), .A4(n20066), .ZN(
        n20075) );
  NOR4_X1 U22959 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20073) );
  AOI211_X1 U22960 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20072) );
  NOR4_X1 U22961 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20071) );
  NOR4_X1 U22962 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20070) );
  NAND4_X1 U22963 ( .A1(n20073), .A2(n20072), .A3(n20071), .A4(n20070), .ZN(
        n20074) );
  NOR2_X1 U22964 ( .A1(n20075), .A2(n20074), .ZN(n20946) );
  INV_X1 U22965 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20077) );
  NOR3_X1 U22966 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20078) );
  OAI21_X1 U22967 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20078), .A(n20946), .ZN(
        n20076) );
  OAI21_X1 U22968 ( .B1(n20946), .B2(n20077), .A(n20076), .ZN(P1_U2807) );
  INV_X1 U22969 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20937) );
  AOI21_X1 U22970 ( .B1(n20939), .B2(n20937), .A(n20078), .ZN(n20080) );
  INV_X1 U22971 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20079) );
  INV_X1 U22972 ( .A(n20946), .ZN(n20941) );
  AOI22_X1 U22973 ( .A1(n20946), .A2(n20080), .B1(n20079), .B2(n20941), .ZN(
        P1_U2808) );
  AOI22_X1 U22974 ( .A1(n20140), .A2(n20081), .B1(n20143), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n20092) );
  AOI22_X1 U22975 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n20139), .B1(
        n20145), .B2(n20082), .ZN(n20091) );
  NOR2_X1 U22976 ( .A1(n20102), .A2(n20083), .ZN(n20085) );
  AOI21_X1 U22977 ( .B1(n20085), .B2(n20084), .A(n16236), .ZN(n20090) );
  INV_X1 U22978 ( .A(n20086), .ZN(n20088) );
  AOI22_X1 U22979 ( .A1(n20088), .A2(n20119), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n20087), .ZN(n20089) );
  NAND4_X1 U22980 ( .A1(n20092), .A2(n20091), .A3(n20090), .A4(n20089), .ZN(
        P1_U2831) );
  INV_X1 U22981 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20112) );
  NAND2_X1 U22982 ( .A1(n20094), .A2(n20093), .ZN(n20125) );
  NOR3_X1 U22983 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20100), .A3(n20125), .ZN(
        n20097) );
  NAND2_X1 U22984 ( .A1(n20143), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n20095) );
  NAND2_X1 U22985 ( .A1(n20095), .A2(n20227), .ZN(n20096) );
  NOR2_X1 U22986 ( .A1(n20097), .A2(n20096), .ZN(n20110) );
  NOR2_X1 U22987 ( .A1(n20099), .A2(n20098), .ZN(n20107) );
  INV_X1 U22988 ( .A(n20100), .ZN(n20101) );
  NOR2_X1 U22989 ( .A1(n20102), .A2(n20101), .ZN(n20103) );
  NOR2_X1 U22990 ( .A1(n20113), .A2(n20103), .ZN(n20123) );
  OAI22_X1 U22991 ( .A1(n20105), .A2(n20104), .B1(n20898), .B2(n20123), .ZN(
        n20106) );
  AOI211_X1 U22992 ( .C1(n20108), .C2(n20145), .A(n20107), .B(n20106), .ZN(
        n20109) );
  OAI211_X1 U22993 ( .C1(n20112), .C2(n20111), .A(n20110), .B(n20109), .ZN(
        P1_U2833) );
  NOR2_X1 U22994 ( .A1(n20896), .A2(n20113), .ZN(n20124) );
  NOR2_X1 U22995 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20124), .ZN(n20122) );
  INV_X1 U22996 ( .A(n20114), .ZN(n20115) );
  AOI22_X1 U22997 ( .A1(n20115), .A2(n20140), .B1(n20145), .B2(n20155), .ZN(
        n20121) );
  AOI21_X1 U22998 ( .B1(n20139), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16236), .ZN(n20116) );
  OAI21_X1 U22999 ( .B1(n20117), .B2(n20160), .A(n20116), .ZN(n20118) );
  AOI21_X1 U23000 ( .B1(n20158), .B2(n20119), .A(n20118), .ZN(n20120) );
  OAI211_X1 U23001 ( .C1(n20123), .C2(n20122), .A(n20121), .B(n20120), .ZN(
        P1_U2834) );
  AOI22_X1 U23002 ( .A1(n20143), .A2(P1_EBX_REG_5__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20139), .ZN(n20137) );
  AOI21_X1 U23003 ( .B1(n20896), .B2(n20125), .A(n20124), .ZN(n20131) );
  NAND2_X1 U23004 ( .A1(n20140), .A2(n20126), .ZN(n20127) );
  OAI21_X1 U23005 ( .B1(n20129), .B2(n20128), .A(n20127), .ZN(n20130) );
  OR2_X1 U23006 ( .A1(n20131), .A2(n20130), .ZN(n20135) );
  NOR2_X1 U23007 ( .A1(n20133), .A2(n20132), .ZN(n20134) );
  NOR2_X1 U23008 ( .A1(n20135), .A2(n20134), .ZN(n20136) );
  NAND3_X1 U23009 ( .A1(n20137), .A2(n20136), .A3(n20227), .ZN(P1_U2835) );
  INV_X1 U23010 ( .A(n20138), .ZN(n20141) );
  AOI222_X1 U23011 ( .A1(n20541), .A2(n20142), .B1(n20141), .B2(n20140), .C1(
        n20139), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20154) );
  AOI22_X1 U23012 ( .A1(n20145), .A2(n20144), .B1(n20143), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n20153) );
  AOI22_X1 U23013 ( .A1(n20148), .A2(n20147), .B1(P1_REIP_REG_3__SCAN_IN), 
        .B2(n20146), .ZN(n20152) );
  NAND2_X1 U23014 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20149) );
  OAI211_X1 U23015 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n20150), .B(n20149), .ZN(n20151) );
  NAND4_X1 U23016 ( .A1(n20154), .A2(n20153), .A3(n20152), .A4(n20151), .ZN(
        P1_U2837) );
  AOI22_X1 U23017 ( .A1(n20158), .A2(n20157), .B1(n20156), .B2(n20155), .ZN(
        n20159) );
  OAI21_X1 U23018 ( .B1(n20161), .B2(n20160), .A(n20159), .ZN(P1_U2866) );
  AOI22_X1 U23019 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20167), .B1(n20184), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20162) );
  OAI21_X1 U23020 ( .B1(n20163), .B2(n20165), .A(n20162), .ZN(P1_U2921) );
  INV_X1 U23021 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n20166) );
  AOI22_X1 U23022 ( .A1(P1_EAX_REG_14__SCAN_IN), .A2(n20167), .B1(n20184), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20164) );
  OAI21_X1 U23023 ( .B1(n20166), .B2(n20165), .A(n20164), .ZN(P1_U2922) );
  AOI22_X1 U23024 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20168) );
  OAI21_X1 U23025 ( .B1(n14386), .B2(n20187), .A(n20168), .ZN(P1_U2923) );
  AOI22_X1 U23026 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20169) );
  OAI21_X1 U23027 ( .B1(n14387), .B2(n20187), .A(n20169), .ZN(P1_U2924) );
  AOI22_X1 U23028 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20170) );
  OAI21_X1 U23029 ( .B1(n14390), .B2(n20187), .A(n20170), .ZN(P1_U2925) );
  AOI22_X1 U23030 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20171) );
  OAI21_X1 U23031 ( .B1(n14392), .B2(n20187), .A(n20171), .ZN(P1_U2926) );
  INV_X1 U23032 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20173) );
  AOI22_X1 U23033 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20172) );
  OAI21_X1 U23034 ( .B1(n20173), .B2(n20187), .A(n20172), .ZN(P1_U2927) );
  AOI22_X1 U23035 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20174) );
  OAI21_X1 U23036 ( .B1(n13625), .B2(n20187), .A(n20174), .ZN(P1_U2928) );
  AOI22_X1 U23037 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20175) );
  OAI21_X1 U23038 ( .B1(n11346), .B2(n20187), .A(n20175), .ZN(P1_U2929) );
  AOI22_X1 U23039 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20176) );
  OAI21_X1 U23040 ( .B1(n11334), .B2(n20187), .A(n20176), .ZN(P1_U2930) );
  AOI22_X1 U23041 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20177) );
  OAI21_X1 U23042 ( .B1(n20178), .B2(n20187), .A(n20177), .ZN(P1_U2931) );
  AOI22_X1 U23043 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20179) );
  OAI21_X1 U23044 ( .B1(n20180), .B2(n20187), .A(n20179), .ZN(P1_U2932) );
  AOI22_X1 U23045 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20181) );
  OAI21_X1 U23046 ( .B1(n11244), .B2(n20187), .A(n20181), .ZN(P1_U2933) );
  AOI22_X1 U23047 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20182) );
  OAI21_X1 U23048 ( .B1(n11191), .B2(n20187), .A(n20182), .ZN(P1_U2934) );
  AOI22_X1 U23049 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20183) );
  OAI21_X1 U23050 ( .B1(n11197), .B2(n20187), .A(n20183), .ZN(P1_U2935) );
  AOI22_X1 U23051 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20185), .B1(n20184), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20186) );
  OAI21_X1 U23052 ( .B1(n20982), .B2(n20187), .A(n20186), .ZN(P1_U2936) );
  AOI22_X1 U23053 ( .A1(n20217), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20220), .ZN(n20190) );
  INV_X1 U23054 ( .A(n20188), .ZN(n20189) );
  NAND2_X1 U23055 ( .A1(n20205), .A2(n20189), .ZN(n20207) );
  NAND2_X1 U23056 ( .A1(n20190), .A2(n20207), .ZN(P1_U2945) );
  AOI22_X1 U23057 ( .A1(n20217), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20220), .ZN(n20193) );
  INV_X1 U23058 ( .A(n20191), .ZN(n20192) );
  NAND2_X1 U23059 ( .A1(n20205), .A2(n20192), .ZN(n20209) );
  NAND2_X1 U23060 ( .A1(n20193), .A2(n20209), .ZN(P1_U2946) );
  AOI22_X1 U23061 ( .A1(n20217), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20220), .ZN(n20196) );
  INV_X1 U23062 ( .A(n20194), .ZN(n20195) );
  NAND2_X1 U23063 ( .A1(n20205), .A2(n20195), .ZN(n20213) );
  NAND2_X1 U23064 ( .A1(n20196), .A2(n20213), .ZN(P1_U2948) );
  AOI22_X1 U23065 ( .A1(n20217), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20220), .ZN(n20199) );
  INV_X1 U23066 ( .A(n20197), .ZN(n20198) );
  NAND2_X1 U23067 ( .A1(n20205), .A2(n20198), .ZN(n20215) );
  NAND2_X1 U23068 ( .A1(n20199), .A2(n20215), .ZN(P1_U2949) );
  AOI22_X1 U23069 ( .A1(n20217), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20220), .ZN(n20202) );
  INV_X1 U23070 ( .A(n20200), .ZN(n20201) );
  NAND2_X1 U23071 ( .A1(n20205), .A2(n20201), .ZN(n20218) );
  NAND2_X1 U23072 ( .A1(n20202), .A2(n20218), .ZN(P1_U2950) );
  AOI22_X1 U23073 ( .A1(n20217), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20220), .ZN(n20206) );
  INV_X1 U23074 ( .A(n20203), .ZN(n20204) );
  NAND2_X1 U23075 ( .A1(n20205), .A2(n20204), .ZN(n20221) );
  NAND2_X1 U23076 ( .A1(n20206), .A2(n20221), .ZN(P1_U2951) );
  AOI22_X1 U23077 ( .A1(n20217), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20220), .ZN(n20208) );
  NAND2_X1 U23078 ( .A1(n20208), .A2(n20207), .ZN(P1_U2960) );
  AOI22_X1 U23079 ( .A1(n20217), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20220), .ZN(n20210) );
  NAND2_X1 U23080 ( .A1(n20210), .A2(n20209), .ZN(P1_U2961) );
  AOI22_X1 U23081 ( .A1(n20217), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20220), .ZN(n20212) );
  NAND2_X1 U23082 ( .A1(n20212), .A2(n20211), .ZN(P1_U2962) );
  AOI22_X1 U23083 ( .A1(n20217), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20220), .ZN(n20214) );
  NAND2_X1 U23084 ( .A1(n20214), .A2(n20213), .ZN(P1_U2963) );
  AOI22_X1 U23085 ( .A1(n20217), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20220), .ZN(n20216) );
  NAND2_X1 U23086 ( .A1(n20216), .A2(n20215), .ZN(P1_U2964) );
  AOI22_X1 U23087 ( .A1(n20217), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20220), .ZN(n20219) );
  NAND2_X1 U23088 ( .A1(n20219), .A2(n20218), .ZN(P1_U2965) );
  AOI22_X1 U23089 ( .A1(n20217), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20220), .ZN(n20222) );
  NAND2_X1 U23090 ( .A1(n20222), .A2(n20221), .ZN(P1_U2966) );
  NAND2_X1 U23091 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20223), .ZN(
        n20238) );
  INV_X1 U23092 ( .A(n20224), .ZN(n20225) );
  AOI21_X1 U23093 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20226), .A(
        n20225), .ZN(n20228) );
  OAI22_X1 U23094 ( .A1(n20229), .A2(n20228), .B1(n20892), .B2(n20227), .ZN(
        n20233) );
  NOR2_X1 U23095 ( .A1(n20231), .A2(n20230), .ZN(n20232) );
  AOI211_X1 U23096 ( .C1(n16243), .C2(n20234), .A(n20233), .B(n20232), .ZN(
        n20235) );
  OAI221_X1 U23097 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20238), .C1(
        n20237), .C2(n20236), .A(n20235), .ZN(P1_U3029) );
  NOR2_X1 U23098 ( .A1(n20240), .A2(n20239), .ZN(P1_U3032) );
  INV_X1 U23099 ( .A(n20328), .ZN(n20244) );
  AOI22_X1 U23100 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n9637), .B1(DATAI_24_), 
        .B2(n9636), .ZN(n20747) );
  NAND2_X1 U23101 ( .A1(n20293), .A2(n20246), .ZN(n20802) );
  NOR3_X1 U23102 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20305) );
  NAND2_X1 U23103 ( .A1(n20696), .A2(n20305), .ZN(n20294) );
  OAI22_X1 U23104 ( .A1(n20865), .A2(n20747), .B1(n20802), .B2(n20294), .ZN(
        n20247) );
  INV_X1 U23105 ( .A(n20247), .ZN(n20261) );
  INV_X1 U23106 ( .A(n20596), .ZN(n20248) );
  NOR2_X1 U23107 ( .A1(n20248), .A2(n20542), .ZN(n20257) );
  INV_X1 U23108 ( .A(n20249), .ZN(n20256) );
  NAND2_X1 U23109 ( .A1(n20256), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20731) );
  INV_X1 U23110 ( .A(n20731), .ZN(n20250) );
  AOI21_X1 U23111 ( .B1(n20327), .B2(n20865), .A(n20736), .ZN(n20251) );
  NOR2_X1 U23112 ( .A1(n20251), .A2(n20706), .ZN(n20255) );
  NAND2_X1 U23113 ( .A1(n10215), .A2(n20667), .ZN(n20258) );
  AOI22_X1 U23114 ( .A1(n20255), .A2(n20258), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20294), .ZN(n20253) );
  OAI211_X1 U23115 ( .C1(n20257), .C2(n20870), .A(n20598), .B(n20253), .ZN(
        n20298) );
  NOR2_X2 U23116 ( .A1(n20254), .A2(n20413), .ZN(n20732) );
  INV_X1 U23117 ( .A(n20255), .ZN(n20259) );
  NOR2_X1 U23118 ( .A1(n20256), .A2(n20870), .ZN(n20414) );
  INV_X1 U23119 ( .A(n20414), .ZN(n20600) );
  INV_X1 U23120 ( .A(n20257), .ZN(n20408) );
  AOI22_X1 U23121 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20298), .B1(
        n20732), .B2(n20297), .ZN(n20260) );
  OAI211_X1 U23122 ( .C1(n20812), .C2(n20327), .A(n20261), .B(n20260), .ZN(
        P1_U3033) );
  AOI22_X1 U23123 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9637), .B1(DATAI_25_), 
        .B2(n9636), .ZN(n20753) );
  NAND2_X1 U23124 ( .A1(n20293), .A2(n20262), .ZN(n20814) );
  OAI22_X1 U23125 ( .A1(n20865), .A2(n20753), .B1(n20814), .B2(n20294), .ZN(
        n20263) );
  INV_X1 U23126 ( .A(n20263), .ZN(n20266) );
  NOR2_X2 U23127 ( .A1(n20264), .A2(n20413), .ZN(n20748) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20298), .B1(
        n20748), .B2(n20297), .ZN(n20265) );
  OAI211_X1 U23129 ( .C1(n20819), .C2(n20327), .A(n20266), .B(n20265), .ZN(
        P1_U3034) );
  AOI22_X1 U23130 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n9637), .B1(DATAI_18_), 
        .B2(n9636), .ZN(n20826) );
  NAND2_X1 U23131 ( .A1(n20293), .A2(n20267), .ZN(n20821) );
  OAI22_X1 U23132 ( .A1(n20865), .A2(n20759), .B1(n20821), .B2(n20294), .ZN(
        n20268) );
  INV_X1 U23133 ( .A(n20268), .ZN(n20271) );
  NOR2_X2 U23134 ( .A1(n20269), .A2(n20413), .ZN(n20754) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20298), .B1(
        n20754), .B2(n20297), .ZN(n20270) );
  OAI211_X1 U23136 ( .C1(n20826), .C2(n20327), .A(n20271), .B(n20270), .ZN(
        P1_U3035) );
  AOI22_X1 U23137 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9637), .B1(DATAI_27_), 
        .B2(n9636), .ZN(n20765) );
  NAND2_X1 U23138 ( .A1(n20293), .A2(n20272), .ZN(n20828) );
  OAI22_X1 U23139 ( .A1(n20865), .A2(n20765), .B1(n20828), .B2(n20294), .ZN(
        n20273) );
  INV_X1 U23140 ( .A(n20273), .ZN(n20276) );
  NOR2_X2 U23141 ( .A1(n20274), .A2(n20413), .ZN(n20760) );
  AOI22_X1 U23142 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20298), .B1(
        n20760), .B2(n20297), .ZN(n20275) );
  OAI211_X1 U23143 ( .C1(n20833), .C2(n20327), .A(n20276), .B(n20275), .ZN(
        P1_U3036) );
  AOI22_X1 U23144 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9637), .B1(DATAI_28_), 
        .B2(n9636), .ZN(n20771) );
  NAND2_X1 U23145 ( .A1(n20293), .A2(n11047), .ZN(n20835) );
  OAI22_X1 U23146 ( .A1(n20865), .A2(n20771), .B1(n20835), .B2(n20294), .ZN(
        n20277) );
  INV_X1 U23147 ( .A(n20277), .ZN(n20280) );
  NOR2_X2 U23148 ( .A1(n20278), .A2(n20413), .ZN(n20766) );
  AOI22_X1 U23149 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20298), .B1(
        n20766), .B2(n20297), .ZN(n20279) );
  OAI211_X1 U23150 ( .C1(n20840), .C2(n20327), .A(n20280), .B(n20279), .ZN(
        P1_U3037) );
  AOI22_X1 U23151 ( .A1(DATAI_21_), .A2(n9636), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n9637), .ZN(n20847) );
  NAND2_X1 U23152 ( .A1(n20293), .A2(n11965), .ZN(n20842) );
  OAI22_X1 U23153 ( .A1(n20865), .A2(n20777), .B1(n20842), .B2(n20294), .ZN(
        n20281) );
  INV_X1 U23154 ( .A(n20281), .ZN(n20284) );
  NOR2_X2 U23155 ( .A1(n20282), .A2(n20413), .ZN(n20772) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20298), .B1(
        n20772), .B2(n20297), .ZN(n20283) );
  OAI211_X1 U23157 ( .C1(n20847), .C2(n20327), .A(n20284), .B(n20283), .ZN(
        P1_U3038) );
  AOI22_X1 U23158 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9637), .B1(DATAI_30_), 
        .B2(n9636), .ZN(n20783) );
  NAND2_X1 U23159 ( .A1(n20293), .A2(n20285), .ZN(n20849) );
  OAI22_X1 U23160 ( .A1(n20865), .A2(n20783), .B1(n20849), .B2(n20294), .ZN(
        n20286) );
  INV_X1 U23161 ( .A(n20286), .ZN(n20289) );
  NOR2_X2 U23162 ( .A1(n20287), .A2(n20413), .ZN(n20778) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20298), .B1(
        n20778), .B2(n20297), .ZN(n20288) );
  OAI211_X1 U23164 ( .C1(n20854), .C2(n20327), .A(n20289), .B(n20288), .ZN(
        P1_U3039) );
  AOI22_X1 U23165 ( .A1(DATAI_31_), .A2(n9636), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n9637), .ZN(n20793) );
  NAND2_X1 U23166 ( .A1(n20293), .A2(n20292), .ZN(n20858) );
  OAI22_X1 U23167 ( .A1(n20865), .A2(n20793), .B1(n20858), .B2(n20294), .ZN(
        n20295) );
  INV_X1 U23168 ( .A(n20295), .ZN(n20300) );
  NOR2_X2 U23169 ( .A1(n20296), .A2(n20413), .ZN(n20785) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20298), .B1(
        n20785), .B2(n20297), .ZN(n20299) );
  OAI211_X1 U23171 ( .C1(n20866), .C2(n20327), .A(n20300), .B(n20299), .ZN(
        P1_U3040) );
  INV_X1 U23172 ( .A(n20305), .ZN(n20302) );
  NOR2_X1 U23173 ( .A1(n20696), .A2(n20302), .ZN(n20322) );
  INV_X1 U23174 ( .A(n20301), .ZN(n20697) );
  AOI21_X1 U23175 ( .B1(n10215), .B2(n20697), .A(n20322), .ZN(n20303) );
  OAI22_X1 U23176 ( .A1(n20303), .A2(n20706), .B1(n20302), .B2(n20870), .ZN(
        n20321) );
  AOI22_X1 U23177 ( .A1(n20733), .A2(n20322), .B1(n20321), .B2(n20732), .ZN(
        n20307) );
  OAI21_X1 U23178 ( .B1(n20371), .B2(n20704), .A(n20303), .ZN(n20304) );
  OAI221_X1 U23179 ( .B1(n20797), .B2(n20305), .C1(n20706), .C2(n20304), .A(
        n20806), .ZN(n20324) );
  INV_X1 U23180 ( .A(n20812), .ZN(n20744) );
  AOI22_X1 U23181 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20324), .B1(
        n20323), .B2(n20744), .ZN(n20306) );
  OAI211_X1 U23182 ( .C1(n20747), .C2(n20327), .A(n20307), .B(n20306), .ZN(
        P1_U3041) );
  AOI22_X1 U23183 ( .A1(n20749), .A2(n20322), .B1(n20321), .B2(n20748), .ZN(
        n20309) );
  INV_X1 U23184 ( .A(n20819), .ZN(n20750) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20324), .B1(
        n20323), .B2(n20750), .ZN(n20308) );
  OAI211_X1 U23186 ( .C1(n20753), .C2(n20327), .A(n20309), .B(n20308), .ZN(
        P1_U3042) );
  AOI22_X1 U23187 ( .A1(n20755), .A2(n20322), .B1(n20321), .B2(n20754), .ZN(
        n20311) );
  INV_X1 U23188 ( .A(n20826), .ZN(n20756) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20324), .B1(
        n20323), .B2(n20756), .ZN(n20310) );
  OAI211_X1 U23190 ( .C1(n20759), .C2(n20327), .A(n20311), .B(n20310), .ZN(
        P1_U3043) );
  AOI22_X1 U23191 ( .A1(n20761), .A2(n20322), .B1(n20321), .B2(n20760), .ZN(
        n20314) );
  INV_X1 U23192 ( .A(n20327), .ZN(n20312) );
  INV_X1 U23193 ( .A(n20765), .ZN(n20830) );
  AOI22_X1 U23194 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20324), .B1(
        n20312), .B2(n20830), .ZN(n20313) );
  OAI211_X1 U23195 ( .C1(n20833), .C2(n20364), .A(n20314), .B(n20313), .ZN(
        P1_U3044) );
  AOI22_X1 U23196 ( .A1(n20767), .A2(n20322), .B1(n20321), .B2(n20766), .ZN(
        n20316) );
  INV_X1 U23197 ( .A(n20840), .ZN(n20768) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20324), .B1(
        n20323), .B2(n20768), .ZN(n20315) );
  OAI211_X1 U23199 ( .C1(n20771), .C2(n20327), .A(n20316), .B(n20315), .ZN(
        P1_U3045) );
  AOI22_X1 U23200 ( .A1(n20773), .A2(n20322), .B1(n20321), .B2(n20772), .ZN(
        n20318) );
  INV_X1 U23201 ( .A(n20847), .ZN(n20774) );
  AOI22_X1 U23202 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20324), .B1(
        n20323), .B2(n20774), .ZN(n20317) );
  OAI211_X1 U23203 ( .C1(n20777), .C2(n20327), .A(n20318), .B(n20317), .ZN(
        P1_U3046) );
  AOI22_X1 U23204 ( .A1(n20779), .A2(n20322), .B1(n20321), .B2(n20778), .ZN(
        n20320) );
  INV_X1 U23205 ( .A(n20854), .ZN(n20780) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20324), .B1(
        n20323), .B2(n20780), .ZN(n20319) );
  OAI211_X1 U23207 ( .C1(n20783), .C2(n20327), .A(n20320), .B(n20319), .ZN(
        P1_U3047) );
  AOI22_X1 U23208 ( .A1(n20787), .A2(n20322), .B1(n20321), .B2(n20785), .ZN(
        n20326) );
  INV_X1 U23209 ( .A(n20866), .ZN(n20788) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20324), .B1(
        n20323), .B2(n20788), .ZN(n20325) );
  OAI211_X1 U23211 ( .C1(n20793), .C2(n20327), .A(n20326), .B(n20325), .ZN(
        P1_U3048) );
  INV_X1 U23212 ( .A(n20734), .ZN(n20329) );
  NAND3_X1 U23213 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20662), .A3(
        n20663), .ZN(n20375) );
  NOR2_X1 U23214 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20375), .ZN(
        n20332) );
  INV_X1 U23215 ( .A(n20332), .ZN(n20358) );
  OAI22_X1 U23216 ( .A1(n20399), .A2(n20812), .B1(n20802), .B2(n20358), .ZN(
        n20330) );
  INV_X1 U23217 ( .A(n20330), .ZN(n20339) );
  NAND2_X1 U23218 ( .A1(n20399), .A2(n20364), .ZN(n20331) );
  AOI21_X1 U23219 ( .B1(n20331), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20706), 
        .ZN(n20335) );
  NAND2_X1 U23220 ( .A1(n10215), .A2(n20739), .ZN(n20336) );
  NOR2_X1 U23221 ( .A1(n20332), .A2(n20669), .ZN(n20333) );
  AOI21_X1 U23222 ( .B1(n20335), .B2(n20336), .A(n20333), .ZN(n20334) );
  OR2_X1 U23223 ( .A1(n20596), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20472) );
  NAND2_X1 U23224 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20472), .ZN(n20469) );
  NAND3_X1 U23225 ( .A1(n20598), .A2(n20334), .A3(n20469), .ZN(n20361) );
  INV_X1 U23226 ( .A(n20335), .ZN(n20337) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20361), .B1(
        n20732), .B2(n20360), .ZN(n20338) );
  OAI211_X1 U23228 ( .C1(n20747), .C2(n20364), .A(n20339), .B(n20338), .ZN(
        P1_U3049) );
  OAI22_X1 U23229 ( .A1(n20364), .A2(n20753), .B1(n20358), .B2(n20814), .ZN(
        n20340) );
  INV_X1 U23230 ( .A(n20340), .ZN(n20342) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20361), .B1(
        n20748), .B2(n20360), .ZN(n20341) );
  OAI211_X1 U23232 ( .C1(n20819), .C2(n20399), .A(n20342), .B(n20341), .ZN(
        P1_U3050) );
  OAI22_X1 U23233 ( .A1(n20399), .A2(n20826), .B1(n20358), .B2(n20821), .ZN(
        n20343) );
  INV_X1 U23234 ( .A(n20343), .ZN(n20345) );
  AOI22_X1 U23235 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20361), .B1(
        n20754), .B2(n20360), .ZN(n20344) );
  OAI211_X1 U23236 ( .C1(n20759), .C2(n20364), .A(n20345), .B(n20344), .ZN(
        P1_U3051) );
  OAI22_X1 U23237 ( .A1(n20364), .A2(n20765), .B1(n20358), .B2(n20828), .ZN(
        n20346) );
  INV_X1 U23238 ( .A(n20346), .ZN(n20348) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20361), .B1(
        n20760), .B2(n20360), .ZN(n20347) );
  OAI211_X1 U23240 ( .C1(n20833), .C2(n20399), .A(n20348), .B(n20347), .ZN(
        P1_U3052) );
  OAI22_X1 U23241 ( .A1(n20399), .A2(n20840), .B1(n20358), .B2(n20835), .ZN(
        n20349) );
  INV_X1 U23242 ( .A(n20349), .ZN(n20351) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20361), .B1(
        n20766), .B2(n20360), .ZN(n20350) );
  OAI211_X1 U23244 ( .C1(n20771), .C2(n20364), .A(n20351), .B(n20350), .ZN(
        P1_U3053) );
  OAI22_X1 U23245 ( .A1(n20364), .A2(n20777), .B1(n20358), .B2(n20842), .ZN(
        n20352) );
  INV_X1 U23246 ( .A(n20352), .ZN(n20354) );
  AOI22_X1 U23247 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20361), .B1(
        n20772), .B2(n20360), .ZN(n20353) );
  OAI211_X1 U23248 ( .C1(n20847), .C2(n20399), .A(n20354), .B(n20353), .ZN(
        P1_U3054) );
  OAI22_X1 U23249 ( .A1(n20399), .A2(n20854), .B1(n20358), .B2(n20849), .ZN(
        n20355) );
  INV_X1 U23250 ( .A(n20355), .ZN(n20357) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20361), .B1(
        n20778), .B2(n20360), .ZN(n20356) );
  OAI211_X1 U23252 ( .C1(n20783), .C2(n20364), .A(n20357), .B(n20356), .ZN(
        P1_U3055) );
  OAI22_X1 U23253 ( .A1(n20399), .A2(n20866), .B1(n20358), .B2(n20858), .ZN(
        n20359) );
  INV_X1 U23254 ( .A(n20359), .ZN(n20363) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20361), .B1(
        n20785), .B2(n20360), .ZN(n20362) );
  OAI211_X1 U23256 ( .C1(n20793), .C2(n20364), .A(n20363), .B(n20362), .ZN(
        P1_U3056) );
  INV_X1 U23257 ( .A(n20630), .ZN(n20365) );
  INV_X1 U23258 ( .A(n20632), .ZN(n20366) );
  NAND2_X1 U23259 ( .A1(n20366), .A2(n20662), .ZN(n20398) );
  OAI22_X1 U23260 ( .A1(n20399), .A2(n20747), .B1(n20802), .B2(n20398), .ZN(
        n20367) );
  INV_X1 U23261 ( .A(n20367), .ZN(n20379) );
  AND2_X1 U23262 ( .A1(n20369), .A2(n20368), .ZN(n20794) );
  INV_X1 U23263 ( .A(n20398), .ZN(n20370) );
  AOI21_X1 U23264 ( .B1(n10215), .B2(n20794), .A(n20370), .ZN(n20377) );
  OR2_X1 U23265 ( .A1(n20371), .A2(n20636), .ZN(n20372) );
  AOI22_X1 U23266 ( .A1(n20377), .A2(n20374), .B1(n20706), .B2(n20375), .ZN(
        n20373) );
  NAND2_X1 U23267 ( .A1(n20806), .A2(n20373), .ZN(n20402) );
  INV_X1 U23268 ( .A(n20374), .ZN(n20376) );
  OAI22_X1 U23269 ( .A1(n20377), .A2(n20376), .B1(n20870), .B2(n20375), .ZN(
        n20401) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20402), .B1(
        n20732), .B2(n20401), .ZN(n20378) );
  OAI211_X1 U23271 ( .C1(n20812), .C2(n20409), .A(n20379), .B(n20378), .ZN(
        P1_U3057) );
  OAI22_X1 U23272 ( .A1(n20399), .A2(n20753), .B1(n20398), .B2(n20814), .ZN(
        n20380) );
  INV_X1 U23273 ( .A(n20380), .ZN(n20382) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20402), .B1(
        n20748), .B2(n20401), .ZN(n20381) );
  OAI211_X1 U23275 ( .C1(n20819), .C2(n20409), .A(n20382), .B(n20381), .ZN(
        P1_U3058) );
  OAI22_X1 U23276 ( .A1(n20399), .A2(n20759), .B1(n20821), .B2(n20398), .ZN(
        n20383) );
  INV_X1 U23277 ( .A(n20383), .ZN(n20385) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20402), .B1(
        n20754), .B2(n20401), .ZN(n20384) );
  OAI211_X1 U23279 ( .C1(n20826), .C2(n20409), .A(n20385), .B(n20384), .ZN(
        P1_U3059) );
  OAI22_X1 U23280 ( .A1(n20409), .A2(n20833), .B1(n20398), .B2(n20828), .ZN(
        n20386) );
  INV_X1 U23281 ( .A(n20386), .ZN(n20388) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20402), .B1(
        n20760), .B2(n20401), .ZN(n20387) );
  OAI211_X1 U23283 ( .C1(n20765), .C2(n20399), .A(n20388), .B(n20387), .ZN(
        P1_U3060) );
  OAI22_X1 U23284 ( .A1(n20399), .A2(n20771), .B1(n20835), .B2(n20398), .ZN(
        n20389) );
  INV_X1 U23285 ( .A(n20389), .ZN(n20391) );
  AOI22_X1 U23286 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20402), .B1(
        n20766), .B2(n20401), .ZN(n20390) );
  OAI211_X1 U23287 ( .C1(n20840), .C2(n20409), .A(n20391), .B(n20390), .ZN(
        P1_U3061) );
  OAI22_X1 U23288 ( .A1(n20409), .A2(n20847), .B1(n20398), .B2(n20842), .ZN(
        n20392) );
  INV_X1 U23289 ( .A(n20392), .ZN(n20394) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20402), .B1(
        n20772), .B2(n20401), .ZN(n20393) );
  OAI211_X1 U23291 ( .C1(n20777), .C2(n20399), .A(n20394), .B(n20393), .ZN(
        P1_U3062) );
  OAI22_X1 U23292 ( .A1(n20399), .A2(n20783), .B1(n20849), .B2(n20398), .ZN(
        n20395) );
  INV_X1 U23293 ( .A(n20395), .ZN(n20397) );
  AOI22_X1 U23294 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20402), .B1(
        n20778), .B2(n20401), .ZN(n20396) );
  OAI211_X1 U23295 ( .C1(n20854), .C2(n20409), .A(n20397), .B(n20396), .ZN(
        P1_U3063) );
  OAI22_X1 U23296 ( .A1(n20399), .A2(n20793), .B1(n20858), .B2(n20398), .ZN(
        n20400) );
  INV_X1 U23297 ( .A(n20400), .ZN(n20404) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20402), .B1(
        n20785), .B2(n20401), .ZN(n20403) );
  OAI211_X1 U23299 ( .C1(n20866), .C2(n20409), .A(n20404), .B(n20403), .ZN(
        P1_U3064) );
  NOR3_X1 U23300 ( .A1(n20663), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20444) );
  INV_X1 U23301 ( .A(n20444), .ZN(n20436) );
  NOR2_X1 U23302 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20436), .ZN(
        n20431) );
  NOR2_X1 U23303 ( .A1(n13162), .A2(n20406), .ZN(n20503) );
  NAND3_X1 U23304 ( .A1(n20503), .A2(n20797), .A3(n20667), .ZN(n20407) );
  OAI21_X1 U23305 ( .B1(n20731), .B2(n20408), .A(n20407), .ZN(n20430) );
  AOI22_X1 U23306 ( .A1(n20733), .A2(n20431), .B1(n20732), .B2(n20430), .ZN(
        n20417) );
  INV_X1 U23307 ( .A(n20503), .ZN(n20412) );
  INV_X1 U23308 ( .A(n20466), .ZN(n20410) );
  OAI21_X1 U23309 ( .B1(n20432), .B2(n20410), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20411) );
  OAI21_X1 U23310 ( .B1(n20739), .B2(n20412), .A(n20411), .ZN(n20415) );
  INV_X1 U23311 ( .A(n20747), .ZN(n20809) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n20809), .ZN(n20416) );
  OAI211_X1 U23313 ( .C1(n20812), .C2(n20466), .A(n20417), .B(n20416), .ZN(
        P1_U3065) );
  AOI22_X1 U23314 ( .A1(n20749), .A2(n20431), .B1(n20748), .B2(n20430), .ZN(
        n20419) );
  INV_X1 U23315 ( .A(n20753), .ZN(n20816) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n20816), .ZN(n20418) );
  OAI211_X1 U23317 ( .C1(n20819), .C2(n20466), .A(n20419), .B(n20418), .ZN(
        P1_U3066) );
  AOI22_X1 U23318 ( .A1(n20755), .A2(n20431), .B1(n20754), .B2(n20430), .ZN(
        n20421) );
  INV_X1 U23319 ( .A(n20759), .ZN(n20823) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n20823), .ZN(n20420) );
  OAI211_X1 U23321 ( .C1(n20826), .C2(n20466), .A(n20421), .B(n20420), .ZN(
        P1_U3067) );
  AOI22_X1 U23322 ( .A1(n20761), .A2(n20431), .B1(n20760), .B2(n20430), .ZN(
        n20423) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n20830), .ZN(n20422) );
  OAI211_X1 U23324 ( .C1(n20833), .C2(n20466), .A(n20423), .B(n20422), .ZN(
        P1_U3068) );
  AOI22_X1 U23325 ( .A1(n20767), .A2(n20431), .B1(n20766), .B2(n20430), .ZN(
        n20425) );
  INV_X1 U23326 ( .A(n20771), .ZN(n20837) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n20837), .ZN(n20424) );
  OAI211_X1 U23328 ( .C1(n20840), .C2(n20466), .A(n20425), .B(n20424), .ZN(
        P1_U3069) );
  AOI22_X1 U23329 ( .A1(n20773), .A2(n20431), .B1(n20772), .B2(n20430), .ZN(
        n20427) );
  INV_X1 U23330 ( .A(n20777), .ZN(n20844) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n20844), .ZN(n20426) );
  OAI211_X1 U23332 ( .C1(n20847), .C2(n20466), .A(n20427), .B(n20426), .ZN(
        P1_U3070) );
  AOI22_X1 U23333 ( .A1(n20779), .A2(n20431), .B1(n20778), .B2(n20430), .ZN(
        n20429) );
  INV_X1 U23334 ( .A(n20783), .ZN(n20851) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n20851), .ZN(n20428) );
  OAI211_X1 U23336 ( .C1(n20854), .C2(n20466), .A(n20429), .B(n20428), .ZN(
        P1_U3071) );
  AOI22_X1 U23337 ( .A1(n20787), .A2(n20431), .B1(n20785), .B2(n20430), .ZN(
        n20435) );
  INV_X1 U23338 ( .A(n20793), .ZN(n20860) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n20860), .ZN(n20434) );
  OAI211_X1 U23340 ( .C1(n20866), .C2(n20466), .A(n20435), .B(n20434), .ZN(
        P1_U3072) );
  NOR2_X1 U23341 ( .A1(n20696), .A2(n20436), .ZN(n20461) );
  NAND2_X1 U23342 ( .A1(n20503), .A2(n20697), .ZN(n20438) );
  INV_X1 U23343 ( .A(n20461), .ZN(n20437) );
  NAND2_X1 U23344 ( .A1(n20438), .A2(n20437), .ZN(n20441) );
  NAND2_X1 U23345 ( .A1(n20441), .A2(n20797), .ZN(n20440) );
  NAND2_X1 U23346 ( .A1(n20444), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20439) );
  NAND2_X1 U23347 ( .A1(n20440), .A2(n20439), .ZN(n20460) );
  AOI22_X1 U23348 ( .A1(n20733), .A2(n20461), .B1(n20732), .B2(n20460), .ZN(
        n20447) );
  INV_X1 U23349 ( .A(n20502), .ZN(n20510) );
  INV_X1 U23350 ( .A(n20441), .ZN(n20442) );
  OAI21_X1 U23351 ( .B1(n20510), .B2(n20704), .A(n20442), .ZN(n20443) );
  OAI221_X1 U23352 ( .B1(n20797), .B2(n20444), .C1(n20706), .C2(n20443), .A(
        n20806), .ZN(n20463) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20463), .B1(
        n20462), .B2(n20744), .ZN(n20446) );
  OAI211_X1 U23354 ( .C1(n20747), .C2(n20466), .A(n20447), .B(n20446), .ZN(
        P1_U3073) );
  AOI22_X1 U23355 ( .A1(n20749), .A2(n20461), .B1(n20748), .B2(n20460), .ZN(
        n20449) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20463), .B1(
        n20462), .B2(n20750), .ZN(n20448) );
  OAI211_X1 U23357 ( .C1(n20753), .C2(n20466), .A(n20449), .B(n20448), .ZN(
        P1_U3074) );
  AOI22_X1 U23358 ( .A1(n20755), .A2(n20461), .B1(n20754), .B2(n20460), .ZN(
        n20451) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20463), .B1(
        n20462), .B2(n20756), .ZN(n20450) );
  OAI211_X1 U23360 ( .C1(n20759), .C2(n20466), .A(n20451), .B(n20450), .ZN(
        P1_U3075) );
  AOI22_X1 U23361 ( .A1(n20761), .A2(n20461), .B1(n20760), .B2(n20460), .ZN(
        n20453) );
  INV_X1 U23362 ( .A(n20833), .ZN(n20762) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20463), .B1(
        n20462), .B2(n20762), .ZN(n20452) );
  OAI211_X1 U23364 ( .C1(n20765), .C2(n20466), .A(n20453), .B(n20452), .ZN(
        P1_U3076) );
  AOI22_X1 U23365 ( .A1(n20767), .A2(n20461), .B1(n20766), .B2(n20460), .ZN(
        n20455) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20463), .B1(
        n20462), .B2(n20768), .ZN(n20454) );
  OAI211_X1 U23367 ( .C1(n20771), .C2(n20466), .A(n20455), .B(n20454), .ZN(
        P1_U3077) );
  AOI22_X1 U23368 ( .A1(n20773), .A2(n20461), .B1(n20772), .B2(n20460), .ZN(
        n20457) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20463), .B1(
        n20462), .B2(n20774), .ZN(n20456) );
  OAI211_X1 U23370 ( .C1(n20777), .C2(n20466), .A(n20457), .B(n20456), .ZN(
        P1_U3078) );
  AOI22_X1 U23371 ( .A1(n20779), .A2(n20461), .B1(n20778), .B2(n20460), .ZN(
        n20459) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20463), .B1(
        n20462), .B2(n20780), .ZN(n20458) );
  OAI211_X1 U23373 ( .C1(n20783), .C2(n20466), .A(n20459), .B(n20458), .ZN(
        P1_U3079) );
  AOI22_X1 U23374 ( .A1(n20787), .A2(n20461), .B1(n20785), .B2(n20460), .ZN(
        n20465) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20463), .B1(
        n20462), .B2(n20788), .ZN(n20464) );
  OAI211_X1 U23376 ( .C1(n20793), .C2(n20466), .A(n20465), .B(n20464), .ZN(
        P1_U3080) );
  NAND2_X1 U23377 ( .A1(n20696), .A2(n10233), .ZN(n20495) );
  OAI22_X1 U23378 ( .A1(n20529), .A2(n20812), .B1(n20802), .B2(n20495), .ZN(
        n20467) );
  INV_X1 U23379 ( .A(n20467), .ZN(n20476) );
  AOI21_X1 U23380 ( .B1(n20529), .B2(n20501), .A(n20736), .ZN(n20468) );
  NOR2_X1 U23381 ( .A1(n20468), .A2(n20706), .ZN(n20471) );
  NAND2_X1 U23382 ( .A1(n20503), .A2(n20739), .ZN(n20473) );
  AOI22_X1 U23383 ( .A1(n20471), .A2(n20473), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20495), .ZN(n20470) );
  NAND3_X1 U23384 ( .A1(n20742), .A2(n20470), .A3(n20469), .ZN(n20498) );
  INV_X1 U23385 ( .A(n20471), .ZN(n20474) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20498), .B1(
        n20732), .B2(n20497), .ZN(n20475) );
  OAI211_X1 U23387 ( .C1(n20747), .C2(n20501), .A(n20476), .B(n20475), .ZN(
        P1_U3081) );
  OAI22_X1 U23388 ( .A1(n20529), .A2(n20819), .B1(n20814), .B2(n20495), .ZN(
        n20477) );
  INV_X1 U23389 ( .A(n20477), .ZN(n20479) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20498), .B1(
        n20748), .B2(n20497), .ZN(n20478) );
  OAI211_X1 U23391 ( .C1(n20753), .C2(n20501), .A(n20479), .B(n20478), .ZN(
        P1_U3082) );
  OAI22_X1 U23392 ( .A1(n20501), .A2(n20759), .B1(n20821), .B2(n20495), .ZN(
        n20480) );
  INV_X1 U23393 ( .A(n20480), .ZN(n20482) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20498), .B1(
        n20754), .B2(n20497), .ZN(n20481) );
  OAI211_X1 U23395 ( .C1(n20826), .C2(n20529), .A(n20482), .B(n20481), .ZN(
        P1_U3083) );
  OAI22_X1 U23396 ( .A1(n20501), .A2(n20765), .B1(n20828), .B2(n20495), .ZN(
        n20483) );
  INV_X1 U23397 ( .A(n20483), .ZN(n20485) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20498), .B1(
        n20760), .B2(n20497), .ZN(n20484) );
  OAI211_X1 U23399 ( .C1(n20833), .C2(n20529), .A(n20485), .B(n20484), .ZN(
        P1_U3084) );
  OAI22_X1 U23400 ( .A1(n20501), .A2(n20771), .B1(n20835), .B2(n20495), .ZN(
        n20486) );
  INV_X1 U23401 ( .A(n20486), .ZN(n20488) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20498), .B1(
        n20766), .B2(n20497), .ZN(n20487) );
  OAI211_X1 U23403 ( .C1(n20840), .C2(n20529), .A(n20488), .B(n20487), .ZN(
        P1_U3085) );
  OAI22_X1 U23404 ( .A1(n20529), .A2(n20847), .B1(n20842), .B2(n20495), .ZN(
        n20489) );
  INV_X1 U23405 ( .A(n20489), .ZN(n20491) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20498), .B1(
        n20772), .B2(n20497), .ZN(n20490) );
  OAI211_X1 U23407 ( .C1(n20777), .C2(n20501), .A(n20491), .B(n20490), .ZN(
        P1_U3086) );
  OAI22_X1 U23408 ( .A1(n20501), .A2(n20783), .B1(n20849), .B2(n20495), .ZN(
        n20492) );
  INV_X1 U23409 ( .A(n20492), .ZN(n20494) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20498), .B1(
        n20778), .B2(n20497), .ZN(n20493) );
  OAI211_X1 U23411 ( .C1(n20854), .C2(n20529), .A(n20494), .B(n20493), .ZN(
        P1_U3087) );
  OAI22_X1 U23412 ( .A1(n20529), .A2(n20866), .B1(n20858), .B2(n20495), .ZN(
        n20496) );
  INV_X1 U23413 ( .A(n20496), .ZN(n20500) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20498), .B1(
        n20785), .B2(n20497), .ZN(n20499) );
  OAI211_X1 U23415 ( .C1(n20793), .C2(n20501), .A(n20500), .B(n20499), .ZN(
        P1_U3088) );
  NAND2_X1 U23416 ( .A1(n20502), .A2(n20630), .ZN(n20540) );
  NAND2_X1 U23417 ( .A1(n20503), .A2(n20794), .ZN(n20504) );
  NAND2_X1 U23418 ( .A1(n20504), .A2(n20534), .ZN(n20505) );
  NAND2_X1 U23419 ( .A1(n20505), .A2(n20797), .ZN(n20507) );
  NAND2_X1 U23420 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n10233), .ZN(n20506) );
  INV_X1 U23421 ( .A(n20732), .ZN(n20801) );
  OAI22_X1 U23422 ( .A1(n20802), .A2(n20534), .B1(n20533), .B2(n20801), .ZN(
        n20508) );
  INV_X1 U23423 ( .A(n20508), .ZN(n20513) );
  INV_X1 U23424 ( .A(n20636), .ZN(n20509) );
  NAND2_X1 U23425 ( .A1(n20509), .A2(n20797), .ZN(n20804) );
  NOR2_X1 U23426 ( .A1(n20510), .A2(n20804), .ZN(n20511) );
  OAI21_X1 U23427 ( .B1(n20511), .B2(n10233), .A(n20806), .ZN(n20537) );
  INV_X1 U23428 ( .A(n20529), .ZN(n20536) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20809), .ZN(n20512) );
  OAI211_X1 U23430 ( .C1(n20812), .C2(n20540), .A(n20513), .B(n20512), .ZN(
        P1_U3089) );
  INV_X1 U23431 ( .A(n20748), .ZN(n20813) );
  OAI22_X1 U23432 ( .A1(n20814), .A2(n20534), .B1(n20533), .B2(n20813), .ZN(
        n20514) );
  INV_X1 U23433 ( .A(n20514), .ZN(n20516) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20816), .ZN(n20515) );
  OAI211_X1 U23435 ( .C1(n20819), .C2(n20540), .A(n20516), .B(n20515), .ZN(
        P1_U3090) );
  INV_X1 U23436 ( .A(n20754), .ZN(n20820) );
  OAI22_X1 U23437 ( .A1(n20821), .A2(n20534), .B1(n20533), .B2(n20820), .ZN(
        n20517) );
  INV_X1 U23438 ( .A(n20517), .ZN(n20519) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20537), .B1(
        n20563), .B2(n20756), .ZN(n20518) );
  OAI211_X1 U23440 ( .C1(n20759), .C2(n20529), .A(n20519), .B(n20518), .ZN(
        P1_U3091) );
  INV_X1 U23441 ( .A(n20760), .ZN(n20827) );
  OAI22_X1 U23442 ( .A1(n20828), .A2(n20534), .B1(n20533), .B2(n20827), .ZN(
        n20520) );
  INV_X1 U23443 ( .A(n20520), .ZN(n20522) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20537), .B1(
        n20563), .B2(n20762), .ZN(n20521) );
  OAI211_X1 U23445 ( .C1(n20765), .C2(n20529), .A(n20522), .B(n20521), .ZN(
        P1_U3092) );
  INV_X1 U23446 ( .A(n20766), .ZN(n20834) );
  OAI22_X1 U23447 ( .A1(n20835), .A2(n20534), .B1(n20533), .B2(n20834), .ZN(
        n20523) );
  INV_X1 U23448 ( .A(n20523), .ZN(n20525) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20837), .ZN(n20524) );
  OAI211_X1 U23450 ( .C1(n20840), .C2(n20540), .A(n20525), .B(n20524), .ZN(
        P1_U3093) );
  INV_X1 U23451 ( .A(n20772), .ZN(n20841) );
  OAI22_X1 U23452 ( .A1(n20842), .A2(n20534), .B1(n20533), .B2(n20841), .ZN(
        n20526) );
  INV_X1 U23453 ( .A(n20526), .ZN(n20528) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20537), .B1(
        n20563), .B2(n20774), .ZN(n20527) );
  OAI211_X1 U23455 ( .C1(n20777), .C2(n20529), .A(n20528), .B(n20527), .ZN(
        P1_U3094) );
  INV_X1 U23456 ( .A(n20778), .ZN(n20848) );
  OAI22_X1 U23457 ( .A1(n20849), .A2(n20534), .B1(n20533), .B2(n20848), .ZN(
        n20530) );
  INV_X1 U23458 ( .A(n20530), .ZN(n20532) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20851), .ZN(n20531) );
  OAI211_X1 U23460 ( .C1(n20854), .C2(n20540), .A(n20532), .B(n20531), .ZN(
        P1_U3095) );
  INV_X1 U23461 ( .A(n20785), .ZN(n20855) );
  OAI22_X1 U23462 ( .A1(n20858), .A2(n20534), .B1(n20533), .B2(n20855), .ZN(
        n20535) );
  INV_X1 U23463 ( .A(n20535), .ZN(n20539) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20860), .ZN(n20538) );
  OAI211_X1 U23465 ( .C1(n20866), .C2(n20540), .A(n20539), .B(n20538), .ZN(
        P1_U3096) );
  NOR3_X1 U23466 ( .A1(n20662), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20570) );
  INV_X1 U23467 ( .A(n20570), .ZN(n20567) );
  NOR2_X1 U23468 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20567), .ZN(
        n20562) );
  NAND2_X1 U23469 ( .A1(n20541), .A2(n13162), .ZN(n20595) );
  INV_X1 U23470 ( .A(n20595), .ZN(n20633) );
  AOI21_X1 U23471 ( .B1(n20633), .B2(n20667), .A(n20562), .ZN(n20544) );
  NAND2_X1 U23472 ( .A1(n20542), .A2(n20596), .ZN(n20671) );
  OAI22_X1 U23473 ( .A1(n20544), .A2(n20706), .B1(n20600), .B2(n20671), .ZN(
        n20561) );
  AOI22_X1 U23474 ( .A1(n20733), .A2(n20562), .B1(n20561), .B2(n20732), .ZN(
        n20548) );
  INV_X1 U23475 ( .A(n20591), .ZN(n20543) );
  OAI21_X1 U23476 ( .B1(n20543), .B2(n20563), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20545) );
  NAND2_X1 U23477 ( .A1(n20545), .A2(n20544), .ZN(n20546) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20809), .ZN(n20547) );
  OAI211_X1 U23479 ( .C1(n20812), .C2(n20591), .A(n20548), .B(n20547), .ZN(
        P1_U3097) );
  AOI22_X1 U23480 ( .A1(n20749), .A2(n20562), .B1(n20561), .B2(n20748), .ZN(
        n20550) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20816), .ZN(n20549) );
  OAI211_X1 U23482 ( .C1(n20819), .C2(n20591), .A(n20550), .B(n20549), .ZN(
        P1_U3098) );
  AOI22_X1 U23483 ( .A1(n20755), .A2(n20562), .B1(n20561), .B2(n20754), .ZN(
        n20552) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20823), .ZN(n20551) );
  OAI211_X1 U23485 ( .C1(n20826), .C2(n20591), .A(n20552), .B(n20551), .ZN(
        P1_U3099) );
  AOI22_X1 U23486 ( .A1(n20761), .A2(n20562), .B1(n20561), .B2(n20760), .ZN(
        n20554) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20830), .ZN(n20553) );
  OAI211_X1 U23488 ( .C1(n20833), .C2(n20591), .A(n20554), .B(n20553), .ZN(
        P1_U3100) );
  AOI22_X1 U23489 ( .A1(n20767), .A2(n20562), .B1(n20561), .B2(n20766), .ZN(
        n20556) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20837), .ZN(n20555) );
  OAI211_X1 U23491 ( .C1(n20840), .C2(n20591), .A(n20556), .B(n20555), .ZN(
        P1_U3101) );
  AOI22_X1 U23492 ( .A1(n20773), .A2(n20562), .B1(n20561), .B2(n20772), .ZN(
        n20558) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20844), .ZN(n20557) );
  OAI211_X1 U23494 ( .C1(n20847), .C2(n20591), .A(n20558), .B(n20557), .ZN(
        P1_U3102) );
  AOI22_X1 U23495 ( .A1(n20779), .A2(n20562), .B1(n20561), .B2(n20778), .ZN(
        n20560) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20851), .ZN(n20559) );
  OAI211_X1 U23497 ( .C1(n20854), .C2(n20591), .A(n20560), .B(n20559), .ZN(
        P1_U3103) );
  AOI22_X1 U23498 ( .A1(n20787), .A2(n20562), .B1(n20561), .B2(n20785), .ZN(
        n20566) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20860), .ZN(n20565) );
  OAI211_X1 U23500 ( .C1(n20866), .C2(n20591), .A(n20566), .B(n20565), .ZN(
        P1_U3104) );
  NOR2_X1 U23501 ( .A1(n20696), .A2(n20567), .ZN(n20586) );
  AOI21_X1 U23502 ( .B1(n20633), .B2(n20697), .A(n20586), .ZN(n20568) );
  OAI22_X1 U23503 ( .A1(n20568), .A2(n20706), .B1(n20567), .B2(n20870), .ZN(
        n20585) );
  AOI22_X1 U23504 ( .A1(n20733), .A2(n20586), .B1(n20585), .B2(n20732), .ZN(
        n20572) );
  OAI21_X1 U23505 ( .B1(n20637), .B2(n20704), .A(n20568), .ZN(n20569) );
  OAI221_X1 U23506 ( .B1(n20797), .B2(n20570), .C1(n20706), .C2(n20569), .A(
        n20806), .ZN(n20588) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20744), .ZN(n20571) );
  OAI211_X1 U23508 ( .C1(n20747), .C2(n20591), .A(n20572), .B(n20571), .ZN(
        P1_U3105) );
  AOI22_X1 U23509 ( .A1(n20749), .A2(n20586), .B1(n20585), .B2(n20748), .ZN(
        n20574) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20750), .ZN(n20573) );
  OAI211_X1 U23511 ( .C1(n20753), .C2(n20591), .A(n20574), .B(n20573), .ZN(
        P1_U3106) );
  AOI22_X1 U23512 ( .A1(n20755), .A2(n20586), .B1(n20585), .B2(n20754), .ZN(
        n20576) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20756), .ZN(n20575) );
  OAI211_X1 U23514 ( .C1(n20759), .C2(n20591), .A(n20576), .B(n20575), .ZN(
        P1_U3107) );
  AOI22_X1 U23515 ( .A1(n20761), .A2(n20586), .B1(n20585), .B2(n20760), .ZN(
        n20578) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20762), .ZN(n20577) );
  OAI211_X1 U23517 ( .C1(n20765), .C2(n20591), .A(n20578), .B(n20577), .ZN(
        P1_U3108) );
  AOI22_X1 U23518 ( .A1(n20767), .A2(n20586), .B1(n20585), .B2(n20766), .ZN(
        n20580) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20768), .ZN(n20579) );
  OAI211_X1 U23520 ( .C1(n20771), .C2(n20591), .A(n20580), .B(n20579), .ZN(
        P1_U3109) );
  AOI22_X1 U23521 ( .A1(n20773), .A2(n20586), .B1(n20585), .B2(n20772), .ZN(
        n20582) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20774), .ZN(n20581) );
  OAI211_X1 U23523 ( .C1(n20777), .C2(n20591), .A(n20582), .B(n20581), .ZN(
        P1_U3110) );
  AOI22_X1 U23524 ( .A1(n20779), .A2(n20586), .B1(n20585), .B2(n20778), .ZN(
        n20584) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20780), .ZN(n20583) );
  OAI211_X1 U23526 ( .C1(n20783), .C2(n20591), .A(n20584), .B(n20583), .ZN(
        P1_U3111) );
  AOI22_X1 U23527 ( .A1(n20787), .A2(n20586), .B1(n20585), .B2(n20785), .ZN(
        n20590) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20788), .ZN(n20589) );
  OAI211_X1 U23529 ( .C1(n20793), .C2(n20591), .A(n20590), .B(n20589), .ZN(
        P1_U3112) );
  NOR3_X1 U23530 ( .A1(n20662), .A2(n20592), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20639) );
  NAND2_X1 U23531 ( .A1(n20696), .A2(n20639), .ZN(n20623) );
  OAI22_X1 U23532 ( .A1(n20640), .A2(n20812), .B1(n20802), .B2(n20623), .ZN(
        n20593) );
  INV_X1 U23533 ( .A(n20593), .ZN(n20604) );
  AOI21_X1 U23534 ( .B1(n20640), .B2(n20629), .A(n20736), .ZN(n20594) );
  NOR2_X1 U23535 ( .A1(n20594), .A2(n20706), .ZN(n20599) );
  OR2_X1 U23536 ( .A1(n20595), .A2(n20667), .ZN(n20601) );
  AOI22_X1 U23537 ( .A1(n20599), .A2(n20601), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20623), .ZN(n20597) );
  OR2_X1 U23538 ( .A1(n20596), .A2(n20662), .ZN(n20730) );
  NAND2_X1 U23539 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20730), .ZN(n20741) );
  NAND3_X1 U23540 ( .A1(n20598), .A2(n20597), .A3(n20741), .ZN(n20626) );
  INV_X1 U23541 ( .A(n20599), .ZN(n20602) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20626), .B1(
        n20732), .B2(n20625), .ZN(n20603) );
  OAI211_X1 U23543 ( .C1(n20747), .C2(n20629), .A(n20604), .B(n20603), .ZN(
        P1_U3113) );
  OAI22_X1 U23544 ( .A1(n20640), .A2(n20819), .B1(n20814), .B2(n20623), .ZN(
        n20605) );
  INV_X1 U23545 ( .A(n20605), .ZN(n20607) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20626), .B1(
        n20748), .B2(n20625), .ZN(n20606) );
  OAI211_X1 U23547 ( .C1(n20753), .C2(n20629), .A(n20607), .B(n20606), .ZN(
        P1_U3114) );
  OAI22_X1 U23548 ( .A1(n20640), .A2(n20826), .B1(n20821), .B2(n20623), .ZN(
        n20608) );
  INV_X1 U23549 ( .A(n20608), .ZN(n20610) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20626), .B1(
        n20754), .B2(n20625), .ZN(n20609) );
  OAI211_X1 U23551 ( .C1(n20759), .C2(n20629), .A(n20610), .B(n20609), .ZN(
        P1_U3115) );
  OAI22_X1 U23552 ( .A1(n20629), .A2(n20765), .B1(n20828), .B2(n20623), .ZN(
        n20611) );
  INV_X1 U23553 ( .A(n20611), .ZN(n20613) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20626), .B1(
        n20760), .B2(n20625), .ZN(n20612) );
  OAI211_X1 U23555 ( .C1(n20833), .C2(n20640), .A(n20613), .B(n20612), .ZN(
        P1_U3116) );
  OAI22_X1 U23556 ( .A1(n20640), .A2(n20840), .B1(n20835), .B2(n20623), .ZN(
        n20614) );
  INV_X1 U23557 ( .A(n20614), .ZN(n20616) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20626), .B1(
        n20766), .B2(n20625), .ZN(n20615) );
  OAI211_X1 U23559 ( .C1(n20771), .C2(n20629), .A(n20616), .B(n20615), .ZN(
        P1_U3117) );
  OAI22_X1 U23560 ( .A1(n20640), .A2(n20847), .B1(n20842), .B2(n20623), .ZN(
        n20617) );
  INV_X1 U23561 ( .A(n20617), .ZN(n20619) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20626), .B1(
        n20772), .B2(n20625), .ZN(n20618) );
  OAI211_X1 U23563 ( .C1(n20777), .C2(n20629), .A(n20619), .B(n20618), .ZN(
        P1_U3118) );
  OAI22_X1 U23564 ( .A1(n20629), .A2(n20783), .B1(n20849), .B2(n20623), .ZN(
        n20620) );
  INV_X1 U23565 ( .A(n20620), .ZN(n20622) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20626), .B1(
        n20778), .B2(n20625), .ZN(n20621) );
  OAI211_X1 U23567 ( .C1(n20854), .C2(n20640), .A(n20622), .B(n20621), .ZN(
        P1_U3119) );
  OAI22_X1 U23568 ( .A1(n20640), .A2(n20866), .B1(n20858), .B2(n20623), .ZN(
        n20624) );
  INV_X1 U23569 ( .A(n20624), .ZN(n20628) );
  AOI22_X1 U23570 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20626), .B1(
        n20785), .B2(n20625), .ZN(n20627) );
  OAI211_X1 U23571 ( .C1(n20793), .C2(n20629), .A(n20628), .B(n20627), .ZN(
        P1_U3120) );
  NOR2_X1 U23572 ( .A1(n20632), .A2(n20662), .ZN(n20656) );
  AOI21_X1 U23573 ( .B1(n20633), .B2(n20794), .A(n20656), .ZN(n20635) );
  INV_X1 U23574 ( .A(n20639), .ZN(n20634) );
  OAI22_X1 U23575 ( .A1(n20635), .A2(n20706), .B1(n20634), .B2(n20870), .ZN(
        n20655) );
  AOI22_X1 U23576 ( .A1(n20733), .A2(n20656), .B1(n20655), .B2(n20732), .ZN(
        n20642) );
  OAI21_X1 U23577 ( .B1(n20637), .B2(n20636), .A(n20635), .ZN(n20638) );
  OAI221_X1 U23578 ( .B1(n20797), .B2(n20639), .C1(n20706), .C2(n20638), .A(
        n20806), .ZN(n20658) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20809), .ZN(n20641) );
  OAI211_X1 U23580 ( .C1(n20812), .C2(n20693), .A(n20642), .B(n20641), .ZN(
        P1_U3121) );
  AOI22_X1 U23581 ( .A1(n20749), .A2(n20656), .B1(n20655), .B2(n20748), .ZN(
        n20644) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20816), .ZN(n20643) );
  OAI211_X1 U23583 ( .C1(n20819), .C2(n20693), .A(n20644), .B(n20643), .ZN(
        P1_U3122) );
  AOI22_X1 U23584 ( .A1(n20755), .A2(n20656), .B1(n20655), .B2(n20754), .ZN(
        n20646) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20823), .ZN(n20645) );
  OAI211_X1 U23586 ( .C1(n20826), .C2(n20693), .A(n20646), .B(n20645), .ZN(
        P1_U3123) );
  AOI22_X1 U23587 ( .A1(n20761), .A2(n20656), .B1(n20655), .B2(n20760), .ZN(
        n20648) );
  AOI22_X1 U23588 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20830), .ZN(n20647) );
  OAI211_X1 U23589 ( .C1(n20833), .C2(n20693), .A(n20648), .B(n20647), .ZN(
        P1_U3124) );
  AOI22_X1 U23590 ( .A1(n20767), .A2(n20656), .B1(n20655), .B2(n20766), .ZN(
        n20650) );
  AOI22_X1 U23591 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20837), .ZN(n20649) );
  OAI211_X1 U23592 ( .C1(n20840), .C2(n20693), .A(n20650), .B(n20649), .ZN(
        P1_U3125) );
  AOI22_X1 U23593 ( .A1(n20773), .A2(n20656), .B1(n20655), .B2(n20772), .ZN(
        n20652) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20844), .ZN(n20651) );
  OAI211_X1 U23595 ( .C1(n20847), .C2(n20693), .A(n20652), .B(n20651), .ZN(
        P1_U3126) );
  AOI22_X1 U23596 ( .A1(n20779), .A2(n20656), .B1(n20655), .B2(n20778), .ZN(
        n20654) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20851), .ZN(n20653) );
  OAI211_X1 U23598 ( .C1(n20854), .C2(n20693), .A(n20654), .B(n20653), .ZN(
        P1_U3127) );
  AOI22_X1 U23599 ( .A1(n20787), .A2(n20656), .B1(n20655), .B2(n20785), .ZN(
        n20660) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20860), .ZN(n20659) );
  OAI211_X1 U23601 ( .C1(n20866), .C2(n20693), .A(n20660), .B(n20659), .ZN(
        P1_U3128) );
  NOR3_X1 U23602 ( .A1(n20663), .A2(n20662), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20707) );
  INV_X1 U23603 ( .A(n20707), .ZN(n20695) );
  NOR2_X1 U23604 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20695), .ZN(
        n20688) );
  AOI22_X1 U23605 ( .A1(n20724), .A2(n20744), .B1(n20733), .B2(n20688), .ZN(
        n20675) );
  INV_X1 U23606 ( .A(n20724), .ZN(n20664) );
  AOI21_X1 U23607 ( .B1(n20664), .B2(n20693), .A(n20736), .ZN(n20665) );
  NOR2_X1 U23608 ( .A1(n20665), .A2(n20706), .ZN(n20670) );
  NOR2_X1 U23609 ( .A1(n13162), .A2(n20666), .ZN(n20795) );
  NAND2_X1 U23610 ( .A1(n20795), .A2(n20667), .ZN(n20672) );
  AOI22_X1 U23611 ( .A1(n20670), .A2(n20672), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20671), .ZN(n20668) );
  INV_X1 U23612 ( .A(n20670), .ZN(n20673) );
  AOI22_X1 U23613 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20690), .B1(
        n20732), .B2(n20689), .ZN(n20674) );
  OAI211_X1 U23614 ( .C1(n20747), .C2(n20693), .A(n20675), .B(n20674), .ZN(
        P1_U3129) );
  AOI22_X1 U23615 ( .A1(n20724), .A2(n20750), .B1(n20749), .B2(n20688), .ZN(
        n20677) );
  AOI22_X1 U23616 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20690), .B1(
        n20748), .B2(n20689), .ZN(n20676) );
  OAI211_X1 U23617 ( .C1(n20753), .C2(n20693), .A(n20677), .B(n20676), .ZN(
        P1_U3130) );
  AOI22_X1 U23618 ( .A1(n20724), .A2(n20756), .B1(n20755), .B2(n20688), .ZN(
        n20679) );
  AOI22_X1 U23619 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20690), .B1(
        n20754), .B2(n20689), .ZN(n20678) );
  OAI211_X1 U23620 ( .C1(n20759), .C2(n20693), .A(n20679), .B(n20678), .ZN(
        P1_U3131) );
  AOI22_X1 U23621 ( .A1(n20724), .A2(n20762), .B1(n20761), .B2(n20688), .ZN(
        n20681) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20690), .B1(
        n20760), .B2(n20689), .ZN(n20680) );
  OAI211_X1 U23623 ( .C1(n20765), .C2(n20693), .A(n20681), .B(n20680), .ZN(
        P1_U3132) );
  AOI22_X1 U23624 ( .A1(n20724), .A2(n20768), .B1(n20767), .B2(n20688), .ZN(
        n20683) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20690), .B1(
        n20766), .B2(n20689), .ZN(n20682) );
  OAI211_X1 U23626 ( .C1(n20771), .C2(n20693), .A(n20683), .B(n20682), .ZN(
        P1_U3133) );
  AOI22_X1 U23627 ( .A1(n20724), .A2(n20774), .B1(n20773), .B2(n20688), .ZN(
        n20685) );
  AOI22_X1 U23628 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20690), .B1(
        n20772), .B2(n20689), .ZN(n20684) );
  OAI211_X1 U23629 ( .C1(n20777), .C2(n20693), .A(n20685), .B(n20684), .ZN(
        P1_U3134) );
  AOI22_X1 U23630 ( .A1(n20724), .A2(n20780), .B1(n20779), .B2(n20688), .ZN(
        n20687) );
  AOI22_X1 U23631 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20690), .B1(
        n20778), .B2(n20689), .ZN(n20686) );
  OAI211_X1 U23632 ( .C1(n20783), .C2(n20693), .A(n20687), .B(n20686), .ZN(
        P1_U3135) );
  AOI22_X1 U23633 ( .A1(n20724), .A2(n20788), .B1(n20787), .B2(n20688), .ZN(
        n20692) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20690), .B1(
        n20785), .B2(n20689), .ZN(n20691) );
  OAI211_X1 U23635 ( .C1(n20793), .C2(n20693), .A(n20692), .B(n20691), .ZN(
        P1_U3136) );
  NOR2_X1 U23636 ( .A1(n20696), .A2(n20695), .ZN(n20723) );
  NAND2_X1 U23637 ( .A1(n20795), .A2(n20697), .ZN(n20699) );
  INV_X1 U23638 ( .A(n20723), .ZN(n20698) );
  NAND2_X1 U23639 ( .A1(n20699), .A2(n20698), .ZN(n20702) );
  NAND2_X1 U23640 ( .A1(n20702), .A2(n20797), .ZN(n20701) );
  NAND2_X1 U23641 ( .A1(n20707), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20700) );
  NAND2_X1 U23642 ( .A1(n20701), .A2(n20700), .ZN(n20722) );
  AOI22_X1 U23643 ( .A1(n20733), .A2(n20723), .B1(n20732), .B2(n20722), .ZN(
        n20709) );
  INV_X1 U23644 ( .A(n20735), .ZN(n20805) );
  INV_X1 U23645 ( .A(n20702), .ZN(n20703) );
  OAI21_X1 U23646 ( .B1(n20805), .B2(n20704), .A(n20703), .ZN(n20705) );
  OAI221_X1 U23647 ( .B1(n20797), .B2(n20707), .C1(n20706), .C2(n20705), .A(
        n20806), .ZN(n20725) );
  AOI22_X1 U23648 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20809), .ZN(n20708) );
  OAI211_X1 U23649 ( .C1(n20812), .C2(n20792), .A(n20709), .B(n20708), .ZN(
        P1_U3137) );
  AOI22_X1 U23650 ( .A1(n20749), .A2(n20723), .B1(n20748), .B2(n20722), .ZN(
        n20711) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20816), .ZN(n20710) );
  OAI211_X1 U23652 ( .C1(n20819), .C2(n20792), .A(n20711), .B(n20710), .ZN(
        P1_U3138) );
  AOI22_X1 U23653 ( .A1(n20755), .A2(n20723), .B1(n20754), .B2(n20722), .ZN(
        n20713) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20823), .ZN(n20712) );
  OAI211_X1 U23655 ( .C1(n20826), .C2(n20792), .A(n20713), .B(n20712), .ZN(
        P1_U3139) );
  AOI22_X1 U23656 ( .A1(n20761), .A2(n20723), .B1(n20760), .B2(n20722), .ZN(
        n20715) );
  AOI22_X1 U23657 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20830), .ZN(n20714) );
  OAI211_X1 U23658 ( .C1(n20833), .C2(n20792), .A(n20715), .B(n20714), .ZN(
        P1_U3140) );
  AOI22_X1 U23659 ( .A1(n20767), .A2(n20723), .B1(n20766), .B2(n20722), .ZN(
        n20717) );
  AOI22_X1 U23660 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20837), .ZN(n20716) );
  OAI211_X1 U23661 ( .C1(n20840), .C2(n20792), .A(n20717), .B(n20716), .ZN(
        P1_U3141) );
  AOI22_X1 U23662 ( .A1(n20773), .A2(n20723), .B1(n20772), .B2(n20722), .ZN(
        n20719) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20844), .ZN(n20718) );
  OAI211_X1 U23664 ( .C1(n20847), .C2(n20792), .A(n20719), .B(n20718), .ZN(
        P1_U3142) );
  AOI22_X1 U23665 ( .A1(n20779), .A2(n20723), .B1(n20778), .B2(n20722), .ZN(
        n20721) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20851), .ZN(n20720) );
  OAI211_X1 U23667 ( .C1(n20854), .C2(n20792), .A(n20721), .B(n20720), .ZN(
        P1_U3143) );
  AOI22_X1 U23668 ( .A1(n20787), .A2(n20723), .B1(n20785), .B2(n20722), .ZN(
        n20727) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20860), .ZN(n20726) );
  OAI211_X1 U23670 ( .C1(n20866), .C2(n20792), .A(n20727), .B(n20726), .ZN(
        P1_U3144) );
  INV_X1 U23671 ( .A(n20807), .ZN(n20728) );
  NOR2_X1 U23672 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20728), .ZN(
        n20786) );
  NAND3_X1 U23673 ( .A1(n20795), .A2(n20739), .A3(n20797), .ZN(n20729) );
  OAI21_X1 U23674 ( .B1(n20731), .B2(n20730), .A(n20729), .ZN(n20784) );
  AOI22_X1 U23675 ( .A1(n20733), .A2(n20786), .B1(n20732), .B2(n20784), .ZN(
        n20746) );
  INV_X1 U23676 ( .A(n20861), .ZN(n20737) );
  AOI21_X1 U23677 ( .B1(n20737), .B2(n20792), .A(n20736), .ZN(n20738) );
  AOI21_X1 U23678 ( .B1(n20795), .B2(n20739), .A(n20738), .ZN(n20740) );
  NOR2_X1 U23679 ( .A1(n20740), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20743) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20789), .B1(
        n20861), .B2(n20744), .ZN(n20745) );
  OAI211_X1 U23681 ( .C1(n20747), .C2(n20792), .A(n20746), .B(n20745), .ZN(
        P1_U3145) );
  AOI22_X1 U23682 ( .A1(n20749), .A2(n20786), .B1(n20748), .B2(n20784), .ZN(
        n20752) );
  AOI22_X1 U23683 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20789), .B1(
        n20861), .B2(n20750), .ZN(n20751) );
  OAI211_X1 U23684 ( .C1(n20753), .C2(n20792), .A(n20752), .B(n20751), .ZN(
        P1_U3146) );
  AOI22_X1 U23685 ( .A1(n20755), .A2(n20786), .B1(n20754), .B2(n20784), .ZN(
        n20758) );
  AOI22_X1 U23686 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20789), .B1(
        n20861), .B2(n20756), .ZN(n20757) );
  OAI211_X1 U23687 ( .C1(n20759), .C2(n20792), .A(n20758), .B(n20757), .ZN(
        P1_U3147) );
  AOI22_X1 U23688 ( .A1(n20761), .A2(n20786), .B1(n20760), .B2(n20784), .ZN(
        n20764) );
  AOI22_X1 U23689 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20789), .B1(
        n20861), .B2(n20762), .ZN(n20763) );
  OAI211_X1 U23690 ( .C1(n20765), .C2(n20792), .A(n20764), .B(n20763), .ZN(
        P1_U3148) );
  AOI22_X1 U23691 ( .A1(n20767), .A2(n20786), .B1(n20766), .B2(n20784), .ZN(
        n20770) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20789), .B1(
        n20861), .B2(n20768), .ZN(n20769) );
  OAI211_X1 U23693 ( .C1(n20771), .C2(n20792), .A(n20770), .B(n20769), .ZN(
        P1_U3149) );
  AOI22_X1 U23694 ( .A1(n20773), .A2(n20786), .B1(n20772), .B2(n20784), .ZN(
        n20776) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20789), .B1(
        n20861), .B2(n20774), .ZN(n20775) );
  OAI211_X1 U23696 ( .C1(n20777), .C2(n20792), .A(n20776), .B(n20775), .ZN(
        P1_U3150) );
  AOI22_X1 U23697 ( .A1(n20779), .A2(n20786), .B1(n20778), .B2(n20784), .ZN(
        n20782) );
  AOI22_X1 U23698 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20789), .B1(
        n20861), .B2(n20780), .ZN(n20781) );
  OAI211_X1 U23699 ( .C1(n20783), .C2(n20792), .A(n20782), .B(n20781), .ZN(
        P1_U3151) );
  AOI22_X1 U23700 ( .A1(n20787), .A2(n20786), .B1(n20785), .B2(n20784), .ZN(
        n20791) );
  AOI22_X1 U23701 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20789), .B1(
        n20861), .B2(n20788), .ZN(n20790) );
  OAI211_X1 U23702 ( .C1(n20793), .C2(n20792), .A(n20791), .B(n20790), .ZN(
        P1_U3152) );
  NAND2_X1 U23703 ( .A1(n20795), .A2(n20794), .ZN(n20796) );
  NAND2_X1 U23704 ( .A1(n20796), .A2(n20857), .ZN(n20798) );
  NAND2_X1 U23705 ( .A1(n20798), .A2(n20797), .ZN(n20800) );
  NAND2_X1 U23706 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20807), .ZN(n20799) );
  AND2_X1 U23707 ( .A1(n20800), .A2(n20799), .ZN(n20856) );
  OAI22_X1 U23708 ( .A1(n20802), .A2(n20857), .B1(n20856), .B2(n20801), .ZN(
        n20803) );
  INV_X1 U23709 ( .A(n20803), .ZN(n20811) );
  NOR2_X1 U23710 ( .A1(n20805), .A2(n20804), .ZN(n20808) );
  OAI21_X1 U23711 ( .B1(n20808), .B2(n20807), .A(n20806), .ZN(n20862) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20862), .B1(
        n20861), .B2(n20809), .ZN(n20810) );
  OAI211_X1 U23713 ( .C1(n20812), .C2(n20865), .A(n20811), .B(n20810), .ZN(
        P1_U3153) );
  OAI22_X1 U23714 ( .A1(n20814), .A2(n20857), .B1(n20856), .B2(n20813), .ZN(
        n20815) );
  INV_X1 U23715 ( .A(n20815), .ZN(n20818) );
  AOI22_X1 U23716 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20862), .B1(
        n20861), .B2(n20816), .ZN(n20817) );
  OAI211_X1 U23717 ( .C1(n20819), .C2(n20865), .A(n20818), .B(n20817), .ZN(
        P1_U3154) );
  OAI22_X1 U23718 ( .A1(n20821), .A2(n20857), .B1(n20856), .B2(n20820), .ZN(
        n20822) );
  INV_X1 U23719 ( .A(n20822), .ZN(n20825) );
  AOI22_X1 U23720 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20862), .B1(
        n20861), .B2(n20823), .ZN(n20824) );
  OAI211_X1 U23721 ( .C1(n20826), .C2(n20865), .A(n20825), .B(n20824), .ZN(
        P1_U3155) );
  OAI22_X1 U23722 ( .A1(n20828), .A2(n20857), .B1(n20856), .B2(n20827), .ZN(
        n20829) );
  INV_X1 U23723 ( .A(n20829), .ZN(n20832) );
  AOI22_X1 U23724 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20862), .B1(
        n20861), .B2(n20830), .ZN(n20831) );
  OAI211_X1 U23725 ( .C1(n20833), .C2(n20865), .A(n20832), .B(n20831), .ZN(
        P1_U3156) );
  OAI22_X1 U23726 ( .A1(n20835), .A2(n20857), .B1(n20856), .B2(n20834), .ZN(
        n20836) );
  INV_X1 U23727 ( .A(n20836), .ZN(n20839) );
  AOI22_X1 U23728 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20862), .B1(
        n20861), .B2(n20837), .ZN(n20838) );
  OAI211_X1 U23729 ( .C1(n20840), .C2(n20865), .A(n20839), .B(n20838), .ZN(
        P1_U3157) );
  OAI22_X1 U23730 ( .A1(n20842), .A2(n20857), .B1(n20856), .B2(n20841), .ZN(
        n20843) );
  INV_X1 U23731 ( .A(n20843), .ZN(n20846) );
  AOI22_X1 U23732 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20862), .B1(
        n20861), .B2(n20844), .ZN(n20845) );
  OAI211_X1 U23733 ( .C1(n20847), .C2(n20865), .A(n20846), .B(n20845), .ZN(
        P1_U3158) );
  OAI22_X1 U23734 ( .A1(n20849), .A2(n20857), .B1(n20856), .B2(n20848), .ZN(
        n20850) );
  INV_X1 U23735 ( .A(n20850), .ZN(n20853) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20862), .B1(
        n20861), .B2(n20851), .ZN(n20852) );
  OAI211_X1 U23737 ( .C1(n20854), .C2(n20865), .A(n20853), .B(n20852), .ZN(
        P1_U3159) );
  OAI22_X1 U23738 ( .A1(n20858), .A2(n20857), .B1(n20856), .B2(n20855), .ZN(
        n20859) );
  INV_X1 U23739 ( .A(n20859), .ZN(n20864) );
  AOI22_X1 U23740 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20862), .B1(
        n20861), .B2(n20860), .ZN(n20863) );
  OAI211_X1 U23741 ( .C1(n20866), .C2(n20865), .A(n20864), .B(n20863), .ZN(
        P1_U3160) );
  NOR2_X1 U23742 ( .A1(n20868), .A2(n20867), .ZN(n20871) );
  OAI21_X1 U23743 ( .B1(n20871), .B2(n20870), .A(n20869), .ZN(P1_U3163) );
  AND2_X1 U23744 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20872), .ZN(
        P1_U3164) );
  AND2_X1 U23745 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20872), .ZN(
        P1_U3165) );
  AND2_X1 U23746 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20872), .ZN(
        P1_U3166) );
  AND2_X1 U23747 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20872), .ZN(
        P1_U3167) );
  AND2_X1 U23748 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20872), .ZN(
        P1_U3168) );
  AND2_X1 U23749 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20872), .ZN(
        P1_U3169) );
  AND2_X1 U23750 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20872), .ZN(
        P1_U3170) );
  AND2_X1 U23751 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20872), .ZN(
        P1_U3171) );
  AND2_X1 U23752 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20872), .ZN(
        P1_U3172) );
  AND2_X1 U23753 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20872), .ZN(
        P1_U3173) );
  AND2_X1 U23754 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20872), .ZN(
        P1_U3174) );
  AND2_X1 U23755 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20872), .ZN(
        P1_U3175) );
  AND2_X1 U23756 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20872), .ZN(
        P1_U3176) );
  AND2_X1 U23757 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20872), .ZN(
        P1_U3177) );
  AND2_X1 U23758 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20872), .ZN(
        P1_U3178) );
  AND2_X1 U23759 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20872), .ZN(
        P1_U3179) );
  AND2_X1 U23760 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20872), .ZN(
        P1_U3180) );
  AND2_X1 U23761 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20872), .ZN(
        P1_U3181) );
  AND2_X1 U23762 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20872), .ZN(
        P1_U3182) );
  AND2_X1 U23763 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20872), .ZN(
        P1_U3183) );
  AND2_X1 U23764 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20872), .ZN(
        P1_U3184) );
  AND2_X1 U23765 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20872), .ZN(
        P1_U3185) );
  AND2_X1 U23766 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20872), .ZN(P1_U3186) );
  AND2_X1 U23767 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20872), .ZN(P1_U3187) );
  AND2_X1 U23768 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20872), .ZN(P1_U3188) );
  AND2_X1 U23769 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20872), .ZN(P1_U3189) );
  AND2_X1 U23770 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20872), .ZN(P1_U3190) );
  AND2_X1 U23771 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20872), .ZN(P1_U3191) );
  AND2_X1 U23772 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20872), .ZN(P1_U3192) );
  AND2_X1 U23773 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20872), .ZN(P1_U3193) );
  INV_X1 U23774 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20879) );
  NOR2_X1 U23775 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20874) );
  OAI22_X1 U23776 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20883), .B1(n20874), 
        .B2(n20873), .ZN(n20875) );
  OAI21_X1 U23777 ( .B1(n20879), .B2(n20875), .A(n20960), .ZN(n20876) );
  OAI211_X1 U23778 ( .C1(n20878), .C2(n20951), .A(n20877), .B(n20876), .ZN(
        P1_U3194) );
  OAI221_X1 U23779 ( .B1(n20878), .B2(n20881), .C1(n20878), .C2(n20883), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n20888) );
  OAI21_X1 U23780 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20879), .A(HOLD), .ZN(
        n20887) );
  NOR2_X1 U23781 ( .A1(NA), .A2(n20884), .ZN(n20880) );
  AOI21_X1 U23782 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20880), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n20886) );
  AND2_X1 U23783 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20881), .ZN(n20882) );
  AOI221_X1 U23784 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20884), .C1(n20883), 
        .C2(n20884), .A(n20882), .ZN(n20885) );
  OAI22_X1 U23785 ( .A1(n20888), .A2(n20887), .B1(n20886), .B2(n20885), .ZN(
        P1_U3196) );
  OR2_X1 U23786 ( .A1(n20960), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20923) );
  OR2_X1 U23787 ( .A1(n20889), .A2(n20960), .ZN(n20920) );
  INV_X1 U23788 ( .A(n20920), .ZN(n20928) );
  AOI222_X1 U23789 ( .A1(n9647), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20928), .ZN(n20890) );
  INV_X1 U23790 ( .A(n20890), .ZN(P1_U3197) );
  AOI22_X1 U23791 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20960), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n9647), .ZN(n20891) );
  OAI21_X1 U23792 ( .B1(n20892), .B2(n20920), .A(n20891), .ZN(P1_U3198) );
  AOI222_X1 U23793 ( .A1(n20928), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n9647), .ZN(n20893) );
  INV_X1 U23794 ( .A(n20893), .ZN(P1_U3199) );
  AOI222_X1 U23795 ( .A1(n9647), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20928), .ZN(n20894) );
  INV_X1 U23796 ( .A(n20894), .ZN(P1_U3200) );
  AOI22_X1 U23797 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20960), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n9647), .ZN(n20895) );
  OAI21_X1 U23798 ( .B1(n20896), .B2(n20920), .A(n20895), .ZN(P1_U3201) );
  AOI22_X1 U23799 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20960), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20928), .ZN(n20897) );
  OAI21_X1 U23800 ( .B1(n20898), .B2(n20923), .A(n20897), .ZN(P1_U3202) );
  AOI222_X1 U23801 ( .A1(n20928), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n9647), .ZN(n20899) );
  INV_X1 U23802 ( .A(n20899), .ZN(P1_U3203) );
  AOI222_X1 U23803 ( .A1(n9647), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20960), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20928), .ZN(n20900) );
  INV_X1 U23804 ( .A(n20900), .ZN(P1_U3204) );
  AOI222_X1 U23805 ( .A1(n20928), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n9647), .ZN(n20901) );
  INV_X1 U23806 ( .A(n20901), .ZN(P1_U3205) );
  AOI222_X1 U23807 ( .A1(n20928), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n9647), .ZN(n20902) );
  INV_X1 U23808 ( .A(n20902), .ZN(P1_U3206) );
  AOI222_X1 U23809 ( .A1(n20928), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n9647), .ZN(n20903) );
  INV_X1 U23810 ( .A(n20903), .ZN(P1_U3207) );
  AOI222_X1 U23811 ( .A1(n20928), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n9647), .ZN(n20904) );
  INV_X1 U23812 ( .A(n20904), .ZN(P1_U3208) );
  AOI222_X1 U23813 ( .A1(n20928), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n9647), .ZN(n20905) );
  INV_X1 U23814 ( .A(n20905), .ZN(P1_U3209) );
  AOI222_X1 U23815 ( .A1(n9647), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20928), .ZN(n20906) );
  INV_X1 U23816 ( .A(n20906), .ZN(P1_U3210) );
  AOI222_X1 U23817 ( .A1(n9647), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20928), .ZN(n20907) );
  INV_X1 U23818 ( .A(n20907), .ZN(P1_U3211) );
  AOI22_X1 U23819 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20960), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n9647), .ZN(n20908) );
  OAI21_X1 U23820 ( .B1(n14577), .B2(n20920), .A(n20908), .ZN(P1_U3212) );
  AOI22_X1 U23821 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20960), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20928), .ZN(n20909) );
  OAI21_X1 U23822 ( .B1(n14563), .B2(n20923), .A(n20909), .ZN(P1_U3213) );
  AOI222_X1 U23823 ( .A1(n20928), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n9647), .ZN(n20910) );
  INV_X1 U23824 ( .A(n20910), .ZN(P1_U3214) );
  AOI222_X1 U23825 ( .A1(n9647), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20928), .ZN(n20911) );
  INV_X1 U23826 ( .A(n20911), .ZN(P1_U3215) );
  AOI222_X1 U23827 ( .A1(n20928), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n9647), .ZN(n20912) );
  INV_X1 U23828 ( .A(n20912), .ZN(P1_U3216) );
  AOI22_X1 U23829 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20960), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n9647), .ZN(n20913) );
  OAI21_X1 U23830 ( .B1(n20914), .B2(n20920), .A(n20913), .ZN(P1_U3217) );
  AOI22_X1 U23831 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20960), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20928), .ZN(n20915) );
  OAI21_X1 U23832 ( .B1(n20916), .B2(n20923), .A(n20915), .ZN(P1_U3218) );
  AOI222_X1 U23833 ( .A1(n20928), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n9647), .ZN(n20917) );
  INV_X1 U23834 ( .A(n20917), .ZN(P1_U3219) );
  AOI222_X1 U23835 ( .A1(n20928), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n9647), .ZN(n20918) );
  INV_X1 U23836 ( .A(n20918), .ZN(P1_U3220) );
  AOI22_X1 U23837 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n9647), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20932), .ZN(n20919) );
  OAI21_X1 U23838 ( .B1(n20921), .B2(n20920), .A(n20919), .ZN(P1_U3221) );
  AOI22_X1 U23839 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20928), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20932), .ZN(n20922) );
  OAI21_X1 U23840 ( .B1(n20924), .B2(n20923), .A(n20922), .ZN(P1_U3222) );
  AOI222_X1 U23841 ( .A1(n9647), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20928), .ZN(n20925) );
  INV_X1 U23842 ( .A(n20925), .ZN(P1_U3223) );
  AOI222_X1 U23843 ( .A1(n20928), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n9647), .ZN(n20926) );
  INV_X1 U23844 ( .A(n20926), .ZN(P1_U3224) );
  AOI222_X1 U23845 ( .A1(n9647), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20928), .ZN(n20927) );
  INV_X1 U23846 ( .A(n20927), .ZN(P1_U3225) );
  AOI222_X1 U23847 ( .A1(n20928), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20932), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n9647), .ZN(n20929) );
  INV_X1 U23848 ( .A(n20929), .ZN(P1_U3226) );
  OAI22_X1 U23849 ( .A1(n20960), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20948), .ZN(n20930) );
  INV_X1 U23850 ( .A(n20930), .ZN(P1_U3458) );
  OAI22_X1 U23851 ( .A1(n20960), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20948), .ZN(n20931) );
  INV_X1 U23852 ( .A(n20931), .ZN(P1_U3459) );
  OAI22_X1 U23853 ( .A1(n20932), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20948), .ZN(n20933) );
  INV_X1 U23854 ( .A(n20933), .ZN(P1_U3460) );
  OAI22_X1 U23855 ( .A1(n20960), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20948), .ZN(n20934) );
  INV_X1 U23856 ( .A(n20934), .ZN(P1_U3461) );
  OAI21_X1 U23857 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20938), .A(n20936), 
        .ZN(n20935) );
  INV_X1 U23858 ( .A(n20935), .ZN(P1_U3464) );
  OAI21_X1 U23859 ( .B1(n20938), .B2(n20937), .A(n20936), .ZN(P1_U3465) );
  AOI21_X1 U23860 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20940) );
  AOI22_X1 U23861 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20940), .B2(n20939), .ZN(n20943) );
  INV_X1 U23862 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20942) );
  AOI22_X1 U23863 ( .A1(n20946), .A2(n20943), .B1(n20942), .B2(n20941), .ZN(
        P1_U3481) );
  INV_X1 U23864 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20945) );
  OAI21_X1 U23865 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20946), .ZN(n20944) );
  OAI21_X1 U23866 ( .B1(n20946), .B2(n20945), .A(n20944), .ZN(P1_U3482) );
  AOI22_X1 U23867 ( .A1(n20948), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20947), 
        .B2(n20960), .ZN(P1_U3483) );
  AOI211_X1 U23868 ( .C1(n20185), .C2(n20951), .A(n20950), .B(n20949), .ZN(
        n20959) );
  INV_X1 U23869 ( .A(n20952), .ZN(n20953) );
  OAI211_X1 U23870 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20954), .A(n20953), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20956) );
  AOI21_X1 U23871 ( .B1(n20956), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20955), 
        .ZN(n20958) );
  NAND2_X1 U23872 ( .A1(n20959), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20957) );
  OAI21_X1 U23873 ( .B1(n20959), .B2(n20958), .A(n20957), .ZN(P1_U3485) );
  MUX2_X1 U23874 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20960), .Z(P1_U3486) );
  INV_X1 U23875 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n21103) );
  AOI22_X1 U23876 ( .A1(n21103), .A2(keyinput87), .B1(keyinput90), .B2(n21109), 
        .ZN(n20961) );
  OAI221_X1 U23877 ( .B1(n21103), .B2(keyinput87), .C1(n21109), .C2(keyinput90), .A(n20961), .ZN(n20971) );
  INV_X1 U23878 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n20963) );
  AOI22_X1 U23879 ( .A1(n20963), .A2(keyinput95), .B1(n21128), .B2(keyinput117), .ZN(n20962) );
  OAI221_X1 U23880 ( .B1(n20963), .B2(keyinput95), .C1(n21128), .C2(
        keyinput117), .A(n20962), .ZN(n20970) );
  INV_X1 U23881 ( .A(DATAI_2_), .ZN(n21099) );
  AOI22_X1 U23882 ( .A1(n21099), .A2(keyinput78), .B1(n20965), .B2(keyinput124), .ZN(n20964) );
  OAI221_X1 U23883 ( .B1(n21099), .B2(keyinput78), .C1(n20965), .C2(
        keyinput124), .A(n20964), .ZN(n20969) );
  INV_X1 U23884 ( .A(P3_UWORD_REG_4__SCAN_IN), .ZN(n20967) );
  AOI22_X1 U23885 ( .A1(n11164), .A2(keyinput106), .B1(keyinput72), .B2(n20967), .ZN(n20966) );
  OAI221_X1 U23886 ( .B1(n11164), .B2(keyinput106), .C1(n20967), .C2(
        keyinput72), .A(n20966), .ZN(n20968) );
  NOR4_X1 U23887 ( .A1(n20971), .A2(n20970), .A3(n20969), .A4(n20968), .ZN(
        n21006) );
  AOI22_X1 U23888 ( .A1(n21123), .A2(keyinput80), .B1(n11811), .B2(keyinput77), 
        .ZN(n20972) );
  OAI221_X1 U23889 ( .B1(n21123), .B2(keyinput80), .C1(n11811), .C2(keyinput77), .A(n20972), .ZN(n20980) );
  AOI22_X1 U23890 ( .A1(BUF1_REG_28__SCAN_IN), .A2(keyinput103), .B1(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .B2(keyinput86), .ZN(n20973) );
  OAI221_X1 U23891 ( .B1(BUF1_REG_28__SCAN_IN), .B2(keyinput103), .C1(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .C2(keyinput86), .A(n20973), .ZN(
        n20979) );
  AOI22_X1 U23892 ( .A1(n21094), .A2(keyinput102), .B1(keyinput91), .B2(n20975), .ZN(n20974) );
  OAI221_X1 U23893 ( .B1(n21094), .B2(keyinput102), .C1(n20975), .C2(
        keyinput91), .A(n20974), .ZN(n20978) );
  AOI22_X1 U23894 ( .A1(n21115), .A2(keyinput121), .B1(keyinput120), .B2(
        n11641), .ZN(n20976) );
  OAI221_X1 U23895 ( .B1(n21115), .B2(keyinput121), .C1(n11641), .C2(
        keyinput120), .A(n20976), .ZN(n20977) );
  NOR4_X1 U23896 ( .A1(n20980), .A2(n20979), .A3(n20978), .A4(n20977), .ZN(
        n21005) );
  AOI22_X1 U23897 ( .A1(n20982), .A2(keyinput92), .B1(keyinput116), .B2(n18253), .ZN(n20981) );
  OAI221_X1 U23898 ( .B1(n20982), .B2(keyinput92), .C1(n18253), .C2(
        keyinput116), .A(n20981), .ZN(n20992) );
  AOI22_X1 U23899 ( .A1(n11846), .A2(keyinput79), .B1(n20984), .B2(keyinput126), .ZN(n20983) );
  OAI221_X1 U23900 ( .B1(n11846), .B2(keyinput79), .C1(n20984), .C2(
        keyinput126), .A(n20983), .ZN(n20991) );
  AOI22_X1 U23901 ( .A1(n21132), .A2(keyinput127), .B1(n20986), .B2(keyinput84), .ZN(n20985) );
  OAI221_X1 U23902 ( .B1(n21132), .B2(keyinput127), .C1(n20986), .C2(
        keyinput84), .A(n20985), .ZN(n20990) );
  XNOR2_X1 U23903 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B(keyinput74), .ZN(
        n20988) );
  XNOR2_X1 U23904 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput73), .ZN(n20987) );
  NAND2_X1 U23905 ( .A1(n20988), .A2(n20987), .ZN(n20989) );
  NOR4_X1 U23906 ( .A1(n20992), .A2(n20991), .A3(n20990), .A4(n20989), .ZN(
        n21004) );
  INV_X1 U23907 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n21080) );
  AOI22_X1 U23908 ( .A1(n21080), .A2(keyinput109), .B1(keyinput125), .B2(
        n20994), .ZN(n20993) );
  OAI221_X1 U23909 ( .B1(n21080), .B2(keyinput109), .C1(n20994), .C2(
        keyinput125), .A(n20993), .ZN(n21002) );
  AOI22_X1 U23910 ( .A1(n21096), .A2(keyinput75), .B1(n11626), .B2(keyinput70), 
        .ZN(n20995) );
  OAI221_X1 U23911 ( .B1(n21096), .B2(keyinput75), .C1(n11626), .C2(keyinput70), .A(n20995), .ZN(n21001) );
  AOI22_X1 U23912 ( .A1(n21118), .A2(keyinput98), .B1(keyinput107), .B2(n21129), .ZN(n20996) );
  OAI221_X1 U23913 ( .B1(n21118), .B2(keyinput98), .C1(n21129), .C2(
        keyinput107), .A(n20996), .ZN(n21000) );
  AOI22_X1 U23914 ( .A1(n20998), .A2(keyinput71), .B1(n21125), .B2(keyinput108), .ZN(n20997) );
  OAI221_X1 U23915 ( .B1(n20998), .B2(keyinput71), .C1(n21125), .C2(
        keyinput108), .A(n20997), .ZN(n20999) );
  NOR4_X1 U23916 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21003) );
  AND4_X1 U23917 ( .A1(n21006), .A2(n21005), .A3(n21004), .A4(n21003), .ZN(
        n21144) );
  OAI22_X1 U23918 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput85), 
        .B1(P2_REIP_REG_18__SCAN_IN), .B2(keyinput123), .ZN(n21007) );
  AOI221_X1 U23919 ( .B1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput85), 
        .C1(keyinput123), .C2(P2_REIP_REG_18__SCAN_IN), .A(n21007), .ZN(n21014) );
  OAI22_X1 U23920 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(keyinput66), .B1(keyinput69), .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n21008) );
  AOI221_X1 U23921 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(keyinput66), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput69), .A(n21008), .ZN(n21013) );
  OAI22_X1 U23922 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(keyinput68), 
        .B1(keyinput100), .B2(P1_EAX_REG_26__SCAN_IN), .ZN(n21009) );
  AOI221_X1 U23923 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput68), 
        .C1(P1_EAX_REG_26__SCAN_IN), .C2(keyinput100), .A(n21009), .ZN(n21012)
         );
  OAI22_X1 U23924 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(keyinput114), 
        .B1(keyinput112), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n21010) );
  AOI221_X1 U23925 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput114), 
        .C1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .C2(keyinput112), .A(n21010), 
        .ZN(n21011) );
  NAND4_X1 U23926 ( .A1(n21014), .A2(n21013), .A3(n21012), .A4(n21011), .ZN(
        n21042) );
  OAI22_X1 U23927 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput111), 
        .B1(P1_LWORD_REG_14__SCAN_IN), .B2(keyinput89), .ZN(n21015) );
  AOI221_X1 U23928 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput111), 
        .C1(keyinput89), .C2(P1_LWORD_REG_14__SCAN_IN), .A(n21015), .ZN(n21022) );
  OAI22_X1 U23929 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(keyinput99), .B1(
        keyinput83), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n21016) );
  AOI221_X1 U23930 ( .B1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B2(keyinput99), 
        .C1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .C2(keyinput83), .A(n21016), .ZN(
        n21021) );
  OAI22_X1 U23931 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(keyinput67), .B1(
        P2_DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput82), .ZN(n21017) );
  AOI221_X1 U23932 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(keyinput67), .C1(
        keyinput82), .C2(P2_DATAWIDTH_REG_20__SCAN_IN), .A(n21017), .ZN(n21020) );
  OAI22_X1 U23933 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(keyinput119), 
        .B1(keyinput104), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n21018) );
  AOI221_X1 U23934 ( .B1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B2(keyinput119), 
        .C1(P1_REIP_REG_6__SCAN_IN), .C2(keyinput104), .A(n21018), .ZN(n21019)
         );
  NAND4_X1 U23935 ( .A1(n21022), .A2(n21021), .A3(n21020), .A4(n21019), .ZN(
        n21041) );
  OAI22_X1 U23936 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(keyinput94), .B1(
        keyinput76), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n21023) );
  AOI221_X1 U23937 ( .B1(P2_REIP_REG_15__SCAN_IN), .B2(keyinput94), .C1(
        P3_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput76), .A(n21023), .ZN(n21030)
         );
  OAI22_X1 U23938 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(keyinput105), 
        .B1(keyinput64), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n21024) );
  AOI221_X1 U23939 ( .B1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B2(keyinput105), 
        .C1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .C2(keyinput64), .A(n21024), .ZN(
        n21029) );
  OAI22_X1 U23940 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(keyinput93), 
        .B1(keyinput97), .B2(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n21025) );
  AOI221_X1 U23941 ( .B1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B2(keyinput93), 
        .C1(P2_ADDRESS_REG_10__SCAN_IN), .C2(keyinput97), .A(n21025), .ZN(
        n21028) );
  OAI22_X1 U23942 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(keyinput118), 
        .B1(keyinput88), .B2(P3_STATE_REG_2__SCAN_IN), .ZN(n21026) );
  AOI221_X1 U23943 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput118), 
        .C1(P3_STATE_REG_2__SCAN_IN), .C2(keyinput88), .A(n21026), .ZN(n21027)
         );
  NAND4_X1 U23944 ( .A1(n21030), .A2(n21029), .A3(n21028), .A4(n21027), .ZN(
        n21040) );
  OAI22_X1 U23945 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(keyinput65), .B1(
        P3_EBX_REG_1__SCAN_IN), .B2(keyinput122), .ZN(n21031) );
  AOI221_X1 U23946 ( .B1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput65), 
        .C1(keyinput122), .C2(P3_EBX_REG_1__SCAN_IN), .A(n21031), .ZN(n21038)
         );
  OAI22_X1 U23947 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(keyinput96), 
        .B1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B2(keyinput81), .ZN(n21032) );
  AOI221_X1 U23948 ( .B1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B2(keyinput96), 
        .C1(keyinput81), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(n21032), .ZN(
        n21037) );
  OAI22_X1 U23949 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(keyinput113), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(keyinput115), .ZN(n21033) );
  AOI221_X1 U23950 ( .B1(P3_DATAO_REG_28__SCAN_IN), .B2(keyinput113), .C1(
        keyinput115), .C2(P3_LWORD_REG_14__SCAN_IN), .A(n21033), .ZN(n21036)
         );
  OAI22_X1 U23951 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(keyinput110), 
        .B1(P3_LWORD_REG_10__SCAN_IN), .B2(keyinput101), .ZN(n21034) );
  AOI221_X1 U23952 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput110), 
        .C1(keyinput101), .C2(P3_LWORD_REG_10__SCAN_IN), .A(n21034), .ZN(
        n21035) );
  NAND4_X1 U23953 ( .A1(n21038), .A2(n21037), .A3(n21036), .A4(n21035), .ZN(
        n21039) );
  NOR4_X1 U23954 ( .A1(n21042), .A2(n21041), .A3(n21040), .A4(n21039), .ZN(
        n21143) );
  AOI22_X1 U23955 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput18), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(keyinput51), .ZN(n21043) );
  OAI221_X1 U23956 ( .B1(P2_DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput18), .C1(
        P3_LWORD_REG_14__SCAN_IN), .C2(keyinput51), .A(n21043), .ZN(n21050) );
  AOI22_X1 U23957 ( .A1(P3_LWORD_REG_10__SCAN_IN), .A2(keyinput37), .B1(
        P3_INSTQUEUE_REG_7__2__SCAN_IN), .B2(keyinput0), .ZN(n21044) );
  OAI221_X1 U23958 ( .B1(P3_LWORD_REG_10__SCAN_IN), .B2(keyinput37), .C1(
        P3_INSTQUEUE_REG_7__2__SCAN_IN), .C2(keyinput0), .A(n21044), .ZN(
        n21049) );
  AOI22_X1 U23959 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(keyinput48), 
        .B1(P1_EAX_REG_21__SCAN_IN), .B2(keyinput9), .ZN(n21045) );
  OAI221_X1 U23960 ( .B1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B2(keyinput48), 
        .C1(P1_EAX_REG_21__SCAN_IN), .C2(keyinput9), .A(n21045), .ZN(n21048)
         );
  AOI22_X1 U23961 ( .A1(P3_UWORD_REG_4__SCAN_IN), .A2(keyinput8), .B1(
        P1_INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput1), .ZN(n21046) );
  OAI221_X1 U23962 ( .B1(P3_UWORD_REG_4__SCAN_IN), .B2(keyinput8), .C1(
        P1_INSTQUEUE_REG_8__6__SCAN_IN), .C2(keyinput1), .A(n21046), .ZN(
        n21047) );
  NOR4_X1 U23963 ( .A1(n21050), .A2(n21049), .A3(n21048), .A4(n21047), .ZN(
        n21078) );
  AOI22_X1 U23964 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(keyinput7), .B1(
        P3_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput12), .ZN(n21051) );
  OAI221_X1 U23965 ( .B1(P2_BE_N_REG_0__SCAN_IN), .B2(keyinput7), .C1(
        P3_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput12), .A(n21051), .ZN(n21058)
         );
  AOI22_X1 U23966 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(keyinput58), .B1(
        P1_EAX_REG_0__SCAN_IN), .B2(keyinput28), .ZN(n21052) );
  OAI221_X1 U23967 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(keyinput58), .C1(
        P1_EAX_REG_0__SCAN_IN), .C2(keyinput28), .A(n21052), .ZN(n21057) );
  AOI22_X1 U23968 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(keyinput19), .B1(
        P2_FLUSH_REG_SCAN_IN), .B2(keyinput2), .ZN(n21053) );
  OAI221_X1 U23969 ( .B1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B2(keyinput19), 
        .C1(P2_FLUSH_REG_SCAN_IN), .C2(keyinput2), .A(n21053), .ZN(n21056) );
  AOI22_X1 U23970 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(keyinput25), .B1(
        P1_INSTQUEUE_REG_12__0__SCAN_IN), .B2(keyinput32), .ZN(n21054) );
  OAI221_X1 U23971 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(keyinput25), .C1(
        P1_INSTQUEUE_REG_12__0__SCAN_IN), .C2(keyinput32), .A(n21054), .ZN(
        n21055) );
  NOR4_X1 U23972 ( .A1(n21058), .A2(n21057), .A3(n21056), .A4(n21055), .ZN(
        n21077) );
  AOI22_X1 U23973 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(keyinput24), .B1(
        P1_INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput13), .ZN(n21059) );
  OAI221_X1 U23974 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(keyinput24), .C1(
        P1_INSTQUEUE_REG_14__4__SCAN_IN), .C2(keyinput13), .A(n21059), .ZN(
        n21066) );
  AOI22_X1 U23975 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(keyinput61), .B1(
        P2_REIP_REG_7__SCAN_IN), .B2(keyinput62), .ZN(n21060) );
  OAI221_X1 U23976 ( .B1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput61), 
        .C1(P2_REIP_REG_7__SCAN_IN), .C2(keyinput62), .A(n21060), .ZN(n21065)
         );
  AOI22_X1 U23977 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(keyinput50), 
        .B1(P2_ADDRESS_REG_10__SCAN_IN), .B2(keyinput33), .ZN(n21061) );
  OAI221_X1 U23978 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput50), 
        .C1(P2_ADDRESS_REG_10__SCAN_IN), .C2(keyinput33), .A(n21061), .ZN(
        n21064) );
  AOI22_X1 U23979 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(keyinput40), .B1(
        P1_INSTQUEUE_REG_1__5__SCAN_IN), .B2(keyinput6), .ZN(n21062) );
  OAI221_X1 U23980 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(keyinput40), .C1(
        P1_INSTQUEUE_REG_1__5__SCAN_IN), .C2(keyinput6), .A(n21062), .ZN(
        n21063) );
  NOR4_X1 U23981 ( .A1(n21066), .A2(n21065), .A3(n21064), .A4(n21063), .ZN(
        n21076) );
  AOI22_X1 U23982 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(keyinput49), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(keyinput31), .ZN(n21067) );
  OAI221_X1 U23983 ( .B1(P3_DATAO_REG_28__SCAN_IN), .B2(keyinput49), .C1(
        P1_LWORD_REG_5__SCAN_IN), .C2(keyinput31), .A(n21067), .ZN(n21074) );
  AOI22_X1 U23984 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(keyinput27), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(keyinput60), .ZN(n21068) );
  OAI221_X1 U23985 ( .B1(P2_DATAWIDTH_REG_7__SCAN_IN), .B2(keyinput27), .C1(
        P2_EAX_REG_8__SCAN_IN), .C2(keyinput60), .A(n21068), .ZN(n21073) );
  AOI22_X1 U23986 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(keyinput15), .B1(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput46), .ZN(n21069) );
  OAI221_X1 U23987 ( .B1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B2(keyinput15), 
        .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(keyinput46), .A(n21069), 
        .ZN(n21072) );
  AOI22_X1 U23988 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(keyinput20), .B1(
        P1_INSTQUEUE_REG_14__6__SCAN_IN), .B2(keyinput56), .ZN(n21070) );
  OAI221_X1 U23989 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(keyinput20), .C1(
        P1_INSTQUEUE_REG_14__6__SCAN_IN), .C2(keyinput56), .A(n21070), .ZN(
        n21071) );
  NOR4_X1 U23990 ( .A1(n21074), .A2(n21073), .A3(n21072), .A4(n21071), .ZN(
        n21075) );
  NAND4_X1 U23991 ( .A1(n21078), .A2(n21077), .A3(n21076), .A4(n21075), .ZN(
        n21142) );
  AOI22_X1 U23992 ( .A1(n21081), .A2(keyinput3), .B1(n21080), .B2(keyinput45), 
        .ZN(n21079) );
  OAI221_X1 U23993 ( .B1(n21081), .B2(keyinput3), .C1(n21080), .C2(keyinput45), 
        .A(n21079), .ZN(n21092) );
  AOI22_X1 U23994 ( .A1(n21084), .A2(keyinput22), .B1(keyinput17), .B2(n21083), 
        .ZN(n21082) );
  OAI221_X1 U23995 ( .B1(n21084), .B2(keyinput22), .C1(n21083), .C2(keyinput17), .A(n21082), .ZN(n21091) );
  INV_X1 U23996 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n21086) );
  AOI22_X1 U23997 ( .A1(n21086), .A2(keyinput5), .B1(n11837), .B2(keyinput35), 
        .ZN(n21085) );
  OAI221_X1 U23998 ( .B1(n21086), .B2(keyinput5), .C1(n11837), .C2(keyinput35), 
        .A(n21085), .ZN(n21090) );
  XOR2_X1 U23999 ( .A(n10834), .B(keyinput59), .Z(n21088) );
  XNOR2_X1 U24000 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B(keyinput41), .ZN(
        n21087) );
  NAND2_X1 U24001 ( .A1(n21088), .A2(n21087), .ZN(n21089) );
  NOR4_X1 U24002 ( .A1(n21092), .A2(n21091), .A3(n21090), .A4(n21089), .ZN(
        n21140) );
  AOI22_X1 U24003 ( .A1(n21094), .A2(keyinput38), .B1(keyinput52), .B2(n18253), 
        .ZN(n21093) );
  OAI221_X1 U24004 ( .B1(n21094), .B2(keyinput38), .C1(n18253), .C2(keyinput52), .A(n21093), .ZN(n21107) );
  AOI22_X1 U24005 ( .A1(n21097), .A2(keyinput4), .B1(keyinput11), .B2(n21096), 
        .ZN(n21095) );
  OAI221_X1 U24006 ( .B1(n21097), .B2(keyinput4), .C1(n21096), .C2(keyinput11), 
        .A(n21095), .ZN(n21106) );
  AOI22_X1 U24007 ( .A1(n21100), .A2(keyinput47), .B1(keyinput14), .B2(n21099), 
        .ZN(n21098) );
  OAI221_X1 U24008 ( .B1(n21100), .B2(keyinput47), .C1(n21099), .C2(keyinput14), .A(n21098), .ZN(n21105) );
  INV_X1 U24009 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n21102) );
  AOI22_X1 U24010 ( .A1(n21103), .A2(keyinput23), .B1(keyinput55), .B2(n21102), 
        .ZN(n21101) );
  OAI221_X1 U24011 ( .B1(n21103), .B2(keyinput23), .C1(n21102), .C2(keyinput55), .A(n21101), .ZN(n21104) );
  NOR4_X1 U24012 ( .A1(n21107), .A2(n21106), .A3(n21105), .A4(n21104), .ZN(
        n21139) );
  AOI22_X1 U24013 ( .A1(n21109), .A2(keyinput26), .B1(n12136), .B2(keyinput29), 
        .ZN(n21108) );
  OAI221_X1 U24014 ( .B1(n21109), .B2(keyinput26), .C1(n12136), .C2(keyinput29), .A(n21108), .ZN(n21113) );
  XOR2_X1 U24015 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B(keyinput10), .Z(
        n21112) );
  XNOR2_X1 U24016 ( .A(n21110), .B(keyinput54), .ZN(n21111) );
  OR3_X1 U24017 ( .A1(n21113), .A2(n21112), .A3(n21111), .ZN(n21121) );
  AOI22_X1 U24018 ( .A1(n21116), .A2(keyinput30), .B1(keyinput57), .B2(n21115), 
        .ZN(n21114) );
  OAI221_X1 U24019 ( .B1(n21116), .B2(keyinput30), .C1(n21115), .C2(keyinput57), .A(n21114), .ZN(n21120) );
  AOI22_X1 U24020 ( .A1(n21118), .A2(keyinput34), .B1(keyinput36), .B2(n14330), 
        .ZN(n21117) );
  OAI221_X1 U24021 ( .B1(n21118), .B2(keyinput34), .C1(n14330), .C2(keyinput36), .A(n21117), .ZN(n21119) );
  NOR3_X1 U24022 ( .A1(n21121), .A2(n21120), .A3(n21119), .ZN(n21138) );
  AOI22_X1 U24023 ( .A1(n21123), .A2(keyinput16), .B1(n11164), .B2(keyinput42), 
        .ZN(n21122) );
  OAI221_X1 U24024 ( .B1(n21123), .B2(keyinput16), .C1(n11164), .C2(keyinput42), .A(n21122), .ZN(n21136) );
  AOI22_X1 U24025 ( .A1(n21126), .A2(keyinput21), .B1(keyinput44), .B2(n21125), 
        .ZN(n21124) );
  OAI221_X1 U24026 ( .B1(n21126), .B2(keyinput21), .C1(n21125), .C2(keyinput44), .A(n21124), .ZN(n21135) );
  AOI22_X1 U24027 ( .A1(n21129), .A2(keyinput43), .B1(n21128), .B2(keyinput53), 
        .ZN(n21127) );
  OAI221_X1 U24028 ( .B1(n21129), .B2(keyinput43), .C1(n21128), .C2(keyinput53), .A(n21127), .ZN(n21134) );
  AOI22_X1 U24029 ( .A1(n21132), .A2(keyinput63), .B1(n21131), .B2(keyinput39), 
        .ZN(n21130) );
  OAI221_X1 U24030 ( .B1(n21132), .B2(keyinput63), .C1(n21131), .C2(keyinput39), .A(n21130), .ZN(n21133) );
  NOR4_X1 U24031 ( .A1(n21136), .A2(n21135), .A3(n21134), .A4(n21133), .ZN(
        n21137) );
  NAND4_X1 U24032 ( .A1(n21140), .A2(n21139), .A3(n21138), .A4(n21137), .ZN(
        n21141) );
  AOI211_X1 U24033 ( .C1(n21144), .C2(n21143), .A(n21142), .B(n21141), .ZN(
        n21147) );
  NAND2_X1 U24034 ( .A1(n21145), .A2(P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n21146) );
  XNOR2_X1 U24035 ( .A(n21147), .B(n21146), .ZN(P3_U3009) );
  INV_X1 U13979 ( .A(n11906), .ZN(n11138) );
  INV_X1 U12824 ( .A(n10412), .ZN(n10394) );
  CLKBUF_X2 U11329 ( .A(n10393), .Z(n9661) );
  NAND2_X1 U11161 ( .A1(n11236), .A2(n11189), .ZN(n13368) );
  NAND2_X1 U11225 ( .A1(n14531), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14493) );
  BUF_X2 U11089 ( .A(n15796), .Z(n9645) );
  CLKBUF_X1 U11092 ( .A(n11839), .Z(n11784) );
  OAI22_X1 U11117 ( .A1(n13161), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13275), 
        .B2(n11126), .ZN(n11103) );
  NAND2_X1 U11124 ( .A1(n12447), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10431) );
  CLKBUF_X1 U11145 ( .A(n10643), .Z(n13811) );
  CLKBUF_X1 U11341 ( .A(n10432), .Z(n9654) );
  INV_X1 U11432 ( .A(n10393), .ZN(n10584) );
  CLKBUF_X1 U11474 ( .A(n12949), .Z(n14053) );
  CLKBUF_X1 U11550 ( .A(n14137), .Z(n14138) );
  CLKBUF_X2 U12235 ( .A(n10401), .Z(n19422) );
  CLKBUF_X1 U12336 ( .A(n13369), .Z(n9665) );
  CLKBUF_X1 U12458 ( .A(n19331), .Z(n19344) );
  CLKBUF_X1 U12690 ( .A(n15179), .Z(n15180) );
  XNOR2_X1 U12848 ( .A(n12205), .B(n12444), .ZN(n12536) );
  AND2_X1 U12854 ( .A1(n13578), .A2(n10194), .ZN(n21148) );
  CLKBUF_X1 U12941 ( .A(n17565), .Z(n17575) );
endmodule

