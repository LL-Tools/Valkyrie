

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, 
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, 
        keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, 
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, 
        keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060;

  INV_X1 U3527 ( .A(n5647), .ZN(n4317) );
  INV_X2 U3528 ( .A(n4601), .ZN(n4427) );
  BUF_X2 U3529 ( .A(n3461), .Z(n4350) );
  CLKBUF_X2 U3530 ( .A(n3441), .Z(n4383) );
  AND4_X1 U3531 ( .A1(n4744), .A2(n3421), .A3(n6707), .A4(
        STATE2_REG_0__SCAN_IN), .ZN(n3422) );
  CLKBUF_X2 U3532 ( .A(n3462), .Z(n3442) );
  CLKBUF_X2 U3533 ( .A(n3427), .Z(n4384) );
  CLKBUF_X2 U3534 ( .A(n3523), .Z(n4386) );
  CLKBUF_X2 U3535 ( .A(n3448), .Z(n4388) );
  CLKBUF_X2 U3536 ( .A(n3370), .Z(n3079) );
  CLKBUF_X2 U3537 ( .A(n3491), .Z(n3440) );
  CLKBUF_X2 U3538 ( .A(n4349), .Z(n4387) );
  CLKBUF_X2 U3539 ( .A(n3304), .Z(n4264) );
  CLKBUF_X1 U3540 ( .A(n3419), .Z(n4815) );
  NAND2_X1 U3541 ( .A1(n3729), .A2(n3391), .ZN(n3221) );
  CLKBUF_X2 U3542 ( .A(n3380), .Z(n4827) );
  CLKBUF_X1 U3543 ( .A(n3384), .Z(n4843) );
  AND2_X2 U3544 ( .A1(n4613), .A2(n4758), .ZN(n4349) );
  AND2_X2 U3545 ( .A1(n3186), .A2(n4740), .ZN(n4385) );
  AND3_X1 U3546 ( .A1(n3121), .A2(n3761), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3688) );
  AND2_X1 U3547 ( .A1(n3137), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3273)
         );
  NOR2_X1 U3548 ( .A1(n3417), .A2(n3761), .ZN(n5778) );
  NOR2_X1 U3549 ( .A1(n3412), .A2(n3391), .ZN(n4584) );
  BUF_X1 U3550 ( .A(n3386), .Z(n4823) );
  NOR2_X1 U3551 ( .A1(n3748), .A2(n4827), .ZN(n4421) );
  AND2_X1 U3552 ( .A1(n3380), .A2(n3417), .ZN(n5774) );
  INV_X2 U3553 ( .A(n4455), .ZN(n3080) );
  INV_X2 U3554 ( .A(n3080), .ZN(n4300) );
  INV_X1 U3555 ( .A(n5694), .ZN(n6364) );
  NAND2_X1 U3556 ( .A1(n3919), .A2(n3918), .ZN(n4867) );
  AND2_X2 U3558 ( .A1(n4717), .A2(n4740), .ZN(n3441) );
  OR2_X2 U3559 ( .A1(n4803), .A2(n3187), .ZN(n3581) );
  NAND2_X2 U3560 ( .A1(n3131), .A2(n3530), .ZN(n4804) );
  NAND2_X2 U3561 ( .A1(n6067), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3570)
         );
  XNOR2_X2 U3562 ( .A(n3589), .B(n3588), .ZN(n4914) );
  NAND2_X2 U3563 ( .A1(n3587), .A2(n3586), .ZN(n3589) );
  NAND2_X1 U3564 ( .A1(n3223), .A2(n3408), .ZN(n3458) );
  NAND2_X2 U3565 ( .A1(n3517), .A2(n5527), .ZN(n3720) );
  CLKBUF_X1 U3566 ( .A(n3546), .Z(n5521) );
  INV_X2 U3568 ( .A(n4836), .ZN(n3121) );
  INV_X2 U3569 ( .A(n3380), .ZN(n3761) );
  CLKBUF_X2 U3571 ( .A(n4356), .Z(n4378) );
  AND2_X2 U3572 ( .A1(n3274), .A2(n4717), .ZN(n3468) );
  INV_X2 U3573 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4603) );
  OAI21_X1 U3574 ( .B1(n4472), .B2(n4303), .A(n3120), .ZN(n3119) );
  XNOR2_X1 U3575 ( .A(n3142), .B(n5899), .ZN(n3881) );
  OR2_X1 U3576 ( .A1(n5900), .A2(n5901), .ZN(n3142) );
  NAND2_X1 U3577 ( .A1(n3157), .A2(n3155), .ZN(n5926) );
  NAND2_X1 U3578 ( .A1(n3130), .A2(n3129), .ZN(n5963) );
  AOI21_X1 U3579 ( .B1(n3247), .B2(n3245), .A(n3108), .ZN(n3244) );
  NOR2_X1 U3580 ( .A1(n3658), .A2(n3123), .ZN(n3261) );
  OAI21_X1 U3581 ( .B1(n3933), .B2(n3187), .A(n3613), .ZN(n3615) );
  AND2_X1 U3582 ( .A1(n4699), .A2(n3571), .ZN(n6426) );
  NAND2_X1 U3583 ( .A1(n3902), .A2(n4581), .ZN(n4598) );
  NAND2_X1 U3584 ( .A1(n3509), .A2(n3508), .ZN(n3125) );
  AND2_X1 U3585 ( .A1(n6479), .A2(n6181), .ZN(n5153) );
  OR2_X1 U3586 ( .A1(n3868), .A2(n3859), .ZN(n6181) );
  NAND2_X1 U3587 ( .A1(n3756), .A2(n5533), .ZN(n3868) );
  OR3_X2 U3588 ( .A1(n5529), .A2(n6457), .A3(n4425), .ZN(n6373) );
  NAND2_X1 U3589 ( .A1(n3458), .A2(n3457), .ZN(n3482) );
  NAND2_X1 U3590 ( .A1(n3138), .A2(n3389), .ZN(n3486) );
  AND2_X1 U3591 ( .A1(n3378), .A2(n3377), .ZN(n3409) );
  CLKBUF_X1 U3592 ( .A(n3748), .Z(n4607) );
  NOR2_X2 U3593 ( .A1(n3415), .A2(n3387), .ZN(n3725) );
  AND2_X1 U3594 ( .A1(n3382), .A2(n3383), .ZN(n3423) );
  AND2_X1 U3595 ( .A1(n3384), .A2(n3761), .ZN(n3546) );
  INV_X1 U3596 ( .A(n3678), .ZN(n5833) );
  BUF_X2 U3597 ( .A(n3381), .Z(n4836) );
  CLKBUF_X1 U3598 ( .A(n3390), .Z(n3412) );
  NAND2_X1 U3599 ( .A1(n3288), .A2(n3287), .ZN(n3393) );
  NAND3_X1 U3600 ( .A1(n3149), .A2(n3263), .A3(n3269), .ZN(n3390) );
  AND4_X1 U3601 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3355)
         );
  AND4_X1 U3602 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3356)
         );
  AND4_X1 U3603 ( .A1(n3341), .A2(n3340), .A3(n3339), .A4(n3338), .ZN(n3357)
         );
  AND4_X1 U3604 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3320)
         );
  AND4_X1 U3605 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3319)
         );
  AND4_X1 U3606 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3318)
         );
  AND4_X1 U3607 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3287)
         );
  AND4_X1 U3608 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3317)
         );
  AND4_X1 U3609 ( .A1(n3282), .A2(n3281), .A3(n3280), .A4(n3279), .ZN(n3288)
         );
  AND3_X1 U3610 ( .A1(n3272), .A2(n3271), .A3(n3270), .ZN(n3149) );
  BUF_X2 U3611 ( .A(n4385), .Z(n4216) );
  AND2_X2 U3612 ( .A1(n3273), .A2(n4717), .ZN(n3370) );
  NAND2_X2 U3613 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6742), .ZN(n4541) );
  AND2_X2 U3614 ( .A1(n3224), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4613)
         );
  AND2_X2 U3615 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4758) );
  INV_X1 U3616 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3224) );
  XNOR2_X2 U3617 ( .A(n3208), .B(n4410), .ZN(n4447) );
  OAI21_X2 U3618 ( .B1(n5150), .B2(n3128), .A(n3107), .ZN(n6017) );
  NAND2_X2 U3619 ( .A1(n3647), .A2(n3646), .ZN(n5150) );
  NOR2_X4 U3620 ( .A1(n5593), .A2(n4209), .ZN(n5466) );
  OAI21_X1 U3621 ( .B1(n3419), .B2(n3390), .A(n3385), .ZN(n3299) );
  NAND2_X1 U3622 ( .A1(n3402), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3403) );
  AOI21_X1 U3623 ( .B1(n3244), .B2(n3144), .A(n3143), .ZN(n3129) );
  AOI22_X1 U3625 ( .A1(n3514), .A2(n5177), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3513), .ZN(n3404) );
  XNOR2_X1 U3626 ( .A(n4742), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3708)
         );
  NAND2_X1 U3627 ( .A1(n3701), .A2(n3700), .ZN(n3711) );
  CLKBUF_X1 U3628 ( .A(n3492), .Z(n3467) );
  CLKBUF_X1 U3629 ( .A(n3493), .Z(n3459) );
  INV_X1 U3630 ( .A(n3674), .ZN(n3255) );
  NAND2_X1 U3631 ( .A1(n3628), .A2(n3627), .ZN(n3648) );
  INV_X1 U3632 ( .A(n3630), .ZN(n3628) );
  INV_X1 U3633 ( .A(n5481), .ZN(n3675) );
  INV_X1 U3634 ( .A(n3677), .ZN(n3124) );
  NAND2_X1 U3635 ( .A1(n5451), .A2(n5450), .ZN(n5917) );
  INV_X1 U3636 ( .A(n5954), .ZN(n5451) );
  INV_X1 U3637 ( .A(n3261), .ZN(n3128) );
  NOR2_X1 U3638 ( .A1(n4927), .A2(n3198), .ZN(n5156) );
  NAND2_X1 U3639 ( .A1(n3200), .A2(n3199), .ZN(n3198) );
  INV_X1 U3640 ( .A(n3201), .ZN(n3200) );
  NOR2_X1 U3641 ( .A1(n3203), .A2(n5157), .ZN(n3199) );
  AND2_X1 U3642 ( .A1(n3264), .A2(n4843), .ZN(n3150) );
  NAND2_X1 U3643 ( .A1(n6365), .A2(EBX_REG_16__SCAN_IN), .ZN(n3218) );
  AND2_X1 U3644 ( .A1(n6373), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U3645 ( .A1(n5547), .A2(n4316), .ZN(n4417) );
  CLKBUF_X1 U3646 ( .A(n3896), .Z(n4405) );
  OR2_X1 U3647 ( .A1(n4208), .A2(n5665), .ZN(n4209) );
  NOR2_X1 U3648 ( .A1(n5593), .A2(n5665), .ZN(n5664) );
  NOR2_X1 U3649 ( .A1(n3211), .A2(n3210), .ZN(n3209) );
  INV_X1 U3650 ( .A(n4077), .ZN(n4078) );
  NAND2_X1 U3651 ( .A1(n4061), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4077)
         );
  INV_X1 U3652 ( .A(n4060), .ZN(n4061) );
  NAND2_X1 U3653 ( .A1(n3923), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3927)
         );
  NAND2_X1 U3654 ( .A1(n4317), .A2(n3779), .ZN(n4589) );
  NOR2_X2 U3655 ( .A1(n3091), .A2(n5548), .ZN(n5547) );
  NAND2_X1 U3656 ( .A1(n4774), .A2(n3417), .ZN(n4746) );
  NAND2_X1 U3657 ( .A1(n3174), .A2(n3739), .ZN(n3723) );
  OAI21_X1 U3658 ( .B1(n3159), .B2(n3103), .A(n3086), .ZN(n3158) );
  AOI21_X1 U3659 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6541), .A(n5178), .ZN(
        n6648) );
  AND2_X1 U3660 ( .A1(n3755), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U3661 ( .A1(n3850), .A2(n5521), .ZN(n4788) );
  AND2_X1 U3662 ( .A1(n6373), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U3663 ( .A1(n3177), .A2(n3176), .ZN(n3175) );
  INV_X1 U3664 ( .A(n3682), .ZN(n3176) );
  AND2_X1 U3665 ( .A1(n4385), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U3666 ( .A1(n3523), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        INSTQUEUE_REG_8__6__SCAN_IN), .B2(n4385), .ZN(n3279) );
  INV_X1 U3667 ( .A(n3385), .ZN(n3379) );
  NAND2_X1 U3668 ( .A1(n3153), .A2(n3102), .ZN(n3630) );
  INV_X1 U3669 ( .A(n3605), .ZN(n3604) );
  NAND2_X1 U3670 ( .A1(n3261), .A2(n3127), .ZN(n3126) );
  INV_X1 U3671 ( .A(n5151), .ZN(n3127) );
  NAND2_X1 U3672 ( .A1(n3221), .A2(n3546), .ZN(n3421) );
  OR2_X1 U3673 ( .A1(n3437), .A2(n3436), .ZN(n3554) );
  NAND3_X1 U3674 ( .A1(n3134), .A2(n3404), .A3(n3403), .ZN(n3484) );
  INV_X1 U3675 ( .A(n4286), .ZN(n3514) );
  CLKBUF_X1 U3676 ( .A(n3486), .Z(n3487) );
  OR2_X1 U3677 ( .A1(n3454), .A2(n3453), .ZN(n3651) );
  NAND2_X1 U3678 ( .A1(n3461), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3322)
         );
  AND2_X1 U3679 ( .A1(n5623), .A2(n5620), .ZN(n5604) );
  NOR2_X1 U3680 ( .A1(n6935), .A2(n3205), .ZN(n3204) );
  INV_X1 U3681 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U3682 ( .A1(n3232), .A2(n5760), .ZN(n3231) );
  INV_X1 U3683 ( .A(n5352), .ZN(n3232) );
  NOR2_X1 U3684 ( .A1(n3392), .A2(n5179), .ZN(n3896) );
  AND2_X1 U3685 ( .A1(n4300), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4296)
         );
  AOI21_X1 U3686 ( .B1(n3256), .B2(n3254), .A(n3104), .ZN(n3253) );
  NAND2_X1 U3687 ( .A1(n5917), .A2(n3259), .ZN(n3157) );
  NOR2_X1 U3688 ( .A1(n5454), .A2(n3260), .ZN(n3259) );
  INV_X1 U3689 ( .A(n5453), .ZN(n3260) );
  OR2_X1 U3690 ( .A1(n4300), .A2(n5452), .ZN(n5453) );
  INV_X1 U3691 ( .A(n4589), .ZN(n4313) );
  AND2_X1 U3692 ( .A1(n3815), .A2(n5822), .ZN(n3196) );
  AND2_X1 U3693 ( .A1(n3814), .A2(n5814), .ZN(n3815) );
  NAND2_X1 U3694 ( .A1(n3663), .A2(n6037), .ZN(n3251) );
  OR2_X1 U3695 ( .A1(n5168), .A2(n5167), .ZN(n3203) );
  AND2_X1 U3696 ( .A1(n4601), .A2(n4317), .ZN(n3784) );
  NAND2_X1 U3697 ( .A1(n5647), .A2(n4601), .ZN(n4309) );
  NOR2_X1 U3698 ( .A1(n5153), .A2(n3164), .ZN(n3163) );
  NOR2_X1 U3699 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n3165), .ZN(n3164)
         );
  INV_X1 U3700 ( .A(n6479), .ZN(n3165) );
  INV_X1 U3701 ( .A(n3688), .ZN(n3713) );
  AND4_X2 U3702 ( .A1(n3357), .A2(n3356), .A3(n3355), .A4(n3354), .ZN(n3380)
         );
  AND2_X1 U3703 ( .A1(n3747), .A2(n3746), .ZN(n4773) );
  AND2_X1 U3704 ( .A1(n3396), .A2(n3110), .ZN(n4774) );
  INV_X1 U3705 ( .A(n4225), .ZN(n4404) );
  CLKBUF_X1 U3706 ( .A(n4345), .Z(n4284) );
  NAND2_X1 U3707 ( .A1(n4078), .A2(n3087), .ZN(n4192) );
  AND2_X1 U3708 ( .A1(n3235), .A2(n4098), .ZN(n3234) );
  INV_X1 U3709 ( .A(n5678), .ZN(n4098) );
  AND2_X1 U3710 ( .A1(n3974), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3989)
         );
  NOR2_X1 U3711 ( .A1(n3944), .A2(n6881), .ZN(n3974) );
  AND2_X1 U3712 ( .A1(n3606), .A2(n3545), .ZN(n3926) );
  NAND2_X1 U3713 ( .A1(n4770), .A2(n5533), .ZN(n4662) );
  NAND2_X1 U3714 ( .A1(n3189), .A2(n3193), .ZN(n3188) );
  INV_X1 U3715 ( .A(n3848), .ZN(n3193) );
  INV_X1 U3716 ( .A(n3190), .ZN(n3189) );
  NAND2_X1 U3717 ( .A1(n6122), .A2(n3090), .ZN(n3185) );
  NAND2_X1 U3718 ( .A1(n3157), .A2(n5457), .ZN(n5462) );
  NAND2_X1 U3719 ( .A1(n5917), .A2(n5453), .ZN(n5947) );
  INV_X1 U3720 ( .A(n3148), .ZN(n3147) );
  OAI21_X1 U3721 ( .B1(n3244), .B2(n3085), .A(n3256), .ZN(n3148) );
  NAND2_X1 U3722 ( .A1(n3163), .A2(n3162), .ZN(n3161) );
  INV_X1 U3723 ( .A(n3870), .ZN(n3162) );
  INV_X1 U3724 ( .A(n6017), .ZN(n3250) );
  INV_X1 U3725 ( .A(n3251), .ZN(n3246) );
  NOR2_X1 U3726 ( .A1(n3251), .A2(n3248), .ZN(n3247) );
  INV_X1 U3727 ( .A(n6012), .ZN(n3248) );
  NAND2_X1 U3728 ( .A1(n3655), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3656)
         );
  NAND2_X1 U3729 ( .A1(n5150), .A2(n5151), .ZN(n3657) );
  NAND2_X1 U3730 ( .A1(n3778), .A2(n3777), .ZN(n4927) );
  INV_X1 U3731 ( .A(n4868), .ZN(n3778) );
  INV_X1 U3732 ( .A(n3163), .ZN(n6455) );
  XNOR2_X1 U3733 ( .A(n4804), .B(n3583), .ZN(n3910) );
  CLKBUF_X1 U3734 ( .A(n4734), .Z(n4735) );
  INV_X1 U3735 ( .A(n5216), .ZN(n5267) );
  NOR2_X1 U3736 ( .A1(n6589), .A2(n6227), .ZN(n6500) );
  AND3_X1 U3737 ( .A1(n6731), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6593) );
  INV_X1 U3738 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6541) );
  OR2_X1 U3739 ( .A1(n6231), .A2(n4874), .ZN(n4878) );
  NAND2_X1 U3740 ( .A1(n4814), .A2(n4813), .ZN(n5178) );
  NAND2_X1 U3741 ( .A1(n6236), .A2(n4812), .ZN(n4814) );
  OR2_X1 U3742 ( .A1(n6231), .A2(n4806), .ZN(n4817) );
  INV_X1 U3743 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5179) );
  OR2_X2 U3744 ( .A1(n3376), .A2(n3375), .ZN(n3417) );
  INV_X1 U3745 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U3746 ( .A1(n6311), .A2(n5988), .ZN(n3220) );
  NOR3_X1 U3747 ( .A1(n3219), .A2(n5698), .A3(n3217), .ZN(n3216) );
  OAI21_X1 U3748 ( .B1(n6151), .B2(n6350), .A(n3218), .ZN(n3217) );
  INV_X1 U3749 ( .A(n5704), .ZN(n3219) );
  INV_X1 U3750 ( .A(n5780), .ZN(n6311) );
  INV_X1 U3751 ( .A(n6365), .ZN(n6306) );
  OR2_X1 U3752 ( .A1(n6714), .A2(n5023), .ZN(n4425) );
  NAND2_X1 U3753 ( .A1(n4409), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3208)
         );
  NAND2_X1 U3754 ( .A1(n4078), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4082)
         );
  OR2_X1 U3755 ( .A1(n4662), .A2(n4780), .ZN(n6245) );
  INV_X1 U3756 ( .A(n6056), .ZN(n6422) );
  INV_X1 U3757 ( .A(n6245), .ZN(n6428) );
  XNOR2_X1 U3758 ( .A(n4328), .B(n4327), .ZN(n5789) );
  NAND2_X1 U3759 ( .A1(n4419), .A2(n4325), .ZN(n4328) );
  XNOR2_X1 U3760 ( .A(n3119), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3136)
         );
  NAND2_X1 U3761 ( .A1(n5479), .A2(n4458), .ZN(n3120) );
  NAND2_X1 U3762 ( .A1(n4477), .A2(n3096), .ZN(n4452) );
  AOI21_X1 U3763 ( .B1(n4454), .B2(n6470), .A(n5893), .ZN(n3179) );
  NAND2_X1 U3764 ( .A1(n4453), .A2(n6837), .ZN(n3180) );
  OR2_X1 U3765 ( .A1(n3868), .A2(n3765), .ZN(n6473) );
  AND2_X1 U3766 ( .A1(n3852), .A2(n3851), .ZN(n6470) );
  INV_X1 U3767 ( .A(n4807), .ZN(n6499) );
  CLKBUF_X1 U3768 ( .A(n4803), .Z(n6231) );
  INV_X1 U3769 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6731) );
  INV_X1 U3770 ( .A(n5397), .ZN(n6728) );
  NAND2_X1 U3771 ( .A1(n6500), .A2(n6499), .ZN(n6551) );
  AND2_X1 U3772 ( .A1(n4300), .A2(n3671), .ZN(n3674) );
  AOI21_X1 U3773 ( .B1(n3575), .B2(n3388), .A(n5774), .ZN(n3377) );
  NAND2_X1 U3774 ( .A1(n3174), .A2(n3169), .ZN(n3168) );
  INV_X1 U3775 ( .A(n3741), .ZN(n3169) );
  NAND2_X1 U3776 ( .A1(n3172), .A2(n3171), .ZN(n3170) );
  NAND2_X1 U3777 ( .A1(n3714), .A2(n3686), .ZN(n3172) );
  AND2_X1 U3778 ( .A1(n3175), .A2(n3166), .ZN(n3171) );
  NAND2_X1 U3779 ( .A1(n3684), .A2(n3685), .ZN(n3167) );
  CLKBUF_X1 U3780 ( .A(n4375), .Z(n4355) );
  NOR2_X1 U3781 ( .A1(n3669), .A2(n3674), .ZN(n3254) );
  OR2_X1 U3782 ( .A1(n4300), .A2(n3664), .ZN(n3665) );
  OR2_X1 U3783 ( .A1(n3603), .A2(n3602), .ZN(n3611) );
  OR2_X1 U3784 ( .A1(n3503), .A2(n3502), .ZN(n3504) );
  OR2_X1 U3785 ( .A1(n3529), .A2(n3528), .ZN(n3585) );
  OR2_X1 U3786 ( .A1(n3729), .A2(n3724), .ZN(n4612) );
  NOR2_X1 U3787 ( .A1(n3268), .A2(n3267), .ZN(n3269) );
  NAND4_X1 U3788 ( .A1(n3399), .A2(n3398), .A3(n3391), .A4(n3392), .ZN(n3748)
         );
  NAND2_X1 U3789 ( .A1(n3379), .A2(n3393), .ZN(n4582) );
  AND2_X1 U3790 ( .A1(n3240), .A2(n4285), .ZN(n3239) );
  NOR2_X1 U3791 ( .A1(n3241), .A2(n5568), .ZN(n3240) );
  INV_X1 U3792 ( .A(n3242), .ZN(n3241) );
  AND2_X1 U3793 ( .A1(n5491), .A2(n5467), .ZN(n3242) );
  NOR2_X1 U3794 ( .A1(n4223), .A2(n6973), .ZN(n3214) );
  AND2_X1 U3795 ( .A1(n4190), .A2(n5604), .ZN(n5594) );
  NOR2_X1 U3796 ( .A1(n4186), .A2(n3213), .ZN(n3212) );
  INV_X1 U3797 ( .A(n4192), .ZN(n4099) );
  NAND2_X1 U3798 ( .A1(n5707), .A2(n4065), .ZN(n3237) );
  NOR2_X1 U3799 ( .A1(n4064), .A2(n3236), .ZN(n3235) );
  INV_X1 U3800 ( .A(n5691), .ZN(n3236) );
  INV_X1 U3801 ( .A(n5737), .ZN(n3230) );
  XNOR2_X1 U3802 ( .A(n3648), .B(n3638), .ZN(n3888) );
  INV_X1 U3803 ( .A(n3896), .ZN(n4402) );
  INV_X1 U3804 ( .A(n3153), .ZN(n3544) );
  NAND2_X1 U3805 ( .A1(n3153), .A2(n3542), .ZN(n3606) );
  INV_X1 U3806 ( .A(n3894), .ZN(n3922) );
  OAI21_X1 U3807 ( .B1(n4803), .B2(n3972), .A(n4225), .ZN(n3907) );
  AND2_X1 U3808 ( .A1(n3889), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3894) );
  OR2_X1 U3809 ( .A1(n3474), .A2(n3473), .ZN(n3566) );
  OR2_X1 U3810 ( .A1(n3114), .A2(n3191), .ZN(n3190) );
  NAND2_X1 U3811 ( .A1(n3192), .A2(n5569), .ZN(n3191) );
  INV_X1 U3812 ( .A(n5596), .ZN(n3192) );
  INV_X1 U3813 ( .A(n3257), .ZN(n3256) );
  OAI21_X1 U3814 ( .B1(n3258), .B2(n3667), .A(n3670), .ZN(n3257) );
  AND2_X1 U3815 ( .A1(n3196), .A2(n3195), .ZN(n3194) );
  INV_X1 U3816 ( .A(n5705), .ZN(n3195) );
  INV_X1 U3817 ( .A(n3784), .ZN(n3836) );
  INV_X1 U3818 ( .A(n3656), .ZN(n3123) );
  NAND2_X1 U3819 ( .A1(n3202), .A2(n4933), .ZN(n3201) );
  INV_X1 U3820 ( .A(n4926), .ZN(n3202) );
  OR2_X1 U3821 ( .A1(n3857), .A2(n3856), .ZN(n3860) );
  NAND2_X1 U3822 ( .A1(n3425), .A2(n3426), .ZN(n3457) );
  OAI21_X1 U3823 ( .B1(n3415), .B2(n3418), .A(n3417), .ZN(n3424) );
  NAND2_X1 U3824 ( .A1(n3563), .A2(n3478), .ZN(n3551) );
  OAI211_X1 U3825 ( .C1(n3713), .C2(n5250), .A(n3456), .B(n3455), .ZN(n3550)
         );
  NAND2_X1 U3826 ( .A1(n3484), .A2(n3407), .ZN(n3481) );
  NAND2_X1 U3827 ( .A1(n3572), .A2(n3125), .ZN(n3583) );
  AND2_X2 U3828 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4717) );
  INV_X1 U3829 ( .A(n3860), .ZN(n4609) );
  NAND2_X1 U3830 ( .A1(n3420), .A2(n4584), .ZN(n4744) );
  AND4_X1 U3831 ( .A1(n4827), .A2(n4815), .A3(n3121), .A4(n3392), .ZN(n3420)
         );
  AND2_X1 U3832 ( .A1(n3719), .A2(n3718), .ZN(n3739) );
  OR2_X1 U3833 ( .A1(n3717), .A2(n3716), .ZN(n3719) );
  NOR2_X1 U3834 ( .A1(n3707), .A2(n3706), .ZN(n3159) );
  NAND2_X1 U3835 ( .A1(n3490), .A2(n3489), .ZN(n3511) );
  AND2_X1 U3836 ( .A1(n3735), .A2(n3734), .ZN(n4569) );
  INV_X1 U3837 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4726) );
  NAND2_X1 U3838 ( .A1(n3893), .A2(n4813), .ZN(n3563) );
  INV_X1 U3839 ( .A(n3417), .ZN(n3384) );
  INV_X1 U3840 ( .A(n3390), .ZN(n3386) );
  INV_X1 U3841 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4984) );
  AND2_X1 U3842 ( .A1(n6704), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U3843 ( .A1(n4836), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3517) );
  INV_X1 U3844 ( .A(n4773), .ZN(n4552) );
  AND2_X1 U3845 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5724), .ZN(n5701) );
  NAND2_X1 U3846 ( .A1(n3393), .A2(n3392), .ZN(n5515) );
  OR2_X1 U3847 ( .A1(n3760), .A2(n4566), .ZN(n4567) );
  NAND2_X1 U3848 ( .A1(n3227), .A2(n3900), .ZN(n4581) );
  INV_X1 U3849 ( .A(n4579), .ZN(n3227) );
  OR2_X1 U3850 ( .A1(n4661), .A2(READY_N), .ZN(n4663) );
  OR2_X1 U3851 ( .A1(n4368), .A2(n5537), .ZN(n4408) );
  OR2_X1 U3852 ( .A1(n4280), .A2(n5559), .ZN(n4366) );
  NOR2_X1 U3853 ( .A1(n4262), .A2(n6849), .ZN(n4279) );
  NAND2_X1 U3854 ( .A1(n5466), .A2(n3242), .ZN(n5567) );
  NAND2_X1 U3855 ( .A1(n3214), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4262)
         );
  INV_X1 U3856 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6973) );
  INV_X1 U3857 ( .A(n3214), .ZN(n4244) );
  NOR2_X1 U3858 ( .A1(n4143), .A2(n5930), .ZN(n4100) );
  NAND2_X1 U3859 ( .A1(n4100), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4223)
         );
  OR2_X1 U3860 ( .A1(n4171), .A2(n5940), .ZN(n4143) );
  INV_X1 U3861 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4186) );
  NAND2_X1 U3862 ( .A1(n4099), .A2(n3212), .ZN(n4188) );
  NAND2_X1 U3863 ( .A1(n4099), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4194)
         );
  NAND2_X1 U3864 ( .A1(n3989), .A2(n3116), .ZN(n4060) );
  AND2_X1 U3865 ( .A1(n4019), .A2(n4018), .ZN(n5819) );
  CLKBUF_X1 U3866 ( .A(n5736), .Z(n5820) );
  AND2_X1 U3867 ( .A1(n3959), .A2(n3958), .ZN(n5352) );
  AND3_X1 U3868 ( .A1(n3957), .A2(n3956), .A3(n3955), .ZN(n3958) );
  OR2_X1 U3869 ( .A1(n3936), .A2(n3884), .ZN(n3944) );
  NAND2_X1 U3870 ( .A1(n3934), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3936)
         );
  NOR2_X1 U3871 ( .A1(n3927), .A2(n3930), .ZN(n3934) );
  INV_X1 U3872 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3930) );
  INV_X1 U3873 ( .A(n4922), .ZN(n3229) );
  AND2_X1 U3874 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3882), .ZN(n3923)
         );
  NAND2_X1 U3875 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U3876 ( .A1(n3228), .A2(n3226), .ZN(n4908) );
  INV_X1 U3877 ( .A(n3907), .ZN(n3228) );
  INV_X1 U3878 ( .A(n3226), .ZN(n3906) );
  OR3_X1 U3879 ( .A1(n4300), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n4299), 
        .ZN(n4468) );
  AND2_X1 U3880 ( .A1(n4312), .A2(n4311), .ZN(n5548) );
  AND2_X1 U3881 ( .A1(n4296), .A2(n3676), .ZN(n3141) );
  NAND2_X1 U3882 ( .A1(n3185), .A2(n3183), .ZN(n6071) );
  AND2_X1 U3883 ( .A1(n6107), .A2(n3181), .ZN(n3183) );
  NOR2_X1 U3884 ( .A1(n3872), .A2(n3105), .ZN(n3181) );
  NOR3_X1 U3885 ( .A1(n5611), .A2(n3114), .A3(n5596), .ZN(n5570) );
  AND2_X1 U3886 ( .A1(n3841), .A2(n3840), .ZN(n5482) );
  NOR2_X1 U3887 ( .A1(n3080), .A2(n5458), .ZN(n5459) );
  AND2_X1 U3888 ( .A1(n5461), .A2(n6094), .ZN(n3152) );
  OR2_X1 U3889 ( .A1(n5609), .A2(n5608), .ZN(n5611) );
  NOR2_X1 U3890 ( .A1(n3156), .A2(n3117), .ZN(n3155) );
  INV_X1 U3891 ( .A(n5457), .ZN(n3156) );
  AND2_X1 U3892 ( .A1(n3810), .A2(n3809), .ZN(n5730) );
  NAND2_X1 U3893 ( .A1(n5823), .A2(n3196), .ZN(n5732) );
  INV_X1 U3894 ( .A(n3266), .ZN(n3245) );
  AND2_X1 U3895 ( .A1(n5823), .A2(n5822), .ZN(n5825) );
  AND2_X1 U3896 ( .A1(n5741), .A2(n3804), .ZN(n5823) );
  INV_X1 U3897 ( .A(n5742), .ZN(n3804) );
  AND2_X1 U3898 ( .A1(n3801), .A2(n3800), .ZN(n5749) );
  OR2_X1 U3899 ( .A1(n4455), .A2(n3661), .ZN(n6037) );
  NAND2_X1 U3900 ( .A1(n3657), .A2(n3261), .ZN(n3154) );
  AND2_X1 U3901 ( .A1(n3796), .A2(n3795), .ZN(n5157) );
  OR2_X1 U3902 ( .A1(n3197), .A2(n4927), .ZN(n5170) );
  OR2_X1 U3903 ( .A1(n3203), .A2(n3201), .ZN(n3197) );
  AND2_X1 U3904 ( .A1(n3790), .A2(n3789), .ZN(n5168) );
  OR2_X1 U3905 ( .A1(n4927), .A2(n3201), .ZN(n5169) );
  NOR2_X1 U3906 ( .A1(n4916), .A2(n6160), .ZN(n6216) );
  NOR2_X1 U3907 ( .A1(n3776), .A2(n3775), .ZN(n4869) );
  INV_X1 U3908 ( .A(n5153), .ZN(n4916) );
  XNOR2_X1 U3909 ( .A(n3458), .B(n3222), .ZN(n3893) );
  INV_X1 U3910 ( .A(n3457), .ZN(n3222) );
  XNOR2_X1 U3911 ( .A(n3481), .B(n3482), .ZN(n4604) );
  CLKBUF_X1 U3912 ( .A(n4713), .Z(n4714) );
  INV_X1 U3913 ( .A(n6230), .ZN(n6638) );
  INV_X1 U3914 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3895) );
  INV_X1 U3915 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3122) );
  INV_X1 U3916 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4742) );
  OR2_X1 U3917 ( .A1(n6727), .A2(n5214), .ZN(n5308) );
  OR2_X1 U3918 ( .A1(n6722), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5397) );
  OR2_X1 U3919 ( .A1(n6727), .A2(n4987), .ZN(n4988) );
  OR2_X1 U3920 ( .A1(n6231), .A2(n5101), .ZN(n6589) );
  OR2_X1 U3921 ( .A1(n5064), .A2(n6227), .ZN(n5068) );
  AND2_X1 U3922 ( .A1(n6727), .A2(n6231), .ZN(n6639) );
  AND2_X1 U3923 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4810), .ZN(n4808)
         );
  NAND2_X1 U3924 ( .A1(n5179), .A2(n6244), .ZN(n4423) );
  OR2_X1 U3925 ( .A1(n4662), .A2(n4554), .ZN(n4661) );
  NAND2_X1 U3926 ( .A1(n4661), .A2(n4558), .ZN(n5529) );
  NAND2_X1 U3927 ( .A1(n4827), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U3928 ( .A1(n3417), .A2(n5522), .ZN(n5528) );
  NAND2_X1 U3929 ( .A1(n4448), .A2(n6373), .ZN(n5780) );
  NOR2_X1 U3930 ( .A1(n4447), .A2(n6704), .ZN(n4448) );
  AND2_X1 U3931 ( .A1(n5779), .A2(n4428), .ZN(n6361) );
  AND2_X1 U3932 ( .A1(n5779), .A2(n4431), .ZN(n6359) );
  INV_X1 U3933 ( .A(n6324), .ZN(n6369) );
  INV_X1 U3934 ( .A(n6358), .ZN(n6347) );
  AND2_X1 U3935 ( .A1(n5779), .A2(n4435), .ZN(n6365) );
  AOI22_X1 U3936 ( .A1(n4420), .A2(n4419), .B1(n4418), .B2(n4417), .ZN(n5500)
         );
  INV_X1 U3937 ( .A(n5829), .ZN(n6375) );
  INV_X1 U3938 ( .A(n6379), .ZN(n5830) );
  NAND2_X1 U3939 ( .A1(n4587), .A2(n4586), .ZN(n6379) );
  OR2_X1 U3940 ( .A1(n4794), .A2(n4427), .ZN(n4586) );
  OR3_X1 U3941 ( .A1(n4770), .A2(n6711), .A3(n4771), .ZN(n4587) );
  INV_X1 U3942 ( .A(n3392), .ZN(n5513) );
  NOR2_X2 U3943 ( .A1(n5885), .A2(n5515), .ZN(n5873) );
  AND2_X1 U3944 ( .A1(n5889), .A2(n5834), .ZN(n5874) );
  INV_X1 U3945 ( .A(n5889), .ZN(n5885) );
  NAND2_X1 U3946 ( .A1(n5889), .A2(n4800), .ZN(n5891) );
  OR3_X1 U3947 ( .A1(n4662), .A2(n4591), .A3(n5522), .ZN(n6402) );
  AND2_X1 U3948 ( .A1(n6402), .A2(n4786), .ZN(n6743) );
  INV_X1 U3949 ( .A(n4798), .ZN(n6419) );
  INV_X1 U3950 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6849) );
  OR2_X1 U3951 ( .A1(n5465), .A2(n5468), .ZN(n5854) );
  INV_X1 U3952 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5930) );
  INV_X1 U3953 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5940) );
  OAI21_X1 U3954 ( .B1(n5624), .B2(n5623), .A(n5622), .ZN(n5945) );
  NAND2_X1 U3955 ( .A1(n4078), .A2(n3209), .ZN(n4083) );
  AND2_X1 U3956 ( .A1(n3989), .A2(n3088), .ZN(n4046) );
  NAND2_X1 U3957 ( .A1(n3989), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3990)
         );
  INV_X1 U3958 ( .A(n6218), .ZN(n6457) );
  NAND2_X1 U3959 ( .A1(n6245), .A2(n4287), .ZN(n6056) );
  NOR2_X1 U3960 ( .A1(n3182), .A2(n3106), .ZN(n6086) );
  INV_X1 U3961 ( .A(n3185), .ZN(n3182) );
  NOR2_X1 U3962 ( .A1(n6129), .A2(n3873), .ZN(n6092) );
  AOI22_X1 U3963 ( .A1(n5462), .A2(n5461), .B1(n5918), .B2(n5955), .ZN(n5919)
         );
  INV_X1 U3964 ( .A(n5462), .ZN(n5936) );
  NOR3_X1 U3965 ( .A1(n3867), .A2(n6205), .A3(n6759), .ZN(n6122) );
  INV_X1 U3966 ( .A(n3161), .ZN(n6119) );
  NAND2_X1 U3967 ( .A1(n3250), .A2(n3266), .ZN(n3249) );
  OR2_X1 U3968 ( .A1(n4286), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U3969 ( .A1(n3657), .A2(n3656), .ZN(n6048) );
  OR2_X1 U3970 ( .A1(n5155), .A2(n5154), .ZN(n6215) );
  INV_X1 U3971 ( .A(n6460), .ZN(n6160) );
  CLKBUF_X1 U3972 ( .A(n4941), .Z(n4942) );
  OR2_X1 U3973 ( .A1(n3868), .A2(n4771), .ZN(n6460) );
  OR2_X1 U3974 ( .A1(n3868), .A2(n4746), .ZN(n6479) );
  AND2_X1 U3975 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n4860) );
  CLKBUF_X1 U3977 ( .A(n4604), .Z(n4605) );
  INV_X1 U3978 ( .A(n4735), .ZN(n6721) );
  AND2_X1 U3979 ( .A1(n4862), .A2(n5178), .ZN(n6732) );
  NAND2_X1 U3980 ( .A1(n4770), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6236) );
  NOR2_X2 U3981 ( .A1(n4988), .A2(n6499), .ZN(n5433) );
  OAI211_X1 U3982 ( .C1(n6550), .C2(n6584), .A(n6549), .B(n6548), .ZN(n6579)
         );
  NAND2_X1 U3983 ( .A1(n5272), .A2(n5271), .ZN(n5297) );
  INV_X1 U3984 ( .A(n5303), .ZN(n5266) );
  INV_X1 U3985 ( .A(n6696), .ZN(n5391) );
  OAI21_X1 U3986 ( .B1(n5366), .B2(n6640), .A(n5365), .ZN(n5389) );
  NOR2_X1 U3987 ( .A1(n5064), .A2(n5265), .ZN(n6695) );
  AOI22_X1 U3988 ( .A1(n6647), .A2(n6645), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6650), .ZN(n6702) );
  OR3_X1 U3989 ( .A1(n4980), .A2(n6722), .A3(n4879), .ZN(n4880) );
  NOR2_X2 U3990 ( .A1(n4878), .A2(n6499), .ZN(n5060) );
  AND2_X1 U3991 ( .A1(n6065), .A2(DATAI_24_), .ZN(n6652) );
  AND2_X1 U3992 ( .A1(n6065), .A2(DATAI_25_), .ZN(n6658) );
  AND2_X1 U3993 ( .A1(n6065), .A2(DATAI_27_), .ZN(n6669) );
  INV_X1 U3994 ( .A(n6670), .ZN(n6607) );
  INV_X1 U3995 ( .A(n6612), .ZN(n6675) );
  AND2_X1 U3996 ( .A1(n6065), .A2(DATAI_29_), .ZN(n6681) );
  INV_X1 U3997 ( .A(n5173), .ZN(n5209) );
  AND2_X1 U3998 ( .A1(n6065), .A2(DATAI_31_), .ZN(n6697) );
  OR2_X1 U3999 ( .A1(n5178), .A2(n4801), .ZN(n6661) );
  AND2_X1 U4000 ( .A1(n6065), .A2(DATAI_17_), .ZN(n6657) );
  OR2_X1 U4001 ( .A1(n4849), .A2(n4823), .ZN(n6601) );
  OR2_X1 U4002 ( .A1(n5178), .A2(n4910), .ZN(n6667) );
  AND2_X1 U4003 ( .A1(n6065), .A2(DATAI_18_), .ZN(n6664) );
  OR2_X1 U4004 ( .A1(n4849), .A2(n4848), .ZN(n6606) );
  OR2_X1 U4005 ( .A1(n5178), .A2(n4847), .ZN(n6673) );
  OR2_X1 U4006 ( .A1(n5178), .A2(n4835), .ZN(n6679) );
  AND2_X1 U4007 ( .A1(n6065), .A2(DATAI_20_), .ZN(n6676) );
  OR2_X1 U4008 ( .A1(n4849), .A2(n5833), .ZN(n6616) );
  AND2_X1 U4009 ( .A1(n6065), .A2(DATAI_21_), .ZN(n6682) );
  OR2_X1 U4010 ( .A1(n4849), .A2(n4815), .ZN(n6621) );
  OR2_X1 U4011 ( .A1(n5178), .A2(n5324), .ZN(n6691) );
  AND2_X1 U4012 ( .A1(n6065), .A2(DATAI_22_), .ZN(n6688) );
  OR2_X1 U4013 ( .A1(n4849), .A2(n5513), .ZN(n6628) );
  OR2_X1 U4014 ( .A1(n5178), .A2(n4831), .ZN(n6701) );
  INV_X1 U4015 ( .A(n5253), .ZN(n4853) );
  AND2_X1 U4016 ( .A1(n6065), .A2(DATAI_23_), .ZN(n6694) );
  OAI21_X1 U4017 ( .B1(n4820), .B2(n4819), .A(n4818), .ZN(n4854) );
  OR2_X1 U4018 ( .A1(n4817), .A2(n6499), .ZN(n5212) );
  AND2_X1 U4019 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4424), .ZN(n5023) );
  NOR2_X1 U4020 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6707) );
  OR2_X1 U4021 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n5525) );
  AND2_X1 U4022 ( .A1(n4509), .A2(n6740), .ZN(n6719) );
  INV_X1 U4023 ( .A(READY_N), .ZN(n6706) );
  INV_X1 U4024 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U4025 ( .A1(n3720), .A2(n3417), .ZN(n3679) );
  OR2_X1 U4026 ( .A1(n5699), .A2(n3215), .ZN(U2811) );
  NAND2_X1 U4027 ( .A1(n3220), .A2(n3216), .ZN(n3215) );
  OAI21_X1 U4028 ( .B1(n5839), .B2(n6057), .A(n4490), .ZN(n4491) );
  OAI21_X1 U4029 ( .B1(n5845), .B2(n6057), .A(n4292), .ZN(n4293) );
  OAI21_X1 U4030 ( .B1(n3136), .B2(n6473), .A(n3135), .ZN(U2987) );
  NOR2_X1 U4031 ( .A1(n3084), .A2(n3100), .ZN(n3135) );
  NAND2_X1 U4032 ( .A1(n4467), .A2(n3097), .ZN(U2988) );
  NAND2_X1 U4033 ( .A1(n4452), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3178) );
  AND2_X1 U4034 ( .A1(n4481), .A2(n4480), .ZN(n4482) );
  OR2_X1 U4035 ( .A1(n5792), .A2(n6221), .ZN(n4481) );
  NAND2_X1 U4036 ( .A1(n3679), .A2(n3678), .ZN(n3684) );
  AND2_X1 U4037 ( .A1(n3194), .A2(n5693), .ZN(n3081) );
  OR2_X2 U4038 ( .A1(n3333), .A2(n3332), .ZN(n3392) );
  OR2_X1 U4039 ( .A1(n5166), .A2(n3231), .ZN(n3082) );
  AND3_X1 U4040 ( .A1(n3364), .A2(n3363), .A3(n3362), .ZN(n3083) );
  OR2_X1 U4041 ( .A1(n4308), .A2(n4307), .ZN(n3084) );
  AND2_X1 U4042 ( .A1(n3233), .A2(n3238), .ZN(n5690) );
  NAND2_X1 U4043 ( .A1(n3665), .A2(n3669), .ZN(n3085) );
  NAND2_X1 U4044 ( .A1(n3249), .A2(n3247), .ZN(n6011) );
  INV_X1 U4045 ( .A(n3872), .ZN(n3184) );
  AND2_X1 U4046 ( .A1(n3722), .A2(n3721), .ZN(n3086) );
  NAND2_X1 U4047 ( .A1(n3133), .A2(n3593), .ZN(n4931) );
  AND2_X1 U4048 ( .A1(n3209), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3087)
         );
  AND2_X1 U4049 ( .A1(n3204), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3088)
         );
  AND2_X1 U4050 ( .A1(n3212), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3089)
         );
  AND2_X1 U4051 ( .A1(n6099), .A2(n3865), .ZN(n3090) );
  OR2_X1 U4052 ( .A1(n5611), .A2(n3188), .ZN(n3091) );
  AND2_X1 U4053 ( .A1(n5466), .A2(n5467), .ZN(n5465) );
  AND2_X1 U4054 ( .A1(n5466), .A2(n3240), .ZN(n4283) );
  AND2_X1 U4055 ( .A1(n6122), .A2(n3865), .ZN(n3092) );
  AND2_X1 U4056 ( .A1(n3185), .A2(n6107), .ZN(n3093) );
  NAND2_X1 U4057 ( .A1(n3233), .A2(n3235), .ZN(n5676) );
  NOR2_X1 U4058 ( .A1(n5166), .A2(n5352), .ZN(n5353) );
  AND4_X1 U4059 ( .A1(n3361), .A2(n3360), .A3(n3359), .A4(n3358), .ZN(n3094)
         );
  NAND2_X1 U4060 ( .A1(n3154), .A2(n3659), .ZN(n6040) );
  OR2_X1 U4061 ( .A1(n3231), .A2(n3988), .ZN(n3095) );
  NOR2_X1 U4062 ( .A1(n5611), .A2(n5596), .ZN(n5473) );
  INV_X1 U4063 ( .A(n3714), .ZN(n3174) );
  OR2_X2 U4064 ( .A1(n3391), .A2(n4827), .ZN(n3779) );
  AOI21_X1 U4065 ( .B1(n3761), .B2(n5833), .A(n3417), .ZN(n3697) );
  INV_X1 U4066 ( .A(n3697), .ZN(n3177) );
  AND2_X1 U4067 ( .A1(n3249), .A2(n3246), .ZN(n6010) );
  OR2_X1 U4068 ( .A1(n6216), .A2(n4460), .ZN(n3096) );
  AND3_X1 U4069 ( .A1(n3180), .A2(n3179), .A3(n3178), .ZN(n3097) );
  OR2_X1 U4070 ( .A1(n5611), .A2(n3190), .ZN(n3098) );
  AND2_X2 U4071 ( .A1(n4613), .A2(n3274), .ZN(n3491) );
  OR2_X1 U4072 ( .A1(n4589), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3099)
         );
  AND2_X1 U4073 ( .A1(n5789), .A2(n6470), .ZN(n3100) );
  AND2_X1 U4074 ( .A1(n3660), .A2(n3659), .ZN(n3101) );
  AND2_X1 U4075 ( .A1(n3604), .A2(n3542), .ZN(n3102) );
  INV_X1 U4076 ( .A(n3685), .ZN(n3173) );
  INV_X1 U4077 ( .A(n3669), .ZN(n3258) );
  AND2_X1 U4078 ( .A1(n3713), .A2(n3745), .ZN(n3103) );
  NOR2_X1 U4079 ( .A1(n4300), .A2(n3673), .ZN(n3104) );
  INV_X1 U4080 ( .A(n3393), .ZN(n3419) );
  NOR2_X1 U4081 ( .A1(n6216), .A2(n3875), .ZN(n3105) );
  NAND2_X1 U4082 ( .A1(n6107), .A2(n3184), .ZN(n3106) );
  AND2_X1 U4083 ( .A1(n3126), .A2(n3101), .ZN(n3107) );
  AND2_X1 U4084 ( .A1(n4300), .A2(n6189), .ZN(n3108) );
  AND2_X1 U4085 ( .A1(n3678), .A2(n3173), .ZN(n3109) );
  AND2_X1 U4086 ( .A1(n3221), .A2(n3264), .ZN(n3110) );
  AND2_X1 U4087 ( .A1(n3256), .A2(n3255), .ZN(n3111) );
  AND2_X1 U4088 ( .A1(n4582), .A2(n3392), .ZN(n3112) );
  OR2_X1 U4089 ( .A1(n3095), .A2(n3230), .ZN(n3113) );
  INV_X1 U4090 ( .A(n3160), .ZN(n6205) );
  NAND2_X1 U4091 ( .A1(n3115), .A2(n3161), .ZN(n3160) );
  INV_X1 U4092 ( .A(n6473), .ZN(n6462) );
  NOR2_X1 U4093 ( .A1(n4927), .A2(n4926), .ZN(n4925) );
  INV_X1 U4094 ( .A(n3187), .ZN(n3687) );
  NAND2_X1 U4095 ( .A1(n3678), .A2(n3417), .ZN(n3187) );
  NOR2_X1 U4096 ( .A1(n5748), .A2(n5749), .ZN(n5741) );
  NAND2_X1 U4097 ( .A1(n4865), .A2(n4867), .ZN(n4866) );
  OR2_X1 U4098 ( .A1(n5485), .A2(n5482), .ZN(n3114) );
  NAND2_X1 U4099 ( .A1(n3132), .A2(n3616), .ZN(n4955) );
  NOR2_X1 U4100 ( .A1(n5634), .A2(n3829), .ZN(n5628) );
  AND3_X1 U4101 ( .A1(n4865), .A2(n3229), .A3(n4867), .ZN(n4923) );
  NAND2_X1 U4102 ( .A1(n3225), .A2(n3892), .ZN(n4597) );
  OR2_X1 U4103 ( .A1(n6460), .A2(n6159), .ZN(n3115) );
  NOR2_X1 U4104 ( .A1(n5679), .A2(n5681), .ZN(n5646) );
  NAND2_X1 U4105 ( .A1(n3989), .A2(n3204), .ZN(n3206) );
  AND2_X1 U4106 ( .A1(n3088), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3116)
         );
  AND2_X1 U4107 ( .A1(n4300), .A2(n6110), .ZN(n3117) );
  INV_X1 U4108 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5976) );
  AND2_X1 U4109 ( .A1(n5823), .A2(n3194), .ZN(n3118) );
  INV_X1 U4110 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3210) );
  INV_X1 U4111 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5578) );
  AND2_X1 U4112 ( .A1(n3761), .A2(n3417), .ZN(n4601) );
  INV_X1 U4113 ( .A(n4064), .ZN(n3238) );
  AND2_X1 U4114 ( .A1(n4506), .A2(STATE_REG_1__SCAN_IN), .ZN(n6742) );
  INV_X1 U4115 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3213) );
  AND2_X2 U4116 ( .A1(n4603), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4611)
         );
  AND2_X2 U4117 ( .A1(n3531), .A2(n4804), .ZN(n3153) );
  OAI21_X1 U4118 ( .B1(n3388), .B2(n3121), .A(n3112), .ZN(n3415) );
  NAND2_X1 U4119 ( .A1(n3419), .A2(n3385), .ZN(n3388) );
  NOR2_X4 U4120 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3186) );
  AND2_X2 U4121 ( .A1(n3122), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4740)
         );
  NAND2_X1 U4122 ( .A1(n4455), .A2(n3654), .ZN(n3655) );
  AND2_X2 U4123 ( .A1(n4298), .A2(n3676), .ZN(n4457) );
  NAND2_X2 U4124 ( .A1(n3124), .A2(n3675), .ZN(n4298) );
  NAND2_X1 U4125 ( .A1(n3252), .A2(n3253), .ZN(n3677) );
  XNOR2_X1 U4126 ( .A(n3572), .B(n3125), .ZN(n4803) );
  OR2_X2 U4127 ( .A1(n3145), .A2(n6017), .ZN(n3130) );
  NAND2_X1 U4128 ( .A1(n3910), .A2(n3687), .ZN(n3587) );
  NAND2_X1 U4129 ( .A1(n3480), .A2(n3479), .ZN(n3572) );
  NAND2_X1 U4130 ( .A1(n4734), .A2(n4813), .ZN(n3131) );
  NAND2_X1 U4131 ( .A1(n4931), .A2(n4930), .ZN(n3132) );
  NAND2_X1 U4132 ( .A1(n4941), .A2(n4940), .ZN(n3133) );
  INV_X1 U4133 ( .A(n3481), .ZN(n3483) );
  NAND2_X1 U4134 ( .A1(n3486), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3134) );
  OAI21_X1 U4135 ( .B1(n3136), .B2(n6245), .A(n4414), .ZN(U2955) );
  INV_X1 U4136 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3137) );
  AND2_X2 U4137 ( .A1(n3186), .A2(n3273), .ZN(n3493) );
  NAND2_X1 U4138 ( .A1(n3139), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3138) );
  NAND4_X1 U4139 ( .A1(n3423), .A2(n3409), .A3(n3725), .A4(n3140), .ZN(n3139)
         );
  NAND2_X1 U4140 ( .A1(n3400), .A2(n5833), .ZN(n3140) );
  AND2_X1 U4141 ( .A1(n4298), .A2(n3141), .ZN(n5901) );
  INV_X1 U4142 ( .A(n3665), .ZN(n3143) );
  INV_X1 U4143 ( .A(n3247), .ZN(n3144) );
  INV_X1 U4144 ( .A(n3244), .ZN(n3145) );
  NAND2_X1 U4145 ( .A1(n3243), .A2(n3244), .ZN(n6001) );
  NAND2_X1 U4146 ( .A1(n6017), .A2(n3247), .ZN(n3243) );
  OR2_X1 U4147 ( .A1(n3243), .A2(n3085), .ZN(n3146) );
  NAND2_X1 U4148 ( .A1(n3146), .A2(n3147), .ZN(n5954) );
  NAND3_X1 U4149 ( .A1(n3396), .A2(n3221), .A3(n3150), .ZN(n3760) );
  NAND2_X1 U4150 ( .A1(n5462), .A2(n3152), .ZN(n3151) );
  NAND2_X1 U4151 ( .A1(n5463), .A2(n3151), .ZN(n5464) );
  NAND2_X2 U4152 ( .A1(n3648), .A2(n3650), .ZN(n4455) );
  OAI21_X2 U4153 ( .B1(n4604), .B2(STATE2_REG_0__SCAN_IN), .A(n3438), .ZN(
        n3552) );
  NAND2_X2 U4154 ( .A1(n3158), .A2(n3723), .ZN(n4770) );
  NAND2_X1 U4155 ( .A1(n3679), .A2(n3109), .ZN(n3166) );
  NAND3_X1 U4156 ( .A1(n3170), .A2(n3168), .A3(n3167), .ZN(n3696) );
  AND2_X2 U4157 ( .A1(n3274), .A2(n3186), .ZN(n3304) );
  INV_X1 U4158 ( .A(n3186), .ZN(n4858) );
  AND2_X2 U4159 ( .A1(n4758), .A2(n3186), .ZN(n3461) );
  NAND2_X1 U4160 ( .A1(n5823), .A2(n3081), .ZN(n5679) );
  INV_X1 U4161 ( .A(n3206), .ZN(n4022) );
  NAND2_X2 U4162 ( .A1(n4447), .A2(n3207), .ZN(n5694) );
  INV_X1 U4163 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4164 ( .A1(n4099), .A2(n3089), .ZN(n4171) );
  NAND2_X1 U4165 ( .A1(n3486), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4166 ( .A1(n4805), .A2(n4057), .ZN(n3225) );
  NAND2_X1 U4167 ( .A1(n4598), .A2(n4597), .ZN(n3226) );
  NAND2_X1 U4168 ( .A1(n4923), .A2(n4963), .ZN(n4962) );
  NAND2_X2 U4169 ( .A1(n3909), .A2(n3908), .ZN(n4865) );
  NOR2_X1 U4170 ( .A1(n5166), .A2(n3095), .ZN(n5735) );
  OR2_X2 U4171 ( .A1(n5166), .A2(n3113), .ZN(n5736) );
  CLKBUF_X1 U4172 ( .A(n3237), .Z(n3233) );
  NAND2_X2 U4173 ( .A1(n3237), .A2(n3234), .ZN(n5593) );
  NAND2_X1 U4174 ( .A1(n5466), .A2(n3239), .ZN(n4345) );
  NAND2_X1 U4175 ( .A1(n5963), .A2(n3111), .ZN(n3252) );
  NAND3_X1 U4176 ( .A1(n3606), .A2(n3545), .A3(n3687), .ZN(n3549) );
  AND2_X1 U4177 ( .A1(n6541), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3690)
         );
  OR2_X1 U4178 ( .A1(n3906), .A2(n4599), .ZN(n6368) );
  NAND2_X1 U4179 ( .A1(n4457), .A2(n4297), .ZN(n4472) );
  NAND2_X1 U4180 ( .A1(n4472), .A2(n4471), .ZN(n4473) );
  NAND2_X1 U4181 ( .A1(n4021), .A2(n4020), .ZN(n5707) );
  INV_X1 U4182 ( .A(n5736), .ZN(n4021) );
  AND2_X2 U4183 ( .A1(n4611), .A2(n4740), .ZN(n3523) );
  AND2_X2 U4184 ( .A1(n4611), .A2(n3273), .ZN(n3492) );
  AND2_X1 U4185 ( .A1(n3370), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3267) );
  CLKBUF_X1 U4186 ( .A(n4804), .Z(n5101) );
  NAND2_X1 U4187 ( .A1(n4385), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4188 ( .A1(n4385), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3293) );
  CLKBUF_X1 U4189 ( .A(n4485), .Z(n5545) );
  OAI21_X1 U4190 ( .B1(n3730), .B2(n5513), .A(n3546), .ZN(n3383) );
  NAND2_X1 U4191 ( .A1(n4582), .A2(n4836), .ZN(n3730) );
  BUF_X1 U4192 ( .A(n3677), .Z(n5480) );
  INV_X1 U4193 ( .A(n5164), .ZN(n3942) );
  XNOR2_X1 U4194 ( .A(n4407), .B(n4406), .ZN(n5514) );
  AOI22_X1 U4195 ( .A1(n4356), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3296) );
  NAND2_X1 U4196 ( .A1(n4503), .A2(n6651), .ZN(n6057) );
  INV_X2 U4197 ( .A(n6057), .ZN(n6065) );
  AOI21_X1 U4198 ( .B1(n3888), .B2(n4057), .A(n3887), .ZN(n5165) );
  INV_X1 U4199 ( .A(n5165), .ZN(n3943) );
  NAND2_X2 U4200 ( .A1(n3563), .A2(n3562), .ZN(n4807) );
  OR2_X1 U4201 ( .A1(n3405), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3262)
         );
  AND4_X1 U4202 ( .A1(n3278), .A2(n3277), .A3(n3276), .A4(n3275), .ZN(n3263)
         );
  AND2_X1 U4203 ( .A1(n3395), .A2(n4827), .ZN(n3264) );
  INV_X1 U4204 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6881) );
  INV_X1 U4205 ( .A(n6722), .ZN(n6651) );
  NAND2_X1 U4206 ( .A1(n5217), .A2(n5179), .ZN(n6722) );
  INV_X1 U4207 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3903) );
  OR2_X1 U4208 ( .A1(n4606), .A2(n5515), .ZN(n3265) );
  AND2_X1 U4209 ( .A1(n6026), .A2(n6018), .ZN(n3266) );
  INV_X1 U4210 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6482) );
  INV_X1 U4211 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4764) );
  AND4_X2 U4212 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3381)
         );
  INV_X1 U4213 ( .A(n5747), .ZN(n3988) );
  NAND2_X2 U4214 ( .A1(n5889), .A2(n4799), .ZN(n5892) );
  OR2_X1 U4215 ( .A1(n5456), .A2(n5934), .ZN(n5457) );
  AOI22_X1 U4216 ( .A1(n4349), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3491), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3278) );
  INV_X1 U4217 ( .A(n3708), .ZN(n3710) );
  OR2_X1 U4218 ( .A1(n3541), .A2(n3540), .ZN(n3608) );
  INV_X1 U4219 ( .A(n3504), .ZN(n3574) );
  AND2_X1 U4220 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6482), .ZN(n3716)
         );
  NAND2_X1 U4221 ( .A1(n4349), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3303)
         );
  AOI21_X1 U4222 ( .B1(n3711), .B2(n3710), .A(n3709), .ZN(n3715) );
  BUF_X1 U4223 ( .A(n3492), .Z(n4348) );
  OR2_X1 U4224 ( .A1(n4258), .A2(n4257), .ZN(n4275) );
  OR2_X1 U4225 ( .A1(n3626), .A2(n3625), .ZN(n3640) );
  AND2_X1 U4226 ( .A1(n3380), .A2(n3391), .ZN(n3575) );
  NAND2_X1 U4227 ( .A1(n3688), .A2(n3687), .ZN(n3714) );
  INV_X1 U4228 ( .A(n3755), .ZN(n3513) );
  AND2_X1 U4229 ( .A1(n3715), .A2(n3712), .ZN(n3745) );
  INV_X1 U4230 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4314) );
  AND2_X1 U4231 ( .A1(n3323), .A2(n3322), .ZN(n3324) );
  NAND2_X1 U4232 ( .A1(n4349), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3345)
         );
  NOR2_X1 U4233 ( .A1(n4612), .A2(n4813), .ZN(n4397) );
  INV_X1 U4234 ( .A(n5819), .ZN(n4020) );
  AND2_X1 U4235 ( .A1(n4296), .A2(n4301), .ZN(n4297) );
  NAND2_X1 U4236 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5458) );
  INV_X1 U4237 ( .A(n5956), .ZN(n5450) );
  AND2_X1 U4238 ( .A1(n3813), .A2(n3812), .ZN(n5814) );
  NOR2_X1 U4239 ( .A1(n3187), .A2(n3649), .ZN(n3650) );
  AOI22_X1 U4240 ( .A1(n3174), .A2(n3745), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4813), .ZN(n3722) );
  AND4_X1 U4241 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n3354)
         );
  INV_X1 U4242 ( .A(n4397), .ZN(n4364) );
  INV_X1 U4243 ( .A(n3972), .ZN(n4057) );
  NAND2_X1 U4244 ( .A1(n4324), .A2(n4323), .ZN(n4325) );
  NAND2_X1 U4245 ( .A1(n4470), .A2(n4469), .ZN(n4471) );
  AND2_X1 U4246 ( .A1(n3833), .A2(n3832), .ZN(n5608) );
  INV_X1 U4247 ( .A(n5649), .ZN(n3825) );
  AND2_X1 U4248 ( .A1(n4911), .A2(n4869), .ZN(n3777) );
  NAND2_X1 U4249 ( .A1(n3516), .A2(n3515), .ZN(n6544) );
  OR2_X1 U4250 ( .A1(n5178), .A2(n5217), .ZN(n4849) );
  INV_X1 U4251 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6935) );
  INV_X1 U4252 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3884) );
  INV_X1 U4253 ( .A(n6359), .ZN(n6321) );
  INV_X1 U4254 ( .A(n4423), .ZN(n4370) );
  AND2_X1 U4255 ( .A1(n4057), .A2(n4035), .ZN(n5812) );
  NAND2_X1 U4256 ( .A1(n4815), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3972) );
  INV_X1 U4257 ( .A(n4326), .ZN(n4327) );
  OR2_X1 U4258 ( .A1(n4300), .A2(n6152), .ZN(n5992) );
  NAND2_X1 U4259 ( .A1(n6707), .A2(n4813), .ZN(n4286) );
  NAND2_X1 U4260 ( .A1(n4568), .A2(n4567), .ZN(n4796) );
  INV_X1 U4261 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n5217) );
  OR2_X1 U4262 ( .A1(n5401), .A2(n5784), .ZN(n4983) );
  NAND2_X1 U4263 ( .A1(n4989), .A2(n6499), .ZN(n5146) );
  AOI21_X1 U4264 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5402), .A(n5178), .ZN(
        n6549) );
  OR2_X1 U4265 ( .A1(n6589), .A2(n5265), .ZN(n6623) );
  INV_X1 U4266 ( .A(n6639), .ZN(n5064) );
  OR2_X1 U4267 ( .A1(n4849), .A2(n4843), .ZN(n6596) );
  INV_X1 U4268 ( .A(n6312), .ZN(n6333) );
  AND2_X1 U4269 ( .A1(n6373), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U4270 ( .A1(n4417), .A2(n4317), .ZN(n4419) );
  AND2_X1 U4271 ( .A1(n6379), .A2(n3392), .ZN(n6376) );
  AOI21_X1 U4272 ( .B1(n4796), .B2(n5533), .A(n4795), .ZN(n4797) );
  INV_X1 U4273 ( .A(n4786), .ZN(n6744) );
  AND2_X1 U4274 ( .A1(n4746), .A2(n4788), .ZN(n4591) );
  OR2_X1 U4275 ( .A1(n4663), .A2(n4843), .ZN(n4798) );
  INV_X2 U4276 ( .A(n6421), .ZN(n6415) );
  AND2_X2 U4277 ( .A1(n4663), .A2(n6421), .ZN(n6418) );
  AND2_X1 U4278 ( .A1(n4173), .A2(n4172), .ZN(n5638) );
  OR2_X1 U4279 ( .A1(n3758), .A2(n3757), .ZN(n4780) );
  INV_X1 U4280 ( .A(n6432), .ZN(n6060) );
  OR2_X1 U4281 ( .A1(n5794), .A2(n6221), .ZN(n3878) );
  AND2_X1 U4282 ( .A1(n3824), .A2(n3823), .ZN(n5649) );
  XNOR2_X1 U4283 ( .A(n3570), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4700)
         );
  OR3_X1 U4284 ( .A1(n4573), .A2(n4796), .A3(n4572), .ZN(n4763) );
  NOR2_X2 U4285 ( .A1(n5308), .A2(n6499), .ZN(n6490) );
  OAI211_X1 U4286 ( .C1(n5400), .C2(n5404), .A(n6549), .B(n6539), .ZN(n5429)
         );
  OAI211_X1 U4287 ( .C1(n4993), .C2(n4992), .A(n6648), .B(n4991), .ZN(n5016)
         );
  AND2_X1 U4288 ( .A1(n6500), .A2(n4807), .ZN(n6529) );
  INV_X1 U4289 ( .A(n6551), .ZN(n6578) );
  INV_X1 U4290 ( .A(n6631), .ZN(n6625) );
  INV_X1 U4291 ( .A(n6623), .ZN(n6633) );
  OAI211_X1 U4292 ( .C1(n5074), .C2(n5073), .A(n6648), .B(n5072), .ZN(n5097)
         );
  INV_X1 U4293 ( .A(n5367), .ZN(n5393) );
  AND2_X1 U4294 ( .A1(n5359), .A2(n4735), .ZN(n6640) );
  AND2_X1 U4295 ( .A1(n6639), .A2(n6534), .ZN(n6696) );
  NAND2_X1 U4296 ( .A1(n5033), .A2(n5032), .ZN(n5056) );
  OAI211_X1 U4297 ( .C1(n6651), .C2(n5031), .A(n4880), .B(n6648), .ZN(n4904)
         );
  INV_X1 U4298 ( .A(n6602), .ZN(n6663) );
  NAND2_X1 U4299 ( .A1(n5181), .A2(n5180), .ZN(n5205) );
  AND2_X1 U4300 ( .A1(n6065), .A2(DATAI_19_), .ZN(n6670) );
  AND2_X1 U4301 ( .A1(n6065), .A2(DATAI_30_), .ZN(n6687) );
  INV_X1 U4302 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6704) );
  INV_X1 U4303 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6244) );
  INV_X1 U4304 ( .A(n6361), .ZN(n6350) );
  NAND2_X1 U4305 ( .A1(n4798), .A2(n4797), .ZN(n5889) );
  OR2_X1 U4306 ( .A1(n6402), .A2(n4827), .ZN(n6747) );
  NAND2_X1 U4307 ( .A1(n4860), .A2(n4813), .ZN(n4786) );
  INV_X1 U4308 ( .A(n6743), .ZN(n6385) );
  OR2_X1 U4309 ( .A1(n4662), .A2(n4788), .ZN(n6421) );
  INV_X1 U4310 ( .A(n4491), .ZN(n4492) );
  INV_X1 U4311 ( .A(n6265), .ZN(n6016) );
  NAND2_X1 U4312 ( .A1(n6056), .A2(n6063), .ZN(n6432) );
  AND2_X1 U4313 ( .A1(n3878), .A2(n3877), .ZN(n3879) );
  INV_X1 U4314 ( .A(n6470), .ZN(n6221) );
  INV_X1 U4315 ( .A(n6215), .ZN(n6449) );
  INV_X1 U4316 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5250) );
  AOI211_X2 U4317 ( .C1(n5220), .C2(n5304), .A(n5219), .B(n5218), .ZN(n5258)
         );
  AOI211_X2 U4318 ( .C1(n5307), .C2(n6722), .A(n5306), .B(n5305), .ZN(n6495)
         );
  INV_X1 U4319 ( .A(n6491), .ZN(n5437) );
  AOI22_X1 U4320 ( .A1(n4986), .A2(n4992), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4985), .ZN(n5019) );
  AOI22_X1 U4321 ( .A1(n6504), .A2(n6498), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6506), .ZN(n6533) );
  OR2_X1 U4322 ( .A1(n6589), .A2(n6535), .ZN(n6631) );
  OR2_X1 U4323 ( .A1(n5068), .A2(n6499), .ZN(n5303) );
  AOI22_X1 U4324 ( .A1(n5070), .A2(n5073), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5269), .ZN(n5100) );
  AOI22_X1 U4325 ( .A1(n5361), .A2(n6640), .B1(n5360), .B2(n6546), .ZN(n5396)
         );
  OR2_X1 U4326 ( .A1(n5178), .A2(n4802), .ZN(n6655) );
  OR2_X1 U4327 ( .A1(n5178), .A2(n4965), .ZN(n6685) );
  INV_X1 U4328 ( .A(n6695), .ZN(n5063) );
  OR2_X1 U4329 ( .A1(n4878), .A2(n4807), .ZN(n5173) );
  INV_X1 U4330 ( .A(n6657), .ZN(n6557) );
  INV_X1 U4331 ( .A(n6682), .ZN(n6617) );
  INV_X1 U4332 ( .A(n6697), .ZN(n6630) );
  INV_X1 U4333 ( .A(n6719), .ZN(n6715) );
  OR2_X1 U4334 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6740), .ZN(n4519) );
  AND2_X2 U4335 ( .A1(n4611), .A2(n4758), .ZN(n3448) );
  NOR2_X4 U4336 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4337 ( .A1(n3448), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3272) );
  AND2_X4 U4338 ( .A1(n4613), .A2(n3273), .ZN(n4356) );
  AND2_X4 U4339 ( .A1(n4717), .A2(n4758), .ZN(n3462) );
  AOI22_X1 U4340 ( .A1(n4356), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4341 ( .A1(n3523), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3270) );
  AND2_X2 U4342 ( .A1(n4613), .A2(n4740), .ZN(n3427) );
  AOI22_X1 U4343 ( .A1(n3427), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3492), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4344 ( .A1(n3441), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3493), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3276) );
  AND2_X4 U4345 ( .A1(n4611), .A2(n3274), .ZN(n4375) );
  AOI22_X1 U4346 ( .A1(n4375), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4347 ( .A1(n4375), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4348 ( .A1(n3427), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3492), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U4349 ( .A1(n3448), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4350 ( .A1(n4356), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4351 ( .A1(n3441), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3493), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4352 ( .A1(n3370), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4353 ( .A1(n4349), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3491), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4354 ( .A1(n4349), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3491), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4355 ( .A1(n3427), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3492), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4356 ( .A1(n3441), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3493), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4357 ( .A1(n4375), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3289) );
  NAND4_X1 U4358 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3298)
         );
  AOI22_X1 U4359 ( .A1(n3523), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4360 ( .A1(n3448), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3294) );
  NAND4_X1 U4361 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(n3297)
         );
  OR2_X2 U4362 ( .A1(n3298), .A2(n3297), .ZN(n3385) );
  NAND2_X1 U4363 ( .A1(n3379), .A2(n3386), .ZN(n3397) );
  NAND2_X1 U4364 ( .A1(n3299), .A2(n3397), .ZN(n3337) );
  NAND2_X1 U4365 ( .A1(n3491), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3302) );
  NAND2_X1 U4366 ( .A1(n4375), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4367 ( .A1(n3468), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3300) );
  NAND2_X1 U4368 ( .A1(n4356), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U4369 ( .A1(n3448), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3307)
         );
  NAND2_X1 U4370 ( .A1(n3304), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3306) );
  NAND2_X1 U4371 ( .A1(n3462), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3305)
         );
  NAND2_X1 U4372 ( .A1(n4385), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U4373 ( .A1(n3523), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3311) );
  NAND2_X1 U4374 ( .A1(n3370), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U4375 ( .A1(n3461), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3309)
         );
  NAND2_X1 U4376 ( .A1(n3492), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4377 ( .A1(n3427), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3315)
         );
  NAND2_X1 U4378 ( .A1(n3441), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3314)
         );
  NAND2_X1 U4379 ( .A1(n3493), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3313) );
  INV_X1 U4380 ( .A(n3381), .ZN(n3321) );
  NAND2_X1 U4381 ( .A1(n3321), .A2(n3390), .ZN(n3334) );
  AOI22_X1 U4382 ( .A1(n3493), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4383 ( .A1(n3492), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4384 ( .A1(n3523), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3325) );
  NAND4_X1 U4385 ( .A1(n3327), .A2(n3326), .A3(n3325), .A4(n3324), .ZN(n3333)
         );
  AOI22_X1 U4386 ( .A1(n4349), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3491), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4387 ( .A1(n3427), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4388 ( .A1(n4375), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4389 ( .A1(n4356), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3328) );
  NAND4_X1 U4390 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3332)
         );
  OAI211_X1 U4391 ( .C1(n3321), .C2(n3393), .A(n3334), .B(n3392), .ZN(n3335)
         );
  INV_X1 U4392 ( .A(n3335), .ZN(n3336) );
  NAND2_X1 U4393 ( .A1(n3337), .A2(n3336), .ZN(n3394) );
  NAND2_X1 U4394 ( .A1(n3523), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3341) );
  NAND2_X1 U4395 ( .A1(n4385), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U4396 ( .A1(n3370), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4397 ( .A1(n3461), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3338)
         );
  NAND2_X1 U4398 ( .A1(n3491), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4399 ( .A1(n4375), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4400 ( .A1(n3468), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3342) );
  NAND2_X1 U4401 ( .A1(n3448), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3349)
         );
  NAND2_X1 U4402 ( .A1(n4356), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3348) );
  NAND2_X1 U4403 ( .A1(n3304), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3347) );
  NAND2_X1 U4404 ( .A1(n3462), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3346)
         );
  NAND2_X1 U4405 ( .A1(n3492), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4406 ( .A1(n3427), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3352)
         );
  NAND2_X1 U4407 ( .A1(n3441), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3351)
         );
  NAND2_X1 U4408 ( .A1(n3493), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U4409 ( .A1(n3394), .A2(n4827), .ZN(n3378) );
  AOI22_X1 U4410 ( .A1(n3523), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4411 ( .A1(n3441), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3493), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4412 ( .A1(n4375), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4413 ( .A1(n3448), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4414 ( .A1(n4349), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3491), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4415 ( .A1(n4356), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4416 ( .A1(n4385), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4417 ( .A1(n3427), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3492), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3362) );
  NAND3_X2 U4418 ( .A1(n3094), .A2(n3365), .A3(n3083), .ZN(n3391) );
  AOI22_X1 U4419 ( .A1(n3427), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4385), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4420 ( .A1(n3491), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4375), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4421 ( .A1(n3523), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4422 ( .A1(n4356), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3366) );
  NAND4_X1 U4423 ( .A1(n3369), .A2(n3368), .A3(n3367), .A4(n3366), .ZN(n3376)
         );
  AOI22_X1 U4424 ( .A1(n4349), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4425 ( .A1(n3493), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4426 ( .A1(n3492), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4427 ( .A1(n3448), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3371) );
  NAND4_X1 U4428 ( .A1(n3374), .A2(n3373), .A3(n3372), .A4(n3371), .ZN(n3375)
         );
  NAND2_X1 U4429 ( .A1(n3381), .A2(n3385), .ZN(n3757) );
  INV_X1 U4430 ( .A(n3757), .ZN(n3395) );
  AND2_X4 U4431 ( .A1(n3391), .A2(n3417), .ZN(n5647) );
  NAND2_X1 U4432 ( .A1(n3395), .A2(n5647), .ZN(n3382) );
  XNOR2_X1 U4433 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n3737) );
  NAND2_X1 U4434 ( .A1(n4843), .A2(n3737), .ZN(n3400) );
  NAND2_X1 U4435 ( .A1(n4823), .A2(n3391), .ZN(n3387) );
  NAND2_X1 U4436 ( .A1(n3688), .A2(n3729), .ZN(n3389) );
  NAND3_X1 U4437 ( .A1(n5778), .A2(n5833), .A3(n4584), .ZN(n4606) );
  INV_X1 U4438 ( .A(n3394), .ZN(n3396) );
  INV_X1 U4439 ( .A(n3730), .ZN(n3399) );
  INV_X1 U4440 ( .A(n3397), .ZN(n3398) );
  NAND2_X1 U4441 ( .A1(n4421), .A2(n3400), .ZN(n3401) );
  NAND3_X1 U4442 ( .A1(n3265), .A2(n3760), .A3(n3401), .ZN(n3402) );
  XNOR2_X1 U4443 ( .A(n6541), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5177)
         );
  INV_X1 U4444 ( .A(n3403), .ZN(n3406) );
  INV_X1 U4445 ( .A(n3404), .ZN(n3405) );
  NAND2_X1 U4446 ( .A1(n3406), .A2(n3262), .ZN(n3407) );
  MUX2_X1 U4447 ( .A(n4286), .B(n3755), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3408) );
  INV_X1 U4448 ( .A(n3409), .ZN(n3411) );
  OR2_X1 U4449 ( .A1(n3757), .A2(n4843), .ZN(n3410) );
  NAND2_X1 U4450 ( .A1(n3411), .A2(n3410), .ZN(n3414) );
  NAND2_X1 U4451 ( .A1(n3761), .A2(n3412), .ZN(n3413) );
  NAND2_X1 U4452 ( .A1(n3414), .A2(n3413), .ZN(n3856) );
  INV_X1 U4453 ( .A(n3856), .ZN(n3426) );
  NAND2_X1 U4454 ( .A1(n3121), .A2(n3729), .ZN(n3416) );
  NAND2_X1 U4455 ( .A1(n3416), .A2(n3391), .ZN(n3418) );
  AND3_X2 U4456 ( .A1(n3424), .A2(n3423), .A3(n3422), .ZN(n3425) );
  INV_X1 U4457 ( .A(n3517), .ZN(n3505) );
  AOI22_X1 U4458 ( .A1(n4384), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4459 ( .A1(n4386), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4460 ( .A1(n4376), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4461 ( .A1(n4216), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3428) );
  NAND4_X1 U4462 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .ZN(n3437)
         );
  AOI22_X1 U4463 ( .A1(n4387), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4464 ( .A1(n4375), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4465 ( .A1(n4383), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4466 ( .A1(n4378), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3432) );
  NAND4_X1 U4467 ( .A1(n3435), .A2(n3434), .A3(n3433), .A4(n3432), .ZN(n3436)
         );
  NAND2_X1 U4468 ( .A1(n3505), .A2(n3554), .ZN(n3438) );
  INV_X1 U4469 ( .A(n5527), .ZN(n3439) );
  NAND2_X1 U4470 ( .A1(n3439), .A2(n3554), .ZN(n3456) );
  AOI22_X1 U4471 ( .A1(n4387), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4472 ( .A1(n3467), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4473 ( .A1(n4386), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4474 ( .A1(n4378), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3443) );
  NAND4_X1 U4475 ( .A1(n3446), .A2(n3445), .A3(n3444), .A4(n3443), .ZN(n3454)
         );
  AOI22_X1 U4476 ( .A1(n4384), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4477 ( .A1(n4216), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4479 ( .A1(n4375), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4480 ( .A1(n4388), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3449) );
  NAND4_X1 U4481 ( .A1(n3452), .A2(n3451), .A3(n3450), .A4(n3449), .ZN(n3453)
         );
  OR2_X1 U4482 ( .A1(n3517), .A2(n3651), .ZN(n3455) );
  AOI22_X1 U4483 ( .A1(n4387), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4484 ( .A1(n4383), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4485 ( .A1(n4216), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4486 ( .A1(n4388), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3463) );
  NAND4_X1 U4487 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3474)
         );
  AOI22_X1 U4488 ( .A1(n4384), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4489 ( .A1(n4386), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4490 ( .A1(n4378), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3470) );
  BUF_X1 U4491 ( .A(n3468), .Z(n3518) );
  AOI22_X1 U4492 ( .A1(n4375), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3469) );
  NAND4_X1 U4493 ( .A1(n3472), .A2(n3471), .A3(n3470), .A4(n3469), .ZN(n3473)
         );
  XNOR2_X1 U4494 ( .A(n3651), .B(n3566), .ZN(n3475) );
  NOR2_X1 U4495 ( .A1(n3475), .A2(n3517), .ZN(n3559) );
  INV_X1 U4496 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5238) );
  AOI21_X1 U4497 ( .B1(n4836), .B2(n3651), .A(n4813), .ZN(n3477) );
  NAND2_X1 U4498 ( .A1(n4827), .A2(n3566), .ZN(n3476) );
  OAI211_X1 U4499 ( .C1(n3713), .C2(n5238), .A(n3477), .B(n3476), .ZN(n3561)
         );
  AOI22_X1 U4500 ( .A1(n3559), .A2(n3561), .B1(n3505), .B2(n3651), .ZN(n3478)
         );
  OAI21_X1 U4501 ( .B1(n3552), .B2(n3550), .A(n3551), .ZN(n3480) );
  NAND2_X1 U4502 ( .A1(n3552), .A2(n3550), .ZN(n3479) );
  NAND2_X1 U4503 ( .A1(n3483), .A2(n3482), .ZN(n3485) );
  NAND2_X1 U4504 ( .A1(n3485), .A2(n3484), .ZN(n3510) );
  NAND2_X1 U4505 ( .A1(n3487), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3490) );
  NAND2_X1 U4506 ( .A1(n4984), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5362) );
  MUX2_X1 U4507 ( .A(n5362), .B(n4984), .S(n6541), .Z(n3488) );
  NAND2_X1 U4508 ( .A1(n4726), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U4509 ( .A1(n3488), .A2(n5104), .ZN(n5034) );
  AOI22_X1 U4510 ( .A1(n5034), .A2(n3514), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3513), .ZN(n3489) );
  XNOR2_X1 U4511 ( .A(n3510), .B(n3511), .ZN(n4713) );
  NAND2_X1 U4512 ( .A1(n4713), .A2(n4813), .ZN(n3509) );
  AOI22_X1 U4513 ( .A1(n4387), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3497) );
  AOI22_X1 U4514 ( .A1(n4384), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3496) );
  BUF_X1 U4515 ( .A(n3493), .Z(n4376) );
  AOI22_X1 U4516 ( .A1(n4383), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4517 ( .A1(n4375), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3494) );
  NAND4_X1 U4518 ( .A1(n3497), .A2(n3496), .A3(n3495), .A4(n3494), .ZN(n3503)
         );
  AOI22_X1 U4519 ( .A1(n4216), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3501) );
  AOI22_X1 U4520 ( .A1(n4388), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4521 ( .A1(n4386), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4522 ( .A1(n4378), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3498) );
  NAND4_X1 U4523 ( .A1(n3501), .A2(n3500), .A3(n3499), .A4(n3498), .ZN(n3502)
         );
  INV_X1 U4524 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5257) );
  OAI22_X1 U4525 ( .A1(n5527), .A2(n3574), .B1(n3713), .B2(n5257), .ZN(n3507)
         );
  AND2_X1 U4526 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  XNOR2_X1 U4527 ( .A(n3507), .B(n3506), .ZN(n3508) );
  INV_X1 U4528 ( .A(n3583), .ZN(n3531) );
  INV_X1 U4529 ( .A(n3510), .ZN(n3512) );
  NAND2_X1 U4530 ( .A1(n3512), .A2(n3511), .ZN(n4574) );
  NAND2_X1 U4531 ( .A1(n3487), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3516) );
  NAND2_X1 U4532 ( .A1(n6593), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6629) );
  NAND3_X1 U4533 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5176) );
  INV_X1 U4534 ( .A(n5176), .ZN(n4810) );
  AOI21_X1 U4535 ( .B1(n6629), .B2(n6731), .A(n4808), .ZN(n5110) );
  AOI22_X1 U4536 ( .A1(n5110), .A2(n3514), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3513), .ZN(n3515) );
  XNOR2_X1 U4537 ( .A(n4574), .B(n6544), .ZN(n4734) );
  INV_X1 U4538 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6804) );
  AOI22_X1 U4539 ( .A1(n4387), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4540 ( .A1(n4384), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4541 ( .A1(n4383), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4542 ( .A1(n4375), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3519) );
  NAND4_X1 U4543 ( .A1(n3522), .A2(n3521), .A3(n3520), .A4(n3519), .ZN(n3529)
         );
  AOI22_X1 U4544 ( .A1(n4216), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4545 ( .A1(n4388), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4546 ( .A1(n4386), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4547 ( .A1(n4378), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3524) );
  NAND4_X1 U4548 ( .A1(n3527), .A2(n3526), .A3(n3525), .A4(n3524), .ZN(n3528)
         );
  AOI22_X1 U4549 ( .A1(n3720), .A2(n3585), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3688), .ZN(n3530) );
  AOI22_X1 U4550 ( .A1(n4387), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4551 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n4355), .B1(n4348), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4552 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4386), .B1(n4356), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4553 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4376), .B1(n4350), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3532) );
  NAND4_X1 U4554 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3541)
         );
  AOI22_X1 U4555 ( .A1(n4383), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4556 ( .A1(n4216), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4557 ( .A1(n4384), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4558 ( .A1(n4388), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3536) );
  NAND4_X1 U4559 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3540)
         );
  AOI22_X1 U4560 ( .A1(n3720), .A2(n3608), .B1(INSTQUEUE_REG_0__4__SCAN_IN), 
        .B2(n3688), .ZN(n3543) );
  INV_X1 U4561 ( .A(n3543), .ZN(n3542) );
  NAND2_X1 U4562 ( .A1(n3544), .A2(n3543), .ZN(n3545) );
  NAND2_X1 U4563 ( .A1(n3554), .A2(n3566), .ZN(n3573) );
  NAND2_X1 U4564 ( .A1(n3573), .A2(n3574), .ZN(n3584) );
  NAND2_X1 U4565 ( .A1(n3584), .A2(n3585), .ZN(n3610) );
  XNOR2_X1 U4566 ( .A(n3610), .B(n3608), .ZN(n3547) );
  NAND2_X1 U4567 ( .A1(n3547), .A2(n5521), .ZN(n3548) );
  NAND2_X1 U4568 ( .A1(n3549), .A2(n3548), .ZN(n3592) );
  INV_X1 U4569 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3780) );
  XNOR2_X1 U4570 ( .A(n3592), .B(n3780), .ZN(n4940) );
  XNOR2_X1 U4571 ( .A(n3551), .B(n3550), .ZN(n3553) );
  XNOR2_X1 U4572 ( .A(n3553), .B(n3552), .ZN(n4805) );
  NAND2_X1 U4573 ( .A1(n4805), .A2(n3687), .ZN(n3558) );
  OAI21_X1 U4574 ( .B1(n3554), .B2(n3566), .A(n3573), .ZN(n3555) );
  INV_X1 U4575 ( .A(n5521), .ZN(n3728) );
  OAI211_X1 U4576 ( .C1(n3555), .C2(n3728), .A(n3678), .B(n3391), .ZN(n3556)
         );
  INV_X1 U4577 ( .A(n3556), .ZN(n3557) );
  NAND2_X1 U4578 ( .A1(n3558), .A2(n3557), .ZN(n4701) );
  INV_X1 U4579 ( .A(n3559), .ZN(n3560) );
  XNOR2_X1 U4580 ( .A(n3561), .B(n3560), .ZN(n3562) );
  INV_X1 U4581 ( .A(n4807), .ZN(n3564) );
  NAND2_X1 U4582 ( .A1(n3564), .A2(n3687), .ZN(n3569) );
  INV_X1 U4583 ( .A(n3575), .ZN(n3565) );
  OAI21_X1 U4584 ( .B1(n3728), .B2(n3566), .A(n3565), .ZN(n3567) );
  INV_X1 U4585 ( .A(n3567), .ZN(n3568) );
  NAND2_X1 U4586 ( .A1(n3569), .A2(n3568), .ZN(n6067) );
  NAND2_X1 U4587 ( .A1(n4701), .A2(n4700), .ZN(n4699) );
  INV_X1 U4588 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6454) );
  OR2_X1 U4589 ( .A1(n3570), .A2(n6454), .ZN(n3571) );
  OAI21_X1 U4590 ( .B1(n3574), .B2(n3573), .A(n3584), .ZN(n3576) );
  AOI21_X1 U4591 ( .B1(n3576), .B2(n5521), .A(n3575), .ZN(n3578) );
  NAND2_X1 U4592 ( .A1(n3581), .A2(n3578), .ZN(n3577) );
  NAND2_X1 U4593 ( .A1(n3577), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6423)
         );
  NAND2_X1 U4594 ( .A1(n6426), .A2(n6423), .ZN(n3582) );
  INV_X1 U4595 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3579) );
  AND2_X1 U4596 ( .A1(n3579), .A2(n3578), .ZN(n3580) );
  NAND2_X1 U4597 ( .A1(n3581), .A2(n3580), .ZN(n6424) );
  AND2_X1 U4598 ( .A1(n3582), .A2(n6424), .ZN(n4915) );
  OAI211_X1 U4599 ( .C1(n3585), .C2(n3584), .A(n3610), .B(n5521), .ZN(n3586)
         );
  INV_X1 U4600 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3588) );
  NAND2_X1 U4601 ( .A1(n4915), .A2(n4914), .ZN(n3591) );
  NAND2_X1 U4602 ( .A1(n3589), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3590)
         );
  NAND2_X1 U4603 ( .A1(n3591), .A2(n3590), .ZN(n4941) );
  NAND2_X1 U4604 ( .A1(n3592), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3593)
         );
  AOI22_X1 U4605 ( .A1(n4387), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4606 ( .A1(n4384), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4607 ( .A1(n4383), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4608 ( .A1(n4375), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3594) );
  NAND4_X1 U4609 ( .A1(n3597), .A2(n3596), .A3(n3595), .A4(n3594), .ZN(n3603)
         );
  AOI22_X1 U4610 ( .A1(n4216), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4611 ( .A1(n4388), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4612 ( .A1(n4386), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4613 ( .A1(n4378), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3598) );
  NAND4_X1 U4614 ( .A1(n3601), .A2(n3600), .A3(n3599), .A4(n3598), .ZN(n3602)
         );
  AOI22_X1 U4615 ( .A1(n3720), .A2(n3611), .B1(INSTQUEUE_REG_0__5__SCAN_IN), 
        .B2(n3688), .ZN(n3605) );
  NAND2_X1 U4616 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  NAND2_X1 U4617 ( .A1(n3630), .A2(n3607), .ZN(n3933) );
  INV_X1 U4618 ( .A(n3608), .ZN(n3609) );
  NOR2_X1 U4619 ( .A1(n3610), .A2(n3609), .ZN(n3612) );
  NAND2_X1 U4620 ( .A1(n3612), .A2(n3611), .ZN(n3639) );
  OAI211_X1 U4621 ( .C1(n3612), .C2(n3611), .A(n3639), .B(n5521), .ZN(n3613)
         );
  INV_X1 U4622 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3614) );
  XNOR2_X1 U4623 ( .A(n3615), .B(n3614), .ZN(n4930) );
  NAND2_X1 U4624 ( .A1(n3615), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3616)
         );
  AOI22_X1 U4625 ( .A1(n4384), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4626 ( .A1(n4216), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4627 ( .A1(n4388), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4628 ( .A1(n4378), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3617) );
  NAND4_X1 U4629 ( .A1(n3620), .A2(n3619), .A3(n3618), .A4(n3617), .ZN(n3626)
         );
  AOI22_X1 U4630 ( .A1(n4387), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4631 ( .A1(n4348), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4632 ( .A1(n4355), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4633 ( .A1(n4386), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3621) );
  NAND4_X1 U4634 ( .A1(n3624), .A2(n3623), .A3(n3622), .A4(n3621), .ZN(n3625)
         );
  AOI22_X1 U4635 ( .A1(n3720), .A2(n3640), .B1(n3688), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3629) );
  INV_X1 U4636 ( .A(n3629), .ZN(n3627) );
  NAND2_X1 U4637 ( .A1(n3630), .A2(n3629), .ZN(n3939) );
  NAND3_X1 U4638 ( .A1(n3648), .A2(n3687), .A3(n3939), .ZN(n3633) );
  XNOR2_X1 U4639 ( .A(n3639), .B(n3640), .ZN(n3631) );
  NAND2_X1 U4640 ( .A1(n3631), .A2(n5521), .ZN(n3632) );
  NAND2_X1 U4641 ( .A1(n3633), .A2(n3632), .ZN(n3634) );
  INV_X1 U4642 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3787) );
  XNOR2_X1 U4643 ( .A(n3634), .B(n3787), .ZN(n4956) );
  NAND2_X1 U4644 ( .A1(n4955), .A2(n4956), .ZN(n3636) );
  NAND2_X1 U4645 ( .A1(n3634), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3635)
         );
  NAND2_X1 U4646 ( .A1(n3636), .A2(n3635), .ZN(n5259) );
  INV_X1 U4647 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U4648 ( .A1(n3720), .A2(n3651), .ZN(n3637) );
  OAI21_X1 U4649 ( .B1(n5230), .B2(n3713), .A(n3637), .ZN(n3638) );
  NAND2_X1 U4650 ( .A1(n3888), .A2(n3687), .ZN(n3644) );
  INV_X1 U4651 ( .A(n3639), .ZN(n3641) );
  NAND2_X1 U4652 ( .A1(n3641), .A2(n3640), .ZN(n3653) );
  XNOR2_X1 U4653 ( .A(n3653), .B(n3651), .ZN(n3642) );
  NAND2_X1 U4654 ( .A1(n3642), .A2(n5521), .ZN(n3643) );
  NAND2_X1 U4655 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  XNOR2_X1 U4656 ( .A(n3645), .B(n6930), .ZN(n5260) );
  NAND2_X1 U4657 ( .A1(n5259), .A2(n5260), .ZN(n3647) );
  NAND2_X1 U4658 ( .A1(n3645), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3646)
         );
  INV_X1 U4659 ( .A(n3651), .ZN(n3649) );
  NAND2_X1 U4660 ( .A1(n5521), .A2(n3651), .ZN(n3652) );
  OR2_X1 U4661 ( .A1(n3653), .A2(n3652), .ZN(n3654) );
  INV_X1 U4662 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3793) );
  XNOR2_X1 U4663 ( .A(n3655), .B(n3793), .ZN(n5151) );
  INV_X1 U4664 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7025) );
  NOR2_X1 U4665 ( .A1(n4455), .A2(n7025), .ZN(n3658) );
  NAND2_X1 U4666 ( .A1(n4455), .A2(n7025), .ZN(n3659) );
  INV_X1 U4667 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3661) );
  AND2_X1 U4668 ( .A1(n4455), .A2(n3661), .ZN(n6038) );
  INV_X1 U4669 ( .A(n6038), .ZN(n3660) );
  INV_X1 U4670 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U4671 ( .A1(n4455), .A2(n6206), .ZN(n6026) );
  INV_X1 U4672 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U4673 ( .A1(n4455), .A2(n6019), .ZN(n6018) );
  NOR2_X1 U4674 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3662) );
  OR2_X1 U4675 ( .A1(n4455), .A2(n3662), .ZN(n3663) );
  XNOR2_X1 U4676 ( .A(n4455), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6012)
         );
  INV_X1 U4677 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6189) );
  INV_X1 U4678 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3664) );
  NAND2_X1 U4679 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3666) );
  NAND2_X1 U4680 ( .A1(n4300), .A2(n3666), .ZN(n3667) );
  INV_X1 U4681 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6962) );
  INV_X1 U4682 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6959) );
  INV_X1 U4683 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5972) );
  INV_X1 U4684 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6152) );
  NAND4_X1 U4685 ( .A1(n6962), .A2(n6959), .A3(n5972), .A4(n6152), .ZN(n3668)
         );
  NAND2_X1 U4686 ( .A1(n3080), .A2(n3668), .ZN(n3669) );
  NAND2_X1 U4687 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6759) );
  OAI21_X1 U4688 ( .B1(n6759), .B2(n5972), .A(n4300), .ZN(n3670) );
  NAND2_X1 U4689 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U4690 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6099) );
  NOR2_X1 U4691 ( .A1(n6121), .A2(n6099), .ZN(n5918) );
  AND2_X1 U4692 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3874) );
  NAND2_X1 U4693 ( .A1(n5918), .A2(n3874), .ZN(n3671) );
  INV_X1 U4694 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6855) );
  INV_X1 U4695 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6110) );
  INV_X1 U4696 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6961) );
  INV_X1 U4697 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6094) );
  NAND4_X1 U4698 ( .A1(n6855), .A2(n6110), .A3(n6961), .A4(n6094), .ZN(n3672)
         );
  INV_X1 U4699 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5452) );
  INV_X1 U4700 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U4701 ( .A1(n5452), .A2(n5455), .ZN(n6120) );
  NOR2_X1 U4702 ( .A1(n3672), .A2(n6120), .ZN(n3673) );
  INV_X1 U4703 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5488) );
  XNOR2_X1 U4704 ( .A(n4300), .B(n5488), .ZN(n5481) );
  NAND2_X1 U4705 ( .A1(n4300), .A2(n5488), .ZN(n3676) );
  INV_X1 U4706 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U4707 ( .A1(n5488), .A2(n6085), .ZN(n6080) );
  NOR3_X1 U4708 ( .A1(n5480), .A2(n4300), .A3(n6080), .ZN(n5900) );
  XNOR2_X1 U4709 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3689) );
  INV_X1 U4710 ( .A(n3689), .ZN(n3680) );
  XNOR2_X1 U4711 ( .A(n3680), .B(n3690), .ZN(n3741) );
  AND2_X1 U4712 ( .A1(n3741), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3685) );
  NOR2_X1 U4713 ( .A1(n6541), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3681)
         );
  NOR2_X1 U4714 ( .A1(n3690), .A2(n3681), .ZN(n3683) );
  AOI21_X1 U4715 ( .B1(n3757), .B2(n3683), .A(n4827), .ZN(n3682) );
  NAND2_X1 U4716 ( .A1(n3720), .A2(n3683), .ZN(n3686) );
  NAND2_X1 U4717 ( .A1(n3690), .A2(n3689), .ZN(n3692) );
  NAND2_X1 U4718 ( .A1(n4726), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3691) );
  NAND2_X1 U4719 ( .A1(n3692), .A2(n3691), .ZN(n3699) );
  XNOR2_X1 U4720 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3698) );
  INV_X1 U4721 ( .A(n3698), .ZN(n3693) );
  XNOR2_X1 U4722 ( .A(n3699), .B(n3693), .ZN(n3740) );
  NAND2_X1 U4723 ( .A1(n3720), .A2(n3740), .ZN(n3694) );
  OAI211_X1 U4724 ( .C1(n3740), .C2(n3713), .A(n3694), .B(n3177), .ZN(n3695)
         );
  NAND2_X1 U4725 ( .A1(n3696), .A2(n3695), .ZN(n3705) );
  NAND3_X1 U4726 ( .A1(n3720), .A2(n3697), .A3(n3740), .ZN(n3704) );
  NAND2_X1 U4727 ( .A1(n3699), .A2(n3698), .ZN(n3701) );
  NAND2_X1 U4728 ( .A1(n4984), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3700) );
  XNOR2_X1 U4729 ( .A(n3711), .B(n3708), .ZN(n3742) );
  INV_X1 U4730 ( .A(n3742), .ZN(n3702) );
  AND2_X1 U4731 ( .A1(n3713), .A2(n3702), .ZN(n3703) );
  AOI21_X1 U4732 ( .B1(n3705), .B2(n3704), .A(n3703), .ZN(n3707) );
  NOR2_X1 U4733 ( .A1(n3714), .A2(n3742), .ZN(n3706) );
  NOR2_X1 U4734 ( .A1(n4742), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3709)
         );
  NOR2_X1 U4735 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6482), .ZN(n3712)
         );
  INV_X1 U4736 ( .A(n3715), .ZN(n3717) );
  NAND2_X1 U4737 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4764), .ZN(n3718) );
  NAND2_X1 U4738 ( .A1(n3720), .A2(n3739), .ZN(n3721) );
  INV_X1 U4739 ( .A(n4770), .ZN(n3736) );
  NAND2_X1 U4740 ( .A1(n3121), .A2(n3392), .ZN(n3724) );
  NOR2_X1 U4741 ( .A1(n4612), .A2(n4843), .ZN(n3861) );
  NAND2_X1 U4742 ( .A1(n4612), .A2(n4827), .ZN(n3726) );
  NAND2_X1 U4743 ( .A1(n3725), .A2(n3726), .ZN(n3758) );
  NAND2_X1 U4744 ( .A1(n3729), .A2(n3761), .ZN(n3727) );
  NAND2_X1 U4745 ( .A1(n3728), .A2(n3727), .ZN(n3732) );
  NAND2_X1 U4746 ( .A1(n3729), .A2(n3392), .ZN(n4799) );
  OR2_X1 U4747 ( .A1(n4799), .A2(n3730), .ZN(n3731) );
  NAND2_X1 U4748 ( .A1(n3732), .A2(n3731), .ZN(n3853) );
  INV_X1 U4749 ( .A(n3853), .ZN(n3733) );
  OR2_X1 U4750 ( .A1(n3758), .A2(n3733), .ZN(n3735) );
  INV_X1 U4751 ( .A(n4774), .ZN(n3734) );
  AOI21_X1 U4752 ( .B1(n3736), .B2(n3861), .A(n4569), .ZN(n3754) );
  INV_X1 U4753 ( .A(n3737), .ZN(n3738) );
  NAND2_X1 U4754 ( .A1(n3738), .A2(n4506), .ZN(n5522) );
  INV_X1 U4755 ( .A(n3739), .ZN(n3744) );
  NAND3_X1 U4756 ( .A1(n3742), .A2(n3741), .A3(n3740), .ZN(n3743) );
  NAND2_X1 U4757 ( .A1(n3744), .A2(n3743), .ZN(n3747) );
  INV_X1 U4758 ( .A(n3745), .ZN(n3746) );
  NOR2_X1 U4759 ( .A1(n4773), .A2(READY_N), .ZN(n4565) );
  NAND2_X1 U4760 ( .A1(n5528), .A2(n4565), .ZN(n3752) );
  NAND2_X1 U4761 ( .A1(n4843), .A2(n5522), .ZN(n4429) );
  NAND2_X1 U4762 ( .A1(n4429), .A2(n6706), .ZN(n3749) );
  OAI211_X1 U4763 ( .C1(n4607), .C2(n3749), .A(n3761), .B(n5515), .ZN(n3750)
         );
  NAND2_X1 U4764 ( .A1(n4770), .A2(n3750), .ZN(n3751) );
  MUX2_X1 U4765 ( .A(n3752), .B(n3751), .S(n4823), .Z(n3753) );
  NAND2_X1 U4766 ( .A1(n3754), .A2(n3753), .ZN(n3756) );
  INV_X1 U4767 ( .A(n4780), .ZN(n3759) );
  INV_X1 U4768 ( .A(n5778), .ZN(n4793) );
  NOR2_X1 U4769 ( .A1(n3758), .A2(n4793), .ZN(n4715) );
  OR2_X1 U4770 ( .A1(n3759), .A2(n4715), .ZN(n4769) );
  OAI22_X1 U4771 ( .A1(n3265), .A2(n4836), .B1(n4607), .B2(n4427), .ZN(n3762)
         );
  INV_X1 U4772 ( .A(n3762), .ZN(n3763) );
  NAND2_X1 U4773 ( .A1(n3760), .A2(n3763), .ZN(n3764) );
  NOR2_X1 U4774 ( .A1(n4769), .A2(n3764), .ZN(n3765) );
  NAND2_X1 U4775 ( .A1(n3881), .A2(n6462), .ZN(n3880) );
  OR2_X1 U4776 ( .A1(n4309), .A2(EBX_REG_1__SCAN_IN), .ZN(n3768) );
  NAND2_X1 U4777 ( .A1(n3779), .A2(n6454), .ZN(n3766) );
  OAI211_X1 U4778 ( .C1(n4427), .C2(EBX_REG_1__SCAN_IN), .A(n4317), .B(n3766), 
        .ZN(n3767) );
  NAND2_X1 U4779 ( .A1(n3768), .A2(n3767), .ZN(n3770) );
  NAND2_X1 U4780 ( .A1(n3779), .A2(EBX_REG_0__SCAN_IN), .ZN(n3769) );
  OAI21_X1 U4781 ( .B1(n5647), .B2(EBX_REG_0__SCAN_IN), .A(n3769), .ZN(n4588)
         );
  XNOR2_X1 U4782 ( .A(n3770), .B(n4588), .ZN(n6360) );
  NAND2_X1 U4783 ( .A1(n6360), .A2(n4601), .ZN(n4600) );
  NAND2_X1 U4784 ( .A1(n4600), .A2(n3770), .ZN(n4868) );
  MUX2_X1 U4785 ( .A(n4309), .B(n3779), .S(EBX_REG_2__SCAN_IN), .Z(n3774) );
  INV_X1 U4786 ( .A(n3779), .ZN(n3771) );
  NAND2_X1 U4787 ( .A1(n3771), .A2(n4427), .ZN(n3806) );
  NAND2_X1 U4788 ( .A1(n4427), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3772)
         );
  AND2_X1 U4789 ( .A1(n3806), .A2(n3772), .ZN(n3773) );
  NAND2_X1 U4790 ( .A1(n3774), .A2(n3773), .ZN(n4911) );
  MUX2_X1 U4791 ( .A(n3784), .B(n5647), .S(EBX_REG_3__SCAN_IN), .Z(n3776) );
  NOR2_X1 U4792 ( .A1(n4589), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3775)
         );
  OR2_X1 U4793 ( .A1(n4309), .A2(EBX_REG_4__SCAN_IN), .ZN(n3783) );
  NAND2_X1 U4794 ( .A1(n3779), .A2(n3780), .ZN(n3781) );
  OAI211_X1 U4795 ( .C1(n4427), .C2(EBX_REG_4__SCAN_IN), .A(n4317), .B(n3781), 
        .ZN(n3782) );
  AND2_X1 U4796 ( .A1(n3783), .A2(n3782), .ZN(n4926) );
  MUX2_X1 U4797 ( .A(n3784), .B(n5647), .S(EBX_REG_5__SCAN_IN), .Z(n3786) );
  NOR2_X1 U4798 ( .A1(n4589), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3785)
         );
  NOR2_X1 U4799 ( .A1(n3786), .A2(n3785), .ZN(n4933) );
  OR2_X1 U4800 ( .A1(n4309), .A2(EBX_REG_6__SCAN_IN), .ZN(n3790) );
  NAND2_X1 U4801 ( .A1(n3779), .A2(n3787), .ZN(n3788) );
  OAI211_X1 U4802 ( .C1(n4427), .C2(EBX_REG_6__SCAN_IN), .A(n4317), .B(n3788), 
        .ZN(n3789) );
  MUX2_X1 U4803 ( .A(n3784), .B(n5647), .S(EBX_REG_7__SCAN_IN), .Z(n3791) );
  INV_X1 U4804 ( .A(n3791), .ZN(n3792) );
  NAND2_X1 U4805 ( .A1(n3792), .A2(n3099), .ZN(n5167) );
  OR2_X1 U4806 ( .A1(n4309), .A2(EBX_REG_8__SCAN_IN), .ZN(n3796) );
  NAND2_X1 U4807 ( .A1(n3779), .A2(n3793), .ZN(n3794) );
  OAI211_X1 U4808 ( .C1(n4427), .C2(EBX_REG_8__SCAN_IN), .A(n4317), .B(n3794), 
        .ZN(n3795) );
  MUX2_X1 U4809 ( .A(n3784), .B(n5647), .S(EBX_REG_9__SCAN_IN), .Z(n3798) );
  NOR2_X1 U4810 ( .A1(n4589), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3797)
         );
  NOR2_X1 U4811 ( .A1(n3798), .A2(n3797), .ZN(n5762) );
  NAND2_X1 U4812 ( .A1(n5156), .A2(n5762), .ZN(n5748) );
  MUX2_X1 U4813 ( .A(n4309), .B(n3779), .S(EBX_REG_10__SCAN_IN), .Z(n3801) );
  NAND2_X1 U4814 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4427), .ZN(n3799) );
  AND2_X1 U4815 ( .A1(n3806), .A2(n3799), .ZN(n3800) );
  NAND2_X1 U4816 ( .A1(n4317), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3802) );
  OAI211_X1 U4817 ( .C1(n4427), .C2(EBX_REG_11__SCAN_IN), .A(n3779), .B(n3802), 
        .ZN(n3803) );
  OAI21_X1 U4818 ( .B1(n3836), .B2(EBX_REG_11__SCAN_IN), .A(n3803), .ZN(n5742)
         );
  MUX2_X1 U4819 ( .A(n4309), .B(n3779), .S(EBX_REG_12__SCAN_IN), .Z(n3808) );
  NAND2_X1 U4820 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4427), .ZN(n3805) );
  AND2_X1 U4821 ( .A1(n3806), .A2(n3805), .ZN(n3807) );
  NAND2_X1 U4822 ( .A1(n3808), .A2(n3807), .ZN(n5822) );
  MUX2_X1 U4823 ( .A(n4309), .B(n3779), .S(EBX_REG_14__SCAN_IN), .Z(n3810) );
  NAND2_X1 U4824 ( .A1(n4427), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3809) );
  INV_X1 U4825 ( .A(n5730), .ZN(n3814) );
  INV_X1 U4826 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U4827 ( .A1(n3784), .A2(n6261), .ZN(n3813) );
  NAND2_X1 U4828 ( .A1(n4317), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3811) );
  OAI211_X1 U4829 ( .C1(n4427), .C2(EBX_REG_13__SCAN_IN), .A(n3779), .B(n3811), 
        .ZN(n3812) );
  NAND2_X1 U4830 ( .A1(n4317), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3816) );
  OAI211_X1 U4831 ( .C1(n4427), .C2(EBX_REG_15__SCAN_IN), .A(n3779), .B(n3816), 
        .ZN(n3817) );
  OAI21_X1 U4832 ( .B1(n3836), .B2(EBX_REG_15__SCAN_IN), .A(n3817), .ZN(n5705)
         );
  MUX2_X1 U4833 ( .A(n4309), .B(n3779), .S(EBX_REG_16__SCAN_IN), .Z(n3819) );
  NAND2_X1 U4834 ( .A1(n4427), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U4835 ( .A1(n3819), .A2(n3818), .ZN(n5693) );
  NAND2_X1 U4836 ( .A1(n4317), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3820) );
  OAI211_X1 U4837 ( .C1(n4427), .C2(EBX_REG_17__SCAN_IN), .A(n3779), .B(n3820), 
        .ZN(n3821) );
  OAI21_X1 U4838 ( .B1(n3836), .B2(EBX_REG_17__SCAN_IN), .A(n3821), .ZN(n5681)
         );
  OR2_X1 U4839 ( .A1(n4309), .A2(EBX_REG_19__SCAN_IN), .ZN(n3824) );
  NAND2_X1 U4840 ( .A1(n3779), .A2(n5452), .ZN(n3822) );
  OAI211_X1 U4841 ( .C1(n4427), .C2(EBX_REG_19__SCAN_IN), .A(n4317), .B(n3822), 
        .ZN(n3823) );
  NAND2_X1 U4842 ( .A1(n5646), .A2(n3825), .ZN(n5634) );
  INV_X1 U4843 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5805) );
  AOI22_X1 U4844 ( .A1(n4313), .A2(n5455), .B1(n4601), .B2(n5805), .ZN(n5635)
         );
  NAND2_X1 U4845 ( .A1(n4589), .A2(EBX_REG_18__SCAN_IN), .ZN(n3827) );
  NAND2_X1 U4846 ( .A1(n4427), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3826) );
  NAND2_X1 U4847 ( .A1(n3827), .A2(n3826), .ZN(n5648) );
  MUX2_X1 U4848 ( .A(n5647), .B(n5635), .S(n5648), .Z(n3828) );
  OAI21_X1 U4849 ( .B1(n5805), .B2(n4317), .A(n3828), .ZN(n3829) );
  MUX2_X1 U4850 ( .A(n3784), .B(n5647), .S(EBX_REG_21__SCAN_IN), .Z(n3831) );
  NOR2_X1 U4851 ( .A1(n4589), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3830)
         );
  NOR2_X1 U4852 ( .A1(n3831), .A2(n3830), .ZN(n5629) );
  NAND2_X1 U4853 ( .A1(n5628), .A2(n5629), .ZN(n5609) );
  MUX2_X1 U4854 ( .A(n4309), .B(n3779), .S(EBX_REG_22__SCAN_IN), .Z(n3833) );
  NAND2_X1 U4855 ( .A1(n4427), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4856 ( .A1(n4317), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3834) );
  OAI211_X1 U4857 ( .C1(n4427), .C2(EBX_REG_23__SCAN_IN), .A(n3779), .B(n3834), 
        .ZN(n3835) );
  OAI21_X1 U4858 ( .B1(n3836), .B2(EBX_REG_23__SCAN_IN), .A(n3835), .ZN(n5596)
         );
  MUX2_X1 U4859 ( .A(n3784), .B(n5647), .S(EBX_REG_25__SCAN_IN), .Z(n3837) );
  INV_X1 U4860 ( .A(n3837), .ZN(n3839) );
  NAND2_X1 U4861 ( .A1(n4313), .A2(n5488), .ZN(n3838) );
  NAND2_X1 U4862 ( .A1(n3839), .A2(n3838), .ZN(n5485) );
  MUX2_X1 U4863 ( .A(n4309), .B(n3779), .S(EBX_REG_24__SCAN_IN), .Z(n3841) );
  NAND2_X1 U4864 ( .A1(n4427), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3840) );
  OR2_X1 U4865 ( .A1(n4309), .A2(EBX_REG_26__SCAN_IN), .ZN(n3844) );
  NAND2_X1 U4866 ( .A1(n3779), .A2(n6085), .ZN(n3842) );
  OAI211_X1 U4867 ( .C1(n4427), .C2(EBX_REG_26__SCAN_IN), .A(n4317), .B(n3842), 
        .ZN(n3843) );
  NAND2_X1 U4868 ( .A1(n3844), .A2(n3843), .ZN(n5569) );
  MUX2_X1 U4869 ( .A(n3784), .B(n5647), .S(EBX_REG_27__SCAN_IN), .Z(n3845) );
  INV_X1 U4870 ( .A(n3845), .ZN(n3847) );
  INV_X1 U4871 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U4872 ( .A1(n4313), .A2(n5899), .ZN(n3846) );
  NAND2_X1 U4873 ( .A1(n3847), .A2(n3846), .ZN(n3848) );
  NAND2_X1 U4874 ( .A1(n3098), .A2(n3848), .ZN(n3849) );
  NAND2_X1 U4875 ( .A1(n3091), .A2(n3849), .ZN(n5794) );
  INV_X1 U4876 ( .A(n3868), .ZN(n3852) );
  INV_X1 U4877 ( .A(n4607), .ZN(n3850) );
  OAI21_X1 U4878 ( .B1(n3265), .B2(n3121), .A(n4788), .ZN(n3851) );
  AND2_X1 U4879 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3875) );
  INV_X1 U4880 ( .A(n5515), .ZN(n3889) );
  NAND2_X1 U4881 ( .A1(n5774), .A2(n4823), .ZN(n4570) );
  OAI211_X1 U4882 ( .C1(n4823), .C2(n3889), .A(n3853), .B(n4570), .ZN(n3854)
         );
  INV_X1 U4883 ( .A(n3854), .ZN(n3855) );
  OAI21_X1 U4884 ( .B1(n3725), .B2(n4313), .A(n3855), .ZN(n3857) );
  INV_X1 U4885 ( .A(n4744), .ZN(n3858) );
  NOR2_X1 U4886 ( .A1(n3860), .A2(n3858), .ZN(n3859) );
  NAND2_X1 U4887 ( .A1(n4609), .A2(n3861), .ZN(n4771) );
  AND3_X1 U4888 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n6180) );
  AND2_X1 U4889 ( .A1(n6180), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6162)
         );
  AND2_X1 U4890 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3862) );
  NAND2_X1 U4891 ( .A1(n6162), .A2(n3862), .ZN(n3867) );
  NAND2_X1 U4892 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4917) );
  INV_X1 U4893 ( .A(n4917), .ZN(n6452) );
  NAND3_X1 U4894 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n6452), .ZN(n4934) );
  NAND2_X1 U4895 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3863) );
  NOR2_X1 U4896 ( .A1(n4934), .A2(n3863), .ZN(n5152) );
  INV_X1 U4897 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6930) );
  NOR2_X1 U4898 ( .A1(n6930), .A2(n3793), .ZN(n6217) );
  INV_X1 U4899 ( .A(n6217), .ZN(n6213) );
  NAND2_X1 U4900 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6214) );
  NOR2_X1 U4901 ( .A1(n6213), .A2(n6214), .ZN(n3864) );
  NAND2_X1 U4902 ( .A1(n5152), .A2(n3864), .ZN(n3870) );
  INV_X1 U4903 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6481) );
  OAI21_X1 U4904 ( .B1(n6454), .B2(n6481), .A(n3579), .ZN(n6459) );
  NAND3_X1 U4905 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6459), .ZN(n4957) );
  NOR2_X1 U4906 ( .A1(n3863), .A2(n4957), .ZN(n5160) );
  NAND2_X1 U4907 ( .A1(n3864), .A2(n5160), .ZN(n6159) );
  INV_X1 U4908 ( .A(n6121), .ZN(n3865) );
  INV_X1 U4909 ( .A(n6216), .ZN(n4304) );
  INV_X1 U4910 ( .A(n6759), .ZN(n3866) );
  NOR2_X1 U4911 ( .A1(n3867), .A2(n6159), .ZN(n6115) );
  NAND3_X1 U4912 ( .A1(n3866), .A2(n3865), .A3(n6115), .ZN(n3871) );
  INV_X1 U4913 ( .A(n3867), .ZN(n6143) );
  OR2_X1 U4914 ( .A1(n6181), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3869)
         );
  NAND2_X1 U4915 ( .A1(n3868), .A2(n6218), .ZN(n6480) );
  NAND2_X1 U4916 ( .A1(n3869), .A2(n6480), .ZN(n5154) );
  AOI21_X1 U4917 ( .B1(n4916), .B2(n3870), .A(n5154), .ZN(n6157) );
  OAI21_X1 U4918 ( .B1(n6143), .B2(n5153), .A(n6157), .ZN(n6117) );
  AOI21_X1 U4919 ( .B1(n4304), .B2(n3871), .A(n6117), .ZN(n6107) );
  AOI21_X1 U4920 ( .B1(n6455), .B2(n6460), .A(n3874), .ZN(n3872) );
  INV_X1 U4921 ( .A(REIP_REG_27__SCAN_IN), .ZN(n4548) );
  NOR2_X1 U4922 ( .A1(n6218), .A2(n4548), .ZN(n4291) );
  INV_X1 U4923 ( .A(n6122), .ZN(n6129) );
  INV_X1 U4924 ( .A(n5918), .ZN(n3873) );
  NAND2_X1 U4925 ( .A1(n6092), .A2(n3874), .ZN(n5486) );
  INV_X1 U4926 ( .A(n3875), .ZN(n6081) );
  NOR2_X1 U4927 ( .A1(n5486), .A2(n6081), .ZN(n4302) );
  INV_X1 U4928 ( .A(n4302), .ZN(n6075) );
  NOR2_X1 U4929 ( .A1(n6075), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3876)
         );
  AOI211_X1 U4930 ( .C1(n6071), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n4291), .B(n3876), .ZN(n3877) );
  NAND2_X1 U4931 ( .A1(n3880), .A2(n3879), .ZN(U2991) );
  NAND2_X1 U4932 ( .A1(n3881), .A2(n6428), .ZN(n4295) );
  INV_X1 U4933 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6784) );
  INV_X1 U4934 ( .A(n3911), .ZN(n3882) );
  NAND2_X1 U4935 ( .A1(n3936), .A2(n3884), .ZN(n3883) );
  NAND2_X1 U4936 ( .A1(n3944), .A2(n3883), .ZN(n6305) );
  NAND2_X1 U4937 ( .A1(n5179), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4225) );
  NOR2_X1 U4938 ( .A1(n4225), .A2(n3884), .ZN(n3885) );
  AOI21_X1 U4939 ( .B1(n6305), .B2(n4370), .A(n3885), .ZN(n3886) );
  OAI21_X1 U4940 ( .B1(n4402), .B2(n6784), .A(n3886), .ZN(n3887) );
  AOI22_X1 U4941 ( .A1(n4405), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5179), .ZN(n3891) );
  NAND2_X1 U4942 ( .A1(n3894), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3890) );
  AND2_X1 U4943 ( .A1(n3891), .A2(n3890), .ZN(n3892) );
  NAND2_X1 U4945 ( .A1(n3896), .A2(EAX_REG_0__SCAN_IN), .ZN(n3898) );
  NAND2_X1 U4946 ( .A1(n5179), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3897)
         );
  OAI211_X1 U4947 ( .C1(n3922), .C2(n3895), .A(n3898), .B(n3897), .ZN(n3899)
         );
  AOI21_X1 U4948 ( .B1(n4623), .B2(n4057), .A(n3899), .ZN(n4578) );
  INV_X1 U4949 ( .A(n4578), .ZN(n3900) );
  OR2_X1 U4950 ( .A1(n3900), .A2(n4423), .ZN(n3902) );
  NAND2_X1 U4951 ( .A1(n4807), .A2(n4815), .ZN(n3901) );
  NAND2_X1 U4952 ( .A1(n3901), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4579) );
  OAI21_X1 U4953 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3911), .ZN(n6431) );
  AOI22_X1 U4954 ( .A1(n4404), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4370), 
        .B2(n6431), .ZN(n3905) );
  NAND2_X1 U4955 ( .A1(n4405), .A2(EAX_REG_2__SCAN_IN), .ZN(n3904) );
  OAI211_X1 U4956 ( .C1(n3922), .C2(n3903), .A(n3905), .B(n3904), .ZN(n4907)
         );
  NAND2_X1 U4957 ( .A1(n4908), .A2(n4907), .ZN(n3909) );
  NAND2_X1 U4958 ( .A1(n3906), .A2(n3907), .ZN(n3908) );
  BUF_X2 U4959 ( .A(n3910), .Z(n6727) );
  NAND2_X1 U4960 ( .A1(n6727), .A2(n4057), .ZN(n3919) );
  INV_X1 U4961 ( .A(n3923), .ZN(n3914) );
  INV_X1 U4962 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3912) );
  NAND2_X1 U4963 ( .A1(n3912), .A2(n3911), .ZN(n3913) );
  NAND2_X1 U4964 ( .A1(n3914), .A2(n3913), .ZN(n6351) );
  AOI22_X1 U4965 ( .A1(n6351), .A2(n4370), .B1(n4404), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3916) );
  NAND2_X1 U4966 ( .A1(n4405), .A2(EAX_REG_3__SCAN_IN), .ZN(n3915) );
  OAI211_X1 U4967 ( .C1(n3922), .C2(n4742), .A(n3916), .B(n3915), .ZN(n3917)
         );
  INV_X1 U4968 ( .A(n3917), .ZN(n3918) );
  NAND2_X1 U4969 ( .A1(n5179), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3921)
         );
  NAND2_X1 U4970 ( .A1(n4405), .A2(EAX_REG_4__SCAN_IN), .ZN(n3920) );
  OAI211_X1 U4971 ( .C1(n3922), .C2(n4764), .A(n3921), .B(n3920), .ZN(n3924)
         );
  OAI21_X1 U4972 ( .B1(n3923), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3927), 
        .ZN(n6344) );
  MUX2_X1 U4973 ( .A(n3924), .B(n6344), .S(n4370), .Z(n3925) );
  AOI21_X1 U4974 ( .B1(n3926), .B2(n4057), .A(n3925), .ZN(n4922) );
  AND2_X1 U4975 ( .A1(n3927), .A2(n3930), .ZN(n3928) );
  OR2_X1 U4976 ( .A1(n3928), .A2(n3934), .ZN(n6328) );
  NAND2_X1 U4977 ( .A1(n6328), .A2(n4370), .ZN(n3929) );
  OAI21_X1 U4978 ( .B1(n3930), .B2(n4225), .A(n3929), .ZN(n3931) );
  AOI21_X1 U4979 ( .B1(n3896), .B2(EAX_REG_5__SCAN_IN), .A(n3931), .ZN(n3932)
         );
  OAI21_X1 U4980 ( .B1(n3933), .B2(n3972), .A(n3932), .ZN(n4963) );
  INV_X1 U4981 ( .A(n4962), .ZN(n3941) );
  INV_X1 U4982 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5325) );
  OR2_X1 U4983 ( .A1(n3934), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3935) );
  NAND2_X1 U4984 ( .A1(n3936), .A2(n3935), .ZN(n6309) );
  AOI22_X1 U4985 ( .A1(n6309), .A2(n4370), .B1(n4404), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3937) );
  OAI21_X1 U4986 ( .B1(n4402), .B2(n5325), .A(n3937), .ZN(n3938) );
  AOI21_X1 U4987 ( .B1(n3939), .B2(n4057), .A(n3938), .ZN(n5323) );
  INV_X1 U4988 ( .A(n5323), .ZN(n3940) );
  NAND2_X1 U4989 ( .A1(n3941), .A2(n3940), .ZN(n5164) );
  NAND2_X1 U4990 ( .A1(n3943), .A2(n3942), .ZN(n5166) );
  AOI21_X1 U4991 ( .B1(n6881), .B2(n3944), .A(n3974), .ZN(n6289) );
  OR2_X1 U4992 ( .A1(n6289), .A2(n4423), .ZN(n3959) );
  AOI22_X1 U4993 ( .A1(n4384), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4387), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4994 ( .A1(n4383), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4995 ( .A1(n4386), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4996 ( .A1(n4388), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4997 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3954)
         );
  AOI22_X1 U4998 ( .A1(n4355), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4999 ( .A1(n4216), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U5000 ( .A1(n3440), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U5001 ( .A1(n4378), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3949) );
  NAND4_X1 U5002 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(n3953)
         );
  OAI21_X1 U5003 ( .B1(n3954), .B2(n3953), .A(n4057), .ZN(n3957) );
  NAND2_X1 U5004 ( .A1(n4405), .A2(EAX_REG_8__SCAN_IN), .ZN(n3956) );
  NAND2_X1 U5005 ( .A1(n4404), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3955)
         );
  AOI22_X1 U5006 ( .A1(n4387), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U5007 ( .A1(n4348), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U5008 ( .A1(n4388), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U5009 ( .A1(n4355), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U5010 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3969)
         );
  AOI22_X1 U5011 ( .A1(n4384), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U5012 ( .A1(n4216), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U5013 ( .A1(n4386), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U5014 ( .A1(n4264), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3964) );
  NAND4_X1 U5015 ( .A1(n3967), .A2(n3966), .A3(n3965), .A4(n3964), .ZN(n3968)
         );
  NOR2_X1 U5016 ( .A1(n3969), .A2(n3968), .ZN(n3973) );
  XNOR2_X1 U5017 ( .A(n3974), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U5018 ( .A1(n6050), .A2(n4370), .ZN(n3971) );
  AOI22_X1 U5019 ( .A1(n4405), .A2(EAX_REG_9__SCAN_IN), .B1(n4404), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3970) );
  OAI211_X1 U5020 ( .C1(n3973), .C2(n3972), .A(n3971), .B(n3970), .ZN(n5760)
         );
  XOR2_X1 U5021 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3989), .Z(n6042) );
  AOI22_X1 U5022 ( .A1(n3440), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U5023 ( .A1(n4384), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U5024 ( .A1(n4386), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U5025 ( .A1(n4388), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U5026 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3984)
         );
  AOI22_X1 U5027 ( .A1(n4348), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U5028 ( .A1(n4387), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U5029 ( .A1(n4216), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U5030 ( .A1(n4378), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U5031 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3983)
         );
  OR2_X1 U5032 ( .A1(n3984), .A2(n3983), .ZN(n3985) );
  AOI22_X1 U5033 ( .A1(n4057), .A2(n3985), .B1(n4404), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3987) );
  NAND2_X1 U5034 ( .A1(n3896), .A2(EAX_REG_10__SCAN_IN), .ZN(n3986) );
  OAI211_X1 U5035 ( .C1(n6042), .C2(n4423), .A(n3987), .B(n3986), .ZN(n5747)
         );
  NAND2_X1 U5036 ( .A1(n3990), .A2(n6935), .ZN(n3991) );
  NAND2_X1 U5037 ( .A1(n3991), .A2(n3206), .ZN(n6033) );
  NAND2_X1 U5038 ( .A1(n6033), .A2(n4370), .ZN(n4006) );
  AOI22_X1 U5039 ( .A1(n4387), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U5040 ( .A1(n4383), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U5041 ( .A1(n4216), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U5042 ( .A1(n4388), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3992) );
  NAND4_X1 U5043 ( .A1(n3995), .A2(n3994), .A3(n3993), .A4(n3992), .ZN(n4001)
         );
  AOI22_X1 U5044 ( .A1(n4384), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U5045 ( .A1(n3440), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U5046 ( .A1(n4378), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U5047 ( .A1(n4386), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3996) );
  NAND4_X1 U5048 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(n4000)
         );
  OAI21_X1 U5049 ( .B1(n4001), .B2(n4000), .A(n4057), .ZN(n4004) );
  NAND2_X1 U5050 ( .A1(n4405), .A2(EAX_REG_11__SCAN_IN), .ZN(n4003) );
  NAND2_X1 U5051 ( .A1(n4404), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4002)
         );
  AND3_X1 U5052 ( .A1(n4004), .A2(n4003), .A3(n4002), .ZN(n4005) );
  NAND2_X1 U5053 ( .A1(n4006), .A2(n4005), .ZN(n5737) );
  XOR2_X1 U5054 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n4022), .Z(n6022) );
  AOI22_X1 U5055 ( .A1(n3896), .A2(EAX_REG_12__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5179), .ZN(n4007) );
  MUX2_X1 U5056 ( .A(n6022), .B(n4007), .S(n4423), .Z(n4019) );
  AOI22_X1 U5057 ( .A1(n4348), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U5058 ( .A1(n3459), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U5059 ( .A1(n4384), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U5060 ( .A1(n4388), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4008) );
  NAND4_X1 U5061 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), .ZN(n4017)
         );
  AOI22_X1 U5062 ( .A1(n4387), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5063 ( .A1(n4355), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U5064 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4386), .B1(n4264), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U5065 ( .A1(n4378), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U5066 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4016)
         );
  OAI21_X1 U5067 ( .B1(n4017), .B2(n4016), .A(n4057), .ZN(n4018) );
  NAND2_X1 U5068 ( .A1(n4405), .A2(EAX_REG_13__SCAN_IN), .ZN(n4024) );
  XNOR2_X1 U5069 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n4046), .ZN(n6263)
         );
  AOI22_X1 U5070 ( .A1(n4370), .A2(n6263), .B1(n4404), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4023) );
  NAND2_X1 U5071 ( .A1(n4024), .A2(n4023), .ZN(n5708) );
  AOI22_X1 U5072 ( .A1(n4387), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U5073 ( .A1(n4384), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U5074 ( .A1(n4383), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U5075 ( .A1(n4355), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4025) );
  NAND4_X1 U5076 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(n4034)
         );
  AOI22_X1 U5077 ( .A1(n4216), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5078 ( .A1(n4388), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5079 ( .A1(n4386), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5080 ( .A1(n4378), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U5081 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4033)
         );
  OR2_X1 U5082 ( .A1(n4034), .A2(n4033), .ZN(n4035) );
  NAND2_X1 U5083 ( .A1(n5708), .A2(n5812), .ZN(n4065) );
  INV_X1 U5084 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5881) );
  AOI22_X1 U5085 ( .A1(n4387), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5086 ( .A1(n4386), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U5087 ( .A1(n3459), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5088 ( .A1(n4378), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4036) );
  NAND4_X1 U5089 ( .A1(n4039), .A2(n4038), .A3(n4037), .A4(n4036), .ZN(n4045)
         );
  AOI22_X1 U5090 ( .A1(n4384), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5091 ( .A1(n4348), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5092 ( .A1(n4216), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5093 ( .A1(n3440), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4040) );
  NAND4_X1 U5094 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4044)
         );
  OAI21_X1 U5095 ( .B1(n4045), .B2(n4044), .A(n4057), .ZN(n4048) );
  INV_X1 U5096 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6005) );
  XNOR2_X1 U5097 ( .A(n4060), .B(n6005), .ZN(n6004) );
  AOI22_X1 U5098 ( .A1(n6004), .A2(n4370), .B1(n4404), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4047) );
  OAI211_X1 U5099 ( .C1(n4402), .C2(n5881), .A(n4048), .B(n4047), .ZN(n5720)
         );
  INV_X1 U5100 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6997) );
  AOI22_X1 U5101 ( .A1(n4386), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5102 ( .A1(n4383), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U5103 ( .A1(n4388), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U5104 ( .A1(n4387), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4049) );
  NAND4_X1 U5105 ( .A1(n4052), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(n4059)
         );
  AOI22_X1 U5106 ( .A1(n3440), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5107 ( .A1(n4384), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5108 ( .A1(n3459), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5109 ( .A1(n4378), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4053) );
  NAND4_X1 U5110 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), .ZN(n4058)
         );
  OAI21_X1 U5111 ( .B1(n4059), .B2(n4058), .A(n4057), .ZN(n4063) );
  XNOR2_X1 U5112 ( .A(n4077), .B(n3210), .ZN(n5997) );
  AOI22_X1 U5113 ( .A1(n5997), .A2(n4370), .B1(n4404), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4062) );
  OAI211_X1 U5114 ( .C1(n4402), .C2(n6997), .A(n4063), .B(n4062), .ZN(n5711)
         );
  OAI211_X1 U5115 ( .C1(n5708), .C2(n5812), .A(n5720), .B(n5711), .ZN(n4064)
         );
  AOI22_X1 U5116 ( .A1(n4384), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5117 ( .A1(n4216), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5118 ( .A1(n4387), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5119 ( .A1(n4378), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4066) );
  NAND4_X1 U5120 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4075)
         );
  AOI22_X1 U5121 ( .A1(n3440), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U5122 ( .A1(n4383), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5123 ( .A1(n4386), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5124 ( .A1(n4388), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4070) );
  NAND4_X1 U5125 ( .A1(n4073), .A2(n4072), .A3(n4071), .A4(n4070), .ZN(n4074)
         );
  OR2_X1 U5126 ( .A1(n4075), .A2(n4074), .ZN(n4076) );
  NAND2_X1 U5127 ( .A1(n4397), .A2(n4076), .ZN(n4081) );
  XNOR2_X1 U5128 ( .A(n4082), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5987)
         );
  OAI22_X1 U5129 ( .A1(n5987), .A2(n4423), .B1(n4225), .B2(n3211), .ZN(n4079)
         );
  AOI21_X1 U5130 ( .B1(n4405), .B2(EAX_REG_16__SCAN_IN), .A(n4079), .ZN(n4080)
         );
  NAND2_X1 U5131 ( .A1(n4081), .A2(n4080), .ZN(n5691) );
  NAND2_X1 U5132 ( .A1(n4083), .A2(n5976), .ZN(n4084) );
  AND2_X1 U5133 ( .A1(n4192), .A2(n4084), .ZN(n5974) );
  AOI22_X1 U5134 ( .A1(n4387), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5135 ( .A1(n4384), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5136 ( .A1(n4386), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5137 ( .A1(n4388), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4085) );
  NAND4_X1 U5138 ( .A1(n4088), .A2(n4087), .A3(n4086), .A4(n4085), .ZN(n4094)
         );
  AOI22_X1 U5139 ( .A1(n4383), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5140 ( .A1(n4348), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5141 ( .A1(n4216), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5142 ( .A1(n4378), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4089) );
  NAND4_X1 U5143 ( .A1(n4092), .A2(n4091), .A3(n4090), .A4(n4089), .ZN(n4093)
         );
  OR2_X1 U5144 ( .A1(n4094), .A2(n4093), .ZN(n4096) );
  INV_X1 U5145 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4659) );
  OAI22_X1 U5146 ( .A1(n4402), .A2(n4659), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5976), .ZN(n4095) );
  AOI21_X1 U5147 ( .B1(n4397), .B2(n4096), .A(n4095), .ZN(n4097) );
  MUX2_X1 U5148 ( .A(n5974), .B(n4097), .S(n4423), .Z(n5678) );
  INV_X1 U5149 ( .A(n4100), .ZN(n4101) );
  INV_X1 U5150 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4123) );
  NAND2_X1 U5151 ( .A1(n4101), .A2(n4123), .ZN(n4102) );
  NAND2_X1 U5152 ( .A1(n4223), .A2(n4102), .ZN(n5921) );
  OR2_X1 U5153 ( .A1(n5921), .A2(n4423), .ZN(n4128) );
  AOI22_X1 U5154 ( .A1(n4387), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5155 ( .A1(n4384), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5156 ( .A1(n4383), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5157 ( .A1(n4355), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4103) );
  NAND4_X1 U5158 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4112)
         );
  AOI22_X1 U5159 ( .A1(n4216), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5160 ( .A1(n4388), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5161 ( .A1(n4386), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5162 ( .A1(n4378), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4107) );
  NAND4_X1 U5163 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4111)
         );
  NOR2_X1 U5164 ( .A1(n4112), .A2(n4111), .ZN(n4211) );
  AOI22_X1 U5165 ( .A1(n4376), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5166 ( .A1(n4348), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5167 ( .A1(n4356), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5168 ( .A1(n4216), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4113) );
  NAND4_X1 U5169 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(n4122)
         );
  AOI22_X1 U5170 ( .A1(n4349), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5171 ( .A1(n4384), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5172 ( .A1(n4386), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5173 ( .A1(n4388), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4117) );
  NAND4_X1 U5174 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4121)
         );
  NOR2_X1 U5175 ( .A1(n4122), .A2(n4121), .ZN(n4210) );
  XNOR2_X1 U5176 ( .A(n4211), .B(n4210), .ZN(n4126) );
  AOI21_X1 U5177 ( .B1(n4123), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4124) );
  AOI21_X1 U5178 ( .B1(n3896), .B2(EAX_REG_23__SCAN_IN), .A(n4124), .ZN(n4125)
         );
  OAI21_X1 U5179 ( .B1(n4364), .B2(n4126), .A(n4125), .ZN(n4127) );
  NAND2_X1 U5180 ( .A1(n4128), .A2(n4127), .ZN(n5595) );
  INV_X1 U5181 ( .A(n5595), .ZN(n4191) );
  XNOR2_X1 U5182 ( .A(n4143), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5928)
         );
  AOI22_X1 U5183 ( .A1(n4384), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5184 ( .A1(n4383), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5185 ( .A1(n4386), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5186 ( .A1(n4378), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4129) );
  NAND4_X1 U5187 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4138)
         );
  AOI22_X1 U5188 ( .A1(n4387), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5189 ( .A1(n4216), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5190 ( .A1(n4388), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5191 ( .A1(n4375), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4133) );
  NAND4_X1 U5192 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4137)
         );
  OR2_X1 U5193 ( .A1(n4138), .A2(n4137), .ZN(n4140) );
  INV_X1 U5194 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4653) );
  OAI22_X1 U5195 ( .A1(n4402), .A2(n4653), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5930), .ZN(n4139) );
  AOI21_X1 U5196 ( .B1(n4397), .B2(n4140), .A(n4139), .ZN(n4141) );
  MUX2_X1 U5197 ( .A(n5928), .B(n4141), .S(n4423), .Z(n5607) );
  INV_X1 U5198 ( .A(n5607), .ZN(n4190) );
  NAND2_X1 U5199 ( .A1(n4171), .A2(n5940), .ZN(n4142) );
  AND2_X1 U5200 ( .A1(n4143), .A2(n4142), .ZN(n5942) );
  AOI22_X1 U5201 ( .A1(n4384), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4387), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5202 ( .A1(n4383), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5203 ( .A1(n4388), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5204 ( .A1(n4216), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4144) );
  NAND4_X1 U5205 ( .A1(n4147), .A2(n4146), .A3(n4145), .A4(n4144), .ZN(n4153)
         );
  AOI22_X1 U5206 ( .A1(n4355), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5207 ( .A1(n4386), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5208 ( .A1(n3440), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5209 ( .A1(n4378), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4148) );
  NAND4_X1 U5210 ( .A1(n4151), .A2(n4150), .A3(n4149), .A4(n4148), .ZN(n4152)
         );
  OR2_X1 U5211 ( .A1(n4153), .A2(n4152), .ZN(n4155) );
  INV_X1 U5212 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6748) );
  OAI22_X1 U5213 ( .A1(n4402), .A2(n6748), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5940), .ZN(n4154) );
  AOI21_X1 U5214 ( .B1(n4397), .B2(n4155), .A(n4154), .ZN(n4156) );
  MUX2_X1 U5215 ( .A(n5942), .B(n4156), .S(n4423), .Z(n5621) );
  AOI22_X1 U5216 ( .A1(n4387), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U5217 ( .A1(n4384), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5218 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4383), .B1(n4376), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5219 ( .A1(n4355), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4157) );
  NAND4_X1 U5220 ( .A1(n4160), .A2(n4159), .A3(n4158), .A4(n4157), .ZN(n4166)
         );
  AOI22_X1 U5221 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4216), .B1(n3079), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U5222 ( .A1(n4388), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5223 ( .A1(n4386), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U5224 ( .A1(n4378), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4161) );
  NAND4_X1 U5225 ( .A1(n4164), .A2(n4163), .A3(n4162), .A4(n4161), .ZN(n4165)
         );
  NOR2_X1 U5226 ( .A1(n4166), .A2(n4165), .ZN(n4169) );
  INV_X1 U5227 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n7019) );
  AOI21_X1 U5228 ( .B1(n7019), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4167) );
  AOI21_X1 U5229 ( .B1(n4405), .B2(EAX_REG_20__SCAN_IN), .A(n4167), .ZN(n4168)
         );
  OAI21_X1 U5230 ( .B1(n4364), .B2(n4169), .A(n4168), .ZN(n4173) );
  NAND2_X1 U5231 ( .A1(n4188), .A2(n7019), .ZN(n4170) );
  NAND2_X1 U5232 ( .A1(n4171), .A2(n4170), .ZN(n5949) );
  OR2_X1 U5233 ( .A1(n5949), .A2(n4423), .ZN(n4172) );
  AOI22_X1 U5234 ( .A1(n4387), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5235 ( .A1(n4384), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5236 ( .A1(n3467), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5237 ( .A1(n4264), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4174) );
  NAND4_X1 U5238 ( .A1(n4177), .A2(n4176), .A3(n4175), .A4(n4174), .ZN(n4183)
         );
  AOI22_X1 U5239 ( .A1(n4386), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U5240 ( .A1(n4388), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5241 ( .A1(n3459), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5242 ( .A1(n4383), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4178) );
  NAND4_X1 U5243 ( .A1(n4181), .A2(n4180), .A3(n4179), .A4(n4178), .ZN(n4182)
         );
  NOR2_X1 U5244 ( .A1(n4183), .A2(n4182), .ZN(n4185) );
  AOI22_X1 U5245 ( .A1(n3896), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5179), .ZN(n4184) );
  OAI21_X1 U5246 ( .B1(n4364), .B2(n4185), .A(n4184), .ZN(n4189) );
  NAND2_X1 U5247 ( .A1(n4194), .A2(n4186), .ZN(n4187) );
  NAND2_X1 U5248 ( .A1(n4188), .A2(n4187), .ZN(n5958) );
  MUX2_X1 U5249 ( .A(n4189), .B(n5958), .S(n4370), .Z(n5652) );
  AND2_X1 U5250 ( .A1(n5638), .A2(n5652), .ZN(n5620) );
  NAND2_X1 U5251 ( .A1(n4191), .A2(n5594), .ZN(n4208) );
  NAND2_X1 U5252 ( .A1(n4192), .A2(n3213), .ZN(n4193) );
  AND2_X1 U5253 ( .A1(n4194), .A2(n4193), .ZN(n5967) );
  AOI22_X1 U5254 ( .A1(n4387), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5255 ( .A1(n4383), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4197) );
  AOI22_X1 U5256 ( .A1(n4386), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4196) );
  AOI22_X1 U5257 ( .A1(n4355), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4195) );
  NAND4_X1 U5258 ( .A1(n4198), .A2(n4197), .A3(n4196), .A4(n4195), .ZN(n4204)
         );
  AOI22_X1 U5259 ( .A1(n4384), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U5260 ( .A1(n4376), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U5261 ( .A1(n3304), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U5262 ( .A1(n4388), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4199) );
  NAND4_X1 U5263 ( .A1(n4202), .A2(n4201), .A3(n4200), .A4(n4199), .ZN(n4203)
         );
  OR2_X1 U5264 ( .A1(n4204), .A2(n4203), .ZN(n4206) );
  INV_X1 U5265 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4655) );
  OAI22_X1 U5266 ( .A1(n4402), .A2(n4655), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3213), .ZN(n4205) );
  AOI21_X1 U5267 ( .B1(n4397), .B2(n4206), .A(n4205), .ZN(n4207) );
  MUX2_X1 U5268 ( .A(n5967), .B(n4207), .S(n4423), .Z(n5665) );
  OR2_X1 U5269 ( .A1(n4211), .A2(n4210), .ZN(n4231) );
  AOI22_X1 U5270 ( .A1(n3440), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U5271 ( .A1(n4384), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4387), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U5272 ( .A1(n4348), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U5273 ( .A1(n4355), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4212) );
  NAND4_X1 U5274 ( .A1(n4215), .A2(n4214), .A3(n4213), .A4(n4212), .ZN(n4222)
         );
  INV_X1 U5275 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n7013) );
  AOI22_X1 U5276 ( .A1(n4386), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5277 ( .A1(n3079), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U5278 ( .A1(n4376), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U5279 ( .A1(n4388), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4217) );
  NAND4_X1 U5280 ( .A1(n4220), .A2(n4219), .A3(n4218), .A4(n4217), .ZN(n4221)
         );
  NOR2_X1 U5281 ( .A1(n4222), .A2(n4221), .ZN(n4230) );
  XNOR2_X1 U5282 ( .A(n4231), .B(n4230), .ZN(n4229) );
  NAND2_X1 U5283 ( .A1(n4223), .A2(n6973), .ZN(n4224) );
  NAND2_X1 U5284 ( .A1(n4244), .A2(n4224), .ZN(n5586) );
  NAND2_X1 U5285 ( .A1(n5586), .A2(n4370), .ZN(n4228) );
  NOR2_X1 U5286 ( .A1(n4225), .A2(n6973), .ZN(n4226) );
  AOI21_X1 U5287 ( .B1(n4405), .B2(EAX_REG_24__SCAN_IN), .A(n4226), .ZN(n4227)
         );
  OAI211_X1 U5288 ( .C1(n4229), .C2(n4364), .A(n4228), .B(n4227), .ZN(n5467)
         );
  OR2_X1 U5289 ( .A1(n4231), .A2(n4230), .ZN(n4247) );
  AOI22_X1 U5290 ( .A1(n4387), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U5291 ( .A1(n4376), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4234) );
  AOI22_X1 U5292 ( .A1(n4355), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U5293 ( .A1(n4350), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4232) );
  NAND4_X1 U5294 ( .A1(n4235), .A2(n4234), .A3(n4233), .A4(n4232), .ZN(n4241)
         );
  AOI22_X1 U5295 ( .A1(n4384), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4239) );
  AOI22_X1 U5296 ( .A1(n4383), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4385), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4238) );
  AOI22_X1 U5297 ( .A1(n4388), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U5298 ( .A1(n4386), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4236) );
  NAND4_X1 U5299 ( .A1(n4239), .A2(n4238), .A3(n4237), .A4(n4236), .ZN(n4240)
         );
  NOR2_X1 U5300 ( .A1(n4241), .A2(n4240), .ZN(n4248) );
  XNOR2_X1 U5301 ( .A(n4247), .B(n4248), .ZN(n4243) );
  AOI22_X1 U5302 ( .A1(n4405), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5179), .ZN(n4242) );
  OAI21_X1 U5303 ( .B1(n4243), .B2(n4364), .A(n4242), .ZN(n4246) );
  NAND2_X1 U5304 ( .A1(n4244), .A2(n5578), .ZN(n4245) );
  NAND2_X1 U5305 ( .A1(n4262), .A2(n4245), .ZN(n5577) );
  MUX2_X1 U5306 ( .A(n4246), .B(n5577), .S(n4370), .Z(n5491) );
  NOR2_X1 U5307 ( .A1(n4248), .A2(n4247), .ZN(n4276) );
  AOI22_X1 U5308 ( .A1(n4349), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U5309 ( .A1(n4384), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U5310 ( .A1(n4383), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U5311 ( .A1(n4375), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4249) );
  NAND4_X1 U5312 ( .A1(n4252), .A2(n4251), .A3(n4250), .A4(n4249), .ZN(n4258)
         );
  AOI22_X1 U5313 ( .A1(n4216), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U5314 ( .A1(n4388), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U5315 ( .A1(n4386), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U5316 ( .A1(n4356), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4253) );
  NAND4_X1 U5317 ( .A1(n4256), .A2(n4255), .A3(n4254), .A4(n4253), .ZN(n4257)
         );
  XOR2_X1 U5318 ( .A(n4276), .B(n4275), .Z(n4261) );
  INV_X1 U5319 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4259) );
  OAI22_X1 U5320 ( .A1(n4402), .A2(n4259), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6849), .ZN(n4260) );
  AOI21_X1 U5321 ( .B1(n4261), .B2(n4397), .A(n4260), .ZN(n4263) );
  AOI21_X1 U5322 ( .B1(n6849), .B2(n4262), .A(n4279), .ZN(n5912) );
  MUX2_X1 U5323 ( .A(n4263), .B(n5912), .S(n4370), .Z(n5568) );
  AOI22_X1 U5324 ( .A1(n4383), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4385), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4268) );
  AOI22_X1 U5325 ( .A1(n4384), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U5326 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4388), .B1(n4264), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4266) );
  AOI22_X1 U5327 ( .A1(n4356), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4265) );
  NAND4_X1 U5328 ( .A1(n4268), .A2(n4267), .A3(n4266), .A4(n4265), .ZN(n4274)
         );
  AOI22_X1 U5329 ( .A1(n4349), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U5330 ( .A1(n4375), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U5331 ( .A1(n4376), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4270) );
  AOI22_X1 U5332 ( .A1(n4386), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4269) );
  NAND4_X1 U5333 ( .A1(n4272), .A2(n4271), .A3(n4270), .A4(n4269), .ZN(n4273)
         );
  NOR2_X1 U5334 ( .A1(n4274), .A2(n4273), .ZN(n4330) );
  NAND2_X1 U5335 ( .A1(n4276), .A2(n4275), .ZN(n4329) );
  XNOR2_X1 U5336 ( .A(n4330), .B(n4329), .ZN(n4278) );
  AOI22_X1 U5337 ( .A1(n4405), .A2(EAX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5179), .ZN(n4277) );
  OAI21_X1 U5338 ( .B1(n4278), .B2(n4364), .A(n4277), .ZN(n4282) );
  INV_X1 U5339 ( .A(n4279), .ZN(n4280) );
  INV_X1 U5340 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U5341 ( .A1(n4280), .A2(n5559), .ZN(n4281) );
  NAND2_X1 U5342 ( .A1(n4366), .A2(n4281), .ZN(n5558) );
  MUX2_X1 U5343 ( .A(n4282), .B(n5558), .S(n4370), .Z(n4285) );
  OAI21_X1 U5344 ( .B1(n4283), .B2(n4285), .A(n4284), .ZN(n5845) );
  AND3_X1 U5345 ( .A1(n4813), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U5346 ( .A1(n4286), .A2(n6722), .ZN(n5530) );
  NAND2_X1 U5347 ( .A1(n5530), .A2(n4813), .ZN(n4287) );
  NAND2_X1 U5348 ( .A1(n4813), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4289) );
  NAND2_X1 U5349 ( .A1(n6244), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4288) );
  NAND2_X1 U5350 ( .A1(n4289), .A2(n4288), .ZN(n6063) );
  NOR2_X1 U5351 ( .A1(n6432), .A2(n5558), .ZN(n4290) );
  AOI211_X1 U5352 ( .C1(n6422), .C2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4291), 
        .B(n4290), .ZN(n4292) );
  INV_X1 U5353 ( .A(n4293), .ZN(n4294) );
  NAND2_X1 U5354 ( .A1(n4295), .A2(n4294), .ZN(U2959) );
  NAND2_X1 U5355 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4305) );
  AND2_X1 U5356 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4460) );
  INV_X1 U5357 ( .A(n4298), .ZN(n5479) );
  INV_X1 U5358 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U5359 ( .A1(n5902), .A2(n5899), .ZN(n4299) );
  NOR3_X1 U5360 ( .A1(n4468), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4458) );
  INV_X1 U5361 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4618) );
  INV_X1 U5362 ( .A(n4305), .ZN(n4301) );
  NAND2_X1 U5363 ( .A1(n4302), .A2(n4301), .ZN(n4476) );
  INV_X1 U5364 ( .A(n4460), .ZN(n4303) );
  NOR2_X1 U5365 ( .A1(n4476), .A2(n4303), .ZN(n4306) );
  AOI21_X1 U5366 ( .B1(n4305), .B2(n4304), .A(n6071), .ZN(n4477) );
  MUX2_X1 U5367 ( .A(n4306), .B(n4452), .S(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .Z(n4308) );
  NAND2_X1 U5368 ( .A1(n6457), .A2(REIP_REG_31__SCAN_IN), .ZN(n4412) );
  INV_X1 U5369 ( .A(n4412), .ZN(n4307) );
  OR2_X1 U5370 ( .A1(n4309), .A2(EBX_REG_28__SCAN_IN), .ZN(n4312) );
  NAND2_X1 U5371 ( .A1(n3779), .A2(n5902), .ZN(n4310) );
  OAI211_X1 U5372 ( .C1(n4427), .C2(EBX_REG_28__SCAN_IN), .A(n4317), .B(n4310), 
        .ZN(n4311) );
  INV_X1 U5373 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6978) );
  NAND2_X1 U5374 ( .A1(n4313), .A2(n6978), .ZN(n4318) );
  NAND2_X1 U5375 ( .A1(n4601), .A2(n4314), .ZN(n4315) );
  AND2_X1 U5376 ( .A1(n4318), .A2(n4315), .ZN(n4316) );
  INV_X1 U5377 ( .A(n4318), .ZN(n4319) );
  MUX2_X1 U5378 ( .A(n4319), .B(EBX_REG_29__SCAN_IN), .S(n5647), .Z(n4320) );
  AOI21_X1 U5379 ( .B1(n3784), .B2(n4314), .A(n4320), .ZN(n4475) );
  NAND2_X1 U5380 ( .A1(n5547), .A2(n4475), .ZN(n4474) );
  INV_X1 U5381 ( .A(n4474), .ZN(n4324) );
  NAND2_X1 U5382 ( .A1(n4589), .A2(EBX_REG_30__SCAN_IN), .ZN(n4322) );
  NAND2_X1 U5383 ( .A1(n4427), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4321) );
  NAND2_X1 U5384 ( .A1(n4322), .A2(n4321), .ZN(n4415) );
  INV_X1 U5385 ( .A(n4415), .ZN(n4323) );
  OAI22_X1 U5386 ( .A1(n4589), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4427), .B2(EBX_REG_31__SCAN_IN), .ZN(n4326) );
  NOR2_X1 U5387 ( .A1(n4330), .A2(n4329), .ZN(n4347) );
  AOI22_X1 U5388 ( .A1(n4349), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4334) );
  AOI22_X1 U5389 ( .A1(n4384), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4333) );
  AOI22_X1 U5390 ( .A1(n4383), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4332) );
  AOI22_X1 U5391 ( .A1(n4375), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4331) );
  NAND4_X1 U5392 ( .A1(n4334), .A2(n4333), .A3(n4332), .A4(n4331), .ZN(n4340)
         );
  AOI22_X1 U5393 ( .A1(n4216), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4338) );
  AOI22_X1 U5394 ( .A1(n4388), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4337) );
  AOI22_X1 U5395 ( .A1(n4386), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4336) );
  AOI22_X1 U5396 ( .A1(n4356), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4335) );
  NAND4_X1 U5397 ( .A1(n4338), .A2(n4337), .A3(n4336), .A4(n4335), .ZN(n4339)
         );
  OR2_X1 U5398 ( .A1(n4340), .A2(n4339), .ZN(n4346) );
  XOR2_X1 U5399 ( .A(n4347), .B(n4346), .Z(n4343) );
  INV_X1 U5400 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4341) );
  INV_X1 U5401 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5905) );
  OAI22_X1 U5402 ( .A1(n4402), .A2(n4341), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5905), .ZN(n4342) );
  AOI21_X1 U5403 ( .B1(n4343), .B2(n4397), .A(n4342), .ZN(n4344) );
  XNOR2_X1 U5404 ( .A(n4366), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5907)
         );
  MUX2_X1 U5405 ( .A(n4344), .B(n5907), .S(n4370), .Z(n5546) );
  NOR2_X2 U5406 ( .A1(n4345), .A2(n5546), .ZN(n4485) );
  NAND2_X1 U5407 ( .A1(n4347), .A2(n4346), .ZN(n4373) );
  AOI22_X1 U5408 ( .A1(n4349), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4348), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U5409 ( .A1(n4383), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3079), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4353) );
  AOI22_X1 U5410 ( .A1(n4386), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4352) );
  AOI22_X1 U5411 ( .A1(n4216), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4351) );
  NAND4_X1 U5412 ( .A1(n4354), .A2(n4353), .A3(n4352), .A4(n4351), .ZN(n4362)
         );
  AOI22_X1 U5413 ( .A1(n4384), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4360) );
  AOI22_X1 U5414 ( .A1(n4388), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4359) );
  AOI22_X1 U5415 ( .A1(n3440), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U5416 ( .A1(n4356), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4357) );
  NAND4_X1 U5417 ( .A1(n4360), .A2(n4359), .A3(n4358), .A4(n4357), .ZN(n4361)
         );
  NOR2_X1 U5418 ( .A1(n4362), .A2(n4361), .ZN(n4374) );
  XNOR2_X1 U5419 ( .A(n4373), .B(n4374), .ZN(n4365) );
  AOI22_X1 U5420 ( .A1(n4405), .A2(EAX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n5179), .ZN(n4363) );
  OAI21_X1 U5421 ( .B1(n4365), .B2(n4364), .A(n4363), .ZN(n4371) );
  INV_X1 U5422 ( .A(n4366), .ZN(n4367) );
  NAND2_X1 U5423 ( .A1(n4367), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4368)
         );
  INV_X1 U5424 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U5425 ( .A1(n4368), .A2(n5537), .ZN(n4369) );
  NAND2_X1 U5426 ( .A1(n4408), .A2(n4369), .ZN(n5536) );
  MUX2_X1 U5427 ( .A(n4371), .B(n5536), .S(n4370), .Z(n4487) );
  NAND2_X1 U5428 ( .A1(n4485), .A2(n4487), .ZN(n4486) );
  INV_X1 U5429 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4372) );
  XNOR2_X1 U5430 ( .A(n4408), .B(n4372), .ZN(n5895) );
  INV_X1 U5431 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4401) );
  NOR2_X1 U5432 ( .A1(n4374), .A2(n4373), .ZN(n4396) );
  AOI22_X1 U5433 ( .A1(n3440), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4375), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U5434 ( .A1(n3467), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4376), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4381) );
  AOI22_X1 U5435 ( .A1(n3079), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4380) );
  AOI22_X1 U5436 ( .A1(n4378), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4379) );
  NAND4_X1 U5437 ( .A1(n4382), .A2(n4381), .A3(n4380), .A4(n4379), .ZN(n4394)
         );
  AOI22_X1 U5438 ( .A1(n4384), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U5439 ( .A1(n4386), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4385), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U5440 ( .A1(n4387), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4390) );
  AOI22_X1 U5441 ( .A1(n4388), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4389) );
  NAND4_X1 U5442 ( .A1(n4392), .A2(n4391), .A3(n4390), .A4(n4389), .ZN(n4393)
         );
  NOR2_X1 U5443 ( .A1(n4394), .A2(n4393), .ZN(n4395) );
  XNOR2_X1 U5444 ( .A(n4396), .B(n4395), .ZN(n4398) );
  NAND2_X1 U5445 ( .A1(n4398), .A2(n4397), .ZN(n4400) );
  OAI21_X1 U5446 ( .B1(n6244), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5179), 
        .ZN(n4399) );
  OAI211_X1 U5447 ( .C1(n4402), .C2(n4401), .A(n4400), .B(n4399), .ZN(n4403)
         );
  OAI21_X1 U5448 ( .B1(n5895), .B2(n4423), .A(n4403), .ZN(n4446) );
  NOR2_X2 U5449 ( .A1(n4486), .A2(n4446), .ZN(n4407) );
  AOI22_X1 U5450 ( .A1(n4405), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4404), .ZN(n4406) );
  INV_X1 U5451 ( .A(n4408), .ZN(n4409) );
  INV_X1 U5452 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4410) );
  NAND2_X1 U5453 ( .A1(n6422), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4411)
         );
  OAI211_X1 U5454 ( .C1(n6432), .C2(n4447), .A(n4412), .B(n4411), .ZN(n4413)
         );
  AOI21_X1 U5455 ( .B1(n5514), .B2(n6065), .A(n4413), .ZN(n4414) );
  AOI21_X1 U5456 ( .B1(n4417), .B2(n5547), .A(n4415), .ZN(n4420) );
  INV_X1 U5457 ( .A(n5547), .ZN(n4416) );
  AOI21_X1 U5458 ( .B1(n4416), .B2(n5647), .A(n4323), .ZN(n4418) );
  INV_X1 U5459 ( .A(n5500), .ZN(n4454) );
  INV_X1 U5460 ( .A(n4421), .ZN(n4554) );
  NAND3_X1 U5461 ( .A1(n4774), .A2(n5533), .A3(n4552), .ZN(n4558) );
  NAND2_X1 U5462 ( .A1(n4813), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4422) );
  NOR2_X1 U5463 ( .A1(n4423), .A2(n4422), .ZN(n6714) );
  NOR2_X1 U5464 ( .A1(n5525), .A2(n5217), .ZN(n4424) );
  NAND2_X1 U5465 ( .A1(n6706), .A2(n6244), .ZN(n4432) );
  NAND2_X1 U5466 ( .A1(n4432), .A2(EBX_REG_31__SCAN_IN), .ZN(n4426) );
  NOR2_X1 U5467 ( .A1(n4427), .A2(n4426), .ZN(n4428) );
  NOR2_X1 U5468 ( .A1(n4827), .A2(n4432), .ZN(n4430) );
  AND2_X1 U5469 ( .A1(n4430), .A2(n4429), .ZN(n4431) );
  INV_X1 U5470 ( .A(REIP_REG_17__SCAN_IN), .ZN(n4512) );
  INV_X1 U5471 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5984) );
  INV_X1 U5472 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6199) );
  INV_X1 U5473 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7009) );
  INV_X1 U5474 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6319) );
  INV_X1 U5475 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6331) );
  NAND3_X1 U5476 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6335) );
  OR2_X1 U5477 ( .A1(n6331), .A2(n6335), .ZN(n6320) );
  NOR2_X1 U5478 ( .A1(n6319), .A2(n6320), .ZN(n6302) );
  NAND2_X1 U5479 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6302), .ZN(n6296) );
  NOR2_X1 U5480 ( .A1(n7009), .A2(n6296), .ZN(n5754) );
  NAND2_X1 U5481 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5754), .ZN(n5753) );
  NAND2_X1 U5482 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n5755) );
  NOR2_X1 U5483 ( .A1(n5753), .A2(n5755), .ZN(n5739) );
  NAND2_X1 U5484 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5739), .ZN(n6266) );
  NOR2_X1 U5485 ( .A1(n6199), .A2(n6266), .ZN(n6268) );
  AND2_X1 U5486 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6268), .ZN(n5724) );
  NAND2_X1 U5487 ( .A1(n5701), .A2(REIP_REG_15__SCAN_IN), .ZN(n5697) );
  NOR3_X1 U5488 ( .A1(n4512), .A2(n5984), .A3(n5697), .ZN(n5670) );
  NAND3_X1 U5489 ( .A1(n6359), .A2(REIP_REG_18__SCAN_IN), .A3(n5670), .ZN(
        n5657) );
  INV_X1 U5490 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5948) );
  INV_X1 U5491 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5957) );
  NOR3_X1 U5492 ( .A1(n5657), .A2(n5948), .A3(n5957), .ZN(n5632) );
  AND3_X1 U5493 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5494 ( .A1(n5632), .A2(n4436), .ZN(n5590) );
  INV_X1 U5495 ( .A(REIP_REG_24__SCAN_IN), .ZN(n4544) );
  INV_X1 U5496 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7040) );
  NOR3_X1 U5497 ( .A1(n5590), .A2(n4544), .A3(n7040), .ZN(n5572) );
  NAND2_X1 U5498 ( .A1(n5572), .A2(REIP_REG_26__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U5499 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4439) );
  NOR2_X1 U5500 ( .A1(n5563), .A2(n4439), .ZN(n5439) );
  INV_X1 U5501 ( .A(n5439), .ZN(n5541) );
  INV_X1 U5502 ( .A(REIP_REG_29__SCAN_IN), .ZN(n4551) );
  NOR3_X1 U5503 ( .A1(n5541), .A2(REIP_REG_30__SCAN_IN), .A3(n4551), .ZN(n4445) );
  INV_X1 U5504 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5499) );
  INV_X1 U5505 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U5506 ( .A1(n4432), .A2(n5790), .ZN(n4434) );
  OR2_X1 U5507 ( .A1(n5522), .A2(n4432), .ZN(n4787) );
  AND2_X1 U5508 ( .A1(n5521), .A2(n4787), .ZN(n5442) );
  INV_X1 U5509 ( .A(n5442), .ZN(n4433) );
  OAI21_X1 U5510 ( .B1(n4827), .B2(n4434), .A(n4433), .ZN(n4435) );
  NAND2_X1 U5511 ( .A1(n6321), .A2(n6373), .ZN(n6329) );
  INV_X1 U5512 ( .A(n4436), .ZN(n4437) );
  INV_X1 U5513 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U5514 ( .A1(n5670), .A2(n6373), .ZN(n5666) );
  NOR3_X1 U5515 ( .A1(n5957), .A2(n5669), .A3(n5666), .ZN(n5656) );
  NAND2_X1 U5516 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5656), .ZN(n5625) );
  NOR2_X1 U5517 ( .A1(n4437), .A2(n5625), .ZN(n5580) );
  NAND4_X1 U5518 ( .A1(n5580), .A2(REIP_REG_24__SCAN_IN), .A3(
        REIP_REG_26__SCAN_IN), .A4(REIP_REG_25__SCAN_IN), .ZN(n4438) );
  NAND2_X1 U5519 ( .A1(n6329), .A2(n4438), .ZN(n5557) );
  NAND2_X1 U5520 ( .A1(n6359), .A2(n4439), .ZN(n4440) );
  NAND2_X1 U5521 ( .A1(n5557), .A2(n4440), .ZN(n5550) );
  OR2_X1 U5522 ( .A1(n5550), .A2(n4551), .ZN(n5441) );
  NAND3_X1 U5523 ( .A1(n5441), .A2(REIP_REG_30__SCAN_IN), .A3(n6329), .ZN(
        n4443) );
  INV_X1 U5524 ( .A(n5895), .ZN(n4441) );
  AOI22_X1 U5525 ( .A1(n6364), .A2(n4441), .B1(n6358), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4442) );
  OAI211_X1 U5526 ( .C1(n5499), .C2(n6306), .A(n4443), .B(n4442), .ZN(n4444)
         );
  AOI211_X1 U5527 ( .C1(n4454), .C2(n6361), .A(n4445), .B(n4444), .ZN(n4451)
         );
  XNOR2_X1 U5528 ( .A(n4486), .B(n4446), .ZN(n5498) );
  INV_X1 U5529 ( .A(n5498), .ZN(n4449) );
  NAND2_X1 U5530 ( .A1(n4449), .A2(n6311), .ZN(n4450) );
  NAND2_X1 U5531 ( .A1(n4451), .A2(n4450), .ZN(U2797) );
  INV_X1 U5532 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5440) );
  NOR2_X1 U5533 ( .A1(n6218), .A2(n5440), .ZN(n5893) );
  NOR2_X1 U5534 ( .A1(n4476), .A2(n6978), .ZN(n4453) );
  INV_X1 U5535 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6837) );
  NOR2_X1 U5536 ( .A1(n6837), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4459)
         );
  NAND3_X1 U5537 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A3(INSTADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n4461) );
  NOR4_X1 U5538 ( .A1(n3080), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6978), 
        .A4(n4461), .ZN(n4456) );
  OAI21_X1 U5539 ( .B1(n4459), .B2(n4456), .A(n5911), .ZN(n4466) );
  INV_X1 U5540 ( .A(n4457), .ZN(n4470) );
  OAI21_X1 U5541 ( .B1(n4458), .B2(n4460), .A(n4470), .ZN(n4465) );
  NAND2_X1 U5542 ( .A1(n4468), .A2(n4459), .ZN(n4463) );
  OAI21_X1 U5543 ( .B1(n3080), .B2(n4461), .A(n4460), .ZN(n4462) );
  AND2_X1 U5544 ( .A1(n4463), .A2(n4462), .ZN(n4464) );
  NAND3_X1 U5545 ( .A1(n4466), .A2(n4465), .A3(n4464), .ZN(n5897) );
  NAND2_X1 U5546 ( .A1(n5897), .A2(n6462), .ZN(n4467) );
  INV_X1 U5547 ( .A(n4468), .ZN(n4469) );
  XNOR2_X2 U5548 ( .A(n4473), .B(n6978), .ZN(n4484) );
  NAND2_X1 U5549 ( .A1(n4484), .A2(n6462), .ZN(n4483) );
  OAI21_X1 U5550 ( .B1(n5547), .B2(n4475), .A(n4474), .ZN(n5792) );
  INV_X1 U5551 ( .A(n4476), .ZN(n4479) );
  NOR2_X1 U5552 ( .A1(n6218), .A2(n4551), .ZN(n4489) );
  NOR2_X1 U5553 ( .A1(n4477), .A2(n6978), .ZN(n4478) );
  AOI211_X1 U5554 ( .C1(n4479), .C2(n6978), .A(n4489), .B(n4478), .ZN(n4480)
         );
  NAND2_X1 U5555 ( .A1(n4483), .A2(n4482), .ZN(U2989) );
  NAND2_X1 U5556 ( .A1(n4484), .A2(n6428), .ZN(n4493) );
  OAI21_X1 U5557 ( .B1(n5545), .B2(n4487), .A(n4486), .ZN(n5839) );
  NOR2_X1 U5558 ( .A1(n6432), .A2(n5536), .ZN(n4488) );
  AOI211_X1 U5559 ( .C1(n6422), .C2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4489), 
        .B(n4488), .ZN(n4490) );
  NAND2_X1 U5560 ( .A1(n4493), .A2(n4492), .ZN(U2957) );
  INV_X1 U5561 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4496) );
  INV_X1 U5562 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4514) );
  NOR2_X1 U5563 ( .A1(n4506), .A2(n4514), .ZN(n4498) );
  AND2_X1 U5564 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n4515) );
  NAND2_X1 U5565 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4494) );
  OAI21_X1 U5566 ( .B1(n4498), .B2(n4515), .A(n4494), .ZN(n4495) );
  OAI211_X1 U5567 ( .C1(n6706), .C2(n4496), .A(n4495), .B(n5522), .ZN(U3182)
         );
  INV_X1 U5568 ( .A(NA_N), .ZN(n4499) );
  AOI221_X1 U5569 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n4499), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n4513) );
  AOI221_X1 U5570 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6706), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4497) );
  AOI221_X1 U5571 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n4497), .C2(HOLD), .A(n4506), .ZN(n4501) );
  AOI22_X1 U5572 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .B1(
        STATE_REG_1__SCAN_IN), .B2(READY_N), .ZN(n4518) );
  AND2_X1 U5573 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n4517) );
  AOI21_X1 U5574 ( .B1(n4499), .B2(n4498), .A(n4517), .ZN(n4500) );
  OAI22_X1 U5575 ( .A1(n4513), .A2(n4501), .B1(n4518), .B2(n4500), .ZN(U3183)
         );
  AND2_X1 U5576 ( .A1(n4860), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5024) );
  INV_X1 U5577 ( .A(n5024), .ZN(n4791) );
  NAND2_X1 U5578 ( .A1(n5179), .A2(READY_N), .ZN(n5021) );
  NOR2_X1 U5579 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6703) );
  INV_X1 U5580 ( .A(n6703), .ZN(n4502) );
  NAND4_X1 U5581 ( .A1(n4791), .A2(n5525), .A3(n5021), .A4(n4502), .ZN(n4505)
         );
  INV_X1 U5582 ( .A(n4503), .ZN(n4504) );
  NAND2_X1 U5583 ( .A1(n4505), .A2(n4504), .ZN(U3150) );
  INV_X1 U5584 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4510) );
  INV_X1 U5585 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4507) );
  NAND2_X1 U5586 ( .A1(n4507), .A2(STATE_REG_1__SCAN_IN), .ZN(n4508) );
  NAND2_X1 U5587 ( .A1(STATE_REG_0__SCAN_IN), .A2(n4508), .ZN(n4509) );
  INV_X2 U5588 ( .A(n6742), .ZN(n6740) );
  OAI21_X1 U5589 ( .B1(n6742), .B2(n4510), .A(n6715), .ZN(U2789) );
  INV_X1 U5590 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6269) );
  INV_X1 U5591 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6802) );
  OAI222_X1 U5592 ( .A1(n4541), .A2(n6199), .B1(n4519), .B2(n6269), .C1(n6742), 
        .C2(n6802), .ZN(U3195) );
  INV_X1 U5593 ( .A(REIP_REG_14__SCAN_IN), .ZN(n4511) );
  INV_X1 U5594 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n7010) );
  INV_X1 U5595 ( .A(REIP_REG_15__SCAN_IN), .ZN(n4535) );
  OAI222_X1 U5596 ( .A1(n4541), .A2(n4511), .B1(n6742), .B2(n7010), .C1(n4535), 
        .C2(n4519), .ZN(U3197) );
  INV_X1 U5597 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6964) );
  INV_X1 U5598 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6977) );
  OAI222_X1 U5599 ( .A1(n4541), .A2(n6964), .B1(n6742), .B2(n6977), .C1(n4551), 
        .C2(n4519), .ZN(U3211) );
  INV_X1 U5600 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6822) );
  OAI222_X1 U5601 ( .A1(n4541), .A2(n5669), .B1(n6742), .B2(n6822), .C1(n4519), 
        .C2(n5957), .ZN(U3201) );
  INV_X1 U5602 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6911) );
  OAI222_X1 U5603 ( .A1(n4541), .A2(n4512), .B1(n6742), .B2(n6911), .C1(n5669), 
        .C2(n4519), .ZN(U3200) );
  INV_X1 U5604 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6846) );
  INV_X1 U5605 ( .A(REIP_REG_26__SCAN_IN), .ZN(n4546) );
  OAI222_X1 U5606 ( .A1(n4541), .A2(n7040), .B1(n6742), .B2(n6846), .C1(n4546), 
        .C2(n4519), .ZN(U3208) );
  AOI221_X1 U5607 ( .B1(n4515), .B2(n6740), .C1(n4514), .C2(n6740), .A(n4513), 
        .ZN(n4516) );
  OAI21_X1 U5608 ( .B1(n4518), .B2(n4517), .A(n4516), .ZN(U3181) );
  INV_X1 U5609 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6301) );
  INV_X1 U5610 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6900) );
  OAI222_X1 U5611 ( .A1(n4519), .A2(n7009), .B1(n4541), .B2(n6301), .C1(n6742), 
        .C2(n6900), .ZN(U3189) );
  INV_X1 U5612 ( .A(n4519), .ZN(n4549) );
  AOI22_X1 U5613 ( .A1(n4549), .A2(REIP_REG_23__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_21__SCAN_IN), .ZN(n4520) );
  OAI21_X1 U5614 ( .B1(n6956), .B2(n4541), .A(n4520), .ZN(U3205) );
  INV_X1 U5615 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6996) );
  AOI22_X1 U5616 ( .A1(n4549), .A2(REIP_REG_2__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_0__SCAN_IN), .ZN(n4521) );
  OAI21_X1 U5617 ( .B1(n6996), .B2(n4541), .A(n4521), .ZN(U3184) );
  INV_X1 U5618 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6989) );
  AOI22_X1 U5619 ( .A1(n4549), .A2(REIP_REG_3__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_1__SCAN_IN), .ZN(n4522) );
  OAI21_X1 U5620 ( .B1(n6989), .B2(n4541), .A(n4522), .ZN(U3185) );
  INV_X1 U5621 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7022) );
  AOI22_X1 U5622 ( .A1(n4549), .A2(REIP_REG_4__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_2__SCAN_IN), .ZN(n4523) );
  OAI21_X1 U5623 ( .B1(n7022), .B2(n4541), .A(n4523), .ZN(U3186) );
  AOI22_X1 U5624 ( .A1(n4549), .A2(REIP_REG_5__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_3__SCAN_IN), .ZN(n4524) );
  OAI21_X1 U5625 ( .B1(n6331), .B2(n4541), .A(n4524), .ZN(U3187) );
  AOI22_X1 U5626 ( .A1(n4549), .A2(REIP_REG_6__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_4__SCAN_IN), .ZN(n4525) );
  OAI21_X1 U5627 ( .B1(n6319), .B2(n4541), .A(n4525), .ZN(U3188) );
  AOI22_X1 U5628 ( .A1(n4549), .A2(REIP_REG_8__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_6__SCAN_IN), .ZN(n4526) );
  OAI21_X1 U5629 ( .B1(n7009), .B2(n4541), .A(n4526), .ZN(U3190) );
  INV_X1 U5630 ( .A(REIP_REG_8__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5631 ( .A1(n4549), .A2(REIP_REG_9__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_7__SCAN_IN), .ZN(n4527) );
  OAI21_X1 U5632 ( .B1(n4528), .B2(n4541), .A(n4527), .ZN(U3191) );
  AOI22_X1 U5633 ( .A1(n4549), .A2(REIP_REG_10__SCAN_IN), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6740), .ZN(n4529) );
  OAI21_X1 U5634 ( .B1(n6838), .B2(n4541), .A(n4529), .ZN(U3192) );
  INV_X1 U5635 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6219) );
  AOI22_X1 U5636 ( .A1(n4549), .A2(REIP_REG_11__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_9__SCAN_IN), .ZN(n4530) );
  OAI21_X1 U5637 ( .B1(n6219), .B2(n4541), .A(n4530), .ZN(U3193) );
  INV_X1 U5638 ( .A(REIP_REG_11__SCAN_IN), .ZN(n4532) );
  AOI22_X1 U5639 ( .A1(n4549), .A2(REIP_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6740), .ZN(n4531) );
  OAI21_X1 U5640 ( .B1(n4532), .B2(n4541), .A(n4531), .ZN(U3194) );
  AOI22_X1 U5641 ( .A1(n4549), .A2(REIP_REG_14__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_12__SCAN_IN), .ZN(n4533) );
  OAI21_X1 U5642 ( .B1(n6269), .B2(n4541), .A(n4533), .ZN(U3196) );
  AOI22_X1 U5643 ( .A1(n4549), .A2(REIP_REG_16__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_14__SCAN_IN), .ZN(n4534) );
  OAI21_X1 U5644 ( .B1(n4535), .B2(n4541), .A(n4534), .ZN(U3198) );
  AOI22_X1 U5645 ( .A1(n4549), .A2(REIP_REG_17__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_15__SCAN_IN), .ZN(n4536) );
  OAI21_X1 U5646 ( .B1(n5984), .B2(n4541), .A(n4536), .ZN(U3199) );
  AOI22_X1 U5647 ( .A1(n4549), .A2(REIP_REG_20__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_18__SCAN_IN), .ZN(n4537) );
  OAI21_X1 U5648 ( .B1(n5957), .B2(n4541), .A(n4537), .ZN(U3202) );
  AOI22_X1 U5649 ( .A1(n4549), .A2(REIP_REG_21__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_19__SCAN_IN), .ZN(n4538) );
  OAI21_X1 U5650 ( .B1(n5948), .B2(n4541), .A(n4538), .ZN(U3203) );
  INV_X1 U5651 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5939) );
  AOI22_X1 U5652 ( .A1(n4549), .A2(REIP_REG_22__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_20__SCAN_IN), .ZN(n4539) );
  OAI21_X1 U5653 ( .B1(n5939), .B2(n4541), .A(n4539), .ZN(U3204) );
  AOI22_X1 U5654 ( .A1(n4549), .A2(REIP_REG_31__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_29__SCAN_IN), .ZN(n4540) );
  OAI21_X1 U5655 ( .B1(n5440), .B2(n4541), .A(n4540), .ZN(U3213) );
  INV_X1 U5656 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6958) );
  AOI22_X1 U5657 ( .A1(n4549), .A2(REIP_REG_24__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_22__SCAN_IN), .ZN(n4542) );
  OAI21_X1 U5658 ( .B1(n6958), .B2(n4541), .A(n4542), .ZN(U3206) );
  AOI22_X1 U5659 ( .A1(n4549), .A2(REIP_REG_25__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_23__SCAN_IN), .ZN(n4543) );
  OAI21_X1 U5660 ( .B1(n4544), .B2(n4541), .A(n4543), .ZN(U3207) );
  AOI22_X1 U5661 ( .A1(n4549), .A2(REIP_REG_27__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_25__SCAN_IN), .ZN(n4545) );
  OAI21_X1 U5662 ( .B1(n4546), .B2(n4541), .A(n4545), .ZN(U3209) );
  AOI22_X1 U5663 ( .A1(n4549), .A2(REIP_REG_28__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_26__SCAN_IN), .ZN(n4547) );
  OAI21_X1 U5664 ( .B1(n4548), .B2(n4541), .A(n4547), .ZN(U3210) );
  AOI22_X1 U5665 ( .A1(n4549), .A2(REIP_REG_30__SCAN_IN), .B1(n6740), .B2(
        ADDRESS_REG_28__SCAN_IN), .ZN(n4550) );
  OAI21_X1 U5666 ( .B1(n4551), .B2(n4541), .A(n4550), .ZN(U3212) );
  OR2_X1 U5667 ( .A1(n4770), .A2(n5778), .ZN(n4556) );
  NAND2_X1 U5668 ( .A1(n4774), .A2(n4552), .ZN(n4553) );
  NAND2_X1 U5669 ( .A1(n4554), .A2(n4553), .ZN(n4555) );
  NAND2_X1 U5670 ( .A1(n4556), .A2(n4555), .ZN(n4778) );
  INV_X1 U5671 ( .A(n5533), .ZN(n6711) );
  NOR2_X1 U5672 ( .A1(n4778), .A2(n6711), .ZN(n4557) );
  INV_X1 U5673 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6871) );
  NOR2_X1 U5674 ( .A1(n6722), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5654) );
  INV_X1 U5675 ( .A(n5654), .ZN(n4559) );
  OAI22_X1 U5676 ( .A1(n4557), .A2(n6871), .B1(n4813), .B2(n4559), .ZN(U2790)
         );
  INV_X1 U5677 ( .A(n4558), .ZN(n4560) );
  INV_X1 U5678 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6741) );
  OAI211_X1 U5679 ( .C1(n4560), .C2(n6741), .A(n4661), .B(n4559), .ZN(U2788)
         );
  INV_X1 U5680 ( .A(n4771), .ZN(n4564) );
  NAND2_X1 U5681 ( .A1(n4427), .A2(n5522), .ZN(n4561) );
  NAND2_X1 U5682 ( .A1(n4561), .A2(n6706), .ZN(n4562) );
  AOI21_X1 U5683 ( .B1(n4746), .B2(n4607), .A(n4562), .ZN(n4563) );
  MUX2_X1 U5684 ( .A(n4564), .B(n4563), .S(n4770), .Z(n4573) );
  NAND2_X1 U5685 ( .A1(n4770), .A2(n4715), .ZN(n4568) );
  INV_X1 U5686 ( .A(n4565), .ZN(n4566) );
  INV_X1 U5687 ( .A(n4569), .ZN(n4571) );
  NAND2_X1 U5688 ( .A1(n4571), .A2(n4570), .ZN(n4572) );
  AOI22_X1 U5689 ( .A1(n4763), .A2(n5533), .B1(n5024), .B2(FLUSH_REG_SCAN_IN), 
        .ZN(n4577) );
  NAND2_X1 U5690 ( .A1(n4813), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U5691 ( .A1(n4577), .A2(n4792), .ZN(n6240) );
  INV_X1 U5692 ( .A(n6544), .ZN(n5029) );
  NOR2_X1 U5693 ( .A1(n4574), .A2(n5029), .ZN(n4575) );
  XNOR2_X1 U5694 ( .A(n4575), .B(n4764), .ZN(n6334) );
  INV_X1 U5695 ( .A(n3760), .ZN(n4761) );
  NAND3_X1 U5696 ( .A1(n6334), .A2(n4761), .A3(n6707), .ZN(n4576) );
  OAI22_X1 U5697 ( .A1(n6240), .A2(n4764), .B1(n4577), .B2(n4576), .ZN(U3455)
         );
  NAND2_X1 U5698 ( .A1(n4579), .A2(n4578), .ZN(n4580) );
  NAND2_X1 U5699 ( .A1(n4581), .A2(n4580), .ZN(n6064) );
  INV_X1 U5700 ( .A(n4582), .ZN(n4585) );
  AND3_X1 U5701 ( .A1(n4836), .A2(n5513), .A3(n5533), .ZN(n4583) );
  NAND3_X1 U5702 ( .A1(n4585), .A2(n4584), .A3(n4583), .ZN(n4794) );
  INV_X2 U5703 ( .A(n6376), .ZN(n5832) );
  INV_X1 U5704 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4590) );
  OAI21_X1 U5705 ( .B1(n4589), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4588), 
        .ZN(n6468) );
  NAND2_X1 U5706 ( .A1(n6379), .A2(n5513), .ZN(n5829) );
  OAI222_X1 U5707 ( .A1(n6064), .A2(n5832), .B1(n6379), .B2(n4590), .C1(n6468), 
        .C2(n5829), .ZN(U2859) );
  INV_X1 U5708 ( .A(n6402), .ZN(n6383) );
  AOI222_X1 U5709 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6744), .B1(n6743), .B2(
        DATAO_REG_8__SCAN_IN), .C1(EAX_REG_8__SCAN_IN), .C2(n6383), .ZN(n4592)
         );
  INV_X1 U5710 ( .A(n4592), .ZN(U2915) );
  INV_X1 U5711 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4594) );
  AOI22_X1 U5712 ( .A1(n6383), .A2(EAX_REG_11__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n4593) );
  OAI21_X1 U5713 ( .B1(n6385), .B2(n4594), .A(n4593), .ZN(U2912) );
  INV_X1 U5714 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4596) );
  AOI22_X1 U5715 ( .A1(n6383), .A2(EAX_REG_3__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n4595) );
  OAI21_X1 U5716 ( .B1(n6385), .B2(n4596), .A(n4595), .ZN(U2920) );
  NOR2_X1 U5717 ( .A1(n4597), .A2(n4598), .ZN(n4599) );
  OAI21_X1 U5718 ( .B1(n6360), .B2(n4601), .A(n4600), .ZN(n4709) );
  AOI22_X1 U5719 ( .A1(n6375), .A2(n4709), .B1(n5830), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4602) );
  OAI21_X1 U5720 ( .B1(n6368), .B2(n5832), .A(n4602), .ZN(U2858) );
  OAI21_X1 U5721 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6236), .A(n6240), 
        .ZN(n4629) );
  INV_X1 U5722 ( .A(n4629), .ZN(n4622) );
  INV_X1 U5723 ( .A(n6240), .ZN(n5511) );
  AND3_X1 U5724 ( .A1(n3760), .A2(n4607), .A3(n4606), .ZN(n4608) );
  NAND2_X1 U5725 ( .A1(n4609), .A2(n4608), .ZN(n4736) );
  INV_X1 U5726 ( .A(n4736), .ZN(n4610) );
  OR2_X1 U5727 ( .A1(n4605), .A2(n4610), .ZN(n4617) );
  INV_X1 U5728 ( .A(n4612), .ZN(n4624) );
  OAI21_X1 U5729 ( .B1(n4613), .B2(n4611), .A(n4624), .ZN(n4614) );
  OAI21_X1 U5730 ( .B1(n4746), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4614), 
        .ZN(n4615) );
  INV_X1 U5731 ( .A(n4615), .ZN(n4616) );
  NAND2_X1 U5732 ( .A1(n4617), .A2(n4616), .ZN(n4723) );
  INV_X1 U5733 ( .A(n4611), .ZN(n4619) );
  OAI22_X1 U5734 ( .A1(n6454), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4618), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U5735 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5506) );
  OAI22_X1 U5736 ( .A1(n6236), .A2(n4619), .B1(n5504), .B2(n5506), .ZN(n4620)
         );
  AOI21_X1 U5737 ( .B1(n6707), .B2(n4723), .A(n4620), .ZN(n4621) );
  OAI22_X1 U5738 ( .A1(n4622), .A2(n4603), .B1(n5511), .B2(n4621), .ZN(U3460)
         );
  NOR2_X1 U5739 ( .A1(n4746), .A2(n3895), .ZN(n4724) );
  INV_X1 U5740 ( .A(n4724), .ZN(n4631) );
  INV_X1 U5741 ( .A(n6707), .ZN(n6238) );
  NAND2_X1 U5742 ( .A1(n4623), .A2(n4736), .ZN(n4626) );
  NAND2_X1 U5743 ( .A1(n4624), .A2(n3895), .ZN(n4625) );
  NAND2_X1 U5744 ( .A1(n4626), .A2(n4625), .ZN(n4725) );
  INV_X1 U5745 ( .A(n4725), .ZN(n4627) );
  OAI22_X1 U5746 ( .A1(n4627), .A2(n6238), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6704), .ZN(n4628) );
  OAI22_X1 U5747 ( .A1(n4629), .A2(n4628), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6240), .ZN(n4630) );
  OAI21_X1 U5748 ( .B1(n4631), .B2(n6238), .A(n4630), .ZN(U3461) );
  INV_X1 U5749 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4634) );
  INV_X1 U5750 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4633) );
  INV_X1 U5751 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n4632) );
  OAI222_X1 U5752 ( .A1(n4634), .A2(n6385), .B1(n6747), .B2(n4633), .C1(n4786), 
        .C2(n4632), .ZN(U2898) );
  INV_X1 U5753 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4637) );
  INV_X1 U5754 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4636) );
  INV_X1 U5755 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n4635) );
  OAI222_X1 U5756 ( .A1(n4637), .A2(n6385), .B1(n6747), .B2(n4636), .C1(n4786), 
        .C2(n4635), .ZN(U2899) );
  INV_X1 U5757 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4639) );
  INV_X1 U5758 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n4638) );
  OAI222_X1 U5759 ( .A1(n4639), .A2(n6385), .B1(n6747), .B2(n4259), .C1(n4786), 
        .C2(n4638), .ZN(U2897) );
  INV_X1 U5760 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4642) );
  INV_X1 U5761 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4641) );
  INV_X1 U5762 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n4640) );
  OAI222_X1 U5763 ( .A1(n4642), .A2(n6385), .B1(n6747), .B2(n4641), .C1(n4786), 
        .C2(n4640), .ZN(U2896) );
  INV_X1 U5764 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4645) );
  INV_X1 U5765 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4644) );
  INV_X1 U5766 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4643) );
  OAI222_X1 U5767 ( .A1(n4645), .A2(n6385), .B1(n6747), .B2(n4644), .C1(n4786), 
        .C2(n4643), .ZN(U2903) );
  INV_X1 U5768 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4647) );
  INV_X1 U5769 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n4646) );
  OAI222_X1 U5770 ( .A1(n4647), .A2(n6385), .B1(n6747), .B2(n4341), .C1(n4786), 
        .C2(n4646), .ZN(U2895) );
  INV_X1 U5771 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4649) );
  INV_X1 U5772 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6955) );
  INV_X1 U5773 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4648) );
  OAI222_X1 U5774 ( .A1(n4649), .A2(n6385), .B1(n4786), .B2(n6955), .C1(n4648), 
        .C2(n6747), .ZN(U2894) );
  INV_X1 U5775 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4652) );
  INV_X1 U5776 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4651) );
  INV_X1 U5777 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n4650) );
  OAI222_X1 U5778 ( .A1(n4652), .A2(n6385), .B1(n6747), .B2(n4651), .C1(n4786), 
        .C2(n4650), .ZN(U2907) );
  INV_X1 U5779 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4654) );
  INV_X1 U5780 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n7037) );
  OAI222_X1 U5781 ( .A1(n4654), .A2(n6385), .B1(n4786), .B2(n7037), .C1(n4653), 
        .C2(n6747), .ZN(U2901) );
  INV_X1 U5782 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4656) );
  INV_X1 U5783 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n6835) );
  OAI222_X1 U5784 ( .A1(n4656), .A2(n6385), .B1(n4786), .B2(n6835), .C1(n4655), 
        .C2(n6747), .ZN(U2905) );
  INV_X1 U5785 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4657) );
  INV_X1 U5786 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6850) );
  OAI222_X1 U5787 ( .A1(n4657), .A2(n6385), .B1(n4786), .B2(n6850), .C1(n5325), 
        .C2(n6402), .ZN(U2917) );
  INV_X1 U5788 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4660) );
  INV_X1 U5789 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4658) );
  OAI222_X1 U5790 ( .A1(n4786), .A2(n4660), .B1(n6747), .B2(n4659), .C1(n6385), 
        .C2(n4658), .ZN(U2906) );
  INV_X1 U5791 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n6834) );
  INV_X1 U5792 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n6945) );
  OAI222_X1 U5793 ( .A1(n6402), .A2(n6997), .B1(n6385), .B2(n6834), .C1(n4786), 
        .C2(n6945), .ZN(U2908) );
  AOI22_X1 U5794 ( .A1(n6418), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6415), .ZN(n4664) );
  NAND2_X1 U5795 ( .A1(n6419), .A2(DATAI_3_), .ZN(n4695) );
  NAND2_X1 U5796 ( .A1(n4664), .A2(n4695), .ZN(U2942) );
  AOI22_X1 U5797 ( .A1(n6418), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6415), .ZN(n4665) );
  NAND2_X1 U5798 ( .A1(n6419), .A2(DATAI_6_), .ZN(n4672) );
  NAND2_X1 U5799 ( .A1(n4665), .A2(n4672), .ZN(U2945) );
  AOI22_X1 U5800 ( .A1(n6418), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6415), .ZN(n4666) );
  NAND2_X1 U5801 ( .A1(n6419), .A2(DATAI_13_), .ZN(n4677) );
  NAND2_X1 U5802 ( .A1(n4666), .A2(n4677), .ZN(U2937) );
  AOI22_X1 U5803 ( .A1(n6418), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6415), .ZN(n4667) );
  INV_X1 U5804 ( .A(DATAI_0_), .ZN(n4802) );
  OR2_X1 U5805 ( .A1(n4798), .A2(n4802), .ZN(n4668) );
  NAND2_X1 U5806 ( .A1(n4667), .A2(n4668), .ZN(U2924) );
  AOI22_X1 U5807 ( .A1(n6418), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6415), .ZN(n4669) );
  NAND2_X1 U5808 ( .A1(n4669), .A2(n4668), .ZN(U2939) );
  AOI22_X1 U5809 ( .A1(n6418), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6415), .ZN(n4670) );
  INV_X1 U5810 ( .A(DATAI_1_), .ZN(n4801) );
  OR2_X1 U5811 ( .A1(n4798), .A2(n4801), .ZN(n4679) );
  NAND2_X1 U5812 ( .A1(n4670), .A2(n4679), .ZN(U2940) );
  AOI22_X1 U5813 ( .A1(n6418), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6415), .ZN(n4671) );
  INV_X1 U5814 ( .A(DATAI_5_), .ZN(n4965) );
  OR2_X1 U5815 ( .A1(n4798), .A2(n4965), .ZN(n4686) );
  NAND2_X1 U5816 ( .A1(n4671), .A2(n4686), .ZN(U2944) );
  AOI22_X1 U5817 ( .A1(n6418), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6415), .ZN(n4673) );
  NAND2_X1 U5818 ( .A1(n4673), .A2(n4672), .ZN(U2930) );
  AOI22_X1 U5819 ( .A1(n6418), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6415), .ZN(n4674) );
  NAND2_X1 U5820 ( .A1(n6419), .A2(DATAI_7_), .ZN(n4690) );
  NAND2_X1 U5821 ( .A1(n4674), .A2(n4690), .ZN(U2946) );
  AOI22_X1 U5822 ( .A1(n6418), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n6415), .ZN(n4675) );
  NAND2_X1 U5823 ( .A1(n6419), .A2(DATAI_12_), .ZN(n4681) );
  NAND2_X1 U5824 ( .A1(n4675), .A2(n4681), .ZN(U2936) );
  AOI22_X1 U5825 ( .A1(n6418), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6415), .ZN(n4676) );
  NAND2_X1 U5826 ( .A1(n6419), .A2(DATAI_4_), .ZN(n4688) );
  NAND2_X1 U5827 ( .A1(n4676), .A2(n4688), .ZN(U2943) );
  AOI22_X1 U5828 ( .A1(n6418), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6415), .ZN(n4678) );
  NAND2_X1 U5829 ( .A1(n4678), .A2(n4677), .ZN(U2952) );
  AOI22_X1 U5830 ( .A1(n6418), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6415), .ZN(n4680) );
  NAND2_X1 U5831 ( .A1(n4680), .A2(n4679), .ZN(U2925) );
  AOI22_X1 U5832 ( .A1(n6418), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n6415), .ZN(n4682) );
  NAND2_X1 U5833 ( .A1(n4682), .A2(n4681), .ZN(U2951) );
  AOI22_X1 U5834 ( .A1(n6418), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6415), .ZN(n4683) );
  INV_X1 U5835 ( .A(DATAI_2_), .ZN(n4910) );
  OR2_X1 U5836 ( .A1(n4798), .A2(n4910), .ZN(n4684) );
  NAND2_X1 U5837 ( .A1(n4683), .A2(n4684), .ZN(U2941) );
  AOI22_X1 U5838 ( .A1(n6418), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6415), .ZN(n4685) );
  NAND2_X1 U5839 ( .A1(n4685), .A2(n4684), .ZN(U2926) );
  AOI22_X1 U5840 ( .A1(n6418), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6415), .ZN(n4687) );
  NAND2_X1 U5841 ( .A1(n4687), .A2(n4686), .ZN(U2929) );
  AOI22_X1 U5842 ( .A1(n6418), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6415), .ZN(n4689) );
  NAND2_X1 U5843 ( .A1(n4689), .A2(n4688), .ZN(U2928) );
  AOI22_X1 U5844 ( .A1(n6418), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6415), .ZN(n4691) );
  NAND2_X1 U5845 ( .A1(n4691), .A2(n4690), .ZN(U2931) );
  AOI22_X1 U5846 ( .A1(n6418), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6415), .ZN(n4692) );
  INV_X1 U5847 ( .A(DATAI_9_), .ZN(n5890) );
  OR2_X1 U5848 ( .A1(n4798), .A2(n5890), .ZN(n4693) );
  NAND2_X1 U5849 ( .A1(n4692), .A2(n4693), .ZN(U2948) );
  AOI22_X1 U5850 ( .A1(n6418), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n6415), .ZN(n4694) );
  NAND2_X1 U5851 ( .A1(n4694), .A2(n4693), .ZN(U2933) );
  AOI22_X1 U5852 ( .A1(n6418), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6415), .ZN(n4696) );
  NAND2_X1 U5853 ( .A1(n4696), .A2(n4695), .ZN(U2927) );
  INV_X1 U5854 ( .A(n6747), .ZN(n6381) );
  AOI222_X1 U5855 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6381), .B1(n6743), .B2(
        DATAO_REG_30__SCAN_IN), .C1(n6744), .C2(UWORD_REG_14__SCAN_IN), .ZN(
        n4697) );
  INV_X1 U5856 ( .A(n4697), .ZN(U2893) );
  AOI222_X1 U5857 ( .A1(EAX_REG_23__SCAN_IN), .A2(n6381), .B1(n6743), .B2(
        DATAO_REG_23__SCAN_IN), .C1(n6744), .C2(UWORD_REG_7__SCAN_IN), .ZN(
        n4698) );
  INV_X1 U5858 ( .A(n4698), .ZN(U2900) );
  INV_X1 U5859 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6928) );
  NAND2_X1 U5860 ( .A1(n6457), .A2(REIP_REG_1__SCAN_IN), .ZN(n4706) );
  OAI21_X1 U5861 ( .B1(n6056), .B2(n6928), .A(n4706), .ZN(n4703) );
  OAI21_X1 U5862 ( .B1(n4701), .B2(n4700), .A(n4699), .ZN(n4712) );
  NOR2_X1 U5863 ( .A1(n4712), .A2(n6245), .ZN(n4702) );
  AOI211_X1 U5864 ( .C1(n6060), .C2(n6928), .A(n4703), .B(n4702), .ZN(n4704)
         );
  OAI21_X1 U5865 ( .B1(n6057), .B2(n6368), .A(n4704), .ZN(U2985) );
  NOR2_X1 U5866 ( .A1(n6460), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4705)
         );
  OAI21_X1 U5867 ( .B1(n5154), .B2(n4705), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4711) );
  INV_X1 U5868 ( .A(n4706), .ZN(n4708) );
  NAND2_X1 U5869 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n6160), .ZN(n6450)
         );
  AOI21_X1 U5870 ( .B1(n6455), .B2(n6450), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4707) );
  AOI211_X1 U5871 ( .C1(n6470), .C2(n4709), .A(n4708), .B(n4707), .ZN(n4710)
         );
  OAI211_X1 U5872 ( .C1(n4712), .C2(n6473), .A(n4711), .B(n4710), .ZN(U3017)
         );
  NAND2_X1 U5873 ( .A1(n4714), .A2(n4736), .ZN(n4722) );
  INV_X1 U5874 ( .A(n4715), .ZN(n4716) );
  NAND2_X1 U5875 ( .A1(n4771), .A2(n4716), .ZN(n4749) );
  XNOR2_X1 U5876 ( .A(n4717), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4720)
         );
  XNOR2_X1 U5877 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4718) );
  OAI22_X1 U5878 ( .A1(n4746), .A2(n4718), .B1(n4744), .B2(n4720), .ZN(n4719)
         );
  AOI21_X1 U5879 ( .B1(n4749), .B2(n4720), .A(n4719), .ZN(n4721) );
  AND2_X1 U5880 ( .A1(n4722), .A2(n4721), .ZN(n5503) );
  MUX2_X1 U5881 ( .A(n3903), .B(n5503), .S(n4763), .Z(n4731) );
  NAND2_X1 U5882 ( .A1(n4731), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4733) );
  NAND2_X1 U5883 ( .A1(n4763), .A2(n4723), .ZN(n4730) );
  OR3_X1 U5884 ( .A1(n4725), .A2(n4724), .A3(n6541), .ZN(n4727) );
  NAND2_X1 U5885 ( .A1(n4727), .A2(n4726), .ZN(n4729) );
  NOR2_X1 U5886 ( .A1(n4727), .A2(n4726), .ZN(n4728) );
  AOI21_X1 U5887 ( .B1(n4730), .B2(n4729), .A(n4728), .ZN(n4732) );
  INV_X1 U5888 ( .A(n4731), .ZN(n4757) );
  AOI22_X1 U5889 ( .A1(n4733), .A2(n4732), .B1(n4757), .B2(n4984), .ZN(n4754)
         );
  NAND2_X1 U5890 ( .A1(n4735), .A2(n4736), .ZN(n4751) );
  MUX2_X1 U5891 ( .A(n3274), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4717), 
        .Z(n4737) );
  NOR2_X1 U5892 ( .A1(n4737), .A2(n4758), .ZN(n4748) );
  NAND2_X1 U5893 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4739) );
  INV_X1 U5894 ( .A(n4739), .ZN(n4738) );
  MUX2_X1 U5895 ( .A(n4739), .B(n4738), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4745) );
  INV_X1 U5896 ( .A(n4740), .ZN(n4741) );
  OAI21_X1 U5897 ( .B1(n4717), .B2(n4742), .A(n4741), .ZN(n4743) );
  NOR2_X1 U5898 ( .A1(n4743), .A2(n3079), .ZN(n6237) );
  OAI22_X1 U5899 ( .A1(n4746), .A2(n4745), .B1(n6237), .B2(n4744), .ZN(n4747)
         );
  AOI21_X1 U5900 ( .B1(n4749), .B2(n4748), .A(n4747), .ZN(n4750) );
  NAND2_X1 U5901 ( .A1(n4751), .A2(n4750), .ZN(n6235) );
  MUX2_X1 U5902 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6235), .S(n4763), 
        .Z(n4756) );
  NOR2_X1 U5903 ( .A1(n4756), .A2(n6731), .ZN(n4753) );
  INV_X1 U5904 ( .A(n4756), .ZN(n4752) );
  OAI22_X1 U5905 ( .A1(n4754), .A2(n4753), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4752), .ZN(n4755) );
  NAND2_X1 U5906 ( .A1(n4755), .A2(n6482), .ZN(n4785) );
  NAND3_X1 U5907 ( .A1(n4757), .A2(n4756), .A3(n6704), .ZN(n4760) );
  NOR2_X1 U5908 ( .A1(FLUSH_REG_SCAN_IN), .A2(n6704), .ZN(n4766) );
  NAND2_X1 U5909 ( .A1(n4766), .A2(n4758), .ZN(n4759) );
  NAND2_X1 U5910 ( .A1(n4760), .A2(n4759), .ZN(n4859) );
  NAND2_X1 U5911 ( .A1(n6334), .A2(n4761), .ZN(n4762) );
  OAI21_X1 U5912 ( .B1(n4764), .B2(n4763), .A(n4762), .ZN(n4765) );
  NAND2_X1 U5913 ( .A1(n4765), .A2(n6704), .ZN(n4768) );
  NAND2_X1 U5914 ( .A1(n4766), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4767) );
  NAND2_X1 U5915 ( .A1(n4768), .A2(n4767), .ZN(n4857) );
  NOR2_X1 U5916 ( .A1(n4769), .A2(n4421), .ZN(n4772) );
  MUX2_X1 U5917 ( .A(n4772), .B(n4771), .S(n4770), .Z(n4776) );
  NAND2_X1 U5918 ( .A1(n4774), .A2(n4773), .ZN(n4775) );
  NAND2_X1 U5919 ( .A1(n4776), .A2(n4775), .ZN(n5535) );
  OR2_X1 U5920 ( .A1(n5774), .A2(n5521), .ZN(n5518) );
  AOI21_X1 U5921 ( .B1(n5518), .B2(n5522), .A(READY_N), .ZN(n4777) );
  OR2_X1 U5922 ( .A1(n4778), .A2(n4777), .ZN(n5534) );
  INV_X1 U5923 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6943) );
  INV_X1 U5924 ( .A(MORE_REG_SCAN_IN), .ZN(n4779) );
  AND2_X1 U5925 ( .A1(n6943), .A2(n4779), .ZN(n4781) );
  OAI21_X1 U5926 ( .B1(n5534), .B2(n4781), .A(n4780), .ZN(n4782) );
  OR3_X1 U5927 ( .A1(n4857), .A2(n5535), .A3(n4782), .ZN(n4783) );
  NOR2_X1 U5928 ( .A1(n4859), .A2(n4783), .ZN(n4784) );
  NAND2_X1 U5929 ( .A1(n4785), .A2(n4784), .ZN(n5020) );
  OAI22_X1 U5930 ( .A1(n5020), .A2(n6711), .B1(n6706), .B2(n4786), .ZN(n4790)
         );
  OR2_X1 U5931 ( .A1(n4788), .A2(n4787), .ZN(n4789) );
  NAND2_X1 U5932 ( .A1(n4790), .A2(n4789), .ZN(n6708) );
  OAI211_X1 U5933 ( .C1(n6708), .C2(n5217), .A(n4792), .B(n4791), .ZN(U3453)
         );
  NOR2_X1 U5934 ( .A1(n4794), .A2(n4793), .ZN(n4795) );
  INV_X1 U5935 ( .A(n4799), .ZN(n4800) );
  INV_X1 U5936 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6823) );
  OAI222_X1 U5937 ( .A1(n6368), .A2(n5892), .B1(n5891), .B2(n4801), .C1(n5889), 
        .C2(n6823), .ZN(U2890) );
  INV_X1 U5938 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6403) );
  OAI222_X1 U5939 ( .A1(n6064), .A2(n5892), .B1(n5891), .B2(n4802), .C1(n5889), 
        .C2(n6403), .ZN(U2891) );
  NAND2_X1 U5940 ( .A1(n5101), .A2(n6227), .ZN(n4806) );
  INV_X1 U5941 ( .A(n6687), .ZN(n5411) );
  OR2_X1 U5942 ( .A1(n4817), .A2(n4807), .ZN(n5253) );
  NAND2_X1 U5943 ( .A1(n4735), .A2(n4623), .ZN(n5067) );
  INV_X1 U5944 ( .A(n4605), .ZN(n6363) );
  NAND2_X1 U5945 ( .A1(n4714), .A2(n6363), .ZN(n6545) );
  OR2_X1 U5946 ( .A1(n5067), .A2(n6545), .ZN(n4809) );
  INV_X1 U5947 ( .A(n4808), .ZN(n4850) );
  NAND2_X1 U5948 ( .A1(n4809), .A2(n4850), .ZN(n4819) );
  AOI22_X1 U5949 ( .A1(n4819), .A2(n6651), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4810), .ZN(n4851) );
  INV_X1 U5950 ( .A(n4860), .ZN(n4811) );
  NAND2_X1 U5951 ( .A1(n4811), .A2(n5525), .ZN(n4812) );
  INV_X1 U5952 ( .A(DATAI_6_), .ZN(n5324) );
  OAI22_X1 U5953 ( .A1(n4851), .A2(n6691), .B1(n4850), .B2(n6621), .ZN(n4816)
         );
  AOI21_X1 U5954 ( .B1(n6688), .B2(n4853), .A(n4816), .ZN(n4822) );
  AOI21_X1 U5955 ( .B1(n4817), .B2(n6065), .A(n6728), .ZN(n4820) );
  INV_X1 U5956 ( .A(n6648), .ZN(n5306) );
  AOI21_X1 U5957 ( .B1(n5176), .B2(n6722), .A(n5306), .ZN(n4818) );
  NAND2_X1 U5958 ( .A1(n4854), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4821)
         );
  OAI211_X1 U5959 ( .C1(n5212), .C2(n5411), .A(n4822), .B(n4821), .ZN(U3146)
         );
  NAND2_X1 U5960 ( .A1(n6065), .A2(DATAI_26_), .ZN(n6602) );
  OAI22_X1 U5961 ( .A1(n4851), .A2(n6667), .B1(n4850), .B2(n6601), .ZN(n4824)
         );
  AOI21_X1 U5962 ( .B1(n6664), .B2(n4853), .A(n4824), .ZN(n4826) );
  NAND2_X1 U5963 ( .A1(n4854), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4825)
         );
  OAI211_X1 U5964 ( .C1(n5212), .C2(n6602), .A(n4826), .B(n4825), .ZN(U3142)
         );
  INV_X1 U5965 ( .A(n6652), .ZN(n5436) );
  NAND2_X1 U5966 ( .A1(n6065), .A2(DATAI_16_), .ZN(n6587) );
  INV_X1 U5967 ( .A(n6587), .ZN(n6644) );
  OR2_X1 U5968 ( .A1(n4849), .A2(n4827), .ZN(n6586) );
  OAI22_X1 U5969 ( .A1(n4851), .A2(n6655), .B1(n4850), .B2(n6586), .ZN(n4828)
         );
  AOI21_X1 U5970 ( .B1(n6644), .B2(n4853), .A(n4828), .ZN(n4830) );
  NAND2_X1 U5971 ( .A1(n4854), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4829)
         );
  OAI211_X1 U5972 ( .C1(n5212), .C2(n5436), .A(n4830), .B(n4829), .ZN(U3140)
         );
  INV_X1 U5973 ( .A(DATAI_7_), .ZN(n4831) );
  OAI22_X1 U5974 ( .A1(n4851), .A2(n6701), .B1(n4850), .B2(n6628), .ZN(n4832)
         );
  AOI21_X1 U5975 ( .B1(n6694), .B2(n4853), .A(n4832), .ZN(n4834) );
  NAND2_X1 U5976 ( .A1(n4854), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4833)
         );
  OAI211_X1 U5977 ( .C1(n5212), .C2(n6630), .A(n4834), .B(n4833), .ZN(U3147)
         );
  NAND2_X1 U5978 ( .A1(n6065), .A2(DATAI_28_), .ZN(n6612) );
  INV_X1 U5979 ( .A(DATAI_4_), .ZN(n4835) );
  OR2_X1 U5980 ( .A1(n4849), .A2(n4836), .ZN(n6611) );
  OAI22_X1 U5981 ( .A1(n4851), .A2(n6679), .B1(n4850), .B2(n6611), .ZN(n4837)
         );
  AOI21_X1 U5982 ( .B1(n6676), .B2(n4853), .A(n4837), .ZN(n4839) );
  NAND2_X1 U5983 ( .A1(n4854), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4838)
         );
  OAI211_X1 U5984 ( .C1(n5212), .C2(n6612), .A(n4839), .B(n4838), .ZN(U3144)
         );
  INV_X1 U5985 ( .A(n6681), .ZN(n5415) );
  OAI22_X1 U5986 ( .A1(n4851), .A2(n6685), .B1(n4850), .B2(n6616), .ZN(n4840)
         );
  AOI21_X1 U5987 ( .B1(n6682), .B2(n4853), .A(n4840), .ZN(n4842) );
  NAND2_X1 U5988 ( .A1(n4854), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4841)
         );
  OAI211_X1 U5989 ( .C1(n5212), .C2(n5415), .A(n4842), .B(n4841), .ZN(U3145)
         );
  INV_X1 U5990 ( .A(n6658), .ZN(n6597) );
  OAI22_X1 U5991 ( .A1(n4851), .A2(n6661), .B1(n4850), .B2(n6596), .ZN(n4844)
         );
  AOI21_X1 U5992 ( .B1(n6657), .B2(n4853), .A(n4844), .ZN(n4846) );
  NAND2_X1 U5993 ( .A1(n4854), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4845)
         );
  OAI211_X1 U5994 ( .C1(n5212), .C2(n6597), .A(n4846), .B(n4845), .ZN(U3141)
         );
  INV_X1 U5995 ( .A(n6669), .ZN(n5422) );
  INV_X1 U5996 ( .A(DATAI_3_), .ZN(n4847) );
  INV_X1 U5997 ( .A(n3391), .ZN(n4848) );
  OAI22_X1 U5998 ( .A1(n4851), .A2(n6673), .B1(n4850), .B2(n6606), .ZN(n4852)
         );
  AOI21_X1 U5999 ( .B1(n6670), .B2(n4853), .A(n4852), .ZN(n4856) );
  NAND2_X1 U6000 ( .A1(n4854), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4855)
         );
  OAI211_X1 U6001 ( .C1(n5212), .C2(n5422), .A(n4856), .B(n4855), .ZN(U3143)
         );
  AOI21_X1 U6002 ( .B1(n4859), .B2(n4858), .A(n4857), .ZN(n5025) );
  NAND2_X1 U6003 ( .A1(n5217), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6226) );
  AOI222_X1 U6004 ( .A1(n5025), .A2(n4860), .B1(n4623), .B2(n6226), .C1(n6499), 
        .C2(n6651), .ZN(n4864) );
  NAND2_X1 U6005 ( .A1(n5025), .A2(n6943), .ZN(n4861) );
  NAND2_X1 U6006 ( .A1(n4861), .A2(n5024), .ZN(n4862) );
  NAND2_X1 U6007 ( .A1(n6732), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4863) );
  OAI21_X1 U6008 ( .B1(n4864), .B2(n6732), .A(n4863), .ZN(U3465) );
  OAI21_X1 U6009 ( .B1(n4865), .B2(n4867), .A(n4866), .ZN(n6352) );
  INV_X1 U6010 ( .A(n4911), .ZN(n4871) );
  INV_X1 U6011 ( .A(n4869), .ZN(n4870) );
  OAI21_X1 U6012 ( .B1(n4868), .B2(n4871), .A(n4870), .ZN(n4872) );
  AND2_X1 U6013 ( .A1(n4872), .A2(n4927), .ZN(n6346) );
  AOI22_X1 U6014 ( .A1(n6375), .A2(n6346), .B1(EBX_REG_3__SCAN_IN), .B2(n5830), 
        .ZN(n4873) );
  OAI21_X1 U6015 ( .B1(n6352), .B2(n5832), .A(n4873), .ZN(U2856) );
  INV_X1 U6016 ( .A(n6227), .ZN(n5213) );
  NAND2_X1 U6017 ( .A1(n5213), .A2(n5101), .ZN(n4874) );
  NAND2_X1 U6018 ( .A1(n4714), .A2(n4605), .ZN(n5102) );
  NOR2_X1 U6019 ( .A1(n5104), .A2(n6731), .ZN(n5031) );
  NAND2_X1 U6020 ( .A1(n5031), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4901) );
  OAI21_X1 U6021 ( .B1(n5067), .B2(n5102), .A(n4901), .ZN(n4879) );
  NAND2_X1 U6022 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4875) );
  NOR2_X1 U6023 ( .A1(n5104), .A2(n4875), .ZN(n4876) );
  AOI21_X1 U6024 ( .B1(n4879), .B2(n6651), .A(n4876), .ZN(n4902) );
  OAI22_X1 U6025 ( .A1(n4902), .A2(n6661), .B1(n6596), .B2(n4901), .ZN(n4877)
         );
  AOI21_X1 U6026 ( .B1(n6658), .B2(n5060), .A(n4877), .ZN(n4882) );
  NOR2_X1 U6027 ( .A1(n4878), .A2(n6244), .ZN(n4980) );
  NAND2_X1 U6028 ( .A1(n4904), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4881)
         );
  OAI211_X1 U6029 ( .C1(n5173), .C2(n6557), .A(n4882), .B(n4881), .ZN(U3125)
         );
  OAI22_X1 U6030 ( .A1(n4902), .A2(n6673), .B1(n6606), .B2(n4901), .ZN(n4883)
         );
  AOI21_X1 U6031 ( .B1(n6669), .B2(n5060), .A(n4883), .ZN(n4885) );
  NAND2_X1 U6032 ( .A1(n4904), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4884)
         );
  OAI211_X1 U6033 ( .C1(n5173), .C2(n6607), .A(n4885), .B(n4884), .ZN(U3127)
         );
  INV_X1 U6034 ( .A(n6694), .ZN(n6582) );
  OAI22_X1 U6035 ( .A1(n4902), .A2(n6701), .B1(n6628), .B2(n4901), .ZN(n4886)
         );
  AOI21_X1 U6036 ( .B1(n6697), .B2(n5060), .A(n4886), .ZN(n4888) );
  NAND2_X1 U6037 ( .A1(n4904), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4887)
         );
  OAI211_X1 U6038 ( .C1(n5173), .C2(n6582), .A(n4888), .B(n4887), .ZN(U3131)
         );
  OAI22_X1 U6039 ( .A1(n4902), .A2(n6655), .B1(n6586), .B2(n4901), .ZN(n4889)
         );
  AOI21_X1 U6040 ( .B1(n6652), .B2(n5060), .A(n4889), .ZN(n4891) );
  NAND2_X1 U6041 ( .A1(n4904), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4890)
         );
  OAI211_X1 U6042 ( .C1(n5173), .C2(n6587), .A(n4891), .B(n4890), .ZN(U3124)
         );
  OAI22_X1 U6043 ( .A1(n4902), .A2(n6685), .B1(n6616), .B2(n4901), .ZN(n4892)
         );
  AOI21_X1 U6044 ( .B1(n6681), .B2(n5060), .A(n4892), .ZN(n4894) );
  NAND2_X1 U6045 ( .A1(n4904), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4893)
         );
  OAI211_X1 U6046 ( .C1(n5173), .C2(n6617), .A(n4894), .B(n4893), .ZN(U3129)
         );
  INV_X1 U6047 ( .A(n6676), .ZN(n6568) );
  OAI22_X1 U6048 ( .A1(n4902), .A2(n6679), .B1(n6611), .B2(n4901), .ZN(n4895)
         );
  AOI21_X1 U6049 ( .B1(n6675), .B2(n5060), .A(n4895), .ZN(n4897) );
  NAND2_X1 U6050 ( .A1(n4904), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4896)
         );
  OAI211_X1 U6051 ( .C1(n5173), .C2(n6568), .A(n4897), .B(n4896), .ZN(U3128)
         );
  INV_X1 U6052 ( .A(n6664), .ZN(n6561) );
  OAI22_X1 U6053 ( .A1(n4902), .A2(n6667), .B1(n6601), .B2(n4901), .ZN(n4898)
         );
  AOI21_X1 U6054 ( .B1(n6663), .B2(n5060), .A(n4898), .ZN(n4900) );
  NAND2_X1 U6055 ( .A1(n4904), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4899)
         );
  OAI211_X1 U6056 ( .C1(n5173), .C2(n6561), .A(n4900), .B(n4899), .ZN(U3126)
         );
  INV_X1 U6057 ( .A(n6688), .ZN(n6622) );
  OAI22_X1 U6058 ( .A1(n4902), .A2(n6691), .B1(n6621), .B2(n4901), .ZN(n4903)
         );
  AOI21_X1 U6059 ( .B1(n6687), .B2(n5060), .A(n4903), .ZN(n4906) );
  NAND2_X1 U6060 ( .A1(n4904), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4905)
         );
  OAI211_X1 U6061 ( .C1(n5173), .C2(n6622), .A(n4906), .B(n4905), .ZN(U3130)
         );
  NOR2_X1 U6062 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  NOR2_X1 U6063 ( .A1(n4865), .A2(n4909), .ZN(n6427) );
  INV_X1 U6064 ( .A(n6427), .ZN(n4913) );
  INV_X1 U6065 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6399) );
  OAI222_X1 U6066 ( .A1(n4913), .A2(n5892), .B1(n5891), .B2(n4910), .C1(n5889), 
        .C2(n6399), .ZN(U2889) );
  XNOR2_X1 U6067 ( .A(n4868), .B(n4911), .ZN(n6453) );
  INV_X1 U6068 ( .A(n6453), .ZN(n4912) );
  INV_X1 U6069 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5775) );
  OAI222_X1 U6070 ( .A1(n4913), .A2(n5832), .B1(n5829), .B2(n4912), .C1(n6379), 
        .C2(n5775), .ZN(U2857) );
  XNOR2_X1 U6071 ( .A(n4915), .B(n4914), .ZN(n4954) );
  AOI21_X1 U6072 ( .B1(n4916), .B2(n4917), .A(n5154), .ZN(n6466) );
  OAI21_X1 U6073 ( .B1(n6460), .B2(n6459), .A(n6466), .ZN(n4947) );
  OAI21_X1 U6074 ( .B1(n6455), .B2(n4917), .A(n6460), .ZN(n5159) );
  AND2_X1 U6075 ( .A1(n5159), .A2(n6459), .ZN(n4918) );
  AOI22_X1 U6076 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4947), .B1(n4918), 
        .B2(n3588), .ZN(n4920) );
  NOR2_X1 U6077 ( .A1(n6218), .A2(n7022), .ZN(n4949) );
  AOI21_X1 U6078 ( .B1(n6470), .B2(n6346), .A(n4949), .ZN(n4919) );
  OAI211_X1 U6079 ( .C1(n4954), .C2(n6473), .A(n4920), .B(n4919), .ZN(U3015)
         );
  INV_X1 U6080 ( .A(EAX_REG_3__SCAN_IN), .ZN(n4921) );
  OAI222_X1 U6081 ( .A1(n6352), .A2(n5892), .B1(n5891), .B2(n4847), .C1(n5889), 
        .C2(n4921), .ZN(U2888) );
  AND2_X1 U6082 ( .A1(n4866), .A2(n4922), .ZN(n4924) );
  OR2_X1 U6083 ( .A1(n4924), .A2(n4923), .ZN(n6340) );
  AND2_X1 U6084 ( .A1(n4927), .A2(n4926), .ZN(n4928) );
  NOR2_X1 U6085 ( .A1(n4925), .A2(n4928), .ZN(n6337) );
  AOI22_X1 U6086 ( .A1(n6375), .A2(n6337), .B1(n5830), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4929) );
  OAI21_X1 U6087 ( .B1(n6340), .B2(n5832), .A(n4929), .ZN(U2855) );
  CLKBUF_X1 U6088 ( .A(n4931), .Z(n4932) );
  XNOR2_X1 U6089 ( .A(n4930), .B(n4932), .ZN(n4979) );
  OAI21_X1 U6090 ( .B1(n4925), .B2(n4933), .A(n5169), .ZN(n4966) );
  INV_X1 U6091 ( .A(n4966), .ZN(n6316) );
  NOR2_X1 U6092 ( .A1(n6218), .A2(n6319), .ZN(n4975) );
  NOR3_X1 U6093 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6455), .A3(n4934), 
        .ZN(n4935) );
  AOI211_X1 U6094 ( .C1(n6470), .C2(n6316), .A(n4975), .B(n4935), .ZN(n4939)
         );
  INV_X1 U6095 ( .A(n4957), .ZN(n4937) );
  NOR2_X1 U6096 ( .A1(n3614), .A2(n4957), .ZN(n4936) );
  OAI21_X1 U6097 ( .B1(n6216), .B2(n4936), .A(n6466), .ZN(n4959) );
  OAI221_X1 U6098 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n6160), .C1(
        INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n4937), .A(n4959), .ZN(n4938) );
  OAI211_X1 U6099 ( .C1(n6473), .C2(n4979), .A(n4939), .B(n4938), .ZN(U3013)
         );
  XNOR2_X1 U6100 ( .A(n4940), .B(n4942), .ZN(n4974) );
  OAI211_X1 U6101 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5159), .B(n6459), .ZN(n4945) );
  NOR2_X1 U6102 ( .A1(n3588), .A2(n3780), .ZN(n4944) );
  NOR2_X1 U6103 ( .A1(n6218), .A2(n6331), .ZN(n4969) );
  AOI21_X1 U6104 ( .B1(n6470), .B2(n6337), .A(n4969), .ZN(n4943) );
  OAI21_X1 U6105 ( .B1(n4945), .B2(n4944), .A(n4943), .ZN(n4946) );
  AOI21_X1 U6106 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n4947), .A(n4946), 
        .ZN(n4948) );
  OAI21_X1 U6107 ( .B1(n6473), .B2(n4974), .A(n4948), .ZN(U3014) );
  INV_X1 U6108 ( .A(n6352), .ZN(n4952) );
  AOI21_X1 U6109 ( .B1(n6422), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4949), 
        .ZN(n4950) );
  OAI21_X1 U6110 ( .B1(n6351), .B2(n6432), .A(n4950), .ZN(n4951) );
  AOI21_X1 U6111 ( .B1(n4952), .B2(n6065), .A(n4951), .ZN(n4953) );
  OAI21_X1 U6112 ( .B1(n4954), .B2(n6245), .A(n4953), .ZN(U2983) );
  XNOR2_X1 U6113 ( .A(n4955), .B(n4956), .ZN(n5351) );
  NOR3_X1 U6114 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n3614), .A3(n4957), 
        .ZN(n4958) );
  AOI22_X1 U6115 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4959), .B1(n5159), 
        .B2(n4958), .ZN(n4961) );
  XOR2_X1 U6116 ( .A(n5168), .B(n5169), .Z(n6374) );
  NOR2_X1 U6117 ( .A1(n6218), .A2(n6301), .ZN(n5347) );
  AOI21_X1 U6118 ( .B1(n6470), .B2(n6374), .A(n5347), .ZN(n4960) );
  OAI211_X1 U6119 ( .C1(n6473), .C2(n5351), .A(n4961), .B(n4960), .ZN(U3012)
         );
  OR2_X1 U6120 ( .A1(n4923), .A2(n4963), .ZN(n4964) );
  AND2_X1 U6121 ( .A1(n4962), .A2(n4964), .ZN(n6325) );
  INV_X1 U6122 ( .A(n6325), .ZN(n4968) );
  INV_X1 U6123 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6395) );
  OAI222_X1 U6124 ( .A1(n4968), .A2(n5892), .B1(n5891), .B2(n4965), .C1(n5889), 
        .C2(n6395), .ZN(U2886) );
  INV_X1 U6125 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4967) );
  OAI222_X1 U6126 ( .A1(n4968), .A2(n5832), .B1(n6379), .B2(n4967), .C1(n4966), 
        .C2(n5829), .ZN(U2854) );
  INV_X1 U6127 ( .A(n6340), .ZN(n4972) );
  AOI21_X1 U6128 ( .B1(n6422), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4969), 
        .ZN(n4970) );
  OAI21_X1 U6129 ( .B1(n6344), .B2(n6432), .A(n4970), .ZN(n4971) );
  AOI21_X1 U6130 ( .B1(n4972), .B2(n6065), .A(n4971), .ZN(n4973) );
  OAI21_X1 U6131 ( .B1(n6245), .B2(n4974), .A(n4973), .ZN(U2982) );
  AOI21_X1 U6132 ( .B1(n6422), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4975), 
        .ZN(n4976) );
  OAI21_X1 U6133 ( .B1(n6328), .B2(n6432), .A(n4976), .ZN(n4977) );
  AOI21_X1 U6134 ( .B1(n6325), .B2(n6065), .A(n4977), .ZN(n4978) );
  OAI21_X1 U6135 ( .B1(n4979), .B2(n6245), .A(n4978), .ZN(U2981) );
  NOR2_X1 U6136 ( .A1(n4980), .A2(n6639), .ZN(n6724) );
  NAND2_X1 U6137 ( .A1(n6227), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6230) );
  NAND3_X1 U6138 ( .A1(n6724), .A2(n6638), .A3(n6231), .ZN(n4981) );
  NAND2_X1 U6139 ( .A1(n4981), .A2(n6651), .ZN(n4993) );
  INV_X1 U6140 ( .A(n4993), .ZN(n4986) );
  NOR2_X1 U6141 ( .A1(n4714), .A2(n4605), .ZN(n5359) );
  NAND2_X1 U6142 ( .A1(n6721), .A2(n5359), .ZN(n5401) );
  INV_X1 U6143 ( .A(n4623), .ZN(n5784) );
  NAND2_X1 U6144 ( .A1(n6731), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4982) );
  OR2_X1 U6145 ( .A1(n5362), .A2(n4982), .ZN(n5014) );
  NAND2_X1 U6146 ( .A1(n4983), .A2(n5014), .ZN(n4992) );
  NAND3_X1 U6147 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6731), .A3(n4984), .ZN(n5399) );
  INV_X1 U6148 ( .A(n5399), .ZN(n4985) );
  NAND2_X1 U6149 ( .A1(n6231), .A2(n6227), .ZN(n4987) );
  INV_X1 U6150 ( .A(n4988), .ZN(n4989) );
  OAI22_X1 U6151 ( .A1(n5146), .A2(n6587), .B1(n6586), .B2(n5014), .ZN(n4990)
         );
  AOI21_X1 U6152 ( .B1(n6652), .B2(n5433), .A(n4990), .ZN(n4995) );
  NAND2_X1 U6153 ( .A1(n6722), .A2(n5399), .ZN(n4991) );
  NAND2_X1 U6154 ( .A1(n5016), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4994) );
  OAI211_X1 U6155 ( .C1(n5019), .C2(n6655), .A(n4995), .B(n4994), .ZN(U3044)
         );
  OAI22_X1 U6156 ( .A1(n5146), .A2(n6622), .B1(n6621), .B2(n5014), .ZN(n4996)
         );
  AOI21_X1 U6157 ( .B1(n6687), .B2(n5433), .A(n4996), .ZN(n4998) );
  NAND2_X1 U6158 ( .A1(n5016), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4997) );
  OAI211_X1 U6159 ( .C1(n5019), .C2(n6691), .A(n4998), .B(n4997), .ZN(U3050)
         );
  OAI22_X1 U6160 ( .A1(n5146), .A2(n6607), .B1(n6606), .B2(n5014), .ZN(n4999)
         );
  AOI21_X1 U6161 ( .B1(n6669), .B2(n5433), .A(n4999), .ZN(n5001) );
  NAND2_X1 U6162 ( .A1(n5016), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5000) );
  OAI211_X1 U6163 ( .C1(n5019), .C2(n6673), .A(n5001), .B(n5000), .ZN(U3047)
         );
  OAI22_X1 U6164 ( .A1(n5146), .A2(n6561), .B1(n6601), .B2(n5014), .ZN(n5002)
         );
  AOI21_X1 U6165 ( .B1(n6663), .B2(n5433), .A(n5002), .ZN(n5004) );
  NAND2_X1 U6166 ( .A1(n5016), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5003) );
  OAI211_X1 U6167 ( .C1(n5019), .C2(n6667), .A(n5004), .B(n5003), .ZN(U3046)
         );
  OAI22_X1 U6168 ( .A1(n5146), .A2(n6568), .B1(n6611), .B2(n5014), .ZN(n5005)
         );
  AOI21_X1 U6169 ( .B1(n6675), .B2(n5433), .A(n5005), .ZN(n5007) );
  NAND2_X1 U6170 ( .A1(n5016), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5006) );
  OAI211_X1 U6171 ( .C1(n5019), .C2(n6679), .A(n5007), .B(n5006), .ZN(U3048)
         );
  OAI22_X1 U6172 ( .A1(n5146), .A2(n6557), .B1(n6596), .B2(n5014), .ZN(n5008)
         );
  AOI21_X1 U6173 ( .B1(n6658), .B2(n5433), .A(n5008), .ZN(n5010) );
  NAND2_X1 U6174 ( .A1(n5016), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5009) );
  OAI211_X1 U6175 ( .C1(n5019), .C2(n6661), .A(n5010), .B(n5009), .ZN(U3045)
         );
  OAI22_X1 U6176 ( .A1(n5146), .A2(n6617), .B1(n6616), .B2(n5014), .ZN(n5011)
         );
  AOI21_X1 U6177 ( .B1(n6681), .B2(n5433), .A(n5011), .ZN(n5013) );
  NAND2_X1 U6178 ( .A1(n5016), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5012) );
  OAI211_X1 U6179 ( .C1(n5019), .C2(n6685), .A(n5013), .B(n5012), .ZN(U3049)
         );
  OAI22_X1 U6180 ( .A1(n5146), .A2(n6582), .B1(n6628), .B2(n5014), .ZN(n5015)
         );
  AOI21_X1 U6181 ( .B1(n6697), .B2(n5433), .A(n5015), .ZN(n5018) );
  NAND2_X1 U6182 ( .A1(n5016), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5017) );
  OAI211_X1 U6183 ( .C1(n5019), .C2(n6701), .A(n5018), .B(n5017), .ZN(U3051)
         );
  INV_X1 U6184 ( .A(n5020), .ZN(n5028) );
  OAI21_X1 U6185 ( .B1(n6236), .B2(n5525), .A(n6708), .ZN(n5022) );
  AND2_X1 U6186 ( .A1(n6708), .A2(n5021), .ZN(n6705) );
  MUX2_X1 U6187 ( .A(n5022), .B(n6705), .S(STATE2_REG_0__SCAN_IN), .Z(n5027)
         );
  AOI21_X1 U6188 ( .B1(n5025), .B2(n5024), .A(n5023), .ZN(n5026) );
  OAI211_X1 U6189 ( .C1(n5028), .C2(n6711), .A(n5027), .B(n5026), .ZN(U3148)
         );
  NAND2_X1 U6190 ( .A1(n6227), .A2(n6499), .ZN(n5265) );
  NOR3_X1 U6191 ( .A1(n6695), .A2(n5060), .A3(n6722), .ZN(n5030) );
  OAI22_X1 U6192 ( .A1(n5030), .A2(n6728), .B1(n5029), .B2(n5102), .ZN(n5033)
         );
  NAND2_X1 U6193 ( .A1(n5031), .A2(n6541), .ZN(n5057) );
  NOR2_X1 U6194 ( .A1(n5034), .A2(n5179), .ZN(n6546) );
  AOI21_X1 U6195 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5177), .A(n5178), .ZN(
        n5105) );
  OAI21_X1 U6196 ( .B1(n5110), .B2(n5179), .A(n5105), .ZN(n5270) );
  AOI211_X1 U6197 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5057), .A(n6546), .B(
        n5270), .ZN(n5032) );
  NAND2_X1 U6198 ( .A1(n5056), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5037)
         );
  NOR2_X1 U6199 ( .A1(n6721), .A2(n6722), .ZN(n5183) );
  INV_X1 U6200 ( .A(n5102), .ZN(n5109) );
  NAND2_X1 U6201 ( .A1(n5034), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6539) );
  INV_X1 U6202 ( .A(n6539), .ZN(n5364) );
  INV_X1 U6203 ( .A(n5110), .ZN(n5106) );
  NOR2_X1 U6204 ( .A1(n5106), .A2(n5177), .ZN(n5274) );
  AOI22_X1 U6205 ( .A1(n5183), .A2(n5109), .B1(n5364), .B2(n5274), .ZN(n5058)
         );
  OAI22_X1 U6206 ( .A1(n5058), .A2(n6701), .B1(n6628), .B2(n5057), .ZN(n5035)
         );
  AOI21_X1 U6207 ( .B1(n6694), .B2(n5060), .A(n5035), .ZN(n5036) );
  OAI211_X1 U6208 ( .C1(n5063), .C2(n6630), .A(n5037), .B(n5036), .ZN(U3123)
         );
  NAND2_X1 U6209 ( .A1(n5056), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5040)
         );
  OAI22_X1 U6210 ( .A1(n5058), .A2(n6679), .B1(n6611), .B2(n5057), .ZN(n5038)
         );
  AOI21_X1 U6211 ( .B1(n6676), .B2(n5060), .A(n5038), .ZN(n5039) );
  OAI211_X1 U6212 ( .C1(n5063), .C2(n6612), .A(n5040), .B(n5039), .ZN(U3120)
         );
  NAND2_X1 U6213 ( .A1(n5056), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5043)
         );
  OAI22_X1 U6214 ( .A1(n5058), .A2(n6655), .B1(n6586), .B2(n5057), .ZN(n5041)
         );
  AOI21_X1 U6215 ( .B1(n6644), .B2(n5060), .A(n5041), .ZN(n5042) );
  OAI211_X1 U6216 ( .C1(n5063), .C2(n5436), .A(n5043), .B(n5042), .ZN(U3116)
         );
  NAND2_X1 U6217 ( .A1(n5056), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5046)
         );
  OAI22_X1 U6218 ( .A1(n5058), .A2(n6691), .B1(n6621), .B2(n5057), .ZN(n5044)
         );
  AOI21_X1 U6219 ( .B1(n6688), .B2(n5060), .A(n5044), .ZN(n5045) );
  OAI211_X1 U6220 ( .C1(n5063), .C2(n5411), .A(n5046), .B(n5045), .ZN(U3122)
         );
  NAND2_X1 U6221 ( .A1(n5056), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5049)
         );
  OAI22_X1 U6222 ( .A1(n5058), .A2(n6685), .B1(n6616), .B2(n5057), .ZN(n5047)
         );
  AOI21_X1 U6223 ( .B1(n6682), .B2(n5060), .A(n5047), .ZN(n5048) );
  OAI211_X1 U6224 ( .C1(n5063), .C2(n5415), .A(n5049), .B(n5048), .ZN(U3121)
         );
  NAND2_X1 U6225 ( .A1(n5056), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5052)
         );
  OAI22_X1 U6226 ( .A1(n5058), .A2(n6661), .B1(n6596), .B2(n5057), .ZN(n5050)
         );
  AOI21_X1 U6227 ( .B1(n6657), .B2(n5060), .A(n5050), .ZN(n5051) );
  OAI211_X1 U6228 ( .C1(n5063), .C2(n6597), .A(n5052), .B(n5051), .ZN(U3117)
         );
  NAND2_X1 U6229 ( .A1(n5056), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5055)
         );
  OAI22_X1 U6230 ( .A1(n5058), .A2(n6673), .B1(n6606), .B2(n5057), .ZN(n5053)
         );
  AOI21_X1 U6231 ( .B1(n6670), .B2(n5060), .A(n5053), .ZN(n5054) );
  OAI211_X1 U6232 ( .C1(n5063), .C2(n5422), .A(n5055), .B(n5054), .ZN(U3119)
         );
  NAND2_X1 U6233 ( .A1(n5056), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5062)
         );
  OAI22_X1 U6234 ( .A1(n5058), .A2(n6667), .B1(n6601), .B2(n5057), .ZN(n5059)
         );
  AOI21_X1 U6235 ( .B1(n6664), .B2(n5060), .A(n5059), .ZN(n5061) );
  OAI211_X1 U6236 ( .C1(n5063), .C2(n6602), .A(n5062), .B(n5061), .ZN(U3118)
         );
  INV_X1 U6237 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6397) );
  OAI222_X1 U6238 ( .A1(n6340), .A2(n5892), .B1(n5891), .B2(n4835), .C1(n5889), 
        .C2(n6397), .ZN(U2887) );
  INV_X1 U6239 ( .A(n5068), .ZN(n5065) );
  AOI21_X1 U6240 ( .B1(n5065), .B2(STATEBS16_REG_SCAN_IN), .A(n6722), .ZN(
        n5070) );
  OR2_X1 U6241 ( .A1(n4714), .A2(n6363), .ZN(n5216) );
  NOR2_X1 U6242 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6243 ( .A1(n5066), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5071) );
  OR2_X1 U6244 ( .A1(n5071), .A2(n6541), .ZN(n5095) );
  OAI21_X1 U6245 ( .B1(n5067), .B2(n5216), .A(n5095), .ZN(n5073) );
  INV_X1 U6246 ( .A(n5071), .ZN(n5269) );
  OR2_X1 U6247 ( .A1(n5068), .A2(n4807), .ZN(n5367) );
  OAI22_X1 U6248 ( .A1(n5367), .A2(n6568), .B1(n6611), .B2(n5095), .ZN(n5069)
         );
  AOI21_X1 U6249 ( .B1(n6675), .B2(n5266), .A(n5069), .ZN(n5076) );
  INV_X1 U6250 ( .A(n5070), .ZN(n5074) );
  NAND2_X1 U6251 ( .A1(n5071), .A2(n6722), .ZN(n5072) );
  NAND2_X1 U6252 ( .A1(n5097), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n5075) );
  OAI211_X1 U6253 ( .C1(n5100), .C2(n6679), .A(n5076), .B(n5075), .ZN(U3096)
         );
  OAI22_X1 U6254 ( .A1(n5367), .A2(n6617), .B1(n6616), .B2(n5095), .ZN(n5077)
         );
  AOI21_X1 U6255 ( .B1(n6681), .B2(n5266), .A(n5077), .ZN(n5079) );
  NAND2_X1 U6256 ( .A1(n5097), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5078) );
  OAI211_X1 U6257 ( .C1(n5100), .C2(n6685), .A(n5079), .B(n5078), .ZN(U3097)
         );
  OAI22_X1 U6258 ( .A1(n5367), .A2(n6557), .B1(n6596), .B2(n5095), .ZN(n5080)
         );
  AOI21_X1 U6259 ( .B1(n6658), .B2(n5266), .A(n5080), .ZN(n5082) );
  NAND2_X1 U6260 ( .A1(n5097), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n5081) );
  OAI211_X1 U6261 ( .C1(n5100), .C2(n6661), .A(n5082), .B(n5081), .ZN(U3093)
         );
  OAI22_X1 U6262 ( .A1(n5367), .A2(n6587), .B1(n6586), .B2(n5095), .ZN(n5083)
         );
  AOI21_X1 U6263 ( .B1(n6652), .B2(n5266), .A(n5083), .ZN(n5085) );
  NAND2_X1 U6264 ( .A1(n5097), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n5084) );
  OAI211_X1 U6265 ( .C1(n5100), .C2(n6655), .A(n5085), .B(n5084), .ZN(U3092)
         );
  OAI22_X1 U6266 ( .A1(n5367), .A2(n6622), .B1(n6621), .B2(n5095), .ZN(n5086)
         );
  AOI21_X1 U6267 ( .B1(n6687), .B2(n5266), .A(n5086), .ZN(n5088) );
  NAND2_X1 U6268 ( .A1(n5097), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n5087) );
  OAI211_X1 U6269 ( .C1(n5100), .C2(n6691), .A(n5088), .B(n5087), .ZN(U3098)
         );
  OAI22_X1 U6270 ( .A1(n5367), .A2(n6582), .B1(n6628), .B2(n5095), .ZN(n5089)
         );
  AOI21_X1 U6271 ( .B1(n6697), .B2(n5266), .A(n5089), .ZN(n5091) );
  NAND2_X1 U6272 ( .A1(n5097), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n5090) );
  OAI211_X1 U6273 ( .C1(n5100), .C2(n6701), .A(n5091), .B(n5090), .ZN(U3099)
         );
  OAI22_X1 U6274 ( .A1(n5367), .A2(n6607), .B1(n6606), .B2(n5095), .ZN(n5092)
         );
  AOI21_X1 U6275 ( .B1(n6669), .B2(n5266), .A(n5092), .ZN(n5094) );
  NAND2_X1 U6276 ( .A1(n5097), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5093) );
  OAI211_X1 U6277 ( .C1(n5100), .C2(n6673), .A(n5094), .B(n5093), .ZN(U3095)
         );
  OAI22_X1 U6278 ( .A1(n5367), .A2(n6561), .B1(n6601), .B2(n5095), .ZN(n5096)
         );
  AOI21_X1 U6279 ( .B1(n6663), .B2(n5266), .A(n5096), .ZN(n5099) );
  NAND2_X1 U6280 ( .A1(n5097), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n5098) );
  OAI211_X1 U6281 ( .C1(n5100), .C2(n6667), .A(n5099), .B(n5098), .ZN(U3094)
         );
  OAI21_X1 U6282 ( .B1(n6500), .B2(n6722), .A(n5397), .ZN(n6504) );
  NOR2_X1 U6283 ( .A1(n5102), .A2(n6544), .ZN(n6497) );
  INV_X1 U6284 ( .A(n6497), .ZN(n5103) );
  OAI211_X1 U6285 ( .C1(n6728), .C2(n5146), .A(n6504), .B(n5103), .ZN(n5108)
         );
  OR2_X1 U6286 ( .A1(n5104), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6496)
         );
  INV_X1 U6287 ( .A(n6496), .ZN(n6506) );
  NAND2_X1 U6288 ( .A1(n6506), .A2(n6541), .ZN(n5113) );
  OAI21_X1 U6289 ( .B1(n5106), .B2(n5179), .A(n5105), .ZN(n5219) );
  AOI211_X1 U6290 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5113), .A(n6546), .B(
        n5219), .ZN(n5107) );
  NAND2_X1 U6291 ( .A1(n5108), .A2(n5107), .ZN(n5148) );
  NAND2_X1 U6292 ( .A1(n6529), .A2(n6670), .ZN(n5115) );
  NOR2_X1 U6293 ( .A1(n4735), .A2(n6722), .ZN(n6536) );
  NAND2_X1 U6294 ( .A1(n6536), .A2(n5109), .ZN(n5112) );
  NOR2_X1 U6295 ( .A1(n5110), .A2(n5177), .ZN(n5221) );
  NAND2_X1 U6296 ( .A1(n5221), .A2(n5364), .ZN(n5111) );
  NAND2_X1 U6297 ( .A1(n5112), .A2(n5111), .ZN(n5143) );
  INV_X1 U6298 ( .A(n6673), .ZN(n6562) );
  INV_X1 U6299 ( .A(n6606), .ZN(n6668) );
  INV_X1 U6300 ( .A(n5113), .ZN(n5142) );
  AOI22_X1 U6301 ( .A1(n5143), .A2(n6562), .B1(n6668), .B2(n5142), .ZN(n5114)
         );
  OAI211_X1 U6302 ( .C1(n5146), .C2(n5422), .A(n5115), .B(n5114), .ZN(n5116)
         );
  AOI21_X1 U6303 ( .B1(n5148), .B2(INSTQUEUE_REG_4__3__SCAN_IN), .A(n5116), 
        .ZN(n5117) );
  INV_X1 U6304 ( .A(n5117), .ZN(U3055) );
  NAND2_X1 U6305 ( .A1(n6529), .A2(n6682), .ZN(n5119) );
  INV_X1 U6306 ( .A(n6685), .ZN(n6569) );
  INV_X1 U6307 ( .A(n6616), .ZN(n6680) );
  AOI22_X1 U6308 ( .A1(n5143), .A2(n6569), .B1(n6680), .B2(n5142), .ZN(n5118)
         );
  OAI211_X1 U6309 ( .C1(n5146), .C2(n5415), .A(n5119), .B(n5118), .ZN(n5120)
         );
  AOI21_X1 U6310 ( .B1(n5148), .B2(INSTQUEUE_REG_4__5__SCAN_IN), .A(n5120), 
        .ZN(n5121) );
  INV_X1 U6311 ( .A(n5121), .ZN(U3057) );
  NAND2_X1 U6312 ( .A1(n6529), .A2(n6657), .ZN(n5123) );
  INV_X1 U6313 ( .A(n6661), .ZN(n6554) );
  INV_X1 U6314 ( .A(n6596), .ZN(n6656) );
  AOI22_X1 U6315 ( .A1(n5143), .A2(n6554), .B1(n6656), .B2(n5142), .ZN(n5122)
         );
  OAI211_X1 U6316 ( .C1(n5146), .C2(n6597), .A(n5123), .B(n5122), .ZN(n5124)
         );
  AOI21_X1 U6317 ( .B1(n5148), .B2(INSTQUEUE_REG_4__1__SCAN_IN), .A(n5124), 
        .ZN(n5125) );
  INV_X1 U6318 ( .A(n5125), .ZN(U3053) );
  NAND2_X1 U6319 ( .A1(n6529), .A2(n6694), .ZN(n5127) );
  INV_X1 U6320 ( .A(n6701), .ZN(n6576) );
  INV_X1 U6321 ( .A(n6628), .ZN(n6693) );
  AOI22_X1 U6322 ( .A1(n5143), .A2(n6576), .B1(n6693), .B2(n5142), .ZN(n5126)
         );
  OAI211_X1 U6323 ( .C1(n5146), .C2(n6630), .A(n5127), .B(n5126), .ZN(n5128)
         );
  AOI21_X1 U6324 ( .B1(n5148), .B2(INSTQUEUE_REG_4__7__SCAN_IN), .A(n5128), 
        .ZN(n5129) );
  INV_X1 U6325 ( .A(n5129), .ZN(U3059) );
  NAND2_X1 U6326 ( .A1(n6529), .A2(n6644), .ZN(n5131) );
  INV_X1 U6327 ( .A(n6655), .ZN(n6542) );
  INV_X1 U6328 ( .A(n6586), .ZN(n6643) );
  AOI22_X1 U6329 ( .A1(n5143), .A2(n6542), .B1(n6643), .B2(n5142), .ZN(n5130)
         );
  OAI211_X1 U6330 ( .C1(n5146), .C2(n5436), .A(n5131), .B(n5130), .ZN(n5132)
         );
  AOI21_X1 U6331 ( .B1(n5148), .B2(INSTQUEUE_REG_4__0__SCAN_IN), .A(n5132), 
        .ZN(n5133) );
  INV_X1 U6332 ( .A(n5133), .ZN(U3052) );
  NAND2_X1 U6333 ( .A1(n6529), .A2(n6688), .ZN(n5135) );
  INV_X1 U6334 ( .A(n6691), .ZN(n6572) );
  INV_X1 U6335 ( .A(n6621), .ZN(n6686) );
  AOI22_X1 U6336 ( .A1(n5143), .A2(n6572), .B1(n6686), .B2(n5142), .ZN(n5134)
         );
  OAI211_X1 U6337 ( .C1(n5146), .C2(n5411), .A(n5135), .B(n5134), .ZN(n5136)
         );
  AOI21_X1 U6338 ( .B1(n5148), .B2(INSTQUEUE_REG_4__6__SCAN_IN), .A(n5136), 
        .ZN(n5137) );
  INV_X1 U6339 ( .A(n5137), .ZN(U3058) );
  NAND2_X1 U6340 ( .A1(n6529), .A2(n6676), .ZN(n5139) );
  INV_X1 U6341 ( .A(n6679), .ZN(n6565) );
  INV_X1 U6342 ( .A(n6611), .ZN(n6674) );
  AOI22_X1 U6343 ( .A1(n5143), .A2(n6565), .B1(n6674), .B2(n5142), .ZN(n5138)
         );
  OAI211_X1 U6344 ( .C1(n5146), .C2(n6612), .A(n5139), .B(n5138), .ZN(n5140)
         );
  AOI21_X1 U6345 ( .B1(n5148), .B2(INSTQUEUE_REG_4__4__SCAN_IN), .A(n5140), 
        .ZN(n5141) );
  INV_X1 U6346 ( .A(n5141), .ZN(U3056) );
  NAND2_X1 U6347 ( .A1(n6529), .A2(n6664), .ZN(n5145) );
  INV_X1 U6348 ( .A(n6667), .ZN(n6558) );
  INV_X1 U6349 ( .A(n6601), .ZN(n6662) );
  AOI22_X1 U6350 ( .A1(n5143), .A2(n6558), .B1(n6662), .B2(n5142), .ZN(n5144)
         );
  OAI211_X1 U6351 ( .C1(n5146), .C2(n6602), .A(n5145), .B(n5144), .ZN(n5147)
         );
  AOI21_X1 U6352 ( .B1(n5148), .B2(INSTQUEUE_REG_4__2__SCAN_IN), .A(n5147), 
        .ZN(n5149) );
  INV_X1 U6353 ( .A(n5149), .ZN(U3054) );
  XNOR2_X1 U6354 ( .A(n5150), .B(n5151), .ZN(n6062) );
  OAI22_X1 U6355 ( .A1(n5153), .A2(n5152), .B1(n5160), .B2(n6460), .ZN(n5155)
         );
  INV_X1 U6356 ( .A(n5156), .ZN(n5764) );
  NAND2_X1 U6357 ( .A1(n5170), .A2(n5157), .ZN(n5158) );
  NAND2_X1 U6358 ( .A1(n5764), .A2(n5158), .ZN(n6286) );
  NAND2_X1 U6359 ( .A1(n6457), .A2(REIP_REG_8__SCAN_IN), .ZN(n6055) );
  OAI21_X1 U6360 ( .B1(n6221), .B2(n6286), .A(n6055), .ZN(n5162) );
  NAND2_X1 U6361 ( .A1(n5160), .A2(n5159), .ZN(n6446) );
  AOI211_X1 U6362 ( .C1(n6930), .C2(n3793), .A(n6217), .B(n6446), .ZN(n5161)
         );
  AOI211_X1 U6363 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n6215), .A(n5162), 
        .B(n5161), .ZN(n5163) );
  OAI21_X1 U6364 ( .B1(n6473), .B2(n6062), .A(n5163), .ZN(U3010) );
  INV_X1 U6365 ( .A(n5164), .ZN(n5322) );
  OAI21_X1 U6366 ( .B1(n5322), .B2(n3943), .A(n5166), .ZN(n6295) );
  OAI21_X1 U6367 ( .B1(n5169), .B2(n5168), .A(n5167), .ZN(n5171) );
  AND2_X1 U6368 ( .A1(n5171), .A2(n5170), .ZN(n6442) );
  AOI22_X1 U6369 ( .A1(n6375), .A2(n6442), .B1(EBX_REG_7__SCAN_IN), .B2(n5830), 
        .ZN(n5172) );
  OAI21_X1 U6370 ( .B1(n6295), .B2(n5832), .A(n5172), .ZN(U2852) );
  INV_X1 U6371 ( .A(n5212), .ZN(n5174) );
  NOR3_X1 U6372 ( .A1(n5174), .A2(n5209), .A3(n6722), .ZN(n5175) );
  OAI22_X1 U6373 ( .A1(n5175), .A2(n6728), .B1(n6721), .B2(n6545), .ZN(n5181)
         );
  OR2_X1 U6374 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5176), .ZN(n5206)
         );
  INV_X1 U6375 ( .A(n5177), .ZN(n5402) );
  OAI21_X1 U6376 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n5179), .A(n6549), 
        .ZN(n5363) );
  AOI211_X1 U6377 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5206), .A(n6546), .B(
        n5363), .ZN(n5180) );
  NAND2_X1 U6378 ( .A1(n5205), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5186)
         );
  INV_X1 U6379 ( .A(n6545), .ZN(n5182) );
  NOR2_X1 U6380 ( .A1(n5402), .A2(n6731), .ZN(n5360) );
  AOI22_X1 U6381 ( .A1(n5183), .A2(n5182), .B1(n5364), .B2(n5360), .ZN(n5207)
         );
  OAI22_X1 U6382 ( .A1(n5207), .A2(n6685), .B1(n6616), .B2(n5206), .ZN(n5184)
         );
  AOI21_X1 U6383 ( .B1(n6681), .B2(n5209), .A(n5184), .ZN(n5185) );
  OAI211_X1 U6384 ( .C1(n5212), .C2(n6617), .A(n5186), .B(n5185), .ZN(U3137)
         );
  NAND2_X1 U6385 ( .A1(n5205), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5189)
         );
  OAI22_X1 U6386 ( .A1(n5207), .A2(n6667), .B1(n6601), .B2(n5206), .ZN(n5187)
         );
  AOI21_X1 U6387 ( .B1(n6663), .B2(n5209), .A(n5187), .ZN(n5188) );
  OAI211_X1 U6388 ( .C1(n5212), .C2(n6561), .A(n5189), .B(n5188), .ZN(U3134)
         );
  NAND2_X1 U6389 ( .A1(n5205), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5192)
         );
  OAI22_X1 U6390 ( .A1(n5207), .A2(n6661), .B1(n6596), .B2(n5206), .ZN(n5190)
         );
  AOI21_X1 U6391 ( .B1(n6658), .B2(n5209), .A(n5190), .ZN(n5191) );
  OAI211_X1 U6392 ( .C1(n5212), .C2(n6557), .A(n5192), .B(n5191), .ZN(U3133)
         );
  NAND2_X1 U6393 ( .A1(n5205), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5195)
         );
  OAI22_X1 U6394 ( .A1(n5207), .A2(n6701), .B1(n6628), .B2(n5206), .ZN(n5193)
         );
  AOI21_X1 U6395 ( .B1(n6697), .B2(n5209), .A(n5193), .ZN(n5194) );
  OAI211_X1 U6396 ( .C1(n5212), .C2(n6582), .A(n5195), .B(n5194), .ZN(U3139)
         );
  NAND2_X1 U6397 ( .A1(n5205), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5198)
         );
  OAI22_X1 U6398 ( .A1(n5207), .A2(n6679), .B1(n6611), .B2(n5206), .ZN(n5196)
         );
  AOI21_X1 U6399 ( .B1(n6675), .B2(n5209), .A(n5196), .ZN(n5197) );
  OAI211_X1 U6400 ( .C1(n5212), .C2(n6568), .A(n5198), .B(n5197), .ZN(U3136)
         );
  NAND2_X1 U6401 ( .A1(n5205), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5201)
         );
  OAI22_X1 U6402 ( .A1(n5207), .A2(n6691), .B1(n6621), .B2(n5206), .ZN(n5199)
         );
  AOI21_X1 U6403 ( .B1(n6687), .B2(n5209), .A(n5199), .ZN(n5200) );
  OAI211_X1 U6404 ( .C1(n5212), .C2(n6622), .A(n5201), .B(n5200), .ZN(U3138)
         );
  NAND2_X1 U6405 ( .A1(n5205), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5204)
         );
  OAI22_X1 U6406 ( .A1(n5207), .A2(n6655), .B1(n6586), .B2(n5206), .ZN(n5202)
         );
  AOI21_X1 U6407 ( .B1(n6652), .B2(n5209), .A(n5202), .ZN(n5203) );
  OAI211_X1 U6408 ( .C1(n5212), .C2(n6587), .A(n5204), .B(n5203), .ZN(U3132)
         );
  NAND2_X1 U6409 ( .A1(n5205), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5211)
         );
  OAI22_X1 U6410 ( .A1(n5207), .A2(n6673), .B1(n6606), .B2(n5206), .ZN(n5208)
         );
  AOI21_X1 U6411 ( .B1(n6669), .B2(n5209), .A(n5208), .ZN(n5210) );
  OAI211_X1 U6412 ( .C1(n5212), .C2(n6607), .A(n5211), .B(n5210), .ZN(U3135)
         );
  NAND2_X1 U6413 ( .A1(n6231), .A2(n5213), .ZN(n5214) );
  NAND2_X1 U6414 ( .A1(n5253), .A2(n6651), .ZN(n5215) );
  OAI21_X1 U6415 ( .B1(n6490), .B2(n5215), .A(n5397), .ZN(n5220) );
  NAND2_X1 U6416 ( .A1(n6721), .A2(n5267), .ZN(n5304) );
  NOR3_X1 U6417 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5311) );
  AND2_X1 U6418 ( .A1(n6541), .A2(n5311), .ZN(n5222) );
  OAI21_X1 U6419 ( .B1(n5222), .B2(n5217), .A(n6539), .ZN(n5218) );
  INV_X1 U6420 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5226) );
  AOI22_X1 U6421 ( .A1(n6536), .A2(n5267), .B1(n6546), .B2(n5221), .ZN(n5252)
         );
  INV_X1 U6422 ( .A(n5222), .ZN(n5251) );
  OAI22_X1 U6423 ( .A1(n5252), .A2(n6679), .B1(n6611), .B2(n5251), .ZN(n5224)
         );
  NOR2_X1 U6424 ( .A1(n5253), .A2(n6612), .ZN(n5223) );
  AOI211_X1 U6425 ( .C1(n6490), .C2(n6676), .A(n5224), .B(n5223), .ZN(n5225)
         );
  OAI21_X1 U6426 ( .B1(n5258), .B2(n5226), .A(n5225), .ZN(U3024) );
  OAI22_X1 U6427 ( .A1(n5252), .A2(n6701), .B1(n6628), .B2(n5251), .ZN(n5228)
         );
  NOR2_X1 U6428 ( .A1(n5253), .A2(n6630), .ZN(n5227) );
  AOI211_X1 U6429 ( .C1(n6490), .C2(n6694), .A(n5228), .B(n5227), .ZN(n5229)
         );
  OAI21_X1 U6430 ( .B1(n5258), .B2(n5230), .A(n5229), .ZN(U3027) );
  INV_X1 U6431 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5234) );
  OAI22_X1 U6432 ( .A1(n5252), .A2(n6691), .B1(n6621), .B2(n5251), .ZN(n5232)
         );
  NOR2_X1 U6433 ( .A1(n5253), .A2(n5411), .ZN(n5231) );
  AOI211_X1 U6434 ( .C1(n6490), .C2(n6688), .A(n5232), .B(n5231), .ZN(n5233)
         );
  OAI21_X1 U6435 ( .B1(n5258), .B2(n5234), .A(n5233), .ZN(U3026) );
  OAI22_X1 U6436 ( .A1(n5252), .A2(n6655), .B1(n6586), .B2(n5251), .ZN(n5236)
         );
  NOR2_X1 U6437 ( .A1(n5253), .A2(n5436), .ZN(n5235) );
  AOI211_X1 U6438 ( .C1(n6490), .C2(n6644), .A(n5236), .B(n5235), .ZN(n5237)
         );
  OAI21_X1 U6439 ( .B1(n5258), .B2(n5238), .A(n5237), .ZN(U3020) );
  INV_X1 U6440 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5242) );
  OAI22_X1 U6441 ( .A1(n5252), .A2(n6685), .B1(n6616), .B2(n5251), .ZN(n5240)
         );
  NOR2_X1 U6442 ( .A1(n5253), .A2(n5415), .ZN(n5239) );
  AOI211_X1 U6443 ( .C1(n6490), .C2(n6682), .A(n5240), .B(n5239), .ZN(n5241)
         );
  OAI21_X1 U6444 ( .B1(n5258), .B2(n5242), .A(n5241), .ZN(U3025) );
  INV_X1 U6445 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5246) );
  OAI22_X1 U6446 ( .A1(n5252), .A2(n6673), .B1(n6606), .B2(n5251), .ZN(n5244)
         );
  NOR2_X1 U6447 ( .A1(n5253), .A2(n5422), .ZN(n5243) );
  AOI211_X1 U6448 ( .C1(n6490), .C2(n6670), .A(n5244), .B(n5243), .ZN(n5245)
         );
  OAI21_X1 U6449 ( .B1(n5258), .B2(n5246), .A(n5245), .ZN(U3023) );
  OAI22_X1 U6450 ( .A1(n5252), .A2(n6661), .B1(n6596), .B2(n5251), .ZN(n5248)
         );
  NOR2_X1 U6451 ( .A1(n5253), .A2(n6597), .ZN(n5247) );
  AOI211_X1 U6452 ( .C1(n6490), .C2(n6657), .A(n5248), .B(n5247), .ZN(n5249)
         );
  OAI21_X1 U6453 ( .B1(n5258), .B2(n5250), .A(n5249), .ZN(U3021) );
  OAI22_X1 U6454 ( .A1(n5252), .A2(n6667), .B1(n6601), .B2(n5251), .ZN(n5255)
         );
  NOR2_X1 U6455 ( .A1(n5253), .A2(n6602), .ZN(n5254) );
  AOI211_X1 U6456 ( .C1(n6490), .C2(n6664), .A(n5255), .B(n5254), .ZN(n5256)
         );
  OAI21_X1 U6457 ( .B1(n5258), .B2(n5257), .A(n5256), .ZN(U3022) );
  INV_X1 U6458 ( .A(n5260), .ZN(n5261) );
  XNOR2_X1 U6459 ( .A(n5259), .B(n5261), .ZN(n6443) );
  NAND2_X1 U6460 ( .A1(n6443), .A2(n6428), .ZN(n5264) );
  NOR2_X1 U6461 ( .A1(n6218), .A2(n7009), .ZN(n6441) );
  NOR2_X1 U6462 ( .A1(n6432), .A2(n6305), .ZN(n5262) );
  AOI211_X1 U6463 ( .C1(n6422), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6441), 
        .B(n5262), .ZN(n5263) );
  OAI211_X1 U6464 ( .C1(n6057), .C2(n6295), .A(n5264), .B(n5263), .ZN(U2979)
         );
  OAI222_X1 U6465 ( .A1(n6295), .A2(n5892), .B1(n5891), .B2(n4831), .C1(n5889), 
        .C2(n6784), .ZN(U2884) );
  OAI21_X1 U6466 ( .B1(n5266), .B2(n6633), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5268) );
  NAND2_X1 U6467 ( .A1(n5267), .A2(n4735), .ZN(n5273) );
  NAND3_X1 U6468 ( .A1(n5268), .A2(n6651), .A3(n5273), .ZN(n5272) );
  NAND2_X1 U6469 ( .A1(n5269), .A2(n6541), .ZN(n5298) );
  AOI211_X1 U6470 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5298), .A(n5364), .B(
        n5270), .ZN(n5271) );
  NAND2_X1 U6471 ( .A1(n5297), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5278) );
  INV_X1 U6472 ( .A(n5273), .ZN(n5275) );
  AOI22_X1 U6473 ( .A1(n5275), .A2(n6651), .B1(n6546), .B2(n5274), .ZN(n5299)
         );
  OAI22_X1 U6474 ( .A1(n5299), .A2(n6673), .B1(n6606), .B2(n5298), .ZN(n5276)
         );
  AOI21_X1 U6475 ( .B1(n6633), .B2(n6669), .A(n5276), .ZN(n5277) );
  OAI211_X1 U6476 ( .C1(n5303), .C2(n6607), .A(n5278), .B(n5277), .ZN(U3087)
         );
  NAND2_X1 U6477 ( .A1(n5297), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5281) );
  OAI22_X1 U6478 ( .A1(n5299), .A2(n6679), .B1(n6611), .B2(n5298), .ZN(n5279)
         );
  AOI21_X1 U6479 ( .B1(n6633), .B2(n6675), .A(n5279), .ZN(n5280) );
  OAI211_X1 U6480 ( .C1(n5303), .C2(n6568), .A(n5281), .B(n5280), .ZN(U3088)
         );
  NAND2_X1 U6481 ( .A1(n5297), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5284) );
  OAI22_X1 U6482 ( .A1(n5299), .A2(n6685), .B1(n6616), .B2(n5298), .ZN(n5282)
         );
  AOI21_X1 U6483 ( .B1(n6633), .B2(n6681), .A(n5282), .ZN(n5283) );
  OAI211_X1 U6484 ( .C1(n5303), .C2(n6617), .A(n5284), .B(n5283), .ZN(U3089)
         );
  NAND2_X1 U6485 ( .A1(n5297), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5287) );
  OAI22_X1 U6486 ( .A1(n5299), .A2(n6655), .B1(n6586), .B2(n5298), .ZN(n5285)
         );
  AOI21_X1 U6487 ( .B1(n6633), .B2(n6652), .A(n5285), .ZN(n5286) );
  OAI211_X1 U6488 ( .C1(n5303), .C2(n6587), .A(n5287), .B(n5286), .ZN(U3084)
         );
  NAND2_X1 U6489 ( .A1(n5297), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5290) );
  OAI22_X1 U6490 ( .A1(n5299), .A2(n6691), .B1(n6621), .B2(n5298), .ZN(n5288)
         );
  AOI21_X1 U6491 ( .B1(n6633), .B2(n6687), .A(n5288), .ZN(n5289) );
  OAI211_X1 U6492 ( .C1(n5303), .C2(n6622), .A(n5290), .B(n5289), .ZN(U3090)
         );
  NAND2_X1 U6493 ( .A1(n5297), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5293) );
  OAI22_X1 U6494 ( .A1(n5299), .A2(n6661), .B1(n6596), .B2(n5298), .ZN(n5291)
         );
  AOI21_X1 U6495 ( .B1(n6633), .B2(n6658), .A(n5291), .ZN(n5292) );
  OAI211_X1 U6496 ( .C1(n5303), .C2(n6557), .A(n5293), .B(n5292), .ZN(U3085)
         );
  NAND2_X1 U6497 ( .A1(n5297), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5296) );
  OAI22_X1 U6498 ( .A1(n5299), .A2(n6667), .B1(n6601), .B2(n5298), .ZN(n5294)
         );
  AOI21_X1 U6499 ( .B1(n6633), .B2(n6663), .A(n5294), .ZN(n5295) );
  OAI211_X1 U6500 ( .C1(n5303), .C2(n6561), .A(n5296), .B(n5295), .ZN(U3086)
         );
  NAND2_X1 U6501 ( .A1(n5297), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5302) );
  OAI22_X1 U6502 ( .A1(n5299), .A2(n6701), .B1(n6628), .B2(n5298), .ZN(n5300)
         );
  AOI21_X1 U6503 ( .B1(n6633), .B2(n6697), .A(n5300), .ZN(n5301) );
  OAI211_X1 U6504 ( .C1(n5303), .C2(n6582), .A(n5302), .B(n5301), .ZN(U3091)
         );
  INV_X1 U6505 ( .A(n5311), .ZN(n5307) );
  OAI21_X1 U6506 ( .B1(n5308), .B2(n6244), .A(n6651), .ZN(n5310) );
  NAND2_X1 U6507 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5311), .ZN(n6488) );
  OAI21_X1 U6508 ( .B1(n5304), .B2(n5784), .A(n6488), .ZN(n5312) );
  NOR2_X1 U6509 ( .A1(n5310), .A2(n5312), .ZN(n5305) );
  INV_X1 U6510 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n6783) );
  NOR2_X1 U6511 ( .A1(n5308), .A2(n4807), .ZN(n6491) );
  NAND2_X1 U6512 ( .A1(n6491), .A2(n6644), .ZN(n5309) );
  OAI21_X1 U6513 ( .B1(n6488), .B2(n6586), .A(n5309), .ZN(n5315) );
  INV_X1 U6514 ( .A(n5310), .ZN(n5313) );
  AOI22_X1 U6515 ( .A1(n5313), .A2(n5312), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5311), .ZN(n6484) );
  NOR2_X1 U6516 ( .A1(n6484), .A2(n6655), .ZN(n5314) );
  AOI211_X1 U6517 ( .C1(n6490), .C2(n6652), .A(n5315), .B(n5314), .ZN(n5316)
         );
  OAI21_X1 U6518 ( .B1(n6495), .B2(n6783), .A(n5316), .ZN(U3028) );
  INV_X1 U6519 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6520 ( .A1(n6491), .A2(n6676), .ZN(n5317) );
  OAI21_X1 U6521 ( .B1(n6488), .B2(n6611), .A(n5317), .ZN(n5319) );
  NOR2_X1 U6522 ( .A1(n6484), .A2(n6679), .ZN(n5318) );
  AOI211_X1 U6523 ( .C1(n6490), .C2(n6675), .A(n5319), .B(n5318), .ZN(n5320)
         );
  OAI21_X1 U6524 ( .B1(n6495), .B2(n5321), .A(n5320), .ZN(U3032) );
  AOI21_X1 U6525 ( .B1(n5323), .B2(n4962), .A(n5322), .ZN(n6377) );
  INV_X1 U6526 ( .A(n6377), .ZN(n5326) );
  OAI222_X1 U6527 ( .A1(n5326), .A2(n5892), .B1(n5889), .B2(n5325), .C1(n5891), 
        .C2(n5324), .ZN(U2885) );
  INV_X1 U6528 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6529 ( .A1(n6491), .A2(n6682), .ZN(n5327) );
  OAI21_X1 U6530 ( .B1(n6488), .B2(n6616), .A(n5327), .ZN(n5329) );
  NOR2_X1 U6531 ( .A1(n6484), .A2(n6685), .ZN(n5328) );
  AOI211_X1 U6532 ( .C1(n6490), .C2(n6681), .A(n5329), .B(n5328), .ZN(n5330)
         );
  OAI21_X1 U6533 ( .B1(n6495), .B2(n5331), .A(n5330), .ZN(U3033) );
  INV_X1 U6534 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6535 ( .A1(n6491), .A2(n6670), .ZN(n5332) );
  OAI21_X1 U6536 ( .B1(n6488), .B2(n6606), .A(n5332), .ZN(n5334) );
  NOR2_X1 U6537 ( .A1(n6484), .A2(n6673), .ZN(n5333) );
  AOI211_X1 U6538 ( .C1(n6490), .C2(n6669), .A(n5334), .B(n5333), .ZN(n5335)
         );
  OAI21_X1 U6539 ( .B1(n6495), .B2(n5336), .A(n5335), .ZN(U3031) );
  INV_X1 U6540 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6541 ( .A1(n6491), .A2(n6694), .ZN(n5337) );
  OAI21_X1 U6542 ( .B1(n6488), .B2(n6628), .A(n5337), .ZN(n5339) );
  NOR2_X1 U6543 ( .A1(n6484), .A2(n6701), .ZN(n5338) );
  AOI211_X1 U6544 ( .C1(n6490), .C2(n6697), .A(n5339), .B(n5338), .ZN(n5340)
         );
  OAI21_X1 U6545 ( .B1(n6495), .B2(n5341), .A(n5340), .ZN(U3035) );
  INV_X1 U6546 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6547 ( .A1(n6491), .A2(n6688), .ZN(n5342) );
  OAI21_X1 U6548 ( .B1(n6488), .B2(n6621), .A(n5342), .ZN(n5344) );
  NOR2_X1 U6549 ( .A1(n6484), .A2(n6691), .ZN(n5343) );
  AOI211_X1 U6550 ( .C1(n6490), .C2(n6687), .A(n5344), .B(n5343), .ZN(n5345)
         );
  OAI21_X1 U6551 ( .B1(n6495), .B2(n5346), .A(n5345), .ZN(U3034) );
  AOI21_X1 U6552 ( .B1(n6422), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5347), 
        .ZN(n5348) );
  OAI21_X1 U6553 ( .B1(n6309), .B2(n6432), .A(n5348), .ZN(n5349) );
  AOI21_X1 U6554 ( .B1(n6377), .B2(n6065), .A(n5349), .ZN(n5350) );
  OAI21_X1 U6555 ( .B1(n6245), .B2(n5351), .A(n5350), .ZN(U2980) );
  AND2_X1 U6556 ( .A1(n5166), .A2(n5352), .ZN(n5354) );
  OR2_X1 U6557 ( .A1(n5354), .A2(n5353), .ZN(n6288) );
  INV_X1 U6558 ( .A(n5891), .ZN(n5886) );
  AOI22_X1 U6559 ( .A1(n5886), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n5885), .ZN(n5355) );
  OAI21_X1 U6560 ( .B1(n6288), .B2(n5892), .A(n5355), .ZN(U2883) );
  INV_X1 U6561 ( .A(n6286), .ZN(n5356) );
  AOI22_X1 U6562 ( .A1(n5356), .A2(n6375), .B1(n5830), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5357) );
  OAI21_X1 U6563 ( .B1(n6288), .B2(n5832), .A(n5357), .ZN(U2851) );
  AND2_X1 U6564 ( .A1(n6227), .A2(n4807), .ZN(n6534) );
  NOR2_X1 U6565 ( .A1(n6696), .A2(n6722), .ZN(n5358) );
  AOI21_X1 U6566 ( .B1(n5358), .B2(n5367), .A(n6728), .ZN(n5366) );
  INV_X1 U6567 ( .A(n5366), .ZN(n5361) );
  NOR2_X1 U6568 ( .A1(n5362), .A2(n6731), .ZN(n6650) );
  NAND2_X1 U6569 ( .A1(n6650), .A2(n6541), .ZN(n5390) );
  AOI211_X1 U6570 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5390), .A(n5364), .B(
        n5363), .ZN(n5365) );
  NAND2_X1 U6571 ( .A1(n5389), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5370)
         );
  OAI22_X1 U6572 ( .A1(n5391), .A2(n6622), .B1(n5390), .B2(n6621), .ZN(n5368)
         );
  AOI21_X1 U6573 ( .B1(n5393), .B2(n6687), .A(n5368), .ZN(n5369) );
  OAI211_X1 U6574 ( .C1(n5396), .C2(n6691), .A(n5370), .B(n5369), .ZN(U3106)
         );
  NAND2_X1 U6575 ( .A1(n5389), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5373)
         );
  OAI22_X1 U6576 ( .A1(n5391), .A2(n6561), .B1(n5390), .B2(n6601), .ZN(n5371)
         );
  AOI21_X1 U6577 ( .B1(n5393), .B2(n6663), .A(n5371), .ZN(n5372) );
  OAI211_X1 U6578 ( .C1(n5396), .C2(n6667), .A(n5373), .B(n5372), .ZN(U3102)
         );
  NAND2_X1 U6579 ( .A1(n5389), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5376)
         );
  OAI22_X1 U6580 ( .A1(n5391), .A2(n6607), .B1(n5390), .B2(n6606), .ZN(n5374)
         );
  AOI21_X1 U6581 ( .B1(n5393), .B2(n6669), .A(n5374), .ZN(n5375) );
  OAI211_X1 U6582 ( .C1(n5396), .C2(n6673), .A(n5376), .B(n5375), .ZN(U3103)
         );
  NAND2_X1 U6583 ( .A1(n5389), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5379)
         );
  OAI22_X1 U6584 ( .A1(n5391), .A2(n6582), .B1(n5390), .B2(n6628), .ZN(n5377)
         );
  AOI21_X1 U6585 ( .B1(n5393), .B2(n6697), .A(n5377), .ZN(n5378) );
  OAI211_X1 U6586 ( .C1(n5396), .C2(n6701), .A(n5379), .B(n5378), .ZN(U3107)
         );
  NAND2_X1 U6587 ( .A1(n5389), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5382)
         );
  OAI22_X1 U6588 ( .A1(n5391), .A2(n6557), .B1(n5390), .B2(n6596), .ZN(n5380)
         );
  AOI21_X1 U6589 ( .B1(n5393), .B2(n6658), .A(n5380), .ZN(n5381) );
  OAI211_X1 U6590 ( .C1(n5396), .C2(n6661), .A(n5382), .B(n5381), .ZN(U3101)
         );
  NAND2_X1 U6591 ( .A1(n5389), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5385)
         );
  OAI22_X1 U6592 ( .A1(n5391), .A2(n6587), .B1(n5390), .B2(n6586), .ZN(n5383)
         );
  AOI21_X1 U6593 ( .B1(n5393), .B2(n6652), .A(n5383), .ZN(n5384) );
  OAI211_X1 U6594 ( .C1(n5396), .C2(n6655), .A(n5385), .B(n5384), .ZN(U3100)
         );
  NAND2_X1 U6595 ( .A1(n5389), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5388)
         );
  OAI22_X1 U6596 ( .A1(n5391), .A2(n6617), .B1(n5390), .B2(n6616), .ZN(n5386)
         );
  AOI21_X1 U6597 ( .B1(n5393), .B2(n6681), .A(n5386), .ZN(n5387) );
  OAI211_X1 U6598 ( .C1(n5396), .C2(n6685), .A(n5388), .B(n5387), .ZN(U3105)
         );
  NAND2_X1 U6599 ( .A1(n5389), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5395)
         );
  OAI22_X1 U6600 ( .A1(n5391), .A2(n6568), .B1(n5390), .B2(n6611), .ZN(n5392)
         );
  AOI21_X1 U6601 ( .B1(n5393), .B2(n6675), .A(n5392), .ZN(n5394) );
  OAI211_X1 U6602 ( .C1(n5396), .C2(n6679), .A(n5395), .B(n5394), .ZN(U3104)
         );
  OAI21_X1 U6603 ( .B1(n6491), .B2(n5433), .A(n5397), .ZN(n5398) );
  AOI21_X1 U6604 ( .B1(n5398), .B2(n5401), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5400) );
  NOR2_X1 U6605 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5399), .ZN(n5404)
         );
  NAND2_X1 U6606 ( .A1(n5429), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5407) );
  INV_X1 U6607 ( .A(n5401), .ZN(n5403) );
  NOR2_X1 U6608 ( .A1(n5402), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6537)
         );
  AOI22_X1 U6609 ( .A1(n5403), .A2(n6651), .B1(n6546), .B2(n6537), .ZN(n5431)
         );
  INV_X1 U6610 ( .A(n5404), .ZN(n5430) );
  OAI22_X1 U6611 ( .A1(n5431), .A2(n6701), .B1(n6628), .B2(n5430), .ZN(n5405)
         );
  AOI21_X1 U6612 ( .B1(n5433), .B2(n6694), .A(n5405), .ZN(n5406) );
  OAI211_X1 U6613 ( .C1(n5437), .C2(n6630), .A(n5407), .B(n5406), .ZN(U3043)
         );
  NAND2_X1 U6614 ( .A1(n5429), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5410) );
  OAI22_X1 U6615 ( .A1(n5431), .A2(n6691), .B1(n6621), .B2(n5430), .ZN(n5408)
         );
  AOI21_X1 U6616 ( .B1(n5433), .B2(n6688), .A(n5408), .ZN(n5409) );
  OAI211_X1 U6617 ( .C1(n5437), .C2(n5411), .A(n5410), .B(n5409), .ZN(U3042)
         );
  NAND2_X1 U6618 ( .A1(n5429), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5414) );
  OAI22_X1 U6619 ( .A1(n5431), .A2(n6685), .B1(n6616), .B2(n5430), .ZN(n5412)
         );
  AOI21_X1 U6620 ( .B1(n5433), .B2(n6682), .A(n5412), .ZN(n5413) );
  OAI211_X1 U6621 ( .C1(n5437), .C2(n5415), .A(n5414), .B(n5413), .ZN(U3041)
         );
  NAND2_X1 U6622 ( .A1(n5429), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5418) );
  OAI22_X1 U6623 ( .A1(n5431), .A2(n6679), .B1(n6611), .B2(n5430), .ZN(n5416)
         );
  AOI21_X1 U6624 ( .B1(n5433), .B2(n6676), .A(n5416), .ZN(n5417) );
  OAI211_X1 U6625 ( .C1(n5437), .C2(n6612), .A(n5418), .B(n5417), .ZN(U3040)
         );
  NAND2_X1 U6626 ( .A1(n5429), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5421) );
  OAI22_X1 U6627 ( .A1(n5431), .A2(n6673), .B1(n6606), .B2(n5430), .ZN(n5419)
         );
  AOI21_X1 U6628 ( .B1(n5433), .B2(n6670), .A(n5419), .ZN(n5420) );
  OAI211_X1 U6629 ( .C1(n5437), .C2(n5422), .A(n5421), .B(n5420), .ZN(U3039)
         );
  NAND2_X1 U6630 ( .A1(n5429), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5425) );
  OAI22_X1 U6631 ( .A1(n5431), .A2(n6667), .B1(n6601), .B2(n5430), .ZN(n5423)
         );
  AOI21_X1 U6632 ( .B1(n5433), .B2(n6664), .A(n5423), .ZN(n5424) );
  OAI211_X1 U6633 ( .C1(n5437), .C2(n6602), .A(n5425), .B(n5424), .ZN(U3038)
         );
  NAND2_X1 U6634 ( .A1(n5429), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5428) );
  OAI22_X1 U6635 ( .A1(n5431), .A2(n6661), .B1(n6596), .B2(n5430), .ZN(n5426)
         );
  AOI21_X1 U6636 ( .B1(n5433), .B2(n6657), .A(n5426), .ZN(n5427) );
  OAI211_X1 U6637 ( .C1(n5437), .C2(n6597), .A(n5428), .B(n5427), .ZN(U3037)
         );
  NAND2_X1 U6638 ( .A1(n5429), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5435) );
  OAI22_X1 U6639 ( .A1(n5431), .A2(n6655), .B1(n6586), .B2(n5430), .ZN(n5432)
         );
  AOI21_X1 U6640 ( .B1(n5433), .B2(n6644), .A(n5432), .ZN(n5434) );
  OAI211_X1 U6641 ( .C1(n5437), .C2(n5436), .A(n5435), .B(n5434), .ZN(U3036)
         );
  INV_X1 U6642 ( .A(n5514), .ZN(n5449) );
  INV_X1 U6643 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5438) );
  NAND4_X1 U6644 ( .A1(n5439), .A2(REIP_REG_29__SCAN_IN), .A3(
        REIP_REG_30__SCAN_IN), .A4(n5438), .ZN(n5446) );
  OAI211_X1 U6645 ( .C1(n5441), .C2(n5440), .A(REIP_REG_31__SCAN_IN), .B(n6329), .ZN(n5445) );
  NAND2_X1 U6646 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5444)
         );
  NAND3_X1 U6647 ( .A1(n5779), .A2(EBX_REG_31__SCAN_IN), .A3(n5442), .ZN(n5443) );
  NAND4_X1 U6648 ( .A1(n5446), .A2(n5445), .A3(n5444), .A4(n5443), .ZN(n5447)
         );
  AOI21_X1 U6649 ( .B1(n5789), .B2(n6361), .A(n5447), .ZN(n5448) );
  OAI21_X1 U6650 ( .B1(n5449), .B2(n5780), .A(n5448), .ZN(U2796) );
  XNOR2_X1 U6651 ( .A(n4300), .B(n5452), .ZN(n5956) );
  XNOR2_X1 U6652 ( .A(n4300), .B(n5455), .ZN(n5946) );
  XNOR2_X1 U6653 ( .A(n4300), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5937)
         );
  INV_X1 U6654 ( .A(n5937), .ZN(n5456) );
  OR2_X1 U6655 ( .A1(n5946), .A2(n5456), .ZN(n5454) );
  NAND2_X1 U6656 ( .A1(n4300), .A2(n5455), .ZN(n5934) );
  INV_X1 U6657 ( .A(n5926), .ZN(n5460) );
  NAND2_X1 U6658 ( .A1(n5460), .A2(n5459), .ZN(n5463) );
  NAND2_X1 U6659 ( .A1(n3080), .A2(n6855), .ZN(n5925) );
  INV_X1 U6660 ( .A(n5925), .ZN(n5461) );
  XNOR2_X1 U6661 ( .A(n5464), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5478)
         );
  NOR2_X1 U6662 ( .A1(n5466), .A2(n5467), .ZN(n5468) );
  INV_X1 U6663 ( .A(n5854), .ZN(n5471) );
  NAND2_X1 U6664 ( .A1(n6457), .A2(REIP_REG_24__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6665 ( .A1(n6422), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5469)
         );
  OAI211_X1 U6666 ( .C1(n6432), .C2(n5586), .A(n5474), .B(n5469), .ZN(n5470)
         );
  AOI21_X1 U6667 ( .B1(n5471), .B2(n6065), .A(n5470), .ZN(n5472) );
  OAI21_X1 U6668 ( .B1(n5478), .B2(n6245), .A(n5472), .ZN(U2962) );
  XNOR2_X1 U6669 ( .A(n5473), .B(n5482), .ZN(n5799) );
  AOI21_X1 U6670 ( .B1(n6092), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5475) );
  OAI21_X1 U6671 ( .B1(n6086), .B2(n5475), .A(n5474), .ZN(n5476) );
  AOI21_X1 U6672 ( .B1(n5799), .B2(n6470), .A(n5476), .ZN(n5477) );
  OAI21_X1 U6673 ( .B1(n5478), .B2(n6473), .A(n5477), .ZN(U2994) );
  AOI21_X1 U6674 ( .B1(n5481), .B2(n5480), .A(n5479), .ZN(n5497) );
  INV_X1 U6675 ( .A(n5482), .ZN(n5483) );
  NAND2_X1 U6676 ( .A1(n5473), .A2(n5483), .ZN(n5484) );
  AOI21_X1 U6677 ( .B1(n5485), .B2(n5484), .A(n5570), .ZN(n5797) );
  INV_X1 U6678 ( .A(n5486), .ZN(n6082) );
  NOR2_X1 U6679 ( .A1(n6218), .A2(n7040), .ZN(n5492) );
  AOI21_X1 U6680 ( .B1(n6082), .B2(n5488), .A(n5492), .ZN(n5487) );
  OAI21_X1 U6681 ( .B1(n6086), .B2(n5488), .A(n5487), .ZN(n5489) );
  AOI21_X1 U6682 ( .B1(n5797), .B2(n6470), .A(n5489), .ZN(n5490) );
  OAI21_X1 U6683 ( .B1(n5497), .B2(n6473), .A(n5490), .ZN(U2993) );
  OAI21_X1 U6684 ( .B1(n5465), .B2(n5491), .A(n5567), .ZN(n5851) );
  INV_X1 U6685 ( .A(n5851), .ZN(n5495) );
  AOI21_X1 U6686 ( .B1(n6422), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5492), 
        .ZN(n5493) );
  OAI21_X1 U6687 ( .B1(n5577), .B2(n6432), .A(n5493), .ZN(n5494) );
  AOI21_X1 U6688 ( .B1(n5495), .B2(n6065), .A(n5494), .ZN(n5496) );
  OAI21_X1 U6689 ( .B1(n5497), .B2(n6245), .A(n5496), .ZN(U2961) );
  OAI222_X1 U6690 ( .A1(n5832), .A2(n5498), .B1(n5829), .B2(n5500), .C1(n5499), 
        .C2(n6379), .ZN(U2829) );
  INV_X1 U6691 ( .A(n6236), .ZN(n5502) );
  INV_X1 U6692 ( .A(n4717), .ZN(n5501) );
  AOI21_X1 U6693 ( .B1(n5502), .B2(n5501), .A(n5511), .ZN(n5512) );
  INV_X1 U6694 ( .A(n5503), .ZN(n5509) );
  NAND2_X1 U6695 ( .A1(n4717), .A2(n3903), .ZN(n5507) );
  INV_X1 U6696 ( .A(n5504), .ZN(n5505) );
  OAI22_X1 U6697 ( .A1(n6236), .A2(n5507), .B1(n5506), .B2(n5505), .ZN(n5508)
         );
  AOI21_X1 U6698 ( .B1(n5509), .B2(n6707), .A(n5508), .ZN(n5510) );
  OAI22_X1 U6699 ( .A1(n5512), .A2(n3903), .B1(n5511), .B2(n5510), .ZN(U3459)
         );
  NAND3_X1 U6700 ( .A1(n5514), .A2(n5513), .A3(n5889), .ZN(n5517) );
  AOI22_X1 U6701 ( .A1(n5873), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5885), .ZN(n5516) );
  NAND2_X1 U6702 ( .A1(n5517), .A2(n5516), .ZN(U2860) );
  OR2_X1 U6703 ( .A1(n5654), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5520) );
  INV_X1 U6704 ( .A(n5518), .ZN(n5519) );
  MUX2_X1 U6705 ( .A(n5520), .B(n5519), .S(n5529), .Z(U3474) );
  OAI21_X1 U6706 ( .B1(n5522), .B2(n6244), .A(n5521), .ZN(n5523) );
  NAND3_X1 U6707 ( .A1(n5523), .A2(STATE2_REG_2__SCAN_IN), .A3(n6706), .ZN(
        n5524) );
  NAND2_X1 U6708 ( .A1(n5524), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5526) );
  OAI211_X1 U6709 ( .C1(n5528), .C2(n5527), .A(n5526), .B(n5525), .ZN(n5532)
         );
  AOI211_X1 U6710 ( .C1(n6744), .C2(n6706), .A(n5530), .B(n5529), .ZN(n5531)
         );
  MUX2_X1 U6711 ( .A(n5532), .B(REQUESTPENDING_REG_SCAN_IN), .S(n5531), .Z(
        U3472) );
  AND2_X1 U6712 ( .A1(n5534), .A2(n5533), .ZN(n6246) );
  MUX2_X1 U6713 ( .A(MORE_REG_SCAN_IN), .B(n5535), .S(n6246), .Z(U3471) );
  INV_X1 U6714 ( .A(n5792), .ZN(n5543) );
  OAI22_X1 U6715 ( .A1(n6347), .A2(n5537), .B1(n5536), .B2(n5694), .ZN(n5539)
         );
  NOR2_X1 U6716 ( .A1(n6306), .A2(n4314), .ZN(n5538) );
  AOI211_X1 U6717 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5550), .A(n5539), .B(n5538), .ZN(n5540) );
  OAI21_X1 U6718 ( .B1(n5541), .B2(REIP_REG_29__SCAN_IN), .A(n5540), .ZN(n5542) );
  AOI21_X1 U6719 ( .B1(n5543), .B2(n6361), .A(n5542), .ZN(n5544) );
  OAI21_X1 U6720 ( .B1(n5839), .B2(n5780), .A(n5544), .ZN(U2798) );
  AOI21_X1 U6721 ( .B1(n5546), .B2(n4284), .A(n5545), .ZN(n5904) );
  INV_X1 U6722 ( .A(n5904), .ZN(n5842) );
  AOI21_X1 U6723 ( .B1(n5548), .B2(n3091), .A(n5547), .ZN(n6077) );
  INV_X1 U6724 ( .A(n5563), .ZN(n5549) );
  AOI21_X1 U6725 ( .B1(n5549), .B2(REIP_REG_27__SCAN_IN), .A(
        REIP_REG_28__SCAN_IN), .ZN(n5554) );
  INV_X1 U6726 ( .A(n5550), .ZN(n5553) );
  AOI22_X1 U6727 ( .A1(n6364), .A2(n5907), .B1(n6358), .B2(
        PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U6728 ( .A1(n6365), .A2(EBX_REG_28__SCAN_IN), .ZN(n5551) );
  OAI211_X1 U6729 ( .C1(n5554), .C2(n5553), .A(n5552), .B(n5551), .ZN(n5555)
         );
  AOI21_X1 U6730 ( .B1(n6077), .B2(n6361), .A(n5555), .ZN(n5556) );
  OAI21_X1 U6731 ( .B1(n5842), .B2(n5780), .A(n5556), .ZN(U2799) );
  INV_X1 U6732 ( .A(n5794), .ZN(n5565) );
  INV_X1 U6733 ( .A(n5557), .ZN(n5571) );
  OAI22_X1 U6734 ( .A1(n6347), .A2(n5559), .B1(n5558), .B2(n5694), .ZN(n5561)
         );
  INV_X1 U6735 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5795) );
  NOR2_X1 U6736 ( .A1(n6306), .A2(n5795), .ZN(n5560) );
  AOI211_X1 U6737 ( .C1(n5571), .C2(REIP_REG_27__SCAN_IN), .A(n5561), .B(n5560), .ZN(n5562) );
  OAI21_X1 U6738 ( .B1(n5563), .B2(REIP_REG_27__SCAN_IN), .A(n5562), .ZN(n5564) );
  AOI21_X1 U6739 ( .B1(n5565), .B2(n6361), .A(n5564), .ZN(n5566) );
  OAI21_X1 U6740 ( .B1(n5845), .B2(n5780), .A(n5566), .ZN(U2800) );
  AOI21_X1 U6741 ( .B1(n5568), .B2(n5567), .A(n4283), .ZN(n5915) );
  INV_X1 U6742 ( .A(n5915), .ZN(n5848) );
  OAI21_X1 U6743 ( .B1(n5570), .B2(n5569), .A(n3098), .ZN(n5796) );
  INV_X1 U6744 ( .A(n5796), .ZN(n6088) );
  INV_X1 U6745 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6875) );
  OAI21_X1 U6746 ( .B1(n5572), .B2(REIP_REG_26__SCAN_IN), .A(n5571), .ZN(n5574) );
  AOI22_X1 U6747 ( .A1(n6364), .A2(n5912), .B1(n6358), .B2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5573) );
  OAI211_X1 U6748 ( .C1(n6306), .C2(n6875), .A(n5574), .B(n5573), .ZN(n5575)
         );
  AOI21_X1 U6749 ( .B1(n6088), .B2(n6361), .A(n5575), .ZN(n5576) );
  OAI21_X1 U6750 ( .B1(n5848), .B2(n5780), .A(n5576), .ZN(U2801) );
  XNOR2_X1 U6751 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n5583) );
  OAI22_X1 U6752 ( .A1(n6347), .A2(n5578), .B1(n5577), .B2(n5694), .ZN(n5579)
         );
  AOI21_X1 U6753 ( .B1(n6365), .B2(EBX_REG_25__SCAN_IN), .A(n5579), .ZN(n5582)
         );
  INV_X1 U6754 ( .A(n6329), .ZN(n5700) );
  NOR2_X1 U6755 ( .A1(n5700), .A2(n5580), .ZN(n5597) );
  NAND2_X1 U6756 ( .A1(n5597), .A2(REIP_REG_25__SCAN_IN), .ZN(n5581) );
  OAI211_X1 U6757 ( .C1(n5590), .C2(n5583), .A(n5582), .B(n5581), .ZN(n5584)
         );
  AOI21_X1 U6758 ( .B1(n5797), .B2(n6361), .A(n5584), .ZN(n5585) );
  OAI21_X1 U6759 ( .B1(n5851), .B2(n5780), .A(n5585), .ZN(U2802) );
  OAI22_X1 U6760 ( .A1(n6347), .A2(n6973), .B1(n5586), .B2(n5694), .ZN(n5587)
         );
  AOI21_X1 U6761 ( .B1(n6365), .B2(EBX_REG_24__SCAN_IN), .A(n5587), .ZN(n5589)
         );
  NAND2_X1 U6762 ( .A1(n5597), .A2(REIP_REG_24__SCAN_IN), .ZN(n5588) );
  OAI211_X1 U6763 ( .C1(n5590), .C2(REIP_REG_24__SCAN_IN), .A(n5589), .B(n5588), .ZN(n5591) );
  AOI21_X1 U6764 ( .B1(n5799), .B2(n6361), .A(n5591), .ZN(n5592) );
  OAI21_X1 U6765 ( .B1(n5854), .B2(n5780), .A(n5592), .ZN(U2803) );
  NAND2_X1 U6766 ( .A1(n5664), .A2(n5594), .ZN(n5605) );
  AOI21_X1 U6767 ( .B1(n5595), .B2(n5605), .A(n5466), .ZN(n5923) );
  INV_X1 U6768 ( .A(n5923), .ZN(n5857) );
  AOI21_X1 U6769 ( .B1(n5596), .B2(n5611), .A(n5473), .ZN(n6096) );
  INV_X1 U6770 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5802) );
  INV_X1 U6771 ( .A(n5632), .ZN(n5617) );
  NOR3_X1 U6772 ( .A1(n5617), .A2(n6956), .A3(n5939), .ZN(n5598) );
  OAI21_X1 U6773 ( .B1(n5598), .B2(REIP_REG_23__SCAN_IN), .A(n5597), .ZN(n5601) );
  INV_X1 U6774 ( .A(n5921), .ZN(n5599) );
  AOI22_X1 U6775 ( .A1(n6364), .A2(n5599), .B1(n6358), .B2(
        PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5600) );
  OAI211_X1 U6776 ( .C1(n6306), .C2(n5802), .A(n5601), .B(n5600), .ZN(n5602)
         );
  AOI21_X1 U6777 ( .B1(n6096), .B2(n6361), .A(n5602), .ZN(n5603) );
  OAI21_X1 U6778 ( .B1(n5857), .B2(n5780), .A(n5603), .ZN(U2804) );
  NAND2_X1 U6779 ( .A1(n5664), .A2(n5604), .ZN(n5622) );
  INV_X1 U6780 ( .A(n5605), .ZN(n5606) );
  AOI21_X1 U6781 ( .B1(n5607), .B2(n5622), .A(n5606), .ZN(n5932) );
  INV_X1 U6782 ( .A(n5932), .ZN(n5860) );
  NAND2_X1 U6783 ( .A1(n5609), .A2(n5608), .ZN(n5610) );
  AND2_X1 U6784 ( .A1(n5611), .A2(n5610), .ZN(n6103) );
  XNOR2_X1 U6785 ( .A(REIP_REG_22__SCAN_IN), .B(REIP_REG_21__SCAN_IN), .ZN(
        n5616) );
  INV_X1 U6786 ( .A(n5928), .ZN(n5612) );
  OAI22_X1 U6787 ( .A1(n6347), .A2(n5930), .B1(n5612), .B2(n5694), .ZN(n5613)
         );
  AOI21_X1 U6788 ( .B1(n6365), .B2(EBX_REG_22__SCAN_IN), .A(n5613), .ZN(n5615)
         );
  NAND3_X1 U6789 ( .A1(n6329), .A2(REIP_REG_22__SCAN_IN), .A3(n5625), .ZN(
        n5614) );
  OAI211_X1 U6790 ( .C1(n5617), .C2(n5616), .A(n5615), .B(n5614), .ZN(n5618)
         );
  AOI21_X1 U6791 ( .B1(n6103), .B2(n6361), .A(n5618), .ZN(n5619) );
  OAI21_X1 U6792 ( .B1(n5860), .B2(n5780), .A(n5619), .ZN(U2805) );
  NAND2_X1 U6793 ( .A1(n5664), .A2(n5620), .ZN(n5637) );
  INV_X1 U6794 ( .A(n5637), .ZN(n5624) );
  INV_X1 U6795 ( .A(n5621), .ZN(n5623) );
  INV_X1 U6796 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5804) );
  AOI22_X1 U6797 ( .A1(n6364), .A2(n5942), .B1(n6358), .B2(
        PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5627) );
  NAND3_X1 U6798 ( .A1(n6329), .A2(REIP_REG_21__SCAN_IN), .A3(n5625), .ZN(
        n5626) );
  OAI211_X1 U6799 ( .C1(n6306), .C2(n5804), .A(n5627), .B(n5626), .ZN(n5631)
         );
  XNOR2_X1 U6800 ( .A(n5628), .B(n5629), .ZN(n6113) );
  NOR2_X1 U6801 ( .A1(n6113), .A2(n6350), .ZN(n5630) );
  AOI211_X1 U6802 ( .C1(n5632), .C2(n5939), .A(n5631), .B(n5630), .ZN(n5633)
         );
  OAI21_X1 U6803 ( .B1(n5945), .B2(n5780), .A(n5633), .ZN(U2806) );
  MUX2_X1 U6804 ( .A(n5648), .B(n5647), .S(n5634), .Z(n5636) );
  XNOR2_X1 U6805 ( .A(n5636), .B(n5635), .ZN(n6127) );
  AND2_X1 U6806 ( .A1(n5664), .A2(n5652), .ZN(n5650) );
  OAI21_X1 U6807 ( .B1(n5650), .B2(n5638), .A(n5637), .ZN(n5953) );
  INV_X1 U6808 ( .A(n5953), .ZN(n5639) );
  NAND2_X1 U6809 ( .A1(n5639), .A2(n6311), .ZN(n5645) );
  OAI22_X1 U6810 ( .A1(n6347), .A2(n7019), .B1(n5949), .B2(n5694), .ZN(n5643)
         );
  INV_X1 U6811 ( .A(n5657), .ZN(n5640) );
  AOI21_X1 U6812 ( .B1(n5640), .B2(REIP_REG_19__SCAN_IN), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5641) );
  AOI211_X1 U6813 ( .C1(REIP_REG_20__SCAN_IN), .C2(n5656), .A(n5700), .B(n5641), .ZN(n5642) );
  AOI211_X1 U6814 ( .C1(n6365), .C2(EBX_REG_20__SCAN_IN), .A(n5643), .B(n5642), 
        .ZN(n5644) );
  OAI211_X1 U6815 ( .C1(n6127), .C2(n6350), .A(n5645), .B(n5644), .ZN(U2807)
         );
  INV_X1 U6816 ( .A(n5646), .ZN(n5680) );
  XNOR2_X1 U6817 ( .A(n5648), .B(n5647), .ZN(n5663) );
  NOR2_X1 U6818 ( .A1(n5680), .A2(n5663), .ZN(n5662) );
  XOR2_X1 U6819 ( .A(n5649), .B(n5662), .Z(n6135) );
  INV_X1 U6820 ( .A(n5650), .ZN(n5651) );
  OAI21_X1 U6821 ( .B1(n5664), .B2(n5652), .A(n5651), .ZN(n5962) );
  INV_X1 U6822 ( .A(n5962), .ZN(n5653) );
  NAND2_X1 U6823 ( .A1(n5653), .A2(n6311), .ZN(n5661) );
  NAND2_X1 U6824 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5655)
         );
  NAND2_X1 U6825 ( .A1(n6373), .A2(n5654), .ZN(n6312) );
  OAI211_X1 U6826 ( .C1(n5694), .C2(n5958), .A(n5655), .B(n6312), .ZN(n5659)
         );
  AOI211_X1 U6827 ( .C1(n5657), .C2(n5957), .A(n5656), .B(n5700), .ZN(n5658)
         );
  AOI211_X1 U6828 ( .C1(EBX_REG_19__SCAN_IN), .C2(n6365), .A(n5659), .B(n5658), 
        .ZN(n5660) );
  OAI211_X1 U6829 ( .C1(n6135), .C2(n6350), .A(n5661), .B(n5660), .ZN(U2808)
         );
  AOI21_X1 U6830 ( .B1(n5663), .B2(n5680), .A(n5662), .ZN(n6140) );
  INV_X1 U6831 ( .A(n6140), .ZN(n5807) );
  AOI21_X1 U6832 ( .B1(n5665), .B2(n5593), .A(n5664), .ZN(n5970) );
  NAND2_X1 U6833 ( .A1(n5970), .A2(n6311), .ZN(n5675) );
  AND2_X1 U6834 ( .A1(n6329), .A2(n5666), .ZN(n5683) );
  INV_X1 U6835 ( .A(n5967), .ZN(n5668) );
  NAND2_X1 U6836 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5667)
         );
  OAI211_X1 U6837 ( .C1(n5694), .C2(n5668), .A(n5667), .B(n6312), .ZN(n5673)
         );
  INV_X1 U6838 ( .A(EBX_REG_18__SCAN_IN), .ZN(n7042) );
  NAND3_X1 U6839 ( .A1(n6359), .A2(n5670), .A3(n5669), .ZN(n5671) );
  OAI21_X1 U6840 ( .B1(n6306), .B2(n7042), .A(n5671), .ZN(n5672) );
  AOI211_X1 U6841 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5683), .A(n5673), .B(n5672), .ZN(n5674) );
  OAI211_X1 U6842 ( .C1(n5807), .C2(n6350), .A(n5675), .B(n5674), .ZN(U2809)
         );
  INV_X1 U6843 ( .A(n5593), .ZN(n5677) );
  AOI21_X1 U6844 ( .B1(n5678), .B2(n5676), .A(n5677), .ZN(n5978) );
  INV_X1 U6845 ( .A(n5978), .ZN(n5872) );
  AOI21_X1 U6846 ( .B1(n5681), .B2(n5679), .A(n5646), .ZN(n6148) );
  INV_X1 U6847 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5687) );
  NOR2_X1 U6848 ( .A1(n6347), .A2(n5976), .ZN(n5682) );
  AOI211_X1 U6849 ( .C1(n6364), .C2(n5974), .A(n6333), .B(n5682), .ZN(n5686)
         );
  NOR3_X1 U6850 ( .A1(n6321), .A2(n5984), .A3(n5697), .ZN(n5684) );
  OAI21_X1 U6851 ( .B1(n5684), .B2(REIP_REG_17__SCAN_IN), .A(n5683), .ZN(n5685) );
  OAI211_X1 U6852 ( .C1(n5687), .C2(n6306), .A(n5686), .B(n5685), .ZN(n5688)
         );
  AOI21_X1 U6853 ( .B1(n6148), .B2(n6361), .A(n5688), .ZN(n5689) );
  OAI21_X1 U6854 ( .B1(n5872), .B2(n5780), .A(n5689), .ZN(U2810) );
  OR2_X1 U6855 ( .A1(n5690), .A2(n5691), .ZN(n5692) );
  AND2_X1 U6856 ( .A1(n5676), .A2(n5692), .ZN(n5988) );
  OAI21_X1 U6857 ( .B1(n3118), .B2(n5693), .A(n5679), .ZN(n6151) );
  INV_X1 U6858 ( .A(n5987), .ZN(n5696) );
  NAND2_X1 U6859 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5695)
         );
  OAI211_X1 U6860 ( .C1(n5694), .C2(n5696), .A(n5695), .B(n6312), .ZN(n5699)
         );
  NOR3_X1 U6861 ( .A1(n6321), .A2(REIP_REG_16__SCAN_IN), .A3(n5697), .ZN(n5698) );
  AOI21_X1 U6862 ( .B1(n5701), .B2(n6373), .A(n5700), .ZN(n5729) );
  INV_X1 U6863 ( .A(n5701), .ZN(n5723) );
  NOR2_X1 U6864 ( .A1(n5723), .A2(REIP_REG_15__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6865 ( .A1(n6359), .A2(n5702), .ZN(n5714) );
  INV_X1 U6866 ( .A(n5714), .ZN(n5703) );
  OAI21_X1 U6867 ( .B1(n5729), .B2(n5703), .A(REIP_REG_16__SCAN_IN), .ZN(n5704) );
  AND2_X1 U6868 ( .A1(n5732), .A2(n5705), .ZN(n5706) );
  OR2_X1 U6869 ( .A1(n5706), .A2(n3118), .ZN(n6169) );
  INV_X1 U6870 ( .A(n5708), .ZN(n5709) );
  XNOR2_X1 U6871 ( .A(n5707), .B(n5709), .ZN(n5813) );
  INV_X1 U6872 ( .A(n5812), .ZN(n5710) );
  OAI22_X1 U6873 ( .A1(n5813), .A2(n5710), .B1(n5709), .B2(n5707), .ZN(n5721)
         );
  NAND2_X1 U6874 ( .A1(n5721), .A2(n5720), .ZN(n5719) );
  INV_X1 U6875 ( .A(n5711), .ZN(n5712) );
  AOI21_X1 U6876 ( .B1(n5719), .B2(n5712), .A(n5690), .ZN(n5999) );
  NAND2_X1 U6877 ( .A1(n5999), .A2(n6311), .ZN(n5718) );
  NAND2_X1 U6878 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5713)
         );
  OAI211_X1 U6879 ( .C1(n5694), .C2(n5997), .A(n5713), .B(n6312), .ZN(n5716)
         );
  INV_X1 U6880 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5810) );
  OAI21_X1 U6881 ( .B1(n6306), .B2(n5810), .A(n5714), .ZN(n5715) );
  AOI211_X1 U6882 ( .C1(n5729), .C2(REIP_REG_15__SCAN_IN), .A(n5716), .B(n5715), .ZN(n5717) );
  OAI211_X1 U6883 ( .C1(n6169), .C2(n6350), .A(n5718), .B(n5717), .ZN(U2812)
         );
  OAI21_X1 U6884 ( .B1(n5721), .B2(n5720), .A(n5719), .ZN(n6003) );
  NAND2_X1 U6885 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5722)
         );
  OAI211_X1 U6886 ( .C1(n5694), .C2(n6004), .A(n5722), .B(n6312), .ZN(n5728)
         );
  INV_X1 U6887 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5726) );
  NAND3_X1 U6888 ( .A1(n6359), .A2(n5724), .A3(n5723), .ZN(n5725) );
  OAI21_X1 U6889 ( .B1(n6306), .B2(n5726), .A(n5725), .ZN(n5727) );
  AOI211_X1 U6890 ( .C1(n5729), .C2(REIP_REG_14__SCAN_IN), .A(n5728), .B(n5727), .ZN(n5734) );
  NAND2_X1 U6891 ( .A1(n5825), .A2(n5814), .ZN(n5816) );
  NAND2_X1 U6892 ( .A1(n5816), .A2(n5730), .ZN(n5731) );
  AND2_X1 U6893 ( .A1(n5732), .A2(n5731), .ZN(n6178) );
  NAND2_X1 U6894 ( .A1(n6178), .A2(n6361), .ZN(n5733) );
  OAI211_X1 U6895 ( .C1(n6003), .C2(n5780), .A(n5734), .B(n5733), .ZN(U2813)
         );
  OAI21_X1 U6896 ( .B1(n5735), .B2(n5737), .A(n5820), .ZN(n6031) );
  INV_X1 U6897 ( .A(n6266), .ZN(n5738) );
  OAI21_X1 U6898 ( .B1(n6321), .B2(n5738), .A(n6373), .ZN(n6276) );
  NAND3_X1 U6899 ( .A1(n6359), .A2(n6266), .A3(n5739), .ZN(n5740) );
  OAI211_X1 U6900 ( .C1(n5694), .C2(n6033), .A(n5740), .B(n6312), .ZN(n5745)
         );
  INV_X1 U6901 ( .A(n5741), .ZN(n5751) );
  AOI21_X1 U6902 ( .B1(n5742), .B2(n5751), .A(n5823), .ZN(n6210) );
  AOI22_X1 U6903 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6365), .B1(n6361), .B2(n6210), .ZN(n5743) );
  OAI21_X1 U6904 ( .B1(n6935), .B2(n6347), .A(n5743), .ZN(n5744) );
  AOI211_X1 U6905 ( .C1(REIP_REG_11__SCAN_IN), .C2(n6276), .A(n5745), .B(n5744), .ZN(n5746) );
  OAI21_X1 U6906 ( .B1(n5780), .B2(n6031), .A(n5746), .ZN(U2816) );
  AOI21_X1 U6907 ( .B1(n3988), .B2(n3082), .A(n5735), .ZN(n6046) );
  INV_X1 U6908 ( .A(n6046), .ZN(n5888) );
  NAND2_X1 U6909 ( .A1(n5748), .A2(n5749), .ZN(n5750) );
  NAND2_X1 U6910 ( .A1(n5751), .A2(n5750), .ZN(n6220) );
  AOI22_X1 U6911 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6365), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6358), .ZN(n5752) );
  OAI211_X1 U6912 ( .C1(n6350), .C2(n6220), .A(n5752), .B(n6312), .ZN(n5758)
         );
  INV_X1 U6913 ( .A(n6373), .ZN(n6330) );
  OAI21_X1 U6914 ( .B1(n6330), .B2(n5753), .A(n6329), .ZN(n6294) );
  AND2_X1 U6915 ( .A1(n6359), .A2(n5754), .ZN(n6285) );
  NAND2_X1 U6916 ( .A1(n6285), .A2(REIP_REG_8__SCAN_IN), .ZN(n5761) );
  OAI21_X1 U6917 ( .B1(REIP_REG_9__SCAN_IN), .B2(REIP_REG_10__SCAN_IN), .A(
        n5755), .ZN(n5756) );
  OAI22_X1 U6918 ( .A1(n6294), .A2(n6219), .B1(n5761), .B2(n5756), .ZN(n5757)
         );
  AOI211_X1 U6919 ( .C1(n6042), .C2(n6364), .A(n5758), .B(n5757), .ZN(n5759)
         );
  OAI21_X1 U6920 ( .B1(n5780), .B2(n5888), .A(n5759), .ZN(U2817) );
  OAI21_X1 U6921 ( .B1(n5353), .B2(n5760), .A(n3082), .ZN(n6054) );
  INV_X1 U6922 ( .A(n6050), .ZN(n5770) );
  INV_X1 U6923 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U6924 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6294), .B1(n5761), .B2(n6838), .ZN(n5769) );
  INV_X1 U6925 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5767) );
  INV_X1 U6926 ( .A(n5762), .ZN(n5765) );
  INV_X1 U6927 ( .A(n5748), .ZN(n5763) );
  AOI21_X1 U6928 ( .B1(n5765), .B2(n5764), .A(n5763), .ZN(n6435) );
  AOI22_X1 U6929 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6365), .B1(n6361), .B2(n6435), 
        .ZN(n5766) );
  OAI211_X1 U6930 ( .C1(n6347), .C2(n5767), .A(n5766), .B(n6312), .ZN(n5768)
         );
  AOI211_X1 U6931 ( .C1(n6364), .C2(n5770), .A(n5769), .B(n5768), .ZN(n5771)
         );
  OAI21_X1 U6932 ( .B1(n5780), .B2(n6054), .A(n5771), .ZN(U2818) );
  AOI21_X1 U6933 ( .B1(n6359), .B2(n6996), .A(n6330), .ZN(n6345) );
  NAND3_X1 U6934 ( .A1(n6359), .A2(REIP_REG_1__SCAN_IN), .A3(n6989), .ZN(n5773) );
  NAND2_X1 U6935 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5772)
         );
  OAI211_X1 U6936 ( .C1(n6431), .C2(n5694), .A(n5773), .B(n5772), .ZN(n5777)
         );
  INV_X1 U6937 ( .A(n4714), .ZN(n6232) );
  AND2_X1 U6938 ( .A1(n5779), .A2(n5774), .ZN(n6362) );
  INV_X1 U6939 ( .A(n6362), .ZN(n6348) );
  OAI22_X1 U6940 ( .A1(n6232), .A2(n6348), .B1(n6306), .B2(n5775), .ZN(n5776)
         );
  AOI211_X1 U6941 ( .C1(n6361), .C2(n6453), .A(n5777), .B(n5776), .ZN(n5783)
         );
  NAND2_X1 U6942 ( .A1(n5779), .A2(n5778), .ZN(n5781) );
  NAND2_X1 U6943 ( .A1(n5781), .A2(n5780), .ZN(n6324) );
  NAND2_X1 U6944 ( .A1(n6427), .A2(n6324), .ZN(n5782) );
  OAI211_X1 U6945 ( .C1(n6345), .C2(n6989), .A(n5783), .B(n5782), .ZN(U2825)
         );
  OAI22_X1 U6946 ( .A1(n5784), .A2(n6348), .B1(n6350), .B2(n6468), .ZN(n5785)
         );
  AOI21_X1 U6947 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6329), .A(n5785), .ZN(n5788)
         );
  NAND2_X1 U6948 ( .A1(n6347), .A2(n5694), .ZN(n5786) );
  AOI22_X1 U6949 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5786), .B1(n6365), 
        .B2(EBX_REG_0__SCAN_IN), .ZN(n5787) );
  OAI211_X1 U6950 ( .C1(n6369), .C2(n6064), .A(n5788), .B(n5787), .ZN(U2827)
         );
  INV_X1 U6951 ( .A(n5789), .ZN(n5791) );
  OAI22_X1 U6952 ( .A1(n5791), .A2(n5829), .B1(n5790), .B2(n6379), .ZN(U2828)
         );
  OAI222_X1 U6953 ( .A1(n4314), .A2(n6379), .B1(n5829), .B2(n5792), .C1(n5839), 
        .C2(n5832), .ZN(U2830) );
  AOI22_X1 U6954 ( .A1(n6077), .A2(n6375), .B1(n5830), .B2(EBX_REG_28__SCAN_IN), .ZN(n5793) );
  OAI21_X1 U6955 ( .B1(n5842), .B2(n5832), .A(n5793), .ZN(U2831) );
  OAI222_X1 U6956 ( .A1(n5795), .A2(n6379), .B1(n5829), .B2(n5794), .C1(n5845), 
        .C2(n5832), .ZN(U2832) );
  OAI222_X1 U6957 ( .A1(n5796), .A2(n5829), .B1(n6875), .B2(n6379), .C1(n5848), 
        .C2(n5832), .ZN(U2833) );
  AOI22_X1 U6958 ( .A1(n5797), .A2(n6375), .B1(n5830), .B2(EBX_REG_25__SCAN_IN), .ZN(n5798) );
  OAI21_X1 U6959 ( .B1(n5851), .B2(n5832), .A(n5798), .ZN(U2834) );
  AOI22_X1 U6960 ( .A1(n5799), .A2(n6375), .B1(EBX_REG_24__SCAN_IN), .B2(n5830), .ZN(n5800) );
  OAI21_X1 U6961 ( .B1(n5854), .B2(n5832), .A(n5800), .ZN(U2835) );
  INV_X1 U6962 ( .A(n6096), .ZN(n5801) );
  OAI222_X1 U6963 ( .A1(n5802), .A2(n6379), .B1(n5829), .B2(n5801), .C1(n5857), 
        .C2(n5832), .ZN(U2836) );
  AOI22_X1 U6964 ( .A1(n6103), .A2(n6375), .B1(n5830), .B2(EBX_REG_22__SCAN_IN), .ZN(n5803) );
  OAI21_X1 U6965 ( .B1(n5860), .B2(n5832), .A(n5803), .ZN(U2837) );
  OAI222_X1 U6966 ( .A1(n6113), .A2(n5829), .B1(n5804), .B2(n6379), .C1(n5945), 
        .C2(n5832), .ZN(U2838) );
  OAI222_X1 U6967 ( .A1(n5953), .A2(n5832), .B1(n5829), .B2(n6127), .C1(n5805), 
        .C2(n6379), .ZN(U2839) );
  INV_X1 U6968 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5806) );
  OAI222_X1 U6969 ( .A1(n5962), .A2(n5832), .B1(n5829), .B2(n6135), .C1(n6379), 
        .C2(n5806), .ZN(U2840) );
  INV_X1 U6970 ( .A(n5970), .ZN(n5869) );
  OAI222_X1 U6971 ( .A1(n5869), .A2(n5832), .B1(n6379), .B2(n7042), .C1(n5807), 
        .C2(n5829), .ZN(U2841) );
  AOI22_X1 U6972 ( .A1(n6148), .A2(n6375), .B1(n5830), .B2(EBX_REG_17__SCAN_IN), .ZN(n5808) );
  OAI21_X1 U6973 ( .B1(n5872), .B2(n5832), .A(n5808), .ZN(U2842) );
  INV_X1 U6974 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5809) );
  INV_X1 U6975 ( .A(n5988), .ZN(n5877) );
  OAI222_X1 U6976 ( .A1(n6151), .A2(n5829), .B1(n5809), .B2(n6379), .C1(n5877), 
        .C2(n5832), .ZN(U2843) );
  INV_X1 U6977 ( .A(n5999), .ZN(n5879) );
  OAI222_X1 U6978 ( .A1(n6169), .A2(n5829), .B1(n5810), .B2(n6379), .C1(n5879), 
        .C2(n5832), .ZN(U2844) );
  INV_X1 U6979 ( .A(n6178), .ZN(n5811) );
  OAI222_X1 U6980 ( .A1(n5811), .A2(n5829), .B1(n6379), .B2(n5726), .C1(n5832), 
        .C2(n6003), .ZN(U2845) );
  XNOR2_X1 U6981 ( .A(n5813), .B(n5812), .ZN(n6265) );
  OR2_X1 U6982 ( .A1(n5825), .A2(n5814), .ZN(n5815) );
  NAND2_X1 U6983 ( .A1(n5816), .A2(n5815), .ZN(n6260) );
  OAI22_X1 U6984 ( .A1(n6260), .A2(n5829), .B1(n6261), .B2(n6379), .ZN(n5817)
         );
  INV_X1 U6985 ( .A(n5817), .ZN(n5818) );
  OAI21_X1 U6986 ( .B1(n6016), .B2(n5832), .A(n5818), .ZN(U2846) );
  NAND2_X1 U6987 ( .A1(n5820), .A2(n5819), .ZN(n5821) );
  AND2_X1 U6988 ( .A1(n5707), .A2(n5821), .ZN(n6279) );
  INV_X1 U6989 ( .A(n6279), .ZN(n5883) );
  INV_X1 U6990 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5826) );
  NOR2_X1 U6991 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  OR2_X1 U6992 ( .A1(n5825), .A2(n5824), .ZN(n6274) );
  OAI222_X1 U6993 ( .A1(n5883), .A2(n5832), .B1(n6379), .B2(n5826), .C1(n5829), 
        .C2(n6274), .ZN(U2847) );
  AOI22_X1 U6994 ( .A1(n6210), .A2(n6375), .B1(n5830), .B2(EBX_REG_11__SCAN_IN), .ZN(n5827) );
  OAI21_X1 U6995 ( .B1(n6031), .B2(n5832), .A(n5827), .ZN(U2848) );
  INV_X1 U6996 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5828) );
  OAI222_X1 U6997 ( .A1(n6220), .A2(n5829), .B1(n6379), .B2(n5828), .C1(n5832), 
        .C2(n5888), .ZN(U2849) );
  AOI22_X1 U6998 ( .A1(n6435), .A2(n6375), .B1(EBX_REG_9__SCAN_IN), .B2(n5830), 
        .ZN(n5831) );
  OAI21_X1 U6999 ( .B1(n6054), .B2(n5832), .A(n5831), .ZN(U2850) );
  AOI22_X1 U7000 ( .A1(n5873), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5885), .ZN(n5836) );
  AND2_X1 U7001 ( .A1(n5833), .A2(n3392), .ZN(n5834) );
  NAND2_X1 U7002 ( .A1(n5874), .A2(DATAI_14_), .ZN(n5835) );
  OAI211_X1 U7003 ( .C1(n5498), .C2(n5892), .A(n5836), .B(n5835), .ZN(U2861)
         );
  AOI22_X1 U7004 ( .A1(n5873), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5885), .ZN(n5838) );
  NAND2_X1 U7005 ( .A1(n5874), .A2(DATAI_13_), .ZN(n5837) );
  OAI211_X1 U7006 ( .C1(n5839), .C2(n5892), .A(n5838), .B(n5837), .ZN(U2862)
         );
  AOI22_X1 U7007 ( .A1(n5873), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5885), .ZN(n5841) );
  NAND2_X1 U7008 ( .A1(n5874), .A2(DATAI_12_), .ZN(n5840) );
  OAI211_X1 U7009 ( .C1(n5842), .C2(n5892), .A(n5841), .B(n5840), .ZN(U2863)
         );
  AOI22_X1 U7010 ( .A1(n5873), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5885), .ZN(n5844) );
  NAND2_X1 U7011 ( .A1(n5874), .A2(DATAI_11_), .ZN(n5843) );
  OAI211_X1 U7012 ( .C1(n5845), .C2(n5892), .A(n5844), .B(n5843), .ZN(U2864)
         );
  AOI22_X1 U7013 ( .A1(n5873), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5885), .ZN(n5847) );
  NAND2_X1 U7014 ( .A1(n5874), .A2(DATAI_10_), .ZN(n5846) );
  OAI211_X1 U7015 ( .C1(n5848), .C2(n5892), .A(n5847), .B(n5846), .ZN(U2865)
         );
  AOI22_X1 U7016 ( .A1(n5873), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5885), .ZN(n5850) );
  NAND2_X1 U7017 ( .A1(n5874), .A2(DATAI_9_), .ZN(n5849) );
  OAI211_X1 U7018 ( .C1(n5851), .C2(n5892), .A(n5850), .B(n5849), .ZN(U2866)
         );
  AOI22_X1 U7019 ( .A1(n5873), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5885), .ZN(n5853) );
  NAND2_X1 U7020 ( .A1(n5874), .A2(DATAI_8_), .ZN(n5852) );
  OAI211_X1 U7021 ( .C1(n5854), .C2(n5892), .A(n5853), .B(n5852), .ZN(U2867)
         );
  AOI22_X1 U7022 ( .A1(n5873), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n5885), .ZN(n5856) );
  NAND2_X1 U7023 ( .A1(n5874), .A2(DATAI_7_), .ZN(n5855) );
  OAI211_X1 U7024 ( .C1(n5857), .C2(n5892), .A(n5856), .B(n5855), .ZN(U2868)
         );
  AOI22_X1 U7025 ( .A1(n5873), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n5885), .ZN(n5859) );
  NAND2_X1 U7026 ( .A1(n5874), .A2(DATAI_6_), .ZN(n5858) );
  OAI211_X1 U7027 ( .C1(n5860), .C2(n5892), .A(n5859), .B(n5858), .ZN(U2869)
         );
  AOI22_X1 U7028 ( .A1(n5873), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n5885), .ZN(n5862) );
  NAND2_X1 U7029 ( .A1(n5874), .A2(DATAI_5_), .ZN(n5861) );
  OAI211_X1 U7030 ( .C1(n5945), .C2(n5892), .A(n5862), .B(n5861), .ZN(U2870)
         );
  AOI22_X1 U7031 ( .A1(n5873), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n5885), .ZN(n5864) );
  NAND2_X1 U7032 ( .A1(n5874), .A2(DATAI_4_), .ZN(n5863) );
  OAI211_X1 U7033 ( .C1(n5953), .C2(n5892), .A(n5864), .B(n5863), .ZN(U2871)
         );
  AOI22_X1 U7034 ( .A1(n5873), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n5885), .ZN(n5866) );
  NAND2_X1 U7035 ( .A1(n5874), .A2(DATAI_3_), .ZN(n5865) );
  OAI211_X1 U7036 ( .C1(n5962), .C2(n5892), .A(n5866), .B(n5865), .ZN(U2872)
         );
  AOI22_X1 U7037 ( .A1(n5873), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n5885), .ZN(n5868) );
  NAND2_X1 U7038 ( .A1(n5874), .A2(DATAI_2_), .ZN(n5867) );
  OAI211_X1 U7039 ( .C1(n5869), .C2(n5892), .A(n5868), .B(n5867), .ZN(U2873)
         );
  AOI22_X1 U7040 ( .A1(n5873), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5885), .ZN(n5871) );
  NAND2_X1 U7041 ( .A1(n5874), .A2(DATAI_1_), .ZN(n5870) );
  OAI211_X1 U7042 ( .C1(n5872), .C2(n5892), .A(n5871), .B(n5870), .ZN(U2874)
         );
  AOI22_X1 U7043 ( .A1(n5873), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n5885), .ZN(n5876) );
  NAND2_X1 U7044 ( .A1(n5874), .A2(DATAI_0_), .ZN(n5875) );
  OAI211_X1 U7045 ( .C1(n5877), .C2(n5892), .A(n5876), .B(n5875), .ZN(U2875)
         );
  INV_X1 U7046 ( .A(DATAI_15_), .ZN(n5878) );
  OAI222_X1 U7047 ( .A1(n5879), .A2(n5892), .B1(n5889), .B2(n6997), .C1(n5891), 
        .C2(n5878), .ZN(U2876) );
  INV_X1 U7048 ( .A(DATAI_14_), .ZN(n5880) );
  OAI222_X1 U7049 ( .A1(n6003), .A2(n5892), .B1(n5889), .B2(n5881), .C1(n5880), 
        .C2(n5891), .ZN(U2877) );
  INV_X1 U7050 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6387) );
  INV_X1 U7051 ( .A(DATAI_13_), .ZN(n6868) );
  OAI222_X1 U7052 ( .A1(n5889), .A2(n6387), .B1(n5891), .B2(n6868), .C1(n5892), 
        .C2(n6016), .ZN(U2878) );
  AOI22_X1 U7053 ( .A1(n5886), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n5885), .ZN(n5882) );
  OAI21_X1 U7054 ( .B1(n5883), .B2(n5892), .A(n5882), .ZN(U2879) );
  AOI22_X1 U7055 ( .A1(n5886), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5885), .ZN(n5884) );
  OAI21_X1 U7056 ( .B1(n6031), .B2(n5892), .A(n5884), .ZN(U2880) );
  AOI22_X1 U7057 ( .A1(n5886), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5885), .ZN(n5887) );
  OAI21_X1 U7058 ( .B1(n5888), .B2(n5892), .A(n5887), .ZN(U2881) );
  INV_X1 U7059 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6965) );
  OAI222_X1 U7060 ( .A1(n6054), .A2(n5892), .B1(n5891), .B2(n5890), .C1(n5889), 
        .C2(n6965), .ZN(U2882) );
  AOI21_X1 U7061 ( .B1(n6422), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5893), 
        .ZN(n5894) );
  OAI21_X1 U7062 ( .B1(n5895), .B2(n6432), .A(n5894), .ZN(n5896) );
  AOI21_X1 U7063 ( .B1(n5897), .B2(n6428), .A(n5896), .ZN(n5898) );
  OAI21_X1 U7064 ( .B1(n5498), .B2(n6057), .A(n5898), .ZN(U2956) );
  AOI22_X1 U7065 ( .A1(n5901), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .B1(n5900), .B2(n5899), .ZN(n5903) );
  XNOR2_X1 U7066 ( .A(n5903), .B(n5902), .ZN(n6079) );
  NAND2_X1 U7067 ( .A1(n5904), .A2(n6065), .ZN(n5909) );
  NAND2_X1 U7068 ( .A1(n6457), .A2(REIP_REG_28__SCAN_IN), .ZN(n6072) );
  OAI21_X1 U7069 ( .B1(n6056), .B2(n5905), .A(n6072), .ZN(n5906) );
  AOI21_X1 U7070 ( .B1(n6060), .B2(n5907), .A(n5906), .ZN(n5908) );
  OAI211_X1 U7071 ( .C1(n6079), .C2(n6245), .A(n5909), .B(n5908), .ZN(U2958)
         );
  XNOR2_X1 U7072 ( .A(n4300), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5910)
         );
  XNOR2_X1 U7073 ( .A(n5911), .B(n5910), .ZN(n6090) );
  NAND2_X1 U7074 ( .A1(n6060), .A2(n5912), .ZN(n5913) );
  NAND2_X1 U7075 ( .A1(n6457), .A2(REIP_REG_26__SCAN_IN), .ZN(n6084) );
  OAI211_X1 U7076 ( .C1(n6056), .C2(n6849), .A(n5913), .B(n6084), .ZN(n5914)
         );
  AOI21_X1 U7077 ( .B1(n5915), .B2(n6065), .A(n5914), .ZN(n5916) );
  OAI21_X1 U7078 ( .B1(n6245), .B2(n6090), .A(n5916), .ZN(U2960) );
  INV_X1 U7079 ( .A(n5917), .ZN(n5955) );
  XNOR2_X1 U7080 ( .A(n5919), .B(n6094), .ZN(n6098) );
  NOR2_X1 U7081 ( .A1(n6218), .A2(n6958), .ZN(n6091) );
  AOI21_X1 U7082 ( .B1(n6422), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6091), 
        .ZN(n5920) );
  OAI21_X1 U7083 ( .B1(n5921), .B2(n6432), .A(n5920), .ZN(n5922) );
  AOI21_X1 U7084 ( .B1(n5923), .B2(n6065), .A(n5922), .ZN(n5924) );
  OAI21_X1 U7085 ( .B1(n6098), .B2(n6245), .A(n5924), .ZN(U2963) );
  OAI21_X1 U7086 ( .B1(n3080), .B2(n6855), .A(n5925), .ZN(n5927) );
  XOR2_X1 U7087 ( .A(n5927), .B(n5926), .Z(n6105) );
  NAND2_X1 U7088 ( .A1(n6060), .A2(n5928), .ZN(n5929) );
  NAND2_X1 U7089 ( .A1(n6457), .A2(REIP_REG_22__SCAN_IN), .ZN(n6101) );
  OAI211_X1 U7090 ( .C1(n6056), .C2(n5930), .A(n5929), .B(n6101), .ZN(n5931)
         );
  AOI21_X1 U7091 ( .B1(n5932), .B2(n6065), .A(n5931), .ZN(n5933) );
  OAI21_X1 U7092 ( .B1(n6105), .B2(n6245), .A(n5933), .ZN(U2964) );
  OR2_X1 U7093 ( .A1(n5947), .A2(n5946), .ZN(n5935) );
  NAND2_X1 U7094 ( .A1(n5935), .A2(n5934), .ZN(n5938) );
  OAI21_X1 U7095 ( .B1(n5938), .B2(n5937), .A(n5936), .ZN(n6106) );
  NAND2_X1 U7096 ( .A1(n6106), .A2(n6428), .ZN(n5944) );
  NOR2_X1 U7097 ( .A1(n6218), .A2(n5939), .ZN(n6109) );
  NOR2_X1 U7098 ( .A1(n6056), .A2(n5940), .ZN(n5941) );
  AOI211_X1 U7099 ( .C1(n6060), .C2(n5942), .A(n6109), .B(n5941), .ZN(n5943)
         );
  OAI211_X1 U7100 ( .C1(n6057), .C2(n5945), .A(n5944), .B(n5943), .ZN(U2965)
         );
  XNOR2_X1 U7101 ( .A(n5947), .B(n5946), .ZN(n6114) );
  NAND2_X1 U7102 ( .A1(n6114), .A2(n6428), .ZN(n5952) );
  NOR2_X1 U7103 ( .A1(n6218), .A2(n5948), .ZN(n6124) );
  NOR2_X1 U7104 ( .A1(n6432), .A2(n5949), .ZN(n5950) );
  AOI211_X1 U7105 ( .C1(n6422), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n6124), 
        .B(n5950), .ZN(n5951) );
  OAI211_X1 U7106 ( .C1(n6057), .C2(n5953), .A(n5952), .B(n5951), .ZN(U2966)
         );
  AOI21_X1 U7107 ( .B1(n5954), .B2(n5956), .A(n5955), .ZN(n6128) );
  NAND2_X1 U7108 ( .A1(n6128), .A2(n6428), .ZN(n5961) );
  NOR2_X1 U7109 ( .A1(n6218), .A2(n5957), .ZN(n6131) );
  NOR2_X1 U7110 ( .A1(n6432), .A2(n5958), .ZN(n5959) );
  AOI211_X1 U7111 ( .C1(n6422), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6131), 
        .B(n5959), .ZN(n5960) );
  OAI211_X1 U7112 ( .C1(n6057), .C2(n5962), .A(n5961), .B(n5960), .ZN(U2967)
         );
  OAI21_X1 U7113 ( .B1(n3080), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5963), 
        .ZN(n5995) );
  NOR2_X1 U7114 ( .A1(n3080), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5991)
         );
  OAI21_X2 U7115 ( .B1(n5995), .B2(n5991), .A(n5992), .ZN(n5982) );
  NOR2_X1 U7116 ( .A1(n4300), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5980)
         );
  NAND2_X1 U7117 ( .A1(n5980), .A2(n6959), .ZN(n5965) );
  NAND4_X1 U7118 ( .A1(n5982), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A4(n4300), .ZN(n5964) );
  OAI21_X1 U7119 ( .B1(n5982), .B2(n5965), .A(n5964), .ZN(n5966) );
  XNOR2_X1 U7120 ( .A(n5966), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6142)
         );
  NAND2_X1 U7121 ( .A1(n6060), .A2(n5967), .ZN(n5968) );
  NAND2_X1 U7122 ( .A1(n6457), .A2(REIP_REG_18__SCAN_IN), .ZN(n6137) );
  OAI211_X1 U7123 ( .C1(n6056), .C2(n3213), .A(n5968), .B(n6137), .ZN(n5969)
         );
  AOI21_X1 U7124 ( .B1(n5970), .B2(n6065), .A(n5969), .ZN(n5971) );
  OAI21_X1 U7125 ( .B1(n6142), .B2(n6245), .A(n5971), .ZN(U2968) );
  NOR2_X1 U7126 ( .A1(n3080), .A2(n5972), .ZN(n5981) );
  MUX2_X1 U7127 ( .A(n5980), .B(n5981), .S(n5982), .Z(n5973) );
  XNOR2_X1 U7128 ( .A(n5973), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6150)
         );
  NAND2_X1 U7129 ( .A1(n6060), .A2(n5974), .ZN(n5975) );
  NAND2_X1 U7130 ( .A1(n6457), .A2(REIP_REG_17__SCAN_IN), .ZN(n6145) );
  OAI211_X1 U7131 ( .C1(n6056), .C2(n5976), .A(n5975), .B(n6145), .ZN(n5977)
         );
  AOI21_X1 U7132 ( .B1(n5978), .B2(n6065), .A(n5977), .ZN(n5979) );
  OAI21_X1 U7133 ( .B1(n6150), .B2(n6245), .A(n5979), .ZN(U2969) );
  NOR2_X1 U7134 ( .A1(n5981), .A2(n5980), .ZN(n5983) );
  XOR2_X1 U7135 ( .A(n5983), .B(n5982), .Z(n6165) );
  NOR2_X1 U7136 ( .A1(n6218), .A2(n5984), .ZN(n6155) );
  INV_X1 U7137 ( .A(n6155), .ZN(n5985) );
  OAI21_X1 U7138 ( .B1(n6056), .B2(n3211), .A(n5985), .ZN(n5986) );
  AOI21_X1 U7139 ( .B1(n6060), .B2(n5987), .A(n5986), .ZN(n5990) );
  NAND2_X1 U7140 ( .A1(n5988), .A2(n6065), .ZN(n5989) );
  OAI211_X1 U7141 ( .C1(n6165), .C2(n6245), .A(n5990), .B(n5989), .ZN(U2970)
         );
  INV_X1 U7142 ( .A(n5991), .ZN(n5993) );
  NAND2_X1 U7143 ( .A1(n5993), .A2(n5992), .ZN(n5994) );
  XNOR2_X1 U7144 ( .A(n5995), .B(n5994), .ZN(n6173) );
  NAND2_X1 U7145 ( .A1(n6457), .A2(REIP_REG_15__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7146 ( .A1(n6422), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5996)
         );
  OAI211_X1 U7147 ( .C1(n6432), .C2(n5997), .A(n6168), .B(n5996), .ZN(n5998)
         );
  AOI21_X1 U7148 ( .B1(n5999), .B2(n6065), .A(n5998), .ZN(n6000) );
  OAI21_X1 U7149 ( .B1(n6173), .B2(n6245), .A(n6000), .ZN(U2971) );
  XNOR2_X1 U7150 ( .A(n3080), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6002)
         );
  XNOR2_X1 U7151 ( .A(n6001), .B(n6002), .ZN(n6185) );
  INV_X1 U7152 ( .A(n6003), .ZN(n6008) );
  NOR2_X1 U7153 ( .A1(n6432), .A2(n6004), .ZN(n6007) );
  NAND2_X1 U7154 ( .A1(n6457), .A2(REIP_REG_14__SCAN_IN), .ZN(n6174) );
  OAI21_X1 U7155 ( .B1(n6056), .B2(n6005), .A(n6174), .ZN(n6006) );
  AOI211_X1 U7156 ( .C1(n6008), .C2(n6065), .A(n6007), .B(n6006), .ZN(n6009)
         );
  OAI21_X1 U7157 ( .B1(n6245), .B2(n6185), .A(n6009), .ZN(U2972) );
  OAI21_X1 U7158 ( .B1(n6010), .B2(n6012), .A(n6011), .ZN(n6186) );
  NAND2_X1 U7159 ( .A1(n6422), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6013)
         );
  NAND2_X1 U7160 ( .A1(n6457), .A2(REIP_REG_13__SCAN_IN), .ZN(n6191) );
  OAI211_X1 U7161 ( .C1(n6432), .C2(n6263), .A(n6013), .B(n6191), .ZN(n6014)
         );
  AOI21_X1 U7162 ( .B1(n6186), .B2(n6428), .A(n6014), .ZN(n6015) );
  OAI21_X1 U7163 ( .B1(n6016), .B2(n6057), .A(n6015), .ZN(U2973) );
  NAND2_X1 U7164 ( .A1(n6017), .A2(n6037), .ZN(n6030) );
  NOR2_X1 U7165 ( .A1(n4300), .A2(n6206), .ZN(n6028) );
  AOI21_X1 U7166 ( .B1(n6030), .B2(n6026), .A(n6028), .ZN(n6021) );
  OAI21_X1 U7167 ( .B1(n4300), .B2(n6019), .A(n6018), .ZN(n6020) );
  XNOR2_X1 U7168 ( .A(n6021), .B(n6020), .ZN(n6203) );
  INV_X1 U7169 ( .A(n6022), .ZN(n6277) );
  AOI22_X1 U7170 ( .A1(n6422), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6457), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n6023) );
  OAI21_X1 U7171 ( .B1(n6277), .B2(n6432), .A(n6023), .ZN(n6024) );
  AOI21_X1 U7172 ( .B1(n6279), .B2(n6065), .A(n6024), .ZN(n6025) );
  OAI21_X1 U7173 ( .B1(n6203), .B2(n6245), .A(n6025), .ZN(U2974) );
  INV_X1 U7174 ( .A(n6026), .ZN(n6027) );
  NOR2_X1 U7175 ( .A1(n6028), .A2(n6027), .ZN(n6029) );
  XNOR2_X1 U7176 ( .A(n6030), .B(n6029), .ZN(n6212) );
  INV_X1 U7177 ( .A(n6031), .ZN(n6035) );
  NAND2_X1 U7178 ( .A1(n6457), .A2(REIP_REG_11__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7179 ( .A1(n6422), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6032)
         );
  OAI211_X1 U7180 ( .C1(n6432), .C2(n6033), .A(n6204), .B(n6032), .ZN(n6034)
         );
  AOI21_X1 U7181 ( .B1(n6035), .B2(n6065), .A(n6034), .ZN(n6036) );
  OAI21_X1 U7182 ( .B1(n6212), .B2(n6245), .A(n6036), .ZN(U2975) );
  INV_X1 U7183 ( .A(n6037), .ZN(n6039) );
  NOR2_X1 U7184 ( .A1(n6039), .A2(n6038), .ZN(n6041) );
  XOR2_X1 U7185 ( .A(n6041), .B(n6040), .Z(n6225) );
  INV_X1 U7186 ( .A(n6042), .ZN(n6044) );
  AOI22_X1 U7187 ( .A1(n6422), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6457), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n6043) );
  OAI21_X1 U7188 ( .B1(n6432), .B2(n6044), .A(n6043), .ZN(n6045) );
  AOI21_X1 U7189 ( .B1(n6046), .B2(n6065), .A(n6045), .ZN(n6047) );
  OAI21_X1 U7190 ( .B1(n6225), .B2(n6245), .A(n6047), .ZN(U2976) );
  XNOR2_X1 U7191 ( .A(n4300), .B(n7025), .ZN(n6049) );
  XNOR2_X1 U7192 ( .A(n6048), .B(n6049), .ZN(n6437) );
  NAND2_X1 U7193 ( .A1(n6437), .A2(n6428), .ZN(n6053) );
  NOR2_X1 U7194 ( .A1(n6218), .A2(n6838), .ZN(n6434) );
  NOR2_X1 U7195 ( .A1(n6432), .A2(n6050), .ZN(n6051) );
  AOI211_X1 U7196 ( .C1(n6422), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6434), 
        .B(n6051), .ZN(n6052) );
  OAI211_X1 U7197 ( .C1(n6057), .C2(n6054), .A(n6053), .B(n6052), .ZN(U2977)
         );
  OAI21_X1 U7198 ( .B1(n6056), .B2(n6881), .A(n6055), .ZN(n6059) );
  NOR2_X1 U7199 ( .A1(n6288), .A2(n6057), .ZN(n6058) );
  AOI211_X1 U7200 ( .C1(n6060), .C2(n6289), .A(n6059), .B(n6058), .ZN(n6061)
         );
  OAI21_X1 U7201 ( .B1(n6245), .B2(n6062), .A(n6061), .ZN(U2978) );
  OAI21_X1 U7202 ( .B1(n6422), .B2(n6063), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6070) );
  INV_X1 U7203 ( .A(n6064), .ZN(n6066) );
  NAND2_X1 U7204 ( .A1(n6066), .A2(n6065), .ZN(n6069) );
  NAND2_X1 U7205 ( .A1(n6457), .A2(REIP_REG_0__SCAN_IN), .ZN(n6475) );
  OR2_X1 U7206 ( .A1(n6067), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6471)
         );
  NAND3_X1 U7207 ( .A1(n6428), .A2(n3570), .A3(n6471), .ZN(n6068) );
  NAND4_X1 U7208 ( .A1(n6070), .A2(n6069), .A3(n6475), .A4(n6068), .ZN(U2986)
         );
  XNOR2_X1 U7209 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7210 ( .A1(n6071), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6073) );
  OAI211_X1 U7211 ( .C1(n6075), .C2(n6074), .A(n6073), .B(n6072), .ZN(n6076)
         );
  AOI21_X1 U7212 ( .B1(n6077), .B2(n6470), .A(n6076), .ZN(n6078) );
  OAI21_X1 U7213 ( .B1(n6079), .B2(n6473), .A(n6078), .ZN(U2990) );
  NAND3_X1 U7214 ( .A1(n6082), .A2(n6081), .A3(n6080), .ZN(n6083) );
  OAI211_X1 U7215 ( .C1(n6086), .C2(n6085), .A(n6084), .B(n6083), .ZN(n6087)
         );
  AOI21_X1 U7216 ( .B1(n6088), .B2(n6470), .A(n6087), .ZN(n6089) );
  OAI21_X1 U7217 ( .B1(n6090), .B2(n6473), .A(n6089), .ZN(U2992) );
  AOI21_X1 U7218 ( .B1(n6092), .B2(n6094), .A(n6091), .ZN(n6093) );
  OAI21_X1 U7219 ( .B1(n3093), .B2(n6094), .A(n6093), .ZN(n6095) );
  AOI21_X1 U7220 ( .B1(n6096), .B2(n6470), .A(n6095), .ZN(n6097) );
  OAI21_X1 U7221 ( .B1(n6098), .B2(n6473), .A(n6097), .ZN(U2995) );
  NAND3_X1 U7222 ( .A1(n3092), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n6099), .ZN(n6100) );
  OAI211_X1 U7223 ( .C1(n3093), .C2(n6855), .A(n6101), .B(n6100), .ZN(n6102)
         );
  AOI21_X1 U7224 ( .B1(n6103), .B2(n6470), .A(n6102), .ZN(n6104) );
  OAI21_X1 U7225 ( .B1(n6105), .B2(n6473), .A(n6104), .ZN(U2996) );
  NAND2_X1 U7226 ( .A1(n6106), .A2(n6462), .ZN(n6112) );
  NOR2_X1 U7227 ( .A1(n6107), .A2(n6110), .ZN(n6108) );
  AOI211_X1 U7228 ( .C1(n3092), .C2(n6110), .A(n6109), .B(n6108), .ZN(n6111)
         );
  OAI211_X1 U7229 ( .C1(n6221), .C2(n6113), .A(n6112), .B(n6111), .ZN(U2997)
         );
  NAND2_X1 U7230 ( .A1(n6114), .A2(n6462), .ZN(n6126) );
  AOI21_X1 U7231 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6115), .A(n6460), 
        .ZN(n6116) );
  NOR2_X1 U7232 ( .A1(n6117), .A2(n6116), .ZN(n6146) );
  INV_X1 U7233 ( .A(n6146), .ZN(n6118) );
  AOI21_X1 U7234 ( .B1(n6119), .B2(n6959), .A(n6118), .ZN(n6138) );
  OAI21_X1 U7235 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6216), .A(n6138), 
        .ZN(n6132) );
  AND3_X1 U7236 ( .A1(n6122), .A2(n6121), .A3(n6120), .ZN(n6123) );
  AOI211_X1 U7237 ( .C1(n6132), .C2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n6124), .B(n6123), .ZN(n6125) );
  OAI211_X1 U7238 ( .C1(n6127), .C2(n6221), .A(n6126), .B(n6125), .ZN(U2998)
         );
  NAND2_X1 U7239 ( .A1(n6128), .A2(n6462), .ZN(n6134) );
  NOR2_X1 U7240 ( .A1(n6129), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6130)
         );
  AOI211_X1 U7241 ( .C1(n6132), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6131), .B(n6130), .ZN(n6133) );
  OAI211_X1 U7242 ( .C1(n6135), .C2(n6221), .A(n6134), .B(n6133), .ZN(U2999)
         );
  NAND4_X1 U7243 ( .A1(n6143), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n6962), .A4(n3160), .ZN(n6136) );
  OAI211_X1 U7244 ( .C1(n6138), .C2(n6962), .A(n6137), .B(n6136), .ZN(n6139)
         );
  AOI21_X1 U7245 ( .B1(n6140), .B2(n6470), .A(n6139), .ZN(n6141) );
  OAI21_X1 U7246 ( .B1(n6142), .B2(n6473), .A(n6141), .ZN(U3000) );
  NAND3_X1 U7247 ( .A1(n6143), .A2(n6959), .A3(n3160), .ZN(n6144) );
  OAI211_X1 U7248 ( .C1(n6146), .C2(n6959), .A(n6145), .B(n6144), .ZN(n6147)
         );
  AOI21_X1 U7249 ( .B1(n6148), .B2(n6470), .A(n6147), .ZN(n6149) );
  OAI21_X1 U7250 ( .B1(n6150), .B2(n6473), .A(n6149), .ZN(U3001) );
  INV_X1 U7251 ( .A(n6151), .ZN(n6156) );
  INV_X1 U7252 ( .A(n6162), .ZN(n6153) );
  NOR4_X1 U7253 ( .A1(n6153), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6205), 
        .A4(n6152), .ZN(n6154) );
  AOI211_X1 U7254 ( .C1(n6156), .C2(n6470), .A(n6155), .B(n6154), .ZN(n6164)
         );
  INV_X1 U7255 ( .A(n6157), .ZN(n6158) );
  AOI21_X1 U7256 ( .B1(n6160), .B2(n6159), .A(n6158), .ZN(n6207) );
  OAI21_X1 U7257 ( .B1(n6162), .B2(n6216), .A(n6207), .ZN(n6171) );
  NOR2_X1 U7258 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6205), .ZN(n6161)
         );
  AND2_X1 U7259 ( .A1(n6162), .A2(n6161), .ZN(n6166) );
  OAI21_X1 U7260 ( .B1(n6171), .B2(n6166), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n6163) );
  OAI211_X1 U7261 ( .C1(n6165), .C2(n6473), .A(n6164), .B(n6163), .ZN(U3002)
         );
  INV_X1 U7262 ( .A(n6166), .ZN(n6167) );
  OAI211_X1 U7263 ( .C1(n6169), .C2(n6221), .A(n6168), .B(n6167), .ZN(n6170)
         );
  AOI21_X1 U7264 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6171), .A(n6170), 
        .ZN(n6172) );
  OAI21_X1 U7265 ( .B1(n6173), .B2(n6473), .A(n6172), .ZN(U3003) );
  INV_X1 U7266 ( .A(n6174), .ZN(n6177) );
  INV_X1 U7267 ( .A(n6180), .ZN(n6175) );
  NOR3_X1 U7268 ( .A1(n6175), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n6205), 
        .ZN(n6176) );
  AOI211_X1 U7269 ( .C1(n6178), .C2(n6470), .A(n6177), .B(n6176), .ZN(n6184)
         );
  NAND2_X1 U7270 ( .A1(n6460), .A2(n6181), .ZN(n6467) );
  NAND2_X1 U7271 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7272 ( .A1(n6467), .A2(n6187), .ZN(n6179) );
  OAI211_X1 U7273 ( .C1(n6180), .C2(n6479), .A(n6207), .B(n6179), .ZN(n6193)
         );
  AOI21_X1 U7274 ( .B1(n3115), .B2(n6181), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n6182) );
  OAI21_X1 U7275 ( .B1(n6193), .B2(n6182), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n6183) );
  OAI211_X1 U7276 ( .C1(n6185), .C2(n6473), .A(n6184), .B(n6183), .ZN(U3004)
         );
  INV_X1 U7277 ( .A(n6186), .ZN(n6195) );
  INV_X1 U7278 ( .A(n6187), .ZN(n6188) );
  NAND3_X1 U7279 ( .A1(n6189), .A2(n3160), .A3(n6188), .ZN(n6190) );
  OAI211_X1 U7280 ( .C1(n6260), .C2(n6221), .A(n6191), .B(n6190), .ZN(n6192)
         );
  AOI21_X1 U7281 ( .B1(n6193), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n6192), 
        .ZN(n6194) );
  OAI21_X1 U7282 ( .B1(n6195), .B2(n6473), .A(n6194), .ZN(U3005) );
  INV_X1 U7283 ( .A(n6274), .ZN(n6201) );
  OAI21_X1 U7284 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6205), .A(n6207), 
        .ZN(n6197) );
  NOR3_X1 U7285 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6205), .A3(n6206), 
        .ZN(n6196) );
  AOI21_X1 U7286 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6197), .A(n6196), 
        .ZN(n6198) );
  OAI21_X1 U7287 ( .B1(n6218), .B2(n6199), .A(n6198), .ZN(n6200) );
  AOI21_X1 U7288 ( .B1(n6201), .B2(n6470), .A(n6200), .ZN(n6202) );
  OAI21_X1 U7289 ( .B1(n6203), .B2(n6473), .A(n6202), .ZN(U3006) );
  OAI21_X1 U7290 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6205), .A(n6204), 
        .ZN(n6209) );
  NOR2_X1 U7291 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  AOI211_X1 U7292 ( .C1(n6470), .C2(n6210), .A(n6209), .B(n6208), .ZN(n6211)
         );
  OAI21_X1 U7293 ( .B1(n6212), .B2(n6473), .A(n6211), .ZN(U3007) );
  NOR2_X1 U7294 ( .A1(n6213), .A2(n6446), .ZN(n6436) );
  OAI211_X1 U7295 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6436), .B(n6214), .ZN(n6224) );
  OAI21_X1 U7296 ( .B1(n6217), .B2(n6216), .A(n6449), .ZN(n6433) );
  OAI22_X1 U7297 ( .A1(n6221), .A2(n6220), .B1(n6219), .B2(n6218), .ZN(n6222)
         );
  AOI21_X1 U7298 ( .B1(n6433), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6222), 
        .ZN(n6223) );
  OAI211_X1 U7299 ( .C1(n6225), .C2(n6473), .A(n6224), .B(n6223), .ZN(U3008)
         );
  INV_X1 U7300 ( .A(n6226), .ZN(n6720) );
  OAI211_X1 U7301 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6227), .A(n6230), .B(
        n6651), .ZN(n6228) );
  OAI21_X1 U7302 ( .B1(n6720), .B2(n4605), .A(n6228), .ZN(n6229) );
  MUX2_X1 U7303 ( .A(n6229), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(n6732), 
        .Z(U3464) );
  XNOR2_X1 U7304 ( .A(n6231), .B(n6230), .ZN(n6233) );
  OAI22_X1 U7305 ( .A1(n6233), .A2(n6722), .B1(n6232), .B2(n6720), .ZN(n6234)
         );
  MUX2_X1 U7306 ( .A(n6234), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(n6732), 
        .Z(U3463) );
  INV_X1 U7307 ( .A(n6235), .ZN(n6239) );
  OAI22_X1 U7308 ( .A1(n6239), .A2(n6238), .B1(n6237), .B2(n6236), .ZN(n6241)
         );
  MUX2_X1 U7309 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6241), .S(n6240), 
        .Z(U3456) );
  AND2_X1 U7310 ( .A1(n6743), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NOR2_X1 U7311 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6243) );
  OAI21_X1 U7312 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6243), .A(n6740), .ZN(n6242)
         );
  OAI21_X1 U7313 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6740), .A(n6242), .ZN(
        U2791) );
  OAI21_X1 U7314 ( .B1(n6243), .B2(BS16_N), .A(n6719), .ZN(n6718) );
  OAI21_X1 U7315 ( .B1(n6719), .B2(n6244), .A(n6718), .ZN(U2792) );
  OAI21_X1 U7316 ( .B1(n6246), .B2(n6943), .A(n6245), .ZN(U2793) );
  INV_X1 U7317 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6716) );
  INV_X1 U7318 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6994) );
  INV_X1 U7319 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7028) );
  NAND2_X1 U7320 ( .A1(n6994), .A2(n7028), .ZN(n6757) );
  INV_X1 U7321 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6866) );
  INV_X1 U7322 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6872) );
  INV_X1 U7323 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6936) );
  INV_X1 U7324 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6853) );
  OAI211_X1 U7325 ( .C1(n6866), .C2(n6872), .A(n6936), .B(n6853), .ZN(n6247)
         );
  NOR4_X1 U7326 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_25__SCAN_IN), .A3(n6757), .A4(n6247), .ZN(n6255) );
  NOR4_X1 U7327 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6254) );
  NOR4_X1 U7328 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n6253) );
  NOR4_X1 U7329 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6251) );
  NOR4_X1 U7330 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6250) );
  NOR4_X1 U7331 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6249) );
  NOR4_X1 U7332 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6248) );
  AND4_X1 U7333 ( .A1(n6251), .A2(n6250), .A3(n6249), .A4(n6248), .ZN(n6252)
         );
  NAND4_X1 U7334 ( .A1(n6255), .A2(n6254), .A3(n6253), .A4(n6252), .ZN(n6736)
         );
  INV_X1 U7335 ( .A(REIP_REG_0__SCAN_IN), .ZN(n7023) );
  NAND3_X1 U7336 ( .A1(n7023), .A2(n6866), .A3(n6872), .ZN(n6257) );
  NOR2_X1 U7337 ( .A1(n6736), .A2(REIP_REG_1__SCAN_IN), .ZN(n6256) );
  AOI22_X1 U7338 ( .A1(n6716), .A2(n6736), .B1(n6257), .B2(n6256), .ZN(U2794)
         );
  INV_X1 U7339 ( .A(n6736), .ZN(n6738) );
  OAI21_X1 U7340 ( .B1(REIP_REG_1__SCAN_IN), .B2(DATAWIDTH_REG_1__SCAN_IN), 
        .A(n6257), .ZN(n6258) );
  INV_X1 U7341 ( .A(n6258), .ZN(n6259) );
  INV_X1 U7342 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6927) );
  AOI22_X1 U7343 ( .A1(n6738), .A2(n6259), .B1(n6927), .B2(n6736), .ZN(U2795)
         );
  OAI22_X1 U7344 ( .A1(n6261), .A2(n6306), .B1(n6350), .B2(n6260), .ZN(n6262)
         );
  AOI211_X1 U7345 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6333), 
        .B(n6262), .ZN(n6273) );
  NOR2_X1 U7346 ( .A1(n5694), .A2(n6263), .ZN(n6264) );
  AOI21_X1 U7347 ( .B1(n6265), .B2(n6311), .A(n6264), .ZN(n6272) );
  NOR2_X1 U7348 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6266), .ZN(n6267) );
  AND2_X1 U7349 ( .A1(n6359), .A2(n6267), .ZN(n6280) );
  OAI21_X1 U7350 ( .B1(n6280), .B2(n6276), .A(REIP_REG_13__SCAN_IN), .ZN(n6271) );
  NAND3_X1 U7351 ( .A1(n6359), .A2(n6269), .A3(n6268), .ZN(n6270) );
  NAND4_X1 U7352 ( .A1(n6273), .A2(n6272), .A3(n6271), .A4(n6270), .ZN(U2814)
         );
  NOR2_X1 U7353 ( .A1(n6350), .A2(n6274), .ZN(n6275) );
  AOI211_X1 U7354 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6333), 
        .B(n6275), .ZN(n6284) );
  AOI22_X1 U7355 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6365), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6276), .ZN(n6283) );
  NOR2_X1 U7356 ( .A1(n5694), .A2(n6277), .ZN(n6278) );
  AOI21_X1 U7357 ( .B1(n6279), .B2(n6311), .A(n6278), .ZN(n6282) );
  INV_X1 U7358 ( .A(n6280), .ZN(n6281) );
  NAND4_X1 U7359 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(U2815)
         );
  NOR2_X1 U7360 ( .A1(n6285), .A2(REIP_REG_8__SCAN_IN), .ZN(n6293) );
  OAI22_X1 U7361 ( .A1(n6881), .A2(n6347), .B1(n6350), .B2(n6286), .ZN(n6287)
         );
  AOI211_X1 U7362 ( .C1(n6365), .C2(EBX_REG_8__SCAN_IN), .A(n6333), .B(n6287), 
        .ZN(n6292) );
  INV_X1 U7363 ( .A(n6288), .ZN(n6290) );
  AOI22_X1 U7364 ( .A1(n6290), .A2(n6311), .B1(n6364), .B2(n6289), .ZN(n6291)
         );
  OAI211_X1 U7365 ( .C1(n6294), .C2(n6293), .A(n6292), .B(n6291), .ZN(U2819)
         );
  INV_X1 U7366 ( .A(n6295), .ZN(n6300) );
  NOR3_X1 U7367 ( .A1(n6321), .A2(REIP_REG_7__SCAN_IN), .A3(n6296), .ZN(n6299)
         );
  AOI22_X1 U7368 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6365), .B1(n6361), .B2(n6442), 
        .ZN(n6297) );
  OAI211_X1 U7369 ( .C1(n6347), .C2(n3884), .A(n6297), .B(n6312), .ZN(n6298)
         );
  AOI211_X1 U7370 ( .C1(n6300), .C2(n6311), .A(n6299), .B(n6298), .ZN(n6304)
         );
  OAI21_X1 U7371 ( .B1(n6321), .B2(n6302), .A(n6373), .ZN(n6323) );
  AND3_X1 U7372 ( .A1(n6359), .A2(n6302), .A3(n6301), .ZN(n6308) );
  OAI21_X1 U7373 ( .B1(n6323), .B2(n6308), .A(REIP_REG_7__SCAN_IN), .ZN(n6303)
         );
  OAI211_X1 U7374 ( .C1(n5694), .C2(n6305), .A(n6304), .B(n6303), .ZN(U2820)
         );
  AOI22_X1 U7375 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6358), .B1(n6361), 
        .B2(n6374), .ZN(n6315) );
  INV_X1 U7376 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6380) );
  NOR2_X1 U7377 ( .A1(n6380), .A2(n6306), .ZN(n6307) );
  AOI211_X1 U7378 ( .C1(n6323), .C2(REIP_REG_6__SCAN_IN), .A(n6308), .B(n6307), 
        .ZN(n6314) );
  INV_X1 U7379 ( .A(n6309), .ZN(n6310) );
  AOI22_X1 U7380 ( .A1(n6377), .A2(n6311), .B1(n6310), .B2(n6364), .ZN(n6313)
         );
  NAND4_X1 U7381 ( .A1(n6315), .A2(n6314), .A3(n6313), .A4(n6312), .ZN(U2821)
         );
  AOI22_X1 U7382 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n6358), .B1(n6361), 
        .B2(n6316), .ZN(n6317) );
  INV_X1 U7383 ( .A(n6317), .ZN(n6318) );
  AOI211_X1 U7384 ( .C1(n6365), .C2(EBX_REG_5__SCAN_IN), .A(n6333), .B(n6318), 
        .ZN(n6327) );
  OAI21_X1 U7385 ( .B1(n6321), .B2(n6320), .A(n6319), .ZN(n6322) );
  AOI22_X1 U7386 ( .A1(n6325), .A2(n6324), .B1(n6323), .B2(n6322), .ZN(n6326)
         );
  OAI211_X1 U7387 ( .C1(n6328), .C2(n5694), .A(n6327), .B(n6326), .ZN(U2822)
         );
  OAI21_X1 U7388 ( .B1(n6330), .B2(n6335), .A(n6329), .ZN(n6357) );
  INV_X1 U7389 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6897) );
  OAI22_X1 U7390 ( .A1(n6357), .A2(n6331), .B1(n6897), .B2(n6347), .ZN(n6332)
         );
  AOI211_X1 U7391 ( .C1(n6334), .C2(n6362), .A(n6333), .B(n6332), .ZN(n6343)
         );
  NOR2_X1 U7392 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6335), .ZN(n6336) );
  AOI22_X1 U7393 ( .A1(n6365), .A2(EBX_REG_4__SCAN_IN), .B1(n6359), .B2(n6336), 
        .ZN(n6339) );
  NAND2_X1 U7394 ( .A1(n6361), .A2(n6337), .ZN(n6338) );
  OAI211_X1 U7395 ( .C1(n6340), .C2(n6369), .A(n6339), .B(n6338), .ZN(n6341)
         );
  INV_X1 U7396 ( .A(n6341), .ZN(n6342) );
  OAI211_X1 U7397 ( .C1(n6344), .C2(n5694), .A(n6343), .B(n6342), .ZN(U2823)
         );
  NAND2_X1 U7398 ( .A1(n6345), .A2(REIP_REG_2__SCAN_IN), .ZN(n6356) );
  INV_X1 U7399 ( .A(n6346), .ZN(n6349) );
  OAI222_X1 U7400 ( .A1(n6350), .A2(n6349), .B1(n6348), .B2(n6721), .C1(n6347), 
        .C2(n3912), .ZN(n6354) );
  OAI22_X1 U7401 ( .A1(n6352), .A2(n6369), .B1(n6351), .B2(n5694), .ZN(n6353)
         );
  AOI211_X1 U7402 ( .C1(EBX_REG_3__SCAN_IN), .C2(n6365), .A(n6354), .B(n6353), 
        .ZN(n6355) );
  OAI221_X1 U7403 ( .B1(n6357), .B2(n7022), .C1(n6357), .C2(n6356), .A(n6355), 
        .ZN(U2824) );
  AOI22_X1 U7404 ( .A1(n6359), .A2(n6996), .B1(PHYADDRPOINTER_REG_1__SCAN_IN), 
        .B2(n6358), .ZN(n6372) );
  AOI22_X1 U7405 ( .A1(n6363), .A2(n6362), .B1(n6361), .B2(n6360), .ZN(n6367)
         );
  AOI22_X1 U7406 ( .A1(n6365), .A2(EBX_REG_1__SCAN_IN), .B1(n6364), .B2(n6928), 
        .ZN(n6366) );
  OAI211_X1 U7407 ( .C1(n6369), .C2(n6368), .A(n6367), .B(n6366), .ZN(n6370)
         );
  INV_X1 U7408 ( .A(n6370), .ZN(n6371) );
  OAI211_X1 U7409 ( .C1(n6373), .C2(n6996), .A(n6372), .B(n6371), .ZN(U2826)
         );
  AOI22_X1 U7410 ( .A1(n6377), .A2(n6376), .B1(n6375), .B2(n6374), .ZN(n6378)
         );
  OAI21_X1 U7411 ( .B1(n6380), .B2(n6379), .A(n6378), .ZN(U2853) );
  INV_X1 U7412 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n6819) );
  AOI22_X1 U7413 ( .A1(n6381), .A2(EAX_REG_19__SCAN_IN), .B1(n6744), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n6382) );
  OAI21_X1 U7414 ( .B1(n6819), .B2(n6385), .A(n6382), .ZN(U2904) );
  INV_X1 U7415 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n6899) );
  AOI22_X1 U7416 ( .A1(n6383), .A2(EAX_REG_14__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6384) );
  OAI21_X1 U7417 ( .B1(n6899), .B2(n6385), .A(n6384), .ZN(U2909) );
  AOI22_X1 U7418 ( .A1(n6743), .A2(DATAO_REG_13__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6386) );
  OAI21_X1 U7419 ( .B1(n6387), .B2(n6402), .A(n6386), .ZN(U2910) );
  INV_X1 U7420 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6389) );
  AOI22_X1 U7421 ( .A1(n6743), .A2(DATAO_REG_12__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6388) );
  OAI21_X1 U7422 ( .B1(n6389), .B2(n6402), .A(n6388), .ZN(U2911) );
  INV_X1 U7423 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6391) );
  AOI22_X1 U7424 ( .A1(n6743), .A2(DATAO_REG_10__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6390) );
  OAI21_X1 U7425 ( .B1(n6391), .B2(n6402), .A(n6390), .ZN(U2913) );
  AOI22_X1 U7426 ( .A1(n6743), .A2(DATAO_REG_9__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6392) );
  OAI21_X1 U7427 ( .B1(n6965), .B2(n6402), .A(n6392), .ZN(U2914) );
  AOI22_X1 U7428 ( .A1(n6743), .A2(DATAO_REG_7__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n6393) );
  OAI21_X1 U7429 ( .B1(n6784), .B2(n6402), .A(n6393), .ZN(U2916) );
  AOI22_X1 U7430 ( .A1(n6743), .A2(DATAO_REG_5__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n6394) );
  OAI21_X1 U7431 ( .B1(n6395), .B2(n6402), .A(n6394), .ZN(U2918) );
  AOI22_X1 U7432 ( .A1(n6743), .A2(DATAO_REG_4__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n6396) );
  OAI21_X1 U7433 ( .B1(n6397), .B2(n6402), .A(n6396), .ZN(U2919) );
  AOI22_X1 U7434 ( .A1(n6743), .A2(DATAO_REG_2__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n6398) );
  OAI21_X1 U7435 ( .B1(n6399), .B2(n6402), .A(n6398), .ZN(U2921) );
  AOI22_X1 U7436 ( .A1(n6743), .A2(DATAO_REG_1__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n6400) );
  OAI21_X1 U7437 ( .B1(n6823), .B2(n6402), .A(n6400), .ZN(U2922) );
  AOI22_X1 U7438 ( .A1(n6743), .A2(DATAO_REG_0__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n6401) );
  OAI21_X1 U7439 ( .B1(n6403), .B2(n6402), .A(n6401), .ZN(U2923) );
  AOI22_X1 U7440 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6415), .B1(n6418), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U7441 ( .A1(n6419), .A2(DATAI_8_), .ZN(n6409) );
  NAND2_X1 U7442 ( .A1(n6404), .A2(n6409), .ZN(U2932) );
  AOI22_X1 U7443 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6415), .B1(n6418), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U7444 ( .A1(n6419), .A2(DATAI_10_), .ZN(n6411) );
  NAND2_X1 U7445 ( .A1(n6405), .A2(n6411), .ZN(U2934) );
  AOI22_X1 U7446 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6415), .B1(n6418), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U7447 ( .A1(n6419), .A2(DATAI_11_), .ZN(n6413) );
  NAND2_X1 U7448 ( .A1(n6406), .A2(n6413), .ZN(U2935) );
  NAND2_X1 U7449 ( .A1(n6419), .A2(DATAI_14_), .ZN(n6416) );
  INV_X1 U7450 ( .A(n6416), .ZN(n6407) );
  AOI21_X1 U7451 ( .B1(n6418), .B2(UWORD_REG_14__SCAN_IN), .A(n6407), .ZN(
        n6408) );
  OAI21_X1 U7452 ( .B1(n4401), .B2(n6421), .A(n6408), .ZN(U2938) );
  AOI22_X1 U7453 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6415), .B1(
        LWORD_REG_8__SCAN_IN), .B2(n6418), .ZN(n6410) );
  NAND2_X1 U7454 ( .A1(n6410), .A2(n6409), .ZN(U2947) );
  AOI22_X1 U7455 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6415), .B1(n6418), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U7456 ( .A1(n6412), .A2(n6411), .ZN(U2949) );
  AOI22_X1 U7457 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6415), .B1(
        LWORD_REG_11__SCAN_IN), .B2(n6418), .ZN(n6414) );
  NAND2_X1 U7458 ( .A1(n6414), .A2(n6413), .ZN(U2950) );
  AOI22_X1 U7459 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6415), .B1(n6418), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U7460 ( .A1(n6417), .A2(n6416), .ZN(U2953) );
  AOI22_X1 U7461 ( .A1(n6419), .A2(DATAI_15_), .B1(n6418), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6420) );
  OAI21_X1 U7462 ( .B1(n6997), .B2(n6421), .A(n6420), .ZN(U2954) );
  AOI22_X1 U7463 ( .A1(n6422), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6457), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U7464 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  XOR2_X1 U7465 ( .A(n6426), .B(n6425), .Z(n6463) );
  AOI22_X1 U7466 ( .A1(n6463), .A2(n6428), .B1(n6427), .B2(n6065), .ZN(n6429)
         );
  OAI211_X1 U7467 ( .C1(n6432), .C2(n6431), .A(n6430), .B(n6429), .ZN(U2984)
         );
  INV_X1 U7468 ( .A(n6433), .ZN(n6440) );
  AOI21_X1 U7469 ( .B1(n6435), .B2(n6470), .A(n6434), .ZN(n6439) );
  AOI22_X1 U7470 ( .A1(n6437), .A2(n6462), .B1(n6436), .B2(n7025), .ZN(n6438)
         );
  OAI211_X1 U7471 ( .C1(n6440), .C2(n7025), .A(n6439), .B(n6438), .ZN(U3009)
         );
  AOI21_X1 U7472 ( .B1(n6470), .B2(n6442), .A(n6441), .ZN(n6445) );
  NAND2_X1 U7473 ( .A1(n6443), .A2(n6462), .ZN(n6444) );
  OAI211_X1 U7474 ( .C1(n6446), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6445), 
        .B(n6444), .ZN(n6447) );
  INV_X1 U7475 ( .A(n6447), .ZN(n6448) );
  OAI21_X1 U7476 ( .B1(n6449), .B2(n6930), .A(n6448), .ZN(U3011) );
  INV_X1 U7477 ( .A(n6450), .ZN(n6451) );
  AOI22_X1 U7478 ( .A1(n6470), .A2(n6453), .B1(n6452), .B2(n6451), .ZN(n6465)
         );
  NOR3_X1 U7479 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n6455), .A3(n6454), 
        .ZN(n6456) );
  AOI21_X1 U7480 ( .B1(n6457), .B2(REIP_REG_2__SCAN_IN), .A(n6456), .ZN(n6458)
         );
  OAI21_X1 U7481 ( .B1(n6460), .B2(n6459), .A(n6458), .ZN(n6461) );
  AOI21_X1 U7482 ( .B1(n6463), .B2(n6462), .A(n6461), .ZN(n6464) );
  OAI211_X1 U7483 ( .C1(n6466), .C2(n3579), .A(n6465), .B(n6464), .ZN(U3016)
         );
  NAND2_X1 U7484 ( .A1(n6467), .A2(n6481), .ZN(n6477) );
  INV_X1 U7485 ( .A(n6468), .ZN(n6469) );
  NAND2_X1 U7486 ( .A1(n6470), .A2(n6469), .ZN(n6476) );
  NAND2_X1 U7487 ( .A1(n6471), .A2(n3570), .ZN(n6472) );
  OR2_X1 U7488 ( .A1(n6473), .A2(n6472), .ZN(n6474) );
  AND4_X1 U7489 ( .A1(n6477), .A2(n6476), .A3(n6475), .A4(n6474), .ZN(n6478)
         );
  OAI221_X1 U7490 ( .B1(n6481), .B2(n6480), .C1(n6481), .C2(n6479), .A(n6478), 
        .ZN(U3018) );
  INV_X1 U7491 ( .A(n6732), .ZN(n6729) );
  NOR2_X1 U7492 ( .A1(n6482), .A2(n6729), .ZN(U3019) );
  INV_X1 U7493 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6487) );
  NOR2_X1 U7494 ( .A1(n6596), .A2(n6488), .ZN(n6483) );
  AOI21_X1 U7495 ( .B1(n6490), .B2(n6658), .A(n6483), .ZN(n6486) );
  INV_X1 U7496 ( .A(n6484), .ZN(n6492) );
  AOI22_X1 U7497 ( .A1(n6492), .A2(n6554), .B1(n6657), .B2(n6491), .ZN(n6485)
         );
  OAI211_X1 U7498 ( .C1(n6495), .C2(n6487), .A(n6486), .B(n6485), .ZN(U3029)
         );
  INV_X1 U7499 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6847) );
  NOR2_X1 U7500 ( .A1(n6601), .A2(n6488), .ZN(n6489) );
  AOI21_X1 U7501 ( .B1(n6490), .B2(n6663), .A(n6489), .ZN(n6494) );
  AOI22_X1 U7502 ( .A1(n6492), .A2(n6558), .B1(n6664), .B2(n6491), .ZN(n6493)
         );
  OAI211_X1 U7503 ( .C1(n6495), .C2(n6847), .A(n6494), .B(n6493), .ZN(U3030)
         );
  NOR2_X1 U7504 ( .A1(n6496), .A2(n6541), .ZN(n6501) );
  AOI21_X1 U7505 ( .B1(n6497), .B2(n4623), .A(n6501), .ZN(n6503) );
  INV_X1 U7506 ( .A(n6503), .ZN(n6498) );
  INV_X1 U7507 ( .A(n6501), .ZN(n6527) );
  OAI22_X1 U7508 ( .A1(n6551), .A2(n6587), .B1(n6586), .B2(n6527), .ZN(n6502)
         );
  INV_X1 U7509 ( .A(n6502), .ZN(n6508) );
  NAND2_X1 U7510 ( .A1(n6504), .A2(n6503), .ZN(n6505) );
  OAI211_X1 U7511 ( .C1(n6651), .C2(n6506), .A(n6505), .B(n6648), .ZN(n6530)
         );
  AOI22_X1 U7512 ( .A1(n6530), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n6652), 
        .B2(n6529), .ZN(n6507) );
  OAI211_X1 U7513 ( .C1(n6533), .C2(n6655), .A(n6508), .B(n6507), .ZN(U3060)
         );
  OAI22_X1 U7514 ( .A1(n6551), .A2(n6557), .B1(n6596), .B2(n6527), .ZN(n6509)
         );
  INV_X1 U7515 ( .A(n6509), .ZN(n6511) );
  AOI22_X1 U7516 ( .A1(n6530), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n6658), 
        .B2(n6529), .ZN(n6510) );
  OAI211_X1 U7517 ( .C1(n6533), .C2(n6661), .A(n6511), .B(n6510), .ZN(U3061)
         );
  OAI22_X1 U7518 ( .A1(n6551), .A2(n6561), .B1(n6601), .B2(n6527), .ZN(n6512)
         );
  INV_X1 U7519 ( .A(n6512), .ZN(n6514) );
  AOI22_X1 U7520 ( .A1(n6530), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n6663), 
        .B2(n6529), .ZN(n6513) );
  OAI211_X1 U7521 ( .C1(n6533), .C2(n6667), .A(n6514), .B(n6513), .ZN(U3062)
         );
  OAI22_X1 U7522 ( .A1(n6551), .A2(n6607), .B1(n6606), .B2(n6527), .ZN(n6515)
         );
  INV_X1 U7523 ( .A(n6515), .ZN(n6517) );
  AOI22_X1 U7524 ( .A1(n6530), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n6669), 
        .B2(n6529), .ZN(n6516) );
  OAI211_X1 U7525 ( .C1(n6533), .C2(n6673), .A(n6517), .B(n6516), .ZN(U3063)
         );
  OAI22_X1 U7526 ( .A1(n6551), .A2(n6568), .B1(n6611), .B2(n6527), .ZN(n6518)
         );
  INV_X1 U7527 ( .A(n6518), .ZN(n6520) );
  AOI22_X1 U7528 ( .A1(n6530), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n6675), 
        .B2(n6529), .ZN(n6519) );
  OAI211_X1 U7529 ( .C1(n6533), .C2(n6679), .A(n6520), .B(n6519), .ZN(U3064)
         );
  OAI22_X1 U7530 ( .A1(n6551), .A2(n6617), .B1(n6616), .B2(n6527), .ZN(n6521)
         );
  INV_X1 U7531 ( .A(n6521), .ZN(n6523) );
  AOI22_X1 U7532 ( .A1(n6530), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n6681), 
        .B2(n6529), .ZN(n6522) );
  OAI211_X1 U7533 ( .C1(n6533), .C2(n6685), .A(n6523), .B(n6522), .ZN(U3065)
         );
  OAI22_X1 U7534 ( .A1(n6551), .A2(n6622), .B1(n6621), .B2(n6527), .ZN(n6524)
         );
  INV_X1 U7535 ( .A(n6524), .ZN(n6526) );
  AOI22_X1 U7536 ( .A1(n6530), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n6687), 
        .B2(n6529), .ZN(n6525) );
  OAI211_X1 U7537 ( .C1(n6533), .C2(n6691), .A(n6526), .B(n6525), .ZN(U3066)
         );
  OAI22_X1 U7538 ( .A1(n6551), .A2(n6582), .B1(n6628), .B2(n6527), .ZN(n6528)
         );
  INV_X1 U7539 ( .A(n6528), .ZN(n6532) );
  AOI22_X1 U7540 ( .A1(n6530), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n6697), 
        .B2(n6529), .ZN(n6531) );
  OAI211_X1 U7541 ( .C1(n6533), .C2(n6701), .A(n6532), .B(n6531), .ZN(U3067)
         );
  INV_X1 U7542 ( .A(n6534), .ZN(n6535) );
  INV_X1 U7543 ( .A(n6536), .ZN(n6540) );
  INV_X1 U7544 ( .A(n6537), .ZN(n6538) );
  OAI22_X1 U7545 ( .A1(n6540), .A2(n6545), .B1(n6539), .B2(n6538), .ZN(n6577)
         );
  NAND2_X1 U7546 ( .A1(n6593), .A2(n6541), .ZN(n6547) );
  INV_X1 U7547 ( .A(n6547), .ZN(n6575) );
  AOI22_X1 U7548 ( .A1(n6577), .A2(n6542), .B1(n6643), .B2(n6575), .ZN(n6553)
         );
  NOR2_X1 U7549 ( .A1(n6625), .A2(n6722), .ZN(n6543) );
  AOI21_X1 U7550 ( .B1(n6543), .B2(n6551), .A(n6728), .ZN(n6550) );
  NOR2_X1 U7551 ( .A1(n6545), .A2(n6544), .ZN(n6584) );
  AOI211_X1 U7552 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6547), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6546), .ZN(n6548) );
  AOI22_X1 U7553 ( .A1(n6579), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6652), 
        .B2(n6578), .ZN(n6552) );
  OAI211_X1 U7554 ( .C1(n6587), .C2(n6631), .A(n6553), .B(n6552), .ZN(U3068)
         );
  AOI22_X1 U7555 ( .A1(n6577), .A2(n6554), .B1(n6656), .B2(n6575), .ZN(n6556)
         );
  AOI22_X1 U7556 ( .A1(n6579), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6658), 
        .B2(n6578), .ZN(n6555) );
  OAI211_X1 U7557 ( .C1(n6557), .C2(n6631), .A(n6556), .B(n6555), .ZN(U3069)
         );
  AOI22_X1 U7558 ( .A1(n6577), .A2(n6558), .B1(n6662), .B2(n6575), .ZN(n6560)
         );
  AOI22_X1 U7559 ( .A1(n6579), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6663), 
        .B2(n6578), .ZN(n6559) );
  OAI211_X1 U7560 ( .C1(n6561), .C2(n6631), .A(n6560), .B(n6559), .ZN(U3070)
         );
  AOI22_X1 U7561 ( .A1(n6577), .A2(n6562), .B1(n6668), .B2(n6575), .ZN(n6564)
         );
  AOI22_X1 U7562 ( .A1(n6579), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6669), 
        .B2(n6578), .ZN(n6563) );
  OAI211_X1 U7563 ( .C1(n6607), .C2(n6631), .A(n6564), .B(n6563), .ZN(U3071)
         );
  AOI22_X1 U7564 ( .A1(n6577), .A2(n6565), .B1(n6674), .B2(n6575), .ZN(n6567)
         );
  AOI22_X1 U7565 ( .A1(n6579), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6675), 
        .B2(n6578), .ZN(n6566) );
  OAI211_X1 U7566 ( .C1(n6568), .C2(n6631), .A(n6567), .B(n6566), .ZN(U3072)
         );
  AOI22_X1 U7567 ( .A1(n6577), .A2(n6569), .B1(n6680), .B2(n6575), .ZN(n6571)
         );
  AOI22_X1 U7568 ( .A1(n6579), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6681), 
        .B2(n6578), .ZN(n6570) );
  OAI211_X1 U7569 ( .C1(n6617), .C2(n6631), .A(n6571), .B(n6570), .ZN(U3073)
         );
  AOI22_X1 U7570 ( .A1(n6577), .A2(n6572), .B1(n6686), .B2(n6575), .ZN(n6574)
         );
  AOI22_X1 U7571 ( .A1(n6579), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6687), 
        .B2(n6578), .ZN(n6573) );
  OAI211_X1 U7572 ( .C1(n6622), .C2(n6631), .A(n6574), .B(n6573), .ZN(U3074)
         );
  AOI22_X1 U7573 ( .A1(n6577), .A2(n6576), .B1(n6693), .B2(n6575), .ZN(n6581)
         );
  AOI22_X1 U7574 ( .A1(n6579), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6697), 
        .B2(n6578), .ZN(n6580) );
  OAI211_X1 U7575 ( .C1(n6582), .C2(n6631), .A(n6581), .B(n6580), .ZN(U3075)
         );
  INV_X1 U7576 ( .A(n6629), .ZN(n6583) );
  AOI21_X1 U7577 ( .B1(n6584), .B2(n4623), .A(n6583), .ZN(n6591) );
  NOR2_X1 U7578 ( .A1(n6591), .A2(n6722), .ZN(n6585) );
  AOI21_X1 U7579 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6593), .A(n6585), .ZN(
        n6637) );
  OAI22_X1 U7580 ( .A1(n6623), .A2(n6587), .B1(n6629), .B2(n6586), .ZN(n6588)
         );
  INV_X1 U7581 ( .A(n6588), .ZN(n6595) );
  INV_X1 U7582 ( .A(n6589), .ZN(n6590) );
  NAND2_X1 U7583 ( .A1(n6590), .A2(n6638), .ZN(n6723) );
  NAND3_X1 U7584 ( .A1(n6723), .A2(n6651), .A3(n6591), .ZN(n6592) );
  OAI211_X1 U7585 ( .C1(n6593), .C2(n6651), .A(n6592), .B(n6648), .ZN(n6634)
         );
  AOI22_X1 U7586 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6634), .B1(n6652), 
        .B2(n6625), .ZN(n6594) );
  OAI211_X1 U7587 ( .C1(n6637), .C2(n6655), .A(n6595), .B(n6594), .ZN(U3076)
         );
  OAI22_X1 U7588 ( .A1(n6631), .A2(n6597), .B1(n6629), .B2(n6596), .ZN(n6598)
         );
  INV_X1 U7589 ( .A(n6598), .ZN(n6600) );
  AOI22_X1 U7590 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6634), .B1(n6657), 
        .B2(n6633), .ZN(n6599) );
  OAI211_X1 U7591 ( .C1(n6637), .C2(n6661), .A(n6600), .B(n6599), .ZN(U3077)
         );
  OAI22_X1 U7592 ( .A1(n6631), .A2(n6602), .B1(n6629), .B2(n6601), .ZN(n6603)
         );
  INV_X1 U7593 ( .A(n6603), .ZN(n6605) );
  AOI22_X1 U7594 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6634), .B1(n6664), 
        .B2(n6633), .ZN(n6604) );
  OAI211_X1 U7595 ( .C1(n6637), .C2(n6667), .A(n6605), .B(n6604), .ZN(U3078)
         );
  OAI22_X1 U7596 ( .A1(n6623), .A2(n6607), .B1(n6629), .B2(n6606), .ZN(n6608)
         );
  INV_X1 U7597 ( .A(n6608), .ZN(n6610) );
  AOI22_X1 U7598 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6634), .B1(n6669), 
        .B2(n6625), .ZN(n6609) );
  OAI211_X1 U7599 ( .C1(n6637), .C2(n6673), .A(n6610), .B(n6609), .ZN(U3079)
         );
  OAI22_X1 U7600 ( .A1(n6631), .A2(n6612), .B1(n6629), .B2(n6611), .ZN(n6613)
         );
  INV_X1 U7601 ( .A(n6613), .ZN(n6615) );
  AOI22_X1 U7602 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6634), .B1(n6676), 
        .B2(n6633), .ZN(n6614) );
  OAI211_X1 U7603 ( .C1(n6637), .C2(n6679), .A(n6615), .B(n6614), .ZN(U3080)
         );
  OAI22_X1 U7604 ( .A1(n6623), .A2(n6617), .B1(n6629), .B2(n6616), .ZN(n6618)
         );
  INV_X1 U7605 ( .A(n6618), .ZN(n6620) );
  AOI22_X1 U7606 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6634), .B1(n6681), 
        .B2(n6625), .ZN(n6619) );
  OAI211_X1 U7607 ( .C1(n6637), .C2(n6685), .A(n6620), .B(n6619), .ZN(U3081)
         );
  OAI22_X1 U7608 ( .A1(n6623), .A2(n6622), .B1(n6629), .B2(n6621), .ZN(n6624)
         );
  INV_X1 U7609 ( .A(n6624), .ZN(n6627) );
  AOI22_X1 U7610 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6634), .B1(n6687), 
        .B2(n6625), .ZN(n6626) );
  OAI211_X1 U7611 ( .C1(n6637), .C2(n6691), .A(n6627), .B(n6626), .ZN(U3082)
         );
  OAI22_X1 U7612 ( .A1(n6631), .A2(n6630), .B1(n6629), .B2(n6628), .ZN(n6632)
         );
  INV_X1 U7613 ( .A(n6632), .ZN(n6636) );
  AOI22_X1 U7614 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6634), .B1(n6694), 
        .B2(n6633), .ZN(n6635) );
  OAI211_X1 U7615 ( .C1(n6637), .C2(n6701), .A(n6636), .B(n6635), .ZN(U3083)
         );
  AOI21_X1 U7616 ( .B1(n6639), .B2(n6638), .A(n6722), .ZN(n6647) );
  NAND2_X1 U7617 ( .A1(n6640), .A2(n4623), .ZN(n6641) );
  NAND2_X1 U7618 ( .A1(n6650), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U7619 ( .A1(n6641), .A2(n6642), .ZN(n6645) );
  INV_X1 U7620 ( .A(n6642), .ZN(n6692) );
  AOI22_X1 U7621 ( .A1(n6695), .A2(n6644), .B1(n6643), .B2(n6692), .ZN(n6654)
         );
  INV_X1 U7622 ( .A(n6645), .ZN(n6646) );
  NAND2_X1 U7623 ( .A1(n6647), .A2(n6646), .ZN(n6649) );
  OAI211_X1 U7624 ( .C1(n6651), .C2(n6650), .A(n6649), .B(n6648), .ZN(n6698)
         );
  AOI22_X1 U7625 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6698), .B1(n6652), 
        .B2(n6696), .ZN(n6653) );
  OAI211_X1 U7626 ( .C1(n6702), .C2(n6655), .A(n6654), .B(n6653), .ZN(U3108)
         );
  AOI22_X1 U7627 ( .A1(n6695), .A2(n6657), .B1(n6656), .B2(n6692), .ZN(n6660)
         );
  AOI22_X1 U7628 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6698), .B1(n6658), 
        .B2(n6696), .ZN(n6659) );
  OAI211_X1 U7629 ( .C1(n6702), .C2(n6661), .A(n6660), .B(n6659), .ZN(U3109)
         );
  AOI22_X1 U7630 ( .A1(n6696), .A2(n6663), .B1(n6662), .B2(n6692), .ZN(n6666)
         );
  AOI22_X1 U7631 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6698), .B1(n6664), 
        .B2(n6695), .ZN(n6665) );
  OAI211_X1 U7632 ( .C1(n6702), .C2(n6667), .A(n6666), .B(n6665), .ZN(U3110)
         );
  AOI22_X1 U7633 ( .A1(n6696), .A2(n6669), .B1(n6668), .B2(n6692), .ZN(n6672)
         );
  AOI22_X1 U7634 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6698), .B1(n6670), 
        .B2(n6695), .ZN(n6671) );
  OAI211_X1 U7635 ( .C1(n6702), .C2(n6673), .A(n6672), .B(n6671), .ZN(U3111)
         );
  AOI22_X1 U7636 ( .A1(n6696), .A2(n6675), .B1(n6674), .B2(n6692), .ZN(n6678)
         );
  AOI22_X1 U7637 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6698), .B1(n6676), 
        .B2(n6695), .ZN(n6677) );
  OAI211_X1 U7638 ( .C1(n6702), .C2(n6679), .A(n6678), .B(n6677), .ZN(U3112)
         );
  AOI22_X1 U7639 ( .A1(n6696), .A2(n6681), .B1(n6680), .B2(n6692), .ZN(n6684)
         );
  AOI22_X1 U7640 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6698), .B1(n6682), 
        .B2(n6695), .ZN(n6683) );
  OAI211_X1 U7641 ( .C1(n6702), .C2(n6685), .A(n6684), .B(n6683), .ZN(U3113)
         );
  AOI22_X1 U7642 ( .A1(n6696), .A2(n6687), .B1(n6686), .B2(n6692), .ZN(n6690)
         );
  AOI22_X1 U7643 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6698), .B1(n6688), 
        .B2(n6695), .ZN(n6689) );
  OAI211_X1 U7644 ( .C1(n6702), .C2(n6691), .A(n6690), .B(n6689), .ZN(U3114)
         );
  AOI22_X1 U7645 ( .A1(n6695), .A2(n6694), .B1(n6693), .B2(n6692), .ZN(n6700)
         );
  AOI22_X1 U7646 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6698), .B1(n6697), 
        .B2(n6696), .ZN(n6699) );
  OAI211_X1 U7647 ( .C1(n6702), .C2(n6701), .A(n6700), .B(n6699), .ZN(U3115)
         );
  NOR3_X1 U7648 ( .A1(n6705), .A2(n6704), .A3(n6703), .ZN(n6713) );
  NAND3_X1 U7649 ( .A1(n6707), .A2(STATE2_REG_0__SCAN_IN), .A3(n6706), .ZN(
        n6710) );
  INV_X1 U7650 ( .A(n6708), .ZN(n6709) );
  AOI21_X1 U7651 ( .B1(n6711), .B2(n6710), .A(n6709), .ZN(n6712) );
  OR3_X1 U7652 ( .A1(n6714), .A2(n6713), .A3(n6712), .ZN(U3149) );
  AND2_X1 U7653 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6715), .ZN(U3151) );
  AND2_X1 U7654 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6715), .ZN(U3152) );
  AND2_X1 U7655 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6715), .ZN(U3153) );
  AND2_X1 U7656 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6715), .ZN(U3154) );
  AND2_X1 U7657 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6715), .ZN(U3155) );
  AND2_X1 U7658 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6715), .ZN(U3156) );
  INV_X1 U7659 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6903) );
  NOR2_X1 U7660 ( .A1(n6719), .A2(n6903), .ZN(U3157) );
  AND2_X1 U7661 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6715), .ZN(U3158) );
  AND2_X1 U7662 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6715), .ZN(U3159) );
  AND2_X1 U7663 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6715), .ZN(U3160) );
  AND2_X1 U7664 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6715), .ZN(U3161) );
  AND2_X1 U7665 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6715), .ZN(U3162) );
  AND2_X1 U7666 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6715), .ZN(U3163) );
  AND2_X1 U7667 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6715), .ZN(U3164) );
  AND2_X1 U7668 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6715), .ZN(U3165) );
  AND2_X1 U7669 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6715), .ZN(U3166) );
  AND2_X1 U7670 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6715), .ZN(U3167) );
  AND2_X1 U7671 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6715), .ZN(U3168) );
  AND2_X1 U7672 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6715), .ZN(U3169) );
  AND2_X1 U7673 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6715), .ZN(U3170) );
  AND2_X1 U7674 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6715), .ZN(U3171) );
  AND2_X1 U7675 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6715), .ZN(U3172) );
  NOR2_X1 U7676 ( .A1(n6719), .A2(n7028), .ZN(U3173) );
  NOR2_X1 U7677 ( .A1(n6719), .A2(n6936), .ZN(U3174) );
  AND2_X1 U7678 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6715), .ZN(U3175) );
  NOR2_X1 U7679 ( .A1(n6719), .A2(n6994), .ZN(U3176) );
  NOR2_X1 U7680 ( .A1(n6719), .A2(n6853), .ZN(U3177) );
  AND2_X1 U7681 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6715), .ZN(U3178) );
  AND2_X1 U7682 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6715), .ZN(U3179) );
  AND2_X1 U7683 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6715), .ZN(U3180) );
  INV_X1 U7684 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n7004) );
  AOI22_X1 U7685 ( .A1(n6742), .A2(n6927), .B1(n7004), .B2(n6740), .ZN(U3445)
         );
  MUX2_X1 U7686 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6740), .Z(U3446) );
  INV_X1 U7687 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6988) );
  AOI22_X1 U7688 ( .A1(n6742), .A2(n6716), .B1(n6988), .B2(n6740), .ZN(U3447)
         );
  MUX2_X1 U7689 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6740), .Z(U3448) );
  OAI21_X1 U7690 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6719), .A(n6718), .ZN(
        n6717) );
  INV_X1 U7691 ( .A(n6717), .ZN(U3451) );
  OAI21_X1 U7692 ( .B1(n6719), .B2(n6872), .A(n6718), .ZN(U3452) );
  NOR2_X1 U7693 ( .A1(n6721), .A2(n6720), .ZN(n6726) );
  AOI21_X1 U7694 ( .B1(n6724), .B2(n6723), .A(n6722), .ZN(n6725) );
  AOI211_X1 U7695 ( .C1(n6728), .C2(n6727), .A(n6726), .B(n6725), .ZN(n6730)
         );
  AOI22_X1 U7696 ( .A1(n6732), .A2(n6731), .B1(n6730), .B2(n6729), .ZN(U3462)
         );
  AOI211_X1 U7697 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(REIP_REG_1__SCAN_IN), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6733) );
  AOI21_X1 U7698 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6733), .ZN(n6735) );
  INV_X1 U7699 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6734) );
  AOI22_X1 U7700 ( .A1(n6738), .A2(n6735), .B1(n6734), .B2(n6736), .ZN(U3468)
         );
  NOR2_X1 U7701 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6737) );
  INV_X1 U7702 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7038) );
  AOI22_X1 U7703 ( .A1(n6738), .A2(n6737), .B1(n7038), .B2(n6736), .ZN(U3469)
         );
  NAND2_X1 U7704 ( .A1(n6740), .A2(W_R_N_REG_SCAN_IN), .ZN(n6739) );
  OAI21_X1 U7705 ( .B1(n6740), .B2(READREQUEST_REG_SCAN_IN), .A(n6739), .ZN(
        U3470) );
  INV_X1 U7706 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6885) );
  AOI22_X1 U7707 ( .A1(n6742), .A2(n6741), .B1(n6885), .B2(n6740), .ZN(U3473)
         );
  NAND2_X1 U7708 ( .A1(n6743), .A2(DATAO_REG_21__SCAN_IN), .ZN(n6746) );
  NAND2_X1 U7709 ( .A1(n6744), .A2(UWORD_REG_5__SCAN_IN), .ZN(n6745) );
  OAI211_X1 U7710 ( .C1(n6748), .C2(n6747), .A(n6746), .B(n6745), .ZN(n6749)
         );
  INV_X1 U7711 ( .A(n6749), .ZN(n7060) );
  INV_X1 U7712 ( .A(keyinput15), .ZN(n7058) );
  NOR4_X1 U7713 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(DATAO_REG_19__SCAN_IN), 
        .A3(ADDRESS_REG_17__SCAN_IN), .A4(n6823), .ZN(n6799) );
  INV_X1 U7714 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6817) );
  NOR4_X1 U7715 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(LWORD_REG_4__SCAN_IN), 
        .A3(LWORD_REG_11__SCAN_IN), .A4(n6817), .ZN(n6798) );
  INV_X1 U7716 ( .A(DATAI_30_), .ZN(n6832) );
  NOR4_X1 U7717 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        REIP_REG_9__SCAN_IN), .A3(DATAO_REG_15__SCAN_IN), .A4(n6832), .ZN(
        n6750) );
  NAND3_X1 U7718 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(UWORD_REG_2__SCAN_IN), 
        .A3(n6750), .ZN(n6756) );
  INV_X1 U7719 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6801) );
  NAND4_X1 U7720 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(ADDRESS_REG_11__SCAN_IN), .A4(
        n6801), .ZN(n6754) );
  INV_X1 U7721 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6807) );
  NAND4_X1 U7722 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n6807), .A3(n5331), .A4(n6804), .ZN(n6753) );
  INV_X1 U7723 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6852) );
  NAND4_X1 U7724 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(LWORD_REG_9__SCAN_IN), 
        .A3(n6852), .A4(n6849), .ZN(n6752) );
  NAND4_X1 U7725 ( .A1(ADDRESS_REG_24__SCAN_IN), .A2(n6847), .A3(n4831), .A4(
        n6850), .ZN(n6751) );
  OR4_X1 U7726 ( .A1(n6754), .A2(n6753), .A3(n6752), .A4(n6751), .ZN(n6755) );
  NOR4_X1 U7727 ( .A1(STATE_REG_2__SCAN_IN), .A2(n5324), .A3(n6756), .A4(n6755), .ZN(n6797) );
  NAND2_X1 U7728 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .ZN(
        n6758) );
  NOR4_X1 U7729 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(n6759), .A3(n6758), 
        .A4(n6757), .ZN(n6767) );
  INV_X1 U7730 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n7034) );
  NOR4_X1 U7731 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_0__SCAN_IN), .A3(n7034), .A4(n7037), .ZN(n6766) );
  NOR4_X1 U7732 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(DATAO_REG_11__SCAN_IN), .A3(BE_N_REG_1__SCAN_IN), .A4(n6997), .ZN(n6765) );
  INV_X1 U7733 ( .A(DATAI_31_), .ZN(n7012) );
  NAND4_X1 U7734 ( .A1(DATAI_27_), .A2(ADDRESS_REG_13__SCAN_IN), .A3(n7012), 
        .A4(n7009), .ZN(n6763) );
  INV_X1 U7735 ( .A(DATAI_17_), .ZN(n7007) );
  NAND4_X1 U7736 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(LWORD_REG_8__SCAN_IN), 
        .A3(n7013), .A4(n7007), .ZN(n6762) );
  INV_X1 U7737 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n7020) );
  NAND4_X1 U7738 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        REIP_REG_0__SCAN_IN), .A3(n7020), .A4(n7022), .ZN(n6761) );
  INV_X1 U7739 ( .A(EBX_REG_24__SCAN_IN), .ZN(n7043) );
  NAND4_X1 U7740 ( .A1(EBX_REG_18__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        DATAO_REG_3__SCAN_IN), .A4(n7043), .ZN(n6760) );
  NOR4_X1 U7741 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(n6764)
         );
  NAND4_X1 U7742 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6795)
         );
  NOR4_X1 U7743 ( .A1(EAX_REG_21__SCAN_IN), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .A3(DATAI_18_), .A4(n6978), .ZN(n6771) );
  INV_X1 U7744 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6932) );
  INV_X1 U7745 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6933) );
  NOR4_X1 U7746 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .A3(n6932), .A4(n6933), .ZN(n6770) );
  NOR4_X1 U7747 ( .A1(EAX_REG_9__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        UWORD_REG_13__SCAN_IN), .A4(n6964), .ZN(n6769) );
  INV_X1 U7748 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6975) );
  NOR4_X1 U7749 ( .A1(ADDRESS_REG_27__SCAN_IN), .A2(n4401), .A3(n6975), .A4(
        n6958), .ZN(n6768) );
  NAND4_X1 U7750 ( .A1(n6771), .A2(n6770), .A3(n6769), .A4(n6768), .ZN(n6794)
         );
  NOR4_X1 U7751 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), .A3(n6928), .A4(n6930), .ZN(n6776) );
  INV_X1 U7752 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n7027) );
  NOR4_X1 U7753 ( .A1(FLUSH_REG_SCAN_IN), .A2(n7025), .A3(n7027), .A4(n4835), 
        .ZN(n6775) );
  NOR4_X1 U7754 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(
        INSTQUEUE_REG_9__5__SCAN_IN), .A3(n3930), .A4(n6945), .ZN(n6774) );
  INV_X1 U7755 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6772) );
  AND4_X1 U7756 ( .A1(n6772), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .A3(
        EBX_REG_23__SCAN_IN), .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6773)
         );
  NAND4_X1 U7757 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(n6793)
         );
  NOR4_X1 U7758 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(
        INSTQUEUE_REG_12__5__SCAN_IN), .A3(DATAI_3_), .A4(n6881), .ZN(n6777)
         );
  NAND3_X1 U7759 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(M_IO_N_REG_SCAN_IN), 
        .A3(n6777), .ZN(n6778) );
  NOR3_X1 U7760 ( .A1(EBX_REG_7__SCAN_IN), .A2(UWORD_REG_5__SCAN_IN), .A3(
        n6778), .ZN(n6791) );
  NOR4_X1 U7761 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(ADDRESS_REG_5__SCAN_IN), .A3(DATAO_REG_14__SCAN_IN), .A4(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6790) );
  NAND4_X1 U7762 ( .A1(DATAI_21_), .A2(DATAWIDTH_REG_0__SCAN_IN), .A3(n6855), 
        .A4(n4659), .ZN(n6788) );
  NAND4_X1 U7763 ( .A1(EBX_REG_26__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(CODEFETCH_REG_SCAN_IN), .A4(n6868), .ZN(n6787) );
  INV_X1 U7764 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6780) );
  NAND4_X1 U7765 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .A3(DATAI_12_), .A4(
        DATAO_REG_17__SCAN_IN), .ZN(n6779) );
  NOR2_X1 U7766 ( .A1(n6780), .A2(n6779), .ZN(n6782) );
  INV_X1 U7767 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6781) );
  NAND4_X1 U7768 ( .A1(n6782), .A2(DATAI_26_), .A3(ADDRESS_REG_16__SCAN_IN), 
        .A4(n6781), .ZN(n6786) );
  NAND4_X1 U7769 ( .A1(n6784), .A2(n6783), .A3(INSTQUEUE_REG_9__3__SCAN_IN), 
        .A4(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6785) );
  NOR4_X1 U7770 ( .A1(n6788), .A2(n6787), .A3(n6786), .A4(n6785), .ZN(n6789)
         );
  NAND3_X1 U7771 ( .A1(n6791), .A2(n6790), .A3(n6789), .ZN(n6792) );
  NOR4_X1 U7772 ( .A1(n6795), .A2(n6794), .A3(n6793), .A4(n6792), .ZN(n6796)
         );
  NAND4_X1 U7773 ( .A1(n6799), .A2(n6798), .A3(n6797), .A4(n6796), .ZN(n7057)
         );
  AOI22_X1 U7774 ( .A1(n6802), .A2(keyinput40), .B1(n6801), .B2(keyinput96), 
        .ZN(n6800) );
  OAI221_X1 U7775 ( .B1(n6802), .B2(keyinput40), .C1(n6801), .C2(keyinput96), 
        .A(n6800), .ZN(n6814) );
  AOI22_X1 U7776 ( .A1(n6804), .A2(keyinput25), .B1(n5331), .B2(keyinput34), 
        .ZN(n6803) );
  OAI221_X1 U7777 ( .B1(n6804), .B2(keyinput25), .C1(n5331), .C2(keyinput34), 
        .A(n6803), .ZN(n6813) );
  INV_X1 U7778 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6806) );
  AOI22_X1 U7779 ( .A1(n6807), .A2(keyinput75), .B1(n6806), .B2(keyinput84), 
        .ZN(n6805) );
  OAI221_X1 U7780 ( .B1(n6807), .B2(keyinput75), .C1(n6806), .C2(keyinput84), 
        .A(n6805), .ZN(n6812) );
  INV_X1 U7781 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n6808) );
  XOR2_X1 U7782 ( .A(n6808), .B(keyinput44), .Z(n6810) );
  XNOR2_X1 U7783 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput73), .ZN(
        n6809) );
  NAND2_X1 U7784 ( .A1(n6810), .A2(n6809), .ZN(n6811) );
  NOR4_X1 U7785 ( .A1(n6814), .A2(n6813), .A3(n6812), .A4(n6811), .ZN(n6864)
         );
  INV_X1 U7786 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6816) );
  AOI22_X1 U7787 ( .A1(n6817), .A2(keyinput81), .B1(n6816), .B2(keyinput37), 
        .ZN(n6815) );
  OAI221_X1 U7788 ( .B1(n6817), .B2(keyinput81), .C1(n6816), .C2(keyinput37), 
        .A(n6815), .ZN(n6830) );
  INV_X1 U7789 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6820) );
  AOI22_X1 U7790 ( .A1(n6820), .A2(keyinput103), .B1(keyinput65), .B2(n6819), 
        .ZN(n6818) );
  OAI221_X1 U7791 ( .B1(n6820), .B2(keyinput103), .C1(n6819), .C2(keyinput65), 
        .A(n6818), .ZN(n6829) );
  AOI22_X1 U7792 ( .A1(n6823), .A2(keyinput95), .B1(keyinput12), .B2(n6822), 
        .ZN(n6821) );
  OAI221_X1 U7793 ( .B1(n6823), .B2(keyinput95), .C1(n6822), .C2(keyinput12), 
        .A(n6821), .ZN(n6828) );
  INV_X1 U7794 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6826) );
  INV_X1 U7795 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6825) );
  AOI22_X1 U7796 ( .A1(n6826), .A2(keyinput27), .B1(n6825), .B2(keyinput117), 
        .ZN(n6824) );
  OAI221_X1 U7797 ( .B1(n6826), .B2(keyinput27), .C1(n6825), .C2(keyinput117), 
        .A(n6824), .ZN(n6827) );
  NOR4_X1 U7798 ( .A1(n6830), .A2(n6829), .A3(n6828), .A4(n6827), .ZN(n6863)
         );
  AOI22_X1 U7799 ( .A1(n6832), .A2(keyinput123), .B1(keyinput83), .B2(n5324), 
        .ZN(n6831) );
  OAI221_X1 U7800 ( .B1(n6832), .B2(keyinput123), .C1(n5324), .C2(keyinput83), 
        .A(n6831), .ZN(n6844) );
  AOI22_X1 U7801 ( .A1(n6835), .A2(keyinput109), .B1(keyinput93), .B2(n6834), 
        .ZN(n6833) );
  OAI221_X1 U7802 ( .B1(n6835), .B2(keyinput109), .C1(n6834), .C2(keyinput93), 
        .A(n6833), .ZN(n6843) );
  AOI22_X1 U7803 ( .A1(n6838), .A2(keyinput11), .B1(n6837), .B2(keyinput66), 
        .ZN(n6836) );
  OAI221_X1 U7804 ( .B1(n6838), .B2(keyinput11), .C1(n6837), .C2(keyinput66), 
        .A(n6836), .ZN(n6842) );
  XNOR2_X1 U7805 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput98), .ZN(n6840) );
  XNOR2_X1 U7806 ( .A(keyinput42), .B(DATAI_7_), .ZN(n6839) );
  NAND2_X1 U7807 ( .A1(n6840), .A2(n6839), .ZN(n6841) );
  NOR4_X1 U7808 ( .A1(n6844), .A2(n6843), .A3(n6842), .A4(n6841), .ZN(n6862)
         );
  AOI22_X1 U7809 ( .A1(n6847), .A2(keyinput9), .B1(keyinput80), .B2(n6846), 
        .ZN(n6845) );
  OAI221_X1 U7810 ( .B1(n6847), .B2(keyinput9), .C1(n6846), .C2(keyinput80), 
        .A(n6845), .ZN(n6860) );
  AOI22_X1 U7811 ( .A1(n6850), .A2(keyinput43), .B1(n6849), .B2(keyinput77), 
        .ZN(n6848) );
  OAI221_X1 U7812 ( .B1(n6850), .B2(keyinput43), .C1(n6849), .C2(keyinput77), 
        .A(n6848), .ZN(n6859) );
  AOI22_X1 U7813 ( .A1(n6853), .A2(keyinput48), .B1(n6852), .B2(keyinput19), 
        .ZN(n6851) );
  OAI221_X1 U7814 ( .B1(n6853), .B2(keyinput48), .C1(n6852), .C2(keyinput19), 
        .A(n6851), .ZN(n6858) );
  INV_X1 U7815 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n6856) );
  AOI22_X1 U7816 ( .A1(n6856), .A2(keyinput124), .B1(n6855), .B2(keyinput23), 
        .ZN(n6854) );
  OAI221_X1 U7817 ( .B1(n6856), .B2(keyinput124), .C1(n6855), .C2(keyinput23), 
        .A(n6854), .ZN(n6857) );
  NOR4_X1 U7818 ( .A1(n6860), .A2(n6859), .A3(n6858), .A4(n6857), .ZN(n6861)
         );
  NAND4_X1 U7819 ( .A1(n6864), .A2(n6863), .A3(n6862), .A4(n6861), .ZN(n7055)
         );
  AOI22_X1 U7820 ( .A1(n6866), .A2(keyinput14), .B1(n4659), .B2(keyinput30), 
        .ZN(n6865) );
  OAI221_X1 U7821 ( .B1(n6866), .B2(keyinput14), .C1(n4659), .C2(keyinput30), 
        .A(n6865), .ZN(n6879) );
  INV_X1 U7822 ( .A(DATAI_21_), .ZN(n6869) );
  AOI22_X1 U7823 ( .A1(n6869), .A2(keyinput59), .B1(n6868), .B2(keyinput122), 
        .ZN(n6867) );
  OAI221_X1 U7824 ( .B1(n6869), .B2(keyinput59), .C1(n6868), .C2(keyinput122), 
        .A(n6867), .ZN(n6878) );
  AOI22_X1 U7825 ( .A1(n6872), .A2(keyinput118), .B1(keyinput6), .B2(n6871), 
        .ZN(n6870) );
  OAI221_X1 U7826 ( .B1(n6872), .B2(keyinput118), .C1(n6871), .C2(keyinput6), 
        .A(n6870), .ZN(n6877) );
  INV_X1 U7827 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6874) );
  AOI22_X1 U7828 ( .A1(n6875), .A2(keyinput18), .B1(keyinput91), .B2(n6874), 
        .ZN(n6873) );
  OAI221_X1 U7829 ( .B1(n6875), .B2(keyinput18), .C1(n6874), .C2(keyinput91), 
        .A(n6873), .ZN(n6876) );
  NOR4_X1 U7830 ( .A1(n6879), .A2(n6878), .A3(n6877), .A4(n6876), .ZN(n6925)
         );
  INV_X1 U7831 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n6882) );
  AOI22_X1 U7832 ( .A1(n6882), .A2(keyinput101), .B1(n6881), .B2(keyinput7), 
        .ZN(n6880) );
  OAI221_X1 U7833 ( .B1(n6882), .B2(keyinput101), .C1(n6881), .C2(keyinput7), 
        .A(n6880), .ZN(n6893) );
  INV_X1 U7834 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6884) );
  AOI22_X1 U7835 ( .A1(n6885), .A2(keyinput125), .B1(n6884), .B2(keyinput89), 
        .ZN(n6883) );
  OAI221_X1 U7836 ( .B1(n6885), .B2(keyinput125), .C1(n6884), .C2(keyinput89), 
        .A(n6883), .ZN(n6892) );
  INV_X1 U7837 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6886) );
  XOR2_X1 U7838 ( .A(n6886), .B(keyinput8), .Z(n6890) );
  XNOR2_X1 U7839 ( .A(keyinput74), .B(DATAI_3_), .ZN(n6889) );
  XNOR2_X1 U7840 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .B(keyinput47), .ZN(n6888)
         );
  XNOR2_X1 U7841 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .B(keyinput56), .ZN(n6887)
         );
  NAND4_X1 U7842 ( .A1(n6890), .A2(n6889), .A3(n6888), .A4(n6887), .ZN(n6891)
         );
  NOR3_X1 U7843 ( .A1(n6893), .A2(n6892), .A3(n6891), .ZN(n6924) );
  AOI22_X1 U7844 ( .A1(n6784), .A2(keyinput92), .B1(n6781), .B2(keyinput54), 
        .ZN(n6894) );
  OAI221_X1 U7845 ( .B1(n6784), .B2(keyinput92), .C1(n6781), .C2(keyinput54), 
        .A(n6894), .ZN(n6907) );
  INV_X1 U7846 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6896) );
  AOI22_X1 U7847 ( .A1(n6897), .A2(keyinput112), .B1(n6896), .B2(keyinput110), 
        .ZN(n6895) );
  OAI221_X1 U7848 ( .B1(n6897), .B2(keyinput112), .C1(n6896), .C2(keyinput110), 
        .A(n6895), .ZN(n6906) );
  AOI22_X1 U7849 ( .A1(n6900), .A2(keyinput126), .B1(keyinput41), .B2(n6899), 
        .ZN(n6898) );
  OAI221_X1 U7850 ( .B1(n6900), .B2(keyinput126), .C1(n6899), .C2(keyinput41), 
        .A(n6898), .ZN(n6905) );
  INV_X1 U7851 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6902) );
  AOI22_X1 U7852 ( .A1(n6903), .A2(keyinput90), .B1(n6902), .B2(keyinput22), 
        .ZN(n6901) );
  OAI221_X1 U7853 ( .B1(n6903), .B2(keyinput90), .C1(n6902), .C2(keyinput22), 
        .A(n6901), .ZN(n6904) );
  NOR4_X1 U7854 ( .A1(n6907), .A2(n6906), .A3(n6905), .A4(n6904), .ZN(n6923)
         );
  INV_X1 U7855 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U7856 ( .A1(n6909), .A2(keyinput20), .B1(keyinput119), .B2(n4658), 
        .ZN(n6908) );
  OAI221_X1 U7857 ( .B1(n6909), .B2(keyinput20), .C1(n4658), .C2(keyinput119), 
        .A(n6908), .ZN(n6921) );
  INV_X1 U7858 ( .A(DATAI_26_), .ZN(n6912) );
  AOI22_X1 U7859 ( .A1(n6912), .A2(keyinput39), .B1(keyinput1), .B2(n6911), 
        .ZN(n6910) );
  OAI221_X1 U7860 ( .B1(n6912), .B2(keyinput39), .C1(n6911), .C2(keyinput1), 
        .A(n6910), .ZN(n6920) );
  INV_X1 U7861 ( .A(DATAI_12_), .ZN(n6915) );
  INV_X1 U7862 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6914) );
  AOI22_X1 U7863 ( .A1(n6915), .A2(keyinput97), .B1(n6914), .B2(keyinput50), 
        .ZN(n6913) );
  OAI221_X1 U7864 ( .B1(n6915), .B2(keyinput97), .C1(n6914), .C2(keyinput50), 
        .A(n6913), .ZN(n6919) );
  XNOR2_X1 U7865 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(keyinput114), .ZN(
        n6917) );
  XNOR2_X1 U7866 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .B(keyinput70), .ZN(n6916)
         );
  NAND2_X1 U7867 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  NOR4_X1 U7868 ( .A1(n6921), .A2(n6920), .A3(n6919), .A4(n6918), .ZN(n6922)
         );
  NAND4_X1 U7869 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(n7054)
         );
  AOI22_X1 U7870 ( .A1(n6928), .A2(keyinput63), .B1(keyinput58), .B2(n6927), 
        .ZN(n6926) );
  OAI221_X1 U7871 ( .B1(n6928), .B2(keyinput63), .C1(n6927), .C2(keyinput58), 
        .A(n6926), .ZN(n6940) );
  AOI22_X1 U7872 ( .A1(n6772), .A2(keyinput72), .B1(keyinput3), .B2(n6930), 
        .ZN(n6929) );
  OAI221_X1 U7873 ( .B1(n6772), .B2(keyinput72), .C1(n6930), .C2(keyinput3), 
        .A(n6929), .ZN(n6939) );
  AOI22_X1 U7874 ( .A1(n6933), .A2(keyinput104), .B1(keyinput113), .B2(n6932), 
        .ZN(n6931) );
  OAI221_X1 U7875 ( .B1(n6933), .B2(keyinput104), .C1(n6932), .C2(keyinput113), 
        .A(n6931), .ZN(n6938) );
  AOI22_X1 U7876 ( .A1(n6936), .A2(keyinput2), .B1(n6935), .B2(keyinput38), 
        .ZN(n6934) );
  OAI221_X1 U7877 ( .B1(n6936), .B2(keyinput2), .C1(n6935), .C2(keyinput38), 
        .A(n6934), .ZN(n6937) );
  NOR4_X1 U7878 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n6986)
         );
  INV_X1 U7879 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6942) );
  AOI22_X1 U7880 ( .A1(n6943), .A2(keyinput29), .B1(n6942), .B2(keyinput94), 
        .ZN(n6941) );
  OAI221_X1 U7881 ( .B1(n6943), .B2(keyinput29), .C1(n6942), .C2(keyinput94), 
        .A(n6941), .ZN(n6953) );
  AOI22_X1 U7882 ( .A1(n6945), .A2(keyinput46), .B1(n3780), .B2(keyinput64), 
        .ZN(n6944) );
  OAI221_X1 U7883 ( .B1(n6945), .B2(keyinput46), .C1(n3780), .C2(keyinput64), 
        .A(n6944), .ZN(n6952) );
  INV_X1 U7884 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6947) );
  AOI22_X1 U7885 ( .A1(n3930), .A2(keyinput99), .B1(n6947), .B2(keyinput69), 
        .ZN(n6946) );
  OAI221_X1 U7886 ( .B1(n3930), .B2(keyinput99), .C1(n6947), .C2(keyinput69), 
        .A(n6946), .ZN(n6951) );
  XNOR2_X1 U7887 ( .A(EBX_REG_23__SCAN_IN), .B(keyinput53), .ZN(n6949) );
  XNOR2_X1 U7888 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .B(keyinput105), .ZN(n6948) );
  NAND2_X1 U7889 ( .A1(n6949), .A2(n6948), .ZN(n6950) );
  NOR4_X1 U7890 ( .A1(n6953), .A2(n6952), .A3(n6951), .A4(n6950), .ZN(n6985)
         );
  INV_X1 U7891 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6956) );
  AOI22_X1 U7892 ( .A1(n6956), .A2(keyinput121), .B1(keyinput60), .B2(n6955), 
        .ZN(n6954) );
  OAI221_X1 U7893 ( .B1(n6956), .B2(keyinput121), .C1(n6955), .C2(keyinput60), 
        .A(n6954), .ZN(n6969) );
  AOI22_X1 U7894 ( .A1(n6959), .A2(keyinput51), .B1(keyinput32), .B2(n6958), 
        .ZN(n6957) );
  OAI221_X1 U7895 ( .B1(n6959), .B2(keyinput51), .C1(n6958), .C2(keyinput32), 
        .A(n6957), .ZN(n6968) );
  AOI22_X1 U7896 ( .A1(n6962), .A2(keyinput33), .B1(n6961), .B2(keyinput45), 
        .ZN(n6960) );
  OAI221_X1 U7897 ( .B1(n6962), .B2(keyinput33), .C1(n6961), .C2(keyinput45), 
        .A(n6960), .ZN(n6967) );
  AOI22_X1 U7898 ( .A1(n6965), .A2(keyinput82), .B1(keyinput120), .B2(n6964), 
        .ZN(n6963) );
  OAI221_X1 U7899 ( .B1(n6965), .B2(keyinput82), .C1(n6964), .C2(keyinput120), 
        .A(n6963), .ZN(n6966) );
  NOR4_X1 U7900 ( .A1(n6969), .A2(n6968), .A3(n6967), .A4(n6966), .ZN(n6984)
         );
  INV_X1 U7901 ( .A(DATAI_18_), .ZN(n6971) );
  AOI22_X1 U7902 ( .A1(n6971), .A2(keyinput62), .B1(n6748), .B2(keyinput0), 
        .ZN(n6970) );
  OAI221_X1 U7903 ( .B1(n6971), .B2(keyinput62), .C1(n6748), .C2(keyinput0), 
        .A(n6970), .ZN(n6982) );
  AOI22_X1 U7904 ( .A1(n3912), .A2(keyinput61), .B1(n6973), .B2(keyinput71), 
        .ZN(n6972) );
  OAI221_X1 U7905 ( .B1(n3912), .B2(keyinput61), .C1(n6973), .C2(keyinput71), 
        .A(n6972), .ZN(n6981) );
  AOI22_X1 U7906 ( .A1(n6975), .A2(keyinput116), .B1(keyinput16), .B2(n4401), 
        .ZN(n6974) );
  OAI221_X1 U7907 ( .B1(n6975), .B2(keyinput116), .C1(n4401), .C2(keyinput16), 
        .A(n6974), .ZN(n6980) );
  AOI22_X1 U7908 ( .A1(n6978), .A2(keyinput115), .B1(keyinput17), .B2(n6977), 
        .ZN(n6976) );
  OAI221_X1 U7909 ( .B1(n6978), .B2(keyinput115), .C1(n6977), .C2(keyinput17), 
        .A(n6976), .ZN(n6979) );
  NOR4_X1 U7910 ( .A1(n6982), .A2(n6981), .A3(n6980), .A4(n6979), .ZN(n6983)
         );
  NAND4_X1 U7911 ( .A1(n6986), .A2(n6985), .A3(n6984), .A4(n6983), .ZN(n7053)
         );
  AOI22_X1 U7912 ( .A1(n6989), .A2(keyinput85), .B1(keyinput57), .B2(n6988), 
        .ZN(n6987) );
  OAI221_X1 U7913 ( .B1(n6989), .B2(keyinput85), .C1(n6988), .C2(keyinput57), 
        .A(n6987), .ZN(n7001) );
  INV_X1 U7914 ( .A(DATAI_27_), .ZN(n6991) );
  AOI22_X1 U7915 ( .A1(n6991), .A2(keyinput31), .B1(keyinput55), .B2(n4594), 
        .ZN(n6990) );
  OAI221_X1 U7916 ( .B1(n6991), .B2(keyinput31), .C1(n4594), .C2(keyinput55), 
        .A(n6990), .ZN(n7000) );
  INV_X1 U7917 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6993) );
  AOI22_X1 U7918 ( .A1(n6994), .A2(keyinput36), .B1(n6993), .B2(keyinput52), 
        .ZN(n6992) );
  OAI221_X1 U7919 ( .B1(n6994), .B2(keyinput36), .C1(n6993), .C2(keyinput52), 
        .A(n6992), .ZN(n6999) );
  AOI22_X1 U7920 ( .A1(n6997), .A2(keyinput4), .B1(keyinput100), .B2(n6996), 
        .ZN(n6995) );
  OAI221_X1 U7921 ( .B1(n6997), .B2(keyinput4), .C1(n6996), .C2(keyinput100), 
        .A(n6995), .ZN(n6998) );
  NOR4_X1 U7922 ( .A1(n7001), .A2(n7000), .A3(n6999), .A4(n6998), .ZN(n7051)
         );
  INV_X1 U7923 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n7003) );
  NAND2_X1 U7924 ( .A1(n7003), .A2(keyinput76), .ZN(n7002) );
  OAI221_X1 U7925 ( .B1(n7004), .B2(keyinput15), .C1(n7003), .C2(keyinput76), 
        .A(n7002), .ZN(n7017) );
  INV_X1 U7926 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n7006) );
  AOI22_X1 U7927 ( .A1(n7007), .A2(keyinput35), .B1(n7006), .B2(keyinput102), 
        .ZN(n7005) );
  OAI221_X1 U7928 ( .B1(n7007), .B2(keyinput35), .C1(n7006), .C2(keyinput102), 
        .A(n7005), .ZN(n7016) );
  AOI22_X1 U7929 ( .A1(n7010), .A2(keyinput28), .B1(n7009), .B2(keyinput87), 
        .ZN(n7008) );
  OAI221_X1 U7930 ( .B1(n7010), .B2(keyinput28), .C1(n7009), .C2(keyinput87), 
        .A(n7008), .ZN(n7015) );
  AOI22_X1 U7931 ( .A1(n7013), .A2(keyinput79), .B1(keyinput67), .B2(n7012), 
        .ZN(n7011) );
  OAI221_X1 U7932 ( .B1(n7013), .B2(keyinput79), .C1(n7012), .C2(keyinput67), 
        .A(n7011), .ZN(n7014) );
  NOR4_X1 U7933 ( .A1(n7017), .A2(n7016), .A3(n7015), .A4(n7014), .ZN(n7050)
         );
  AOI22_X1 U7934 ( .A1(n7020), .A2(keyinput107), .B1(keyinput49), .B2(n7019), 
        .ZN(n7018) );
  OAI221_X1 U7935 ( .B1(n7020), .B2(keyinput107), .C1(n7019), .C2(keyinput49), 
        .A(n7018), .ZN(n7032) );
  AOI22_X1 U7936 ( .A1(n7023), .A2(keyinput24), .B1(n7022), .B2(keyinput86), 
        .ZN(n7021) );
  OAI221_X1 U7937 ( .B1(n7023), .B2(keyinput24), .C1(n7022), .C2(keyinput86), 
        .A(n7021), .ZN(n7031) );
  AOI22_X1 U7938 ( .A1(n7025), .A2(keyinput10), .B1(keyinput88), .B2(n4835), 
        .ZN(n7024) );
  OAI221_X1 U7939 ( .B1(n7025), .B2(keyinput10), .C1(n4835), .C2(keyinput88), 
        .A(n7024), .ZN(n7030) );
  AOI22_X1 U7940 ( .A1(n7028), .A2(keyinput108), .B1(n7027), .B2(keyinput78), 
        .ZN(n7026) );
  OAI221_X1 U7941 ( .B1(n7028), .B2(keyinput108), .C1(n7027), .C2(keyinput78), 
        .A(n7026), .ZN(n7029) );
  NOR4_X1 U7942 ( .A1(n7032), .A2(n7031), .A3(n7030), .A4(n7029), .ZN(n7049)
         );
  INV_X1 U7943 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n7035) );
  AOI22_X1 U7944 ( .A1(n7035), .A2(keyinput127), .B1(n7034), .B2(keyinput111), 
        .ZN(n7033) );
  OAI221_X1 U7945 ( .B1(n7035), .B2(keyinput127), .C1(n7034), .C2(keyinput111), 
        .A(n7033), .ZN(n7047) );
  AOI22_X1 U7946 ( .A1(n7038), .A2(keyinput5), .B1(keyinput21), .B2(n7037), 
        .ZN(n7036) );
  OAI221_X1 U7947 ( .B1(n7038), .B2(keyinput5), .C1(n7037), .C2(keyinput21), 
        .A(n7036), .ZN(n7046) );
  AOI22_X1 U7948 ( .A1(n4596), .A2(keyinput13), .B1(n7040), .B2(keyinput26), 
        .ZN(n7039) );
  OAI221_X1 U7949 ( .B1(n4596), .B2(keyinput13), .C1(n7040), .C2(keyinput26), 
        .A(n7039), .ZN(n7045) );
  AOI22_X1 U7950 ( .A1(n7043), .A2(keyinput68), .B1(keyinput106), .B2(n7042), 
        .ZN(n7041) );
  OAI221_X1 U7951 ( .B1(n7043), .B2(keyinput68), .C1(n7042), .C2(keyinput106), 
        .A(n7041), .ZN(n7044) );
  NOR4_X1 U7952 ( .A1(n7047), .A2(n7046), .A3(n7045), .A4(n7044), .ZN(n7048)
         );
  NAND4_X1 U7953 ( .A1(n7051), .A2(n7050), .A3(n7049), .A4(n7048), .ZN(n7052)
         );
  NOR4_X1 U7954 ( .A1(n7055), .A2(n7054), .A3(n7053), .A4(n7052), .ZN(n7056)
         );
  OAI221_X1 U7955 ( .B1(n7058), .B2(BE_N_REG_3__SCAN_IN), .C1(n7058), .C2(
        n7057), .A(n7056), .ZN(n7059) );
  XOR2_X1 U7956 ( .A(n7060), .B(n7059), .Z(U2902) );
  CLKBUF_X1 U3557 ( .A(n3468), .Z(n3447) );
  CLKBUF_X1 U3567 ( .A(n3385), .Z(n3678) );
  CLKBUF_X2 U3570 ( .A(n3388), .Z(n3729) );
  CLKBUF_X1 U3624 ( .A(n4805), .Z(n6227) );
  CLKBUF_X1 U3976 ( .A(n4457), .Z(n5911) );
  CLKBUF_X1 U4478 ( .A(n3893), .Z(n4623) );
endmodule

