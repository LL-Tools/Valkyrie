

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput127,
         keyinput126, keyinput125, keyinput124, keyinput123, keyinput122,
         keyinput121, keyinput120, keyinput119, keyinput118, keyinput117,
         keyinput116, keyinput115, keyinput114, keyinput113, keyinput112,
         keyinput111, keyinput110, keyinput109, keyinput108, keyinput107,
         keyinput106, keyinput105, keyinput104, keyinput103, keyinput102,
         keyinput101, keyinput100, keyinput99, keyinput98, keyinput97,
         keyinput96, keyinput95, keyinput94, keyinput93, keyinput92,
         keyinput91, keyinput90, keyinput89, keyinput88, keyinput87,
         keyinput86, keyinput85, keyinput84, keyinput83, keyinput82,
         keyinput81, keyinput80, keyinput79, keyinput78, keyinput77,
         keyinput76, keyinput75, keyinput74, keyinput73, keyinput72,
         keyinput71, keyinput70, keyinput69, keyinput68, keyinput67,
         keyinput66, keyinput65, keyinput64, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11452, n11453,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343;

  OAI21_X1 U7264 ( .B1(n12060), .B2(n6657), .A(n7084), .ZN(n7083) );
  NOR2_X1 U7265 ( .A1(n10485), .A2(n10473), .ZN(n10709) );
  INV_X2 U7266 ( .A(n10803), .ZN(n6520) );
  CLKBUF_X2 U7267 ( .A(n8563), .Z(n6518) );
  CLKBUF_X2 U7268 ( .A(n8537), .Z(n9078) );
  INV_X1 U7269 ( .A(n10495), .ZN(n11861) );
  NOR2_X1 U7270 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n8414) );
  AND2_X1 U7271 ( .A1(n9324), .A2(n9323), .ZN(n9536) );
  INV_X1 U7273 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9164) );
  INV_X1 U7274 ( .A(n12095), .ZN(n6517) );
  INV_X2 U7275 ( .A(n12973), .ZN(n12997) );
  NAND2_X1 U7276 ( .A1(n9595), .A2(n9591), .ZN(n13739) );
  OAI21_X1 U7277 ( .B1(n12354), .B2(n11633), .A(n10110), .ZN(n9985) );
  INV_X1 U7278 ( .A(n8814), .ZN(n11764) );
  AND2_X1 U7279 ( .A1(n12309), .A2(n12323), .ZN(n12331) );
  NAND2_X1 U7280 ( .A1(n12292), .A2(n12291), .ZN(n12293) );
  INV_X1 U7281 ( .A(n11736), .ZN(n11755) );
  INV_X1 U7282 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6812) );
  NAND2_X1 U7283 ( .A1(n13201), .A2(n13172), .ZN(n13218) );
  CLKBUF_X2 U7285 ( .A(n10605), .Z(n13697) );
  NAND2_X1 U7286 ( .A1(n10405), .A2(n10374), .ZN(n10021) );
  OAI22_X1 U7287 ( .A1(n12168), .A2(n12023), .B1(n12494), .B2(n12166), .ZN(
        n12084) );
  BUF_X1 U7288 ( .A(n8534), .Z(n6527) );
  OR2_X1 U7290 ( .A1(n14886), .A2(n12210), .ZN(n7043) );
  NAND2_X1 U7291 ( .A1(n11751), .A2(n11750), .ZN(n12373) );
  AND2_X1 U7292 ( .A1(n6516), .A2(n7527), .ZN(n8430) );
  OAI21_X1 U7293 ( .B1(n8805), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8807) );
  OR2_X1 U7294 ( .A1(n8727), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8755) );
  INV_X2 U7295 ( .A(n9650), .ZN(n12959) );
  NAND2_X1 U7296 ( .A1(n8356), .A2(n10018), .ZN(n10009) );
  NOR2_X1 U7297 ( .A1(n14864), .A2(n8686), .ZN(n14863) );
  AOI21_X1 U7298 ( .B1(n12336), .B2(n12335), .A(n12334), .ZN(n12359) );
  INV_X1 U7299 ( .A(n13858), .ZN(n10405) );
  INV_X1 U7300 ( .A(n8005), .ZN(n8346) );
  XNOR2_X1 U7302 ( .A(n13174), .B(n13202), .ZN(n13444) );
  INV_X1 U7303 ( .A(n13049), .ZN(n12968) );
  INV_X1 U7304 ( .A(n10374), .ZN(n14585) );
  NAND4_X1 U7305 ( .A1(n7811), .A2(n7810), .A3(n7809), .A4(n7808), .ZN(n13854)
         );
  AND4_X2 U7306 ( .A1(n7097), .A2(n7098), .A3(n7524), .A4(n7523), .ZN(n6516)
         );
  NAND2_X4 U7307 ( .A1(n7759), .A2(n9343), .ZN(n8005) );
  AND2_X2 U7309 ( .A1(n6921), .A2(n9524), .ZN(n9533) );
  NAND2_X2 U7310 ( .A1(n6982), .A2(n14537), .ZN(n7651) );
  NAND2_X2 U7311 ( .A1(n8490), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8488) );
  AND2_X2 U7312 ( .A1(n12786), .A2(n11973), .ZN(n11985) );
  NAND2_X2 U7313 ( .A1(n12734), .A2(n7250), .ZN(n12786) );
  XNOR2_X2 U7314 ( .A(n7673), .B(n14292), .ZN(n7678) );
  OR2_X1 U7315 ( .A1(n12206), .A2(n10322), .ZN(n11650) );
  XNOR2_X1 U7316 ( .A(n13074), .B(n6534), .ZN(n13006) );
  OAI21_X2 U7317 ( .B1(n13392), .B2(n7116), .A(n7114), .ZN(n13335) );
  OAI222_X1 U7318 ( .A1(n13580), .A2(n15216), .B1(P2_U3088), .B2(n9334), .C1(
        n13578), .C2(n11188), .ZN(P2_U3306) );
  OR2_X4 U7319 ( .A1(n9334), .A2(n9333), .ZN(n6571) );
  NAND2_X2 U7320 ( .A1(n8516), .A2(n8515), .ZN(n9677) );
  OR2_X2 U7321 ( .A1(n8559), .A2(n8444), .ZN(n8446) );
  NOR2_X1 U7322 ( .A1(n15342), .A2(n15343), .ZN(n15341) );
  OAI22_X2 U7323 ( .A1(n14098), .A2(n14097), .B1(n14236), .B2(n13844), .ZN(
        n14088) );
  NAND2_X2 U7324 ( .A1(n14125), .A2(n7532), .ZN(n14098) );
  NAND2_X1 U7325 ( .A1(n8348), .A2(n11295), .ZN(n9511) );
  NAND2_X1 U7326 ( .A1(n8435), .A2(n12686), .ZN(n8563) );
  OAI222_X1 U7327 ( .A1(P3_U3151), .A2(n8434), .B1(n12698), .B2(n12689), .C1(
        n12694), .C2(n12688), .ZN(P3_U3266) );
  OAI22_X2 U7328 ( .A1(n9871), .A2(n6528), .B1(n9883), .B2(n9349), .ZN(n9356)
         );
  OAI211_X2 U7329 ( .C1(n9142), .C2(n9078), .A(n8574), .B(n8573), .ZN(n10322)
         );
  OR2_X2 U7330 ( .A1(n11775), .A2(SI_4_), .ZN(n8573) );
  NOR2_X2 U7331 ( .A1(n6863), .A2(n6637), .ZN(n12414) );
  XNOR2_X2 U7332 ( .A(n6927), .B(n9217), .ZN(n9334) );
  INV_X2 U7333 ( .A(n9216), .ZN(n6927) );
  XNOR2_X2 U7334 ( .A(n12262), .B(n12277), .ZN(n12244) );
  OAI22_X2 U7335 ( .A1(n8086), .A2(n6729), .B1(n9777), .B2(n8084), .ZN(n8136)
         );
  NAND2_X2 U7336 ( .A1(n8077), .A2(n8076), .ZN(n8086) );
  OR2_X1 U7337 ( .A1(n14796), .A2(n9333), .ZN(n6519) );
  OAI21_X2 U7338 ( .B1(n7641), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n14322), .ZN(
        n14328) );
  NAND2_X1 U7339 ( .A1(n6767), .A2(n7542), .ZN(n12381) );
  CLKBUF_X1 U7340 ( .A(n14050), .Z(n6836) );
  NOR2_X1 U7341 ( .A1(n7541), .A2(n6733), .ZN(n6732) );
  NAND2_X1 U7342 ( .A1(n6797), .A2(n12940), .ZN(n13141) );
  NAND2_X1 U7343 ( .A1(n13187), .A2(n13186), .ZN(n13337) );
  OAI21_X1 U7344 ( .B1(n6763), .B2(n6762), .A(n6760), .ZN(n8724) );
  INV_X1 U7345 ( .A(n11189), .ZN(n11101) );
  NOR2_X1 U7346 ( .A1(n13601), .A2(n13847), .ZN(n11196) );
  CLKBUF_X2 U7348 ( .A(P2_U3947), .Z(n6523) );
  INV_X2 U7349 ( .A(n14945), .ZN(n10425) );
  NAND2_X1 U7350 ( .A1(n9642), .A2(n6742), .ZN(n12820) );
  INV_X1 U7351 ( .A(n10415), .ZN(n7725) );
  INV_X1 U7352 ( .A(n6823), .ZN(n8522) );
  INV_X2 U7353 ( .A(n8298), .ZN(n8180) );
  BUF_X2 U7354 ( .A(n11764), .Z(n6532) );
  NAND2_X2 U7355 ( .A1(n9602), .A2(n10973), .ZN(n9590) );
  CLKBUF_X2 U7356 ( .A(n7771), .Z(n8298) );
  NAND2_X1 U7357 ( .A1(n7759), .A2(n6967), .ZN(n8002) );
  BUF_X4 U7358 ( .A(n12965), .Z(n6521) );
  OR2_X1 U7359 ( .A1(n8489), .A2(n7074), .ZN(n7073) );
  XNOR2_X1 U7360 ( .A(n7692), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8348) );
  INV_X1 U7361 ( .A(n11295), .ZN(n10792) );
  BUF_X1 U7362 ( .A(n7677), .Z(n14299) );
  NOR2_X1 U7363 ( .A1(n7690), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n8389) );
  XNOR2_X1 U7364 ( .A(n7613), .B(n6839), .ZN(n7616) );
  NAND4_X1 U7365 ( .A1(n9084), .A2(n8583), .A3(n8415), .A4(n8414), .ZN(n8604)
         );
  AND2_X2 U7366 ( .A1(n6811), .A2(n6812), .ZN(n9084) );
  INV_X1 U7367 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8429) );
  NOR2_X1 U7368 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8417) );
  INV_X1 U7369 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6811) );
  INV_X1 U7370 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8910) );
  NOR2_X1 U7371 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8422) );
  NOR2_X1 U7372 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8415) );
  OAI21_X1 U7373 ( .B1(n8991), .B2(n15029), .A(n9003), .ZN(n9004) );
  OAI21_X1 U7374 ( .B1(n6696), .B2(n6759), .A(n7363), .ZN(n8387) );
  AND2_X1 U7375 ( .A1(n6734), .A2(n6732), .ZN(n13443) );
  NOR2_X1 U7376 ( .A1(n12550), .A2(n6594), .ZN(n7040) );
  OAI21_X1 U7377 ( .B1(n6750), .B2(n6749), .A(n7341), .ZN(n8266) );
  AND2_X1 U7378 ( .A1(n11832), .A2(n8946), .ZN(n6810) );
  AND2_X1 U7379 ( .A1(n11929), .A2(n7246), .ZN(n7245) );
  OR2_X1 U7380 ( .A1(n6589), .A2(n12385), .ZN(n12555) );
  NAND2_X1 U7381 ( .A1(n6913), .A2(n11928), .ZN(n11929) );
  AND2_X1 U7382 ( .A1(n7034), .A2(n7035), .ZN(n7033) );
  OR2_X1 U7383 ( .A1(n13036), .A2(n12945), .ZN(n12985) );
  OR4_X1 U7384 ( .A1(n13036), .A2(n13202), .A3(n13035), .A4(n13034), .ZN(
        n13037) );
  OR2_X1 U7385 ( .A1(n12159), .A2(n12444), .ZN(n12157) );
  NAND2_X1 U7386 ( .A1(n7023), .A2(n7021), .ZN(n12441) );
  NAND2_X1 U7387 ( .A1(n12478), .A2(n7027), .ZN(n7023) );
  AND2_X1 U7388 ( .A1(n13242), .A2(n7233), .ZN(n13209) );
  NAND2_X1 U7389 ( .A1(n13337), .A2(n13338), .ZN(n13336) );
  NAND2_X1 U7390 ( .A1(n12726), .A2(n11898), .ZN(n11912) );
  OAI21_X1 U7391 ( .B1(n12486), .B2(n7515), .A(n7512), .ZN(n12440) );
  CLKBUF_X1 U7392 ( .A(n7417), .Z(n6862) );
  NAND2_X1 U7393 ( .A1(n6915), .A2(n6914), .ZN(n12726) );
  AOI22_X1 U7394 ( .A1(n14297), .A2(n6539), .B1(n8346), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n14171) );
  NOR2_X1 U7395 ( .A1(n14029), .A2(n14195), .ZN(n14011) );
  NAND2_X1 U7396 ( .A1(n11471), .A2(n7418), .ZN(n7417) );
  XNOR2_X1 U7397 ( .A(n8345), .B(n8344), .ZN(n14297) );
  NAND2_X1 U7398 ( .A1(n12778), .A2(n6916), .ZN(n6915) );
  OAI21_X1 U7399 ( .B1(n8342), .B2(n8341), .A(n8340), .ZN(n8345) );
  OAI21_X1 U7400 ( .B1(n12504), .B2(n8935), .A(n11724), .ZN(n12484) );
  NAND2_X1 U7401 ( .A1(n8327), .A2(n8326), .ZN(n8342) );
  NAND2_X1 U7402 ( .A1(n8327), .A2(n8311), .ZN(n13568) );
  NAND2_X1 U7403 ( .A1(n8868), .A2(n8867), .ZN(n12047) );
  OR2_X1 U7404 ( .A1(n8310), .A2(n8309), .ZN(n8311) );
  NAND2_X1 U7405 ( .A1(n11413), .A2(n6792), .ZN(n11459) );
  AOI21_X1 U7406 ( .B1(n6916), .B2(n6918), .A(n6627), .ZN(n6914) );
  NAND2_X1 U7407 ( .A1(n6801), .A2(n6800), .ZN(n8305) );
  NAND2_X1 U7408 ( .A1(n8264), .A2(n8263), .ZN(n14195) );
  AOI21_X1 U7409 ( .B1(n6890), .B2(n6893), .A(n6623), .ZN(n6889) );
  NAND2_X1 U7410 ( .A1(n8191), .A2(n8190), .ZN(n14074) );
  OAI21_X1 U7411 ( .B1(n8286), .B2(n8285), .A(n8284), .ZN(n8291) );
  NAND2_X1 U7412 ( .A1(n8738), .A2(n8737), .ZN(n11509) );
  NAND2_X1 U7413 ( .A1(n11135), .A2(n11134), .ZN(n11138) );
  AND2_X1 U7414 ( .A1(n14307), .A2(n7759), .ZN(n14228) );
  XNOR2_X1 U7415 ( .A(n8189), .B(n8188), .ZN(n11914) );
  NAND2_X1 U7416 ( .A1(n11901), .A2(n11900), .ZN(n13482) );
  NAND2_X1 U7417 ( .A1(n11322), .A2(n11691), .ZN(n14365) );
  NAND2_X1 U7418 ( .A1(n8113), .A2(n8112), .ZN(n14249) );
  NAND2_X1 U7419 ( .A1(n7063), .A2(n6606), .ZN(n7062) );
  OAI21_X1 U7420 ( .B1(n10806), .B2(n7141), .A(n7138), .ZN(n10998) );
  AOI21_X1 U7421 ( .B1(n7392), .B2(n7389), .A(n6593), .ZN(n7388) );
  NAND2_X1 U7422 ( .A1(n11243), .A2(n11242), .ZN(n11244) );
  NAND2_X1 U7423 ( .A1(n8138), .A2(n8137), .ZN(n14244) );
  NAND2_X1 U7424 ( .A1(n11871), .A2(n11870), .ZN(n13493) );
  XNOR2_X1 U7425 ( .A(n8111), .B(n8110), .ZN(n11860) );
  NAND2_X1 U7426 ( .A1(n10807), .A2(n13017), .ZN(n10806) );
  NAND2_X1 U7427 ( .A1(n8028), .A2(n8027), .ZN(n13622) );
  NAND2_X1 U7428 ( .A1(n8092), .A2(n8091), .ZN(n14254) );
  NAND2_X1 U7429 ( .A1(n8008), .A2(n8007), .ZN(n14436) );
  OAI21_X1 U7430 ( .B1(n8173), .B2(n8172), .A(n8171), .ZN(n8205) );
  NAND2_X1 U7431 ( .A1(n11379), .A2(n11378), .ZN(n13521) );
  OR2_X1 U7432 ( .A1(n11048), .A2(n8932), .ZN(n8933) );
  INV_X1 U7433 ( .A(n13208), .ZN(n6733) );
  OR2_X1 U7434 ( .A1(n11125), .A2(n11124), .ZN(n11242) );
  NAND2_X1 U7435 ( .A1(n8478), .A2(n8477), .ZN(n8840) );
  OR2_X1 U7436 ( .A1(n8000), .A2(n8050), .ZN(n8020) );
  NAND2_X1 U7437 ( .A1(n10889), .A2(n10888), .ZN(n12880) );
  NAND2_X1 U7438 ( .A1(n7962), .A2(n7961), .ZN(n13601) );
  NAND2_X1 U7439 ( .A1(n9966), .A2(n9965), .ZN(n10059) );
  NAND2_X1 U7440 ( .A1(n10750), .A2(n10749), .ZN(n14844) );
  NAND2_X1 U7441 ( .A1(n6832), .A2(SI_14_), .ZN(n8019) );
  NAND2_X1 U7442 ( .A1(n7925), .A2(n7924), .ZN(n11345) );
  NAND2_X1 U7443 ( .A1(n7988), .A2(n7987), .ZN(n13610) );
  AND2_X1 U7444 ( .A1(n7044), .A2(n6635), .ZN(n10135) );
  OR2_X1 U7445 ( .A1(n10148), .A2(n10149), .ZN(n6678) );
  NAND2_X1 U7446 ( .A1(n10499), .A2(n10498), .ZN(n13424) );
  NAND2_X1 U7447 ( .A1(n7902), .A2(n7901), .ZN(n14616) );
  NOR2_X1 U7448 ( .A1(n9646), .A2(n9645), .ZN(n9740) );
  AOI21_X1 U7449 ( .B1(n14929), .B2(n8924), .A(n8552), .ZN(n10422) );
  NAND2_X1 U7450 ( .A1(n7834), .A2(n7833), .ZN(n10612) );
  NAND2_X2 U7451 ( .A1(n9917), .A2(n14803), .ZN(n14809) );
  NAND2_X1 U7452 ( .A1(n7857), .A2(n7856), .ZN(n10689) );
  NAND2_X1 U7453 ( .A1(n7877), .A2(n7894), .ZN(n10276) );
  NAND2_X1 U7454 ( .A1(n7804), .A2(n7803), .ZN(n10579) );
  NAND2_X1 U7455 ( .A1(n8465), .A2(n8464), .ZN(n8726) );
  NOR2_X1 U7456 ( .A1(n9096), .A2(n9095), .ZN(n10044) );
  AND2_X1 U7457 ( .A1(n7057), .A2(n7056), .ZN(n9076) );
  AND2_X1 U7458 ( .A1(n6720), .A2(n6719), .ZN(n7852) );
  NAND2_X1 U7459 ( .A1(n7052), .A2(n7050), .ZN(n7057) );
  NAND2_X1 U7460 ( .A1(n15326), .A2(n7625), .ZN(n7627) );
  NAND2_X1 U7461 ( .A1(n7725), .A2(n7724), .ZN(n10018) );
  AND2_X1 U7462 ( .A1(n7053), .A2(n6563), .ZN(n7050) );
  INV_X2 U7463 ( .A(n12820), .ZN(n6522) );
  OAI211_X1 U7464 ( .C1(n9136), .C2(n9078), .A(n8550), .B(n8549), .ZN(n14924)
         );
  NAND2_X2 U7465 ( .A1(n6669), .A2(n6878), .ZN(n13740) );
  NAND3_X1 U7466 ( .A1(n8512), .A2(n7540), .A3(n8513), .ZN(n6823) );
  OAI211_X1 U7467 ( .C1(n7759), .C2(n13884), .A(n7750), .B(n7749), .ZN(n10374)
         );
  NAND2_X1 U7468 ( .A1(n6679), .A2(n9834), .ZN(n9839) );
  NAND4_X1 U7469 ( .A1(n8556), .A2(n8555), .A3(n8554), .A4(n8553), .ZN(n14911)
         );
  NAND4_X1 U7470 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n12206)
         );
  NAND4_X1 U7471 ( .A1(n8598), .A2(n8597), .A3(n8596), .A4(n8595), .ZN(n12205)
         );
  INV_X1 U7472 ( .A(n13739), .ZN(n6878) );
  INV_X1 U7473 ( .A(n10400), .ZN(n10312) );
  NAND2_X2 U7474 ( .A1(n9595), .A2(n9592), .ZN(n13741) );
  NOR2_X1 U7475 ( .A1(n9767), .A2(n9044), .ZN(n9831) );
  INV_X2 U7476 ( .A(n12886), .ZN(n12833) );
  NAND2_X1 U7477 ( .A1(n7244), .A2(n13412), .ZN(n9875) );
  OR2_X1 U7478 ( .A1(n15331), .A2(n15330), .ZN(n6977) );
  CLKBUF_X1 U7479 ( .A(n8002), .Z(n6531) );
  XNOR2_X1 U7480 ( .A(n8909), .B(P3_IR_REG_21__SCAN_IN), .ZN(n11633) );
  CLKBUF_X3 U7481 ( .A(n11764), .Z(n6533) );
  CLKBUF_X1 U7482 ( .A(n7971), .Z(n8268) );
  NAND2_X1 U7483 ( .A1(n9766), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9837) );
  MUX2_X1 U7484 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14308), .S(n7759), .Z(n10400)
         );
  AND2_X1 U7485 ( .A1(n9591), .A2(n9511), .ZN(n7544) );
  NAND4_X1 U7486 ( .A1(n9380), .A2(n9379), .A3(n9378), .A4(n9377), .ZN(n13074)
         );
  CLKBUF_X2 U7487 ( .A(n8540), .Z(n6537) );
  NOR2_X1 U7488 ( .A1(n7560), .A2(n7561), .ZN(n7563) );
  NAND2_X1 U7489 ( .A1(n11833), .A2(n8912), .ZN(n8537) );
  NOR2_X1 U7490 ( .A1(n7874), .A2(n6721), .ZN(n7171) );
  INV_X1 U7491 ( .A(n8324), .ZN(n7971) );
  AND2_X1 U7492 ( .A1(n8759), .A2(n8758), .ZN(n8778) );
  INV_X1 U7493 ( .A(n11375), .ZN(n12963) );
  INV_X1 U7494 ( .A(n11375), .ZN(n6524) );
  NAND2_X2 U7495 ( .A1(n7681), .A2(n14299), .ZN(n8269) );
  XNOR2_X1 U7496 ( .A(n8911), .B(n8910), .ZN(n10110) );
  NAND2_X1 U7497 ( .A1(n7681), .A2(n7680), .ZN(n7771) );
  NAND2_X1 U7498 ( .A1(n7075), .A2(n7073), .ZN(n8912) );
  INV_X2 U7499 ( .A(n7865), .ZN(n8320) );
  INV_X1 U7500 ( .A(n9601), .ZN(n10973) );
  INV_X1 U7501 ( .A(n7678), .ZN(n7681) );
  OAI21_X1 U7502 ( .B1(n8396), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8398) );
  AND2_X1 U7503 ( .A1(n9219), .A2(n6575), .ZN(n13049) );
  XNOR2_X1 U7504 ( .A(n6757), .B(n7693), .ZN(n11295) );
  XNOR2_X1 U7505 ( .A(n7686), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9601) );
  OR2_X1 U7506 ( .A1(n8389), .A2(n7691), .ZN(n7692) );
  XNOR2_X1 U7507 ( .A(n7697), .B(n7696), .ZN(n14306) );
  NAND2_X1 U7508 ( .A1(n12678), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U7509 ( .A1(n8089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6757) );
  XNOR2_X1 U7510 ( .A(n9332), .B(P2_IR_REG_20__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U7511 ( .A1(n8404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U7512 ( .A1(n14291), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U7513 ( .A1(n6545), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9321) );
  XNOR2_X1 U7514 ( .A(n7676), .B(n7675), .ZN(n7677) );
  NAND2_X1 U7515 ( .A1(n6741), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6740) );
  OR2_X1 U7516 ( .A1(n7674), .A2(n7691), .ZN(n7676) );
  XNOR2_X1 U7517 ( .A(n7616), .B(n7617), .ZN(n15342) );
  BUF_X2 U7518 ( .A(n8022), .Z(n8025) );
  INV_X1 U7519 ( .A(n8605), .ZN(n7099) );
  AND2_X2 U7520 ( .A1(n7709), .A2(n7708), .ZN(n9345) );
  NOR2_X1 U7521 ( .A1(n8604), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n7097) );
  INV_X1 U7522 ( .A(n8418), .ZN(n7524) );
  AND2_X1 U7523 ( .A1(n7539), .A2(n8416), .ZN(n7098) );
  NOR2_X1 U7524 ( .A1(n7529), .A2(n7528), .ZN(n7527) );
  NOR2_X1 U7525 ( .A1(n9214), .A2(n9013), .ZN(n7131) );
  AND2_X1 U7526 ( .A1(n6980), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n7614) );
  NOR2_X1 U7527 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n15265), .ZN(n15041) );
  AND4_X1 U7528 ( .A1(n8426), .A2(n8905), .A3(n8910), .A4(n8425), .ZN(n7539)
         );
  NAND4_X1 U7529 ( .A1(n8417), .A2(n8633), .A3(n8666), .A4(n8680), .ZN(n8418)
         );
  AND2_X1 U7530 ( .A1(n8440), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8533) );
  AND2_X1 U7531 ( .A1(n7666), .A2(n7667), .ZN(n6877) );
  AND4_X1 U7532 ( .A1(n9008), .A2(n9007), .A3(n9145), .A4(n9006), .ZN(n9011)
         );
  NAND2_X1 U7533 ( .A1(n7332), .A2(n9213), .ZN(n7330) );
  INV_X4 U7534 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7535 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8633) );
  NOR2_X1 U7536 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n9330) );
  NOR2_X1 U7537 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n9329) );
  INV_X1 U7538 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10079) );
  NOR2_X1 U7539 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n9007) );
  NOR2_X1 U7540 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n9008) );
  INV_X1 U7541 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8583) );
  NOR2_X1 U7542 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n6704) );
  NOR2_X1 U7543 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6706) );
  NOR2_X1 U7544 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6705) );
  INV_X1 U7545 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15265) );
  INV_X1 U7546 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8666) );
  INV_X1 U7547 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9285) );
  NOR2_X1 U7548 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n7669) );
  INV_X1 U7549 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6980) );
  XNOR2_X1 U7550 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n7613) );
  INV_X1 U7551 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8680) );
  INV_X1 U7552 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9145) );
  INV_X1 U7553 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6707) );
  INV_X4 U7554 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7555 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8390) );
  NOR2_X1 U7556 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7661) );
  INV_X1 U7557 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9005) );
  XNOR2_X2 U7558 ( .A(n11927), .B(n11928), .ZN(n12706) );
  NOR2_X4 U7559 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7699) );
  NAND2_X1 U7560 ( .A1(n6877), .A2(n7699), .ZN(n7782) );
  NOR2_X2 U7561 ( .A1(n13386), .A2(n13504), .ZN(n7238) );
  INV_X1 U7562 ( .A(n12834), .ZN(n7205) );
  OAI21_X1 U7563 ( .B1(n6824), .B2(n14949), .A(n12389), .ZN(n12554) );
  NAND3_X2 U7564 ( .A1(n8542), .A2(n8541), .A3(n6794), .ZN(n14945) );
  NAND3_X2 U7565 ( .A1(n9342), .A2(n9340), .A3(n9341), .ZN(n13075) );
  OAI22_X2 U7566 ( .A1(n10059), .A2(n10058), .B1(n10057), .B2(n10056), .ZN(
        n10283) );
  NOR2_X2 U7567 ( .A1(n11301), .A2(n11300), .ZN(n11302) );
  OAI21_X2 U7568 ( .B1(n11459), .B2(n11458), .A(n6822), .ZN(n11461) );
  XNOR2_X1 U7569 ( .A(n8807), .B(n8806), .ZN(n12354) );
  OAI22_X2 U7570 ( .A1(n8601), .A2(n8599), .B1(P1_DATAO_REG_6__SCAN_IN), .B2(
        n9162), .ZN(n8621) );
  INV_X1 U7571 ( .A(n8005), .ZN(n6526) );
  NOR2_X2 U7572 ( .A1(n8949), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n8489) );
  OAI21_X2 U7573 ( .B1(n11509), .B2(n6654), .A(n8751), .ZN(n12535) );
  INV_X1 U7574 ( .A(n9459), .ZN(n6528) );
  OR2_X4 U7575 ( .A1(n14796), .A2(n9333), .ZN(n9459) );
  BUF_X2 U7576 ( .A(n8530), .Z(n6529) );
  CLKBUF_X1 U7577 ( .A(n14306), .Z(n6530) );
  NAND2_X1 U7578 ( .A1(n9346), .A2(n6967), .ZN(n12965) );
  XNOR2_X2 U7579 ( .A(n6739), .B(n9212), .ZN(n9223) );
  NAND2_X2 U7580 ( .A1(n8923), .A2(n11629), .ZN(n9983) );
  CLKBUF_X2 U7581 ( .A(n12813), .Z(n6534) );
  OAI211_X1 U7582 ( .C1(n10495), .C2(n14666), .A(n9529), .B(n9528), .ZN(n12813) );
  AND2_X1 U7583 ( .A1(n7709), .A2(n7708), .ZN(n6535) );
  AND2_X1 U7584 ( .A1(n7709), .A2(n7708), .ZN(n6536) );
  BUF_X8 U7585 ( .A(n9345), .Z(n6967) );
  OR2_X1 U7586 ( .A1(n12686), .A2(n8434), .ZN(n8540) );
  INV_X1 U7587 ( .A(n8002), .ZN(n6539) );
  INV_X2 U7588 ( .A(n6531), .ZN(n8347) );
  OAI21_X1 U7589 ( .B1(n8136), .B2(n8135), .A(n8134), .ZN(n8156) );
  OAI21_X1 U7590 ( .B1(n14383), .B2(n14351), .A(n11783), .ZN(n11815) );
  OR2_X1 U7591 ( .A1(n12627), .A2(n12386), .ZN(n7542) );
  NAND2_X1 U7592 ( .A1(n12401), .A2(n8878), .ZN(n6767) );
  OR2_X1 U7593 ( .A1(n12047), .A2(n12415), .ZN(n8878) );
  NOR2_X1 U7594 ( .A1(n7030), .A2(n7028), .ZN(n7027) );
  INV_X1 U7595 ( .A(n8850), .ZN(n7030) );
  NOR2_X1 U7596 ( .A1(n6543), .A2(n7167), .ZN(n7159) );
  OAI21_X1 U7597 ( .B1(n8248), .B2(n7191), .A(n7190), .ZN(n8286) );
  OR2_X1 U7598 ( .A1(n6667), .A2(n7194), .ZN(n7190) );
  NAND2_X1 U7599 ( .A1(n7193), .A2(n7192), .ZN(n7191) );
  NAND2_X1 U7600 ( .A1(n14340), .A2(n14339), .ZN(n11493) );
  INV_X1 U7601 ( .A(n6537), .ZN(n8897) );
  INV_X1 U7602 ( .A(n6518), .ZN(n8913) );
  INV_X1 U7603 ( .A(n12686), .ZN(n8433) );
  INV_X2 U7604 ( .A(n6527), .ZN(n11774) );
  NAND2_X1 U7605 ( .A1(n13336), .A2(n7137), .ZN(n13322) );
  NOR2_X1 U7606 ( .A1(n13326), .A2(n6802), .ZN(n7137) );
  INV_X1 U7607 ( .A(n13189), .ZN(n6802) );
  INV_X1 U7608 ( .A(n9819), .ZN(n6860) );
  INV_X1 U7609 ( .A(n12415), .ZN(n12386) );
  NAND2_X1 U7610 ( .A1(n7770), .A2(n7769), .ZN(n6710) );
  NOR2_X1 U7611 ( .A1(n7862), .A2(n7859), .ZN(n7349) );
  NAND2_X1 U7612 ( .A1(n6687), .A2(n6686), .ZN(n7860) );
  NAND2_X1 U7613 ( .A1(n6688), .A2(n7835), .ZN(n6687) );
  NAND2_X1 U7614 ( .A1(n7325), .A2(n12877), .ZN(n7324) );
  INV_X1 U7615 ( .A(n12878), .ZN(n7325) );
  NAND2_X1 U7616 ( .A1(n7305), .A2(n7304), .ZN(n7303) );
  NAND2_X1 U7617 ( .A1(n6873), .A2(n6871), .ZN(n8177) );
  NAND2_X1 U7618 ( .A1(n8161), .A2(n6872), .ZN(n6871) );
  AND2_X1 U7619 ( .A1(n12928), .A2(n7316), .ZN(n7315) );
  NAND2_X1 U7620 ( .A1(n7319), .A2(n7317), .ZN(n7316) );
  NAND2_X1 U7621 ( .A1(n6838), .A2(n6604), .ZN(n12989) );
  INV_X1 U7622 ( .A(n12985), .ZN(n6838) );
  INV_X1 U7623 ( .A(n8265), .ZN(n6813) );
  NAND2_X1 U7624 ( .A1(n14195), .A2(n13582), .ZN(n7220) );
  NAND2_X1 U7625 ( .A1(n9839), .A2(n9090), .ZN(n9092) );
  NAND2_X1 U7626 ( .A1(n12208), .A2(n12207), .ZN(n6829) );
  OR2_X1 U7627 ( .A1(n12102), .A2(n12387), .ZN(n11751) );
  OR2_X1 U7628 ( .A1(n12511), .A2(n12494), .ZN(n11714) );
  NAND2_X1 U7629 ( .A1(n7505), .A2(n7507), .ZN(n7503) );
  INV_X1 U7630 ( .A(n8708), .ZN(n6762) );
  NAND2_X1 U7631 ( .A1(n7531), .A2(n7530), .ZN(n7529) );
  INV_X1 U7632 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7531) );
  INV_X1 U7633 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7530) );
  INV_X1 U7634 ( .A(n8490), .ZN(n7077) );
  NOR2_X1 U7635 ( .A1(n8479), .A2(n7430), .ZN(n8480) );
  AND2_X1 U7636 ( .A1(n11915), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7430) );
  INV_X1 U7637 ( .A(n8456), .ZN(n7458) );
  AND2_X1 U7638 ( .A1(n8665), .A2(n8454), .ZN(n7459) );
  NAND2_X1 U7639 ( .A1(n6631), .A2(n7264), .ZN(n7257) );
  INV_X1 U7640 ( .A(n11948), .ZN(n7249) );
  AOI21_X1 U7641 ( .B1(n7338), .B2(n7336), .A(n7335), .ZN(n7334) );
  INV_X1 U7642 ( .A(n12936), .ZN(n7335) );
  NOR2_X1 U7643 ( .A1(n6572), .A2(n7148), .ZN(n7147) );
  INV_X1 U7644 ( .A(n13196), .ZN(n7148) );
  INV_X1 U7645 ( .A(n11138), .ZN(n11140) );
  NAND2_X1 U7646 ( .A1(n10766), .A2(n10765), .ZN(n10801) );
  INV_X1 U7647 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9018) );
  INV_X1 U7648 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9029) );
  INV_X1 U7649 ( .A(n13701), .ZN(n7387) );
  INV_X1 U7650 ( .A(n8314), .ZN(n6697) );
  INV_X1 U7651 ( .A(n7677), .ZN(n7680) );
  OR2_X1 U7652 ( .A1(n14023), .A2(n11595), .ZN(n7221) );
  NOR2_X1 U7653 ( .A1(n14047), .A2(n7425), .ZN(n7424) );
  INV_X1 U7654 ( .A(n7428), .ZN(n7425) );
  NOR2_X1 U7655 ( .A1(n11593), .A2(n6727), .ZN(n7223) );
  OR2_X1 U7656 ( .A1(n6964), .A2(n14149), .ZN(n6963) );
  NAND2_X1 U7657 ( .A1(n6959), .A2(n11414), .ZN(n6958) );
  NAND2_X1 U7658 ( .A1(n10549), .A2(n10548), .ZN(n10622) );
  AND2_X1 U7659 ( .A1(n8356), .A2(n8358), .ZN(n10020) );
  NOR2_X1 U7660 ( .A1(n8348), .A2(n7353), .ZN(n9602) );
  NAND2_X1 U7661 ( .A1(n8228), .A2(n8227), .ZN(n8248) );
  NAND2_X1 U7662 ( .A1(n8225), .A2(n8224), .ZN(n8228) );
  OAI21_X1 U7663 ( .B1(n8155), .B2(n8154), .A(n8157), .ZN(n8173) );
  XNOR2_X1 U7664 ( .A(n8075), .B(SI_16_), .ZN(n8073) );
  NAND2_X1 U7665 ( .A1(n7994), .A2(n7993), .ZN(n7998) );
  XNOR2_X1 U7666 ( .A(n7559), .B(n15082), .ZN(n7607) );
  XNOR2_X1 U7667 ( .A(n7563), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n7622) );
  NOR2_X1 U7668 ( .A1(n7570), .A2(n7569), .ZN(n7636) );
  AOI21_X1 U7669 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14865), .A(n7576), .ZN(
        n7598) );
  NOR2_X1 U7670 ( .A1(n7600), .A2(n7599), .ZN(n7576) );
  NAND2_X1 U7671 ( .A1(n10845), .A2(n7081), .ZN(n12071) );
  AND2_X1 U7672 ( .A1(n12126), .A2(n12018), .ZN(n7100) );
  NAND2_X1 U7673 ( .A1(n7088), .A2(n7085), .ZN(n14340) );
  INV_X1 U7674 ( .A(n7086), .ZN(n7085) );
  NAND2_X1 U7675 ( .A1(n11244), .A2(n7089), .ZN(n7088) );
  OAI21_X1 U7676 ( .B1(n7087), .B2(n11488), .A(n11487), .ZN(n7086) );
  NAND2_X1 U7677 ( .A1(n12686), .A2(n8434), .ZN(n8814) );
  INV_X1 U7678 ( .A(n8434), .ZN(n8435) );
  NOR2_X1 U7679 ( .A1(n10046), .A2(n10035), .ZN(n10148) );
  NAND2_X1 U7680 ( .A1(n6678), .A2(n6677), .ZN(n6994) );
  INV_X1 U7681 ( .A(n10151), .ZN(n6677) );
  NOR2_X1 U7682 ( .A1(n10489), .A2(n10472), .ZN(n10702) );
  NAND2_X1 U7683 ( .A1(n7049), .A2(n7048), .ZN(n11075) );
  INV_X1 U7684 ( .A(n10705), .ZN(n7048) );
  NAND2_X1 U7685 ( .A1(n12441), .A2(n6592), .ZN(n12428) );
  INV_X1 U7686 ( .A(n7516), .ZN(n7515) );
  AOI21_X1 U7687 ( .B1(n7516), .B2(n7514), .A(n7513), .ZN(n7512) );
  NOR2_X1 U7688 ( .A1(n11619), .A2(n7517), .ZN(n7516) );
  NAND2_X1 U7689 ( .A1(n6586), .A2(n7025), .ZN(n7024) );
  NAND2_X1 U7690 ( .A1(n11624), .A2(n8850), .ZN(n7025) );
  OR2_X1 U7691 ( .A1(n12650), .A2(n12495), .ZN(n11626) );
  NOR2_X1 U7692 ( .A1(n12507), .A2(n6580), .ZN(n12493) );
  INV_X1 U7693 ( .A(n9078), .ZN(n8808) );
  INV_X1 U7694 ( .A(n11775), .ZN(n8809) );
  AND2_X1 U7695 ( .A1(n8976), .A2(n8959), .ZN(n9178) );
  AOI21_X1 U7696 ( .B1(n7433), .B2(n7435), .A(n6662), .ZN(n7432) );
  OAI21_X1 U7697 ( .B1(n8446), .B2(n7438), .A(n7436), .ZN(n8586) );
  INV_X1 U7698 ( .A(n7437), .ZN(n7436) );
  OAI21_X1 U7699 ( .B1(n7439), .B2(n7438), .A(n8587), .ZN(n7437) );
  INV_X1 U7700 ( .A(n8448), .ZN(n7438) );
  AND2_X1 U7701 ( .A1(n9125), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8444) );
  AOI21_X1 U7702 ( .B1(n7275), .B2(n12700), .A(n6616), .ZN(n7273) );
  NAND2_X1 U7703 ( .A1(n13568), .A2(n12963), .ZN(n7176) );
  XNOR2_X1 U7704 ( .A(n13439), .B(n13001), .ZN(n13202) );
  XNOR2_X1 U7705 ( .A(n13454), .B(n13252), .ZN(n13247) );
  INV_X1 U7706 ( .A(n7162), .ZN(n7161) );
  NAND2_X1 U7707 ( .A1(n10772), .A2(n10771), .ZN(n10807) );
  INV_X1 U7708 ( .A(n10523), .ZN(n7136) );
  NAND2_X1 U7709 ( .A1(n10170), .A2(n7135), .ZN(n6731) );
  AND2_X1 U7710 ( .A1(n10647), .A2(n13012), .ZN(n7135) );
  OR2_X1 U7711 ( .A1(n6520), .A2(n13412), .ZN(n9886) );
  AND2_X1 U7712 ( .A1(n9360), .A2(n9359), .ZN(n14812) );
  XNOR2_X1 U7713 ( .A(n7130), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9323) );
  OR2_X1 U7714 ( .A1(n9319), .A2(n10301), .ZN(n7130) );
  OAI21_X1 U7715 ( .B1(n6903), .B2(n13745), .A(n6899), .ZN(n6898) );
  NAND2_X1 U7716 ( .A1(n6903), .A2(n6900), .ZN(n6899) );
  NAND2_X1 U7717 ( .A1(n6901), .A2(n6905), .ZN(n6900) );
  NAND2_X1 U7718 ( .A1(n13786), .A2(n6605), .ZN(n13751) );
  AND2_X1 U7719 ( .A1(n9954), .A2(n9952), .ZN(n6882) );
  XNOR2_X1 U7720 ( .A(n14195), .B(n13840), .ZN(n14005) );
  OR2_X1 U7721 ( .A1(n13622), .A2(n13845), .ZN(n6822) );
  OR2_X1 U7722 ( .A1(n13622), .A2(n14441), .ZN(n11455) );
  AOI21_X1 U7723 ( .B1(n11101), .B2(n7409), .A(n11196), .ZN(n7408) );
  INV_X1 U7724 ( .A(n11099), .ZN(n7409) );
  AND2_X1 U7725 ( .A1(n7228), .A2(n7227), .ZN(n7226) );
  NOR2_X1 U7726 ( .A1(n7782), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n7228) );
  NAND2_X1 U7727 ( .A1(n7795), .A2(n6554), .ZN(n6720) );
  NAND2_X1 U7728 ( .A1(n6950), .A2(n7847), .ZN(n6719) );
  OAI21_X1 U7729 ( .B1(n6782), .B2(n6785), .A(n6983), .ZN(n6982) );
  INV_X1 U7730 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6983) );
  INV_X1 U7731 ( .A(n6784), .ZN(n6785) );
  OAI21_X1 U7732 ( .B1(n11830), .B2(n11829), .A(n6809), .ZN(n6808) );
  NOR2_X1 U7733 ( .A1(n11831), .A2(n6810), .ZN(n6809) );
  NOR2_X1 U7734 ( .A1(n12380), .A2(n6825), .ZN(n6824) );
  OR2_X1 U7735 ( .A1(n11370), .A2(n9028), .ZN(n9388) );
  OR2_X1 U7736 ( .A1(n12817), .A2(n12816), .ZN(n12818) );
  AND2_X1 U7737 ( .A1(n7766), .A2(n10379), .ZN(n6865) );
  NAND2_X1 U7738 ( .A1(n7763), .A2(n7989), .ZN(n7765) );
  NAND2_X1 U7739 ( .A1(n6709), .A2(n6708), .ZN(n7814) );
  OAI21_X1 U7740 ( .B1(n7860), .B2(n7349), .A(n6620), .ZN(n7884) );
  NAND2_X1 U7741 ( .A1(n7860), .A2(n6684), .ZN(n6746) );
  NOR2_X1 U7742 ( .A1(n6685), .A2(n6747), .ZN(n6684) );
  INV_X1 U7743 ( .A(n7348), .ZN(n6685) );
  INV_X1 U7744 ( .A(n6745), .ZN(n6744) );
  OAI21_X1 U7745 ( .B1(n6549), .B2(n6747), .A(n6621), .ZN(n6745) );
  NAND2_X1 U7746 ( .A1(n7990), .A2(n7992), .ZN(n7359) );
  NOR2_X1 U7747 ( .A1(n12890), .A2(n12887), .ZN(n7305) );
  NAND2_X1 U7748 ( .A1(n12890), .A2(n12887), .ZN(n7304) );
  OAI21_X1 U7749 ( .B1(n12879), .B2(n7326), .A(n6850), .ZN(n12884) );
  AND2_X1 U7750 ( .A1(n7324), .A2(n7323), .ZN(n6850) );
  NAND2_X1 U7751 ( .A1(n14149), .A2(n6590), .ZN(n6804) );
  OAI21_X1 U7752 ( .B1(n12904), .B2(n12903), .A(n12901), .ZN(n12907) );
  NAND2_X1 U7753 ( .A1(n6690), .A2(n8122), .ZN(n8141) );
  NAND2_X1 U7754 ( .A1(n6691), .A2(n14144), .ZN(n6690) );
  NAND2_X1 U7755 ( .A1(n7318), .A2(n12923), .ZN(n7317) );
  INV_X1 U7756 ( .A(n12924), .ZN(n7318) );
  INV_X1 U7757 ( .A(n8192), .ZN(n6826) );
  NAND2_X1 U7758 ( .A1(n6695), .A2(n6694), .ZN(n6693) );
  NAND2_X1 U7759 ( .A1(n6753), .A2(n8175), .ZN(n6752) );
  INV_X1 U7760 ( .A(n8176), .ZN(n6694) );
  NAND2_X1 U7761 ( .A1(n8215), .A2(n7355), .ZN(n7354) );
  INV_X1 U7762 ( .A(n8214), .ZN(n7355) );
  AND2_X1 U7763 ( .A1(n7320), .A2(n12924), .ZN(n7319) );
  INV_X1 U7764 ( .A(n12923), .ZN(n7320) );
  INV_X1 U7765 ( .A(n7317), .ZN(n6852) );
  INV_X1 U7766 ( .A(n12919), .ZN(n6848) );
  INV_X1 U7767 ( .A(n8050), .ZN(n8052) );
  NAND2_X1 U7768 ( .A1(n6819), .A2(n8672), .ZN(n8671) );
  NAND2_X1 U7769 ( .A1(n7351), .A2(n7353), .ZN(n7350) );
  NAND2_X1 U7770 ( .A1(n8296), .A2(n7344), .ZN(n7343) );
  INV_X1 U7771 ( .A(n8295), .ZN(n7344) );
  NAND2_X1 U7772 ( .A1(n7342), .A2(n8253), .ZN(n7341) );
  AOI21_X1 U7773 ( .B1(n8235), .B2(n8236), .A(n6751), .ZN(n6750) );
  NOR2_X1 U7774 ( .A1(n8052), .A2(SI_14_), .ZN(n8055) );
  INV_X1 U7775 ( .A(n7997), .ZN(n7189) );
  INV_X1 U7776 ( .A(n7956), .ZN(n7181) );
  NAND2_X1 U7777 ( .A1(n6771), .A2(n6770), .ZN(n7558) );
  NAND2_X1 U7778 ( .A1(n6772), .A2(n6790), .ZN(n6770) );
  INV_X1 U7779 ( .A(n10848), .ZN(n7082) );
  INV_X1 U7780 ( .A(n11120), .ZN(n7080) );
  NOR2_X1 U7781 ( .A1(n11813), .A2(n11814), .ZN(n7471) );
  NAND2_X1 U7782 ( .A1(n11075), .A2(n11074), .ZN(n6830) );
  OR2_X1 U7783 ( .A1(n12642), .A2(n12470), .ZN(n11620) );
  OR2_X1 U7784 ( .A1(n12655), .A2(n12509), .ZN(n11724) );
  OAI21_X1 U7785 ( .B1(n8707), .B2(n6762), .A(n8722), .ZN(n6761) );
  INV_X1 U7786 ( .A(n11317), .ZN(n6763) );
  OR2_X1 U7787 ( .A1(n14393), .A2(n14372), .ZN(n11691) );
  INV_X1 U7788 ( .A(n14376), .ZN(n7486) );
  OR2_X1 U7789 ( .A1(n12076), .A2(n14378), .ZN(n11682) );
  NAND2_X1 U7790 ( .A1(n10433), .A2(n6607), .ZN(n10910) );
  NAND2_X1 U7791 ( .A1(n6764), .A2(n6766), .ZN(n10433) );
  AND2_X1 U7792 ( .A1(n8575), .A2(n10434), .ZN(n6764) );
  NAND2_X1 U7793 ( .A1(n14945), .A2(n14924), .ZN(n11637) );
  NAND2_X1 U7794 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), 
        .ZN(n7074) );
  AOI21_X1 U7795 ( .B1(n8620), .B2(n8452), .A(n6629), .ZN(n7453) );
  INV_X1 U7796 ( .A(n8452), .ZN(n7451) );
  AND2_X1 U7797 ( .A1(n7440), .A2(n8445), .ZN(n7439) );
  INV_X1 U7798 ( .A(n8569), .ZN(n7440) );
  NAND2_X1 U7799 ( .A1(n6933), .A2(n11524), .ZN(n6932) );
  INV_X1 U7800 ( .A(n7257), .ZN(n6933) );
  XNOR2_X1 U7801 ( .A(n13509), .B(n7249), .ZN(n11844) );
  BUF_X1 U7802 ( .A(n9744), .Z(n11948) );
  INV_X1 U7803 ( .A(n12989), .ZN(n6799) );
  NOR2_X1 U7804 ( .A1(n12988), .A2(n12987), .ZN(n6798) );
  INV_X1 U7805 ( .A(n9534), .ZN(n9970) );
  INV_X1 U7806 ( .A(n9324), .ZN(n9322) );
  NOR2_X1 U7807 ( .A1(n13439), .A2(n13228), .ZN(n7233) );
  OAI21_X1 U7808 ( .B1(n13197), .B2(n6572), .A(n13247), .ZN(n7151) );
  INV_X1 U7809 ( .A(n13247), .ZN(n7112) );
  NOR2_X1 U7810 ( .A1(n13171), .A2(n7111), .ZN(n7110) );
  INV_X1 U7811 ( .A(n13169), .ZN(n7111) );
  NAND2_X1 U7812 ( .A1(n13308), .A2(n13191), .ZN(n13193) );
  NOR2_X1 U7813 ( .A1(n7157), .A2(n13021), .ZN(n7153) );
  INV_X1 U7814 ( .A(n13023), .ZN(n7157) );
  NAND2_X1 U7815 ( .A1(n13023), .A2(n7156), .ZN(n7155) );
  INV_X1 U7816 ( .A(n11212), .ZN(n7156) );
  INV_X1 U7817 ( .A(n10774), .ZN(n7140) );
  NAND2_X1 U7818 ( .A1(n14800), .A2(n9381), .ZN(n9877) );
  XNOR2_X1 U7819 ( .A(n12806), .B(n12968), .ZN(n7244) );
  NAND2_X1 U7820 ( .A1(n9936), .A2(n9872), .ZN(n10115) );
  OR2_X1 U7821 ( .A1(n9207), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9283) );
  AND2_X1 U7822 ( .A1(n7353), .A2(n10973), .ZN(n9592) );
  NOR2_X1 U7823 ( .A1(n13978), .A2(n7007), .ZN(n7006) );
  INV_X1 U7824 ( .A(n7008), .ZN(n7007) );
  NOR2_X1 U7825 ( .A1(n13985), .A2(n13982), .ZN(n7008) );
  INV_X1 U7826 ( .A(n14005), .ZN(n7216) );
  OAI21_X1 U7827 ( .B1(n14144), .B2(n7202), .A(n11589), .ZN(n7201) );
  OR2_X1 U7828 ( .A1(n14244), .A2(n14137), .ZN(n11589) );
  NAND2_X1 U7829 ( .A1(n7012), .A2(n11599), .ZN(n7011) );
  NOR2_X1 U7830 ( .A1(n14249), .A2(n14259), .ZN(n7012) );
  OAI21_X1 U7831 ( .B1(n14162), .B2(n6965), .A(n6966), .ZN(n6964) );
  INV_X1 U7832 ( .A(n11585), .ZN(n6965) );
  NOR2_X1 U7833 ( .A1(n7419), .A2(n11578), .ZN(n7418) );
  INV_X1 U7834 ( .A(n7420), .ZN(n7419) );
  NAND2_X1 U7835 ( .A1(n6814), .A2(n10415), .ZN(n8356) );
  NAND2_X1 U7836 ( .A1(n8305), .A2(n8304), .ZN(n8310) );
  NAND2_X1 U7837 ( .A1(n8310), .A2(n8309), .ZN(n8327) );
  XNOR2_X1 U7838 ( .A(n8156), .B(n10112), .ZN(n8155) );
  AOI21_X1 U7839 ( .B1(n7187), .B2(n7188), .A(n7186), .ZN(n7185) );
  OR2_X1 U7840 ( .A1(n7959), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n7960) );
  NOR2_X1 U7841 ( .A1(n7957), .A2(n7183), .ZN(n7182) );
  INV_X1 U7842 ( .A(n7936), .ZN(n7183) );
  XNOR2_X1 U7843 ( .A(n7979), .B(n15171), .ZN(n7977) );
  NAND2_X1 U7844 ( .A1(n7916), .A2(SI_10_), .ZN(n7936) );
  OAI22_X1 U7845 ( .A1(n7628), .A2(n7567), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n7566), .ZN(n7568) );
  OAI21_X1 U7846 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15304), .A(n7573), .ZN(
        n7574) );
  INV_X1 U7847 ( .A(n14518), .ZN(n6774) );
  AOI21_X1 U7848 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15285), .A(n7577), .ZN(
        n7596) );
  INV_X1 U7849 ( .A(n14943), .ZN(n8922) );
  NAND2_X1 U7850 ( .A1(n10858), .A2(n10837), .ZN(n10845) );
  NOR2_X1 U7851 ( .A1(n8869), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8870) );
  INV_X1 U7852 ( .A(n11815), .ZN(n11825) );
  OAI21_X1 U7853 ( .B1(n9677), .B2(n9678), .A(n9085), .ZN(n9662) );
  NAND2_X1 U7854 ( .A1(n9072), .A2(n6827), .ZN(n9767) );
  OR2_X1 U7855 ( .A1(n9071), .A2(n9774), .ZN(n6827) );
  OAI21_X1 U7856 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n9833) );
  NAND2_X1 U7857 ( .A1(n9837), .A2(n9835), .ZN(n6679) );
  NAND2_X1 U7858 ( .A1(n9808), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9807) );
  INV_X1 U7859 ( .A(n6996), .ZN(n10146) );
  NOR2_X1 U7860 ( .A1(n10709), .A2(n10710), .ZN(n10712) );
  INV_X1 U7861 ( .A(n6992), .ZN(n10707) );
  XNOR2_X1 U7862 ( .A(n6830), .B(n14866), .ZN(n14871) );
  INV_X1 U7863 ( .A(n11078), .ZN(n7061) );
  XNOR2_X1 U7864 ( .A(n6829), .B(n6828), .ZN(n14887) );
  NAND2_X1 U7865 ( .A1(n7043), .A2(n12223), .ZN(n7042) );
  OAI211_X1 U7866 ( .C1(n12255), .C2(n12268), .A(n6990), .B(n6991), .ZN(n12257) );
  OR2_X1 U7867 ( .A1(n12268), .A2(n12256), .ZN(n6991) );
  NOR2_X1 U7868 ( .A1(n11748), .A2(n7494), .ZN(n7493) );
  AND2_X1 U7869 ( .A1(n8884), .A2(n12098), .ZN(n14352) );
  OR2_X1 U7870 ( .A1(n12620), .A2(n12387), .ZN(n7553) );
  OR2_X1 U7871 ( .A1(n12631), .A2(n12145), .ZN(n7552) );
  INV_X1 U7872 ( .A(n7023), .ZN(n7020) );
  AND2_X1 U7873 ( .A1(n12442), .A2(n7022), .ZN(n7021) );
  INV_X1 U7874 ( .A(n7024), .ZN(n7022) );
  NAND2_X1 U7875 ( .A1(n12112), .A2(n12458), .ZN(n7519) );
  NOR2_X1 U7876 ( .A1(n8938), .A2(n7521), .ZN(n7520) );
  INV_X1 U7877 ( .A(n11626), .ZN(n7521) );
  AND2_X1 U7878 ( .A1(n11621), .A2(n11620), .ZN(n12461) );
  OR2_X1 U7879 ( .A1(n11624), .A2(n11623), .ZN(n12472) );
  AND4_X1 U7880 ( .A1(n8829), .A2(n8828), .A3(n8827), .A4(n8826), .ZN(n12495)
         );
  AND2_X1 U7881 ( .A1(n11714), .A2(n11719), .ZN(n11806) );
  NAND2_X1 U7882 ( .A1(n12532), .A2(n12531), .ZN(n7492) );
  INV_X1 U7883 ( .A(n11693), .ZN(n7509) );
  AND2_X1 U7884 ( .A1(n11702), .A2(n11707), .ZN(n11802) );
  AOI21_X1 U7885 ( .B1(n7508), .B2(n11690), .A(n7506), .ZN(n7505) );
  INV_X1 U7886 ( .A(n11699), .ZN(n7506) );
  INV_X1 U7887 ( .A(n12201), .ZN(n11432) );
  NAND2_X1 U7888 ( .A1(n6763), .A2(n8707), .ZN(n11320) );
  AOI21_X1 U7889 ( .B1(n11062), .B2(n7491), .A(n7490), .ZN(n7489) );
  INV_X1 U7890 ( .A(n11672), .ZN(n7491) );
  INV_X1 U7891 ( .A(n11675), .ZN(n7490) );
  INV_X1 U7892 ( .A(n7475), .ZN(n7474) );
  OAI21_X1 U7893 ( .B1(n7546), .B2(n7477), .A(n11669), .ZN(n7475) );
  OR2_X1 U7894 ( .A1(n12205), .A2(n10916), .ZN(n11660) );
  CLKBUF_X1 U7895 ( .A(n10433), .Z(n6795) );
  OR2_X1 U7896 ( .A1(n9993), .A2(n11755), .ZN(n14932) );
  NAND2_X1 U7897 ( .A1(n9993), .A2(n11736), .ZN(n14930) );
  AND2_X1 U7898 ( .A1(n14351), .A2(n14350), .ZN(n14386) );
  NAND2_X1 U7899 ( .A1(n8492), .A2(n8491), .ZN(n12014) );
  NAND2_X1 U7900 ( .A1(n8998), .A2(n10418), .ZN(n15013) );
  AND2_X1 U7901 ( .A1(n9779), .A2(n12673), .ZN(n9794) );
  NAND2_X1 U7902 ( .A1(n8487), .A2(n8427), .ZN(n7528) );
  INV_X1 U7903 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U7904 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n14303), .ZN(n6854) );
  NOR2_X1 U7905 ( .A1(n7529), .A2(P3_IR_REG_25__SCAN_IN), .ZN(n7041) );
  AND2_X1 U7906 ( .A1(n8952), .A2(n8951), .ZN(n8976) );
  XNOR2_X1 U7907 ( .A(n8480), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n8497) );
  AND2_X1 U7908 ( .A1(n15205), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6805) );
  INV_X1 U7909 ( .A(n8839), .ZN(n6806) );
  INV_X1 U7910 ( .A(n8840), .ZN(n6807) );
  OAI21_X1 U7911 ( .B1(n8804), .B2(n8802), .A(n8476), .ZN(n7469) );
  AOI21_X1 U7912 ( .B1(n7434), .B2(n8472), .A(n6665), .ZN(n7433) );
  INV_X1 U7913 ( .A(n8471), .ZN(n7434) );
  INV_X1 U7914 ( .A(n8472), .ZN(n7435) );
  NAND2_X1 U7915 ( .A1(n7460), .A2(n7461), .ZN(n8754) );
  AOI21_X1 U7916 ( .B1(n7463), .B2(n8466), .A(n7462), .ZN(n7461) );
  INV_X1 U7917 ( .A(n8469), .ZN(n7462) );
  AND2_X1 U7918 ( .A1(n8471), .A2(n8470), .ZN(n8753) );
  INV_X1 U7919 ( .A(n8726), .ZN(n7467) );
  INV_X1 U7920 ( .A(n7457), .ZN(n7456) );
  NAND2_X1 U7921 ( .A1(n6568), .A2(n7459), .ZN(n8664) );
  NAND2_X1 U7922 ( .A1(n9169), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U7923 ( .A1(n7455), .A2(n7454), .ZN(n8623) );
  INV_X1 U7924 ( .A(n8620), .ZN(n7454) );
  INV_X1 U7925 ( .A(n8621), .ZN(n7455) );
  NAND2_X1 U7926 ( .A1(n8446), .A2(n7439), .ZN(n8572) );
  NOR2_X1 U7927 ( .A1(n7047), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8584) );
  OAI22_X1 U7928 ( .A1(n8548), .A2(n8443), .B1(P2_DATAO_REG_2__SCAN_IN), .B2(
        n9526), .ZN(n8559) );
  NAND2_X1 U7929 ( .A1(n8546), .A2(n9084), .ZN(n7047) );
  NOR2_X1 U7930 ( .A1(n12789), .A2(n11958), .ZN(n7250) );
  OR2_X1 U7931 ( .A1(n11972), .A2(n11971), .ZN(n11973) );
  AND2_X1 U7932 ( .A1(n10280), .A2(n10281), .ZN(n6928) );
  NAND2_X1 U7933 ( .A1(n10881), .A2(n7266), .ZN(n7265) );
  INV_X1 U7934 ( .A(n10882), .ZN(n7266) );
  NOR2_X1 U7935 ( .A1(n10883), .A2(n7262), .ZN(n7261) );
  NOR2_X1 U7936 ( .A1(n14637), .A2(n7263), .ZN(n7262) );
  AND2_X1 U7937 ( .A1(n11395), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11534) );
  INV_X1 U7938 ( .A(n12741), .ZN(n7283) );
  NAND2_X1 U7939 ( .A1(n12706), .A2(n12707), .ZN(n7247) );
  XNOR2_X1 U7940 ( .A(n6522), .B(n11948), .ZN(n9737) );
  OR2_X1 U7941 ( .A1(n10752), .A2(n10751), .ZN(n10893) );
  NAND2_X1 U7942 ( .A1(n7253), .A2(n7252), .ZN(n7255) );
  NOR2_X1 U7943 ( .A1(n11520), .A2(n7258), .ZN(n7252) );
  INV_X1 U7944 ( .A(n7261), .ZN(n7253) );
  INV_X1 U7945 ( .A(n7265), .ZN(n7258) );
  NAND2_X1 U7946 ( .A1(n7264), .A2(n6663), .ZN(n7256) );
  OR2_X1 U7947 ( .A1(n10733), .A2(n7257), .ZN(n6935) );
  AND2_X1 U7948 ( .A1(n11847), .A2(n7283), .ZN(n7282) );
  XNOR2_X1 U7949 ( .A(n13460), .B(n7249), .ZN(n11972) );
  OR2_X1 U7950 ( .A1(n12937), .A2(n12936), .ZN(n12938) );
  AND2_X1 U7951 ( .A1(n9324), .A2(n13569), .ZN(n9649) );
  NAND2_X1 U7952 ( .A1(n13259), .A2(n13274), .ZN(n7113) );
  AOI21_X1 U7953 ( .B1(n13251), .B2(n13197), .A(n6572), .ZN(n7149) );
  NAND2_X1 U7954 ( .A1(n13237), .A2(n13407), .ZN(n6842) );
  NAND2_X1 U7955 ( .A1(n13289), .A2(n13167), .ZN(n13267) );
  NAND2_X1 U7956 ( .A1(n13299), .A2(n7126), .ZN(n13289) );
  AND2_X1 U7957 ( .A1(n13290), .A2(n13166), .ZN(n7126) );
  INV_X1 U7958 ( .A(n13193), .ZN(n7133) );
  NAND2_X1 U7959 ( .A1(n13480), .A2(n7127), .ZN(n13299) );
  NOR2_X1 U7960 ( .A1(n13307), .A2(n7128), .ZN(n7127) );
  INV_X1 U7961 ( .A(n13165), .ZN(n7128) );
  NOR2_X1 U7962 ( .A1(n13184), .A2(n7164), .ZN(n7163) );
  INV_X1 U7963 ( .A(n13181), .ZN(n7164) );
  NOR2_X1 U7964 ( .A1(n13157), .A2(n7121), .ZN(n7120) );
  INV_X1 U7965 ( .A(n13156), .ZN(n7121) );
  AOI21_X1 U7966 ( .B1(n13027), .B2(n7124), .A(n6553), .ZN(n7122) );
  INV_X1 U7967 ( .A(n7124), .ZN(n7123) );
  NAND2_X1 U7968 ( .A1(n6736), .A2(n7143), .ZN(n13177) );
  INV_X1 U7969 ( .A(n7144), .ZN(n7143) );
  OAI21_X1 U7970 ( .B1(n11544), .B2(n13403), .A(n11546), .ZN(n7144) );
  NAND2_X1 U7971 ( .A1(n11558), .A2(n11557), .ZN(n7125) );
  OR2_X1 U7972 ( .A1(n10893), .A2(n14648), .ZN(n11388) );
  AOI21_X1 U7973 ( .B1(n11211), .B2(n13021), .A(n11210), .ZN(n11404) );
  NAND2_X1 U7974 ( .A1(n11140), .A2(n11139), .ZN(n11213) );
  AND2_X1 U7975 ( .A1(n7134), .A2(n13016), .ZN(n6730) );
  AND2_X1 U7976 ( .A1(n7104), .A2(n10641), .ZN(n7103) );
  NAND2_X1 U7977 ( .A1(n10170), .A2(n13012), .ZN(n10524) );
  NAND2_X1 U7978 ( .A1(n6738), .A2(n13010), .ZN(n10209) );
  NAND2_X1 U7979 ( .A1(n11975), .A2(n11974), .ZN(n13454) );
  NAND2_X1 U7980 ( .A1(n11947), .A2(n11946), .ZN(n13276) );
  NAND2_X1 U7981 ( .A1(n11890), .A2(n11889), .ZN(n13488) );
  NAND2_X1 U7982 ( .A1(n11850), .A2(n11849), .ZN(n13504) );
  INV_X1 U7983 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9017) );
  INV_X1 U7984 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9213) );
  INV_X1 U7985 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7288) );
  NOR2_X1 U7986 ( .A1(n9283), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9286) );
  AOI21_X1 U7987 ( .B1(n7385), .B2(n7387), .A(n6625), .ZN(n7382) );
  AND2_X1 U7988 ( .A1(n13618), .A2(n6891), .ZN(n6890) );
  NAND2_X1 U7989 ( .A1(n6892), .A2(n13795), .ZN(n6891) );
  INV_X1 U7990 ( .A(n7388), .ZN(n6892) );
  NAND2_X1 U7991 ( .A1(n13814), .A2(n13813), .ZN(n7396) );
  AND2_X1 U7992 ( .A1(n13822), .A2(n7386), .ZN(n7385) );
  OR2_X1 U7993 ( .A1(n13771), .A2(n7387), .ZN(n7386) );
  NOR2_X1 U7994 ( .A1(n13760), .A2(n7393), .ZN(n7392) );
  INV_X1 U7995 ( .A(n13599), .ZN(n7393) );
  INV_X1 U7996 ( .A(n6886), .ZN(n6885) );
  OAI21_X1 U7997 ( .B1(n13805), .B2(n6887), .A(n13717), .ZN(n6886) );
  INV_X1 U7998 ( .A(n13679), .ZN(n6887) );
  NOR2_X1 U7999 ( .A1(n7397), .A2(n6909), .ZN(n6908) );
  INV_X1 U8000 ( .A(n11019), .ZN(n6909) );
  NAND2_X1 U8001 ( .A1(n6912), .A2(n7398), .ZN(n7397) );
  NAND2_X1 U8002 ( .A1(n13751), .A2(n13671), .ZN(n13804) );
  NAND2_X1 U8003 ( .A1(n10194), .A2(n10193), .ZN(n7371) );
  NAND2_X1 U8004 ( .A1(n7378), .A2(n10337), .ZN(n7377) );
  NAND2_X1 U8005 ( .A1(n7375), .A2(n10194), .ZN(n6881) );
  NOR2_X1 U8006 ( .A1(n7376), .A2(n6578), .ZN(n7375) );
  OR2_X1 U8007 ( .A1(n8372), .A2(n8373), .ZN(n8383) );
  NAND2_X1 U8008 ( .A1(n7364), .A2(n7365), .ZN(n7363) );
  AOI21_X1 U8009 ( .B1(n8315), .B2(n8316), .A(n6697), .ZN(n6696) );
  OAI21_X1 U8010 ( .B1(n8315), .B2(n8316), .A(n7362), .ZN(n6759) );
  NAND2_X1 U8011 ( .A1(n6880), .A2(n6879), .ZN(n9595) );
  NOR2_X1 U8012 ( .A1(n11450), .A2(n11372), .ZN(n6879) );
  AND2_X1 U8013 ( .A1(n7006), .A2(n7005), .ZN(n7003) );
  INV_X1 U8014 ( .A(n14171), .ZN(n7005) );
  INV_X1 U8015 ( .A(n7006), .ZN(n7001) );
  NAND2_X1 U8016 ( .A1(n6969), .A2(n6728), .ZN(n14023) );
  NAND2_X1 U8017 ( .A1(n6972), .A2(n6970), .ZN(n6728) );
  INV_X1 U8018 ( .A(n7422), .ZN(n7421) );
  OAI22_X1 U8019 ( .A1(n14020), .A2(n7426), .B1(n14031), .B2(n13772), .ZN(
        n7422) );
  NAND2_X1 U8020 ( .A1(n14070), .A2(n7014), .ZN(n14029) );
  AND2_X1 U8021 ( .A1(n6551), .A2(n14031), .ZN(n7014) );
  NAND2_X1 U8022 ( .A1(n14209), .A2(n13841), .ZN(n7426) );
  NAND2_X1 U8023 ( .A1(n6836), .A2(n7424), .ZN(n7427) );
  NAND2_X1 U8024 ( .A1(n14069), .A2(n7223), .ZN(n6973) );
  NAND2_X1 U8025 ( .A1(n6962), .A2(n14144), .ZN(n7203) );
  NOR2_X1 U8026 ( .A1(n6581), .A2(n7416), .ZN(n7415) );
  INV_X1 U8027 ( .A(n11577), .ZN(n7416) );
  INV_X1 U8028 ( .A(n7203), .ZN(n14131) );
  NOR2_X1 U8029 ( .A1(n14259), .A2(n11584), .ZN(n11585) );
  OAI211_X1 U8030 ( .C1(n6956), .C2(n6955), .A(n6954), .B(n6659), .ZN(n11475)
         );
  INV_X1 U8031 ( .A(n6955), .ZN(n6952) );
  NAND2_X1 U8032 ( .A1(n13631), .A2(n13629), .ZN(n7420) );
  AND2_X1 U8033 ( .A1(n6958), .A2(n11458), .ZN(n6956) );
  NAND2_X1 U8034 ( .A1(n11101), .A2(n11308), .ZN(n7406) );
  CLKBUF_X1 U8035 ( .A(n11100), .Z(n6835) );
  AOI21_X1 U8036 ( .B1(n10667), .B2(n10626), .A(n10625), .ZN(n10629) );
  XNOR2_X1 U8037 ( .A(n11030), .B(n10624), .ZN(n10666) );
  NAND2_X1 U8038 ( .A1(n10660), .A2(n10666), .ZN(n10659) );
  NOR2_X1 U8039 ( .A1(n10575), .A2(n10579), .ZN(n10574) );
  XNOR2_X1 U8040 ( .A(n8342), .B(n8337), .ZN(n12964) );
  NAND2_X1 U8041 ( .A1(n7670), .A2(n8025), .ZN(n8402) );
  XNOR2_X1 U8042 ( .A(n8205), .B(n8841), .ZN(n11335) );
  AND2_X1 U8043 ( .A1(n7367), .A2(n7688), .ZN(n7366) );
  OAI21_X1 U8044 ( .B1(n7998), .B2(n7188), .A(n7187), .ZN(n8074) );
  NOR2_X1 U8045 ( .A1(n7851), .A2(n7172), .ZN(n6721) );
  INV_X1 U8046 ( .A(n7871), .ZN(n7172) );
  NAND2_X1 U8047 ( .A1(n7872), .A2(n7871), .ZN(n7876) );
  NAND2_X1 U8048 ( .A1(n7852), .A2(n7851), .ZN(n7872) );
  OR2_X1 U8049 ( .A1(n6723), .A2(SI_5_), .ZN(n6722) );
  NAND2_X1 U8050 ( .A1(n7795), .A2(n7794), .ZN(n7796) );
  INV_X1 U8051 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U8052 ( .A1(n6535), .A2(n8531), .ZN(n6861) );
  NAND2_X1 U8053 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6789), .ZN(n6788) );
  INV_X1 U8054 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6789) );
  AND2_X1 U8055 ( .A1(n15265), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n6790) );
  XNOR2_X1 U8056 ( .A(n7607), .B(n7606), .ZN(n7608) );
  INV_X1 U8057 ( .A(n6976), .ZN(n7623) );
  OR2_X1 U8058 ( .A1(n9467), .A2(n7574), .ZN(n7602) );
  AND2_X1 U8059 ( .A1(n6787), .A2(n14520), .ZN(n7645) );
  AND4_X1 U8060 ( .A1(n8788), .A2(n8787), .A3(n8786), .A4(n8785), .ZN(n12020)
         );
  NOR2_X1 U8061 ( .A1(n11494), .A2(n7102), .ZN(n7101) );
  INV_X1 U8062 ( .A(n11492), .ZN(n7102) );
  NOR2_X1 U8063 ( .A1(n12139), .A2(n6655), .ZN(n7084) );
  AND2_X1 U8064 ( .A1(n8683), .A2(n8682), .ZN(n11130) );
  NAND2_X1 U8065 ( .A1(n8794), .A2(n8793), .ZN(n12511) );
  NAND4_X1 U8066 ( .A1(n8647), .A2(n8646), .A3(n8645), .A4(n8644), .ZN(n12202)
         );
  OR2_X1 U8067 ( .A1(n10702), .A2(n10703), .ZN(n7049) );
  AOI21_X1 U8068 ( .B1(n12681), .B2(n11774), .A(n11763), .ZN(n14383) );
  NAND2_X1 U8069 ( .A1(n11777), .A2(n11776), .ZN(n14387) );
  NAND2_X1 U8070 ( .A1(n12398), .A2(n11613), .ZN(n12384) );
  INV_X1 U8071 ( .A(n12014), .ZN(n12624) );
  NAND2_X1 U8072 ( .A1(n8823), .A2(n8822), .ZN(n12650) );
  NAND2_X1 U8073 ( .A1(n8781), .A2(n8780), .ZN(n12659) );
  INV_X1 U8074 ( .A(n13454), .ZN(n13240) );
  AND2_X1 U8075 ( .A1(n10733), .A2(n10732), .ZN(n14638) );
  NOR2_X1 U8076 ( .A1(n7271), .A2(n14652), .ZN(n7269) );
  AND2_X1 U8077 ( .A1(n7273), .A2(n6652), .ZN(n7271) );
  NAND2_X1 U8078 ( .A1(n7273), .A2(n7274), .ZN(n7272) );
  INV_X1 U8079 ( .A(n7275), .ZN(n7274) );
  NAND2_X1 U8080 ( .A1(n6735), .A2(n14798), .ZN(n6734) );
  NAND2_X1 U8081 ( .A1(n11209), .A2(n11208), .ZN(n14658) );
  NAND2_X1 U8082 ( .A1(n14817), .A2(n9382), .ZN(n14803) );
  OAI21_X1 U8083 ( .B1(n13445), .B2(n13529), .A(n13448), .ZN(n13540) );
  NAND2_X1 U8084 ( .A1(n9371), .A2(n9370), .ZN(n14816) );
  NOR2_X1 U8085 ( .A1(n6557), .A2(n14476), .ZN(n6895) );
  NAND2_X1 U8086 ( .A1(n6898), .A2(n6902), .ZN(n6897) );
  NAND2_X1 U8087 ( .A1(n13745), .A2(n13737), .ZN(n6902) );
  AND4_X1 U8088 ( .A1(n8037), .A2(n8036), .A3(n8035), .A4(n8034), .ZN(n14441)
         );
  NAND2_X1 U8089 ( .A1(n8213), .A2(n8212), .ZN(n14216) );
  NAND2_X1 U8090 ( .A1(n9605), .A2(n14106), .ZN(n14481) );
  AND2_X1 U8091 ( .A1(n9316), .A2(n13878), .ZN(n14154) );
  OR2_X1 U8092 ( .A1(n9606), .A2(n9604), .ZN(n14106) );
  NAND2_X1 U8093 ( .A1(n15339), .A2(n15340), .ZN(n15336) );
  NAND2_X1 U8094 ( .A1(n15338), .A2(n15336), .ZN(n15330) );
  INV_X1 U8095 ( .A(n7639), .ZN(n6984) );
  NAND2_X1 U8096 ( .A1(n14321), .A2(n15086), .ZN(n14320) );
  NAND2_X1 U8097 ( .A1(n7645), .A2(n7644), .ZN(n14526) );
  NAND2_X1 U8098 ( .A1(n14526), .A2(n14527), .ZN(n14523) );
  NAND2_X1 U8099 ( .A1(n6975), .A2(n6974), .ZN(n14525) );
  INV_X1 U8100 ( .A(n7644), .ZN(n6974) );
  INV_X1 U8101 ( .A(n7645), .ZN(n6975) );
  NAND2_X1 U8102 ( .A1(n14330), .A2(n6596), .ZN(n6791) );
  INV_X1 U8103 ( .A(n14311), .ZN(n6779) );
  NAND2_X1 U8104 ( .A1(n14330), .A2(n7652), .ZN(n14310) );
  INV_X1 U8105 ( .A(n6791), .ZN(n14309) );
  NAND2_X1 U8106 ( .A1(n12821), .A2(n12823), .ZN(n7313) );
  AOI21_X1 U8107 ( .B1(n8357), .B2(n9592), .A(n8376), .ZN(n7726) );
  AOI21_X1 U8108 ( .B1(n6683), .B2(n8376), .A(n7725), .ZN(n7730) );
  NAND2_X1 U8109 ( .A1(n6689), .A2(n7837), .ZN(n6688) );
  NAND2_X1 U8110 ( .A1(n7836), .A2(n7838), .ZN(n6689) );
  NAND2_X1 U8111 ( .A1(n7859), .A2(n7862), .ZN(n7348) );
  INV_X1 U8112 ( .A(n7881), .ZN(n6747) );
  OR2_X1 U8113 ( .A1(n7361), .A2(n7904), .ZN(n6874) );
  INV_X1 U8114 ( .A(n7903), .ZN(n7361) );
  OR2_X1 U8115 ( .A1(n7307), .A2(n12867), .ZN(n7306) );
  INV_X1 U8116 ( .A(n12866), .ZN(n7307) );
  NAND2_X1 U8117 ( .A1(n7944), .A2(n7946), .ZN(n6820) );
  AOI21_X1 U8118 ( .B1(n7326), .B2(n7324), .A(n7323), .ZN(n7322) );
  AND2_X1 U8119 ( .A1(n7327), .A2(n12878), .ZN(n7326) );
  INV_X1 U8120 ( .A(n12877), .ZN(n7327) );
  NAND2_X1 U8121 ( .A1(n7360), .A2(n7359), .ZN(n7358) );
  NOR2_X1 U8122 ( .A1(n7992), .A2(n7990), .ZN(n7360) );
  AND2_X1 U8123 ( .A1(n11455), .A2(n11414), .ZN(n8039) );
  NAND2_X1 U8124 ( .A1(n6588), .A2(n6756), .ZN(n6754) );
  INV_X1 U8125 ( .A(n7359), .ZN(n6756) );
  AND2_X1 U8126 ( .A1(n12894), .A2(n7304), .ZN(n6858) );
  NAND2_X1 U8127 ( .A1(n8098), .A2(n6803), .ZN(n6692) );
  NAND2_X1 U8128 ( .A1(n8141), .A2(n8142), .ZN(n8140) );
  NAND2_X1 U8129 ( .A1(n7308), .A2(n7309), .ZN(n12920) );
  NAND2_X1 U8130 ( .A1(n12915), .A2(n7310), .ZN(n7309) );
  NAND2_X1 U8131 ( .A1(n8177), .A2(n8176), .ZN(n6753) );
  INV_X1 U8132 ( .A(n8177), .ZN(n6695) );
  INV_X1 U8133 ( .A(n12920), .ZN(n6849) );
  OAI21_X1 U8134 ( .B1(n13439), .B2(n12997), .A(n7175), .ZN(n12975) );
  NAND2_X1 U8135 ( .A1(n13001), .A2(n12997), .ZN(n7175) );
  NAND2_X1 U8136 ( .A1(n7174), .A2(n7173), .ZN(n12974) );
  NAND2_X1 U8137 ( .A1(n13060), .A2(n12973), .ZN(n7173) );
  NAND2_X1 U8138 ( .A1(n13439), .A2(n12997), .ZN(n7174) );
  NAND2_X1 U8139 ( .A1(n8254), .A2(n7340), .ZN(n7339) );
  INV_X1 U8140 ( .A(n8253), .ZN(n7340) );
  OAI21_X1 U8141 ( .B1(n6869), .B2(n6870), .A(n7356), .ZN(n8235) );
  NAND2_X1 U8142 ( .A1(n7357), .A2(n8214), .ZN(n7356) );
  INV_X1 U8143 ( .A(n8234), .ZN(n6751) );
  NAND2_X1 U8144 ( .A1(n7694), .A2(n9511), .ZN(n8331) );
  OAI21_X1 U8145 ( .B1(n12925), .B2(n7319), .A(n6851), .ZN(n12929) );
  NOR2_X1 U8146 ( .A1(n12928), .A2(n6852), .ZN(n6851) );
  NAND2_X1 U8147 ( .A1(n7337), .A2(n12931), .ZN(n7336) );
  NOR2_X1 U8148 ( .A1(n7337), .A2(n12931), .ZN(n7338) );
  NOR2_X1 U8149 ( .A1(n8260), .A2(n12697), .ZN(n7194) );
  NAND2_X1 U8150 ( .A1(n8260), .A2(n12697), .ZN(n7195) );
  INV_X1 U8151 ( .A(n8247), .ZN(n7193) );
  INV_X1 U8152 ( .A(n7194), .ZN(n7192) );
  NOR2_X1 U8153 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n7662) );
  INV_X1 U8154 ( .A(n8073), .ZN(n7186) );
  INV_X1 U8155 ( .A(n6853), .ZN(n7559) );
  OAI21_X1 U8156 ( .B1(n7610), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6624), .ZN(
        n6853) );
  NOR2_X1 U8157 ( .A1(n11360), .A2(n7096), .ZN(n7095) );
  INV_X1 U8158 ( .A(n11262), .ZN(n7096) );
  NAND2_X1 U8159 ( .A1(n7091), .A2(n7094), .ZN(n7087) );
  AND2_X1 U8160 ( .A1(n7090), .A2(n7091), .ZN(n7089) );
  INV_X1 U8161 ( .A(n11488), .ZN(n7090) );
  OR2_X1 U8162 ( .A1(n9833), .A2(n9091), .ZN(n7052) );
  NAND2_X1 U8163 ( .A1(n7060), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7059) );
  OR2_X1 U8164 ( .A1(n10044), .A2(n6617), .ZN(n6996) );
  NOR2_X1 U8165 ( .A1(n12383), .A2(n7495), .ZN(n7494) );
  NAND2_X1 U8166 ( .A1(n7497), .A2(n11613), .ZN(n7495) );
  INV_X1 U8167 ( .A(n8942), .ZN(n7497) );
  NOR2_X1 U8168 ( .A1(n7038), .A2(n6541), .ZN(n7037) );
  NOR2_X1 U8169 ( .A1(n12383), .A2(n7499), .ZN(n7498) );
  INV_X1 U8170 ( .A(n7519), .ZN(n7517) );
  INV_X1 U8171 ( .A(n7520), .ZN(n7514) );
  INV_X1 U8172 ( .A(n11620), .ZN(n7513) );
  OR2_X1 U8173 ( .A1(n11623), .A2(n7029), .ZN(n7028) );
  INV_X1 U8174 ( .A(n8830), .ZN(n7029) );
  NAND2_X1 U8175 ( .A1(n8671), .A2(n6603), .ZN(n11060) );
  NAND2_X1 U8176 ( .A1(n11791), .A2(n11789), .ZN(n7473) );
  OR2_X1 U8177 ( .A1(n12202), .A2(n10850), .ZN(n11673) );
  AND2_X1 U8178 ( .A1(n10421), .A2(n8927), .ZN(n6765) );
  NAND2_X1 U8179 ( .A1(n6823), .A2(n14941), .ZN(n11629) );
  INV_X1 U8180 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8426) );
  INV_X1 U8181 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8905) );
  NOR2_X1 U8182 ( .A1(n6544), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8907) );
  INV_X1 U8183 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8421) );
  INV_X1 U8184 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8420) );
  INV_X1 U8185 ( .A(n8467), .ZN(n7464) );
  INV_X1 U8186 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U8187 ( .A1(n8461), .A2(n8460), .ZN(n8463) );
  OAI21_X1 U8188 ( .B1(n7459), .B2(n7458), .A(n8457), .ZN(n7457) );
  INV_X1 U8189 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8416) );
  INV_X1 U8190 ( .A(n11986), .ZN(n7276) );
  XNOR2_X1 U8191 ( .A(n13493), .B(n7249), .ZN(n11891) );
  NOR2_X1 U8192 ( .A1(n12716), .A2(n11853), .ZN(n7248) );
  INV_X1 U8193 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9010) );
  AND2_X1 U8194 ( .A1(n11902), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n11918) );
  NOR2_X1 U8195 ( .A1(n13343), .A2(n13482), .ZN(n7230) );
  OAI21_X1 U8196 ( .B1(n7163), .B2(n6543), .A(n13353), .ZN(n7162) );
  INV_X1 U8197 ( .A(n13159), .ZN(n7118) );
  INV_X1 U8198 ( .A(n7120), .ZN(n7115) );
  INV_X1 U8199 ( .A(n13178), .ZN(n7168) );
  AND2_X1 U8200 ( .A1(n13027), .A2(n13413), .ZN(n7142) );
  NAND2_X1 U8201 ( .A1(n13322), .A2(n13190), .ZN(n13308) );
  NOR2_X1 U8202 ( .A1(n13373), .A2(n13493), .ZN(n13359) );
  NAND2_X1 U8203 ( .A1(n7238), .A2(n7237), .ZN(n13373) );
  NAND2_X1 U8204 ( .A1(n10114), .A2(n10115), .ZN(n10113) );
  OR2_X1 U8205 ( .A1(n9575), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n9712) );
  OR2_X1 U8206 ( .A1(n9154), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U8207 ( .A1(n6682), .A2(n6681), .ZN(n9690) );
  NAND2_X1 U8208 ( .A1(n6878), .A2(n10415), .ZN(n6681) );
  INV_X1 U8209 ( .A(n11023), .ZN(n7398) );
  INV_X1 U8210 ( .A(n7378), .ZN(n7376) );
  NAND2_X1 U8211 ( .A1(n8336), .A2(n8335), .ZN(n7362) );
  NAND2_X1 U8212 ( .A1(n7346), .A2(n8295), .ZN(n7345) );
  AOI21_X1 U8213 ( .B1(n8266), .B2(n8267), .A(n6813), .ZN(n6868) );
  INV_X1 U8214 ( .A(n11594), .ZN(n6970) );
  NOR2_X1 U8215 ( .A1(n14074), .A2(n14216), .ZN(n7015) );
  NAND2_X1 U8216 ( .A1(n11455), .A2(n11460), .ZN(n6955) );
  NOR2_X1 U8217 ( .A1(n6540), .A2(n10627), .ZN(n6944) );
  NOR2_X1 U8218 ( .A1(n10945), .A2(n6947), .ZN(n6946) );
  INV_X1 U8219 ( .A(n10784), .ZN(n6947) );
  INV_X1 U8220 ( .A(n10618), .ZN(n7405) );
  NOR2_X1 U8221 ( .A1(n7405), .A2(n7404), .ZN(n7403) );
  INV_X1 U8222 ( .A(n10616), .ZN(n7404) );
  INV_X1 U8223 ( .A(n14004), .ZN(n13772) );
  INV_X1 U8224 ( .A(n8290), .ZN(n6800) );
  INV_X1 U8225 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7706) );
  AND2_X1 U8226 ( .A1(n7685), .A2(n7693), .ZN(n7367) );
  AND2_X1 U8227 ( .A1(n6705), .A2(n6706), .ZN(n7685) );
  NOR2_X1 U8228 ( .A1(n8085), .A2(SI_17_), .ZN(n6729) );
  AOI21_X1 U8229 ( .B1(n6626), .B2(n7545), .A(n6560), .ZN(n7187) );
  INV_X1 U8230 ( .A(n7545), .ZN(n7188) );
  AND2_X1 U8231 ( .A1(n7177), .A2(n6726), .ZN(n6725) );
  NAND2_X1 U8232 ( .A1(n7179), .A2(n7917), .ZN(n6726) );
  AOI21_X1 U8233 ( .B1(n7179), .B2(n7181), .A(n6612), .ZN(n7177) );
  XNOR2_X1 U8234 ( .A(n7996), .B(SI_13_), .ZN(n7993) );
  OR2_X1 U8235 ( .A1(n7854), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n7878) );
  OAI21_X1 U8236 ( .B1(n6967), .B2(n9156), .A(n6724), .ZN(n6723) );
  NAND2_X1 U8237 ( .A1(n7780), .A2(n7779), .ZN(n7793) );
  INV_X1 U8238 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7666) );
  OAI21_X1 U8239 ( .B1(n6536), .B2(n9347), .A(n6968), .ZN(n7711) );
  NAND2_X1 U8240 ( .A1(n6535), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6968) );
  XNOR2_X1 U8241 ( .A(n7558), .B(n7557), .ZN(n7610) );
  AOI22_X1 U8242 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n7579), .B1(n7596), .B2(
        n7578), .ZN(n7646) );
  INV_X1 U8243 ( .A(n14538), .ZN(n6783) );
  INV_X1 U8244 ( .A(n7095), .ZN(n7094) );
  AOI21_X1 U8245 ( .B1(n7093), .B2(n7095), .A(n7092), .ZN(n7091) );
  INV_X1 U8246 ( .A(n11359), .ZN(n7092) );
  INV_X1 U8247 ( .A(n11245), .ZN(n7093) );
  NAND2_X1 U8248 ( .A1(n8642), .A2(n8641), .ZN(n8658) );
  XNOR2_X1 U8249 ( .A(n10229), .B(n6517), .ZN(n10320) );
  NOR2_X1 U8250 ( .A1(n12108), .A2(n7070), .ZN(n7069) );
  INV_X1 U8251 ( .A(n12029), .ZN(n7070) );
  NOR2_X1 U8252 ( .A1(n8824), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8844) );
  OAI21_X1 U8253 ( .B1(n12141), .B2(n12118), .A(n12117), .ZN(n12116) );
  OR2_X1 U8254 ( .A1(n8502), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U8255 ( .A1(n11244), .A2(n11245), .ZN(n11263) );
  OAI21_X1 U8256 ( .B1(n10845), .B2(n7080), .A(n7078), .ZN(n11125) );
  AND2_X1 U8257 ( .A1(n7079), .A2(n11123), .ZN(n7078) );
  OR2_X1 U8258 ( .A1(n7081), .A2(n7080), .ZN(n7079) );
  NOR2_X1 U8259 ( .A1(n11816), .A2(n7470), .ZN(n11818) );
  NAND2_X1 U8260 ( .A1(n11825), .A2(n7471), .ZN(n7470) );
  OR2_X1 U8261 ( .A1(n6537), .A2(n14925), .ZN(n8543) );
  OR2_X1 U8262 ( .A1(n8540), .A2(n9998), .ZN(n8510) );
  AND3_X1 U8263 ( .A1(n6796), .A2(n8525), .A3(n8526), .ZN(n8529) );
  OR2_X1 U8264 ( .A1(n6518), .A2(n8523), .ZN(n6796) );
  NAND2_X1 U8265 ( .A1(n9664), .A2(n9085), .ZN(n9718) );
  AND2_X1 U8266 ( .A1(n9807), .A2(n9093), .ZN(n9096) );
  XNOR2_X1 U8267 ( .A(n6996), .B(n10049), .ZN(n10046) );
  NAND2_X1 U8268 ( .A1(n6831), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7044) );
  INV_X1 U8269 ( .A(n10032), .ZN(n6831) );
  NAND2_X1 U8270 ( .A1(n6994), .A2(n6993), .ZN(n6992) );
  NAND2_X1 U8271 ( .A1(n10487), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6993) );
  AND2_X1 U8272 ( .A1(n11082), .A2(n11081), .ZN(n11083) );
  INV_X1 U8273 ( .A(n6830), .ZN(n11076) );
  INV_X1 U8274 ( .A(n6829), .ZN(n12209) );
  AND2_X1 U8275 ( .A1(n12235), .A2(n12234), .ZN(n12236) );
  NAND2_X1 U8276 ( .A1(n7042), .A2(n12246), .ZN(n12262) );
  NOR2_X1 U8277 ( .A1(n12278), .A2(n12279), .ZN(n12284) );
  NAND2_X1 U8278 ( .A1(n12255), .A2(n12256), .ZN(n12276) );
  AND2_X1 U8279 ( .A1(n6985), .A2(n6591), .ZN(n12295) );
  NAND2_X1 U8280 ( .A1(n12294), .A2(n12310), .ZN(n6985) );
  NAND2_X1 U8281 ( .A1(n12295), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U8282 ( .A1(n7037), .A2(n12382), .ZN(n7034) );
  AOI21_X1 U8283 ( .B1(n7038), .B2(n6541), .A(n14949), .ZN(n7035) );
  NAND2_X1 U8284 ( .A1(n7038), .A2(n12383), .ZN(n7036) );
  AND2_X1 U8285 ( .A1(n12381), .A2(n12382), .ZN(n6825) );
  AOI21_X1 U8286 ( .B1(n12431), .B2(n8940), .A(n6582), .ZN(n12420) );
  AND2_X1 U8287 ( .A1(n11616), .A2(n12418), .ZN(n12430) );
  OAI21_X1 U8288 ( .B1(n7026), .B2(n7028), .A(n11622), .ZN(n12455) );
  INV_X1 U8289 ( .A(n12478), .ZN(n7026) );
  AND4_X1 U8290 ( .A1(n8801), .A2(n8800), .A3(n8799), .A4(n8798), .ZN(n12494)
         );
  NOR2_X1 U8291 ( .A1(n11806), .A2(n6769), .ZN(n6768) );
  INV_X1 U8292 ( .A(n8790), .ZN(n6769) );
  INV_X1 U8293 ( .A(n7505), .ZN(n7504) );
  AND2_X1 U8294 ( .A1(n7503), .A2(n11802), .ZN(n7502) );
  AND2_X1 U8295 ( .A1(n11709), .A2(n11708), .ZN(n12541) );
  NOR2_X1 U8296 ( .A1(n8763), .A2(n8411), .ZN(n8783) );
  INV_X1 U8297 ( .A(n6761), .ZN(n6760) );
  NOR2_X1 U8298 ( .A1(n8702), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8714) );
  AND2_X1 U8299 ( .A1(n11691), .A2(n11688), .ZN(n11799) );
  NAND2_X1 U8300 ( .A1(n7482), .A2(n7483), .ZN(n11323) );
  AOI21_X1 U8301 ( .B1(n7485), .B2(n11677), .A(n7484), .ZN(n7483) );
  INV_X1 U8302 ( .A(n11682), .ZN(n7484) );
  OR2_X1 U8303 ( .A1(n8658), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8684) );
  OR2_X1 U8304 ( .A1(n8684), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8702) );
  INV_X1 U8305 ( .A(n11130), .ZN(n14378) );
  AND2_X1 U8306 ( .A1(n8627), .A2(n10154), .ZN(n8642) );
  NAND2_X1 U8307 ( .A1(n7481), .A2(n7479), .ZN(n10962) );
  NAND2_X1 U8308 ( .A1(n10907), .A2(n6664), .ZN(n7481) );
  OR2_X1 U8309 ( .A1(n8593), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8611) );
  NOR2_X1 U8310 ( .A1(n8611), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8627) );
  INV_X1 U8311 ( .A(n10871), .ZN(n11794) );
  NAND2_X1 U8312 ( .A1(n10907), .A2(n11791), .ZN(n10906) );
  AND3_X1 U8313 ( .A1(n8609), .A2(n8608), .A3(n8607), .ZN(n10916) );
  INV_X1 U8314 ( .A(n10434), .ZN(n11793) );
  NOR2_X1 U8315 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8577) );
  INV_X1 U8316 ( .A(n8927), .ZN(n14908) );
  NAND2_X1 U8317 ( .A1(n11641), .A2(n11646), .ZN(n10421) );
  OR2_X1 U8318 ( .A1(n6529), .A2(n12697), .ZN(n8867) );
  NAND2_X1 U8319 ( .A1(n8857), .A2(n8856), .ZN(n12041) );
  INV_X1 U8320 ( .A(n12617), .ZN(n15011) );
  AND2_X1 U8321 ( .A1(n8947), .A2(n8996), .ZN(n14967) );
  NOR2_X1 U8322 ( .A1(n13566), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7443) );
  AOI21_X1 U8323 ( .B1(n7447), .B2(n7446), .A(n6673), .ZN(n7445) );
  NAND2_X1 U8324 ( .A1(n8485), .A2(n8484), .ZN(n8879) );
  NAND2_X1 U8325 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n8483), .ZN(n8484) );
  NAND2_X1 U8326 ( .A1(n8866), .A2(n8864), .ZN(n8485) );
  NOR2_X1 U8327 ( .A1(n7077), .A2(n7076), .ZN(n7075) );
  NOR2_X1 U8328 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7076) );
  NAND2_X1 U8329 ( .A1(n7429), .A2(n8481), .ZN(n8855) );
  NAND2_X1 U8330 ( .A1(n8497), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7429) );
  INV_X1 U8331 ( .A(n8820), .ZN(n7468) );
  NOR2_X1 U8332 ( .A1(n8618), .A2(n8418), .ZN(n8697) );
  AND2_X1 U8333 ( .A1(n8456), .A2(n8455), .ZN(n8665) );
  AOI21_X1 U8334 ( .B1(n7453), .B2(n7451), .A(n6628), .ZN(n7450) );
  INV_X1 U8335 ( .A(n7453), .ZN(n7452) );
  NAND2_X1 U8336 ( .A1(n8586), .A2(n8450), .ZN(n8601) );
  NAND2_X1 U8337 ( .A1(n6937), .A2(n11524), .ZN(n6930) );
  NAND2_X1 U8338 ( .A1(n7254), .A2(n11524), .ZN(n6934) );
  XNOR2_X1 U8339 ( .A(n12000), .B(n7249), .ZN(n12001) );
  NOR2_X1 U8340 ( .A1(n6567), .A2(n7276), .ZN(n7275) );
  INV_X1 U8341 ( .A(n12753), .ZN(n7246) );
  NOR2_X1 U8342 ( .A1(n10290), .A2(n10289), .ZN(n10508) );
  OR2_X1 U8343 ( .A1(n10064), .A2(n10296), .ZN(n10290) );
  INV_X1 U8344 ( .A(n6917), .ZN(n6916) );
  OAI21_X1 U8345 ( .B1(n7248), .B2(n6918), .A(n12762), .ZN(n6917) );
  INV_X1 U8346 ( .A(n12763), .ZN(n6918) );
  NAND2_X1 U8347 ( .A1(n12778), .A2(n7248), .ZN(n12765) );
  XNOR2_X1 U8348 ( .A(n14658), .B(n7249), .ZN(n11523) );
  INV_X1 U8349 ( .A(n9356), .ZN(n6920) );
  NAND2_X1 U8350 ( .A1(n11550), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n11874) );
  AND2_X1 U8351 ( .A1(n12948), .A2(n13000), .ZN(n7300) );
  NAND2_X1 U8352 ( .A1(n6799), .A2(n6798), .ZN(n12990) );
  NAND2_X1 U8353 ( .A1(n9331), .A2(n6859), .ZN(n10076) );
  INV_X1 U8354 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8355 ( .A1(n9331), .A2(n7543), .ZN(n10637) );
  NOR2_X1 U8356 ( .A1(n13140), .A2(n7232), .ZN(n7231) );
  INV_X1 U8357 ( .A(n7233), .ZN(n7232) );
  INV_X1 U8358 ( .A(n7151), .ZN(n7150) );
  AOI21_X1 U8359 ( .B1(n7107), .B2(n7106), .A(n6599), .ZN(n7105) );
  INV_X1 U8360 ( .A(n7110), .ZN(n7106) );
  NAND2_X1 U8361 ( .A1(n7230), .A2(n7229), .ZN(n13302) );
  INV_X1 U8362 ( .A(n7230), .ZN(n13324) );
  INV_X1 U8363 ( .A(n7117), .ZN(n7116) );
  AOI21_X1 U8364 ( .B1(n7115), .B2(n7117), .A(n6614), .ZN(n7114) );
  NOR2_X1 U8365 ( .A1(n13161), .A2(n7118), .ZN(n7117) );
  NAND2_X1 U8366 ( .A1(n6847), .A2(n6846), .ZN(n13401) );
  AND2_X1 U8367 ( .A1(n11559), .A2(n13403), .ZN(n7124) );
  NOR2_X1 U8368 ( .A1(n11388), .A2(n11387), .ZN(n11395) );
  OR2_X1 U8369 ( .A1(n11222), .A2(n14658), .ZN(n11443) );
  AND2_X1 U8370 ( .A1(n7155), .A2(n11373), .ZN(n7154) );
  NAND2_X1 U8371 ( .A1(n11143), .A2(n11231), .ZN(n11222) );
  OAI21_X1 U8372 ( .B1(n11150), .B2(n11149), .A(n11148), .ZN(n11211) );
  NAND2_X1 U8373 ( .A1(n7242), .A2(n10802), .ZN(n11002) );
  INV_X1 U8374 ( .A(n7243), .ZN(n7242) );
  AND2_X1 U8375 ( .A1(n7139), .A2(n10995), .ZN(n7138) );
  NAND2_X1 U8376 ( .A1(n10801), .A2(n10767), .ZN(n10769) );
  NAND2_X1 U8377 ( .A1(n10802), .A2(n10812), .ZN(n10805) );
  NOR2_X1 U8378 ( .A1(n9858), .A2(n9857), .ZN(n9971) );
  NOR2_X2 U8379 ( .A1(n10217), .A2(n14835), .ZN(n10527) );
  NAND2_X1 U8380 ( .A1(n7206), .A2(n7205), .ZN(n10217) );
  INV_X1 U8381 ( .A(n10215), .ZN(n7206) );
  XNOR2_X1 U8382 ( .A(n13073), .B(n6522), .ZN(n13008) );
  INV_X1 U8383 ( .A(n13008), .ZN(n9908) );
  NAND2_X1 U8384 ( .A1(n10125), .A2(n6522), .ZN(n9915) );
  NAND2_X1 U8385 ( .A1(n7129), .A2(n9871), .ZN(n9936) );
  CLKBUF_X1 U8386 ( .A(n9875), .Z(n10205) );
  NAND2_X1 U8387 ( .A1(n14297), .A2(n12963), .ZN(n6797) );
  NAND2_X1 U8388 ( .A1(n7145), .A2(n11544), .ZN(n13404) );
  NAND2_X1 U8389 ( .A1(n11543), .A2(n13027), .ZN(n7145) );
  INV_X1 U8390 ( .A(n13529), .ZN(n14833) );
  AND2_X1 U8391 ( .A1(n10205), .A2(n14822), .ZN(n13529) );
  NOR2_X1 U8392 ( .A1(n6575), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U8393 ( .A1(n7286), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9332) );
  NOR2_X1 U8394 ( .A1(n9157), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9165) );
  NOR2_X2 U8395 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9110) );
  INV_X1 U8396 ( .A(n13795), .ZN(n6893) );
  INV_X1 U8397 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7906) );
  OR2_X1 U8398 ( .A1(n9951), .A2(n9950), .ZN(n9952) );
  INV_X1 U8399 ( .A(n13745), .ZN(n6901) );
  INV_X1 U8400 ( .A(n6904), .ZN(n6903) );
  OAI21_X1 U8401 ( .B1(n7382), .B2(n6905), .A(n6906), .ZN(n6904) );
  NAND2_X1 U8402 ( .A1(n13736), .A2(n13735), .ZN(n6906) );
  NOR2_X1 U8403 ( .A1(n7840), .A2(n7839), .ZN(n7863) );
  NAND2_X1 U8404 ( .A1(n6876), .A2(n9695), .ZN(n9696) );
  OR2_X1 U8405 ( .A1(n9694), .A2(n7544), .ZN(n9695) );
  NAND2_X1 U8406 ( .A1(n8067), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U8407 ( .A1(n7399), .A2(n7398), .ZN(n11156) );
  INV_X1 U8408 ( .A(n11022), .ZN(n7399) );
  NAND2_X1 U8409 ( .A1(n6912), .A2(n6911), .ZN(n6910) );
  INV_X1 U8410 ( .A(n11155), .ZN(n6911) );
  INV_X1 U8411 ( .A(n13594), .ZN(n7389) );
  INV_X1 U8412 ( .A(n7392), .ZN(n7391) );
  AND2_X1 U8413 ( .A1(n8148), .A2(n8147), .ZN(n8162) );
  NAND2_X1 U8414 ( .A1(n13804), .A2(n13805), .ZN(n13803) );
  OR2_X1 U8415 ( .A1(n7907), .A2(n7906), .ZN(n7931) );
  AND2_X1 U8416 ( .A1(n8378), .A2(n8377), .ZN(n8386) );
  INV_X1 U8417 ( .A(n8269), .ZN(n8319) );
  OR2_X1 U8419 ( .A1(n7878), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U8420 ( .A1(n14189), .A2(n14003), .ZN(n7219) );
  AOI21_X1 U8421 ( .B1(n7215), .B2(n7218), .A(n6611), .ZN(n7213) );
  NAND2_X1 U8422 ( .A1(n7215), .A2(n7211), .ZN(n7210) );
  AND2_X1 U8423 ( .A1(n7219), .A2(n7212), .ZN(n7211) );
  INV_X1 U8424 ( .A(n11595), .ZN(n7212) );
  NAND2_X1 U8425 ( .A1(n8313), .A2(n8312), .ZN(n13985) );
  AOI21_X1 U8426 ( .B1(n13582), .B2(n14012), .A(n14001), .ZN(n11583) );
  XNOR2_X1 U8427 ( .A(n6942), .B(n11596), .ZN(n6941) );
  AOI21_X1 U8428 ( .B1(n7221), .B2(n7217), .A(n7214), .ZN(n6942) );
  NAND2_X1 U8429 ( .A1(n8238), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U8430 ( .A1(n7221), .A2(n6579), .ZN(n14006) );
  NAND2_X1 U8431 ( .A1(n14070), .A2(n6551), .ZN(n14037) );
  INV_X1 U8432 ( .A(n6972), .ZN(n6971) );
  AOI21_X1 U8433 ( .B1(n14068), .B2(n7223), .A(n6619), .ZN(n7222) );
  INV_X1 U8434 ( .A(n8196), .ZN(n8197) );
  NAND2_X1 U8435 ( .A1(n7225), .A2(n7223), .ZN(n14052) );
  NOR2_X1 U8436 ( .A1(n14081), .A2(n14082), .ZN(n14080) );
  NOR2_X1 U8437 ( .A1(n14099), .A2(n14228), .ZN(n14070) );
  NAND2_X1 U8438 ( .A1(n14070), .A2(n11600), .ZN(n14071) );
  AND2_X1 U8439 ( .A1(n14228), .A2(n13718), .ZN(n11590) );
  OR2_X1 U8440 ( .A1(n14069), .A2(n14068), .ZN(n7225) );
  XNOR2_X1 U8441 ( .A(n14090), .B(n14105), .ZN(n14087) );
  NOR3_X1 U8442 ( .A1(n11477), .A2(n7011), .A3(n14244), .ZN(n14101) );
  INV_X1 U8443 ( .A(n7201), .ZN(n7200) );
  NAND2_X1 U8444 ( .A1(n6548), .A2(n6964), .ZN(n6960) );
  NAND2_X1 U8445 ( .A1(n11586), .A2(n6548), .ZN(n6961) );
  AOI21_X1 U8446 ( .B1(n7417), .B2(n7414), .A(n7412), .ZN(n14127) );
  AND2_X1 U8447 ( .A1(n14133), .A2(n7415), .ZN(n7414) );
  NAND2_X1 U8448 ( .A1(n7413), .A2(n6613), .ZN(n7412) );
  NAND2_X1 U8449 ( .A1(n6957), .A2(n6958), .ZN(n11457) );
  NAND2_X1 U8450 ( .A1(n14436), .A2(n6793), .ZN(n6792) );
  OR2_X1 U8451 ( .A1(n8012), .A2(n8011), .ZN(n8029) );
  NOR2_X1 U8452 ( .A1(n13610), .A2(n13846), .ZN(n11300) );
  NAND2_X1 U8453 ( .A1(n11311), .A2(n11310), .ZN(n11416) );
  NOR2_X1 U8454 ( .A1(n7931), .A2(n7930), .ZN(n7948) );
  NAND2_X1 U8455 ( .A1(n7017), .A2(n7016), .ZN(n11200) );
  INV_X1 U8456 ( .A(n11111), .ZN(n7017) );
  NAND2_X1 U8457 ( .A1(n7019), .A2(n7018), .ZN(n11111) );
  INV_X1 U8458 ( .A(n6945), .ZN(n11104) );
  AOI21_X1 U8459 ( .B1(n10785), .B2(n6946), .A(n6540), .ZN(n6945) );
  NOR2_X1 U8460 ( .A1(n10662), .A2(n14616), .ZN(n10790) );
  INV_X1 U8461 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7886) );
  OR2_X1 U8462 ( .A1(n7887), .A2(n7886), .ZN(n7907) );
  OAI21_X1 U8463 ( .B1(n10622), .B2(n10621), .A(n10623), .ZN(n10667) );
  NAND2_X1 U8464 ( .A1(n10617), .A2(n10616), .ZN(n10660) );
  NAND2_X1 U8465 ( .A1(n10555), .A2(n10554), .ZN(n10617) );
  AND2_X1 U8466 ( .A1(n10603), .A2(n10574), .ZN(n10561) );
  AND2_X1 U8467 ( .A1(n10453), .A2(n14591), .ZN(n7013) );
  NAND2_X1 U8468 ( .A1(n10386), .A2(n14591), .ZN(n10385) );
  AND4_X1 U8469 ( .A1(n7775), .A2(n7774), .A3(n7773), .A4(n7772), .ZN(n10585)
         );
  OR2_X1 U8470 ( .A1(n13859), .A2(n10415), .ZN(n10010) );
  INV_X1 U8471 ( .A(n10020), .ZN(n7204) );
  NOR2_X1 U8472 ( .A1(n10020), .A2(n10019), .ZN(n10363) );
  INV_X1 U8473 ( .A(n14154), .ZN(n14136) );
  OR2_X1 U8474 ( .A1(n9588), .A2(n13878), .ZN(n14138) );
  OR3_X1 U8475 ( .A1(n10308), .A2(n10307), .A3(n10306), .ZN(n13989) );
  OR2_X1 U8476 ( .A1(n9587), .A2(n9586), .ZN(n14609) );
  NAND2_X1 U8477 ( .A1(n9595), .A2(n9175), .ZN(n9604) );
  AND3_X1 U8478 ( .A1(n8022), .A2(n7410), .A3(n7670), .ZN(n7674) );
  AND2_X1 U8479 ( .A1(n6555), .A2(n7672), .ZN(n7410) );
  INV_X1 U8480 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7675) );
  XNOR2_X1 U8481 ( .A(n8286), .B(n8262), .ZN(n13576) );
  XNOR2_X1 U8482 ( .A(n8261), .B(n8250), .ZN(n11967) );
  NAND2_X1 U8483 ( .A1(n7196), .A2(n8249), .ZN(n8261) );
  OR2_X1 U8484 ( .A1(n8248), .A2(n8247), .ZN(n7196) );
  INV_X1 U8485 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U8486 ( .A1(n8025), .A2(n7685), .ZN(n8089) );
  XNOR2_X1 U8487 ( .A(n8021), .B(n8051), .ZN(n11383) );
  NAND2_X1 U8488 ( .A1(n7178), .A2(n7956), .ZN(n7978) );
  NAND2_X1 U8489 ( .A1(n7937), .A2(n7182), .ZN(n7178) );
  NAND2_X1 U8490 ( .A1(n7937), .A2(n7936), .ZN(n7958) );
  NAND2_X1 U8491 ( .A1(n7170), .A2(n6837), .ZN(n7898) );
  AOI21_X1 U8492 ( .B1(n7171), .B2(n7172), .A(n7169), .ZN(n6837) );
  NAND2_X1 U8493 ( .A1(n7171), .A2(n7852), .ZN(n7170) );
  INV_X1 U8494 ( .A(n7893), .ZN(n7169) );
  OAI21_X1 U8495 ( .B1(n7900), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7940) );
  INV_X1 U8496 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n9679) );
  XNOR2_X1 U8497 ( .A(n7622), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n7624) );
  NAND2_X1 U8498 ( .A1(n6977), .A2(n6598), .ZN(n6976) );
  NOR2_X1 U8499 ( .A1(n7565), .A2(n7564), .ZN(n7628) );
  AND2_X1 U8500 ( .A1(n9568), .A2(n7622), .ZN(n7564) );
  NOR2_X1 U8501 ( .A1(n14317), .A2(n7630), .ZN(n7633) );
  AOI21_X1 U8502 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n7572), .A(n7571), .ZN(
        n7604) );
  NOR2_X1 U8503 ( .A1(n7636), .A2(n7637), .ZN(n7571) );
  NAND2_X1 U8504 ( .A1(n7601), .A2(n7575), .ZN(n7599) );
  NAND2_X1 U8505 ( .A1(n14327), .A2(n6816), .ZN(n6773) );
  NAND2_X1 U8506 ( .A1(n14328), .A2(n6776), .ZN(n6775) );
  NAND2_X1 U8507 ( .A1(n6777), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6776) );
  INV_X1 U8508 ( .A(n14327), .ZN(n6777) );
  AND2_X1 U8509 ( .A1(n6978), .A2(n14516), .ZN(n7642) );
  NAND2_X1 U8510 ( .A1(n6778), .A2(n6979), .ZN(n6978) );
  INV_X1 U8511 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6979) );
  NAND2_X1 U8512 ( .A1(n6775), .A2(n6609), .ZN(n6778) );
  AND2_X1 U8513 ( .A1(n14523), .A2(n14525), .ZN(n7649) );
  NAND2_X1 U8514 ( .A1(n6780), .A2(n6781), .ZN(n6784) );
  INV_X1 U8515 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6781) );
  INV_X1 U8516 ( .A(n14534), .ZN(n6786) );
  OR2_X1 U8517 ( .A1(n8884), .A2(n8413), .ZN(n12390) );
  OAI21_X1 U8518 ( .B1(n11244), .B2(n7094), .A(n7091), .ZN(n11489) );
  NAND2_X1 U8519 ( .A1(n12071), .A2(n11120), .ZN(n12072) );
  NAND2_X1 U8520 ( .A1(n8883), .A2(n8882), .ZN(n12102) );
  NAND2_X1 U8521 ( .A1(n8921), .A2(n10255), .ZN(n9990) );
  NAND2_X1 U8522 ( .A1(n12030), .A2(n12029), .ZN(n12107) );
  NAND2_X1 U8523 ( .A1(n11493), .A2(n11492), .ZN(n11495) );
  NAND2_X1 U8524 ( .A1(n10537), .A2(n10538), .ZN(n10858) );
  AND2_X1 U8525 ( .A1(n12019), .A2(n12018), .ZN(n12127) );
  NAND2_X1 U8526 ( .A1(n10845), .A2(n10844), .ZN(n10847) );
  NAND2_X1 U8527 ( .A1(n11263), .A2(n11262), .ZN(n11361) );
  OR2_X1 U8528 ( .A1(n9994), .A2(n9799), .ZN(n12192) );
  AND2_X1 U8529 ( .A1(n9787), .A2(n9786), .ZN(n14347) );
  NAND2_X1 U8530 ( .A1(n9796), .A2(n14926), .ZN(n14341) );
  INV_X1 U8531 ( .A(n12174), .ZN(n14343) );
  AND2_X1 U8532 ( .A1(n11770), .A2(n8902), .ZN(n12370) );
  AOI21_X1 U8533 ( .B1(n12375), .B2(n8897), .A(n8889), .ZN(n12387) );
  NAND2_X1 U8534 ( .A1(n8877), .A2(n8876), .ZN(n12415) );
  OR2_X1 U8535 ( .A1(n9662), .A2(n9034), .ZN(n9664) );
  INV_X1 U8536 ( .A(n7044), .ZN(n10132) );
  INV_X1 U8537 ( .A(n6678), .ZN(n10152) );
  INV_X1 U8538 ( .A(n6994), .ZN(n10484) );
  XNOR2_X1 U8539 ( .A(n6992), .B(n10488), .ZN(n10485) );
  XNOR2_X1 U8540 ( .A(n11083), .B(n6995), .ZN(n14864) );
  INV_X1 U8541 ( .A(n7063), .ZN(n14870) );
  INV_X1 U8542 ( .A(n7062), .ZN(n11079) );
  NAND2_X1 U8543 ( .A1(n12235), .A2(n6661), .ZN(n6986) );
  INV_X1 U8544 ( .A(n7042), .ZN(n12243) );
  INV_X1 U8545 ( .A(n7043), .ZN(n12213) );
  OR2_X1 U8546 ( .A1(n12244), .A2(n12610), .ZN(n7067) );
  NOR2_X1 U8547 ( .A1(n9099), .A2(n11834), .ZN(n12362) );
  NOR2_X1 U8548 ( .A1(n7020), .A2(n7024), .ZN(n12443) );
  NAND2_X1 U8549 ( .A1(n7518), .A2(n7519), .ZN(n12462) );
  NAND2_X1 U8550 ( .A1(n12486), .A2(n7520), .ZN(n7518) );
  NAND2_X1 U8551 ( .A1(n12478), .A2(n8830), .ZN(n12468) );
  NAND2_X1 U8552 ( .A1(n12486), .A2(n11626), .ZN(n12471) );
  NAND2_X1 U8553 ( .A1(n7492), .A2(n11712), .ZN(n12518) );
  AND2_X1 U8554 ( .A1(n8762), .A2(n8761), .ZN(n12547) );
  NAND2_X1 U8555 ( .A1(n7501), .A2(n7505), .ZN(n11511) );
  NAND2_X1 U8556 ( .A1(n14365), .A2(n7508), .ZN(n7501) );
  NAND2_X1 U8557 ( .A1(n7510), .A2(n11693), .ZN(n11428) );
  NAND2_X1 U8558 ( .A1(n7511), .A2(n11692), .ZN(n7510) );
  INV_X1 U8559 ( .A(n14365), .ZN(n7511) );
  NAND2_X1 U8560 ( .A1(n11320), .A2(n8708), .ZN(n14359) );
  NAND2_X1 U8561 ( .A1(n7487), .A2(n7489), .ZN(n14377) );
  NAND2_X1 U8562 ( .A1(n7488), .A2(n11062), .ZN(n7487) );
  INV_X1 U8563 ( .A(n8933), .ZN(n7488) );
  NAND2_X1 U8564 ( .A1(n14379), .A2(n14980), .ZN(n14354) );
  NAND2_X1 U8565 ( .A1(n8933), .A2(n11672), .ZN(n11067) );
  NAND2_X1 U8566 ( .A1(n10971), .A2(n10419), .ZN(n14380) );
  NAND2_X1 U8567 ( .A1(n6795), .A2(n8592), .ZN(n10912) );
  INV_X1 U8568 ( .A(n14926), .ZN(n14952) );
  AND2_X1 U8569 ( .A1(n14385), .A2(n14384), .ZN(n14404) );
  NAND2_X1 U8570 ( .A1(n11576), .A2(n8948), .ZN(n8991) );
  OR2_X1 U8571 ( .A1(n11570), .A2(n12617), .ZN(n8948) );
  INV_X1 U8572 ( .A(n12102), .ZN(n12620) );
  INV_X1 U8573 ( .A(n12047), .ZN(n12627) );
  INV_X1 U8574 ( .A(n12041), .ZN(n12631) );
  AND2_X1 U8575 ( .A1(n8499), .A2(n8498), .ZN(n12635) );
  AND2_X1 U8576 ( .A1(n8509), .A2(n8508), .ZN(n12639) );
  NAND2_X1 U8577 ( .A1(n8843), .A2(n8842), .ZN(n12642) );
  NAND2_X1 U8578 ( .A1(n8811), .A2(n8810), .ZN(n12655) );
  INV_X1 U8579 ( .A(n12547), .ZN(n12663) );
  AND2_X1 U8580 ( .A1(n8965), .A2(n8964), .ZN(n12672) );
  AND2_X1 U8581 ( .A1(n8962), .A2(n8961), .ZN(n12674) );
  AND2_X1 U8582 ( .A1(n9778), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12673) );
  NAND2_X1 U8583 ( .A1(n7444), .A2(n7442), .ZN(n11762) );
  AOI21_X1 U8584 ( .B1(n7445), .B2(n6671), .A(n7443), .ZN(n7442) );
  INV_X1 U8585 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12675) );
  NAND2_X1 U8586 ( .A1(n6516), .A2(n6595), .ZN(n12678) );
  NAND2_X1 U8587 ( .A1(n7441), .A2(n7445), .ZN(n11773) );
  NAND2_X1 U8588 ( .A1(n7449), .A2(n8892), .ZN(n11759) );
  XNOR2_X1 U8589 ( .A(n8891), .B(n7446), .ZN(n11605) );
  INV_X1 U8590 ( .A(n8976), .ZN(n12699) );
  INV_X1 U8591 ( .A(SI_20_), .ZN(n10112) );
  INV_X1 U8592 ( .A(n7469), .ZN(n8821) );
  OAI21_X1 U8593 ( .B1(n8752), .B2(n7435), .A(n7433), .ZN(n8791) );
  NAND2_X1 U8594 ( .A1(n8752), .A2(n8471), .ZN(n8774) );
  INV_X1 U8595 ( .A(SI_15_), .ZN(n9523) );
  NAND2_X1 U8596 ( .A1(n7465), .A2(n8467), .ZN(n8741) );
  NAND2_X1 U8597 ( .A1(n7467), .A2(n7466), .ZN(n7465) );
  INV_X1 U8598 ( .A(SI_11_), .ZN(n9161) );
  NAND2_X1 U8599 ( .A1(n8664), .A2(n8456), .ZN(n8678) );
  NAND2_X1 U8600 ( .A1(n8623), .A2(n8452), .ZN(n8638) );
  NAND2_X1 U8601 ( .A1(n8572), .A2(n8448), .ZN(n8588) );
  NAND2_X1 U8602 ( .A1(n8446), .A2(n8445), .ZN(n8570) );
  OR2_X1 U8603 ( .A1(n8584), .A2(n8429), .ZN(n8568) );
  NAND2_X1 U8604 ( .A1(n7047), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U8605 ( .A1(n8546), .A2(n8429), .ZN(n7045) );
  NAND2_X1 U8606 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8514) );
  NOR2_X1 U8607 ( .A1(n12700), .A2(n6926), .ZN(n6925) );
  INV_X1 U8608 ( .A(n11973), .ZN(n6926) );
  AOI21_X1 U8609 ( .B1(n12734), .B2(n6556), .A(n6924), .ZN(n6923) );
  OAI21_X1 U8610 ( .B1(n11984), .B2(n11973), .A(n14644), .ZN(n6924) );
  AND4_X1 U8611 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n14420) );
  NAND2_X1 U8612 ( .A1(n12778), .A2(n11854), .ZN(n12715) );
  NAND2_X1 U8613 ( .A1(n9354), .A2(n9524), .ZN(n9355) );
  NAND2_X1 U8614 ( .A1(n7261), .A2(n7263), .ZN(n7259) );
  NAND2_X1 U8615 ( .A1(n7261), .A2(n14638), .ZN(n7260) );
  NAND2_X1 U8616 ( .A1(n7277), .A2(n7283), .ZN(n7278) );
  NAND2_X1 U8617 ( .A1(n11933), .A2(n11932), .ZN(n13470) );
  AND2_X1 U8618 ( .A1(n9737), .A2(n9738), .ZN(n6815) );
  NAND2_X1 U8619 ( .A1(n6660), .A2(n7255), .ZN(n14654) );
  AND2_X1 U8620 ( .A1(n6929), .A2(n6935), .ZN(n14651) );
  NOR2_X1 U8621 ( .A1(n7254), .A2(n6937), .ZN(n6929) );
  AOI21_X1 U8622 ( .B1(n14638), .B2(n14637), .A(n7263), .ZN(n10884) );
  OR2_X1 U8623 ( .A1(n12740), .A2(n7280), .ZN(n7279) );
  INV_X1 U8624 ( .A(n11847), .ZN(n7280) );
  NOR2_X1 U8625 ( .A1(n9383), .A2(n13042), .ZN(n12783) );
  NAND2_X1 U8626 ( .A1(n12734), .A2(n11959), .ZN(n12788) );
  NAND4_X1 U8627 ( .A1(n9654), .A2(n9653), .A3(n9652), .A4(n9651), .ZN(n13072)
         );
  AND2_X1 U8628 ( .A1(n9338), .A2(n9339), .ZN(n9342) );
  OR2_X1 U8629 ( .A1(n13242), .A2(n13241), .ZN(n13457) );
  NAND2_X1 U8630 ( .A1(n7109), .A2(n7113), .ZN(n13248) );
  NAND2_X1 U8631 ( .A1(n7109), .A2(n7107), .ZN(n13453) );
  AOI21_X1 U8632 ( .B1(n13239), .B2(n14798), .A(n6840), .ZN(n13458) );
  NAND2_X1 U8633 ( .A1(n6842), .A2(n6841), .ZN(n6840) );
  NAND2_X1 U8634 ( .A1(n13238), .A2(n13405), .ZN(n6841) );
  NAND2_X1 U8635 ( .A1(n13170), .A2(n13169), .ZN(n13255) );
  NOR2_X1 U8636 ( .A1(n7133), .A2(n7132), .ZN(n13285) );
  INV_X1 U8637 ( .A(n13192), .ZN(n7132) );
  NAND2_X1 U8638 ( .A1(n13480), .A2(n13165), .ZN(n13301) );
  NAND2_X1 U8639 ( .A1(n13336), .A2(n13189), .ZN(n13317) );
  INV_X1 U8640 ( .A(n7160), .ZN(n13354) );
  AOI21_X1 U8641 ( .B1(n7165), .B2(n7163), .A(n6543), .ZN(n7160) );
  NAND2_X1 U8642 ( .A1(n7119), .A2(n13159), .ZN(n13352) );
  NAND2_X1 U8643 ( .A1(n13392), .A2(n7120), .ZN(n7119) );
  NAND2_X1 U8644 ( .A1(n7165), .A2(n13181), .ZN(n13367) );
  NAND2_X1 U8645 ( .A1(n13392), .A2(n13156), .ZN(n13372) );
  NAND2_X1 U8646 ( .A1(n13179), .A2(n13178), .ZN(n13382) );
  NAND2_X1 U8647 ( .A1(n11549), .A2(n11548), .ZN(n13509) );
  NAND2_X1 U8648 ( .A1(n7125), .A2(n11559), .ZN(n13414) );
  NAND2_X1 U8649 ( .A1(n7125), .A2(n7124), .ZN(n13516) );
  NAND2_X1 U8650 ( .A1(n11519), .A2(n11518), .ZN(n13514) );
  NAND2_X1 U8651 ( .A1(n11214), .A2(n13023), .ZN(n11374) );
  NAND2_X1 U8652 ( .A1(n11213), .A2(n11212), .ZN(n11214) );
  NAND2_X1 U8653 ( .A1(n10775), .A2(n13019), .ZN(n10996) );
  NAND2_X1 U8654 ( .A1(n10806), .A2(n10774), .ZN(n10775) );
  AND2_X1 U8655 ( .A1(n6731), .A2(n7134), .ZN(n10650) );
  NAND2_X1 U8656 ( .A1(n10642), .A2(n10641), .ZN(n10644) );
  NAND2_X1 U8657 ( .A1(n10524), .A2(n10523), .ZN(n10648) );
  OR2_X1 U8658 ( .A1(n9917), .A2(n13052), .ZN(n14789) );
  INV_X1 U8659 ( .A(n13390), .ZN(n14785) );
  INV_X1 U8660 ( .A(n13141), .ZN(n13533) );
  AND2_X1 U8661 ( .A1(n9388), .A2(n9357), .ZN(n14817) );
  INV_X1 U8662 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U8663 ( .A1(n7329), .A2(n9318), .ZN(n7328) );
  INV_X1 U8664 ( .A(n7331), .ZN(n7329) );
  INV_X1 U8665 ( .A(n9323), .ZN(n13569) );
  NAND2_X1 U8666 ( .A1(n9019), .A2(n7234), .ZN(n6741) );
  AND2_X1 U8667 ( .A1(n6583), .A2(n7332), .ZN(n7234) );
  XNOR2_X1 U8668 ( .A(n9027), .B(n7332), .ZN(n11453) );
  INV_X1 U8669 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n15291) );
  INV_X1 U8670 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15205) );
  INV_X1 U8671 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11869) );
  INV_X1 U8672 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n15116) );
  NAND2_X1 U8673 ( .A1(n9331), .A2(n7287), .ZN(n9335) );
  AND2_X1 U8674 ( .A1(n7543), .A2(n7288), .ZN(n7287) );
  INV_X1 U8675 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10244) );
  INV_X1 U8676 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10081) );
  INV_X1 U8677 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9822) );
  INV_X1 U8678 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9577) );
  INV_X1 U8679 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9308) );
  INV_X1 U8680 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10496) );
  OR2_X1 U8681 ( .A1(n9288), .A2(n9287), .ZN(n14705) );
  INV_X1 U8682 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9209) );
  INV_X1 U8683 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9167) );
  INV_X1 U8684 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9148) );
  INV_X1 U8685 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9641) );
  INV_X1 U8686 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9526) );
  OAI21_X1 U8687 ( .B1(n7390), .B2(n6893), .A(n6890), .ZN(n14432) );
  NAND2_X1 U8688 ( .A1(n13803), .A2(n13679), .ZN(n13716) );
  AND2_X1 U8689 ( .A1(n6907), .A2(n6552), .ZN(n11347) );
  NAND2_X1 U8690 ( .A1(n9953), .A2(n9952), .ZN(n9956) );
  INV_X1 U8691 ( .A(n14103), .ZN(n14137) );
  NAND2_X1 U8692 ( .A1(n7396), .A2(n13655), .ZN(n13725) );
  NAND2_X1 U8693 ( .A1(n11020), .A2(n11019), .ZN(n11022) );
  NAND2_X1 U8694 ( .A1(n13786), .A2(n13666), .ZN(n13753) );
  NAND2_X1 U8695 ( .A1(n14477), .A2(n13599), .ZN(n13761) );
  NAND2_X1 U8696 ( .A1(n14477), .A2(n7392), .ZN(n13762) );
  AND2_X1 U8697 ( .A1(n7373), .A2(n7380), .ZN(n10602) );
  NAND2_X1 U8698 ( .A1(n7371), .A2(n10337), .ZN(n7380) );
  OR2_X1 U8699 ( .A1(n9845), .A2(n6531), .ZN(n7804) );
  AOI21_X1 U8700 ( .B1(n6885), .B2(n6887), .A(n6608), .ZN(n6884) );
  OAI211_X1 U8701 ( .C1(n10194), .C2(n10337), .A(n7378), .B(n7374), .ZN(n10339) );
  NAND2_X1 U8702 ( .A1(n10194), .A2(n6578), .ZN(n7374) );
  AND2_X1 U8703 ( .A1(n11156), .A2(n11155), .ZN(n11161) );
  NAND2_X1 U8704 ( .A1(n6907), .A2(n6910), .ZN(n11340) );
  NOR2_X1 U8705 ( .A1(n13808), .A2(n14138), .ZN(n14457) );
  NAND2_X1 U8706 ( .A1(n13796), .A2(n13795), .ZN(n14430) );
  NAND2_X1 U8707 ( .A1(n7390), .A2(n7388), .ZN(n13796) );
  INV_X1 U8708 ( .A(n14228), .ZN(n14090) );
  NAND2_X1 U8709 ( .A1(n13595), .A2(n13594), .ZN(n14477) );
  INV_X1 U8710 ( .A(n13857), .ZN(n10365) );
  OR2_X1 U8711 ( .A1(n9600), .A2(n10306), .ZN(n13808) );
  NAND2_X1 U8712 ( .A1(n7371), .A2(n7370), .ZN(n7372) );
  NOR2_X1 U8713 ( .A1(n10601), .A2(n7381), .ZN(n7370) );
  NAND2_X1 U8714 ( .A1(n7384), .A2(n13701), .ZN(n13821) );
  NAND2_X1 U8715 ( .A1(n13770), .A2(n13771), .ZN(n7384) );
  NAND2_X1 U8716 ( .A1(n13831), .A2(n13830), .ZN(n14442) );
  INV_X1 U8717 ( .A(n10585), .ZN(n13855) );
  INV_X1 U8718 ( .A(n10404), .ZN(n13860) );
  NAND2_X1 U8719 ( .A1(n7001), .A2(n14171), .ZN(n7000) );
  NAND2_X1 U8720 ( .A1(n14011), .A2(n7003), .ZN(n7002) );
  XNOR2_X1 U8721 ( .A(n7208), .B(n7207), .ZN(n14183) );
  INV_X1 U8722 ( .A(n13997), .ZN(n7207) );
  OAI22_X1 U8723 ( .A1(n14023), .A2(n7210), .B1(n7209), .B2(n7213), .ZN(n7208)
         );
  INV_X1 U8724 ( .A(n7219), .ZN(n7209) );
  NAND2_X1 U8725 ( .A1(n6940), .A2(n6938), .ZN(n14188) );
  INV_X1 U8726 ( .A(n6939), .ZN(n6938) );
  NAND2_X1 U8727 ( .A1(n6941), .A2(n14264), .ZN(n6940) );
  OAI22_X1 U8728 ( .A1(n13582), .A2(n14136), .B1(n14138), .B2(n11597), .ZN(
        n6939) );
  AND2_X1 U8729 ( .A1(n7427), .A2(n7426), .ZN(n14021) );
  NAND2_X1 U8730 ( .A1(n6836), .A2(n7428), .ZN(n14046) );
  NAND2_X1 U8731 ( .A1(n8159), .A2(n8158), .ZN(n14236) );
  NAND2_X1 U8732 ( .A1(n7203), .A2(n7199), .ZN(n14117) );
  NOR2_X1 U8733 ( .A1(n14131), .A2(n11588), .ZN(n14119) );
  INV_X1 U8734 ( .A(n7411), .ZN(n14145) );
  AOI21_X1 U8735 ( .B1(n6862), .B2(n7415), .A(n6587), .ZN(n7411) );
  NAND2_X1 U8736 ( .A1(n6862), .A2(n11577), .ZN(n14163) );
  NOR2_X1 U8737 ( .A1(n11586), .A2(n11585), .ZN(n14150) );
  NAND2_X1 U8738 ( .A1(n8081), .A2(n8080), .ZN(n14259) );
  NAND2_X1 U8739 ( .A1(n11471), .A2(n7420), .ZN(n11579) );
  NAND2_X1 U8740 ( .A1(n6957), .A2(n6956), .ZN(n6953) );
  OAI21_X1 U8741 ( .B1(n6835), .B2(n11189), .A(n7408), .ZN(n11198) );
  NAND2_X1 U8742 ( .A1(n11102), .A2(n11101), .ZN(n11197) );
  NAND2_X1 U8743 ( .A1(n6835), .A2(n11099), .ZN(n11102) );
  NAND2_X1 U8744 ( .A1(n10785), .A2(n10784), .ZN(n10946) );
  NAND2_X1 U8745 ( .A1(n10659), .A2(n10618), .ZN(n10619) );
  NAND2_X1 U8746 ( .A1(n7762), .A2(n7761), .ZN(n10388) );
  NAND2_X1 U8747 ( .A1(n14076), .A2(n10311), .ZN(n14161) );
  INV_X1 U8748 ( .A(n14167), .ZN(n14112) );
  AND2_X1 U8749 ( .A1(n14076), .A2(n10316), .ZN(n14114) );
  NAND2_X1 U8750 ( .A1(n6718), .A2(n6717), .ZN(n6716) );
  INV_X1 U8751 ( .A(n14199), .ZN(n6717) );
  INV_X1 U8752 ( .A(n14200), .ZN(n6718) );
  INV_X2 U8753 ( .A(n14625), .ZN(n14627) );
  INV_X1 U8754 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14292) );
  NAND2_X1 U8755 ( .A1(n6817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U8756 ( .A1(n8402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8403) );
  INV_X1 U8757 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15151) );
  INV_X1 U8758 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8397) );
  XNOR2_X1 U8759 ( .A(n8174), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14307) );
  NAND2_X1 U8760 ( .A1(n7690), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7689) );
  INV_X1 U8761 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n15244) );
  INV_X1 U8762 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10300) );
  INV_X1 U8763 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n15126) );
  AND2_X1 U8764 ( .A1(n7986), .A2(n8003), .ZN(n9760) );
  INV_X1 U8765 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9714) );
  INV_X1 U8766 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9309) );
  INV_X1 U8767 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9210) );
  OAI21_X1 U8768 ( .B1(n7852), .B2(n7172), .A(n7171), .ZN(n7894) );
  INV_X1 U8769 ( .A(n7874), .ZN(n7875) );
  INV_X1 U8770 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9169) );
  INV_X1 U8771 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9162) );
  OAI21_X1 U8772 ( .B1(n7796), .B2(n6951), .A(n6949), .ZN(n7848) );
  INV_X1 U8773 ( .A(n6950), .ZN(n6949) );
  INV_X1 U8774 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9153) );
  INV_X1 U8775 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9150) );
  INV_X1 U8776 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9125) );
  NAND2_X1 U8777 ( .A1(n6711), .A2(n7715), .ZN(n7716) );
  INV_X1 U8778 ( .A(n7713), .ZN(n6711) );
  INV_X1 U8779 ( .A(P1_RD_REG_SCAN_IN), .ZN(n15076) );
  NOR2_X1 U8780 ( .A1(n7618), .A2(n15341), .ZN(n14314) );
  NOR2_X1 U8781 ( .A1(n6790), .A2(n15041), .ZN(n7611) );
  NAND2_X1 U8782 ( .A1(n7556), .A2(n6788), .ZN(n7612) );
  OR2_X1 U8783 ( .A1(n7621), .A2(n7620), .ZN(n15339) );
  XNOR2_X1 U8784 ( .A(n7624), .B(n6976), .ZN(n15328) );
  NAND2_X1 U8785 ( .A1(n15328), .A2(n15327), .ZN(n15326) );
  NAND2_X1 U8786 ( .A1(n14320), .A2(n7640), .ZN(n14324) );
  NAND2_X1 U8787 ( .A1(n6775), .A2(n6773), .ZN(n14517) );
  NAND2_X1 U8788 ( .A1(n7642), .A2(n7643), .ZN(n14522) );
  NAND2_X1 U8789 ( .A1(n14522), .A2(n14745), .ZN(n14520) );
  NOR2_X1 U8790 ( .A1(n7649), .A2(n7648), .ZN(n14529) );
  NAND2_X1 U8791 ( .A1(n7649), .A2(n7648), .ZN(n14531) );
  NAND2_X1 U8792 ( .A1(n14531), .A2(n14532), .ZN(n14528) );
  NAND2_X1 U8793 ( .A1(n14533), .A2(n6784), .ZN(n14539) );
  INV_X1 U8794 ( .A(n7650), .ZN(n6981) );
  NAND2_X1 U8795 ( .A1(n14331), .A2(n15226), .ZN(n14330) );
  INV_X1 U8796 ( .A(n6808), .ZN(n11840) );
  INV_X1 U8797 ( .A(n7049), .ZN(n10706) );
  INV_X1 U8798 ( .A(n6844), .ZN(n6843) );
  OAI22_X1 U8799 ( .A1(n12624), .A2(n12612), .B1(n15031), .B2(n12556), .ZN(
        n6844) );
  NAND2_X1 U8800 ( .A1(n7272), .A2(n14644), .ZN(n7270) );
  NAND2_X1 U8801 ( .A1(n6734), .A2(n13208), .ZN(n13442) );
  OAI21_X1 U8802 ( .B1(n13540), .B2(n13539), .A(n7537), .ZN(n13541) );
  NAND2_X1 U8803 ( .A1(n6897), .A2(n14464), .ZN(n6896) );
  NAND2_X1 U8804 ( .A1(n6713), .A2(n6712), .ZN(P1_U3555) );
  NAND2_X1 U8805 ( .A1(n14634), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U8806 ( .A1(n6716), .A2(n14636), .ZN(n6713) );
  NAND2_X1 U8807 ( .A1(n6715), .A2(n6714), .ZN(P1_U3523) );
  OR2_X1 U8808 ( .A1(n14627), .A2(n8255), .ZN(n6714) );
  NAND2_X1 U8809 ( .A1(n6716), .A2(n14627), .ZN(n6715) );
  INV_X1 U8810 ( .A(n6977), .ZN(n15329) );
  NAND2_X1 U8811 ( .A1(n14328), .A2(n14327), .ZN(n14326) );
  INV_X1 U8812 ( .A(n14525), .ZN(n14524) );
  AOI21_X1 U8813 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7653), .A(n14309), .ZN(
        n7660) );
  NAND2_X2 U8814 ( .A1(n7350), .A2(n7352), .ZN(n7858) );
  AND2_X1 U8815 ( .A1(n6948), .A2(n13849), .ZN(n6540) );
  NAND2_X1 U8816 ( .A1(n7099), .A2(n8416), .ZN(n8618) );
  AND2_X1 U8817 ( .A1(n12624), .A2(n12193), .ZN(n6541) );
  OR2_X1 U8818 ( .A1(n6574), .A2(n12265), .ZN(n6542) );
  NAND2_X2 U8819 ( .A1(n12807), .A2(n12968), .ZN(n12886) );
  AND2_X1 U8820 ( .A1(n13375), .A2(n13183), .ZN(n6543) );
  NAND2_X1 U8821 ( .A1(n7525), .A2(n7526), .ZN(n6544) );
  OR2_X1 U8822 ( .A1(n9211), .A2(n7328), .ZN(n6545) );
  XNOR2_X1 U8823 ( .A(n8568), .B(P3_IR_REG_4__SCAN_IN), .ZN(n9142) );
  OR2_X1 U8824 ( .A1(n11477), .A2(n14259), .ZN(n6546) );
  AND2_X1 U8825 ( .A1(n14070), .A2(n7015), .ZN(n6547) );
  INV_X1 U8826 ( .A(n14144), .ZN(n14133) );
  AND2_X1 U8827 ( .A1(n11587), .A2(n8119), .ZN(n14144) );
  AND2_X1 U8828 ( .A1(n7199), .A2(n6963), .ZN(n6548) );
  AND2_X1 U8829 ( .A1(n7347), .A2(n7882), .ZN(n6549) );
  OR2_X1 U8830 ( .A1(n8324), .A2(n9594), .ZN(n6550) );
  AND2_X1 U8831 ( .A1(n7015), .A2(n14042), .ZN(n6551) );
  AND2_X1 U8832 ( .A1(n6910), .A2(n6602), .ZN(n6552) );
  XNOR2_X1 U8833 ( .A(n14216), .B(n13842), .ZN(n14053) );
  INV_X1 U8834 ( .A(n14053), .ZN(n6727) );
  AND2_X1 U8835 ( .A1(n13514), .A2(n13061), .ZN(n6553) );
  INV_X1 U8836 ( .A(n11345), .ZN(n6948) );
  NAND2_X1 U8837 ( .A1(n11969), .A2(n11968), .ZN(n13460) );
  AND3_X1 U8838 ( .A1(n7825), .A2(n7794), .A3(n7847), .ZN(n6554) );
  AND2_X1 U8839 ( .A1(n7671), .A2(n7696), .ZN(n6555) );
  AND2_X1 U8840 ( .A1(n7250), .A2(n12700), .ZN(n6556) );
  AND2_X1 U8841 ( .A1(n6898), .A2(n6610), .ZN(n6557) );
  AND3_X1 U8842 ( .A1(n7065), .A2(n7064), .A3(n7066), .ZN(n6558) );
  INV_X1 U8843 ( .A(n13228), .ZN(n13542) );
  NAND2_X1 U8844 ( .A1(n11990), .A2(n11989), .ZN(n13228) );
  INV_X1 U8845 ( .A(n7218), .ZN(n7217) );
  NAND2_X1 U8846 ( .A1(n6579), .A2(n7220), .ZN(n7218) );
  AND2_X1 U8847 ( .A1(n8520), .A2(n8519), .ZN(n6559) );
  INV_X1 U8848 ( .A(n12112), .ZN(n12647) );
  NAND2_X1 U8849 ( .A1(n8835), .A2(n8834), .ZN(n12112) );
  INV_X1 U8850 ( .A(n13631), .ZN(n14450) );
  AND2_X1 U8851 ( .A1(n8065), .A2(n8064), .ZN(n13631) );
  AND2_X1 U8852 ( .A1(n8058), .A2(n9523), .ZN(n6560) );
  INV_X1 U8853 ( .A(n8336), .ZN(n7364) );
  INV_X1 U8854 ( .A(n8254), .ZN(n7342) );
  INV_X1 U8855 ( .A(n8296), .ZN(n7346) );
  AND2_X1 U8856 ( .A1(n6552), .A2(n11346), .ZN(n6561) );
  AND2_X1 U8857 ( .A1(n11806), .A2(n11712), .ZN(n6562) );
  AND2_X1 U8858 ( .A1(n7054), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n6563) );
  AND2_X1 U8859 ( .A1(n7524), .A2(n8419), .ZN(n6564) );
  INV_X1 U8860 ( .A(n8924), .ZN(n14922) );
  NAND2_X1 U8861 ( .A1(n7943), .A2(n7942), .ZN(n14504) );
  INV_X1 U8862 ( .A(n14504), .ZN(n7018) );
  AND2_X1 U8863 ( .A1(n6988), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6565) );
  INV_X1 U8864 ( .A(n8890), .ZN(n7446) );
  OR2_X1 U8865 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n11771), .ZN(n6566) );
  XOR2_X1 U8866 ( .A(n13228), .B(n12001), .Z(n6567) );
  OR2_X1 U8867 ( .A1(n8654), .A2(n8453), .ZN(n6568) );
  INV_X1 U8868 ( .A(n13019), .ZN(n7141) );
  OR2_X1 U8869 ( .A1(n13302), .A2(n13470), .ZN(n6569) );
  NAND2_X1 U8870 ( .A1(n13179), .A2(n7166), .ZN(n7165) );
  AND2_X1 U8871 ( .A1(n7825), .A2(n6722), .ZN(n6570) );
  INV_X1 U8872 ( .A(n9091), .ZN(n9813) );
  INV_X1 U8873 ( .A(n13859), .ZN(n6683) );
  AND2_X1 U8874 ( .A1(n13460), .A2(n13274), .ZN(n6572) );
  NOR2_X1 U8875 ( .A1(n8642), .A2(n8628), .ZN(n6573) );
  INV_X1 U8876 ( .A(n9970), .ZN(n11977) );
  NAND2_X1 U8877 ( .A1(n12262), .A2(n12277), .ZN(n6574) );
  NAND2_X1 U8878 ( .A1(n8025), .A2(n7367), .ZN(n7687) );
  NAND2_X1 U8879 ( .A1(n7699), .A2(n7666), .ZN(n7739) );
  OR2_X1 U8880 ( .A1(n9015), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n6575) );
  NAND4_X1 U8881 ( .A1(n7523), .A2(n7098), .A3(n7524), .A4(n7099), .ZN(n6576)
         );
  AND4_X1 U8882 ( .A1(n9010), .A2(n9164), .A3(n9285), .A4(n9009), .ZN(n6577)
         );
  AND2_X1 U8883 ( .A1(n10193), .A2(n10337), .ZN(n6578) );
  INV_X1 U8884 ( .A(n13172), .ZN(n13223) );
  OR2_X1 U8885 ( .A1(n14031), .A2(n14004), .ZN(n6579) );
  NOR2_X1 U8886 ( .A1(n12511), .A2(n12525), .ZN(n6580) );
  AND2_X1 U8887 ( .A1(n14254), .A2(n14456), .ZN(n6581) );
  OR2_X1 U8888 ( .A1(n14436), .A2(n13833), .ZN(n11414) );
  INV_X1 U8889 ( .A(n6937), .ZN(n6936) );
  OAI21_X1 U8890 ( .B1(n7257), .B2(n10732), .A(n7256), .ZN(n6937) );
  NOR2_X1 U8891 ( .A1(n12413), .A2(n12418), .ZN(n6582) );
  AND4_X1 U8892 ( .A1(n9018), .A2(n9029), .A3(n9017), .A4(n9016), .ZN(n6583)
         );
  INV_X1 U8893 ( .A(n6962), .ZN(n14132) );
  AOI21_X1 U8894 ( .B1(n11586), .B2(n14149), .A(n6964), .ZN(n6962) );
  AND2_X1 U8895 ( .A1(n7734), .A2(n7736), .ZN(n6584) );
  AND2_X1 U8896 ( .A1(n11414), .A2(n11310), .ZN(n6585) );
  OR2_X1 U8897 ( .A1(n12642), .A2(n12444), .ZN(n6586) );
  NOR2_X1 U8898 ( .A1(n6581), .A2(n11580), .ZN(n6587) );
  AND2_X1 U8899 ( .A1(n11415), .A2(n7358), .ZN(n6588) );
  AND2_X1 U8900 ( .A1(n7788), .A2(n7787), .ZN(n10453) );
  NAND2_X1 U8901 ( .A1(n11660), .A2(n11658), .ZN(n6864) );
  INV_X1 U8902 ( .A(n10337), .ZN(n7381) );
  AND2_X1 U8903 ( .A1(n12398), .A2(n7498), .ZN(n6589) );
  INV_X1 U8904 ( .A(n13737), .ZN(n6905) );
  OR2_X1 U8905 ( .A1(n8099), .A2(n11578), .ZN(n6590) );
  NAND2_X1 U8906 ( .A1(n7247), .A2(n11929), .ZN(n12752) );
  INV_X1 U8907 ( .A(n8160), .ZN(n6872) );
  NAND2_X1 U8908 ( .A1(n12293), .A2(n12323), .ZN(n6591) );
  OR2_X1 U8909 ( .A1(n12639), .A2(n12162), .ZN(n6592) );
  INV_X1 U8910 ( .A(n11520), .ZN(n7264) );
  INV_X1 U8911 ( .A(n13027), .ZN(n11557) );
  XNOR2_X1 U8912 ( .A(n12897), .B(n13406), .ZN(n13027) );
  AND2_X1 U8913 ( .A1(n13605), .A2(n13607), .ZN(n6593) );
  INV_X1 U8914 ( .A(n12932), .ZN(n7337) );
  AND2_X1 U8915 ( .A1(n12551), .A2(n15011), .ZN(n6594) );
  INV_X1 U8916 ( .A(n8335), .ZN(n7365) );
  INV_X1 U8917 ( .A(n13982), .ZN(n14189) );
  NAND2_X1 U8918 ( .A1(n8294), .A2(n8293), .ZN(n13982) );
  AND2_X1 U8919 ( .A1(n7527), .A2(n8431), .ZN(n6595) );
  AND2_X1 U8920 ( .A1(n7652), .A2(n6779), .ZN(n6596) );
  AND2_X1 U8921 ( .A1(n8103), .A2(n8102), .ZN(n6597) );
  OR2_X1 U8922 ( .A1(n7608), .A2(n7609), .ZN(n6598) );
  AND2_X1 U8923 ( .A1(n13454), .A2(n13252), .ZN(n6599) );
  INV_X1 U8924 ( .A(n13439), .ZN(n13212) );
  NAND2_X1 U8925 ( .A1(n7176), .A2(n6670), .ZN(n13439) );
  AND2_X1 U8926 ( .A1(n13830), .A2(n13639), .ZN(n6600) );
  OR2_X1 U8927 ( .A1(n9078), .A2(n9677), .ZN(n6601) );
  NAND2_X1 U8928 ( .A1(n11339), .A2(n11338), .ZN(n6602) );
  NAND2_X1 U8929 ( .A1(n11045), .A2(n8672), .ZN(n6603) );
  NAND2_X1 U8930 ( .A1(n12955), .A2(n12954), .ZN(n6604) );
  AND2_X1 U8931 ( .A1(n13668), .A2(n13666), .ZN(n6605) );
  OR2_X1 U8932 ( .A1(n6995), .A2(n11076), .ZN(n6606) );
  AND2_X1 U8933 ( .A1(n6864), .A2(n8592), .ZN(n6607) );
  INV_X1 U8934 ( .A(n13140), .ZN(n13537) );
  NAND2_X1 U8935 ( .A1(n12967), .A2(n12966), .ZN(n13140) );
  INV_X1 U8936 ( .A(n13978), .ZN(n14175) );
  NAND2_X1 U8937 ( .A1(n8329), .A2(n8328), .ZN(n13978) );
  INV_X1 U8938 ( .A(n7267), .ZN(n7263) );
  NAND2_X1 U8939 ( .A1(n10739), .A2(n10740), .ZN(n7267) );
  INV_X1 U8940 ( .A(n11613), .ZN(n7499) );
  OR2_X1 U8941 ( .A1(n12047), .A2(n12386), .ZN(n11613) );
  AND2_X1 U8942 ( .A1(n13685), .A2(n13684), .ZN(n6608) );
  AND2_X1 U8943 ( .A1(n6774), .A2(n6773), .ZN(n6609) );
  NAND2_X1 U8944 ( .A1(n6903), .A2(n6901), .ZN(n6610) );
  INV_X1 U8945 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7696) );
  AND2_X1 U8946 ( .A1(n13982), .A2(n13994), .ZN(n6611) );
  INV_X1 U8947 ( .A(n7837), .ZN(n6758) );
  NAND2_X1 U8948 ( .A1(n8252), .A2(n8251), .ZN(n14201) );
  INV_X1 U8949 ( .A(n14201), .ZN(n14031) );
  INV_X1 U8950 ( .A(n14209), .ZN(n14042) );
  NAND2_X1 U8951 ( .A1(n8233), .A2(n8232), .ZN(n14209) );
  AND2_X1 U8952 ( .A1(n7980), .A2(n15171), .ZN(n6612) );
  NAND2_X1 U8953 ( .A1(n14143), .A2(n13816), .ZN(n6613) );
  NOR2_X1 U8954 ( .A1(n13493), .A2(n13160), .ZN(n6614) );
  AND2_X1 U8955 ( .A1(n6973), .A2(n6971), .ZN(n6615) );
  AND2_X1 U8956 ( .A1(n6567), .A2(n7276), .ZN(n6616) );
  XNOR2_X1 U8957 ( .A(n7689), .B(n6707), .ZN(n11073) );
  INV_X1 U8958 ( .A(n11073), .ZN(n7353) );
  INV_X1 U8959 ( .A(n11593), .ZN(n7224) );
  AND2_X1 U8960 ( .A1(n14074), .A2(n11592), .ZN(n11593) );
  AND2_X1 U8961 ( .A1(n10045), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6617) );
  AND2_X1 U8962 ( .A1(n14786), .A2(n10649), .ZN(n6618) );
  NOR2_X1 U8963 ( .A1(n14216), .A2(n13773), .ZN(n6619) );
  AND2_X1 U8964 ( .A1(n7348), .A2(n7883), .ZN(n6620) );
  OR2_X1 U8965 ( .A1(n7905), .A2(n7903), .ZN(n6621) );
  AND2_X1 U8966 ( .A1(n13299), .A2(n13166), .ZN(n6622) );
  INV_X1 U8967 ( .A(n7825), .ZN(n6951) );
  NAND2_X1 U8968 ( .A1(n6723), .A2(SI_5_), .ZN(n7825) );
  INV_X1 U8969 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8419) );
  INV_X1 U8970 ( .A(n7167), .ZN(n7166) );
  OR2_X1 U8971 ( .A1(n13182), .A2(n7168), .ZN(n7167) );
  INV_X1 U8972 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7671) );
  INV_X1 U8973 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8427) );
  INV_X1 U8974 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9156) );
  INV_X1 U8975 ( .A(n7108), .ZN(n7107) );
  NAND2_X1 U8976 ( .A1(n7112), .A2(n7113), .ZN(n7108) );
  AND2_X1 U8977 ( .A1(n13621), .A2(n13620), .ZN(n6623) );
  OR2_X1 U8978 ( .A1(n7558), .A2(n7557), .ZN(n6624) );
  AND2_X1 U8979 ( .A1(n13710), .A2(n13709), .ZN(n6625) );
  OR2_X1 U8980 ( .A1(n7189), .A2(n8055), .ZN(n6626) );
  NAND2_X1 U8981 ( .A1(n11894), .A2(n12723), .ZN(n6627) );
  AND2_X1 U8982 ( .A1(n9210), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6628) );
  AND2_X1 U8983 ( .A1(n9209), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n6629) );
  AND2_X1 U8984 ( .A1(n11130), .A2(n12076), .ZN(n6630) );
  AND2_X1 U8985 ( .A1(n7265), .A2(n7267), .ZN(n6631) );
  INV_X1 U8986 ( .A(n6864), .ZN(n11791) );
  NAND2_X1 U8987 ( .A1(n7216), .A2(n7220), .ZN(n7215) );
  INV_X1 U8988 ( .A(n7215), .ZN(n7214) );
  INV_X1 U8989 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8487) );
  INV_X1 U8990 ( .A(n8215), .ZN(n7357) );
  INV_X1 U8991 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15104) );
  INV_X1 U8992 ( .A(n12883), .ZN(n7323) );
  INV_X1 U8993 ( .A(n11456), .ZN(n11458) );
  AND2_X1 U8994 ( .A1(n7223), .A2(n6970), .ZN(n6632) );
  MUX2_X1 U8995 ( .A(n13073), .B(n12820), .S(n12833), .Z(n12822) );
  AND3_X1 U8996 ( .A1(n7543), .A2(n7288), .A3(n9336), .ZN(n6633) );
  AND3_X1 U8997 ( .A1(n13038), .A2(n9334), .A3(n13051), .ZN(n6634) );
  OR2_X1 U8998 ( .A1(n10147), .A2(n10131), .ZN(n6635) );
  AND2_X1 U8999 ( .A1(n7424), .A2(n14022), .ZN(n6636) );
  AND2_X1 U9000 ( .A1(n12635), .A2(n12066), .ZN(n6637) );
  INV_X1 U9001 ( .A(n8521), .ZN(n14941) );
  NAND2_X1 U9002 ( .A1(n6559), .A2(n6601), .ZN(n8521) );
  AND2_X1 U9003 ( .A1(n6568), .A2(n8454), .ZN(n6638) );
  AND2_X1 U9004 ( .A1(n13192), .A2(n13284), .ZN(n6639) );
  AND2_X1 U9005 ( .A1(n11414), .A2(n8038), .ZN(n11415) );
  INV_X1 U9006 ( .A(n11415), .ZN(n6959) );
  AND2_X1 U9007 ( .A1(n12893), .A2(n7303), .ZN(n6640) );
  AND2_X1 U9008 ( .A1(n12999), .A2(n12998), .ZN(n6641) );
  INV_X1 U9009 ( .A(n7180), .ZN(n7179) );
  OAI21_X1 U9010 ( .B1(n7182), .B2(n7181), .A(n7977), .ZN(n7180) );
  AND2_X1 U9011 ( .A1(n11531), .A2(n7285), .ZN(n6642) );
  AND2_X1 U9012 ( .A1(n13657), .A2(n13655), .ZN(n6643) );
  OR2_X1 U9013 ( .A1(n12868), .A2(n12866), .ZN(n6644) );
  OR2_X1 U9014 ( .A1(n7310), .A2(n12915), .ZN(n6645) );
  OR2_X1 U9015 ( .A1(n6872), .A2(n8161), .ZN(n6646) );
  AND2_X1 U9016 ( .A1(n7059), .A2(n9091), .ZN(n6647) );
  NOR2_X1 U9017 ( .A1(n13049), .A2(n13412), .ZN(n6648) );
  AND2_X1 U9018 ( .A1(n7067), .A2(n6574), .ZN(n6649) );
  NOR2_X1 U9019 ( .A1(n12428), .A2(n12430), .ZN(n6863) );
  OR2_X1 U9020 ( .A1(n7946), .A2(n7944), .ZN(n6650) );
  AND2_X1 U9021 ( .A1(n7225), .A2(n7224), .ZN(n6651) );
  AND2_X1 U9022 ( .A1(n11753), .A2(n12371), .ZN(n12382) );
  INV_X1 U9023 ( .A(n12382), .ZN(n12383) );
  INV_X1 U9024 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7332) );
  NAND2_X1 U9025 ( .A1(n11984), .A2(n6567), .ZN(n6652) );
  INV_X1 U9026 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7688) );
  AND2_X1 U9027 ( .A1(n7489), .A2(n7486), .ZN(n7485) );
  NAND2_X1 U9028 ( .A1(n6967), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6653) );
  INV_X1 U9029 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9336) );
  INV_X1 U9030 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9212) );
  AND2_X1 U9031 ( .A1(n14342), .A2(n12537), .ZN(n6654) );
  INV_X1 U9032 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U9033 ( .A1(n11311), .A2(n6585), .ZN(n6957) );
  NAND2_X1 U9034 ( .A1(n6737), .A2(n11382), .ZN(n11543) );
  INV_X1 U9035 ( .A(n13238), .ZN(n13274) );
  INV_X1 U9036 ( .A(n14866), .ZN(n6995) );
  NAND2_X1 U9037 ( .A1(n6953), .A2(n11455), .ZN(n11474) );
  NAND2_X1 U9038 ( .A1(n11917), .A2(n11916), .ZN(n13476) );
  INV_X1 U9039 ( .A(n13476), .ZN(n7229) );
  AND2_X1 U9040 ( .A1(n12061), .A2(n12456), .ZN(n6655) );
  OR2_X1 U9041 ( .A1(n8049), .A2(n8048), .ZN(n14458) );
  NOR2_X1 U9042 ( .A1(n7642), .A2(n7643), .ZN(n14521) );
  INV_X1 U9043 ( .A(n14521), .ZN(n6787) );
  INV_X1 U9044 ( .A(n8466), .ZN(n7466) );
  NAND2_X1 U9045 ( .A1(n14118), .A2(n11587), .ZN(n7202) );
  INV_X1 U9046 ( .A(n7202), .ZN(n7199) );
  AND2_X1 U9047 ( .A1(n12524), .A2(n8790), .ZN(n6656) );
  INV_X1 U9048 ( .A(n6847), .ZN(n11442) );
  NOR2_X1 U9049 ( .A1(n11443), .A2(n13521), .ZN(n6847) );
  INV_X1 U9050 ( .A(n7238), .ZN(n13385) );
  AND2_X1 U9051 ( .A1(n12039), .A2(n12162), .ZN(n6657) );
  INV_X1 U9052 ( .A(n7010), .ZN(n14155) );
  NOR3_X1 U9053 ( .A1(n11477), .A2(n14259), .A3(n14254), .ZN(n7010) );
  AND2_X1 U9054 ( .A1(n7278), .A2(n12740), .ZN(n6658) );
  INV_X1 U9055 ( .A(n7009), .ZN(n14140) );
  NOR2_X1 U9056 ( .A1(n11477), .A2(n7011), .ZN(n7009) );
  OR2_X1 U9057 ( .A1(n13631), .A2(n14458), .ZN(n6659) );
  NOR2_X1 U9058 ( .A1(n11200), .A2(n13610), .ZN(n11305) );
  AND2_X1 U9059 ( .A1(n6935), .A2(n6936), .ZN(n6660) );
  NOR2_X1 U9060 ( .A1(n8739), .A2(n7464), .ZN(n7463) );
  NAND2_X2 U9061 ( .A1(n13989), .A2(n14106), .ZN(n14076) );
  INV_X1 U9062 ( .A(n14652), .ZN(n14644) );
  INV_X2 U9063 ( .A(n12886), .ZN(n12973) );
  NAND2_X1 U9064 ( .A1(n11864), .A2(n11863), .ZN(n13375) );
  INV_X1 U9065 ( .A(n13375), .ZN(n7237) );
  NAND2_X1 U9066 ( .A1(n11385), .A2(n11384), .ZN(n12897) );
  INV_X1 U9067 ( .A(n12897), .ZN(n6846) );
  INV_X1 U9068 ( .A(n13601), .ZN(n7016) );
  NAND2_X1 U9069 ( .A1(n8980), .A2(n11829), .ZN(n14934) );
  INV_X1 U9070 ( .A(n14934), .ZN(n14949) );
  AND2_X1 U9071 ( .A1(n12234), .A2(n14882), .ZN(n6661) );
  XOR2_X1 U9072 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .Z(n6662) );
  AND2_X1 U9073 ( .A1(n10891), .A2(n10890), .ZN(n6663) );
  NAND2_X1 U9074 ( .A1(n9603), .A2(n9589), .ZN(n14476) );
  NAND2_X1 U9075 ( .A1(n10790), .A2(n6948), .ZN(n10955) );
  INV_X1 U9076 ( .A(n10955), .ZN(n7019) );
  NOR2_X1 U9077 ( .A1(n6864), .A2(n7546), .ZN(n6664) );
  INV_X1 U9078 ( .A(n7508), .ZN(n7507) );
  NOR2_X1 U9079 ( .A1(n11430), .A2(n7509), .ZN(n7508) );
  AND2_X1 U9080 ( .A1(n10240), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n6665) );
  AND2_X1 U9081 ( .A1(n11869), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6666) );
  AND2_X1 U9082 ( .A1(n8249), .A2(n7195), .ZN(n6667) );
  OR2_X1 U9083 ( .A1(n12265), .A2(n12610), .ZN(n6668) );
  INV_X1 U9084 ( .A(n8931), .ZN(n7480) );
  INV_X1 U9085 ( .A(n11789), .ZN(n7478) );
  INV_X1 U9086 ( .A(n13833), .ZN(n6793) );
  INV_X2 U9087 ( .A(n14634), .ZN(n14636) );
  OR2_X1 U9088 ( .A1(n9590), .A2(n10792), .ZN(n6669) );
  INV_X1 U9089 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n15117) );
  INV_X1 U9090 ( .A(n11666), .ZN(n6819) );
  INV_X1 U9091 ( .A(n14844), .ZN(n7241) );
  INV_X1 U9092 ( .A(n14639), .ZN(n7239) );
  INV_X1 U9093 ( .A(n7448), .ZN(n7447) );
  NAND2_X1 U9094 ( .A1(n6672), .A2(n8892), .ZN(n7448) );
  AND2_X1 U9095 ( .A1(n9514), .A2(n9513), .ZN(n14275) );
  INV_X1 U9096 ( .A(n14275), .ZN(n14264) );
  OR2_X1 U9097 ( .A1(n6521), .A2(n13570), .ZN(n6670) );
  AND2_X1 U9098 ( .A1(n7448), .A2(n6566), .ZN(n6671) );
  INV_X1 U9099 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6816) );
  OR2_X1 U9100 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13570), .ZN(n6672) );
  AND2_X1 U9101 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13570), .ZN(n6673) );
  INV_X1 U9102 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13579) );
  AND2_X1 U9103 ( .A1(n7445), .A2(n6566), .ZN(n6674) );
  AND2_X1 U9104 ( .A1(n12256), .A2(n12268), .ZN(n6675) );
  AND2_X1 U9105 ( .A1(n6766), .A2(n8575), .ZN(n6676) );
  INV_X1 U9106 ( .A(n12265), .ZN(n7066) );
  OR2_X1 U9107 ( .A1(n12236), .A2(n14882), .ZN(n6680) );
  INV_X1 U9108 ( .A(n14882), .ZN(n6828) );
  OR2_X1 U9109 ( .A1(n12235), .A2(n14882), .ZN(n6987) );
  OR2_X1 U9110 ( .A1(n12234), .A2(n14882), .ZN(n6988) );
  OR2_X2 U9111 ( .A1(n12284), .A2(n12283), .ZN(n12292) );
  OR2_X2 U9112 ( .A1(n10712), .A2(n10711), .ZN(n11082) );
  NOR2_X2 U9113 ( .A1(n12238), .A2(n12237), .ZN(n12254) );
  AND2_X2 U9114 ( .A1(n6989), .A2(n6680), .ZN(n12238) );
  NAND2_X1 U9115 ( .A1(n10605), .A2(n13859), .ZN(n6682) );
  OAI22_X1 U9116 ( .A1(n13740), .A2(n6683), .B1(n7725), .B2(n13741), .ZN(n9691) );
  OAI22_X1 U9117 ( .A1(n14136), .A2(n6683), .B1(n10365), .B2(n14138), .ZN(
        n10366) );
  OAI22_X1 U9118 ( .A1(n14470), .A2(n6683), .B1(n14471), .B2(n10365), .ZN(
        n9707) );
  NAND3_X1 U9119 ( .A1(n7836), .A2(n7838), .A3(n6758), .ZN(n6686) );
  NAND2_X1 U9120 ( .A1(n6692), .A2(n6597), .ZN(n6691) );
  AOI21_X1 U9121 ( .B1(n8193), .B2(n8194), .A(n6826), .ZN(n6870) );
  NAND2_X1 U9122 ( .A1(n6752), .A2(n6693), .ZN(n8193) );
  NAND3_X1 U9123 ( .A1(n6700), .A2(n6650), .A3(n6698), .ZN(n6821) );
  NAND2_X1 U9124 ( .A1(n6699), .A2(n7928), .ZN(n6698) );
  INV_X1 U9125 ( .A(n6702), .ZN(n6699) );
  NAND2_X1 U9126 ( .A1(n6701), .A2(n7926), .ZN(n6700) );
  NAND2_X1 U9127 ( .A1(n6702), .A2(n7927), .ZN(n6701) );
  NAND2_X1 U9128 ( .A1(n6748), .A2(n6874), .ZN(n6702) );
  NOR2_X2 U9129 ( .A1(n8399), .A2(n6703), .ZN(n7670) );
  NAND3_X1 U9130 ( .A1(n6705), .A2(n6706), .A3(n7669), .ZN(n6703) );
  NAND4_X1 U9131 ( .A1(n6704), .A2(n8390), .A3(n6707), .A4(n7688), .ZN(n8399)
         );
  NAND2_X1 U9132 ( .A1(n7814), .A2(n7815), .ZN(n7813) );
  NAND2_X1 U9133 ( .A1(n6710), .A2(n7790), .ZN(n6708) );
  OAI21_X1 U9134 ( .B1(n6710), .B2(n7790), .A(n7789), .ZN(n6709) );
  AND2_X1 U9135 ( .A1(n6833), .A2(n7741), .ZN(n7713) );
  NAND2_X1 U9136 ( .A1(n6967), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U9137 ( .A1(n7919), .A2(n7918), .ZN(n7937) );
  OAI21_X1 U9138 ( .B1(n7919), .B2(n7180), .A(n6725), .ZN(n7994) );
  NAND2_X1 U9139 ( .A1(n6731), .A2(n6730), .ZN(n10772) );
  XNOR2_X1 U9140 ( .A(n13203), .B(n13202), .ZN(n6735) );
  NAND2_X1 U9141 ( .A1(n11543), .A2(n7142), .ZN(n6736) );
  NAND2_X1 U9142 ( .A1(n11440), .A2(n11380), .ZN(n6737) );
  OAI21_X1 U9143 ( .B1(n13010), .B2(n6738), .A(n10209), .ZN(n9913) );
  NAND2_X1 U9144 ( .A1(n9911), .A2(n9910), .ZN(n6738) );
  NAND2_X2 U9145 ( .A1(n13577), .A2(n9223), .ZN(n9346) );
  OAI21_X2 U9146 ( .B1(n9211), .B2(n7330), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6739) );
  XNOR2_X2 U9147 ( .A(n6740), .B(n9213), .ZN(n13577) );
  OR2_X2 U9148 ( .A1(n10998), .A2(n10997), .ZN(n11135) );
  AOI21_X1 U9149 ( .B1(n6524), .B2(n9640), .A(n6743), .ZN(n6742) );
  NOR2_X1 U9150 ( .A1(n10495), .A2(n9643), .ZN(n6743) );
  NOR2_X2 U9151 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n7938) );
  NAND3_X1 U9152 ( .A1(n6746), .A2(n7884), .A3(n6744), .ZN(n6748) );
  OAI21_X1 U9153 ( .B1(n8235), .B2(n8236), .A(n7339), .ZN(n6749) );
  NAND3_X1 U9154 ( .A1(n8041), .A2(n6755), .A3(n6754), .ZN(n8043) );
  NAND3_X1 U9155 ( .A1(n7970), .A2(n6588), .A3(n7969), .ZN(n6755) );
  NAND2_X1 U9156 ( .A1(n6765), .A2(n10422), .ZN(n6766) );
  OR2_X2 U9157 ( .A1(n12381), .A2(n12382), .ZN(n7039) );
  AND2_X2 U9158 ( .A1(n12524), .A2(n6768), .ZN(n12507) );
  NAND2_X1 U9159 ( .A1(n12493), .A2(n12503), .ZN(n12492) );
  NAND3_X1 U9160 ( .A1(n6772), .A2(n7556), .A3(n6788), .ZN(n6771) );
  INV_X1 U9161 ( .A(n15041), .ZN(n6772) );
  NAND2_X1 U9162 ( .A1(n14533), .A2(n6783), .ZN(n6782) );
  NAND2_X1 U9163 ( .A1(n14528), .A2(n14530), .ZN(n14535) );
  NAND3_X1 U9164 ( .A1(n14528), .A2(n14530), .A3(n6786), .ZN(n6780) );
  NOR2_X1 U9165 ( .A1(n15333), .A2(n7635), .ZN(n7638) );
  XNOR2_X1 U9166 ( .A(n7638), .B(n6984), .ZN(n14321) );
  NOR2_X1 U9167 ( .A1(n15335), .A2(n15334), .ZN(n15333) );
  XNOR2_X1 U9168 ( .A(n7651), .B(n6981), .ZN(n14331) );
  NOR2_X1 U9169 ( .A1(n14319), .A2(n14318), .ZN(n14317) );
  NOR2_X1 U9170 ( .A1(n14323), .A2(n14324), .ZN(n7641) );
  INV_X1 U9171 ( .A(n7614), .ZN(n6839) );
  OAI21_X2 U9172 ( .B1(n14370), .B2(n6630), .A(n8692), .ZN(n11317) );
  AOI21_X2 U9173 ( .B1(n8920), .B2(n14934), .A(n8919), .ZN(n11576) );
  NAND2_X1 U9174 ( .A1(n12412), .A2(n7552), .ZN(n12401) );
  NAND2_X1 U9175 ( .A1(n12492), .A2(n8819), .ZN(n12479) );
  NAND2_X1 U9176 ( .A1(n12414), .A2(n12413), .ZN(n12412) );
  NAND2_X1 U9177 ( .A1(n6791), .A2(n6856), .ZN(n6855) );
  NAND2_X1 U9178 ( .A1(n10015), .A2(n10377), .ZN(n10017) );
  NAND2_X1 U9179 ( .A1(n10573), .A2(n10449), .ZN(n10451) );
  NAND2_X1 U9180 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  NAND3_X1 U9181 ( .A1(n6584), .A2(n7735), .A3(n7733), .ZN(n13858) );
  NAND2_X1 U9182 ( .A1(n10358), .A2(n10012), .ZN(n10014) );
  NAND2_X1 U9183 ( .A1(n10021), .A2(n7763), .ZN(n10012) );
  OAI21_X1 U9184 ( .B1(n10446), .B2(n10445), .A(n10444), .ZN(n10571) );
  NAND2_X1 U9185 ( .A1(n10910), .A2(n8610), .ZN(n10872) );
  NAND2_X1 U9186 ( .A1(n8529), .A2(n8528), .ZN(n8921) );
  XNOR2_X2 U9187 ( .A(n8428), .B(n12675), .ZN(n12686) );
  AND2_X1 U9188 ( .A1(n8510), .A2(n8511), .ZN(n7540) );
  AND2_X1 U9189 ( .A1(n8544), .A2(n8543), .ZN(n6794) );
  NAND2_X1 U9190 ( .A1(n8676), .A2(n8675), .ZN(n14370) );
  NAND2_X4 U9191 ( .A1(n8433), .A2(n8434), .ZN(n11767) );
  NAND2_X1 U9192 ( .A1(n8522), .A2(n8521), .ZN(n8923) );
  NAND2_X1 U9193 ( .A1(n10872), .A2(n10871), .ZN(n10870) );
  NAND2_X1 U9194 ( .A1(n7898), .A2(n7897), .ZN(n7915) );
  INV_X1 U9195 ( .A(n8291), .ZN(n6801) );
  OAI21_X1 U9196 ( .B1(n6536), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n6861), .ZN(
        n7712) );
  NAND2_X1 U9197 ( .A1(n7746), .A2(n7747), .ZN(n7757) );
  NAND2_X1 U9198 ( .A1(n7742), .A2(n7741), .ZN(n7746) );
  NOR3_X1 U9199 ( .A1(n8387), .A2(n8386), .A3(n8385), .ZN(n8394) );
  AOI21_X1 U9200 ( .B1(n8083), .B2(n8082), .A(n6804), .ZN(n6803) );
  OAI21_X1 U9201 ( .B1(n8266), .B2(n8267), .A(n7343), .ZN(n6867) );
  NOR2_X1 U9202 ( .A1(n14080), .A2(n11581), .ZN(n14051) );
  OAI22_X1 U9203 ( .A1(n8002), .A2(n9344), .B1(n7759), .B2(n13867), .ZN(n6998)
         );
  AND2_X1 U9204 ( .A1(n7938), .A2(n7663), .ZN(n6999) );
  NAND2_X1 U9205 ( .A1(n14051), .A2(n6727), .ZN(n14050) );
  CLKBUF_X2 U9206 ( .A(n7724), .Z(n13859) );
  AOI21_X2 U9207 ( .B1(n6807), .B2(n6806), .A(n6805), .ZN(n8507) );
  NAND2_X1 U9208 ( .A1(n8855), .A2(n8853), .ZN(n8482) );
  NAND2_X1 U9209 ( .A1(n8754), .A2(n8753), .ZN(n8752) );
  AOI21_X2 U9210 ( .B1(n7469), .B2(n7468), .A(n6666), .ZN(n8833) );
  INV_X1 U9211 ( .A(n7498), .ZN(n7496) );
  OAI21_X1 U9212 ( .B1(n6568), .B2(n7458), .A(n7456), .ZN(n8459) );
  NAND2_X1 U9213 ( .A1(n7500), .A2(n11751), .ZN(n11824) );
  NAND2_X1 U9214 ( .A1(n6849), .A2(n6848), .ZN(n12921) );
  NAND3_X1 U9215 ( .A1(n7297), .A2(n7295), .A3(n7296), .ZN(n12817) );
  NAND2_X1 U9216 ( .A1(n7292), .A2(n7289), .ZN(n12904) );
  NAND2_X1 U9217 ( .A1(n12856), .A2(n12855), .ZN(n12860) );
  OAI21_X1 U9218 ( .B1(n12912), .B2(n12911), .A(n12910), .ZN(n12914) );
  AND2_X2 U9219 ( .A1(n9331), .A2(n7131), .ZN(n9019) );
  NAND2_X1 U9220 ( .A1(n9718), .A2(n9719), .ZN(n9717) );
  OR2_X2 U9221 ( .A1(n12233), .A2(n12232), .ZN(n12235) );
  NAND2_X1 U9222 ( .A1(n7713), .A2(n7714), .ZN(n7742) );
  NAND2_X1 U9223 ( .A1(n7349), .A2(n7348), .ZN(n7347) );
  NAND2_X1 U9224 ( .A1(n11637), .A2(n11636), .ZN(n8924) );
  NAND2_X1 U9225 ( .A1(n13193), .A2(n6639), .ZN(n13283) );
  NAND2_X1 U9226 ( .A1(n13194), .A2(n13266), .ZN(n13271) );
  NAND2_X1 U9227 ( .A1(n7152), .A2(n7154), .ZN(n11440) );
  NAND2_X2 U9228 ( .A1(n6997), .A2(n7717), .ZN(n10415) );
  NAND3_X1 U9229 ( .A1(n12818), .A2(n12819), .A3(n7312), .ZN(n7311) );
  NAND2_X1 U9230 ( .A1(n12817), .A2(n12816), .ZN(n12815) );
  INV_X1 U9231 ( .A(n7724), .ZN(n6814) );
  INV_X1 U9232 ( .A(n6998), .ZN(n6997) );
  NOR2_X2 U9233 ( .A1(n6571), .A2(n13412), .ZN(n12807) );
  NAND2_X1 U9234 ( .A1(n12896), .A2(n12895), .ZN(n7294) );
  NAND2_X1 U9235 ( .A1(n13047), .A2(n13039), .ZN(n6834) );
  NAND2_X1 U9236 ( .A1(n6834), .A2(n6634), .ZN(n13057) );
  OR2_X2 U9237 ( .A1(n10733), .A2(n6932), .ZN(n6931) );
  AOI21_X2 U9238 ( .B1(n9740), .B2(n9739), .A(n6815), .ZN(n9748) );
  NAND2_X2 U9239 ( .A1(n12780), .A2(n12779), .ZN(n12778) );
  NAND2_X1 U9240 ( .A1(n9854), .A2(n9855), .ZN(n9966) );
  NAND2_X1 U9241 ( .A1(n6642), .A2(n12795), .ZN(n7284) );
  NOR2_X1 U9242 ( .A1(n7607), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n7560) );
  XNOR2_X1 U9243 ( .A(n7633), .B(n7634), .ZN(n15334) );
  NAND2_X1 U9244 ( .A1(n9354), .A2(n6919), .ZN(n6921) );
  NAND2_X1 U9245 ( .A1(n7613), .A2(n7614), .ZN(n7556) );
  NAND2_X1 U9246 ( .A1(n7764), .A2(n7765), .ZN(n7766) );
  INV_X4 U9247 ( .A(n7858), .ZN(n8376) );
  OAI21_X1 U9248 ( .B1(n8193), .B2(n8194), .A(n7354), .ZN(n6869) );
  NAND3_X1 U9249 ( .A1(n8022), .A2(n6555), .A3(n7670), .ZN(n6817) );
  NAND3_X1 U9250 ( .A1(n6818), .A2(n7554), .A3(n7684), .ZN(n7724) );
  NAND2_X1 U9251 ( .A1(n7971), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6818) );
  NAND2_X1 U9252 ( .A1(n7039), .A2(n7037), .ZN(n12367) );
  NAND2_X1 U9253 ( .A1(n7915), .A2(n7914), .ZN(n7919) );
  NAND2_X1 U9254 ( .A1(n7999), .A2(n8019), .ZN(n8000) );
  INV_X1 U9255 ( .A(n8056), .ZN(n6832) );
  NAND2_X1 U9256 ( .A1(n6821), .A2(n6820), .ZN(n7965) );
  NAND2_X1 U9257 ( .A1(n7726), .A2(n10020), .ZN(n7727) );
  NAND2_X2 U9258 ( .A1(n11461), .A2(n11473), .ZN(n11471) );
  NAND2_X1 U9259 ( .A1(n10406), .A2(n10009), .ZN(n10011) );
  NAND2_X1 U9260 ( .A1(n7423), .A2(n7421), .ZN(n14002) );
  AOI21_X1 U9261 ( .B1(n14992), .B2(n12555), .A(n12554), .ZN(n12621) );
  NAND2_X1 U9262 ( .A1(n12479), .A2(n12483), .ZN(n12478) );
  OR2_X1 U9263 ( .A1(n10404), .A2(n10312), .ZN(n10406) );
  NOR2_X1 U9264 ( .A1(n14002), .A2(n14005), .ZN(n14001) );
  AND4_X2 U9265 ( .A1(n6550), .A2(n7721), .A3(n7720), .A4(n7719), .ZN(n10404)
         );
  NAND2_X1 U9266 ( .A1(n12125), .A2(n12022), .ZN(n12168) );
  NAND2_X1 U9267 ( .A1(n10451), .A2(n10450), .ZN(n10553) );
  NAND2_X1 U9268 ( .A1(n10953), .A2(n10952), .ZN(n11100) );
  NAND2_X1 U9269 ( .A1(n7402), .A2(n7400), .ZN(n10788) );
  NAND2_X1 U9270 ( .A1(n7072), .A2(n7071), .ZN(n12037) );
  AOI21_X2 U9271 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n10045), .A(n10031), .ZN(
        n10131) );
  XNOR2_X1 U9272 ( .A(n10701), .B(n10708), .ZN(n10489) );
  NOR2_X1 U9273 ( .A1(n14887), .A2(n14888), .ZN(n14886) );
  XNOR2_X1 U9274 ( .A(n9136), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U9275 ( .A1(n7062), .A2(n7061), .ZN(n12208) );
  AOI21_X1 U9276 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10487), .A(n10486), .ZN(
        n10701) );
  OR2_X1 U9277 ( .A1(n7711), .A2(SI_1_), .ZN(n6833) );
  OR2_X1 U9278 ( .A1(n7796), .A2(n6570), .ZN(n7797) );
  AND2_X1 U9279 ( .A1(n12949), .A2(n12947), .ZN(n12948) );
  NAND2_X1 U9280 ( .A1(n7158), .A2(n7161), .ZN(n13187) );
  NAND4_X1 U9281 ( .A1(n13458), .A2(n13456), .A3(n13455), .A4(n13457), .ZN(
        n13543) );
  INV_X1 U9282 ( .A(n7149), .ZN(n13236) );
  NAND2_X1 U9283 ( .A1(n11140), .A2(n7153), .ZN(n7152) );
  NOR2_X2 U9284 ( .A1(n7668), .A2(n7782), .ZN(n8022) );
  NAND3_X1 U9285 ( .A1(n6999), .A2(n7665), .A3(n7664), .ZN(n7668) );
  NAND2_X1 U9286 ( .A1(n6845), .A2(n6843), .ZN(P3_U3486) );
  OR2_X1 U9287 ( .A1(n12621), .A2(n15029), .ZN(n6845) );
  NAND4_X2 U9288 ( .A1(n7755), .A2(n7754), .A3(n7753), .A4(n7752), .ZN(n13857)
         );
  INV_X1 U9289 ( .A(n7039), .ZN(n12380) );
  NAND2_X1 U9290 ( .A1(n11764), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8511) );
  AND2_X2 U9291 ( .A1(n10802), .A2(n7240), .ZN(n11143) );
  XNOR2_X1 U9292 ( .A(n10131), .B(n10147), .ZN(n10032) );
  NAND2_X1 U9293 ( .A1(n13400), .A2(n12751), .ZN(n13386) );
  NAND2_X1 U9294 ( .A1(n8545), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7046) );
  NAND2_X1 U9295 ( .A1(n9721), .A2(n9722), .ZN(n9720) );
  NOR2_X1 U9296 ( .A1(n10135), .A2(n10134), .ZN(n10486) );
  AND2_X1 U9297 ( .A1(n10527), .A2(n10531), .ZN(n10645) );
  NAND2_X2 U9298 ( .A1(n9346), .A2(n9343), .ZN(n11375) );
  NAND3_X2 U9299 ( .A1(n6860), .A2(n7131), .A3(n6583), .ZN(n9211) );
  INV_X1 U9300 ( .A(n9883), .ZN(n14797) );
  NAND2_X1 U9301 ( .A1(n14539), .A2(n14538), .ZN(n14537) );
  NAND2_X1 U9302 ( .A1(n14517), .A2(n14518), .ZN(n14516) );
  NAND3_X1 U9303 ( .A1(n7198), .A2(n6641), .A3(n7197), .ZN(n13053) );
  NAND2_X1 U9304 ( .A1(n8778), .A2(n8777), .ZN(n8805) );
  NAND2_X1 U9305 ( .A1(n12157), .A2(n12038), .ZN(n12060) );
  NAND2_X1 U9306 ( .A1(n12019), .A2(n7100), .ZN(n12125) );
  NAND2_X1 U9307 ( .A1(n12030), .A2(n7069), .ZN(n12105) );
  INV_X1 U9308 ( .A(n7083), .ZN(n12141) );
  NAND2_X1 U9309 ( .A1(n10102), .A2(n10103), .ZN(n7068) );
  NAND2_X1 U9310 ( .A1(n8833), .A2(n8831), .ZN(n8478) );
  NAND2_X1 U9311 ( .A1(n8459), .A2(n8458), .ZN(n8694) );
  MUX2_X2 U9312 ( .A(n11757), .B(n11756), .S(n11755), .Z(n11781) );
  OAI21_X2 U9313 ( .B1(n11781), .B2(n11823), .A(n11821), .ZN(n11786) );
  NAND2_X1 U9314 ( .A1(n8709), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8465) );
  NAND2_X2 U9315 ( .A1(n8881), .A2(n6854), .ZN(n8891) );
  XNOR2_X1 U9316 ( .A(n7608), .B(n7609), .ZN(n15331) );
  XNOR2_X1 U9317 ( .A(n6855), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9318 ( .A1(n14310), .A2(n14311), .ZN(n6856) );
  NAND2_X1 U9319 ( .A1(n6857), .A2(n7306), .ZN(n12871) );
  NAND3_X1 U9320 ( .A1(n12865), .A2(n12864), .A3(n6644), .ZN(n6857) );
  OAI21_X1 U9321 ( .B1(n12888), .B2(n7305), .A(n6858), .ZN(n12895) );
  INV_X1 U9322 ( .A(n13053), .ZN(n13047) );
  NAND2_X1 U9323 ( .A1(n7300), .A2(n7301), .ZN(n7198) );
  NOR2_X2 U9324 ( .A1(n10076), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n10302) );
  OAI21_X1 U9325 ( .B1(n6570), .B2(n6951), .A(n7829), .ZN(n6950) );
  INV_X2 U9326 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7702) );
  NAND2_X1 U9327 ( .A1(n7826), .A2(n7825), .ZN(n7830) );
  NAND2_X1 U9328 ( .A1(n11302), .A2(n6959), .ZN(n11413) );
  OAI22_X1 U9329 ( .A1(n11100), .A2(n7406), .B1(n7408), .B2(n7407), .ZN(n11301) );
  NAND2_X1 U9330 ( .A1(n8349), .A2(n10792), .ZN(n7694) );
  NAND2_X1 U9331 ( .A1(n6866), .A2(n6865), .ZN(n7770) );
  NAND2_X1 U9332 ( .A1(n7751), .A2(n10364), .ZN(n6866) );
  OAI21_X1 U9333 ( .B1(n6868), .B2(n6867), .A(n7345), .ZN(n8315) );
  NAND3_X1 U9334 ( .A1(n8146), .A2(n8145), .A3(n6646), .ZN(n6873) );
  NAND2_X1 U9335 ( .A1(n7965), .A2(n7966), .ZN(n7964) );
  NAND2_X1 U9336 ( .A1(n6876), .A2(n6875), .ZN(n13875) );
  OR2_X1 U9337 ( .A1(n9599), .A2(n9694), .ZN(n6875) );
  NAND2_X1 U9338 ( .A1(n9599), .A2(n9694), .ZN(n6876) );
  INV_X1 U9339 ( .A(n11610), .ZN(n6880) );
  OAI211_X1 U9340 ( .C1(n7377), .C2(n10194), .A(n6881), .B(n10338), .ZN(n7373)
         );
  NAND2_X2 U9341 ( .A1(n6882), .A2(n9953), .ZN(n10194) );
  NAND2_X1 U9342 ( .A1(n13804), .A2(n6885), .ZN(n6883) );
  NAND2_X1 U9343 ( .A1(n6883), .A2(n6884), .ZN(n13778) );
  NAND2_X1 U9344 ( .A1(n7390), .A2(n6890), .ZN(n6888) );
  NAND2_X1 U9345 ( .A1(n6888), .A2(n6889), .ZN(n13628) );
  NAND2_X1 U9346 ( .A1(n7383), .A2(n6895), .ZN(n6894) );
  NAND2_X1 U9347 ( .A1(n7383), .A2(n7382), .ZN(n13738) );
  OAI211_X1 U9348 ( .C1(n7383), .C2(n6896), .A(n13750), .B(n6894), .ZN(
        P1_U3220) );
  NAND2_X1 U9349 ( .A1(n11020), .A2(n6908), .ZN(n6907) );
  NAND2_X1 U9350 ( .A1(n6907), .A2(n6561), .ZN(n13595) );
  INV_X1 U9351 ( .A(n11160), .ZN(n6912) );
  INV_X1 U9352 ( .A(n11927), .ZN(n6913) );
  NAND2_X2 U9353 ( .A1(n12770), .A2(n11913), .ZN(n11927) );
  NAND2_X1 U9354 ( .A1(n12772), .A2(n12771), .ZN(n12770) );
  OAI21_X1 U9355 ( .B1(n12778), .B2(n6918), .A(n6916), .ZN(n12722) );
  AND2_X1 U9356 ( .A1(n9524), .A2(n6920), .ZN(n6919) );
  NAND2_X1 U9357 ( .A1(n9352), .A2(n9353), .ZN(n9524) );
  INV_X1 U9358 ( .A(n6921), .ZN(n9525) );
  NAND2_X1 U9359 ( .A1(n12786), .A2(n6925), .ZN(n6922) );
  NAND2_X1 U9360 ( .A1(n6923), .A2(n6922), .ZN(n12705) );
  AOI21_X2 U9361 ( .B1(n10283), .B2(n10282), .A(n6928), .ZN(n10287) );
  NAND3_X1 U9362 ( .A1(n6934), .A2(n6931), .A3(n6930), .ZN(n14414) );
  NAND3_X2 U9363 ( .A1(n9146), .A2(n9011), .A3(n6577), .ZN(n9819) );
  OAI211_X1 U9364 ( .C1(n6946), .C2(n6540), .A(n6943), .B(n11103), .ZN(n11106)
         );
  NAND2_X1 U9365 ( .A1(n10629), .A2(n6944), .ZN(n6943) );
  NAND2_X1 U9366 ( .A1(n10629), .A2(n10628), .ZN(n10785) );
  NAND2_X1 U9367 ( .A1(n7796), .A2(n6570), .ZN(n7826) );
  NAND3_X1 U9368 ( .A1(n11311), .A2(n6952), .A3(n6585), .ZN(n6954) );
  NAND3_X1 U9369 ( .A1(n6961), .A2(n6960), .A3(n7200), .ZN(n14096) );
  OR2_X1 U9370 ( .A1(n14254), .A2(n14135), .ZN(n6966) );
  MUX2_X1 U9371 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n6536), .Z(n7743) );
  MUX2_X1 U9372 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6536), .Z(n7758) );
  MUX2_X1 U9373 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6967), .Z(n7781) );
  MUX2_X1 U9374 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6967), .Z(n7827) );
  MUX2_X1 U9375 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6967), .Z(n7849) );
  MUX2_X1 U9376 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6967), .Z(n7873) );
  MUX2_X1 U9377 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n6967), .Z(n7895) );
  MUX2_X1 U9378 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6967), .Z(n7954) );
  MUX2_X1 U9379 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6967), .Z(n7916) );
  MUX2_X1 U9380 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6967), .Z(n7979) );
  MUX2_X1 U9381 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6967), .Z(n8057) );
  MUX2_X1 U9382 ( .A(n10078), .B(n15126), .S(n6967), .Z(n8050) );
  MUX2_X1 U9383 ( .A(n9822), .B(n8462), .S(n6967), .Z(n7996) );
  MUX2_X1 U9384 ( .A(n10081), .B(n15244), .S(n6967), .Z(n8075) );
  MUX2_X1 U9385 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n6967), .Z(n8108) );
  MUX2_X1 U9386 ( .A(n10244), .B(n10240), .S(n6967), .Z(n8084) );
  MUX2_X1 U9387 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6967), .Z(n8129) );
  MUX2_X1 U9388 ( .A(n15216), .B(n11072), .S(n6967), .Z(n8169) );
  MUX2_X1 U9389 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6967), .Z(n8154) );
  MUX2_X1 U9390 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n6967), .Z(n8207) );
  MUX2_X1 U9391 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n6967), .Z(n8206) );
  MUX2_X1 U9392 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6967), .Z(n8226) );
  MUX2_X1 U9393 ( .A(n15291), .B(n15151), .S(n6967), .Z(n8229) );
  MUX2_X1 U9394 ( .A(n15117), .B(n8483), .S(n9345), .Z(n8260) );
  MUX2_X1 U9395 ( .A(n13579), .B(n14303), .S(n9345), .Z(n8282) );
  MUX2_X1 U9396 ( .A(n11988), .B(n11568), .S(n9345), .Z(n8287) );
  MUX2_X1 U9397 ( .A(n13570), .B(n14301), .S(n9345), .Z(n8306) );
  NAND2_X1 U9398 ( .A1(n14069), .A2(n6632), .ZN(n6969) );
  NAND2_X1 U9399 ( .A1(n6973), .A2(n7222), .ZN(n14035) );
  NAND2_X1 U9400 ( .A1(n7222), .A2(n14047), .ZN(n6972) );
  OAI21_X2 U9401 ( .B1(n10276), .B2(n6531), .A(n7880), .ZN(n11030) );
  NAND3_X1 U9402 ( .A1(n6987), .A2(n6988), .A3(n6986), .ZN(n14881) );
  NAND3_X1 U9403 ( .A1(n6987), .A2(n6565), .A3(n6986), .ZN(n6989) );
  INV_X1 U9404 ( .A(n6989), .ZN(n14880) );
  NOR2_X2 U9405 ( .A1(n12257), .A2(n15185), .ZN(n12278) );
  NAND2_X1 U9406 ( .A1(n12255), .A2(n6675), .ZN(n6990) );
  AND2_X1 U9407 ( .A1(n14011), .A2(n7008), .ZN(n13983) );
  OR2_X1 U9408 ( .A1(n14011), .A2(n7005), .ZN(n7004) );
  NAND2_X1 U9409 ( .A1(n14011), .A2(n14189), .ZN(n13984) );
  NAND3_X1 U9410 ( .A1(n7004), .A2(n7002), .A3(n7000), .ZN(n14169) );
  NAND2_X1 U9411 ( .A1(n7013), .A2(n10386), .ZN(n10575) );
  OR2_X1 U9412 ( .A1(n12381), .A2(n7036), .ZN(n7032) );
  NAND3_X1 U9413 ( .A1(n7032), .A2(n7031), .A3(n7033), .ZN(n12369) );
  NAND2_X1 U9414 ( .A1(n12381), .A2(n7037), .ZN(n7031) );
  INV_X2 U9415 ( .A(n12373), .ZN(n7038) );
  MUX2_X1 U9416 ( .A(n12552), .B(n7040), .S(n15031), .Z(n12553) );
  MUX2_X1 U9417 ( .A(n12618), .B(n7040), .S(n15019), .Z(n12619) );
  NAND2_X1 U9418 ( .A1(n6516), .A2(n8427), .ZN(n8949) );
  AND3_X2 U9420 ( .A1(n7047), .A2(n7046), .A3(n7045), .ZN(n9136) );
  NAND2_X1 U9421 ( .A1(n7053), .A2(n7051), .ZN(n9811) );
  AND2_X1 U9422 ( .A1(n7052), .A2(n7054), .ZN(n7051) );
  NAND2_X1 U9423 ( .A1(n9833), .A2(n7059), .ZN(n7058) );
  NAND2_X1 U9424 ( .A1(n9833), .A2(n6647), .ZN(n7053) );
  NAND2_X1 U9425 ( .A1(n7055), .A2(n9813), .ZN(n7054) );
  INV_X1 U9426 ( .A(n7059), .ZN(n7055) );
  INV_X1 U9427 ( .A(n7057), .ZN(n9810) );
  NAND2_X1 U9428 ( .A1(n7058), .A2(n9813), .ZN(n7056) );
  INV_X1 U9429 ( .A(n9142), .ZN(n7060) );
  OR2_X2 U9430 ( .A1(n14871), .A2(n8687), .ZN(n7063) );
  OAI211_X1 U9431 ( .C1(n12244), .C2(n6668), .A(n12308), .B(n6542), .ZN(n12309) );
  NAND2_X1 U9432 ( .A1(n6574), .A2(n12610), .ZN(n7064) );
  NAND2_X1 U9433 ( .A1(n6574), .A2(n12244), .ZN(n7065) );
  INV_X1 U9434 ( .A(n7067), .ZN(n12263) );
  NAND2_X1 U9435 ( .A1(n10231), .A2(n7068), .ZN(n10330) );
  OAI21_X1 U9436 ( .B1(n10103), .B2(n10102), .A(n7068), .ZN(n10104) );
  AOI21_X1 U9437 ( .B1(n7068), .B2(n10233), .A(n10232), .ZN(n10234) );
  NAND2_X1 U9438 ( .A1(n12105), .A2(n12034), .ZN(n12036) );
  INV_X1 U9439 ( .A(n12035), .ZN(n7071) );
  INV_X1 U9440 ( .A(n12036), .ZN(n7072) );
  AND2_X1 U9441 ( .A1(n10844), .A2(n7082), .ZN(n7081) );
  NOR2_X2 U9442 ( .A1(n8424), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U9443 ( .A1(n11493), .A2(n7101), .ZN(n12019) );
  INV_X1 U9444 ( .A(n13016), .ZN(n7104) );
  NAND2_X1 U9445 ( .A1(n10642), .A2(n7103), .ZN(n10766) );
  NAND2_X1 U9446 ( .A1(n13170), .A2(n7110), .ZN(n7109) );
  OAI21_X2 U9447 ( .B1(n13170), .B2(n7108), .A(n7105), .ZN(n13224) );
  OAI21_X1 U9448 ( .B1(n11558), .B2(n7123), .A(n7122), .ZN(n11561) );
  INV_X2 U9449 ( .A(n7129), .ZN(n13007) );
  NAND2_X1 U9450 ( .A1(n9877), .A2(n9870), .ZN(n7129) );
  INV_X1 U9451 ( .A(n9019), .ZN(n9015) );
  NAND2_X1 U9452 ( .A1(n13283), .A2(n13268), .ZN(n13194) );
  AOI21_X1 U9453 ( .B1(n10647), .B2(n7136), .A(n6618), .ZN(n7134) );
  NAND2_X1 U9454 ( .A1(n13019), .A2(n7140), .ZN(n7139) );
  NAND2_X1 U9455 ( .A1(n13271), .A2(n13196), .ZN(n13251) );
  NAND2_X1 U9456 ( .A1(n7146), .A2(n7150), .ZN(n13200) );
  NAND2_X1 U9457 ( .A1(n13271), .A2(n7147), .ZN(n7146) );
  NAND2_X1 U9458 ( .A1(n13179), .A2(n7159), .ZN(n7158) );
  NAND2_X1 U9459 ( .A1(n12975), .A2(n12974), .ZN(n12979) );
  NAND2_X1 U9460 ( .A1(n7998), .A2(n7187), .ZN(n7184) );
  NAND2_X1 U9461 ( .A1(n7184), .A2(n7185), .ZN(n8077) );
  NAND2_X1 U9462 ( .A1(n7998), .A2(n7997), .ZN(n8056) );
  NAND2_X1 U9463 ( .A1(n12994), .A2(n13000), .ZN(n7197) );
  NAND2_X1 U9464 ( .A1(n10203), .A2(n10181), .ZN(n10518) );
  NOR2_X1 U9465 ( .A1(n9211), .A2(n7331), .ZN(n9319) );
  AOI21_X2 U9466 ( .B1(n13335), .B2(n13188), .A(n13163), .ZN(n13327) );
  NAND2_X1 U9467 ( .A1(n11011), .A2(n11010), .ZN(n11150) );
  AOI21_X2 U9468 ( .B1(n12311), .B2(n12310), .A(n12331), .ZN(n12312) );
  NAND2_X1 U9469 ( .A1(n8211), .A2(n8210), .ZN(n8225) );
  NAND2_X1 U9470 ( .A1(n7526), .A2(n6564), .ZN(n8727) );
  NAND2_X4 U9471 ( .A1(n9986), .A2(n9985), .ZN(n12095) );
  NAND4_X1 U9472 ( .A1(n7763), .A2(n10018), .A3(n10021), .A4(n7204), .ZN(
        n10362) );
  INV_X1 U9473 ( .A(n10012), .ZN(n10364) );
  NAND2_X1 U9474 ( .A1(n10362), .A2(n10021), .ZN(n10380) );
  OR2_X1 U9475 ( .A1(n9915), .A2(n12824), .ZN(n10215) );
  NOR2_X2 U9476 ( .A1(n10122), .A2(n12813), .ZN(n10125) );
  INV_X1 U9477 ( .A(n7225), .ZN(n14067) );
  INV_X1 U9478 ( .A(n7668), .ZN(n7227) );
  NAND2_X1 U9479 ( .A1(n7226), .A2(n7670), .ZN(n8404) );
  NOR2_X2 U9480 ( .A1(n6569), .A2(n13276), .ZN(n13275) );
  NAND2_X1 U9481 ( .A1(n13242), .A2(n7231), .ZN(n13149) );
  NAND2_X1 U9482 ( .A1(n13242), .A2(n13542), .ZN(n13231) );
  NAND2_X1 U9483 ( .A1(n7536), .A2(n7235), .ZN(n9381) );
  NAND2_X1 U9484 ( .A1(n7236), .A2(n9346), .ZN(n7235) );
  OAI21_X1 U9485 ( .B1(n9344), .B2(n6967), .A(n6653), .ZN(n7236) );
  NOR2_X2 U9486 ( .A1(n13401), .A2(n13514), .ZN(n13400) );
  NAND2_X1 U9487 ( .A1(n7239), .A2(n10812), .ZN(n7243) );
  NOR2_X1 U9488 ( .A1(n7243), .A2(n14844), .ZN(n7240) );
  INV_X1 U9489 ( .A(n9349), .ZN(n9744) );
  NAND2_X2 U9490 ( .A1(n9875), .A2(n6571), .ZN(n9349) );
  NAND2_X1 U9491 ( .A1(n7247), .A2(n7245), .ZN(n12754) );
  NAND2_X2 U9492 ( .A1(n12733), .A2(n12735), .ZN(n12734) );
  NAND2_X1 U9493 ( .A1(n7255), .A2(n7251), .ZN(n7254) );
  INV_X1 U9494 ( .A(n14653), .ZN(n7251) );
  NAND3_X1 U9495 ( .A1(n7260), .A2(n7259), .A3(n7265), .ZN(n11521) );
  NAND2_X1 U9496 ( .A1(n11985), .A2(n7269), .ZN(n7268) );
  OAI211_X1 U9497 ( .C1(n11985), .C2(n7270), .A(n7268), .B(n12013), .ZN(
        P2_U3192) );
  NAND2_X1 U9498 ( .A1(n7284), .A2(n7282), .ZN(n7281) );
  CLKBUF_X1 U9499 ( .A(n7284), .Z(n7277) );
  NAND2_X2 U9500 ( .A1(n7281), .A2(n7279), .ZN(n12780) );
  NAND2_X1 U9501 ( .A1(n12795), .A2(n11531), .ZN(n11532) );
  INV_X1 U9502 ( .A(n7277), .ZN(n12742) );
  INV_X1 U9503 ( .A(n11533), .ZN(n7285) );
  NAND2_X1 U9504 ( .A1(n9331), .A2(n6633), .ZN(n7286) );
  NAND2_X1 U9505 ( .A1(n7291), .A2(n7290), .ZN(n7289) );
  INV_X1 U9506 ( .A(n12899), .ZN(n7290) );
  INV_X1 U9507 ( .A(n7294), .ZN(n7291) );
  NAND2_X1 U9508 ( .A1(n7293), .A2(n12898), .ZN(n7292) );
  NAND2_X1 U9509 ( .A1(n7294), .A2(n12899), .ZN(n7293) );
  NAND2_X1 U9510 ( .A1(n12810), .A2(n12812), .ZN(n7296) );
  NAND3_X1 U9511 ( .A1(n7298), .A2(n12808), .A3(n12810), .ZN(n7295) );
  NAND3_X1 U9512 ( .A1(n12812), .A2(n12808), .A3(n7298), .ZN(n7297) );
  NAND2_X1 U9513 ( .A1(n7299), .A2(n6648), .ZN(n7298) );
  INV_X1 U9514 ( .A(n12809), .ZN(n7299) );
  NAND2_X1 U9515 ( .A1(n12938), .A2(n12939), .ZN(n7301) );
  NAND2_X1 U9516 ( .A1(n7302), .A2(n6640), .ZN(n12892) );
  NAND2_X1 U9517 ( .A1(n12888), .A2(n7304), .ZN(n7302) );
  NAND3_X1 U9518 ( .A1(n12914), .A2(n12913), .A3(n6645), .ZN(n7308) );
  INV_X1 U9519 ( .A(n12916), .ZN(n7310) );
  OR2_X1 U9520 ( .A1(n12821), .A2(n12823), .ZN(n7312) );
  NAND2_X1 U9521 ( .A1(n7311), .A2(n7313), .ZN(n12827) );
  NAND2_X1 U9522 ( .A1(n7314), .A2(n7315), .ZN(n12927) );
  NAND2_X1 U9523 ( .A1(n12925), .A2(n7317), .ZN(n7314) );
  NAND2_X1 U9524 ( .A1(n7321), .A2(n7322), .ZN(n12882) );
  NAND2_X1 U9525 ( .A1(n12879), .A2(n7324), .ZN(n7321) );
  NAND3_X1 U9526 ( .A1(n9213), .A2(n7332), .A3(n9212), .ZN(n7331) );
  NAND2_X1 U9527 ( .A1(n12933), .A2(n7336), .ZN(n7333) );
  OAI21_X1 U9528 ( .B1(n12933), .B2(n7338), .A(n7336), .ZN(n12937) );
  NAND2_X1 U9529 ( .A1(n7333), .A2(n7334), .ZN(n12935) );
  NAND2_X1 U9530 ( .A1(n7694), .A2(n9511), .ZN(n7351) );
  NAND3_X1 U9531 ( .A1(n7694), .A2(n9511), .A3(n10973), .ZN(n7352) );
  NAND2_X1 U9532 ( .A1(n7366), .A2(n8025), .ZN(n7690) );
  NAND2_X1 U9533 ( .A1(n9703), .A2(n7368), .ZN(n9697) );
  OR2_X1 U9534 ( .A1(n9696), .A2(n7369), .ZN(n7368) );
  NAND2_X1 U9535 ( .A1(n7369), .A2(n9696), .ZN(n9703) );
  NOR2_X1 U9536 ( .A1(n9693), .A2(n9701), .ZN(n7369) );
  OAI211_X2 U9537 ( .C1(n7373), .C2(n10601), .A(n10600), .B(n7372), .ZN(n10609) );
  NAND2_X1 U9538 ( .A1(n7379), .A2(n7381), .ZN(n7378) );
  INV_X1 U9539 ( .A(n10193), .ZN(n7379) );
  NAND2_X1 U9540 ( .A1(n13770), .A2(n7385), .ZN(n7383) );
  OR2_X2 U9541 ( .A1(n13595), .A2(n7391), .ZN(n7390) );
  NAND2_X1 U9542 ( .A1(n13831), .A2(n6600), .ZN(n7394) );
  OAI211_X1 U9543 ( .C1(n13634), .C2(n7395), .A(n7394), .B(n14454), .ZN(n13647) );
  INV_X1 U9544 ( .A(n13639), .ZN(n7395) );
  NAND2_X1 U9545 ( .A1(n14446), .A2(n13639), .ZN(n14455) );
  NAND2_X1 U9546 ( .A1(n13634), .A2(n14442), .ZN(n14446) );
  NAND2_X1 U9547 ( .A1(n7396), .A2(n6643), .ZN(n13726) );
  INV_X1 U9548 ( .A(n7401), .ZN(n7400) );
  OAI21_X1 U9549 ( .B1(n7405), .B2(n10666), .A(n10627), .ZN(n7401) );
  NAND2_X1 U9550 ( .A1(n10617), .A2(n7403), .ZN(n7402) );
  INV_X1 U9551 ( .A(n11308), .ZN(n7407) );
  NAND2_X1 U9552 ( .A1(n14133), .A2(n6587), .ZN(n7413) );
  NAND2_X1 U9553 ( .A1(n14050), .A2(n6636), .ZN(n7423) );
  INV_X1 U9554 ( .A(n7427), .ZN(n14045) );
  OR2_X1 U9555 ( .A1(n14216), .A2(n13842), .ZN(n7428) );
  XNOR2_X2 U9556 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8517) );
  NAND2_X1 U9557 ( .A1(n8752), .A2(n7433), .ZN(n7431) );
  NAND2_X1 U9558 ( .A1(n7431), .A2(n7432), .ZN(n8474) );
  OR2_X1 U9559 ( .A1(n8891), .A2(n7448), .ZN(n7441) );
  NAND2_X1 U9560 ( .A1(n8891), .A2(n6674), .ZN(n7444) );
  NAND2_X1 U9561 ( .A1(n8891), .A2(n8890), .ZN(n7449) );
  OAI21_X1 U9562 ( .B1(n8621), .B2(n7452), .A(n7450), .ZN(n8654) );
  NAND2_X1 U9563 ( .A1(n8726), .A2(n7463), .ZN(n7460) );
  NAND2_X1 U9564 ( .A1(n8551), .A2(n10425), .ZN(n11636) );
  NAND2_X1 U9565 ( .A1(n7472), .A2(n10907), .ZN(n7476) );
  NOR2_X1 U9566 ( .A1(n7473), .A2(n7546), .ZN(n7472) );
  NAND2_X1 U9567 ( .A1(n7476), .A2(n7474), .ZN(n11048) );
  OR2_X1 U9568 ( .A1(n7546), .A2(n8931), .ZN(n7479) );
  NAND2_X1 U9569 ( .A1(n7480), .A2(n11789), .ZN(n7477) );
  NAND2_X1 U9570 ( .A1(n8933), .A2(n7485), .ZN(n7482) );
  NAND2_X1 U9571 ( .A1(n7492), .A2(n6562), .ZN(n12516) );
  OAI21_X1 U9572 ( .B1(n12420), .B2(n7496), .A(n7493), .ZN(n7500) );
  NAND2_X1 U9573 ( .A1(n12420), .A2(n8942), .ZN(n12398) );
  OAI21_X1 U9574 ( .B1(n14365), .B2(n7504), .A(n7502), .ZN(n8934) );
  NAND2_X1 U9575 ( .A1(n7522), .A2(n8529), .ZN(n14943) );
  AND2_X1 U9576 ( .A1(n8528), .A2(n10255), .ZN(n7522) );
  AND2_X1 U9577 ( .A1(n7524), .A2(n7523), .ZN(n7525) );
  INV_X1 U9578 ( .A(n8618), .ZN(n7526) );
  NAND2_X1 U9579 ( .A1(n13007), .A2(n9933), .ZN(n9932) );
  INV_X1 U9580 ( .A(n9381), .ZN(n9348) );
  XNOR2_X1 U9581 ( .A(n9349), .B(n9348), .ZN(n9352) );
  INV_X1 U9582 ( .A(n11156), .ZN(n11021) );
  OR2_X1 U9583 ( .A1(n8269), .A2(n9395), .ZN(n7684) );
  XNOR2_X1 U9584 ( .A(n13628), .B(n13626), .ZN(n13831) );
  AND2_X1 U9585 ( .A1(n9536), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7549) );
  OR2_X1 U9586 ( .A1(n14187), .A2(n14623), .ZN(n14194) );
  CLKBUF_X1 U9587 ( .A(n9211), .Z(n9026) );
  NOR2_X1 U9588 ( .A1(n7535), .A2(n7549), .ZN(n9326) );
  NOR2_X2 U9589 ( .A1(n9533), .A2(n9532), .ZN(n9646) );
  AND2_X1 U9590 ( .A1(n9692), .A2(n9691), .ZN(n9693) );
  NAND2_X1 U9591 ( .A1(n7678), .A2(n7677), .ZN(n7865) );
  OAI21_X1 U9592 ( .B1(n8991), .B2(n15018), .A(n8988), .ZN(n8990) );
  INV_X1 U9593 ( .A(n12507), .ZN(n12508) );
  OR2_X1 U9594 ( .A1(n14124), .A2(n14137), .ZN(n7532) );
  OR2_X1 U9595 ( .A1(n11572), .A2(n12612), .ZN(n7533) );
  OR2_X1 U9596 ( .A1(n11572), .A2(n12669), .ZN(n7534) );
  INV_X1 U9597 ( .A(n15031), .ZN(n15029) );
  INV_X2 U9598 ( .A(n15018), .ZN(n15019) );
  INV_X2 U9599 ( .A(n14955), .ZN(n14957) );
  INV_X1 U9600 ( .A(n9649), .ZN(n9650) );
  AND2_X1 U9601 ( .A1(n9534), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7535) );
  OR2_X1 U9602 ( .A1(n9346), .A2(n13082), .ZN(n7536) );
  INV_X1 U9603 ( .A(n11806), .ZN(n12517) );
  OR2_X1 U9604 ( .A1(n14855), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7537) );
  OR2_X1 U9605 ( .A1(n14861), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7538) );
  INV_X1 U9606 ( .A(n14855), .ZN(n13539) );
  INV_X1 U9607 ( .A(n14861), .ZN(n13449) );
  OR2_X2 U9608 ( .A1(n13441), .A2(n13440), .ZN(n7541) );
  AND3_X1 U9609 ( .A1(n9330), .A2(n9329), .A3(n10079), .ZN(n7543) );
  AND2_X1 U9610 ( .A1(n8054), .A2(n8053), .ZN(n7545) );
  NOR2_X1 U9611 ( .A1(n8930), .A2(n11794), .ZN(n7546) );
  AND2_X1 U9612 ( .A1(n9063), .A2(n9056), .ZN(n7547) );
  INV_X1 U9613 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7710) );
  INV_X1 U9614 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11072) );
  AND2_X1 U9615 ( .A1(n9825), .A2(n9047), .ZN(n7548) );
  INV_X1 U9616 ( .A(n14440), .ZN(n11584) );
  INV_X1 U9617 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n15216) );
  AND2_X1 U9618 ( .A1(n9384), .A2(n9387), .ZN(n13405) );
  AND2_X1 U9619 ( .A1(n7931), .A2(n7930), .ZN(n7550) );
  INV_X1 U9620 ( .A(n14074), .ZN(n11600) );
  AND2_X1 U9621 ( .A1(n8702), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7551) );
  INV_X1 U9622 ( .A(n12483), .ZN(n8936) );
  AND2_X1 U9623 ( .A1(n7683), .A2(n7682), .ZN(n7554) );
  AND2_X1 U9624 ( .A1(n8383), .A2(n8382), .ZN(n7555) );
  NAND2_X1 U9625 ( .A1(n8376), .A2(n10021), .ZN(n7764) );
  AND2_X1 U9626 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  INV_X1 U9627 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9009) );
  INV_X1 U9628 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8425) );
  INV_X1 U9629 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9006) );
  INV_X1 U9630 ( .A(n8051), .ZN(n8054) );
  INV_X1 U9631 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9016) );
  INV_X1 U9632 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15082) );
  INV_X1 U9633 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10154) );
  INV_X1 U9634 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8641) );
  INV_X1 U9635 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U9636 ( .A1(n10870), .A2(n8626), .ZN(n10963) );
  INV_X1 U9637 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8483) );
  INV_X1 U9638 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9857) );
  OR2_X1 U9639 ( .A1(n13504), .A2(n13180), .ZN(n13181) );
  AND2_X1 U9640 ( .A1(n13439), .A2(n14843), .ZN(n13440) );
  INV_X1 U9641 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9318) );
  INV_X1 U9642 ( .A(n9957), .ZN(n9954) );
  INV_X1 U9643 ( .A(n13741), .ZN(n10605) );
  INV_X1 U9644 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7839) );
  INV_X1 U9645 ( .A(n13852), .ZN(n10679) );
  AND2_X1 U9646 ( .A1(n8844), .A2(n8412), .ZN(n8846) );
  OR2_X1 U9647 ( .A1(n8812), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8824) );
  OR2_X1 U9648 ( .A1(n14352), .A2(n8885), .ZN(n12375) );
  NAND2_X1 U9649 ( .A1(n8796), .A2(n15188), .ZN(n8812) );
  OR3_X1 U9650 ( .A1(n11817), .A2(n10110), .A3(n8998), .ZN(n8996) );
  NAND2_X1 U9651 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n11568), .ZN(n8892) );
  NAND2_X1 U9652 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n11072), .ZN(n8477) );
  OR2_X1 U9653 ( .A1(n11874), .A2(n11873), .ZN(n11881) );
  NAND2_X1 U9654 ( .A1(n10741), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10752) );
  AND2_X1 U9655 ( .A1(n14428), .A2(n14429), .ZN(n13618) );
  INV_X1 U9656 ( .A(n11017), .ZN(n11018) );
  OR2_X1 U9657 ( .A1(n13598), .A2(n13597), .ZN(n13599) );
  NAND2_X1 U9658 ( .A1(n10192), .A2(n10191), .ZN(n10193) );
  INV_X1 U9659 ( .A(n13606), .ZN(n13607) );
  INV_X1 U9660 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n15138) );
  INV_X1 U9661 ( .A(n8217), .ZN(n8218) );
  INV_X1 U9662 ( .A(n14554), .ZN(n10827) );
  NAND2_X1 U9663 ( .A1(n13982), .A2(n14003), .ZN(n13995) );
  AND2_X1 U9664 ( .A1(n14074), .A2(n13843), .ZN(n11581) );
  INV_X1 U9665 ( .A(n14254), .ZN(n11599) );
  INV_X1 U9666 ( .A(n11103), .ZN(n10952) );
  INV_X1 U9667 ( .A(n9592), .ZN(n9591) );
  NAND2_X1 U9668 ( .A1(n11305), .A2(n14492), .ZN(n11420) );
  INV_X1 U9669 ( .A(n10581), .ZN(n10447) );
  NOR2_X1 U9670 ( .A1(n10402), .A2(n10374), .ZN(n10386) );
  INV_X1 U9671 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8388) );
  NOR2_X1 U9672 ( .A1(n7632), .A2(n7631), .ZN(n7569) );
  NOR2_X1 U9673 ( .A1(n7598), .A2(n7597), .ZN(n7577) );
  NAND2_X1 U9674 ( .A1(n8846), .A2(n8500), .ZN(n8502) );
  OR2_X1 U9675 ( .A1(n8858), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8869) );
  AND2_X1 U9676 ( .A1(n8783), .A2(n12129), .ZN(n8796) );
  INV_X1 U9677 ( .A(n14862), .ZN(n14883) );
  AND2_X1 U9678 ( .A1(n8870), .A2(n12055), .ZN(n8884) );
  INV_X1 U9679 ( .A(n11804), .ZN(n12531) );
  INV_X1 U9680 ( .A(n12537), .ZN(n11490) );
  INV_X1 U9681 ( .A(n11799), .ZN(n8707) );
  INV_X1 U9682 ( .A(n6525), .ZN(n11817) );
  INV_X1 U9683 ( .A(n12672), .ZN(n9000) );
  INV_X1 U9684 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8987) );
  AND2_X1 U9685 ( .A1(n11692), .A2(n11693), .ZN(n14364) );
  INV_X1 U9686 ( .A(n14967), .ZN(n14978) );
  XNOR2_X1 U9687 ( .A(n9162), .B(P1_DATAO_REG_6__SCAN_IN), .ZN(n8599) );
  INV_X1 U9688 ( .A(n12700), .ZN(n11984) );
  INV_X1 U9689 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10296) );
  INV_X1 U9690 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n14648) );
  NOR2_X1 U9691 ( .A1(n11881), .A2(n12729), .ZN(n11902) );
  AND2_X1 U9692 ( .A1(n11534), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11550) );
  INV_X1 U9693 ( .A(n13311), .ZN(n13273) );
  INV_X1 U9694 ( .A(n13405), .ZN(n13318) );
  INV_X1 U9695 ( .A(n13028), .ZN(n11560) );
  INV_X1 U9696 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U9697 ( .A1(n7948), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8012) );
  INV_X1 U9698 ( .A(n13724), .ZN(n13657) );
  NAND2_X1 U9699 ( .A1(n11016), .A2(n11018), .ZN(n11019) );
  NOR2_X1 U9700 ( .A1(n8114), .A2(n15168), .ZN(n8148) );
  INV_X1 U9701 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7930) );
  INV_X1 U9702 ( .A(n14457), .ZN(n14471) );
  OR3_X1 U9703 ( .A1(n9585), .A2(n10306), .A3(n9584), .ZN(n9607) );
  NOR2_X1 U9704 ( .A1(n8029), .A2(n15138), .ZN(n8044) );
  AND2_X1 U9705 ( .A1(n8162), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8178) );
  OR2_X1 U9706 ( .A1(n8094), .A2(n8093), .ZN(n8114) );
  AND2_X1 U9707 ( .A1(n9630), .A2(n9621), .ZN(n9622) );
  INV_X1 U9708 ( .A(n14195), .ZN(n14012) );
  NOR2_X1 U9709 ( .A1(n11475), .A2(n11476), .ZN(n11586) );
  INV_X1 U9710 ( .A(n13846), .ZN(n14427) );
  INV_X1 U9711 ( .A(n14609), .ZN(n14617) );
  OR2_X1 U9712 ( .A1(n10315), .A2(n10792), .ZN(n14010) );
  XNOR2_X1 U9713 ( .A(n7954), .B(SI_11_), .ZN(n7957) );
  OAI21_X1 U9714 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n15294), .A(n7580), .ZN(
        n7593) );
  AND2_X1 U9715 ( .A1(n9078), .A2(n9077), .ZN(n9102) );
  INV_X1 U9716 ( .A(n14347), .ZN(n12195) );
  OR2_X1 U9717 ( .A1(n8731), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8763) );
  AOI21_X1 U9718 ( .B1(n12390), .B2(n8897), .A(n8439), .ZN(n12193) );
  AND4_X1 U9719 ( .A1(n8736), .A2(n8735), .A3(n8734), .A4(n8733), .ZN(n14337)
         );
  INV_X1 U9720 ( .A(n9083), .ZN(n9099) );
  INV_X1 U9721 ( .A(n14903), .ZN(n12307) );
  AND2_X1 U9722 ( .A1(n9102), .A2(n9100), .ZN(n9083) );
  INV_X1 U9723 ( .A(n14932), .ZN(n14946) );
  INV_X1 U9724 ( .A(n11053), .ZN(n14379) );
  INV_X1 U9725 ( .A(n14354), .ZN(n14919) );
  AND3_X1 U9726 ( .A1(n8995), .A2(n8994), .A3(n8993), .ZN(n10251) );
  AND2_X1 U9727 ( .A1(n14967), .A2(n15006), .ZN(n12617) );
  INV_X1 U9728 ( .A(n15013), .ZN(n14980) );
  INV_X1 U9729 ( .A(n15006), .ZN(n14992) );
  INV_X1 U9730 ( .A(n14930), .ZN(n14944) );
  XNOR2_X1 U9731 ( .A(n8906), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11836) );
  NAND2_X1 U9732 ( .A1(n8474), .A2(n8473), .ZN(n8804) );
  AND2_X1 U9733 ( .A1(n8450), .A2(n8449), .ZN(n8587) );
  AND2_X1 U9734 ( .A1(n10508), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10741) );
  INV_X1 U9735 ( .A(n14660), .ZN(n12800) );
  AND3_X1 U9736 ( .A1(n12944), .A2(n12943), .A3(n12942), .ZN(n13145) );
  AND2_X1 U9737 ( .A1(n11909), .A2(n11908), .ZN(n13310) );
  INV_X1 U9738 ( .A(n12004), .ZN(n11887) );
  NOR2_X1 U9739 ( .A1(n10089), .A2(n14730), .ZN(n14753) );
  AND2_X1 U9740 ( .A1(n9248), .A2(n13044), .ZN(n14776) );
  INV_X1 U9741 ( .A(n13188), .ZN(n13338) );
  AND2_X1 U9742 ( .A1(n9223), .A2(n9387), .ZN(n13407) );
  INV_X1 U9743 ( .A(n14789), .ZN(n13425) );
  INV_X1 U9744 ( .A(n13396), .ZN(n14792) );
  INV_X1 U9745 ( .A(n14837), .ZN(n14843) );
  NOR2_X1 U9746 ( .A1(n14818), .A2(n9888), .ZN(n10258) );
  AND2_X1 U9747 ( .A1(n11357), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9357) );
  AND2_X1 U9748 ( .A1(n8044), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8067) );
  AND3_X1 U9749 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n7819) );
  INV_X1 U9750 ( .A(n14476), .ZN(n14464) );
  AND4_X1 U9751 ( .A1(n8018), .A2(n8017), .A3(n8016), .A4(n8015), .ZN(n13833)
         );
  OR2_X1 U9752 ( .A1(n9629), .A2(n9628), .ZN(n9630) );
  INV_X1 U9753 ( .A(n14552), .ZN(n14563) );
  INV_X1 U9754 ( .A(n14138), .ZN(n14152) );
  INV_X1 U9755 ( .A(n10786), .ZN(n10945) );
  INV_X1 U9756 ( .A(n10453), .ZN(n10456) );
  INV_X1 U9757 ( .A(n14161), .ZN(n14110) );
  OR2_X1 U9758 ( .A1(n10307), .A2(n9585), .ZN(n9600) );
  INV_X1 U9759 ( .A(n14615), .ZN(n14623) );
  NAND2_X1 U9760 ( .A1(n14010), .A2(n14219), .ZN(n14615) );
  INV_X1 U9761 ( .A(n9585), .ZN(n10308) );
  XNOR2_X1 U9762 ( .A(n8391), .B(n8390), .ZN(n9315) );
  NAND2_X1 U9763 ( .A1(n9792), .A2(n9794), .ZN(n12174) );
  INV_X1 U9764 ( .A(n12020), .ZN(n12538) );
  INV_X1 U9765 ( .A(n9139), .ZN(n9774) );
  INV_X1 U9766 ( .A(n12362), .ZN(n14897) );
  AND2_X1 U9767 ( .A1(n12527), .A2(n12526), .ZN(n12599) );
  NAND2_X1 U9768 ( .A1(n9795), .A2(n9794), .ZN(n14926) );
  NAND2_X1 U9769 ( .A1(n10252), .A2(n14926), .ZN(n14955) );
  AND2_X2 U9770 ( .A1(n10251), .A2(n9002), .ZN(n15031) );
  AND4_X1 U9771 ( .A1(n14985), .A2(n14984), .A3(n14983), .A4(n14982), .ZN(
        n15024) );
  AND2_X2 U9772 ( .A1(n8986), .A2(n8985), .ZN(n15018) );
  INV_X1 U9773 ( .A(n11633), .ZN(n10418) );
  INV_X1 U9774 ( .A(SI_12_), .ZN(n15171) );
  NAND2_X1 U9775 ( .A1(n9647), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14660) );
  INV_X1 U9776 ( .A(n14657), .ZN(n14415) );
  NAND2_X1 U9777 ( .A1(n9376), .A2(n9375), .ZN(n14652) );
  INV_X1 U9778 ( .A(n14420), .ZN(n13406) );
  INV_X1 U9779 ( .A(n14770), .ZN(n14740) );
  OR2_X1 U9780 ( .A1(n9225), .A2(n13044), .ZN(n14747) );
  NAND2_X1 U9781 ( .A1(n14809), .A2(n9919), .ZN(n13390) );
  NAND2_X1 U9782 ( .A1(n14809), .A2(n9907), .ZN(n13396) );
  AND2_X2 U9783 ( .A1(n10258), .A2(n9889), .ZN(n14861) );
  AND4_X1 U9784 ( .A1(n14853), .A2(n14852), .A3(n14851), .A4(n14850), .ZN(
        n14860) );
  AND3_X1 U9785 ( .A1(n14842), .A2(n14841), .A3(n14840), .ZN(n14859) );
  NOR2_X1 U9786 ( .A1(n14820), .A2(n14812), .ZN(n14813) );
  INV_X1 U9787 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10078) );
  INV_X1 U9788 ( .A(n14249), .ZN(n14143) );
  INV_X1 U9789 ( .A(n14244), .ZN(n14124) );
  INV_X1 U9790 ( .A(n13610), .ZN(n14497) );
  NAND2_X1 U9791 ( .A1(n9958), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14485) );
  OR2_X1 U9792 ( .A1(n14546), .A2(n14542), .ZN(n14557) );
  OR2_X1 U9793 ( .A1(n14546), .A2(n13878), .ZN(n14571) );
  INV_X1 U9794 ( .A(n14544), .ZN(n14575) );
  AND2_X1 U9795 ( .A1(n14121), .A2(n14120), .ZN(n14247) );
  AND2_X1 U9796 ( .A1(n10949), .A2(n10948), .ZN(n14509) );
  INV_X1 U9797 ( .A(n14114), .ZN(n14164) );
  OR2_X1 U9798 ( .A1(n9600), .A2(n9517), .ZN(n14634) );
  AND2_X1 U9799 ( .A1(n14509), .A2(n14508), .ZN(n14515) );
  OR3_X1 U9800 ( .A1(n9517), .A2(n10308), .A3(n10307), .ZN(n14625) );
  AND2_X1 U9801 ( .A1(n9315), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9175) );
  INV_X1 U9802 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10240) );
  INV_X1 U9803 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9580) );
  AND2_X2 U9804 ( .A1(n9032), .A2(n12673), .ZN(P3_U3897) );
  NOR2_X1 U9805 ( .A1(n9388), .A2(n9031), .ZN(P2_U3947) );
  INV_X1 U9806 ( .A(n13856), .ZN(P1_U4016) );
  XNOR2_X1 U9807 ( .A(n7660), .B(n7659), .ZN(SUB_1596_U4) );
  INV_X1 U9808 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15085) );
  XNOR2_X1 U9809 ( .A(n15085), .B(P3_ADDR_REG_15__SCAN_IN), .ZN(n7594) );
  INV_X1 U9810 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15294) );
  XNOR2_X1 U9811 ( .A(P1_ADDR_REG_14__SCAN_IN), .B(P3_ADDR_REG_14__SCAN_IN), 
        .ZN(n7647) );
  INV_X1 U9812 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7579) );
  INV_X1 U9813 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15285) );
  INV_X1 U9814 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14865) );
  XOR2_X1 U9815 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n7600) );
  INV_X1 U9816 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9467) );
  INV_X1 U9817 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15304) );
  INV_X1 U9818 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n7572) );
  INV_X1 U9819 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7557) );
  NOR2_X1 U9820 ( .A1(n7559), .A2(n15082), .ZN(n7561) );
  INV_X1 U9821 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7562) );
  NOR2_X1 U9822 ( .A1(n7563), .A2(n7562), .ZN(n7565) );
  INV_X1 U9823 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9568) );
  INV_X1 U9824 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n13927) );
  NOR2_X1 U9825 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n13927), .ZN(n7567) );
  INV_X1 U9826 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n7566) );
  NOR2_X1 U9827 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n7568), .ZN(n7570) );
  XNOR2_X1 U9828 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n7568), .ZN(n7632) );
  INV_X1 U9829 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7631) );
  INV_X1 U9830 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9449) );
  XOR2_X1 U9831 ( .A(n7572), .B(n9449), .Z(n7637) );
  XNOR2_X1 U9832 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7605) );
  NAND2_X1 U9833 ( .A1(n7604), .A2(n7605), .ZN(n7573) );
  NAND2_X1 U9834 ( .A1(n9467), .A2(n7574), .ZN(n7601) );
  NAND2_X1 U9835 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n7602), .ZN(n7575) );
  XOR2_X1 U9836 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n7597) );
  INV_X1 U9837 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14884) );
  NAND2_X1 U9838 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14884), .ZN(n7578) );
  NAND2_X1 U9839 ( .A1(n7647), .A2(n7646), .ZN(n7580) );
  NOR2_X1 U9840 ( .A1(n7594), .A2(n7593), .ZN(n7581) );
  AOI21_X1 U9841 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n15085), .A(n7581), .ZN(
        n7582) );
  NOR2_X1 U9842 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n7582), .ZN(n7584) );
  INV_X1 U9843 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15271) );
  XNOR2_X1 U9844 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n7582), .ZN(n7592) );
  NOR2_X1 U9845 ( .A1(n15271), .A2(n7592), .ZN(n7583) );
  NOR2_X1 U9846 ( .A1(n7584), .A2(n7583), .ZN(n7585) );
  NOR2_X1 U9847 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n7585), .ZN(n7588) );
  INV_X1 U9848 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n7586) );
  XNOR2_X1 U9849 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n7585), .ZN(n7591) );
  NOR2_X1 U9850 ( .A1(n7586), .A2(n7591), .ZN(n7587) );
  NOR2_X1 U9851 ( .A1(n7588), .A2(n7587), .ZN(n7655) );
  INV_X1 U9852 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12321) );
  NOR2_X1 U9853 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n12321), .ZN(n7589) );
  AOI21_X1 U9854 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n12321), .A(n7589), .ZN(
        n7590) );
  XNOR2_X1 U9855 ( .A(n7655), .B(n7590), .ZN(n14311) );
  XNOR2_X1 U9856 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n7591), .ZN(n7650) );
  XNOR2_X1 U9857 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n7592), .ZN(n14538) );
  XOR2_X1 U9858 ( .A(n7594), .B(n7593), .Z(n14534) );
  XOR2_X1 U9859 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n7595) );
  XOR2_X1 U9860 ( .A(n7596), .B(n7595), .Z(n7644) );
  XOR2_X1 U9861 ( .A(n7598), .B(n7597), .Z(n7643) );
  XNOR2_X1 U9862 ( .A(n7600), .B(n7599), .ZN(n14518) );
  NAND2_X1 U9863 ( .A1(n7602), .A2(n7601), .ZN(n7603) );
  XNOR2_X1 U9864 ( .A(n7603), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14327) );
  XOR2_X1 U9865 ( .A(n7605), .B(n7604), .Z(n14323) );
  INV_X1 U9866 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7606) );
  INV_X1 U9867 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7609) );
  XOR2_X1 U9868 ( .A(n7610), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n7620) );
  XOR2_X1 U9869 ( .A(n7612), .B(n7611), .Z(n14315) );
  INV_X1 U9870 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7617) );
  NOR2_X1 U9871 ( .A1(n7616), .A2(n7617), .ZN(n7618) );
  AOI21_X1 U9872 ( .B1(n9679), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n7614), .ZN(
        n7615) );
  INV_X1 U9873 ( .A(n7615), .ZN(n15332) );
  NAND2_X1 U9874 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15332), .ZN(n15343) );
  NOR2_X1 U9875 ( .A1(n14315), .A2(n14314), .ZN(n7619) );
  NAND2_X1 U9876 ( .A1(n14315), .A2(n14314), .ZN(n14313) );
  OAI21_X1 U9877 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n7619), .A(n14313), .ZN(
        n7621) );
  NAND2_X1 U9878 ( .A1(n7620), .A2(n7621), .ZN(n15338) );
  INV_X1 U9879 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15340) );
  NAND2_X1 U9880 ( .A1(n7623), .A2(n7624), .ZN(n7625) );
  INV_X1 U9881 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15327) );
  INV_X1 U9882 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7626) );
  NOR2_X1 U9883 ( .A1(n7627), .A2(n7626), .ZN(n7630) );
  XNOR2_X1 U9884 ( .A(n7627), .B(n7626), .ZN(n14319) );
  XNOR2_X1 U9885 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n7629) );
  XNOR2_X1 U9886 ( .A(n7629), .B(n7628), .ZN(n14318) );
  INV_X1 U9887 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7634) );
  NOR2_X1 U9888 ( .A1(n7633), .A2(n7634), .ZN(n7635) );
  XNOR2_X1 U9889 ( .A(n7632), .B(n7631), .ZN(n15335) );
  XNOR2_X1 U9890 ( .A(n7637), .B(n7636), .ZN(n7639) );
  NAND2_X1 U9891 ( .A1(n7638), .A2(n7639), .ZN(n7640) );
  INV_X1 U9892 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15086) );
  NAND2_X1 U9893 ( .A1(n14323), .A2(n14324), .ZN(n14322) );
  INV_X1 U9894 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14745) );
  INV_X1 U9895 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14527) );
  XOR2_X1 U9896 ( .A(n7647), .B(n7646), .Z(n7648) );
  INV_X1 U9897 ( .A(n14529), .ZN(n14530) );
  INV_X1 U9898 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14532) );
  NAND2_X1 U9899 ( .A1(n14534), .A2(n14535), .ZN(n14533) );
  NAND2_X1 U9900 ( .A1(n7650), .A2(n7651), .ZN(n7652) );
  INV_X1 U9901 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15226) );
  NAND2_X1 U9902 ( .A1(n14311), .A2(n14310), .ZN(n7653) );
  INV_X1 U9903 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14576) );
  NOR2_X1 U9904 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n14576), .ZN(n7654) );
  OAI22_X1 U9905 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n12321), .B1(n7655), .B2(
        n7654), .ZN(n7658) );
  INV_X2 U9906 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7703) );
  XNOR2_X1 U9907 ( .A(n7703), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7656) );
  XNOR2_X1 U9908 ( .A(n7656), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7657) );
  XNOR2_X1 U9909 ( .A(n7658), .B(n7657), .ZN(n7659) );
  AND2_X1 U9910 ( .A1(n7662), .A2(n7661), .ZN(n7665) );
  NOR3_X2 U9911 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n7664) );
  NOR2_X1 U9912 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7663) );
  INV_X1 U9913 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7672) );
  NAND2_X1 U9914 ( .A1(n7674), .A2(n7675), .ZN(n14291) );
  NAND2_X4 U9916 ( .A1(n11569), .A2(n7680), .ZN(n8324) );
  INV_X1 U9917 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9395) );
  INV_X1 U9918 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7679) );
  OR2_X1 U9919 ( .A1(n7865), .A2(n7679), .ZN(n7683) );
  INV_X1 U9920 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10410) );
  OR2_X1 U9921 ( .A1(n7771), .A2(n10410), .ZN(n7682) );
  NAND2_X1 U9922 ( .A1(n7687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7686) );
  INV_X1 U9923 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7691) );
  INV_X1 U9924 ( .A(n8348), .ZN(n8349) );
  XNOR2_X2 U9925 ( .A(n7695), .B(n7672), .ZN(n13873) );
  NAND2_X1 U9926 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7698) );
  MUX2_X1 U9927 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7698), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n7701) );
  INV_X1 U9928 ( .A(n7699), .ZN(n7700) );
  NAND2_X1 U9929 ( .A1(n7701), .A2(n7700), .ZN(n13867) );
  NAND3_X1 U9930 ( .A1(n7703), .A2(n7702), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7704) );
  NAND2_X1 U9931 ( .A1(n7704), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7709) );
  INV_X1 U9932 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7705) );
  NAND3_X1 U9933 ( .A1(n7706), .A2(n7705), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7707) );
  NAND2_X1 U9934 ( .A1(n7707), .A2(n11299), .ZN(n7708) );
  NAND2_X1 U9935 ( .A1(n7711), .A2(SI_1_), .ZN(n7741) );
  INV_X1 U9936 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8531) );
  INV_X1 U9937 ( .A(SI_0_), .ZN(n9119) );
  NOR2_X1 U9938 ( .A1(n7712), .A2(n9119), .ZN(n7714) );
  INV_X1 U9939 ( .A(n7714), .ZN(n7715) );
  NAND2_X1 U9940 ( .A1(n7742), .A2(n7716), .ZN(n9344) );
  OR2_X1 U9941 ( .A1(n8005), .A2(n7710), .ZN(n7717) );
  AOI21_X1 U9942 ( .B1(n13859), .B2(n7858), .A(n10415), .ZN(n7729) );
  NAND2_X1 U9943 ( .A1(n8320), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7721) );
  INV_X1 U9944 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9594) );
  INV_X1 U9945 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10309) );
  OR2_X1 U9946 ( .A1(n7771), .A2(n10309), .ZN(n7720) );
  INV_X1 U9947 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7718) );
  OR2_X1 U9948 ( .A1(n8269), .A2(n7718), .ZN(n7719) );
  NOR2_X1 U9949 ( .A1(n9343), .A2(n9119), .ZN(n7722) );
  XNOR2_X1 U9950 ( .A(n7722), .B(n8531), .ZN(n14308) );
  NAND2_X1 U9951 ( .A1(n10404), .A2(n10400), .ZN(n8358) );
  INV_X1 U9952 ( .A(n8358), .ZN(n7723) );
  NAND3_X1 U9953 ( .A1(n7723), .A2(n8376), .A3(n10018), .ZN(n7728) );
  NAND2_X1 U9954 ( .A1(n13860), .A2(n10312), .ZN(n8357) );
  OAI211_X1 U9955 ( .C1(n7730), .C2(n7729), .A(n7728), .B(n7727), .ZN(n7751)
         );
  INV_X1 U9956 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7731) );
  OR2_X1 U9957 ( .A1(n7771), .A2(n7731), .ZN(n7736) );
  NAND2_X1 U9958 ( .A1(n7971), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7735) );
  INV_X1 U9959 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7732) );
  OR2_X1 U9960 ( .A1(n7865), .A2(n7732), .ZN(n7734) );
  INV_X1 U9961 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9394) );
  OR2_X1 U9962 ( .A1(n8269), .A2(n9394), .ZN(n7733) );
  NOR2_X1 U9963 ( .A1(n7699), .A2(n7691), .ZN(n7737) );
  MUX2_X1 U9964 ( .A(n7691), .B(n7737), .S(P1_IR_REG_2__SCAN_IN), .Z(n7738) );
  INV_X1 U9965 ( .A(n7738), .ZN(n7740) );
  NAND2_X1 U9966 ( .A1(n7740), .A2(n7739), .ZN(n13884) );
  INV_X1 U9967 ( .A(n7746), .ZN(n7744) );
  NAND2_X1 U9968 ( .A1(n7743), .A2(SI_2_), .ZN(n7756) );
  OAI21_X1 U9969 ( .B1(n7743), .B2(SI_2_), .A(n7756), .ZN(n7745) );
  NAND2_X1 U9970 ( .A1(n7744), .A2(n7745), .ZN(n7748) );
  INV_X1 U9971 ( .A(n7745), .ZN(n7747) );
  NAND2_X1 U9972 ( .A1(n7748), .A2(n7757), .ZN(n9527) );
  OR2_X1 U9973 ( .A1(n9527), .A2(n8002), .ZN(n7750) );
  INV_X1 U9974 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9113) );
  OR2_X1 U9975 ( .A1(n8005), .A2(n9113), .ZN(n7749) );
  NAND2_X1 U9976 ( .A1(n13858), .A2(n14585), .ZN(n7763) );
  NAND2_X1 U9977 ( .A1(n8320), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7755) );
  OR2_X1 U9978 ( .A1(n7771), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7754) );
  INV_X1 U9979 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9415) );
  OR2_X1 U9980 ( .A1(n8324), .A2(n9415), .ZN(n7753) );
  INV_X1 U9981 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10384) );
  OR2_X1 U9982 ( .A1(n8269), .A2(n10384), .ZN(n7752) );
  NAND2_X1 U9983 ( .A1(n7757), .A2(n7756), .ZN(n7778) );
  NAND2_X1 U9984 ( .A1(n7758), .A2(SI_3_), .ZN(n7779) );
  OAI21_X1 U9985 ( .B1(n7758), .B2(SI_3_), .A(n7779), .ZN(n7776) );
  XNOR2_X1 U9986 ( .A(n7778), .B(n7776), .ZN(n9640) );
  NAND2_X1 U9987 ( .A1(n9640), .A2(n6539), .ZN(n7762) );
  INV_X2 U9988 ( .A(n7759), .ZN(n9314) );
  NAND2_X1 U9989 ( .A1(n7739), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7760) );
  XNOR2_X1 U9990 ( .A(n7760), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U9991 ( .A1(n6526), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n9314), .B2(
        n13896), .ZN(n7761) );
  XNOR2_X1 U9992 ( .A(n13857), .B(n10388), .ZN(n10379) );
  CLKBUF_X3 U9993 ( .A(n7858), .Z(n7989) );
  NAND2_X1 U9994 ( .A1(n13857), .A2(n8376), .ZN(n7768) );
  NAND2_X1 U9995 ( .A1(n10365), .A2(n7858), .ZN(n7767) );
  MUX2_X1 U9996 ( .A(n7768), .B(n7767), .S(n10388), .Z(n7769) );
  NAND2_X1 U9997 ( .A1(n8320), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7775) );
  INV_X1 U9998 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9418) );
  OR2_X1 U9999 ( .A1(n8324), .A2(n9418), .ZN(n7774) );
  INV_X1 U10000 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10392) );
  OR2_X1 U10001 ( .A1(n8269), .A2(n10392), .ZN(n7773) );
  XNOR2_X1 U10002 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10395) );
  OR2_X1 U10003 ( .A1(n8298), .A2(n10395), .ZN(n7772) );
  INV_X1 U10004 ( .A(n7776), .ZN(n7777) );
  NAND2_X1 U10005 ( .A1(n7778), .A2(n7777), .ZN(n7780) );
  NAND2_X1 U10006 ( .A1(n7781), .A2(SI_4_), .ZN(n7794) );
  OAI21_X1 U10007 ( .B1(n7781), .B2(SI_4_), .A(n7794), .ZN(n7791) );
  XNOR2_X1 U10008 ( .A(n7793), .B(n7791), .ZN(n9741) );
  NAND2_X1 U10009 ( .A1(n9741), .A2(n8347), .ZN(n7788) );
  NAND2_X1 U10010 ( .A1(n7782), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7783) );
  MUX2_X1 U10011 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7783), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n7786) );
  INV_X1 U10012 ( .A(n7782), .ZN(n7785) );
  INV_X1 U10013 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U10014 ( .A1(n7785), .A2(n7784), .ZN(n7799) );
  NAND2_X1 U10015 ( .A1(n7786), .A2(n7799), .ZN(n13914) );
  INV_X1 U10016 ( .A(n13914), .ZN(n9421) );
  AOI22_X1 U10017 ( .A1(n8346), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9314), .B2(
        n9421), .ZN(n7787) );
  MUX2_X1 U10018 ( .A(n10585), .B(n10453), .S(n8376), .Z(n7790) );
  MUX2_X1 U10019 ( .A(n13855), .B(n10456), .S(n7989), .Z(n7789) );
  INV_X1 U10020 ( .A(n7791), .ZN(n7792) );
  NAND2_X1 U10021 ( .A1(n7793), .A2(n7792), .ZN(n7795) );
  NAND2_X1 U10022 ( .A1(n7797), .A2(n7826), .ZN(n9845) );
  NAND2_X1 U10023 ( .A1(n7799), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7798) );
  MUX2_X1 U10024 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7798), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7802) );
  INV_X1 U10025 ( .A(n7799), .ZN(n7801) );
  INV_X1 U10026 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U10027 ( .A1(n7801), .A2(n7800), .ZN(n7854) );
  AND2_X1 U10028 ( .A1(n7802), .A2(n7854), .ZN(n9566) );
  AOI22_X1 U10029 ( .A1(n8346), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9314), .B2(
        n9566), .ZN(n7803) );
  AOI21_X1 U10030 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7805) );
  NOR2_X1 U10031 ( .A1(n7805), .A2(n7819), .ZN(n10578) );
  NAND2_X1 U10032 ( .A1(n8180), .A2(n10578), .ZN(n7811) );
  INV_X1 U10033 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9398) );
  OR2_X1 U10034 ( .A1(n8269), .A2(n9398), .ZN(n7810) );
  INV_X1 U10035 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7806) );
  OR2_X1 U10036 ( .A1(n8324), .A2(n7806), .ZN(n7809) );
  INV_X1 U10037 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7807) );
  OR2_X1 U10038 ( .A1(n8277), .A2(n7807), .ZN(n7808) );
  MUX2_X1 U10039 ( .A(n10579), .B(n13854), .S(n8376), .Z(n7815) );
  MUX2_X1 U10040 ( .A(n10579), .B(n13854), .S(n7858), .Z(n7812) );
  NAND2_X1 U10041 ( .A1(n7813), .A2(n7812), .ZN(n7836) );
  INV_X1 U10042 ( .A(n7814), .ZN(n7817) );
  INV_X1 U10043 ( .A(n7815), .ZN(n7816) );
  NAND2_X1 U10044 ( .A1(n7817), .A2(n7816), .ZN(n7838) );
  NAND2_X1 U10045 ( .A1(n8319), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7824) );
  INV_X1 U10046 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7818) );
  OR2_X1 U10047 ( .A1(n8324), .A2(n7818), .ZN(n7823) );
  NAND2_X1 U10048 ( .A1(n7819), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7840) );
  OAI21_X1 U10049 ( .B1(n7819), .B2(P1_REG3_REG_6__SCAN_IN), .A(n7840), .ZN(
        n10615) );
  OR2_X1 U10050 ( .A1(n8298), .A2(n10615), .ZN(n7822) );
  INV_X1 U10051 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7820) );
  OR2_X1 U10052 ( .A1(n8277), .A2(n7820), .ZN(n7821) );
  NAND4_X1 U10053 ( .A1(n7824), .A2(n7823), .A3(n7822), .A4(n7821), .ZN(n13853) );
  NAND2_X1 U10054 ( .A1(n7827), .A2(SI_6_), .ZN(n7847) );
  OAI21_X1 U10055 ( .B1(SI_6_), .B2(n7827), .A(n7847), .ZN(n7828) );
  INV_X1 U10056 ( .A(n7828), .ZN(n7829) );
  OR2_X1 U10057 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  NAND2_X1 U10058 ( .A1(n7848), .A2(n7831), .ZN(n9967) );
  OR2_X1 U10059 ( .A1(n9967), .A2(n6531), .ZN(n7834) );
  NAND2_X1 U10060 ( .A1(n7854), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7832) );
  XNOR2_X1 U10061 ( .A(n7832), .B(P1_IR_REG_6__SCAN_IN), .ZN(n13929) );
  AOI22_X1 U10062 ( .A1(n8346), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9314), .B2(
        n13929), .ZN(n7833) );
  MUX2_X1 U10063 ( .A(n13853), .B(n10612), .S(n8376), .Z(n7837) );
  MUX2_X1 U10064 ( .A(n10612), .B(n13853), .S(n8376), .Z(n7835) );
  NAND2_X1 U10065 ( .A1(n8319), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7846) );
  INV_X1 U10066 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9426) );
  OR2_X1 U10067 ( .A1(n8324), .A2(n9426), .ZN(n7845) );
  AND2_X1 U10068 ( .A1(n7840), .A2(n7839), .ZN(n7841) );
  OR2_X1 U10069 ( .A1(n7841), .A2(n7863), .ZN(n10683) );
  OR2_X1 U10070 ( .A1(n8298), .A2(n10683), .ZN(n7844) );
  INV_X1 U10071 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7842) );
  OR2_X1 U10072 ( .A1(n8277), .A2(n7842), .ZN(n7843) );
  NAND4_X1 U10073 ( .A1(n7846), .A2(n7845), .A3(n7844), .A4(n7843), .ZN(n13852) );
  NAND2_X1 U10074 ( .A1(n7849), .A2(SI_7_), .ZN(n7871) );
  OAI21_X1 U10075 ( .B1(n7849), .B2(SI_7_), .A(n7871), .ZN(n7850) );
  INV_X1 U10076 ( .A(n7850), .ZN(n7851) );
  OR2_X1 U10077 ( .A1(n7852), .A2(n7851), .ZN(n7853) );
  NAND2_X1 U10078 ( .A1(n7872), .A2(n7853), .ZN(n10060) );
  OR2_X1 U10079 ( .A1(n10060), .A2(n6531), .ZN(n7857) );
  NAND2_X1 U10080 ( .A1(n7878), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7855) );
  XNOR2_X1 U10081 ( .A(n7855), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9546) );
  AOI22_X1 U10082 ( .A1(n8346), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9314), .B2(
        n9546), .ZN(n7856) );
  MUX2_X1 U10083 ( .A(n13852), .B(n10689), .S(n7858), .Z(n7861) );
  MUX2_X1 U10084 ( .A(n10689), .B(n13852), .S(n7989), .Z(n7859) );
  INV_X1 U10085 ( .A(n7861), .ZN(n7862) );
  NAND2_X1 U10086 ( .A1(n8319), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7870) );
  INV_X1 U10087 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9428) );
  OR2_X1 U10088 ( .A1(n8324), .A2(n9428), .ZN(n7869) );
  NAND2_X1 U10089 ( .A1(n7863), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7887) );
  OR2_X1 U10090 ( .A1(n7863), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U10091 ( .A1(n7887), .A2(n7864), .ZN(n11028) );
  OR2_X1 U10092 ( .A1(n8298), .A2(n11028), .ZN(n7868) );
  INV_X1 U10093 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7866) );
  OR2_X1 U10094 ( .A1(n8277), .A2(n7866), .ZN(n7867) );
  NAND4_X1 U10095 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .ZN(n13851) );
  NAND2_X1 U10096 ( .A1(n7873), .A2(SI_8_), .ZN(n7893) );
  OAI21_X1 U10097 ( .B1(SI_8_), .B2(n7873), .A(n7893), .ZN(n7874) );
  OR2_X1 U10098 ( .A1(n7876), .A2(n7875), .ZN(n7877) );
  NAND2_X1 U10099 ( .A1(n7900), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7879) );
  XNOR2_X1 U10100 ( .A(n7879), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9451) );
  AOI22_X1 U10101 ( .A1(n8346), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9314), .B2(
        n9451), .ZN(n7880) );
  MUX2_X1 U10102 ( .A(n13851), .B(n11030), .S(n8376), .Z(n7882) );
  MUX2_X1 U10103 ( .A(n13851), .B(n11030), .S(n7989), .Z(n7881) );
  INV_X1 U10104 ( .A(n7882), .ZN(n7883) );
  NAND2_X1 U10105 ( .A1(n8320), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7892) );
  INV_X1 U10106 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7885) );
  OR2_X1 U10107 ( .A1(n8324), .A2(n7885), .ZN(n7891) );
  INV_X1 U10108 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10631) );
  OR2_X1 U10109 ( .A1(n8269), .A2(n10631), .ZN(n7890) );
  NAND2_X1 U10110 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  NAND2_X1 U10111 ( .A1(n7907), .A2(n7888), .ZN(n11165) );
  OR2_X1 U10112 ( .A1(n8298), .A2(n11165), .ZN(n7889) );
  NAND4_X1 U10113 ( .A1(n7892), .A2(n7891), .A3(n7890), .A4(n7889), .ZN(n13850) );
  NAND2_X1 U10114 ( .A1(n7895), .A2(SI_9_), .ZN(n7914) );
  OAI21_X1 U10115 ( .B1(n7895), .B2(SI_9_), .A(n7914), .ZN(n7896) );
  INV_X1 U10116 ( .A(n7896), .ZN(n7897) );
  OR2_X1 U10117 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  NAND2_X1 U10118 ( .A1(n7915), .A2(n7899), .ZN(n10494) );
  OR2_X1 U10119 ( .A1(n10494), .A2(n6531), .ZN(n7902) );
  XNOR2_X1 U10120 ( .A(n7940), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9488) );
  AOI22_X1 U10121 ( .A1(n8346), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9314), .B2(
        n9488), .ZN(n7901) );
  MUX2_X1 U10122 ( .A(n13850), .B(n14616), .S(n7989), .Z(n7904) );
  MUX2_X1 U10123 ( .A(n13850), .B(n14616), .S(n8376), .Z(n7903) );
  INV_X1 U10124 ( .A(n7904), .ZN(n7905) );
  NAND2_X1 U10125 ( .A1(n8319), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7913) );
  INV_X1 U10126 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9432) );
  OR2_X1 U10127 ( .A1(n8324), .A2(n9432), .ZN(n7912) );
  NAND2_X1 U10128 ( .A1(n7907), .A2(n7906), .ZN(n7908) );
  NAND2_X1 U10129 ( .A1(n7931), .A2(n7908), .ZN(n11348) );
  OR2_X1 U10130 ( .A1(n8298), .A2(n11348), .ZN(n7911) );
  INV_X1 U10131 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7909) );
  OR2_X1 U10132 ( .A1(n8277), .A2(n7909), .ZN(n7910) );
  NAND4_X1 U10133 ( .A1(n7913), .A2(n7912), .A3(n7911), .A4(n7910), .ZN(n13849) );
  OAI21_X1 U10134 ( .B1(n7916), .B2(SI_10_), .A(n7936), .ZN(n7917) );
  INV_X1 U10135 ( .A(n7917), .ZN(n7918) );
  OR2_X1 U10136 ( .A1(n7919), .A2(n7918), .ZN(n7920) );
  NAND2_X1 U10137 ( .A1(n7937), .A2(n7920), .ZN(n10734) );
  OR2_X1 U10138 ( .A1(n10734), .A2(n6531), .ZN(n7925) );
  INV_X1 U10139 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10140 ( .A1(n7940), .A2(n7921), .ZN(n7922) );
  NAND2_X1 U10141 ( .A1(n7922), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7923) );
  XNOR2_X1 U10142 ( .A(n7923), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9469) );
  AOI22_X1 U10143 ( .A1(n9314), .A2(n9469), .B1(n8346), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n7924) );
  MUX2_X1 U10144 ( .A(n13849), .B(n11345), .S(n8376), .Z(n7927) );
  MUX2_X1 U10145 ( .A(n13849), .B(n11345), .S(n7989), .Z(n7926) );
  INV_X1 U10146 ( .A(n7927), .ZN(n7928) );
  NAND2_X1 U10147 ( .A1(n8320), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7935) );
  INV_X1 U10148 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7929) );
  OR2_X1 U10149 ( .A1(n8324), .A2(n7929), .ZN(n7934) );
  OR2_X1 U10150 ( .A1(n7550), .A2(n7948), .ZN(n14484) );
  OR2_X1 U10151 ( .A1(n8298), .A2(n14484), .ZN(n7933) );
  INV_X1 U10152 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10957) );
  OR2_X1 U10153 ( .A1(n8269), .A2(n10957), .ZN(n7932) );
  NAND4_X1 U10154 ( .A1(n7935), .A2(n7934), .A3(n7933), .A4(n7932), .ZN(n13848) );
  XNOR2_X1 U10155 ( .A(n7958), .B(n7957), .ZN(n10747) );
  NAND2_X1 U10156 ( .A1(n10747), .A2(n8347), .ZN(n7943) );
  OR2_X1 U10157 ( .A1(n7938), .A2(n7691), .ZN(n7939) );
  NAND2_X1 U10158 ( .A1(n7940), .A2(n7939), .ZN(n7959) );
  INV_X1 U10159 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n7941) );
  XNOR2_X1 U10160 ( .A(n7959), .B(n7941), .ZN(n13950) );
  AOI22_X1 U10161 ( .A1(n8346), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n13950), 
        .B2(n9314), .ZN(n7942) );
  MUX2_X1 U10162 ( .A(n13848), .B(n14504), .S(n7989), .Z(n7945) );
  MUX2_X1 U10163 ( .A(n13848), .B(n14504), .S(n8376), .Z(n7944) );
  INV_X1 U10164 ( .A(n7945), .ZN(n7946) );
  NAND2_X1 U10165 ( .A1(n8320), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7953) );
  INV_X1 U10166 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11112) );
  OR2_X1 U10167 ( .A1(n8269), .A2(n11112), .ZN(n7952) );
  INV_X1 U10168 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7947) );
  OR2_X1 U10169 ( .A1(n8324), .A2(n7947), .ZN(n7951) );
  OR2_X1 U10170 ( .A1(n7948), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10171 ( .A1(n8012), .A2(n7949), .ZN(n13764) );
  OR2_X1 U10172 ( .A1(n8298), .A2(n13764), .ZN(n7950) );
  NAND4_X1 U10173 ( .A1(n7953), .A2(n7952), .A3(n7951), .A4(n7950), .ZN(n13847) );
  INV_X1 U10174 ( .A(n7954), .ZN(n7955) );
  NAND2_X1 U10175 ( .A1(n7955), .A2(n9161), .ZN(n7956) );
  XNOR2_X1 U10176 ( .A(n7978), .B(n7977), .ZN(n10885) );
  NAND2_X1 U10177 ( .A1(n10885), .A2(n8347), .ZN(n7962) );
  NAND2_X1 U10178 ( .A1(n7960), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7982) );
  XNOR2_X1 U10179 ( .A(n7982), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9434) );
  AOI22_X1 U10180 ( .A1(n9434), .A2(n9314), .B1(n8346), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n7961) );
  MUX2_X1 U10181 ( .A(n13847), .B(n13601), .S(n8376), .Z(n7966) );
  MUX2_X1 U10182 ( .A(n13847), .B(n13601), .S(n7989), .Z(n7963) );
  NAND2_X1 U10183 ( .A1(n7964), .A2(n7963), .ZN(n7970) );
  INV_X1 U10184 ( .A(n7965), .ZN(n7968) );
  INV_X1 U10185 ( .A(n7966), .ZN(n7967) );
  NAND2_X1 U10186 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  NAND2_X1 U10187 ( .A1(n8268), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7976) );
  INV_X1 U10188 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8010) );
  XNOR2_X1 U10189 ( .A(n8012), .B(n8010), .ZN(n13797) );
  OR2_X1 U10190 ( .A1(n8298), .A2(n13797), .ZN(n7975) );
  INV_X1 U10191 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7972) );
  OR2_X1 U10192 ( .A1(n8277), .A2(n7972), .ZN(n7974) );
  INV_X1 U10193 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11202) );
  OR2_X1 U10194 ( .A1(n8269), .A2(n11202), .ZN(n7973) );
  NAND4_X1 U10195 ( .A1(n7976), .A2(n7975), .A3(n7974), .A4(n7973), .ZN(n13846) );
  INV_X1 U10196 ( .A(n7979), .ZN(n7980) );
  XNOR2_X1 U10197 ( .A(n7994), .B(n7993), .ZN(n11207) );
  NAND2_X1 U10198 ( .A1(n11207), .A2(n8347), .ZN(n7988) );
  INV_X1 U10199 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7981) );
  AOI21_X1 U10200 ( .B1(n7982), .B2(n7981), .A(n7691), .ZN(n7983) );
  NAND2_X1 U10201 ( .A1(n7983), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n7986) );
  INV_X1 U10202 ( .A(n7983), .ZN(n7985) );
  INV_X1 U10203 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U10204 ( .A1(n7985), .A2(n7984), .ZN(n8003) );
  AOI22_X1 U10205 ( .A1(n9760), .A2(n9314), .B1(n8346), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n7987) );
  MUX2_X1 U10206 ( .A(n13846), .B(n13610), .S(n7989), .Z(n7991) );
  MUX2_X1 U10207 ( .A(n13846), .B(n13610), .S(n8376), .Z(n7990) );
  INV_X1 U10208 ( .A(n7991), .ZN(n7992) );
  INV_X1 U10209 ( .A(SI_13_), .ZN(n7995) );
  NAND2_X1 U10210 ( .A1(n7996), .A2(n7995), .ZN(n7997) );
  INV_X1 U10211 ( .A(SI_14_), .ZN(n9312) );
  NAND2_X1 U10212 ( .A1(n8056), .A2(n9312), .ZN(n7999) );
  NAND2_X1 U10213 ( .A1(n8000), .A2(n8050), .ZN(n8001) );
  NAND2_X1 U10214 ( .A1(n8020), .A2(n8001), .ZN(n11376) );
  OR2_X1 U10215 ( .A1(n11376), .A2(n8002), .ZN(n8008) );
  NAND2_X1 U10216 ( .A1(n8003), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8004) );
  XNOR2_X1 U10217 ( .A(n8004), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10823) );
  NOR2_X1 U10218 ( .A1(n8005), .A2(n15126), .ZN(n8006) );
  AOI21_X1 U10219 ( .B1(n10823), .B2(n9314), .A(n8006), .ZN(n8007) );
  NAND2_X1 U10220 ( .A1(n8320), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8018) );
  INV_X1 U10221 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8009) );
  OAI21_X1 U10222 ( .B1(n8012), .B2(n8010), .A(n8009), .ZN(n8013) );
  NAND2_X1 U10223 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n8011) );
  NAND2_X1 U10224 ( .A1(n8013), .A2(n8029), .ZN(n14439) );
  OR2_X1 U10225 ( .A1(n8298), .A2(n14439), .ZN(n8017) );
  INV_X1 U10226 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8014) );
  OR2_X1 U10227 ( .A1(n8324), .A2(n8014), .ZN(n8016) );
  INV_X1 U10228 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11303) );
  OR2_X1 U10229 ( .A1(n8269), .A2(n11303), .ZN(n8015) );
  NAND2_X1 U10230 ( .A1(n14436), .A2(n13833), .ZN(n8038) );
  NAND2_X1 U10231 ( .A1(n8020), .A2(n8019), .ZN(n8021) );
  XNOR2_X1 U10232 ( .A(n8057), .B(SI_15_), .ZN(n8051) );
  NAND2_X1 U10233 ( .A1(n11383), .A2(n8347), .ZN(n8028) );
  NOR2_X1 U10234 ( .A1(n8025), .A2(n7691), .ZN(n8023) );
  MUX2_X1 U10235 ( .A(n7691), .B(n8023), .S(P1_IR_REG_15__SCAN_IN), .Z(n8026)
         );
  INV_X1 U10236 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8024) );
  AND2_X1 U10237 ( .A1(n8025), .A2(n8024), .ZN(n8061) );
  OR2_X1 U10238 ( .A1(n8026), .A2(n8061), .ZN(n14554) );
  AOI22_X1 U10239 ( .A1(n8346), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9314), 
        .B2(n10827), .ZN(n8027) );
  AND2_X1 U10240 ( .A1(n8029), .A2(n15138), .ZN(n8030) );
  NOR2_X1 U10241 ( .A1(n8044), .A2(n8030), .ZN(n13836) );
  NAND2_X1 U10242 ( .A1(n8180), .A2(n13836), .ZN(n8037) );
  INV_X1 U10243 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8031) );
  OR2_X1 U10244 ( .A1(n8269), .A2(n8031), .ZN(n8036) );
  INV_X1 U10245 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8032) );
  OR2_X1 U10246 ( .A1(n8324), .A2(n8032), .ZN(n8035) );
  INV_X1 U10247 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8033) );
  OR2_X1 U10248 ( .A1(n8277), .A2(n8033), .ZN(n8034) );
  NAND2_X1 U10249 ( .A1(n13622), .A2(n14441), .ZN(n8355) );
  AND2_X1 U10250 ( .A1(n8355), .A2(n8038), .ZN(n8040) );
  MUX2_X1 U10251 ( .A(n8040), .B(n8039), .S(n7989), .Z(n8041) );
  MUX2_X1 U10252 ( .A(n8355), .B(n11455), .S(n8376), .Z(n8042) );
  NAND2_X1 U10253 ( .A1(n8043), .A2(n8042), .ZN(n8083) );
  NOR2_X1 U10254 ( .A1(n8044), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8045) );
  OR2_X1 U10255 ( .A1(n8067), .A2(n8045), .ZN(n14453) );
  NAND2_X1 U10256 ( .A1(n8268), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8046) );
  OAI21_X1 U10257 ( .B1(n14453), .B2(n8298), .A(n8046), .ZN(n8049) );
  INV_X1 U10258 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n13964) );
  NAND2_X1 U10259 ( .A1(n8320), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8047) );
  OAI21_X1 U10260 ( .B1(n8269), .B2(n13964), .A(n8047), .ZN(n8048) );
  INV_X1 U10261 ( .A(n14458), .ZN(n13629) );
  NAND2_X1 U10262 ( .A1(n8052), .A2(SI_14_), .ZN(n8053) );
  INV_X1 U10263 ( .A(n8057), .ZN(n8058) );
  XNOR2_X1 U10264 ( .A(n8074), .B(n8073), .ZN(n11516) );
  NAND2_X1 U10265 ( .A1(n11516), .A2(n8347), .ZN(n8065) );
  NOR2_X1 U10266 ( .A1(n8061), .A2(n7691), .ZN(n8059) );
  MUX2_X1 U10267 ( .A(n7691), .B(n8059), .S(P1_IR_REG_16__SCAN_IN), .Z(n8063)
         );
  INV_X1 U10268 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U10269 ( .A1(n8061), .A2(n8060), .ZN(n8087) );
  INV_X1 U10270 ( .A(n8087), .ZN(n8062) );
  OR2_X1 U10271 ( .A1(n8063), .A2(n8062), .ZN(n10822) );
  INV_X1 U10272 ( .A(n10822), .ZN(n13966) );
  AOI22_X1 U10273 ( .A1(n8346), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9314), 
        .B2(n13966), .ZN(n8064) );
  MUX2_X1 U10274 ( .A(n13629), .B(n13631), .S(n8376), .Z(n8082) );
  MUX2_X1 U10275 ( .A(n14458), .B(n14450), .S(n7989), .Z(n8066) );
  OAI21_X1 U10276 ( .B1(n8083), .B2(n8082), .A(n8066), .ZN(n8098) );
  OR2_X1 U10277 ( .A1(n8067), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U10278 ( .A1(n8094), .A2(n8068), .ZN(n14468) );
  INV_X1 U10279 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n15123) );
  OR2_X1 U10280 ( .A1(n8277), .A2(n15123), .ZN(n8070) );
  INV_X1 U10281 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11283) );
  OR2_X1 U10282 ( .A1(n8324), .A2(n11283), .ZN(n8069) );
  AND2_X1 U10283 ( .A1(n8070), .A2(n8069), .ZN(n8072) );
  INV_X1 U10284 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11479) );
  OR2_X1 U10285 ( .A1(n8269), .A2(n11479), .ZN(n8071) );
  OAI211_X1 U10286 ( .C1(n14468), .C2(n8298), .A(n8072), .B(n8071), .ZN(n14440) );
  INV_X1 U10287 ( .A(SI_16_), .ZN(n9581) );
  NAND2_X1 U10288 ( .A1(n8075), .A2(n9581), .ZN(n8076) );
  XNOR2_X1 U10289 ( .A(n8084), .B(SI_17_), .ZN(n8078) );
  XNOR2_X1 U10290 ( .A(n8086), .B(n8078), .ZN(n11547) );
  NAND2_X1 U10291 ( .A1(n11547), .A2(n8347), .ZN(n8081) );
  NAND2_X1 U10292 ( .A1(n8087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8079) );
  XNOR2_X1 U10293 ( .A(n8079), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U10294 ( .A1(n8346), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9314), 
        .B2(n11273), .ZN(n8080) );
  MUX2_X1 U10295 ( .A(n14440), .B(n14259), .S(n8376), .Z(n8099) );
  NOR2_X1 U10296 ( .A1(n14259), .A2(n14440), .ZN(n11578) );
  INV_X1 U10297 ( .A(SI_17_), .ZN(n9777) );
  INV_X1 U10298 ( .A(n8084), .ZN(n8085) );
  XNOR2_X1 U10299 ( .A(n8136), .B(SI_18_), .ZN(n8104) );
  XNOR2_X1 U10300 ( .A(n8104), .B(n8129), .ZN(n11848) );
  NAND2_X1 U10301 ( .A1(n11848), .A2(n8347), .ZN(n8092) );
  OAI21_X1 U10302 ( .B1(n8087), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8088) );
  MUX2_X1 U10303 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8088), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n8090) );
  AND2_X1 U10304 ( .A1(n8090), .A2(n8089), .ZN(n11286) );
  AOI22_X1 U10305 ( .A1(n8346), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9314), 
        .B2(n11286), .ZN(n8091) );
  INV_X1 U10306 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U10307 ( .A1(n8094), .A2(n8093), .ZN(n8095) );
  NAND2_X1 U10308 ( .A1(n8114), .A2(n8095), .ZN(n14156) );
  AOI22_X1 U10309 ( .A1(n8268), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8319), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U10310 ( .A1(n8320), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8096) );
  OAI211_X1 U10311 ( .C1(n14156), .C2(n8298), .A(n8097), .B(n8096), .ZN(n14456) );
  XNOR2_X1 U10312 ( .A(n14254), .B(n14456), .ZN(n14149) );
  NAND2_X1 U10313 ( .A1(n14259), .A2(n14440), .ZN(n11577) );
  NAND3_X1 U10314 ( .A1(n14149), .A2(n11577), .A3(n8099), .ZN(n8103) );
  INV_X1 U10315 ( .A(n14456), .ZN(n14135) );
  OR3_X1 U10316 ( .A1(n14254), .A2(n8376), .A3(n14135), .ZN(n8101) );
  NAND3_X1 U10317 ( .A1(n14254), .A2(n14135), .A3(n8376), .ZN(n8100) );
  INV_X1 U10318 ( .A(n8104), .ZN(n8105) );
  NAND2_X1 U10319 ( .A1(n8105), .A2(n8129), .ZN(n8107) );
  NAND2_X1 U10320 ( .A1(n8136), .A2(SI_18_), .ZN(n8106) );
  NAND2_X1 U10321 ( .A1(n8107), .A2(n8106), .ZN(n8111) );
  NAND2_X1 U10322 ( .A1(n8108), .A2(SI_19_), .ZN(n8132) );
  INV_X1 U10323 ( .A(n8108), .ZN(n8109) );
  INV_X1 U10324 ( .A(SI_19_), .ZN(n9930) );
  NAND2_X1 U10325 ( .A1(n8109), .A2(n9930), .ZN(n8130) );
  NAND2_X1 U10326 ( .A1(n8132), .A2(n8130), .ZN(n8110) );
  NAND2_X1 U10327 ( .A1(n11860), .A2(n8347), .ZN(n8113) );
  AOI22_X1 U10328 ( .A1(n8346), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10792), 
        .B2(n9314), .ZN(n8112) );
  INV_X1 U10329 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n15168) );
  AND2_X1 U10330 ( .A1(n8114), .A2(n15168), .ZN(n8115) );
  NOR2_X1 U10331 ( .A1(n8115), .A2(n8148), .ZN(n14141) );
  INV_X1 U10332 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n11289) );
  NAND2_X1 U10333 ( .A1(n8319), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U10334 ( .A1(n8320), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8116) );
  OAI211_X1 U10335 ( .C1(n8324), .C2(n11289), .A(n8117), .B(n8116), .ZN(n8118)
         );
  AOI21_X1 U10336 ( .B1(n14141), .B2(n8180), .A(n8118), .ZN(n13816) );
  NAND2_X1 U10337 ( .A1(n14249), .A2(n13816), .ZN(n11587) );
  OR2_X1 U10338 ( .A1(n14249), .A2(n13816), .ZN(n8119) );
  INV_X1 U10339 ( .A(n13816), .ZN(n14153) );
  NAND2_X1 U10340 ( .A1(n14153), .A2(n7989), .ZN(n8120) );
  OAI22_X1 U10341 ( .A1(n11587), .A2(n7989), .B1(n14249), .B2(n8120), .ZN(
        n8121) );
  INV_X1 U10342 ( .A(n8121), .ZN(n8122) );
  INV_X1 U10343 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13791) );
  XNOR2_X1 U10344 ( .A(n8148), .B(n13791), .ZN(n14122) );
  NAND2_X1 U10345 ( .A1(n14122), .A2(n8180), .ZN(n8127) );
  INV_X1 U10346 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n15122) );
  NAND2_X1 U10347 ( .A1(n8319), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8124) );
  NAND2_X1 U10348 ( .A1(n8320), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8123) );
  OAI211_X1 U10349 ( .C1(n8324), .C2(n15122), .A(n8124), .B(n8123), .ZN(n8125)
         );
  INV_X1 U10350 ( .A(n8125), .ZN(n8126) );
  NAND2_X1 U10351 ( .A1(n8127), .A2(n8126), .ZN(n14103) );
  INV_X1 U10352 ( .A(SI_18_), .ZN(n9928) );
  INV_X1 U10353 ( .A(n8129), .ZN(n8128) );
  OAI21_X1 U10354 ( .B1(n9928), .B2(n8128), .A(n8132), .ZN(n8135) );
  NOR2_X1 U10355 ( .A1(n8129), .A2(SI_18_), .ZN(n8133) );
  INV_X1 U10356 ( .A(n8130), .ZN(n8131) );
  AOI21_X1 U10357 ( .B1(n8133), .B2(n8132), .A(n8131), .ZN(n8134) );
  XNOR2_X1 U10358 ( .A(n8155), .B(n8154), .ZN(n11868) );
  NAND2_X1 U10359 ( .A1(n11868), .A2(n8347), .ZN(n8138) );
  INV_X1 U10360 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10972) );
  OR2_X1 U10361 ( .A1(n8005), .A2(n10972), .ZN(n8137) );
  MUX2_X1 U10362 ( .A(n14103), .B(n14244), .S(n8376), .Z(n8142) );
  MUX2_X1 U10363 ( .A(n14103), .B(n14244), .S(n7989), .Z(n8139) );
  NAND2_X1 U10364 ( .A1(n8140), .A2(n8139), .ZN(n8146) );
  INV_X1 U10365 ( .A(n8141), .ZN(n8144) );
  INV_X1 U10366 ( .A(n8142), .ZN(n8143) );
  NAND2_X1 U10367 ( .A1(n8144), .A2(n8143), .ZN(n8145) );
  AND2_X1 U10368 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n8147) );
  AOI21_X1 U10369 ( .B1(n8148), .B2(P1_REG3_REG_20__SCAN_IN), .A(
        P1_REG3_REG_21__SCAN_IN), .ZN(n8149) );
  OR2_X1 U10370 ( .A1(n8162), .A2(n8149), .ZN(n14107) );
  INV_X1 U10371 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14102) );
  NAND2_X1 U10372 ( .A1(n8268), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10373 ( .A1(n8320), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8150) );
  OAI211_X1 U10374 ( .C1(n8269), .C2(n14102), .A(n8151), .B(n8150), .ZN(n8152)
         );
  INV_X1 U10375 ( .A(n8152), .ZN(n8153) );
  OAI21_X1 U10376 ( .B1(n14107), .B2(n8298), .A(n8153), .ZN(n13844) );
  NAND2_X1 U10377 ( .A1(n8156), .A2(n10112), .ZN(n8157) );
  XNOR2_X1 U10378 ( .A(n8169), .B(SI_21_), .ZN(n8168) );
  XNOR2_X1 U10379 ( .A(n8173), .B(n8168), .ZN(n11888) );
  NAND2_X1 U10380 ( .A1(n11888), .A2(n8347), .ZN(n8159) );
  OR2_X1 U10381 ( .A1(n8005), .A2(n11072), .ZN(n8158) );
  MUX2_X1 U10382 ( .A(n13844), .B(n14236), .S(n7989), .Z(n8160) );
  MUX2_X1 U10383 ( .A(n13844), .B(n14236), .S(n8376), .Z(n8161) );
  NOR2_X1 U10384 ( .A1(n8162), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8163) );
  OR2_X1 U10385 ( .A1(n8178), .A2(n8163), .ZN(n14089) );
  INV_X1 U10386 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n15263) );
  NAND2_X1 U10387 ( .A1(n8320), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10388 ( .A1(n8319), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8164) );
  OAI211_X1 U10389 ( .C1(n8324), .C2(n15263), .A(n8165), .B(n8164), .ZN(n8166)
         );
  INV_X1 U10390 ( .A(n8166), .ZN(n8167) );
  OAI21_X1 U10391 ( .B1(n14089), .B2(n8298), .A(n8167), .ZN(n14105) );
  INV_X1 U10392 ( .A(n8168), .ZN(n8172) );
  INV_X1 U10393 ( .A(n8169), .ZN(n8170) );
  NAND2_X1 U10394 ( .A1(n8170), .A2(SI_21_), .ZN(n8171) );
  INV_X1 U10395 ( .A(SI_22_), .ZN(n8841) );
  NAND2_X1 U10396 ( .A1(n11335), .A2(n9345), .ZN(n8174) );
  MUX2_X1 U10397 ( .A(n14105), .B(n14228), .S(n8376), .Z(n8176) );
  MUX2_X1 U10398 ( .A(n14105), .B(n14228), .S(n7989), .Z(n8175) );
  OR2_X1 U10399 ( .A1(n8178), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U10400 ( .A1(n8178), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8196) );
  AND2_X1 U10401 ( .A1(n8179), .A2(n8196), .ZN(n14075) );
  NAND2_X1 U10402 ( .A1(n14075), .A2(n8180), .ZN(n8185) );
  INV_X1 U10403 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n15125) );
  NAND2_X1 U10404 ( .A1(n8319), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U10405 ( .A1(n8268), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8181) );
  OAI211_X1 U10406 ( .C1(n15125), .C2(n8277), .A(n8182), .B(n8181), .ZN(n8183)
         );
  INV_X1 U10407 ( .A(n8183), .ZN(n8184) );
  NAND2_X1 U10408 ( .A1(n8185), .A2(n8184), .ZN(n13843) );
  NAND2_X1 U10409 ( .A1(n11335), .A2(n8206), .ZN(n8187) );
  NAND2_X1 U10410 ( .A1(n8205), .A2(SI_22_), .ZN(n8186) );
  NAND2_X1 U10411 ( .A1(n8187), .A2(n8186), .ZN(n8189) );
  XNOR2_X1 U10412 ( .A(n8207), .B(SI_23_), .ZN(n8188) );
  NAND2_X1 U10413 ( .A1(n11914), .A2(n8347), .ZN(n8191) );
  INV_X1 U10414 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11356) );
  OR2_X1 U10415 ( .A1(n8005), .A2(n11356), .ZN(n8190) );
  MUX2_X1 U10416 ( .A(n13843), .B(n14074), .S(n7989), .Z(n8194) );
  MUX2_X1 U10417 ( .A(n13843), .B(n14074), .S(n8376), .Z(n8192) );
  NAND2_X1 U10418 ( .A1(n8268), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8201) );
  INV_X1 U10419 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8195) );
  OR2_X1 U10420 ( .A1(n8277), .A2(n8195), .ZN(n8200) );
  NAND2_X1 U10421 ( .A1(n8197), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8217) );
  OAI21_X1 U10422 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8197), .A(n8217), .ZN(
        n14059) );
  OR2_X1 U10423 ( .A1(n8298), .A2(n14059), .ZN(n8199) );
  INV_X1 U10424 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14060) );
  OR2_X1 U10425 ( .A1(n8269), .A2(n14060), .ZN(n8198) );
  NAND4_X1 U10426 ( .A1(n8201), .A2(n8200), .A3(n8199), .A4(n8198), .ZN(n13842) );
  INV_X1 U10427 ( .A(n8207), .ZN(n8202) );
  INV_X1 U10428 ( .A(SI_23_), .ZN(n10923) );
  NAND2_X1 U10429 ( .A1(n8202), .A2(n10923), .ZN(n8208) );
  OAI21_X1 U10430 ( .B1(SI_22_), .B2(n8206), .A(n8208), .ZN(n8203) );
  INV_X1 U10431 ( .A(n8203), .ZN(n8204) );
  NAND2_X1 U10432 ( .A1(n8205), .A2(n8204), .ZN(n8211) );
  INV_X1 U10433 ( .A(n8206), .ZN(n11334) );
  NOR2_X1 U10434 ( .A1(n11334), .A2(n8841), .ZN(n8209) );
  AOI22_X1 U10435 ( .A1(n8209), .A2(n8208), .B1(n8207), .B2(SI_23_), .ZN(n8210) );
  XNOR2_X1 U10436 ( .A(n8226), .B(SI_24_), .ZN(n8223) );
  XNOR2_X1 U10437 ( .A(n8225), .B(n8223), .ZN(n11930) );
  NAND2_X1 U10438 ( .A1(n11930), .A2(n8347), .ZN(n8213) );
  INV_X1 U10439 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11608) );
  OR2_X1 U10440 ( .A1(n8005), .A2(n11608), .ZN(n8212) );
  MUX2_X1 U10441 ( .A(n13842), .B(n14216), .S(n8376), .Z(n8215) );
  MUX2_X1 U10442 ( .A(n13842), .B(n14216), .S(n7989), .Z(n8214) );
  NAND2_X1 U10443 ( .A1(n8319), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8222) );
  INV_X1 U10444 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8216) );
  OR2_X1 U10445 ( .A1(n8324), .A2(n8216), .ZN(n8221) );
  NAND2_X1 U10446 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8218), .ZN(n8240) );
  OAI21_X1 U10447 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8218), .A(n8240), .ZN(
        n14038) );
  OR2_X1 U10448 ( .A1(n8298), .A2(n14038), .ZN(n8220) );
  INV_X1 U10449 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n15307) );
  OR2_X1 U10450 ( .A1(n8277), .A2(n15307), .ZN(n8219) );
  NAND4_X1 U10451 ( .A1(n8222), .A2(n8221), .A3(n8220), .A4(n8219), .ZN(n13841) );
  INV_X1 U10452 ( .A(n8223), .ZN(n8224) );
  NAND2_X1 U10453 ( .A1(n8226), .A2(SI_24_), .ZN(n8227) );
  INV_X1 U10454 ( .A(SI_25_), .ZN(n15275) );
  NAND2_X1 U10455 ( .A1(n8229), .A2(n15275), .ZN(n8249) );
  INV_X1 U10456 ( .A(n8229), .ZN(n8230) );
  NAND2_X1 U10457 ( .A1(n8230), .A2(SI_25_), .ZN(n8231) );
  NAND2_X1 U10458 ( .A1(n8249), .A2(n8231), .ZN(n8247) );
  XNOR2_X1 U10459 ( .A(n8248), .B(n8247), .ZN(n11945) );
  NAND2_X1 U10460 ( .A1(n11945), .A2(n8347), .ZN(n8233) );
  OR2_X1 U10461 ( .A1(n8005), .A2(n15151), .ZN(n8232) );
  MUX2_X1 U10462 ( .A(n13841), .B(n14209), .S(n7989), .Z(n8236) );
  MUX2_X1 U10463 ( .A(n13841), .B(n14209), .S(n8376), .Z(n8234) );
  NAND2_X1 U10464 ( .A1(n8319), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8246) );
  INV_X1 U10465 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8237) );
  OR2_X1 U10466 ( .A1(n8324), .A2(n8237), .ZN(n8245) );
  INV_X1 U10467 ( .A(n8240), .ZN(n8238) );
  INV_X1 U10468 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U10469 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  NAND2_X1 U10470 ( .A1(n8272), .A2(n8241), .ZN(n14026) );
  OR2_X1 U10471 ( .A1(n8298), .A2(n14026), .ZN(n8244) );
  INV_X1 U10472 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8242) );
  OR2_X1 U10473 ( .A1(n8277), .A2(n8242), .ZN(n8243) );
  NAND4_X1 U10474 ( .A1(n8246), .A2(n8245), .A3(n8244), .A4(n8243), .ZN(n14004) );
  XNOR2_X1 U10475 ( .A(n8260), .B(SI_26_), .ZN(n8250) );
  NAND2_X1 U10476 ( .A1(n11967), .A2(n8347), .ZN(n8252) );
  OR2_X1 U10477 ( .A1(n8005), .A2(n8483), .ZN(n8251) );
  MUX2_X1 U10478 ( .A(n14004), .B(n14201), .S(n8376), .Z(n8254) );
  MUX2_X1 U10479 ( .A(n14004), .B(n14201), .S(n7989), .Z(n8253) );
  NAND2_X1 U10480 ( .A1(n8268), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8259) );
  INV_X1 U10481 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14014) );
  OR2_X1 U10482 ( .A1(n8269), .A2(n14014), .ZN(n8258) );
  INV_X1 U10483 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8271) );
  XNOR2_X1 U10484 ( .A(n8272), .B(n8271), .ZN(n14013) );
  OR2_X1 U10485 ( .A1(n8298), .A2(n14013), .ZN(n8257) );
  INV_X1 U10486 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8255) );
  OR2_X1 U10487 ( .A1(n8277), .A2(n8255), .ZN(n8256) );
  NAND4_X1 U10488 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n13840) );
  INV_X1 U10489 ( .A(SI_26_), .ZN(n12697) );
  INV_X1 U10490 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14303) );
  XNOR2_X1 U10491 ( .A(n8282), .B(SI_27_), .ZN(n8262) );
  NAND2_X1 U10492 ( .A1(n13576), .A2(n8347), .ZN(n8264) );
  OR2_X1 U10493 ( .A1(n8005), .A2(n14303), .ZN(n8263) );
  MUX2_X1 U10494 ( .A(n13840), .B(n14195), .S(n7989), .Z(n8267) );
  MUX2_X1 U10495 ( .A(n13840), .B(n14195), .S(n8376), .Z(n8265) );
  NAND2_X1 U10496 ( .A1(n8268), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8281) );
  INV_X1 U10497 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n11598) );
  OR2_X1 U10498 ( .A1(n8269), .A2(n11598), .ZN(n8280) );
  INV_X1 U10499 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8270) );
  OAI21_X1 U10500 ( .B1(n8272), .B2(n8271), .A(n8270), .ZN(n8275) );
  INV_X1 U10501 ( .A(n8272), .ZN(n8274) );
  AND2_X1 U10502 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n8273) );
  NAND2_X1 U10503 ( .A1(n8274), .A2(n8273), .ZN(n13988) );
  NAND2_X1 U10504 ( .A1(n8275), .A2(n13988), .ZN(n13748) );
  OR2_X1 U10505 ( .A1(n8298), .A2(n13748), .ZN(n8279) );
  INV_X1 U10506 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8276) );
  OR2_X1 U10507 ( .A1(n8277), .A2(n8276), .ZN(n8278) );
  NAND4_X1 U10508 ( .A1(n8281), .A2(n8280), .A3(n8279), .A4(n8278), .ZN(n14003) );
  INV_X1 U10509 ( .A(n8282), .ZN(n8283) );
  NOR2_X1 U10510 ( .A1(n8283), .A2(SI_27_), .ZN(n8285) );
  NAND2_X1 U10511 ( .A1(n8283), .A2(SI_27_), .ZN(n8284) );
  INV_X1 U10512 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11568) );
  INV_X1 U10513 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n11988) );
  INV_X1 U10514 ( .A(SI_28_), .ZN(n11606) );
  NAND2_X1 U10515 ( .A1(n8287), .A2(n11606), .ZN(n8304) );
  INV_X1 U10516 ( .A(n8287), .ZN(n8288) );
  NAND2_X1 U10517 ( .A1(n8288), .A2(SI_28_), .ZN(n8289) );
  NAND2_X1 U10518 ( .A1(n8304), .A2(n8289), .ZN(n8290) );
  NAND2_X1 U10519 ( .A1(n8291), .A2(n8290), .ZN(n8292) );
  NAND2_X1 U10520 ( .A1(n8305), .A2(n8292), .ZN(n11987) );
  NAND2_X1 U10521 ( .A1(n11987), .A2(n6539), .ZN(n8294) );
  OR2_X1 U10522 ( .A1(n8005), .A2(n11568), .ZN(n8293) );
  MUX2_X1 U10523 ( .A(n14003), .B(n13982), .S(n8376), .Z(n8296) );
  MUX2_X1 U10524 ( .A(n14003), .B(n13982), .S(n7989), .Z(n8295) );
  NAND2_X1 U10525 ( .A1(n8319), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8303) );
  INV_X1 U10526 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8297) );
  OR2_X1 U10527 ( .A1(n8324), .A2(n8297), .ZN(n8302) );
  OR2_X1 U10528 ( .A1(n8298), .A2(n13988), .ZN(n8301) );
  INV_X1 U10529 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8299) );
  OR2_X1 U10530 ( .A1(n8277), .A2(n8299), .ZN(n8300) );
  NAND4_X1 U10531 ( .A1(n8303), .A2(n8302), .A3(n8301), .A4(n8300), .ZN(n13839) );
  INV_X1 U10532 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14301) );
  INV_X1 U10533 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13570) );
  INV_X1 U10534 ( .A(SI_29_), .ZN(n12689) );
  NAND2_X1 U10535 ( .A1(n8306), .A2(n12689), .ZN(n8326) );
  INV_X1 U10536 ( .A(n8306), .ZN(n8307) );
  NAND2_X1 U10537 ( .A1(n8307), .A2(SI_29_), .ZN(n8308) );
  AND2_X1 U10538 ( .A1(n8326), .A2(n8308), .ZN(n8309) );
  NAND2_X1 U10539 ( .A1(n13568), .A2(n8347), .ZN(n8313) );
  OR2_X1 U10540 ( .A1(n8005), .A2(n14301), .ZN(n8312) );
  MUX2_X1 U10541 ( .A(n13839), .B(n13985), .S(n7989), .Z(n8316) );
  MUX2_X1 U10542 ( .A(n13839), .B(n13985), .S(n8376), .Z(n8314) );
  INV_X1 U10543 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15170) );
  NAND2_X1 U10544 ( .A1(n8319), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10545 ( .A1(n8320), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8317) );
  OAI211_X1 U10546 ( .C1(n8324), .C2(n15170), .A(n8318), .B(n8317), .ZN(n13975) );
  NAND2_X1 U10547 ( .A1(n7353), .A2(n9601), .ZN(n9513) );
  INV_X1 U10548 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10549 ( .A1(n8319), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U10550 ( .A1(n8320), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8321) );
  OAI211_X1 U10551 ( .C1(n8324), .C2(n8323), .A(n8322), .B(n8321), .ZN(n13987)
         );
  OAI21_X1 U10552 ( .B1(n13975), .B2(n9513), .A(n13987), .ZN(n8325) );
  INV_X1 U10553 ( .A(n8325), .ZN(n8330) );
  INV_X1 U10554 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11771) );
  INV_X1 U10555 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13566) );
  MUX2_X1 U10556 ( .A(n11771), .B(n13566), .S(n9343), .Z(n8338) );
  XNOR2_X1 U10557 ( .A(n8338), .B(SI_30_), .ZN(n8337) );
  NAND2_X1 U10558 ( .A1(n12964), .A2(n8347), .ZN(n8329) );
  OR2_X1 U10559 ( .A1(n8005), .A2(n11771), .ZN(n8328) );
  MUX2_X1 U10560 ( .A(n8330), .B(n13978), .S(n8376), .Z(n8336) );
  NAND2_X1 U10561 ( .A1(n13975), .A2(n8376), .ZN(n8377) );
  NAND2_X1 U10562 ( .A1(n8331), .A2(n11073), .ZN(n8333) );
  INV_X1 U10563 ( .A(n13987), .ZN(n8332) );
  AOI21_X1 U10564 ( .B1(n8377), .B2(n8333), .A(n8332), .ZN(n8334) );
  AOI21_X1 U10565 ( .B1(n13978), .B2(n7989), .A(n8334), .ZN(n8335) );
  INV_X1 U10566 ( .A(n8337), .ZN(n8341) );
  INV_X1 U10567 ( .A(n8338), .ZN(n8339) );
  NAND2_X1 U10568 ( .A1(n8339), .A2(SI_30_), .ZN(n8340) );
  MUX2_X1 U10569 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9343), .Z(n8343) );
  XNOR2_X1 U10570 ( .A(n8343), .B(SI_31_), .ZN(n8344) );
  XOR2_X1 U10571 ( .A(n13975), .B(n14171), .Z(n8354) );
  NAND2_X1 U10572 ( .A1(n8348), .A2(n7353), .ZN(n9588) );
  NAND2_X1 U10573 ( .A1(n8349), .A2(n10973), .ZN(n8350) );
  NAND2_X1 U10574 ( .A1(n9588), .A2(n8350), .ZN(n8351) );
  OR2_X1 U10575 ( .A1(n9591), .A2(n11295), .ZN(n10360) );
  NAND2_X1 U10576 ( .A1(n8351), .A2(n10360), .ZN(n8381) );
  INV_X1 U10577 ( .A(n8381), .ZN(n8352) );
  AND2_X1 U10578 ( .A1(n8354), .A2(n8352), .ZN(n8353) );
  NAND2_X1 U10579 ( .A1(n8387), .A2(n8353), .ZN(n8384) );
  INV_X1 U10580 ( .A(n8354), .ZN(n8375) );
  XNOR2_X1 U10581 ( .A(n14175), .B(n13987), .ZN(n8370) );
  XNOR2_X1 U10582 ( .A(n13985), .B(n13839), .ZN(n13997) );
  NOR2_X1 U10583 ( .A1(n14042), .A2(n13841), .ZN(n11594) );
  AOI21_X1 U10584 ( .B1(n14042), .B2(n13841), .A(n11594), .ZN(n14047) );
  XNOR2_X1 U10585 ( .A(n14244), .B(n14137), .ZN(n14126) );
  INV_X1 U10586 ( .A(n14149), .ZN(n14162) );
  XNOR2_X1 U10587 ( .A(n13610), .B(n14427), .ZN(n11308) );
  NAND2_X1 U10588 ( .A1(n11455), .A2(n8355), .ZN(n11456) );
  XNOR2_X1 U10589 ( .A(n13601), .B(n13847), .ZN(n11189) );
  INV_X1 U10590 ( .A(n13850), .ZN(n11025) );
  XNOR2_X1 U10591 ( .A(n14616), .B(n11025), .ZN(n10627) );
  INV_X1 U10592 ( .A(n13851), .ZN(n10624) );
  XNOR2_X1 U10593 ( .A(n10689), .B(n10679), .ZN(n10554) );
  XNOR2_X1 U10594 ( .A(n10612), .B(n13853), .ZN(n10546) );
  AND2_X1 U10595 ( .A1(n10456), .A2(n13855), .ZN(n10443) );
  NOR2_X1 U10596 ( .A1(n10456), .A2(n13855), .ZN(n10445) );
  NOR2_X1 U10597 ( .A1(n10443), .A2(n10445), .ZN(n10023) );
  NAND2_X1 U10598 ( .A1(n8358), .A2(n8357), .ZN(n10317) );
  NOR4_X1 U10599 ( .A1(n10023), .A2(n10012), .A3(n10009), .A4(n10317), .ZN(
        n8359) );
  XNOR2_X1 U10600 ( .A(n10579), .B(n13854), .ZN(n10581) );
  NAND4_X1 U10601 ( .A1(n10546), .A2(n8359), .A3(n10379), .A4(n10581), .ZN(
        n8360) );
  NOR4_X1 U10602 ( .A1(n10627), .A2(n10666), .A3(n10554), .A4(n8360), .ZN(
        n8361) );
  XNOR2_X1 U10603 ( .A(n14504), .B(n13848), .ZN(n11103) );
  XNOR2_X1 U10604 ( .A(n11345), .B(n13849), .ZN(n10786) );
  NAND4_X1 U10605 ( .A1(n11189), .A2(n8361), .A3(n11103), .A4(n10786), .ZN(
        n8362) );
  NOR4_X1 U10606 ( .A1(n6959), .A2(n11308), .A3(n11456), .A4(n8362), .ZN(n8364) );
  XNOR2_X1 U10607 ( .A(n14450), .B(n14458), .ZN(n11460) );
  INV_X1 U10608 ( .A(n11578), .ZN(n8363) );
  NAND2_X1 U10609 ( .A1(n8363), .A2(n11577), .ZN(n11472) );
  NAND3_X1 U10610 ( .A1(n8364), .A2(n11460), .A3(n11472), .ZN(n8365) );
  NOR4_X1 U10611 ( .A1(n14126), .A2(n14133), .A3(n14162), .A4(n8365), .ZN(
        n8366) );
  XNOR2_X1 U10612 ( .A(n14236), .B(n13844), .ZN(n14097) );
  NAND4_X1 U10613 ( .A1(n14047), .A2(n8366), .A3(n14053), .A4(n14097), .ZN(
        n8367) );
  XOR2_X1 U10614 ( .A(n13843), .B(n14074), .Z(n14068) );
  XNOR2_X1 U10615 ( .A(n14201), .B(n13772), .ZN(n14022) );
  NOR4_X1 U10616 ( .A1(n8367), .A2(n14068), .A3(n14022), .A4(n14087), .ZN(
        n8368) );
  XNOR2_X1 U10617 ( .A(n13982), .B(n14003), .ZN(n11596) );
  NAND4_X1 U10618 ( .A1(n13997), .A2(n8368), .A3(n14005), .A4(n11596), .ZN(
        n8369) );
  NOR3_X1 U10619 ( .A1(n8375), .A2(n8370), .A3(n8369), .ZN(n8371) );
  XNOR2_X1 U10620 ( .A(n8371), .B(n10792), .ZN(n8372) );
  NAND2_X1 U10621 ( .A1(n11073), .A2(n9601), .ZN(n8373) );
  NAND2_X1 U10622 ( .A1(n8381), .A2(n8373), .ZN(n8385) );
  INV_X1 U10623 ( .A(n8385), .ZN(n8374) );
  NAND2_X1 U10624 ( .A1(n8375), .A2(n8374), .ZN(n8380) );
  MUX2_X1 U10625 ( .A(n8376), .B(n13975), .S(n14171), .Z(n8378) );
  INV_X1 U10626 ( .A(n8386), .ZN(n8379) );
  MUX2_X1 U10627 ( .A(n8381), .B(n8380), .S(n8379), .Z(n8382) );
  NAND2_X1 U10628 ( .A1(n8384), .A2(n7555), .ZN(n8395) );
  NAND2_X1 U10629 ( .A1(n8389), .A2(n8388), .ZN(n8396) );
  NAND2_X1 U10630 ( .A1(n8396), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8391) );
  INV_X1 U10631 ( .A(n9315), .ZN(n8392) );
  NAND2_X1 U10632 ( .A1(n8392), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11354) );
  INV_X1 U10633 ( .A(n11354), .ZN(n8393) );
  OAI21_X1 U10634 ( .B1(n8395), .B2(n8394), .A(n8393), .ZN(n8410) );
  XNOR2_X1 U10635 ( .A(n8398), .B(n8397), .ZN(n11610) );
  OAI21_X1 U10636 ( .B1(n7687), .B2(n8399), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8400) );
  MUX2_X1 U10637 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8400), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8401) );
  NAND2_X1 U10638 ( .A1(n8401), .A2(n8402), .ZN(n11372) );
  MUX2_X1 U10639 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8403), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8405) );
  NAND2_X1 U10640 ( .A1(n8405), .A2(n8404), .ZN(n11450) );
  AND2_X1 U10641 ( .A1(n10973), .A2(n11295), .ZN(n9586) );
  OAI21_X1 U10642 ( .B1(n9588), .B2(n9586), .A(n9315), .ZN(n8406) );
  INV_X1 U10643 ( .A(n8406), .ZN(n8407) );
  NAND2_X1 U10644 ( .A1(n9595), .A2(n8407), .ZN(n9608) );
  NOR2_X1 U10645 ( .A1(n9608), .A2(P1_U3086), .ZN(n9505) );
  INV_X1 U10646 ( .A(n6530), .ZN(n14542) );
  INV_X1 U10647 ( .A(n9588), .ZN(n9316) );
  INV_X1 U10648 ( .A(n13873), .ZN(n13878) );
  NAND3_X1 U10649 ( .A1(n9505), .A2(n14542), .A3(n14154), .ZN(n8408) );
  OAI211_X1 U10650 ( .C1(n8348), .C2(n11354), .A(n8408), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8409) );
  NAND2_X1 U10651 ( .A1(n8410), .A2(n8409), .ZN(P1_U3242) );
  NAND2_X1 U10652 ( .A1(n8577), .A2(n8576), .ZN(n8593) );
  INV_X1 U10653 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U10654 ( .A1(n8714), .A2(n8713), .ZN(n8731) );
  INV_X1 U10655 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15228) );
  INV_X1 U10656 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U10657 ( .A1(n15228), .A2(n8746), .ZN(n8411) );
  INV_X1 U10658 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12129) );
  INV_X1 U10659 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15188) );
  NOR2_X1 U10660 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(P3_REG3_REG_22__SCAN_IN), 
        .ZN(n8412) );
  INV_X1 U10661 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n8500) );
  INV_X1 U10662 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n12055) );
  NOR2_X1 U10663 ( .A1(n8870), .A2(n12055), .ZN(n8413) );
  NOR2_X1 U10664 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n8423) );
  NAND4_X1 U10665 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .ZN(n8424)
         );
  XNOR2_X2 U10667 ( .A(n8432), .B(n8431), .ZN(n8434) );
  INV_X1 U10668 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10669 ( .A1(n6533), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U10670 ( .A1(n8913), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8436) );
  OAI211_X1 U10671 ( .C1(n8438), .C2(n11767), .A(n8437), .B(n8436), .ZN(n8439)
         );
  INV_X1 U10672 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11915) );
  NAND2_X1 U10673 ( .A1(n8517), .A2(n8533), .ZN(n8442) );
  INV_X1 U10674 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9347) );
  NAND2_X1 U10675 ( .A1(n9347), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U10676 ( .A1(n8442), .A2(n8441), .ZN(n8548) );
  AND2_X1 U10677 ( .A1(n9526), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U10678 ( .A1(n9641), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10679 ( .A1(n9150), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U10680 ( .A1(n9148), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10681 ( .A1(n8448), .A2(n8447), .ZN(n8569) );
  NAND2_X1 U10682 ( .A1(n9153), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U10683 ( .A1(n9156), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U10684 ( .A1(n9167), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U10685 ( .A1(n8452), .A2(n8451), .ZN(n8620) );
  NOR2_X1 U10686 ( .A1(n10496), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10687 ( .A1(n10496), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U10688 ( .A1(n9309), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10689 ( .A1(n9308), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U10690 ( .A1(n9577), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10691 ( .A1(n9580), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8458) );
  XNOR2_X1 U10692 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8693) );
  NAND2_X1 U10693 ( .A1(n8694), .A2(n8693), .ZN(n8461) );
  NAND2_X1 U10694 ( .A1(n9714), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8460) );
  XNOR2_X2 U10695 ( .A(n8463), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U10696 ( .A1(n8463), .A2(n8462), .ZN(n8464) );
  NOR2_X1 U10697 ( .A1(n10078), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U10698 ( .A1(n10078), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10699 ( .A1(n10300), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8469) );
  INV_X1 U10700 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U10701 ( .A1(n10305), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10702 ( .A1(n8469), .A2(n8468), .ZN(n8739) );
  NAND2_X1 U10703 ( .A1(n15244), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U10704 ( .A1(n10081), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U10705 ( .A1(n10244), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8472) );
  INV_X1 U10706 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10636) );
  NAND2_X1 U10707 ( .A1(n10636), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U10708 ( .A1(n15116), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8476) );
  INV_X1 U10709 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10799) );
  NAND2_X1 U10710 ( .A1(n10799), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10711 ( .A1(n8476), .A2(n8475), .ZN(n8802) );
  AOI22_X1 U10712 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(
        P1_DATAO_REG_20__SCAN_IN), .B1(n11869), .B2(n10972), .ZN(n8820) );
  AOI22_X1 U10713 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n15216), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n11072), .ZN(n8831) );
  INV_X1 U10714 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n15290) );
  AOI22_X1 U10715 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n15205), .B2(n15290), .ZN(n8839) );
  AOI22_X1 U10716 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n11915), .B2(n11356), .ZN(n8506) );
  NOR2_X1 U10717 ( .A1(n8507), .A2(n8506), .ZN(n8479) );
  NAND2_X1 U10718 ( .A1(n8480), .A2(n11608), .ZN(n8481) );
  AOI22_X1 U10719 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n15291), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n15151), .ZN(n8853) );
  OAI21_X2 U10720 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(n15291), .A(n8482), 
        .ZN(n8866) );
  AOI22_X1 U10721 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n15117), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8483), .ZN(n8864) );
  AOI22_X1 U10722 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13579), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n14303), .ZN(n8880) );
  INV_X1 U10723 ( .A(n8880), .ZN(n8486) );
  XNOR2_X1 U10724 ( .A(n8879), .B(n8486), .ZN(n12690) );
  XNOR2_X2 U10725 ( .A(n8488), .B(n8487), .ZN(n11833) );
  NAND2_X1 U10726 ( .A1(n8537), .A2(n6967), .ZN(n8534) );
  NAND2_X1 U10727 ( .A1(n12690), .A2(n11774), .ZN(n8492) );
  NAND2_X1 U10728 ( .A1(n8537), .A2(n9343), .ZN(n8530) );
  BUF_X2 U10729 ( .A(n6529), .Z(n11775) );
  INV_X1 U10730 ( .A(SI_27_), .ZN(n12692) );
  OR2_X1 U10731 ( .A1(n11775), .A2(n12692), .ZN(n8491) );
  INV_X1 U10732 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10733 ( .A1(n8502), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U10734 ( .A1(n8858), .A2(n8493), .ZN(n12435) );
  NAND2_X1 U10735 ( .A1(n12435), .A2(n8897), .ZN(n8495) );
  AOI22_X1 U10736 ( .A1(n6532), .A2(P3_REG0_REG_24__SCAN_IN), .B1(n8913), .B2(
        P3_REG1_REG_24__SCAN_IN), .ZN(n8494) );
  OAI211_X1 U10737 ( .C1(n11767), .C2(n8496), .A(n8495), .B(n8494), .ZN(n12445) );
  INV_X1 U10738 ( .A(n12445), .ZN(n12066) );
  INV_X1 U10739 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11931) );
  XNOR2_X1 U10740 ( .A(n11931), .B(n8497), .ZN(n11329) );
  NAND2_X1 U10741 ( .A1(n11329), .A2(n11774), .ZN(n8499) );
  INV_X1 U10742 ( .A(SI_24_), .ZN(n11331) );
  OR2_X1 U10743 ( .A1(n6529), .A2(n11331), .ZN(n8498) );
  INV_X1 U10744 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n8505) );
  OR2_X1 U10745 ( .A1(n8846), .A2(n8500), .ZN(n8501) );
  NAND2_X1 U10746 ( .A1(n8502), .A2(n8501), .ZN(n12448) );
  NAND2_X1 U10747 ( .A1(n12448), .A2(n8897), .ZN(n8504) );
  AOI22_X1 U10748 ( .A1(n6533), .A2(P3_REG0_REG_23__SCAN_IN), .B1(n8913), .B2(
        P3_REG1_REG_23__SCAN_IN), .ZN(n8503) );
  OAI211_X1 U10749 ( .C1(n11767), .C2(n8505), .A(n8504), .B(n8503), .ZN(n12456) );
  INV_X1 U10750 ( .A(n12456), .ZN(n12162) );
  XNOR2_X1 U10751 ( .A(n8507), .B(n8506), .ZN(n10921) );
  NAND2_X1 U10752 ( .A1(n10921), .A2(n11774), .ZN(n8509) );
  OR2_X1 U10753 ( .A1(n11775), .A2(n10923), .ZN(n8508) );
  INV_X1 U10754 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9033) );
  OR2_X1 U10755 ( .A1(n8563), .A2(n9033), .ZN(n8513) );
  INV_X1 U10756 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9034) );
  OR2_X1 U10757 ( .A1(n11767), .A2(n9034), .ZN(n8512) );
  INV_X1 U10758 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n9998) );
  MUX2_X1 U10759 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8514), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n8516) );
  INV_X1 U10760 ( .A(n9084), .ZN(n8515) );
  INV_X1 U10761 ( .A(n9677), .ZN(n9035) );
  INV_X1 U10762 ( .A(SI_1_), .ZN(n9114) );
  OR2_X1 U10763 ( .A1(n8530), .A2(n9114), .ZN(n8520) );
  INV_X1 U10764 ( .A(n8533), .ZN(n8518) );
  XNOR2_X1 U10765 ( .A(n8518), .B(n8517), .ZN(n9115) );
  OR2_X1 U10766 ( .A1(n8534), .A2(n9115), .ZN(n8519) );
  INV_X1 U10767 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10253) );
  OR2_X1 U10768 ( .A1(n6537), .A2(n10253), .ZN(n8526) );
  INV_X1 U10769 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n8523) );
  INV_X1 U10770 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8524) );
  OR2_X1 U10771 ( .A1(n8814), .A2(n8524), .ZN(n8525) );
  INV_X1 U10772 ( .A(n11767), .ZN(n8527) );
  NAND2_X1 U10773 ( .A1(n8527), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8528) );
  INV_X1 U10774 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9121) );
  OR2_X1 U10775 ( .A1(n6529), .A2(n9119), .ZN(n8536) );
  AND2_X1 U10776 ( .A1(n8531), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8532) );
  NOR2_X1 U10777 ( .A1(n8533), .A2(n8532), .ZN(n9120) );
  OR2_X1 U10778 ( .A1(n6527), .A2(n9120), .ZN(n8535) );
  OAI211_X1 U10779 ( .C1(n9121), .C2(n9078), .A(n8536), .B(n8535), .ZN(n10255)
         );
  NAND2_X1 U10780 ( .A1(n9983), .A2(n9990), .ZN(n8539) );
  OR2_X1 U10781 ( .A1(n6823), .A2(n8521), .ZN(n8538) );
  NAND2_X1 U10782 ( .A1(n8539), .A2(n8538), .ZN(n14929) );
  NAND2_X1 U10783 ( .A1(n6533), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8544) );
  INV_X1 U10784 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n14925) );
  INV_X1 U10785 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9086) );
  OR2_X1 U10786 ( .A1(n11767), .A2(n9086), .ZN(n8542) );
  INV_X1 U10787 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9070) );
  OR2_X1 U10788 ( .A1(n6518), .A2(n9070), .ZN(n8541) );
  NOR2_X1 U10789 ( .A1(n9084), .A2(n8429), .ZN(n8545) );
  INV_X1 U10790 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8546) );
  XNOR2_X1 U10791 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8547) );
  XNOR2_X1 U10792 ( .A(n8548), .B(n8547), .ZN(n9137) );
  OR2_X1 U10793 ( .A1(n6527), .A2(n9137), .ZN(n8550) );
  OR2_X1 U10794 ( .A1(n6529), .A2(SI_2_), .ZN(n8549) );
  INV_X1 U10795 ( .A(n14924), .ZN(n8551) );
  NOR2_X1 U10796 ( .A1(n14945), .A2(n8551), .ZN(n8552) );
  NAND2_X1 U10797 ( .A1(n6532), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8556) );
  OR2_X1 U10798 ( .A1(n6537), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8555) );
  INV_X1 U10799 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10428) );
  OR2_X1 U10800 ( .A1(n11767), .A2(n10428), .ZN(n8554) );
  INV_X1 U10801 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n9044) );
  OR2_X1 U10802 ( .A1(n6518), .A2(n9044), .ZN(n8553) );
  XNOR2_X1 U10803 ( .A(n8557), .B(P3_IR_REG_3__SCAN_IN), .ZN(n9139) );
  XNOR2_X1 U10804 ( .A(n9641), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n8558) );
  XNOR2_X1 U10805 ( .A(n8559), .B(n8558), .ZN(n9140) );
  OR2_X1 U10806 ( .A1(n6527), .A2(n9140), .ZN(n8561) );
  OR2_X1 U10807 ( .A1(n6529), .A2(SI_3_), .ZN(n8560) );
  OAI211_X1 U10808 ( .C1(n9139), .C2(n9078), .A(n8561), .B(n8560), .ZN(n10229)
         );
  OR2_X1 U10809 ( .A1(n14911), .A2(n10229), .ZN(n11641) );
  NAND2_X1 U10810 ( .A1(n14911), .A2(n10229), .ZN(n11646) );
  NAND2_X1 U10811 ( .A1(n6533), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8567) );
  AND2_X1 U10812 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8562) );
  NOR2_X1 U10813 ( .A1(n8577), .A2(n8562), .ZN(n14921) );
  OR2_X1 U10814 ( .A1(n6537), .A2(n14921), .ZN(n8566) );
  INV_X1 U10815 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9048) );
  OR2_X1 U10816 ( .A1(n11767), .A2(n9048), .ZN(n8565) );
  INV_X1 U10817 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9073) );
  OR2_X1 U10818 ( .A1(n8563), .A2(n9073), .ZN(n8564) );
  NAND2_X1 U10819 ( .A1(n8570), .A2(n8569), .ZN(n8571) );
  AND2_X1 U10820 ( .A1(n8572), .A2(n8571), .ZN(n9143) );
  OR2_X1 U10821 ( .A1(n6527), .A2(n9143), .ZN(n8574) );
  NAND2_X1 U10822 ( .A1(n12206), .A2(n10322), .ZN(n11645) );
  NAND2_X1 U10823 ( .A1(n11650), .A2(n11645), .ZN(n8927) );
  INV_X1 U10824 ( .A(n10229), .ZN(n14971) );
  AND2_X1 U10825 ( .A1(n14911), .A2(n14971), .ZN(n14906) );
  INV_X1 U10826 ( .A(n10322), .ZN(n14973) );
  AOI22_X1 U10827 ( .A1(n8927), .A2(n14906), .B1(n14973), .B2(n12206), .ZN(
        n8575) );
  NAND2_X1 U10828 ( .A1(n6533), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8582) );
  INV_X1 U10829 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9053) );
  OR2_X1 U10830 ( .A1(n6518), .A2(n9053), .ZN(n8581) );
  OR2_X1 U10831 ( .A1(n8577), .A2(n8576), .ZN(n8578) );
  AND2_X1 U10832 ( .A1(n8593), .A2(n8578), .ZN(n10542) );
  OR2_X1 U10833 ( .A1(n6538), .A2(n10542), .ZN(n8580) );
  INV_X1 U10834 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10438) );
  OR2_X1 U10835 ( .A1(n11767), .A2(n10438), .ZN(n8579) );
  NAND4_X1 U10836 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(n14910) );
  NAND2_X1 U10837 ( .A1(n8584), .A2(n8583), .ZN(n8602) );
  NAND2_X1 U10838 ( .A1(n8602), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8585) );
  XNOR2_X1 U10839 ( .A(n8585), .B(P3_IR_REG_5__SCAN_IN), .ZN(n9091) );
  OAI21_X1 U10840 ( .B1(n8588), .B2(n8587), .A(n8586), .ZN(n9116) );
  INV_X1 U10841 ( .A(n9116), .ZN(n8589) );
  OR2_X1 U10842 ( .A1(n6527), .A2(n8589), .ZN(n8591) );
  OR2_X1 U10843 ( .A1(n11775), .A2(SI_5_), .ZN(n8590) );
  OAI211_X1 U10844 ( .C1(n9091), .C2(n9078), .A(n8591), .B(n8590), .ZN(n11655)
         );
  XNOR2_X1 U10845 ( .A(n14910), .B(n11655), .ZN(n10434) );
  INV_X1 U10846 ( .A(n11655), .ZN(n14981) );
  OR2_X1 U10847 ( .A1(n14910), .A2(n14981), .ZN(n8592) );
  NAND2_X1 U10848 ( .A1(n6533), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8598) );
  INV_X1 U10849 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9057) );
  OR2_X1 U10850 ( .A1(n6518), .A2(n9057), .ZN(n8597) );
  NAND2_X1 U10851 ( .A1(n8593), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8594) );
  AND2_X1 U10852 ( .A1(n8611), .A2(n8594), .ZN(n12181) );
  OR2_X1 U10853 ( .A1(n6538), .A2(n12181), .ZN(n8596) );
  INV_X1 U10854 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10915) );
  OR2_X1 U10855 ( .A1(n11767), .A2(n10915), .ZN(n8595) );
  INV_X1 U10856 ( .A(SI_6_), .ZN(n9130) );
  OR2_X1 U10857 ( .A1(n6529), .A2(n9130), .ZN(n8609) );
  INV_X1 U10858 ( .A(n8599), .ZN(n8600) );
  XNOR2_X1 U10859 ( .A(n8601), .B(n8600), .ZN(n9131) );
  OR2_X1 U10860 ( .A1(n6527), .A2(n9131), .ZN(n8608) );
  OAI21_X1 U10861 ( .B1(n8602), .B2(P3_IR_REG_5__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8603) );
  MUX2_X1 U10862 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8603), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n8606) );
  BUF_X1 U10863 ( .A(n8604), .Z(n8605) );
  NAND2_X1 U10864 ( .A1(n8606), .A2(n8605), .ZN(n10045) );
  INV_X1 U10865 ( .A(n10045), .ZN(n9058) );
  NAND2_X1 U10866 ( .A1(n8808), .A2(n9058), .ZN(n8607) );
  NAND2_X1 U10867 ( .A1(n12205), .A2(n10916), .ZN(n11658) );
  INV_X1 U10868 ( .A(n10916), .ZN(n12180) );
  NAND2_X1 U10869 ( .A1(n12205), .A2(n12180), .ZN(n8610) );
  NAND2_X1 U10870 ( .A1(n6532), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8616) );
  INV_X1 U10871 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10034) );
  OR2_X1 U10872 ( .A1(n6518), .A2(n10034), .ZN(n8615) );
  AND2_X1 U10873 ( .A1(n8611), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8612) );
  NOR2_X1 U10874 ( .A1(n8627), .A2(n8612), .ZN(n10868) );
  OR2_X1 U10875 ( .A1(n6537), .A2(n10868), .ZN(n8614) );
  INV_X1 U10876 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10035) );
  OR2_X1 U10877 ( .A1(n11767), .A2(n10035), .ZN(n8613) );
  NAND4_X1 U10878 ( .A1(n8616), .A2(n8615), .A3(n8614), .A4(n8613), .ZN(n12204) );
  NAND2_X1 U10879 ( .A1(n8605), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8617) );
  MUX2_X1 U10880 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8617), .S(
        P3_IR_REG_7__SCAN_IN), .Z(n8619) );
  NAND2_X1 U10881 ( .A1(n8619), .A2(n8618), .ZN(n10049) );
  INV_X1 U10882 ( .A(n10049), .ZN(n10147) );
  NAND2_X1 U10883 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  AND2_X1 U10884 ( .A1(n8623), .A2(n8622), .ZN(n9134) );
  OR2_X1 U10885 ( .A1(n6527), .A2(n9134), .ZN(n8625) );
  OR2_X1 U10886 ( .A1(n11775), .A2(SI_7_), .ZN(n8624) );
  OAI211_X1 U10887 ( .C1(n10147), .C2(n9078), .A(n8625), .B(n8624), .ZN(n14994) );
  XNOR2_X1 U10888 ( .A(n12204), .B(n14994), .ZN(n10871) );
  INV_X1 U10889 ( .A(n14994), .ZN(n10862) );
  NAND2_X1 U10890 ( .A1(n12204), .A2(n10862), .ZN(n8626) );
  NAND2_X1 U10891 ( .A1(n6532), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8632) );
  INV_X1 U10892 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10136) );
  OR2_X1 U10893 ( .A1(n6518), .A2(n10136), .ZN(n8631) );
  NOR2_X1 U10894 ( .A1(n8627), .A2(n10154), .ZN(n8628) );
  OR2_X1 U10895 ( .A1(n6537), .A2(n6573), .ZN(n8630) );
  INV_X1 U10896 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10137) );
  OR2_X1 U10897 ( .A1(n11767), .A2(n10137), .ZN(n8629) );
  NAND4_X1 U10898 ( .A1(n8632), .A2(n8631), .A3(n8630), .A4(n8629), .ZN(n12203) );
  NAND2_X1 U10899 ( .A1(n8618), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8634) );
  MUX2_X1 U10900 ( .A(n8634), .B(P3_IR_REG_31__SCAN_IN), .S(n8633), .Z(n8636)
         );
  NOR2_X1 U10901 ( .A1(n8618), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8651) );
  INV_X1 U10902 ( .A(n8651), .ZN(n8635) );
  NAND2_X1 U10903 ( .A1(n8636), .A2(n8635), .ZN(n10487) );
  XNOR2_X1 U10904 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8637) );
  XNOR2_X1 U10905 ( .A(n8638), .B(n8637), .ZN(n9118) );
  OR2_X1 U10906 ( .A1(n6527), .A2(n9118), .ZN(n8640) );
  INV_X1 U10907 ( .A(SI_8_), .ZN(n15203) );
  OR2_X1 U10908 ( .A1(n11775), .A2(n15203), .ZN(n8639) );
  OAI211_X1 U10909 ( .C1(n9078), .C2(n10487), .A(n8640), .B(n8639), .ZN(n11038) );
  OR2_X1 U10910 ( .A1(n12203), .A2(n11038), .ZN(n11044) );
  NAND2_X1 U10911 ( .A1(n6532), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8647) );
  INV_X1 U10912 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10472) );
  OR2_X1 U10913 ( .A1(n6518), .A2(n10472), .ZN(n8646) );
  OR2_X1 U10914 ( .A1(n8642), .A2(n8641), .ZN(n8643) );
  AND2_X1 U10915 ( .A1(n8658), .A2(n8643), .ZN(n11054) );
  OR2_X1 U10916 ( .A1(n6537), .A2(n11054), .ZN(n8645) );
  INV_X1 U10917 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10473) );
  OR2_X1 U10918 ( .A1(n11767), .A2(n10473), .ZN(n8644) );
  NOR2_X1 U10919 ( .A1(n8651), .A2(n8429), .ZN(n8648) );
  MUX2_X1 U10920 ( .A(n8429), .B(n8648), .S(P3_IR_REG_9__SCAN_IN), .Z(n8649)
         );
  INV_X1 U10921 ( .A(n8649), .ZN(n8652) );
  INV_X1 U10922 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U10923 ( .A1(n8651), .A2(n8650), .ZN(n8679) );
  NAND2_X1 U10924 ( .A1(n8652), .A2(n8679), .ZN(n10488) );
  INV_X1 U10925 ( .A(n10488), .ZN(n10708) );
  OR2_X1 U10926 ( .A1(n6529), .A2(SI_9_), .ZN(n8656) );
  XNOR2_X1 U10927 ( .A(n10496), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n8653) );
  XNOR2_X1 U10928 ( .A(n8654), .B(n8653), .ZN(n9132) );
  OR2_X1 U10929 ( .A1(n6527), .A2(n9132), .ZN(n8655) );
  OAI211_X1 U10930 ( .C1(n10708), .C2(n9078), .A(n8656), .B(n8655), .ZN(n10850) );
  INV_X1 U10931 ( .A(n10850), .ZN(n11052) );
  NAND2_X1 U10932 ( .A1(n12202), .A2(n11052), .ZN(n8672) );
  NAND2_X1 U10933 ( .A1(n12202), .A2(n10850), .ZN(n11672) );
  NAND2_X1 U10934 ( .A1(n11673), .A2(n11672), .ZN(n11666) );
  AND2_X1 U10935 ( .A1(n11044), .A2(n8671), .ZN(n11059) );
  NAND2_X1 U10936 ( .A1(n8913), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8663) );
  INV_X1 U10937 ( .A(n6532), .ZN(n8874) );
  INV_X1 U10938 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8657) );
  OR2_X1 U10939 ( .A1(n8874), .A2(n8657), .ZN(n8662) );
  NAND2_X1 U10940 ( .A1(n8658), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8659) );
  AND2_X1 U10941 ( .A1(n8684), .A2(n8659), .ZN(n12078) );
  OR2_X1 U10942 ( .A1(n6538), .A2(n12078), .ZN(n8661) );
  INV_X1 U10943 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10716) );
  OR2_X1 U10944 ( .A1(n11767), .A2(n10716), .ZN(n8660) );
  NAND4_X1 U10945 ( .A1(n8663), .A2(n8662), .A3(n8661), .A4(n8660), .ZN(n14371) );
  OAI21_X1 U10946 ( .B1(n6638), .B2(n8665), .A(n8664), .ZN(n9151) );
  NAND2_X1 U10947 ( .A1(n9151), .A2(n11774), .ZN(n8669) );
  NAND2_X1 U10948 ( .A1(n8679), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8667) );
  XNOR2_X1 U10949 ( .A(n8667), .B(n8666), .ZN(n11080) );
  NAND2_X1 U10950 ( .A1(n8808), .A2(n11080), .ZN(n8668) );
  OAI211_X1 U10951 ( .C1(SI_10_), .C2(n11775), .A(n8669), .B(n8668), .ZN(
        n15014) );
  OR2_X1 U10952 ( .A1(n14371), .A2(n15014), .ZN(n11674) );
  NAND2_X1 U10953 ( .A1(n14371), .A2(n15014), .ZN(n11675) );
  NAND2_X1 U10954 ( .A1(n11674), .A2(n11675), .ZN(n11677) );
  AND2_X1 U10955 ( .A1(n11059), .A2(n11677), .ZN(n8670) );
  NAND2_X1 U10956 ( .A1(n10963), .A2(n8670), .ZN(n8676) );
  INV_X1 U10957 ( .A(n11677), .ZN(n11062) );
  NAND2_X1 U10958 ( .A1(n12203), .A2(n11038), .ZN(n11045) );
  OR2_X1 U10959 ( .A1(n11062), .A2(n11060), .ZN(n8674) );
  INV_X1 U10960 ( .A(n15014), .ZN(n12077) );
  NAND2_X1 U10961 ( .A1(n14371), .A2(n12077), .ZN(n8673) );
  AND2_X1 U10962 ( .A1(n8674), .A2(n8673), .ZN(n8675) );
  XNOR2_X1 U10963 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8677) );
  XNOR2_X1 U10964 ( .A(n8678), .B(n8677), .ZN(n9160) );
  NAND2_X1 U10965 ( .A1(n9160), .A2(n11774), .ZN(n8683) );
  OR2_X1 U10966 ( .A1(n8679), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U10967 ( .A1(n8695), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8681) );
  XNOR2_X1 U10968 ( .A(n8681), .B(n8680), .ZN(n14866) );
  AOI22_X1 U10969 ( .A1(n8809), .A2(n9161), .B1(n8808), .B2(n14866), .ZN(n8682) );
  NAND2_X1 U10970 ( .A1(n6532), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U10971 ( .A1(n8684), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8685) );
  AND2_X1 U10972 ( .A1(n8702), .A2(n8685), .ZN(n14374) );
  OR2_X1 U10973 ( .A1(n6537), .A2(n14374), .ZN(n8690) );
  INV_X1 U10974 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n8686) );
  OR2_X1 U10975 ( .A1(n11767), .A2(n8686), .ZN(n8689) );
  INV_X1 U10976 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8687) );
  OR2_X1 U10977 ( .A1(n6518), .A2(n8687), .ZN(n8688) );
  NAND4_X1 U10978 ( .A1(n8691), .A2(n8690), .A3(n8689), .A4(n8688), .ZN(n12076) );
  INV_X1 U10979 ( .A(n12076), .ZN(n11318) );
  NAND2_X1 U10980 ( .A1(n11318), .A2(n14378), .ZN(n8692) );
  XNOR2_X1 U10981 ( .A(n8694), .B(n8693), .ZN(n9163) );
  NAND2_X1 U10982 ( .A1(n9163), .A2(n11774), .ZN(n8701) );
  OAI21_X1 U10983 ( .B1(n8695), .B2(P3_IR_REG_11__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8696) );
  MUX2_X1 U10984 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8696), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8699) );
  INV_X1 U10985 ( .A(n8697), .ZN(n8698) );
  NAND2_X1 U10986 ( .A1(n8699), .A2(n8698), .ZN(n12216) );
  AOI22_X1 U10987 ( .A1(n8809), .A2(n15171), .B1(n8808), .B2(n12216), .ZN(
        n8700) );
  NAND2_X1 U10988 ( .A1(n8701), .A2(n8700), .ZN(n14393) );
  NAND2_X1 U10989 ( .A1(n6533), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8706) );
  INV_X1 U10990 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14398) );
  OR2_X1 U10991 ( .A1(n8563), .A2(n14398), .ZN(n8705) );
  NOR2_X1 U10992 ( .A1(n8714), .A2(n7551), .ZN(n11324) );
  OR2_X1 U10993 ( .A1(n6538), .A2(n11324), .ZN(n8704) );
  INV_X1 U10994 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11325) );
  OR2_X1 U10995 ( .A1(n11767), .A2(n11325), .ZN(n8703) );
  NAND4_X1 U10996 ( .A1(n8706), .A2(n8705), .A3(n8704), .A4(n8703), .ZN(n14372) );
  NAND2_X1 U10997 ( .A1(n14393), .A2(n14372), .ZN(n11688) );
  INV_X1 U10998 ( .A(n14372), .ZN(n11237) );
  OR2_X1 U10999 ( .A1(n14393), .A2(n11237), .ZN(n8708) );
  XNOR2_X1 U11000 ( .A(n8709), .B(n9822), .ZN(n9259) );
  NAND2_X1 U11001 ( .A1(n9259), .A2(n11774), .ZN(n8712) );
  OR2_X1 U11002 ( .A1(n8697), .A2(n8429), .ZN(n8710) );
  XNOR2_X1 U11003 ( .A(n8710), .B(P3_IR_REG_13__SCAN_IN), .ZN(n14882) );
  AOI22_X1 U11004 ( .A1(n8809), .A2(SI_13_), .B1(n8808), .B2(n14882), .ZN(
        n8711) );
  NAND2_X1 U11005 ( .A1(n8712), .A2(n8711), .ZN(n14366) );
  NAND2_X1 U11006 ( .A1(n8913), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8721) );
  OR2_X1 U11007 ( .A1(n8714), .A2(n8713), .ZN(n8715) );
  AND2_X1 U11008 ( .A1(n8715), .A2(n8731), .ZN(n14362) );
  OR2_X1 U11009 ( .A1(n6538), .A2(n14362), .ZN(n8720) );
  INV_X1 U11010 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8716) );
  OR2_X1 U11011 ( .A1(n11767), .A2(n8716), .ZN(n8719) );
  INV_X1 U11012 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n8717) );
  OR2_X1 U11013 ( .A1(n8874), .A2(n8717), .ZN(n8718) );
  NAND4_X1 U11014 ( .A1(n8721), .A2(n8720), .A3(n8719), .A4(n8718), .ZN(n12201) );
  OR2_X1 U11015 ( .A1(n14366), .A2(n12201), .ZN(n8722) );
  NAND2_X1 U11016 ( .A1(n14366), .A2(n12201), .ZN(n8723) );
  NAND2_X1 U11017 ( .A1(n8724), .A2(n8723), .ZN(n11429) );
  XNOR2_X1 U11018 ( .A(n10078), .B(P2_DATAO_REG_14__SCAN_IN), .ZN(n8725) );
  XNOR2_X1 U11019 ( .A(n8726), .B(n8725), .ZN(n9310) );
  NAND2_X1 U11020 ( .A1(n9310), .A2(n11774), .ZN(n8730) );
  NAND2_X1 U11021 ( .A1(n8727), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8728) );
  XNOR2_X1 U11022 ( .A(n8728), .B(P3_IR_REG_14__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U11023 ( .A1(n8809), .A2(SI_14_), .B1(n8808), .B2(n12231), .ZN(
        n8729) );
  NAND2_X1 U11024 ( .A1(n8730), .A2(n8729), .ZN(n12614) );
  NAND2_X1 U11025 ( .A1(n8913), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8736) );
  INV_X1 U11026 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n15078) );
  OR2_X1 U11027 ( .A1(n8874), .A2(n15078), .ZN(n8735) );
  NAND2_X1 U11028 ( .A1(n8731), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8732) );
  AND2_X1 U11029 ( .A1(n8763), .A2(n8732), .ZN(n11433) );
  OR2_X1 U11030 ( .A1(n6537), .A2(n11433), .ZN(n8734) );
  INV_X1 U11031 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12220) );
  OR2_X1 U11032 ( .A1(n11767), .A2(n12220), .ZN(n8733) );
  OR2_X1 U11033 ( .A1(n12614), .A2(n14337), .ZN(n11698) );
  NAND2_X1 U11034 ( .A1(n12614), .A2(n14337), .ZN(n11699) );
  NAND2_X1 U11035 ( .A1(n11698), .A2(n11699), .ZN(n11430) );
  NAND2_X1 U11036 ( .A1(n11429), .A2(n11430), .ZN(n8738) );
  INV_X1 U11037 ( .A(n14337), .ZN(n14360) );
  NAND2_X1 U11038 ( .A1(n12614), .A2(n14360), .ZN(n8737) );
  INV_X1 U11039 ( .A(n8739), .ZN(n8740) );
  XNOR2_X1 U11040 ( .A(n8741), .B(n8740), .ZN(n9521) );
  NAND2_X1 U11041 ( .A1(n9521), .A2(n11774), .ZN(n8745) );
  NAND2_X1 U11042 ( .A1(n8755), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8743) );
  INV_X1 U11043 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8742) );
  XNOR2_X1 U11044 ( .A(n8743), .B(n8742), .ZN(n12277) );
  INV_X1 U11045 ( .A(n12277), .ZN(n12268) );
  AOI22_X1 U11046 ( .A1(n8809), .A2(SI_15_), .B1(n8808), .B2(n12268), .ZN(
        n8744) );
  NAND2_X1 U11047 ( .A1(n8745), .A2(n8744), .ZN(n14342) );
  NAND2_X1 U11048 ( .A1(n6533), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8750) );
  XNOR2_X1 U11049 ( .A(n8763), .B(n8746), .ZN(n14348) );
  OR2_X1 U11050 ( .A1(n6538), .A2(n14348), .ZN(n8749) );
  INV_X1 U11051 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15185) );
  OR2_X1 U11052 ( .A1(n11767), .A2(n15185), .ZN(n8748) );
  INV_X1 U11053 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12610) );
  OR2_X1 U11054 ( .A1(n8563), .A2(n12610), .ZN(n8747) );
  NAND4_X1 U11055 ( .A1(n8750), .A2(n8749), .A3(n8748), .A4(n8747), .ZN(n12537) );
  OR2_X1 U11056 ( .A1(n14342), .A2(n12537), .ZN(n8751) );
  INV_X1 U11057 ( .A(n12535), .ZN(n8772) );
  OAI21_X1 U11058 ( .B1(n8754), .B2(n8753), .A(n8752), .ZN(n9582) );
  OR2_X1 U11059 ( .A1(n9582), .A2(n6527), .ZN(n8762) );
  NOR2_X2 U11060 ( .A1(n8755), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8759) );
  INV_X1 U11061 ( .A(n8759), .ZN(n8756) );
  NAND2_X1 U11062 ( .A1(n8756), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8757) );
  MUX2_X1 U11063 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8757), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8760) );
  INV_X1 U11064 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8758) );
  INV_X1 U11065 ( .A(n8778), .ZN(n8775) );
  AND2_X1 U11066 ( .A1(n8760), .A2(n8775), .ZN(n12281) );
  AOI22_X1 U11067 ( .A1(n8809), .A2(SI_16_), .B1(n8808), .B2(n12281), .ZN(
        n8761) );
  NAND2_X1 U11068 ( .A1(n6532), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8770) );
  OAI21_X1 U11069 ( .B1(n8763), .B2(P3_REG3_REG_15__SCAN_IN), .A(
        P3_REG3_REG_16__SCAN_IN), .ZN(n8764) );
  INV_X1 U11070 ( .A(n8764), .ZN(n8765) );
  OR2_X1 U11071 ( .A1(n8765), .A2(n8783), .ZN(n12545) );
  INV_X1 U11072 ( .A(n12545), .ZN(n8766) );
  OR2_X1 U11073 ( .A1(n6537), .A2(n8766), .ZN(n8769) );
  INV_X1 U11074 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12280) );
  OR2_X1 U11075 ( .A1(n11767), .A2(n12280), .ZN(n8768) );
  INV_X1 U11076 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12270) );
  OR2_X1 U11077 ( .A1(n6518), .A2(n12270), .ZN(n8767) );
  NAND4_X1 U11078 ( .A1(n8770), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n14332) );
  NAND2_X1 U11079 ( .A1(n12547), .A2(n14332), .ZN(n11709) );
  INV_X1 U11080 ( .A(n14332), .ZN(n12131) );
  NAND2_X1 U11081 ( .A1(n12663), .A2(n12131), .ZN(n11708) );
  INV_X1 U11082 ( .A(n12541), .ZN(n8771) );
  NAND2_X1 U11083 ( .A1(n8772), .A2(n8771), .ZN(n12521) );
  NAND2_X1 U11084 ( .A1(n12663), .A2(n14332), .ZN(n12522) );
  NAND2_X1 U11085 ( .A1(n12521), .A2(n12522), .ZN(n8789) );
  XNOR2_X1 U11086 ( .A(n10244), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n8773) );
  XNOR2_X1 U11087 ( .A(n8774), .B(n8773), .ZN(n9775) );
  NAND2_X1 U11088 ( .A1(n9775), .A2(n11774), .ZN(n8781) );
  NAND2_X1 U11089 ( .A1(n8775), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8776) );
  MUX2_X1 U11090 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8776), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8779) );
  INV_X1 U11091 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U11092 ( .A1(n8779), .A2(n8805), .ZN(n12323) );
  INV_X1 U11093 ( .A(n12323), .ZN(n12310) );
  AOI22_X1 U11094 ( .A1(n8809), .A2(SI_17_), .B1(n8808), .B2(n12310), .ZN(
        n8780) );
  NAND2_X1 U11095 ( .A1(n8913), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8788) );
  INV_X1 U11096 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n8782) );
  OR2_X1 U11097 ( .A1(n8874), .A2(n8782), .ZN(n8787) );
  NOR2_X1 U11098 ( .A1(n8783), .A2(n12129), .ZN(n8784) );
  OR2_X1 U11099 ( .A1(n8796), .A2(n8784), .ZN(n12133) );
  INV_X1 U11100 ( .A(n12133), .ZN(n12528) );
  OR2_X1 U11101 ( .A1(n6538), .A2(n12528), .ZN(n8786) );
  INV_X1 U11102 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12529) );
  OR2_X1 U11103 ( .A1(n11767), .A2(n12529), .ZN(n8785) );
  OR2_X1 U11104 ( .A1(n12659), .A2(n12020), .ZN(n11713) );
  NAND2_X1 U11105 ( .A1(n12659), .A2(n12020), .ZN(n11712) );
  NAND2_X1 U11106 ( .A1(n11713), .A2(n11712), .ZN(n11804) );
  NAND2_X1 U11107 ( .A1(n8789), .A2(n11804), .ZN(n12524) );
  NAND2_X1 U11108 ( .A1(n12659), .A2(n12538), .ZN(n8790) );
  XNOR2_X1 U11109 ( .A(n8791), .B(n6662), .ZN(n9926) );
  NAND2_X1 U11110 ( .A1(n9926), .A2(n11774), .ZN(n8794) );
  NAND2_X1 U11111 ( .A1(n8805), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8792) );
  XNOR2_X1 U11112 ( .A(n8792), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U11113 ( .A1(n8809), .A2(SI_18_), .B1(n8808), .B2(n12347), .ZN(
        n8793) );
  NAND2_X1 U11114 ( .A1(n8913), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8801) );
  INV_X1 U11115 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n8795) );
  OR2_X1 U11116 ( .A1(n8874), .A2(n8795), .ZN(n8800) );
  OR2_X1 U11117 ( .A1(n8796), .A2(n15188), .ZN(n8797) );
  AND2_X1 U11118 ( .A1(n8812), .A2(n8797), .ZN(n12512) );
  OR2_X1 U11119 ( .A1(n6538), .A2(n12512), .ZN(n8799) );
  INV_X1 U11120 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12513) );
  OR2_X1 U11121 ( .A1(n11767), .A2(n12513), .ZN(n8798) );
  NAND2_X1 U11122 ( .A1(n12511), .A2(n12494), .ZN(n11719) );
  INV_X1 U11123 ( .A(n12494), .ZN(n12525) );
  INV_X1 U11124 ( .A(n8802), .ZN(n8803) );
  XNOR2_X1 U11125 ( .A(n8804), .B(n8803), .ZN(n9931) );
  NAND2_X1 U11126 ( .A1(n9931), .A2(n11774), .ZN(n8811) );
  INV_X1 U11127 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8806) );
  AOI22_X1 U11128 ( .A1(n8809), .A2(n9930), .B1(n8808), .B2(n6525), .ZN(n8810)
         );
  NAND2_X1 U11129 ( .A1(n8812), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U11130 ( .A1(n8824), .A2(n8813), .ZN(n12086) );
  NAND2_X1 U11131 ( .A1(n8897), .A2(n12086), .ZN(n8818) );
  INV_X1 U11132 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12591) );
  OR2_X1 U11133 ( .A1(n8563), .A2(n12591), .ZN(n8817) );
  INV_X1 U11134 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12652) );
  OR2_X1 U11135 ( .A1(n8814), .A2(n12652), .ZN(n8816) );
  INV_X1 U11136 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12500) );
  OR2_X1 U11137 ( .A1(n11767), .A2(n12500), .ZN(n8815) );
  NAND4_X1 U11138 ( .A1(n8818), .A2(n8817), .A3(n8816), .A4(n8815), .ZN(n12509) );
  NAND2_X1 U11139 ( .A1(n12655), .A2(n12509), .ZN(n11725) );
  NAND2_X1 U11140 ( .A1(n11724), .A2(n11725), .ZN(n12503) );
  INV_X1 U11141 ( .A(n12509), .ZN(n12169) );
  OR2_X1 U11142 ( .A1(n12655), .A2(n12169), .ZN(n8819) );
  XNOR2_X1 U11143 ( .A(n8821), .B(n8820), .ZN(n10109) );
  NAND2_X1 U11144 ( .A1(n10109), .A2(n11774), .ZN(n8823) );
  OR2_X1 U11145 ( .A1(n6529), .A2(n10112), .ZN(n8822) );
  AND2_X1 U11146 ( .A1(n8824), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8825) );
  OR2_X1 U11147 ( .A1(n8825), .A2(n8844), .ZN(n12487) );
  NAND2_X1 U11148 ( .A1(n12487), .A2(n8897), .ZN(n8829) );
  NAND2_X1 U11149 ( .A1(n8913), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8828) );
  NAND2_X1 U11150 ( .A1(n6533), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U11151 ( .A1(n8527), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U11152 ( .A1(n12650), .A2(n12495), .ZN(n11625) );
  NAND2_X1 U11153 ( .A1(n11626), .A2(n11625), .ZN(n12483) );
  INV_X1 U11154 ( .A(n12495), .ZN(n12200) );
  NAND2_X1 U11155 ( .A1(n12650), .A2(n12200), .ZN(n8830) );
  INV_X1 U11156 ( .A(n8831), .ZN(n8832) );
  XNOR2_X1 U11157 ( .A(n8833), .B(n8832), .ZN(n10355) );
  NAND2_X1 U11158 ( .A1(n10355), .A2(n11774), .ZN(n8835) );
  INV_X1 U11159 ( .A(SI_21_), .ZN(n10356) );
  OR2_X1 U11160 ( .A1(n11775), .A2(n10356), .ZN(n8834) );
  INV_X1 U11161 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n8838) );
  INV_X1 U11162 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12109) );
  XNOR2_X1 U11163 ( .A(n8844), .B(n12109), .ZN(n12473) );
  NAND2_X1 U11164 ( .A1(n12473), .A2(n8897), .ZN(n8837) );
  AOI22_X1 U11165 ( .A1(n6532), .A2(P3_REG0_REG_21__SCAN_IN), .B1(n8913), .B2(
        P3_REG1_REG_21__SCAN_IN), .ZN(n8836) );
  OAI211_X1 U11166 ( .C1(n11767), .C2(n8838), .A(n8837), .B(n8836), .ZN(n12480) );
  AND2_X1 U11167 ( .A1(n12112), .A2(n12480), .ZN(n11623) );
  OR2_X1 U11168 ( .A1(n12112), .A2(n12480), .ZN(n11622) );
  XNOR2_X1 U11169 ( .A(n8840), .B(n8839), .ZN(n10568) );
  NAND2_X1 U11170 ( .A1(n10568), .A2(n11774), .ZN(n8843) );
  OR2_X1 U11171 ( .A1(n6529), .A2(n8841), .ZN(n8842) );
  INV_X1 U11172 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8849) );
  INV_X1 U11173 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15266) );
  AOI21_X1 U11174 ( .B1(n8844), .B2(n12109), .A(n15266), .ZN(n8845) );
  OR2_X1 U11175 ( .A1(n8846), .A2(n8845), .ZN(n12463) );
  NAND2_X1 U11176 ( .A1(n12463), .A2(n8897), .ZN(n8848) );
  AOI22_X1 U11177 ( .A1(n6533), .A2(P3_REG0_REG_22__SCAN_IN), .B1(n8913), .B2(
        P3_REG1_REG_22__SCAN_IN), .ZN(n8847) );
  OAI211_X1 U11178 ( .C1(n11767), .C2(n8849), .A(n8848), .B(n8847), .ZN(n12444) );
  NAND2_X1 U11179 ( .A1(n12642), .A2(n12444), .ZN(n8850) );
  NAND2_X1 U11180 ( .A1(n12639), .A2(n12456), .ZN(n11615) );
  INV_X1 U11181 ( .A(n12639), .ZN(n12449) );
  NAND2_X1 U11182 ( .A1(n12449), .A2(n12162), .ZN(n8851) );
  NAND2_X1 U11183 ( .A1(n11615), .A2(n8851), .ZN(n12442) );
  NAND2_X1 U11184 ( .A1(n12635), .A2(n12445), .ZN(n11616) );
  INV_X1 U11185 ( .A(n12635), .ZN(n8852) );
  NAND2_X1 U11186 ( .A1(n8852), .A2(n12066), .ZN(n12418) );
  INV_X1 U11187 ( .A(n8853), .ZN(n8854) );
  XNOR2_X1 U11188 ( .A(n8855), .B(n8854), .ZN(n11367) );
  NAND2_X1 U11189 ( .A1(n11367), .A2(n11774), .ZN(n8857) );
  OR2_X1 U11190 ( .A1(n11775), .A2(n15275), .ZN(n8856) );
  NAND2_X1 U11191 ( .A1(n8858), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8859) );
  NAND2_X1 U11192 ( .A1(n8869), .A2(n8859), .ZN(n12423) );
  INV_X1 U11193 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U11194 ( .A1(n8913), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U11195 ( .A1(n6532), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8860) );
  OAI211_X1 U11196 ( .C1(n8862), .C2(n11767), .A(n8861), .B(n8860), .ZN(n8863)
         );
  AOI21_X1 U11197 ( .B1(n12423), .B2(n8897), .A(n8863), .ZN(n12145) );
  OR2_X1 U11198 ( .A1(n12041), .A2(n12145), .ZN(n11614) );
  NAND2_X1 U11199 ( .A1(n12041), .A2(n12145), .ZN(n12395) );
  NAND2_X1 U11200 ( .A1(n11614), .A2(n12395), .ZN(n12413) );
  INV_X1 U11201 ( .A(n8864), .ZN(n8865) );
  XNOR2_X1 U11202 ( .A(n8866), .B(n8865), .ZN(n12695) );
  NAND2_X1 U11203 ( .A1(n12695), .A2(n11774), .ZN(n8868) );
  AND2_X1 U11204 ( .A1(n8869), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8871) );
  OR2_X1 U11205 ( .A1(n8871), .A2(n8870), .ZN(n12407) );
  NAND2_X1 U11206 ( .A1(n12407), .A2(n8897), .ZN(n8877) );
  INV_X1 U11207 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n15165) );
  NAND2_X1 U11208 ( .A1(n8913), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U11209 ( .A1(n8527), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8872) );
  OAI211_X1 U11210 ( .C1(n8874), .C2(n15165), .A(n8873), .B(n8872), .ZN(n8875)
         );
  INV_X1 U11211 ( .A(n8875), .ZN(n8876) );
  OR2_X1 U11212 ( .A1(n12014), .A2(n12193), .ZN(n11753) );
  NAND2_X1 U11213 ( .A1(n12014), .A2(n12193), .ZN(n12371) );
  NAND2_X1 U11214 ( .A1(n8880), .A2(n8879), .ZN(n8881) );
  AOI22_X1 U11215 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n11988), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n11568), .ZN(n8890) );
  NAND2_X1 U11216 ( .A1(n11605), .A2(n11774), .ZN(n8883) );
  OR2_X1 U11217 ( .A1(n11775), .A2(n11606), .ZN(n8882) );
  INV_X1 U11218 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12098) );
  NOR2_X1 U11219 ( .A1(n8884), .A2(n12098), .ZN(n8885) );
  INV_X1 U11220 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U11221 ( .A1(n6532), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U11222 ( .A1(n8913), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8886) );
  OAI211_X1 U11223 ( .C1(n8888), .C2(n11767), .A(n8887), .B(n8886), .ZN(n8889)
         );
  NAND2_X1 U11224 ( .A1(n12102), .A2(n12387), .ZN(n11750) );
  NAND2_X1 U11225 ( .A1(n12367), .A2(n7553), .ZN(n8904) );
  AOI22_X1 U11226 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n14301), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n13570), .ZN(n8893) );
  INV_X1 U11227 ( .A(n8893), .ZN(n8894) );
  XNOR2_X1 U11228 ( .A(n11759), .B(n8894), .ZN(n12687) );
  NAND2_X1 U11229 ( .A1(n12687), .A2(n11774), .ZN(n8896) );
  OR2_X1 U11230 ( .A1(n6529), .A2(n12689), .ZN(n8895) );
  NAND2_X1 U11231 ( .A1(n8896), .A2(n8895), .ZN(n8989) );
  NAND2_X1 U11232 ( .A1(n14352), .A2(n8897), .ZN(n11770) );
  INV_X1 U11233 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U11234 ( .A1(n6533), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U11235 ( .A1(n8527), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8898) );
  OAI211_X1 U11236 ( .C1(n8900), .C2(n6518), .A(n8899), .B(n8898), .ZN(n8901)
         );
  INV_X1 U11237 ( .A(n8901), .ZN(n8902) );
  OR2_X1 U11238 ( .A1(n8989), .A2(n12370), .ZN(n11758) );
  NAND2_X1 U11239 ( .A1(n8989), .A2(n12370), .ZN(n11779) );
  NAND2_X1 U11240 ( .A1(n11758), .A2(n11779), .ZN(n11814) );
  INV_X1 U11241 ( .A(n11814), .ZN(n8903) );
  XNOR2_X1 U11242 ( .A(n8904), .B(n8903), .ZN(n8920) );
  NAND2_X1 U11243 ( .A1(n8907), .A2(n8905), .ZN(n8977) );
  NAND2_X1 U11244 ( .A1(n8977), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U11245 ( .A1(n11817), .A2(n11836), .ZN(n8980) );
  INV_X1 U11246 ( .A(n8907), .ZN(n8908) );
  NAND2_X1 U11247 ( .A1(n8908), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8909) );
  NAND2_X1 U11248 ( .A1(n6544), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8911) );
  INV_X1 U11249 ( .A(n10110), .ZN(n8997) );
  NAND2_X1 U11250 ( .A1(n11633), .A2(n8997), .ZN(n11829) );
  INV_X1 U11251 ( .A(n11833), .ZN(n9098) );
  CLKBUF_X3 U11252 ( .A(n8912), .Z(n12691) );
  INV_X1 U11253 ( .A(n12691), .ZN(n11834) );
  NAND2_X1 U11254 ( .A1(n9098), .A2(n11834), .ZN(n9081) );
  NAND2_X1 U11255 ( .A1(n9078), .A2(n9081), .ZN(n9993) );
  AND2_X2 U11256 ( .A1(n11836), .A2(n11633), .ZN(n11736) );
  INV_X1 U11257 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14405) );
  NAND2_X1 U11258 ( .A1(n8913), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U11259 ( .A1(n8527), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8914) );
  OAI211_X1 U11260 ( .C1(n8874), .C2(n14405), .A(n8915), .B(n8914), .ZN(n8916)
         );
  INV_X1 U11261 ( .A(n8916), .ZN(n8917) );
  AND2_X1 U11262 ( .A1(n11770), .A2(n8917), .ZN(n11782) );
  AND2_X1 U11263 ( .A1(n9098), .A2(P3_B_REG_SCAN_IN), .ZN(n8918) );
  OR2_X1 U11264 ( .A1(n14930), .A2(n8918), .ZN(n14349) );
  OAI22_X1 U11265 ( .A1(n12387), .A2(n14932), .B1(n11782), .B2(n14349), .ZN(
        n8919) );
  INV_X1 U11266 ( .A(n10255), .ZN(n9894) );
  NAND2_X1 U11267 ( .A1(n8922), .A2(n11629), .ZN(n9987) );
  NAND2_X1 U11268 ( .A1(n9987), .A2(n8923), .ZN(n14923) );
  NAND2_X1 U11269 ( .A1(n14923), .A2(n14922), .ZN(n8925) );
  NAND2_X1 U11270 ( .A1(n8925), .A2(n11636), .ZN(n10420) );
  INV_X1 U11271 ( .A(n10421), .ZN(n11788) );
  NAND2_X1 U11272 ( .A1(n10420), .A2(n11788), .ZN(n8926) );
  NAND2_X1 U11273 ( .A1(n8926), .A2(n11641), .ZN(n14905) );
  NAND2_X1 U11274 ( .A1(n14905), .A2(n14908), .ZN(n8928) );
  NAND2_X1 U11275 ( .A1(n8928), .A2(n11650), .ZN(n10432) );
  NAND2_X1 U11276 ( .A1(n10432), .A2(n11793), .ZN(n8929) );
  OR2_X1 U11277 ( .A1(n14910), .A2(n11655), .ZN(n11651) );
  NAND2_X1 U11278 ( .A1(n8929), .A2(n11651), .ZN(n10907) );
  OR2_X1 U11279 ( .A1(n12204), .A2(n14994), .ZN(n11661) );
  AND2_X1 U11280 ( .A1(n11660), .A2(n11661), .ZN(n8931) );
  INV_X1 U11281 ( .A(n11661), .ZN(n8930) );
  XNOR2_X1 U11282 ( .A(n12203), .B(n11038), .ZN(n11789) );
  INV_X1 U11283 ( .A(n11038), .ZN(n11667) );
  OR2_X1 U11284 ( .A1(n12203), .A2(n11667), .ZN(n11669) );
  INV_X1 U11285 ( .A(n11673), .ZN(n8932) );
  NAND2_X1 U11286 ( .A1(n14378), .A2(n12076), .ZN(n11686) );
  NAND2_X1 U11287 ( .A1(n11682), .A2(n11686), .ZN(n14376) );
  NAND2_X1 U11288 ( .A1(n11323), .A2(n11799), .ZN(n11322) );
  AND2_X1 U11289 ( .A1(n14366), .A2(n11432), .ZN(n11690) );
  OR2_X1 U11290 ( .A1(n14366), .A2(n11432), .ZN(n11693) );
  OR2_X1 U11291 ( .A1(n14342), .A2(n11490), .ZN(n11702) );
  NAND2_X1 U11292 ( .A1(n14342), .A2(n11490), .ZN(n11707) );
  NAND2_X1 U11293 ( .A1(n8934), .A2(n11707), .ZN(n12542) );
  NAND2_X1 U11294 ( .A1(n12542), .A2(n12541), .ZN(n12544) );
  NAND2_X1 U11295 ( .A1(n12544), .A2(n11708), .ZN(n12532) );
  NAND2_X1 U11296 ( .A1(n12516), .A2(n11714), .ZN(n12504) );
  INV_X1 U11297 ( .A(n11725), .ZN(n8935) );
  INV_X1 U11298 ( .A(n12484), .ZN(n8937) );
  NAND2_X1 U11299 ( .A1(n8937), .A2(n8936), .ZN(n12486) );
  INV_X1 U11300 ( .A(n12480), .ZN(n12458) );
  NOR2_X1 U11301 ( .A1(n12112), .A2(n12458), .ZN(n8938) );
  INV_X1 U11302 ( .A(n12444), .ZN(n12470) );
  AND2_X1 U11303 ( .A1(n12642), .A2(n12470), .ZN(n11619) );
  INV_X1 U11304 ( .A(n12442), .ZN(n11733) );
  INV_X1 U11305 ( .A(n11615), .ZN(n8939) );
  AOI21_X2 U11306 ( .B1(n12440), .B2(n11733), .A(n8939), .ZN(n12431) );
  INV_X1 U11307 ( .A(n12413), .ZN(n12421) );
  AND2_X1 U11308 ( .A1(n12430), .A2(n12421), .ZN(n8940) );
  NAND2_X1 U11309 ( .A1(n12047), .A2(n12386), .ZN(n11612) );
  NAND2_X1 U11310 ( .A1(n11613), .A2(n11612), .ZN(n12396) );
  INV_X1 U11311 ( .A(n12395), .ZN(n8941) );
  NOR2_X1 U11312 ( .A1(n12396), .A2(n8941), .ZN(n8942) );
  NAND2_X1 U11313 ( .A1(n11750), .A2(n12371), .ZN(n11748) );
  XOR2_X1 U11314 ( .A(n11814), .B(n11824), .Z(n11570) );
  NAND2_X1 U11315 ( .A1(n6525), .A2(n10418), .ZN(n8945) );
  NAND2_X1 U11316 ( .A1(n10418), .A2(n10110), .ZN(n8943) );
  XNOR2_X1 U11317 ( .A(n11836), .B(n8943), .ZN(n8944) );
  NAND2_X1 U11318 ( .A1(n8945), .A2(n8944), .ZN(n9788) );
  NAND2_X1 U11319 ( .A1(n6525), .A2(n10110), .ZN(n11611) );
  INV_X1 U11320 ( .A(n11611), .ZN(n8946) );
  INV_X1 U11321 ( .A(n11836), .ZN(n8998) );
  NAND3_X1 U11322 ( .A1(n9788), .A2(n8946), .A3(n15013), .ZN(n8947) );
  NAND2_X1 U11323 ( .A1(n11817), .A2(n10110), .ZN(n14951) );
  OR2_X1 U11324 ( .A1(n14951), .A2(n11836), .ZN(n15006) );
  NAND2_X1 U11325 ( .A1(n8949), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8950) );
  MUX2_X1 U11326 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8950), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8952) );
  INV_X1 U11327 ( .A(n8489), .ZN(n8951) );
  INV_X1 U11328 ( .A(n6516), .ZN(n8956) );
  NAND2_X1 U11329 ( .A1(n8956), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8953) );
  MUX2_X1 U11330 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8953), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8954) );
  NAND2_X1 U11331 ( .A1(n8954), .A2(n8949), .ZN(n11369) );
  NAND2_X1 U11332 ( .A1(n6576), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8955) );
  MUX2_X1 U11333 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8955), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8957) );
  NAND2_X1 U11334 ( .A1(n8957), .A2(n8956), .ZN(n11332) );
  XNOR2_X1 U11335 ( .A(n11332), .B(P3_B_REG_SCAN_IN), .ZN(n8958) );
  NAND2_X1 U11336 ( .A1(n11369), .A2(n8958), .ZN(n8959) );
  INV_X1 U11337 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8960) );
  NAND2_X1 U11338 ( .A1(n9178), .A2(n8960), .ZN(n8962) );
  NAND2_X1 U11339 ( .A1(n12699), .A2(n11332), .ZN(n8961) );
  INV_X1 U11340 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U11341 ( .A1(n9178), .A2(n8963), .ZN(n8965) );
  NAND2_X1 U11342 ( .A1(n12699), .A2(n11369), .ZN(n8964) );
  NAND2_X1 U11343 ( .A1(n12674), .A2(n12672), .ZN(n8995) );
  NOR2_X1 U11344 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .ZN(
        n15032) );
  NOR4_X1 U11345 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n8968) );
  NOR4_X1 U11346 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n8967) );
  NOR4_X1 U11347 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n8966) );
  NAND4_X1 U11348 ( .A1(n15032), .A2(n8968), .A3(n8967), .A4(n8966), .ZN(n8974) );
  NOR4_X1 U11349 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8972) );
  NOR4_X1 U11350 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n8971) );
  NOR4_X1 U11351 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8970) );
  NOR4_X1 U11352 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8969) );
  NAND4_X1 U11353 ( .A1(n8972), .A2(n8971), .A3(n8970), .A4(n8969), .ZN(n8973)
         );
  OAI21_X1 U11354 ( .B1(n8974), .B2(n8973), .A(n9178), .ZN(n8992) );
  INV_X1 U11355 ( .A(n8992), .ZN(n8984) );
  NOR2_X1 U11356 ( .A1(n8995), .A2(n8984), .ZN(n9793) );
  NOR2_X1 U11357 ( .A1(n11611), .A2(n11755), .ZN(n9892) );
  NOR2_X1 U11358 ( .A1(n11369), .A2(n11332), .ZN(n8975) );
  NAND2_X1 U11359 ( .A1(n8976), .A2(n8975), .ZN(n9779) );
  OAI21_X1 U11360 ( .B1(n8977), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8978) );
  MUX2_X1 U11361 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8978), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8979) );
  NAND2_X1 U11362 ( .A1(n8979), .A2(n6576), .ZN(n9778) );
  NAND2_X1 U11363 ( .A1(n9892), .A2(n9794), .ZN(n11835) );
  OR2_X1 U11364 ( .A1(n11633), .A2(n10110), .ZN(n11819) );
  NOR2_X1 U11365 ( .A1(n8980), .A2(n11819), .ZN(n9789) );
  NAND2_X1 U11366 ( .A1(n9789), .A2(n9794), .ZN(n8981) );
  NAND2_X1 U11367 ( .A1(n11835), .A2(n8981), .ZN(n8982) );
  NAND2_X1 U11368 ( .A1(n9793), .A2(n8982), .ZN(n8986) );
  INV_X1 U11369 ( .A(n12674), .ZN(n8983) );
  NAND2_X1 U11370 ( .A1(n8983), .A2(n9000), .ZN(n8993) );
  NOR2_X1 U11371 ( .A1(n8993), .A2(n8984), .ZN(n9798) );
  NAND3_X1 U11372 ( .A1(n9798), .A2(n9794), .A3(n9788), .ZN(n8985) );
  NAND2_X1 U11373 ( .A1(n15018), .A2(n8987), .ZN(n8988) );
  INV_X1 U11374 ( .A(n8989), .ZN(n11572) );
  OR2_X1 U11375 ( .A1(n15018), .A2(n15013), .ZN(n12669) );
  NAND2_X1 U11376 ( .A1(n8990), .A2(n7534), .ZN(P3_U3456) );
  AND2_X1 U11377 ( .A1(n8992), .A2(n9794), .ZN(n8994) );
  NAND2_X1 U11378 ( .A1(n11611), .A2(n11736), .ZN(n9780) );
  NAND2_X1 U11379 ( .A1(n8996), .A2(n11755), .ZN(n10246) );
  AND2_X1 U11380 ( .A1(n9780), .A2(n10246), .ZN(n10248) );
  OAI22_X1 U11381 ( .A1(n11817), .A2(n8998), .B1(n8997), .B2(n15013), .ZN(
        n8999) );
  AOI21_X1 U11382 ( .B1(n8999), .B2(n11611), .A(n11736), .ZN(n9001) );
  MUX2_X1 U11383 ( .A(n10248), .B(n9001), .S(n9000), .Z(n9002) );
  OR2_X1 U11384 ( .A1(n15031), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U11385 ( .A1(n15031), .A2(n14980), .ZN(n12612) );
  NAND2_X1 U11386 ( .A1(n9004), .A2(n7533), .ZN(P3_U3488) );
  AND2_X2 U11387 ( .A1(n9110), .A2(n9005), .ZN(n9146) );
  NOR2_X1 U11388 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n9012) );
  NAND4_X1 U11389 ( .A1(n9330), .A2(n9012), .A3(n9336), .A4(n10079), .ZN(n9214) );
  NAND2_X1 U11390 ( .A1(n9329), .A2(n9217), .ZN(n9013) );
  NAND2_X1 U11391 ( .A1(n9021), .A2(n9018), .ZN(n9024) );
  NAND2_X1 U11392 ( .A1(n9024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9014) );
  MUX2_X1 U11393 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9014), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9020) );
  NAND2_X1 U11394 ( .A1(n9020), .A2(n9026), .ZN(n11370) );
  INV_X1 U11395 ( .A(n9021), .ZN(n9022) );
  NAND2_X1 U11396 ( .A1(n9022), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9023) );
  MUX2_X1 U11397 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9023), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9025) );
  NAND2_X1 U11398 ( .A1(n9025), .A2(n9024), .ZN(n11333) );
  NAND2_X1 U11399 ( .A1(n9026), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9027) );
  OR2_X1 U11400 ( .A1(n11333), .A2(n11453), .ZN(n9028) );
  NAND2_X1 U11401 ( .A1(n6575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9030) );
  XNOR2_X1 U11402 ( .A(n9030), .B(n9029), .ZN(n11357) );
  INV_X1 U11403 ( .A(n9357), .ZN(n9031) );
  INV_X1 U11404 ( .A(n9175), .ZN(n9256) );
  OR2_X2 U11405 ( .A1(n9256), .A2(n9595), .ZN(n13856) );
  INV_X1 U11406 ( .A(n9779), .ZN(n9032) );
  INV_X2 U11407 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  MUX2_X1 U11408 ( .A(n9034), .B(n9033), .S(n12691), .Z(n9036) );
  NAND2_X1 U11409 ( .A1(n9036), .A2(n9035), .ZN(n9731) );
  INV_X1 U11410 ( .A(n9036), .ZN(n9037) );
  NAND2_X1 U11411 ( .A1(n9037), .A2(n9677), .ZN(n9038) );
  NAND2_X1 U11412 ( .A1(n9731), .A2(n9038), .ZN(n9666) );
  INV_X1 U11413 ( .A(n9666), .ZN(n9039) );
  MUX2_X1 U11414 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n12691), .Z(n9683) );
  NOR2_X1 U11415 ( .A1(n9683), .A2(n9121), .ZN(n9665) );
  NAND2_X1 U11416 ( .A1(n9039), .A2(n9665), .ZN(n9732) );
  MUX2_X1 U11417 ( .A(n9086), .B(n9070), .S(n12691), .Z(n9040) );
  NAND2_X1 U11418 ( .A1(n9040), .A2(n9136), .ZN(n9043) );
  INV_X1 U11419 ( .A(n9040), .ZN(n9041) );
  INV_X1 U11420 ( .A(n9136), .ZN(n9726) );
  NAND2_X1 U11421 ( .A1(n9041), .A2(n9726), .ZN(n9042) );
  NAND2_X1 U11422 ( .A1(n9043), .A2(n9042), .ZN(n9730) );
  AOI21_X1 U11423 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(n9763) );
  INV_X1 U11424 ( .A(n9043), .ZN(n9762) );
  MUX2_X1 U11425 ( .A(n10428), .B(n9044), .S(n12691), .Z(n9045) );
  NAND2_X1 U11426 ( .A1(n9045), .A2(n9139), .ZN(n9825) );
  INV_X1 U11427 ( .A(n9045), .ZN(n9046) );
  NAND2_X1 U11428 ( .A1(n9046), .A2(n9774), .ZN(n9047) );
  OAI21_X1 U11429 ( .B1(n9763), .B2(n9762), .A(n7548), .ZN(n9826) );
  MUX2_X1 U11430 ( .A(n9048), .B(n9073), .S(n12691), .Z(n9049) );
  NAND2_X1 U11431 ( .A1(n9049), .A2(n9142), .ZN(n9052) );
  INV_X1 U11432 ( .A(n9049), .ZN(n9050) );
  NAND2_X1 U11433 ( .A1(n9050), .A2(n7060), .ZN(n9051) );
  NAND2_X1 U11434 ( .A1(n9052), .A2(n9051), .ZN(n9824) );
  AOI21_X1 U11435 ( .B1(n9826), .B2(n9825), .A(n9824), .ZN(n9828) );
  INV_X1 U11436 ( .A(n9052), .ZN(n9804) );
  MUX2_X1 U11437 ( .A(n10438), .B(n9053), .S(n12691), .Z(n9054) );
  NAND2_X1 U11438 ( .A1(n9054), .A2(n9091), .ZN(n9063) );
  INV_X1 U11439 ( .A(n9054), .ZN(n9055) );
  NAND2_X1 U11440 ( .A1(n9055), .A2(n9813), .ZN(n9056) );
  OAI21_X1 U11441 ( .B1(n9828), .B2(n9804), .A(n7547), .ZN(n9803) );
  MUX2_X1 U11442 ( .A(n10915), .B(n9057), .S(n12691), .Z(n9059) );
  NAND2_X1 U11443 ( .A1(n9059), .A2(n9058), .ZN(n10033) );
  INV_X1 U11444 ( .A(n9059), .ZN(n9060) );
  NAND2_X1 U11445 ( .A1(n9060), .A2(n10045), .ZN(n9061) );
  NAND2_X1 U11446 ( .A1(n10033), .A2(n9061), .ZN(n9062) );
  AOI21_X1 U11447 ( .B1(n9803), .B2(n9063), .A(n9062), .ZN(n10041) );
  INV_X1 U11448 ( .A(n10041), .ZN(n9065) );
  NAND3_X1 U11449 ( .A1(n9803), .A2(n9063), .A3(n9062), .ZN(n9064) );
  AND2_X1 U11450 ( .A1(P3_U3897), .A2(n11833), .ZN(n14893) );
  INV_X1 U11451 ( .A(n14893), .ZN(n14873) );
  AOI21_X1 U11452 ( .B1(n9065), .B2(n9064), .A(n14873), .ZN(n9108) );
  NAND2_X1 U11453 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n9121), .ZN(n9068) );
  NAND2_X1 U11454 ( .A1(n9677), .A2(n9068), .ZN(n9067) );
  INV_X1 U11455 ( .A(n9068), .ZN(n9682) );
  NAND2_X1 U11456 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9682), .ZN(n9066) );
  NAND2_X1 U11457 ( .A1(n9067), .A2(n9066), .ZN(n9669) );
  NAND2_X1 U11458 ( .A1(n9669), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9668) );
  OR2_X1 U11459 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9068), .ZN(n9069) );
  NAND2_X1 U11460 ( .A1(n9668), .A2(n9069), .ZN(n9721) );
  OAI21_X1 U11461 ( .B1(n9136), .B2(n9070), .A(n9720), .ZN(n9071) );
  NAND2_X1 U11462 ( .A1(n9071), .A2(n9774), .ZN(n9072) );
  INV_X1 U11463 ( .A(n9072), .ZN(n9830) );
  XNOR2_X1 U11464 ( .A(n9142), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n9829) );
  NAND2_X1 U11465 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n10045), .ZN(n9074) );
  OAI21_X1 U11466 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n10045), .A(n9074), .ZN(
        n9075) );
  NOR2_X1 U11467 ( .A1(n9076), .A2(n9075), .ZN(n10031) );
  AOI21_X1 U11468 ( .B1(n9076), .B2(n9075), .A(n10031), .ZN(n9080) );
  NAND2_X1 U11469 ( .A1(n11736), .A2(n9778), .ZN(n9077) );
  OR2_X1 U11470 ( .A1(n9778), .A2(P3_U3151), .ZN(n11839) );
  INV_X1 U11471 ( .A(n11839), .ZN(n9079) );
  OR2_X1 U11472 ( .A1(n9794), .A2(n9079), .ZN(n9100) );
  NOR2_X1 U11473 ( .A1(n9080), .A2(n14897), .ZN(n9107) );
  INV_X1 U11474 ( .A(n9081), .ZN(n9082) );
  NAND2_X1 U11475 ( .A1(n9083), .A2(n9082), .ZN(n14903) );
  XNOR2_X1 U11476 ( .A(n9136), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n9719) );
  INV_X1 U11477 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n15155) );
  NOR2_X1 U11478 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n15155), .ZN(n9678) );
  NAND2_X1 U11479 ( .A1(n9084), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9085) );
  OR2_X1 U11480 ( .A1(n9136), .A2(n9086), .ZN(n9087) );
  NAND2_X1 U11481 ( .A1(n9717), .A2(n9087), .ZN(n9088) );
  NAND2_X1 U11482 ( .A1(n9088), .A2(n9774), .ZN(n9835) );
  OR2_X1 U11483 ( .A1(n9088), .A2(n9774), .ZN(n9089) );
  AND2_X1 U11484 ( .A1(n9835), .A2(n9089), .ZN(n9766) );
  XNOR2_X1 U11485 ( .A(n9142), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U11486 ( .A1(n7060), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9090) );
  XNOR2_X1 U11487 ( .A(n9092), .B(n9091), .ZN(n9808) );
  NAND2_X1 U11488 ( .A1(n9092), .A2(n9813), .ZN(n9093) );
  NAND2_X1 U11489 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n10045), .ZN(n9094) );
  OAI21_X1 U11490 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10045), .A(n9094), .ZN(
        n9095) );
  AOI21_X1 U11491 ( .B1(n9096), .B2(n9095), .A(n10044), .ZN(n9097) );
  NOR2_X1 U11492 ( .A1(n14903), .A2(n9097), .ZN(n9106) );
  INV_X1 U11493 ( .A(P3_U3897), .ZN(n12199) );
  MUX2_X1 U11494 ( .A(n9099), .B(n12199), .S(n9098), .Z(n14885) );
  INV_X1 U11495 ( .A(n9100), .ZN(n9101) );
  NOR2_X1 U11496 ( .A1(n9102), .A2(n9101), .ZN(n14862) );
  INV_X1 U11497 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n9103) );
  NOR2_X1 U11498 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9103), .ZN(n12179) );
  AOI21_X1 U11499 ( .B1(n14862), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n12179), .ZN(
        n9104) );
  OAI21_X1 U11500 ( .B1(n14885), .B2(n10045), .A(n9104), .ZN(n9105) );
  OR4_X1 U11501 ( .A1(n9108), .A2(n9107), .A3(n9106), .A4(n9105), .ZN(P3_U3188) );
  NAND2_X1 U11502 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9109) );
  MUX2_X1 U11503 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9109), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9112) );
  INV_X1 U11504 ( .A(n9110), .ZN(n9111) );
  NAND2_X1 U11505 ( .A1(n9112), .A2(n9111), .ZN(n13082) );
  NAND2_X1 U11506 ( .A1(n9343), .A2(P2_U3088), .ZN(n13574) );
  AND2_X1 U11507 ( .A1(n9345), .A2(P2_U3088), .ZN(n13572) );
  INV_X2 U11508 ( .A(n13572), .ZN(n13580) );
  OAI222_X1 U11509 ( .A1(P2_U3088), .A2(n13082), .B1(n13574), .B2(n9344), .C1(
        n9347), .C2(n13580), .ZN(P2_U3326) );
  NOR2_X1 U11510 ( .A1(n9343), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14296) );
  INV_X2 U11511 ( .A(n14296), .ZN(n14305) );
  AND2_X1 U11512 ( .A1(n9343), .A2(P1_U3086), .ZN(n9759) );
  INV_X2 U11513 ( .A(n9759), .ZN(n14302) );
  OAI222_X1 U11514 ( .A1(P1_U3086), .A2(n13884), .B1(n14305), .B2(n9527), .C1(
        n9113), .C2(n14302), .ZN(P1_U3353) );
  NAND2_X1 U11515 ( .A1(n9345), .A2(P3_U3151), .ZN(n12694) );
  NAND2_X2 U11516 ( .A1(n9343), .A2(P3_U3151), .ZN(n12698) );
  OAI222_X1 U11517 ( .A1(n12694), .A2(n9115), .B1(n12698), .B2(n9114), .C1(
        P3_U3151), .C2(n9677), .ZN(P3_U3294) );
  INV_X1 U11518 ( .A(SI_5_), .ZN(n9117) );
  OAI222_X1 U11519 ( .A1(P3_U3151), .A2(n9813), .B1(n12698), .B2(n9117), .C1(
        n12694), .C2(n9116), .ZN(P3_U3290) );
  OAI222_X1 U11520 ( .A1(P3_U3151), .A2(n10487), .B1(n12698), .B2(n15203), 
        .C1(n12694), .C2(n9118), .ZN(P3_U3287) );
  OAI222_X1 U11521 ( .A1(P3_U3151), .A2(n9121), .B1(n12694), .B2(n9120), .C1(
        n9119), .C2(n12698), .ZN(P3_U3295) );
  OAI222_X1 U11522 ( .A1(P1_U3086), .A2(n13867), .B1(n14305), .B2(n9344), .C1(
        n7710), .C2(n14302), .ZN(P1_U3354) );
  INV_X1 U11523 ( .A(n9640), .ZN(n9124) );
  INV_X1 U11524 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n10301) );
  OR2_X1 U11525 ( .A1(n9146), .A2(n10301), .ZN(n9122) );
  XNOR2_X1 U11526 ( .A(n9122), .B(n9145), .ZN(n9643) );
  OAI222_X1 U11527 ( .A1(n13580), .A2(n9641), .B1(n13574), .B2(n9124), .C1(
        P2_U3088), .C2(n9643), .ZN(P2_U3324) );
  INV_X1 U11528 ( .A(n13896), .ZN(n9123) );
  OAI222_X1 U11529 ( .A1(n14302), .A2(n9125), .B1(n14305), .B2(n9124), .C1(
        n9123), .C2(P1_U3086), .ZN(P1_U3352) );
  NOR2_X1 U11530 ( .A1(n9110), .A2(n10301), .ZN(n9126) );
  MUX2_X1 U11531 ( .A(n10301), .B(n9126), .S(P2_IR_REG_2__SCAN_IN), .Z(n9127)
         );
  INV_X1 U11532 ( .A(n9127), .ZN(n9129) );
  INV_X1 U11533 ( .A(n9146), .ZN(n9128) );
  NAND2_X1 U11534 ( .A1(n9129), .A2(n9128), .ZN(n14666) );
  INV_X1 U11535 ( .A(n13574), .ZN(n13564) );
  INV_X1 U11536 ( .A(n13564), .ZN(n13578) );
  OAI222_X1 U11537 ( .A1(P2_U3088), .A2(n14666), .B1(n13578), .B2(n9527), .C1(
        n9526), .C2(n13580), .ZN(P2_U3325) );
  OAI222_X1 U11538 ( .A1(n12694), .A2(n9131), .B1(n12698), .B2(n9130), .C1(
        P3_U3151), .C2(n10045), .ZN(P3_U3289) );
  INV_X1 U11539 ( .A(n12694), .ZN(n12680) );
  INV_X1 U11540 ( .A(n12698), .ZN(n9258) );
  AOI222_X1 U11541 ( .A1(n9132), .A2(n12680), .B1(SI_9_), .B2(n9258), .C1(
        n10708), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9133) );
  INV_X1 U11542 ( .A(n9133), .ZN(P3_U3286) );
  AOI222_X1 U11543 ( .A1(n9134), .A2(n12680), .B1(SI_7_), .B2(n9258), .C1(
        n10147), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9135) );
  INV_X1 U11544 ( .A(n9135), .ZN(P3_U3288) );
  AOI222_X1 U11545 ( .A1(n9137), .A2(n12680), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9136), .C1(SI_2_), .C2(n9258), .ZN(n9138) );
  INV_X1 U11546 ( .A(n9138), .ZN(P3_U3293) );
  AOI222_X1 U11547 ( .A1(n9140), .A2(n12680), .B1(n9139), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_3_), .C2(n9258), .ZN(n9141) );
  INV_X1 U11548 ( .A(n9141), .ZN(P3_U3292) );
  AOI222_X1 U11549 ( .A1(n9143), .A2(n12680), .B1(SI_4_), .B2(n9258), .C1(
        n9142), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9144) );
  INV_X1 U11550 ( .A(n9144), .ZN(P3_U3291) );
  INV_X1 U11551 ( .A(n9741), .ZN(n9149) );
  NAND2_X1 U11552 ( .A1(n9146), .A2(n9145), .ZN(n9154) );
  NAND2_X1 U11553 ( .A1(n9154), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9147) );
  XNOR2_X1 U11554 ( .A(n9147), .B(P2_IR_REG_4__SCAN_IN), .ZN(n13098) );
  INV_X1 U11555 ( .A(n13098), .ZN(n13092) );
  OAI222_X1 U11556 ( .A1(n13580), .A2(n9148), .B1(n13574), .B2(n9149), .C1(
        P2_U3088), .C2(n13092), .ZN(P2_U3323) );
  OAI222_X1 U11557 ( .A1(n14302), .A2(n9150), .B1(n14305), .B2(n9149), .C1(
        n13914), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U11558 ( .A(SI_10_), .ZN(n9152) );
  OAI222_X1 U11559 ( .A1(P3_U3151), .A2(n11080), .B1(n12698), .B2(n9152), .C1(
        n12694), .C2(n9151), .ZN(P3_U3285) );
  INV_X1 U11560 ( .A(n9566), .ZN(n9423) );
  OAI222_X1 U11561 ( .A1(P1_U3086), .A2(n9423), .B1(n14305), .B2(n9845), .C1(
        n9153), .C2(n14302), .ZN(P1_U3350) );
  NAND2_X1 U11562 ( .A1(n9157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9155) );
  XNOR2_X1 U11563 ( .A(n9155), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9846) );
  INV_X1 U11564 ( .A(n9846), .ZN(n9255) );
  OAI222_X1 U11565 ( .A1(P2_U3088), .A2(n9255), .B1(n13578), .B2(n9845), .C1(
        n9156), .C2(n13580), .ZN(P2_U3322) );
  OR2_X1 U11566 ( .A1(n9165), .A2(n10301), .ZN(n9158) );
  XNOR2_X1 U11567 ( .A(n9158), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14690) );
  AOI22_X1 U11568 ( .A1(n14690), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n13572), .ZN(n9159) );
  OAI21_X1 U11569 ( .B1(n9967), .B2(n13574), .A(n9159), .ZN(P2_U3321) );
  OAI222_X1 U11570 ( .A1(P3_U3151), .A2(n14866), .B1(n12698), .B2(n9161), .C1(
        n12694), .C2(n9160), .ZN(P3_U3284) );
  INV_X1 U11571 ( .A(n13929), .ZN(n9400) );
  OAI222_X1 U11572 ( .A1(P1_U3086), .A2(n9400), .B1(n14305), .B2(n9967), .C1(
        n9162), .C2(n14302), .ZN(P1_U3349) );
  OAI222_X1 U11573 ( .A1(n12216), .A2(P3_U3151), .B1(n12694), .B2(n9163), .C1(
        n12698), .C2(n15171), .ZN(P3_U3283) );
  NAND2_X1 U11574 ( .A1(n9165), .A2(n9164), .ZN(n9207) );
  NAND2_X1 U11575 ( .A1(n9207), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9166) );
  XNOR2_X1 U11576 ( .A(n9166), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10061) );
  INV_X1 U11577 ( .A(n10061), .ZN(n9168) );
  OAI222_X1 U11578 ( .A1(P2_U3088), .A2(n9168), .B1(n13574), .B2(n10060), .C1(
        n9167), .C2(n13580), .ZN(P2_U3320) );
  INV_X1 U11579 ( .A(n9546), .ZN(n9558) );
  OAI222_X1 U11580 ( .A1(P1_U3086), .A2(n9558), .B1(n14305), .B2(n10060), .C1(
        n9169), .C2(n14302), .ZN(P1_U3348) );
  NAND2_X1 U11581 ( .A1(n11372), .A2(P1_B_REG_SCAN_IN), .ZN(n9170) );
  MUX2_X1 U11582 ( .A(P1_B_REG_SCAN_IN), .B(n9170), .S(n11610), .Z(n9172) );
  INV_X1 U11583 ( .A(n11450), .ZN(n9171) );
  NAND2_X1 U11584 ( .A1(n9172), .A2(n9171), .ZN(n9508) );
  INV_X1 U11585 ( .A(n9604), .ZN(n9173) );
  NAND2_X1 U11586 ( .A1(n9508), .A2(n9173), .ZN(n14578) );
  INV_X1 U11587 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9176) );
  NAND2_X1 U11588 ( .A1(n11372), .A2(n11450), .ZN(n9509) );
  INV_X1 U11589 ( .A(n9509), .ZN(n9174) );
  AOI22_X1 U11590 ( .A1(n14578), .A2(n9176), .B1(n9175), .B2(n9174), .ZN(
        P1_U3446) );
  INV_X1 U11591 ( .A(n12673), .ZN(n9177) );
  NOR2_X1 U11592 ( .A1(n9178), .A2(n9177), .ZN(n9181) );
  INV_X1 U11593 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9179) );
  NOR2_X1 U11594 ( .A1(n9203), .A2(n9179), .ZN(P3_U3242) );
  INV_X1 U11595 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9180) );
  NOR2_X1 U11596 ( .A1(n9181), .A2(n9180), .ZN(P3_U3243) );
  INV_X1 U11597 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n15139) );
  NOR2_X1 U11598 ( .A1(n9181), .A2(n15139), .ZN(P3_U3245) );
  CLKBUF_X1 U11599 ( .A(n9181), .Z(n9203) );
  INV_X1 U11600 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9182) );
  NOR2_X1 U11601 ( .A1(n9203), .A2(n9182), .ZN(P3_U3246) );
  INV_X1 U11602 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n15257) );
  NOR2_X1 U11603 ( .A1(n9181), .A2(n15257), .ZN(P3_U3244) );
  INV_X1 U11604 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9183) );
  NOR2_X1 U11605 ( .A1(n9203), .A2(n9183), .ZN(P3_U3248) );
  INV_X1 U11606 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9184) );
  NOR2_X1 U11607 ( .A1(n9203), .A2(n9184), .ZN(P3_U3249) );
  INV_X1 U11608 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9185) );
  NOR2_X1 U11609 ( .A1(n9203), .A2(n9185), .ZN(P3_U3255) );
  INV_X1 U11610 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9186) );
  NOR2_X1 U11611 ( .A1(n9203), .A2(n9186), .ZN(P3_U3254) );
  INV_X1 U11612 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15079) );
  NOR2_X1 U11613 ( .A1(n9203), .A2(n15079), .ZN(P3_U3253) );
  INV_X1 U11614 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9187) );
  NOR2_X1 U11615 ( .A1(n9203), .A2(n9187), .ZN(P3_U3252) );
  INV_X1 U11616 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9188) );
  NOR2_X1 U11617 ( .A1(n9203), .A2(n9188), .ZN(P3_U3251) );
  INV_X1 U11618 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9189) );
  NOR2_X1 U11619 ( .A1(n9203), .A2(n9189), .ZN(P3_U3250) );
  INV_X1 U11620 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9190) );
  NOR2_X1 U11621 ( .A1(n9181), .A2(n9190), .ZN(P3_U3234) );
  INV_X1 U11622 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9191) );
  NOR2_X1 U11623 ( .A1(n9181), .A2(n9191), .ZN(P3_U3235) );
  INV_X1 U11624 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9192) );
  NOR2_X1 U11625 ( .A1(n9203), .A2(n9192), .ZN(P3_U3263) );
  INV_X1 U11626 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9193) );
  NOR2_X1 U11627 ( .A1(n9181), .A2(n9193), .ZN(P3_U3262) );
  INV_X1 U11628 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9194) );
  NOR2_X1 U11629 ( .A1(n9203), .A2(n9194), .ZN(P3_U3261) );
  INV_X1 U11630 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9195) );
  NOR2_X1 U11631 ( .A1(n9181), .A2(n9195), .ZN(P3_U3260) );
  INV_X1 U11632 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9196) );
  NOR2_X1 U11633 ( .A1(n9181), .A2(n9196), .ZN(P3_U3240) );
  INV_X1 U11634 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9197) );
  NOR2_X1 U11635 ( .A1(n9203), .A2(n9197), .ZN(P3_U3259) );
  INV_X1 U11636 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9198) );
  NOR2_X1 U11637 ( .A1(n9181), .A2(n9198), .ZN(P3_U3258) );
  INV_X1 U11638 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9199) );
  NOR2_X1 U11639 ( .A1(n9203), .A2(n9199), .ZN(P3_U3257) );
  INV_X1 U11640 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9200) );
  NOR2_X1 U11641 ( .A1(n9203), .A2(n9200), .ZN(P3_U3256) );
  INV_X1 U11642 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9201) );
  NOR2_X1 U11643 ( .A1(n9181), .A2(n9201), .ZN(P3_U3238) );
  INV_X1 U11644 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n15093) );
  NOR2_X1 U11645 ( .A1(n9181), .A2(n15093), .ZN(P3_U3236) );
  INV_X1 U11646 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9202) );
  NOR2_X1 U11647 ( .A1(n9203), .A2(n9202), .ZN(P3_U3247) );
  INV_X1 U11648 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9204) );
  NOR2_X1 U11649 ( .A1(n9203), .A2(n9204), .ZN(P3_U3241) );
  INV_X1 U11650 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9205) );
  NOR2_X1 U11651 ( .A1(n9203), .A2(n9205), .ZN(P3_U3239) );
  INV_X1 U11652 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9206) );
  NOR2_X1 U11653 ( .A1(n9203), .A2(n9206), .ZN(P3_U3237) );
  NAND2_X1 U11654 ( .A1(n9283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9208) );
  XNOR2_X1 U11655 ( .A(n9208), .B(P2_IR_REG_8__SCAN_IN), .ZN(n13114) );
  INV_X1 U11656 ( .A(n13114), .ZN(n13107) );
  OAI222_X1 U11657 ( .A1(P2_U3088), .A2(n13107), .B1(n13574), .B2(n10276), 
        .C1(n9209), .C2(n13580), .ZN(P2_U3319) );
  INV_X1 U11658 ( .A(n9451), .ZN(n9429) );
  OAI222_X1 U11659 ( .A1(P1_U3086), .A2(n9429), .B1(n14305), .B2(n10276), .C1(
        n9210), .C2(n14302), .ZN(P1_U3347) );
  INV_X1 U11660 ( .A(n11357), .ZN(n9222) );
  INV_X1 U11661 ( .A(n9214), .ZN(n9215) );
  AOI21_X1 U11662 ( .B1(n10302), .B2(n9215), .A(n10301), .ZN(n9216) );
  INV_X1 U11663 ( .A(n9334), .ZN(n13048) );
  NAND2_X1 U11664 ( .A1(n9015), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9218) );
  MUX2_X1 U11665 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9218), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n9219) );
  AND2_X1 U11666 ( .A1(n13048), .A2(n13049), .ZN(n9387) );
  NAND2_X1 U11667 ( .A1(n9387), .A2(n11357), .ZN(n9220) );
  NAND2_X1 U11668 ( .A1(n10495), .A2(n9220), .ZN(n9221) );
  OAI21_X1 U11669 ( .B1(n9388), .B2(n9222), .A(n9221), .ZN(n9240) );
  AND2_X1 U11670 ( .A1(n9223), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9224) );
  AND2_X1 U11671 ( .A1(n9240), .A2(n9224), .ZN(n14770) );
  NOR2_X1 U11672 ( .A1(n9223), .A2(P2_U3088), .ZN(n13571) );
  AND2_X1 U11673 ( .A1(n9240), .A2(n13571), .ZN(n9248) );
  INV_X1 U11674 ( .A(n9248), .ZN(n9225) );
  INV_X1 U11675 ( .A(n13577), .ZN(n13044) );
  INV_X1 U11676 ( .A(n14747), .ZN(n14774) );
  INV_X1 U11677 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9226) );
  MUX2_X1 U11678 ( .A(n9226), .B(P2_REG1_REG_2__SCAN_IN), .S(n14666), .Z(
        n14672) );
  INV_X1 U11679 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9227) );
  MUX2_X1 U11680 ( .A(n9227), .B(P2_REG1_REG_1__SCAN_IN), .S(n13082), .Z(n9229) );
  AND2_X1 U11681 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9228) );
  NAND2_X1 U11682 ( .A1(n9229), .A2(n9228), .ZN(n13081) );
  OAI21_X1 U11683 ( .B1(n9227), .B2(n13082), .A(n13081), .ZN(n14673) );
  NAND2_X1 U11684 ( .A1(n14672), .A2(n14673), .ZN(n14671) );
  OR2_X1 U11685 ( .A1(n14666), .A2(n9226), .ZN(n9230) );
  NAND2_X1 U11686 ( .A1(n14671), .A2(n9230), .ZN(n14682) );
  INV_X1 U11687 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9231) );
  MUX2_X1 U11688 ( .A(n9231), .B(P2_REG1_REG_3__SCAN_IN), .S(n9643), .Z(n14681) );
  NAND2_X1 U11689 ( .A1(n14682), .A2(n14681), .ZN(n14680) );
  INV_X1 U11690 ( .A(n9643), .ZN(n14678) );
  NAND2_X1 U11691 ( .A1(n14678), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n13100) );
  NAND2_X1 U11692 ( .A1(n14680), .A2(n13100), .ZN(n9234) );
  INV_X1 U11693 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9232) );
  MUX2_X1 U11694 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9232), .S(n13098), .Z(n9233) );
  NAND2_X1 U11695 ( .A1(n9234), .A2(n9233), .ZN(n13102) );
  NAND2_X1 U11696 ( .A1(n13098), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U11697 ( .A1(n13102), .A2(n9238), .ZN(n9236) );
  MUX2_X1 U11698 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10226), .S(n9846), .Z(n9235) );
  NAND2_X1 U11699 ( .A1(n9236), .A2(n9235), .ZN(n9262) );
  INV_X1 U11700 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10226) );
  MUX2_X1 U11701 ( .A(n10226), .B(P2_REG1_REG_5__SCAN_IN), .S(n9846), .Z(n9237) );
  NAND3_X1 U11702 ( .A1(n13102), .A2(n9238), .A3(n9237), .ZN(n9239) );
  NAND3_X1 U11703 ( .A1(n14774), .A2(n9262), .A3(n9239), .ZN(n9254) );
  OR2_X1 U11704 ( .A1(n9240), .A2(P2_U3088), .ZN(n14744) );
  INV_X1 U11705 ( .A(n14744), .ZN(n14768) );
  NAND2_X1 U11706 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n9864) );
  INV_X1 U11707 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9241) );
  MUX2_X1 U11708 ( .A(n9241), .B(P2_REG2_REG_2__SCAN_IN), .S(n14666), .Z(
        n14669) );
  INV_X1 U11709 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n13083) );
  MUX2_X1 U11710 ( .A(n13083), .B(P2_REG2_REG_1__SCAN_IN), .S(n13082), .Z(
        n9243) );
  AND2_X1 U11711 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9242) );
  NAND2_X1 U11712 ( .A1(n9243), .A2(n9242), .ZN(n13087) );
  OAI21_X1 U11713 ( .B1(n13083), .B2(n13082), .A(n13087), .ZN(n14670) );
  NAND2_X1 U11714 ( .A1(n14669), .A2(n14670), .ZN(n14668) );
  OR2_X1 U11715 ( .A1(n14666), .A2(n9241), .ZN(n9244) );
  NAND2_X1 U11716 ( .A1(n14668), .A2(n9244), .ZN(n14685) );
  INV_X1 U11717 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10162) );
  MUX2_X1 U11718 ( .A(n10162), .B(P2_REG2_REG_3__SCAN_IN), .S(n9643), .Z(
        n14684) );
  NAND2_X1 U11719 ( .A1(n14685), .A2(n14684), .ZN(n14683) );
  NAND2_X1 U11720 ( .A1(n14678), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n13095) );
  NAND2_X1 U11721 ( .A1(n14683), .A2(n13095), .ZN(n9246) );
  INV_X1 U11722 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9914) );
  MUX2_X1 U11723 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9914), .S(n13098), .Z(n9245) );
  NAND2_X1 U11724 ( .A1(n9246), .A2(n9245), .ZN(n13097) );
  NAND2_X1 U11725 ( .A1(n13098), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U11726 ( .A1(n13097), .A2(n9247), .ZN(n9250) );
  INV_X1 U11727 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10214) );
  MUX2_X1 U11728 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10214), .S(n9846), .Z(n9249) );
  NAND2_X1 U11729 ( .A1(n9250), .A2(n9249), .ZN(n9273) );
  OAI211_X1 U11730 ( .C1(n9250), .C2(n9249), .A(n14776), .B(n9273), .ZN(n9251)
         );
  NAND2_X1 U11731 ( .A1(n9864), .A2(n9251), .ZN(n9252) );
  AOI21_X1 U11732 ( .B1(n14768), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n9252), .ZN(
        n9253) );
  OAI211_X1 U11733 ( .C1(n14740), .C2(n9255), .A(n9254), .B(n9253), .ZN(
        P2_U3219) );
  INV_X1 U11734 ( .A(n14578), .ZN(n14577) );
  NAND2_X1 U11735 ( .A1(n11610), .A2(n11450), .ZN(n9506) );
  OAI22_X1 U11736 ( .A1(n14577), .A2(P1_D_REG_0__SCAN_IN), .B1(n9256), .B2(
        n9506), .ZN(n9257) );
  INV_X1 U11737 ( .A(n9257), .ZN(P1_U3445) );
  AOI222_X1 U11738 ( .A1(n9259), .A2(n12680), .B1(n14882), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_13_), .C2(n9258), .ZN(n9260) );
  INV_X1 U11739 ( .A(n9260), .ZN(P3_U3282) );
  NAND2_X1 U11740 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10070) );
  OAI21_X1 U11741 ( .B1(n14744), .B2(n7634), .A(n10070), .ZN(n9271) );
  NAND2_X1 U11742 ( .A1(n9846), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9261) );
  NAND2_X1 U11743 ( .A1(n9262), .A2(n9261), .ZN(n14693) );
  INV_X1 U11744 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9263) );
  MUX2_X1 U11745 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9263), .S(n14690), .Z(
        n14692) );
  NAND2_X1 U11746 ( .A1(n14693), .A2(n14692), .ZN(n14691) );
  NAND2_X1 U11747 ( .A1(n14690), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U11748 ( .A1(n14691), .A2(n9268), .ZN(n9266) );
  INV_X1 U11749 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9264) );
  MUX2_X1 U11750 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9264), .S(n10061), .Z(n9265) );
  NAND2_X1 U11751 ( .A1(n9266), .A2(n9265), .ZN(n13117) );
  MUX2_X1 U11752 ( .A(n9264), .B(P2_REG1_REG_7__SCAN_IN), .S(n10061), .Z(n9267) );
  NAND3_X1 U11753 ( .A1(n14691), .A2(n9268), .A3(n9267), .ZN(n9269) );
  AND3_X1 U11754 ( .A1(n14774), .A2(n13117), .A3(n9269), .ZN(n9270) );
  AOI211_X1 U11755 ( .C1(n14770), .C2(n10061), .A(n9271), .B(n9270), .ZN(n9281) );
  NAND2_X1 U11756 ( .A1(n9846), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U11757 ( .A1(n9273), .A2(n9272), .ZN(n14696) );
  INV_X1 U11758 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10177) );
  MUX2_X1 U11759 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10177), .S(n14690), .Z(
        n14695) );
  NAND2_X1 U11760 ( .A1(n14696), .A2(n14695), .ZN(n14694) );
  NAND2_X1 U11761 ( .A1(n14690), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11762 ( .A1(n14694), .A2(n9278), .ZN(n9276) );
  INV_X1 U11763 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9274) );
  MUX2_X1 U11764 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9274), .S(n10061), .Z(n9275) );
  NAND2_X1 U11765 ( .A1(n9276), .A2(n9275), .ZN(n13111) );
  MUX2_X1 U11766 ( .A(n9274), .B(P2_REG2_REG_7__SCAN_IN), .S(n10061), .Z(n9277) );
  NAND3_X1 U11767 ( .A1(n14694), .A2(n9278), .A3(n9277), .ZN(n9279) );
  NAND3_X1 U11768 ( .A1(n14776), .A2(n13111), .A3(n9279), .ZN(n9280) );
  NAND2_X1 U11769 ( .A1(n9281), .A2(n9280), .ZN(P2_U3221) );
  INV_X1 U11770 ( .A(n9488), .ZN(n9282) );
  INV_X1 U11771 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n15174) );
  OAI222_X1 U11772 ( .A1(P1_U3086), .A2(n9282), .B1(n14305), .B2(n10494), .C1(
        n15174), .C2(n14302), .ZN(P1_U3346) );
  NOR2_X1 U11773 ( .A1(n9286), .A2(n10301), .ZN(n9284) );
  MUX2_X1 U11774 ( .A(n10301), .B(n9284), .S(P2_IR_REG_9__SCAN_IN), .Z(n9288)
         );
  NAND2_X1 U11775 ( .A1(n9286), .A2(n9285), .ZN(n9575) );
  INV_X1 U11776 ( .A(n9575), .ZN(n9287) );
  OAI222_X1 U11777 ( .A1(P2_U3088), .A2(n14705), .B1(n13574), .B2(n10494), 
        .C1(n10496), .C2(n13580), .ZN(P2_U3318) );
  NAND2_X1 U11778 ( .A1(n9575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9289) );
  XNOR2_X1 U11779 ( .A(n9289), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10735) );
  INV_X1 U11780 ( .A(n10735), .ZN(n10086) );
  INV_X1 U11781 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n15106) );
  NAND2_X1 U11782 ( .A1(n10061), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n13116) );
  NAND2_X1 U11783 ( .A1(n13117), .A2(n13116), .ZN(n9291) );
  MUX2_X1 U11784 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n15262), .S(n13114), .Z(
        n9290) );
  NAND2_X1 U11785 ( .A1(n9291), .A2(n9290), .ZN(n13119) );
  NAND2_X1 U11786 ( .A1(n13114), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U11787 ( .A1(n13119), .A2(n9292), .ZN(n14708) );
  MUX2_X1 U11788 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n15106), .S(n14705), .Z(
        n14707) );
  NOR2_X1 U11789 ( .A1(n14708), .A2(n14707), .ZN(n14710) );
  AOI21_X1 U11790 ( .B1(n15106), .B2(n14705), .A(n14710), .ZN(n9295) );
  INV_X1 U11791 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9293) );
  MUX2_X1 U11792 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9293), .S(n10735), .Z(
        n9294) );
  NAND2_X1 U11793 ( .A1(n9295), .A2(n9294), .ZN(n10083) );
  OAI211_X1 U11794 ( .C1(n9295), .C2(n9294), .A(n10083), .B(n14774), .ZN(n9307) );
  NAND2_X1 U11795 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14640)
         );
  INV_X1 U11796 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n13422) );
  NAND2_X1 U11797 ( .A1(n10061), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13110) );
  NAND2_X1 U11798 ( .A1(n13111), .A2(n13110), .ZN(n9298) );
  INV_X1 U11799 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9296) );
  MUX2_X1 U11800 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9296), .S(n13114), .Z(n9297) );
  NAND2_X1 U11801 ( .A1(n9298), .A2(n9297), .ZN(n13113) );
  NAND2_X1 U11802 ( .A1(n13114), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9299) );
  AND2_X1 U11803 ( .A1(n13113), .A2(n9299), .ZN(n14702) );
  MUX2_X1 U11804 ( .A(n13422), .B(P2_REG2_REG_9__SCAN_IN), .S(n14705), .Z(
        n14701) );
  AND2_X1 U11805 ( .A1(n14702), .A2(n14701), .ZN(n14704) );
  AOI21_X1 U11806 ( .B1(n14705), .B2(n13422), .A(n14704), .ZN(n9303) );
  INV_X1 U11807 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9300) );
  MUX2_X1 U11808 ( .A(n9300), .B(P2_REG2_REG_10__SCAN_IN), .S(n10735), .Z(
        n9301) );
  INV_X1 U11809 ( .A(n9301), .ZN(n9302) );
  NAND2_X1 U11810 ( .A1(n9303), .A2(n9302), .ZN(n10085) );
  OAI211_X1 U11811 ( .C1(n9303), .C2(n9302), .A(n14776), .B(n10085), .ZN(n9304) );
  NAND2_X1 U11812 ( .A1(n14640), .A2(n9304), .ZN(n9305) );
  AOI21_X1 U11813 ( .B1(n14768), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9305), .ZN(
        n9306) );
  OAI211_X1 U11814 ( .C1(n14740), .C2(n10086), .A(n9307), .B(n9306), .ZN(
        P2_U3224) );
  OAI222_X1 U11815 ( .A1(P2_U3088), .A2(n10086), .B1(n13578), .B2(n10734), 
        .C1(n9308), .C2(n13580), .ZN(P2_U3317) );
  INV_X1 U11816 ( .A(n9469), .ZN(n9405) );
  OAI222_X1 U11817 ( .A1(P1_U3086), .A2(n9405), .B1(n14305), .B2(n10734), .C1(
        n9309), .C2(n14302), .ZN(P1_U3345) );
  INV_X1 U11818 ( .A(n12231), .ZN(n9313) );
  INV_X1 U11819 ( .A(n9310), .ZN(n9311) );
  OAI222_X1 U11820 ( .A1(P3_U3151), .A2(n9313), .B1(n12698), .B2(n9312), .C1(
        n12694), .C2(n9311), .ZN(P3_U3281) );
  NAND2_X1 U11821 ( .A1(n9604), .A2(n11354), .ZN(n9409) );
  AOI21_X1 U11822 ( .B1(n9316), .B2(n9315), .A(n9314), .ZN(n9408) );
  INV_X1 U11823 ( .A(n9408), .ZN(n9317) );
  AND2_X1 U11824 ( .A1(n9409), .A2(n9317), .ZN(n14544) );
  NOR2_X1 U11825 ( .A1(n14544), .A2(P1_U4016), .ZN(P1_U3085) );
  XNOR2_X2 U11826 ( .A(n9321), .B(n9320), .ZN(n9324) );
  AND2_X4 U11827 ( .A1(n9323), .A2(n9322), .ZN(n12004) );
  NAND2_X1 U11828 ( .A1(n12004), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9327) );
  AND2_X2 U11829 ( .A1(n9322), .A2(n13569), .ZN(n9534) );
  NAND2_X1 U11830 ( .A1(n9649), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9325) );
  NAND3_X1 U11831 ( .A1(n9327), .A2(n9326), .A3(n9325), .ZN(n9385) );
  NAND2_X1 U11832 ( .A1(n9343), .A2(SI_0_), .ZN(n9328) );
  XNOR2_X1 U11833 ( .A(n9328), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13581) );
  MUX2_X1 U11834 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13581), .S(n9346), .Z(n9883)
         );
  NAND2_X1 U11835 ( .A1(n9385), .A2(n9883), .ZN(n9871) );
  NAND2_X1 U11836 ( .A1(n9334), .A2(n12968), .ZN(n14796) );
  INV_X2 U11837 ( .A(n9819), .ZN(n9331) );
  NAND2_X1 U11838 ( .A1(n9335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9337) );
  XNOR2_X2 U11839 ( .A(n9337), .B(n9336), .ZN(n13412) );
  NAND2_X1 U11840 ( .A1(n9534), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U11841 ( .A1(n9536), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U11842 ( .A1(n9649), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U11843 ( .A1(n12004), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9340) );
  INV_X2 U11844 ( .A(n9459), .ZN(n10803) );
  NAND2_X1 U11845 ( .A1(n13075), .A2(n6519), .ZN(n9353) );
  INV_X1 U11846 ( .A(n9353), .ZN(n9351) );
  INV_X1 U11847 ( .A(n9352), .ZN(n9350) );
  NAND2_X1 U11848 ( .A1(n9351), .A2(n9350), .ZN(n9354) );
  AOI21_X1 U11849 ( .B1(n9356), .B2(n9355), .A(n9525), .ZN(n9393) );
  XNOR2_X1 U11850 ( .A(n11333), .B(P2_B_REG_SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11851 ( .A1(n9358), .A2(n11370), .ZN(n9360) );
  INV_X1 U11852 ( .A(n11453), .ZN(n9359) );
  INV_X1 U11853 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14821) );
  AOI22_X1 U11854 ( .A1(n14812), .A2(n14821), .B1(n11453), .B2(n11370), .ZN(
        n9885) );
  NOR4_X1 U11855 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n9364) );
  NOR4_X1 U11856 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9363) );
  NOR4_X1 U11857 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n9362) );
  NOR4_X1 U11858 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n9361) );
  NAND4_X1 U11859 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(n9369)
         );
  NOR4_X1 U11860 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n15043) );
  NOR2_X1 U11861 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n9367) );
  NOR4_X1 U11862 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n9366) );
  NOR4_X1 U11863 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9365) );
  NAND4_X1 U11864 ( .A1(n15043), .A2(n9367), .A3(n9366), .A4(n9365), .ZN(n9368) );
  OAI21_X1 U11865 ( .B1(n9369), .B2(n9368), .A(n14812), .ZN(n9887) );
  NAND2_X1 U11866 ( .A1(n9885), .A2(n9887), .ZN(n9386) );
  INV_X1 U11867 ( .A(n9386), .ZN(n9904) );
  NAND2_X1 U11868 ( .A1(n14817), .A2(n9904), .ZN(n9372) );
  INV_X1 U11869 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14815) );
  NAND2_X1 U11870 ( .A1(n14812), .A2(n14815), .ZN(n9371) );
  NAND2_X1 U11871 ( .A1(n11333), .A2(n11453), .ZN(n9370) );
  OR2_X1 U11872 ( .A1(n9372), .A2(n14816), .ZN(n9383) );
  INV_X1 U11873 ( .A(n9383), .ZN(n9376) );
  INV_X1 U11874 ( .A(n14796), .ZN(n9373) );
  INV_X1 U11875 ( .A(n9333), .ZN(n13039) );
  NAND2_X1 U11876 ( .A1(n13039), .A2(n13412), .ZN(n13042) );
  NAND2_X1 U11877 ( .A1(n9373), .A2(n13042), .ZN(n14837) );
  INV_X1 U11878 ( .A(n9387), .ZN(n9374) );
  AND2_X1 U11879 ( .A1(n14837), .A2(n9374), .ZN(n9375) );
  NAND2_X1 U11880 ( .A1(n12783), .A2(n13407), .ZN(n14419) );
  INV_X1 U11881 ( .A(n14419), .ZN(n12798) );
  NAND2_X1 U11882 ( .A1(n9534), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9380) );
  NAND2_X1 U11883 ( .A1(n12004), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9379) );
  NAND2_X1 U11884 ( .A1(n9649), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U11885 ( .A1(n9536), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9377) );
  OR2_X1 U11886 ( .A1(n14796), .A2(n13039), .ZN(n9918) );
  INV_X1 U11887 ( .A(n9886), .ZN(n9382) );
  OAI21_X2 U11888 ( .B1(n9383), .B2(n9918), .A(n14803), .ZN(n14657) );
  AOI22_X1 U11889 ( .A1(n12798), .A2(n13074), .B1(n9381), .B2(n14657), .ZN(
        n9392) );
  INV_X1 U11890 ( .A(n9223), .ZN(n9384) );
  NAND2_X1 U11891 ( .A1(n12783), .A2(n13405), .ZN(n14418) );
  INV_X1 U11892 ( .A(n14418), .ZN(n12801) );
  OAI21_X1 U11893 ( .B1(n14816), .B2(n9386), .A(n9886), .ZN(n9390) );
  NAND2_X1 U11894 ( .A1(n9387), .A2(n13042), .ZN(n9903) );
  AND3_X1 U11895 ( .A1(n9388), .A2(n11357), .A3(n9903), .ZN(n9389) );
  NAND2_X1 U11896 ( .A1(n9390), .A2(n9389), .ZN(n9647) );
  OR2_X1 U11897 ( .A1(n9647), .A2(P2_U3088), .ZN(n9541) );
  AOI22_X1 U11898 ( .A1(n12801), .A2(n9385), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9541), .ZN(n9391) );
  OAI211_X1 U11899 ( .C1(n9393), .C2(n14652), .A(n9392), .B(n9391), .ZN(
        P2_U3194) );
  MUX2_X1 U11900 ( .A(n11112), .B(P1_REG2_REG_12__SCAN_IN), .S(n9434), .Z(
        n9407) );
  INV_X1 U11901 ( .A(n13950), .ZN(n9578) );
  MUX2_X1 U11902 ( .A(n9394), .B(P1_REG2_REG_2__SCAN_IN), .S(n13884), .Z(
        n13882) );
  MUX2_X1 U11903 ( .A(n9395), .B(P1_REG2_REG_1__SCAN_IN), .S(n13867), .Z(
        n13866) );
  AND2_X1 U11904 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13877) );
  NAND2_X1 U11905 ( .A1(n13866), .A2(n13877), .ZN(n13865) );
  OAI21_X1 U11906 ( .B1(n9395), .B2(n13867), .A(n13865), .ZN(n13881) );
  NAND2_X1 U11907 ( .A1(n13882), .A2(n13881), .ZN(n13899) );
  OR2_X1 U11908 ( .A1(n13884), .A2(n9394), .ZN(n13898) );
  NAND2_X1 U11909 ( .A1(n13899), .A2(n13898), .ZN(n9397) );
  MUX2_X1 U11910 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10384), .S(n13896), .Z(
        n9396) );
  NAND2_X1 U11911 ( .A1(n9397), .A2(n9396), .ZN(n13919) );
  NAND2_X1 U11912 ( .A1(n13896), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13918) );
  MUX2_X1 U11913 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10392), .S(n13914), .Z(
        n13917) );
  AOI21_X1 U11914 ( .B1(n13919), .B2(n13918), .A(n13917), .ZN(n13916) );
  NOR2_X1 U11915 ( .A1(n13914), .A2(n10392), .ZN(n9563) );
  MUX2_X1 U11916 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9398), .S(n9566), .Z(n9562)
         );
  OAI21_X1 U11917 ( .B1(n13916), .B2(n9563), .A(n9562), .ZN(n13937) );
  NAND2_X1 U11918 ( .A1(n9566), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n13936) );
  INV_X1 U11919 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9399) );
  MUX2_X1 U11920 ( .A(n9399), .B(P1_REG2_REG_6__SCAN_IN), .S(n13929), .Z(
        n13935) );
  AOI21_X1 U11921 ( .B1(n13937), .B2(n13936), .A(n13935), .ZN(n13934) );
  NOR2_X1 U11922 ( .A1(n9400), .A2(n9399), .ZN(n9545) );
  INV_X1 U11923 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9401) );
  MUX2_X1 U11924 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9401), .S(n9546), .Z(n9402)
         );
  OAI21_X1 U11925 ( .B1(n13934), .B2(n9545), .A(n9402), .ZN(n9549) );
  NAND2_X1 U11926 ( .A1(n9546), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9453) );
  INV_X1 U11927 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9403) );
  MUX2_X1 U11928 ( .A(n9403), .B(P1_REG2_REG_8__SCAN_IN), .S(n9451), .Z(n9452)
         );
  AOI21_X1 U11929 ( .B1(n9549), .B2(n9453), .A(n9452), .ZN(n9479) );
  NOR2_X1 U11930 ( .A1(n9429), .A2(n9403), .ZN(n9478) );
  MUX2_X1 U11931 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10631), .S(n9488), .Z(n9477) );
  OAI21_X1 U11932 ( .B1(n9479), .B2(n9478), .A(n9477), .ZN(n9476) );
  NAND2_X1 U11933 ( .A1(n9488), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9465) );
  INV_X1 U11934 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9404) );
  MUX2_X1 U11935 ( .A(n9404), .B(P1_REG2_REG_10__SCAN_IN), .S(n9469), .Z(n9464) );
  AOI21_X1 U11936 ( .B1(n9476), .B2(n9465), .A(n9464), .ZN(n13945) );
  NOR2_X1 U11937 ( .A1(n9405), .A2(n9404), .ZN(n13944) );
  MUX2_X1 U11938 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10957), .S(n13950), .Z(
        n13943) );
  OAI21_X1 U11939 ( .B1(n13945), .B2(n13944), .A(n13943), .ZN(n13947) );
  OAI21_X1 U11940 ( .B1(n9578), .B2(n10957), .A(n13947), .ZN(n9406) );
  NOR2_X1 U11941 ( .A1(n9406), .A2(n9407), .ZN(n9613) );
  AOI21_X1 U11942 ( .B1(n9407), .B2(n9406), .A(n9613), .ZN(n9444) );
  NAND2_X1 U11943 ( .A1(n9409), .A2(n9408), .ZN(n14546) );
  OR3_X1 U11944 ( .A1(n14546), .A2(n6530), .A3(n13873), .ZN(n14552) );
  INV_X1 U11945 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n13765) );
  NOR2_X1 U11946 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13765), .ZN(n9411) );
  INV_X1 U11947 ( .A(n9434), .ZN(n9716) );
  NOR2_X1 U11948 ( .A1(n14571), .A2(n9716), .ZN(n9410) );
  AOI211_X1 U11949 ( .C1(n14544), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9411), .B(
        n9410), .ZN(n9443) );
  INV_X1 U11950 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9412) );
  MUX2_X1 U11951 ( .A(n9412), .B(P1_REG1_REG_2__SCAN_IN), .S(n13884), .Z(
        n13887) );
  INV_X1 U11952 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15154) );
  MUX2_X1 U11953 ( .A(n15154), .B(P1_REG1_REG_1__SCAN_IN), .S(n13867), .Z(
        n9414) );
  AND2_X1 U11954 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9413) );
  NAND2_X1 U11955 ( .A1(n9414), .A2(n9413), .ZN(n13864) );
  OAI21_X1 U11956 ( .B1(n15154), .B2(n13867), .A(n13864), .ZN(n13886) );
  NAND2_X1 U11957 ( .A1(n13887), .A2(n13886), .ZN(n13894) );
  OR2_X1 U11958 ( .A1(n13884), .A2(n9412), .ZN(n13893) );
  NAND2_X1 U11959 ( .A1(n13894), .A2(n13893), .ZN(n9417) );
  MUX2_X1 U11960 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9415), .S(n13896), .Z(n9416) );
  NAND2_X1 U11961 ( .A1(n9417), .A2(n9416), .ZN(n13910) );
  NAND2_X1 U11962 ( .A1(n13896), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n13909) );
  NAND2_X1 U11963 ( .A1(n13910), .A2(n13909), .ZN(n9420) );
  MUX2_X1 U11964 ( .A(n9418), .B(P1_REG1_REG_4__SCAN_IN), .S(n13914), .Z(n9419) );
  NAND2_X1 U11965 ( .A1(n9420), .A2(n9419), .ZN(n13912) );
  NAND2_X1 U11966 ( .A1(n9421), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9422) );
  AND2_X1 U11967 ( .A1(n13912), .A2(n9422), .ZN(n9560) );
  MUX2_X1 U11968 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7806), .S(n9566), .Z(n9561)
         );
  NAND2_X1 U11969 ( .A1(n9560), .A2(n9561), .ZN(n9559) );
  NAND2_X1 U11970 ( .A1(n9423), .A2(n7806), .ZN(n9424) );
  NAND2_X1 U11971 ( .A1(n9559), .A2(n9424), .ZN(n13931) );
  MUX2_X1 U11972 ( .A(n7818), .B(P1_REG1_REG_6__SCAN_IN), .S(n13929), .Z(
        n13930) );
  OR2_X1 U11973 ( .A1(n13931), .A2(n13930), .ZN(n13933) );
  NAND2_X1 U11974 ( .A1(n13929), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U11975 ( .A1(n13933), .A2(n9425), .ZN(n9553) );
  MUX2_X1 U11976 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9426), .S(n9546), .Z(n9552)
         );
  NAND2_X1 U11977 ( .A1(n9553), .A2(n9552), .ZN(n9551) );
  NAND2_X1 U11978 ( .A1(n9546), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U11979 ( .A1(n9551), .A2(n9427), .ZN(n9447) );
  MUX2_X1 U11980 ( .A(n9428), .B(P1_REG1_REG_8__SCAN_IN), .S(n9451), .Z(n9448)
         );
  OR2_X1 U11981 ( .A1(n9447), .A2(n9448), .ZN(n9485) );
  NAND2_X1 U11982 ( .A1(n9429), .A2(n9428), .ZN(n9483) );
  NAND2_X1 U11983 ( .A1(n9485), .A2(n9483), .ZN(n9430) );
  MUX2_X1 U11984 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7885), .S(n9488), .Z(n9482)
         );
  NAND2_X1 U11985 ( .A1(n9430), .A2(n9482), .ZN(n9487) );
  OR2_X1 U11986 ( .A1(n9488), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9431) );
  AND2_X1 U11987 ( .A1(n9487), .A2(n9431), .ZN(n9472) );
  MUX2_X1 U11988 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9432), .S(n9469), .Z(n9471) );
  NAND2_X1 U11989 ( .A1(n9472), .A2(n9471), .ZN(n9470) );
  NAND2_X1 U11990 ( .A1(n9469), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9433) );
  AND2_X1 U11991 ( .A1(n9470), .A2(n9433), .ZN(n13952) );
  MUX2_X1 U11992 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7929), .S(n13950), .Z(
        n13953) );
  NAND2_X1 U11993 ( .A1(n13952), .A2(n13953), .ZN(n13951) );
  INV_X1 U11994 ( .A(n13951), .ZN(n9436) );
  MUX2_X1 U11995 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7947), .S(n9434), .Z(n9438) );
  OR2_X1 U11996 ( .A1(n13950), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9437) );
  INV_X1 U11997 ( .A(n9437), .ZN(n9435) );
  NOR3_X1 U11998 ( .A1(n9436), .A2(n9438), .A3(n9435), .ZN(n9441) );
  NAND2_X1 U11999 ( .A1(n13951), .A2(n9437), .ZN(n9439) );
  NAND2_X1 U12000 ( .A1(n9439), .A2(n9438), .ZN(n9620) );
  INV_X1 U12001 ( .A(n9620), .ZN(n9440) );
  INV_X1 U12002 ( .A(n14557), .ZN(n14566) );
  OAI21_X1 U12003 ( .B1(n9441), .B2(n9440), .A(n14566), .ZN(n9442) );
  OAI211_X1 U12004 ( .C1(n9444), .C2(n14552), .A(n9443), .B(n9442), .ZN(
        P1_U3255) );
  INV_X1 U12005 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U12006 ( .A1(P1_U4016), .A2(n13975), .ZN(n9445) );
  OAI21_X1 U12007 ( .B1(P1_U4016), .B2(n11760), .A(n9445), .ZN(P1_U3591) );
  INV_X1 U12008 ( .A(n9485), .ZN(n9446) );
  AOI21_X1 U12009 ( .B1(n9448), .B2(n9447), .A(n9446), .ZN(n9458) );
  INV_X1 U12010 ( .A(n14571), .ZN(n13963) );
  NAND2_X1 U12011 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11024) );
  OAI21_X1 U12012 ( .B1(n14575), .B2(n9449), .A(n11024), .ZN(n9450) );
  AOI21_X1 U12013 ( .B1(n9451), .B2(n13963), .A(n9450), .ZN(n9457) );
  INV_X1 U12014 ( .A(n9479), .ZN(n9455) );
  NAND3_X1 U12015 ( .A1(n9549), .A2(n9453), .A3(n9452), .ZN(n9454) );
  NAND3_X1 U12016 ( .A1(n9455), .A2(n14563), .A3(n9454), .ZN(n9456) );
  OAI211_X1 U12017 ( .C1(n9458), .C2(n14557), .A(n9457), .B(n9456), .ZN(
        P1_U3251) );
  NAND2_X1 U12018 ( .A1(n9385), .A2(n14797), .ZN(n13004) );
  MUX2_X1 U12019 ( .A(n13004), .B(n14797), .S(n10803), .Z(n9460) );
  INV_X1 U12020 ( .A(n9385), .ZN(n9935) );
  NAND2_X1 U12021 ( .A1(n9935), .A2(n9883), .ZN(n13005) );
  AOI21_X1 U12022 ( .B1(n9460), .B2(n13005), .A(n14652), .ZN(n9462) );
  INV_X2 U12023 ( .A(n13075), .ZN(n14800) );
  OAI22_X1 U12024 ( .A1(n14415), .A2(n14797), .B1(n14419), .B2(n14800), .ZN(
        n9461) );
  AOI211_X1 U12025 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n9541), .A(n9462), .B(
        n9461), .ZN(n9463) );
  INV_X1 U12026 ( .A(n9463), .ZN(P2_U3204) );
  NAND3_X1 U12027 ( .A1(n9476), .A2(n9465), .A3(n9464), .ZN(n9466) );
  NAND2_X1 U12028 ( .A1(n9466), .A2(n14563), .ZN(n9475) );
  AND2_X1 U12029 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11350) );
  NOR2_X1 U12030 ( .A1(n14575), .A2(n9467), .ZN(n9468) );
  AOI211_X1 U12031 ( .C1(n13963), .C2(n9469), .A(n11350), .B(n9468), .ZN(n9474) );
  OAI211_X1 U12032 ( .C1(n9472), .C2(n9471), .A(n9470), .B(n14566), .ZN(n9473)
         );
  OAI211_X1 U12033 ( .C1(n13945), .C2(n9475), .A(n9474), .B(n9473), .ZN(
        P1_U3253) );
  INV_X1 U12034 ( .A(n9476), .ZN(n9481) );
  NOR3_X1 U12035 ( .A1(n9479), .A2(n9478), .A3(n9477), .ZN(n9480) );
  NOR3_X1 U12036 ( .A1(n9481), .A2(n9480), .A3(n14552), .ZN(n9493) );
  INV_X1 U12037 ( .A(n9482), .ZN(n9484) );
  NAND3_X1 U12038 ( .A1(n9485), .A2(n9484), .A3(n9483), .ZN(n9486) );
  AOI21_X1 U12039 ( .B1(n9487), .B2(n9486), .A(n14557), .ZN(n9492) );
  INV_X1 U12040 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U12041 ( .A1(n13963), .A2(n9488), .ZN(n9489) );
  NAND2_X1 U12042 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11162) );
  OAI211_X1 U12043 ( .C1(n9490), .C2(n14575), .A(n9489), .B(n11162), .ZN(n9491) );
  OR3_X1 U12044 ( .A1(n9493), .A2(n9492), .A3(n9491), .ZN(P1_U3252) );
  NOR4_X1 U12045 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n9497) );
  NOR4_X1 U12046 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n9496) );
  NOR4_X1 U12047 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9495) );
  NOR4_X1 U12048 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9494) );
  NAND4_X1 U12049 ( .A1(n9497), .A2(n9496), .A3(n9495), .A4(n9494), .ZN(n9503)
         );
  NOR2_X1 U12050 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .ZN(
        n9501) );
  NOR4_X1 U12051 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9500) );
  NOR4_X1 U12052 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9499) );
  NOR4_X1 U12053 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9498) );
  NAND4_X1 U12054 ( .A1(n9501), .A2(n9500), .A3(n9499), .A4(n9498), .ZN(n9502)
         );
  NOR2_X1 U12055 ( .A1(n9503), .A2(n9502), .ZN(n9504) );
  OR2_X1 U12056 ( .A1(n9508), .A2(n9504), .ZN(n9583) );
  NAND2_X1 U12057 ( .A1(n9583), .A2(n9505), .ZN(n10307) );
  OR2_X1 U12058 ( .A1(n9508), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U12059 ( .A1(n9507), .A2(n9506), .ZN(n9585) );
  OR2_X1 U12060 ( .A1(n9508), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9510) );
  NAND2_X1 U12061 ( .A1(n9510), .A2(n9509), .ZN(n10306) );
  OR2_X1 U12062 ( .A1(n9590), .A2(n11295), .ZN(n9606) );
  NAND2_X1 U12063 ( .A1(n10306), .A2(n9606), .ZN(n9517) );
  INV_X1 U12064 ( .A(n9602), .ZN(n9587) );
  INV_X2 U12065 ( .A(n7544), .ZN(n13705) );
  OAI21_X1 U12066 ( .B1(n9591), .B2(n9511), .A(n13705), .ZN(n10315) );
  NOR2_X1 U12067 ( .A1(n9601), .A2(n11295), .ZN(n9512) );
  NAND2_X1 U12068 ( .A1(n8349), .A2(n9512), .ZN(n14219) );
  NAND2_X1 U12069 ( .A1(n8348), .A2(n10792), .ZN(n9514) );
  OAI21_X1 U12070 ( .B1(n14615), .B2(n14264), .A(n10317), .ZN(n9515) );
  NAND2_X1 U12071 ( .A1(n13859), .A2(n14152), .ZN(n10310) );
  OAI211_X1 U12072 ( .C1(n9587), .C2(n10312), .A(n9515), .B(n10310), .ZN(n9518) );
  NAND2_X1 U12073 ( .A1(n14636), .A2(n9518), .ZN(n9516) );
  OAI21_X1 U12074 ( .B1(n14636), .B2(n9594), .A(n9516), .ZN(P1_U3528) );
  INV_X1 U12075 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9520) );
  NAND2_X1 U12076 ( .A1(n14627), .A2(n9518), .ZN(n9519) );
  OAI21_X1 U12077 ( .B1(n14627), .B2(n9520), .A(n9519), .ZN(P1_U3459) );
  INV_X1 U12078 ( .A(n9521), .ZN(n9522) );
  OAI222_X1 U12079 ( .A1(n12698), .A2(n9523), .B1(n12694), .B2(n9522), .C1(
        n12277), .C2(P3_U3151), .ZN(P3_U3280) );
  NAND2_X1 U12080 ( .A1(n13074), .A2(n9459), .ZN(n9531) );
  OR2_X1 U12081 ( .A1(n12965), .A2(n9526), .ZN(n9529) );
  OR2_X1 U12082 ( .A1(n11375), .A2(n9527), .ZN(n9528) );
  XNOR2_X1 U12083 ( .A(n6534), .B(n9744), .ZN(n9530) );
  NAND2_X1 U12084 ( .A1(n9531), .A2(n9530), .ZN(n9644) );
  OAI21_X1 U12085 ( .B1(n9531), .B2(n9530), .A(n9644), .ZN(n9532) );
  AOI21_X1 U12086 ( .B1(n9533), .B2(n9532), .A(n9646), .ZN(n9544) );
  INV_X2 U12087 ( .A(n9970), .ZN(n12941) );
  NAND2_X1 U12088 ( .A1(n11977), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9540) );
  INV_X1 U12089 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U12090 ( .A1(n12004), .A2(n9535), .ZN(n9539) );
  NAND2_X1 U12091 ( .A1(n9649), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9538) );
  CLKBUF_X3 U12092 ( .A(n9536), .Z(n12958) );
  NAND2_X1 U12093 ( .A1(n12958), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9537) );
  NAND4_X1 U12094 ( .A1(n9540), .A2(n9539), .A3(n9538), .A4(n9537), .ZN(n13073) );
  AOI22_X1 U12095 ( .A1(n12798), .A2(n13073), .B1(n6534), .B2(n14657), .ZN(
        n9543) );
  AOI22_X1 U12096 ( .A1(n12801), .A2(n13075), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n9541), .ZN(n9542) );
  OAI211_X1 U12097 ( .C1(n9544), .C2(n14652), .A(n9543), .B(n9542), .ZN(
        P2_U3209) );
  INV_X1 U12098 ( .A(n9545), .ZN(n9548) );
  MUX2_X1 U12099 ( .A(n9401), .B(P1_REG2_REG_7__SCAN_IN), .S(n9546), .Z(n9547)
         );
  NAND2_X1 U12100 ( .A1(n9548), .A2(n9547), .ZN(n9550) );
  OAI211_X1 U12101 ( .C1(n13934), .C2(n9550), .A(n14563), .B(n9549), .ZN(n9557) );
  NAND2_X1 U12102 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10684) );
  OAI211_X1 U12103 ( .C1(n9553), .C2(n9552), .A(n14566), .B(n9551), .ZN(n9554)
         );
  NAND2_X1 U12104 ( .A1(n10684), .A2(n9554), .ZN(n9555) );
  AOI21_X1 U12105 ( .B1(n14544), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9555), .ZN(
        n9556) );
  OAI211_X1 U12106 ( .C1(n14571), .C2(n9558), .A(n9557), .B(n9556), .ZN(
        P1_U3250) );
  OAI21_X1 U12107 ( .B1(n9561), .B2(n9560), .A(n9559), .ZN(n9571) );
  INV_X1 U12108 ( .A(n13937), .ZN(n9565) );
  NOR3_X1 U12109 ( .A1(n13916), .A2(n9563), .A3(n9562), .ZN(n9564) );
  NOR3_X1 U12110 ( .A1(n14552), .A2(n9565), .A3(n9564), .ZN(n9570) );
  NAND2_X1 U12111 ( .A1(n13963), .A2(n9566), .ZN(n9567) );
  NAND2_X1 U12112 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10350) );
  OAI211_X1 U12113 ( .C1(n9568), .C2(n14575), .A(n9567), .B(n10350), .ZN(n9569) );
  AOI211_X1 U12114 ( .C1(n14566), .C2(n9571), .A(n9570), .B(n9569), .ZN(n9572)
         );
  INV_X1 U12115 ( .A(n9572), .ZN(P1_U3248) );
  INV_X1 U12116 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n15094) );
  NAND2_X1 U12117 ( .A1(n14945), .A2(P3_U3897), .ZN(n9573) );
  OAI21_X1 U12118 ( .B1(P3_U3897), .B2(n15094), .A(n9573), .ZN(P3_U3493) );
  INV_X1 U12119 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n15243) );
  NAND2_X1 U12120 ( .A1(n12076), .A2(P3_U3897), .ZN(n9574) );
  OAI21_X1 U12121 ( .B1(P3_U3897), .B2(n15243), .A(n9574), .ZN(P3_U3502) );
  INV_X1 U12122 ( .A(n10747), .ZN(n9579) );
  NAND2_X1 U12123 ( .A1(n9712), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9576) );
  XNOR2_X1 U12124 ( .A(n9576), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10748) );
  INV_X1 U12125 ( .A(n10748), .ZN(n14721) );
  OAI222_X1 U12126 ( .A1(n13580), .A2(n9577), .B1(n13578), .B2(n9579), .C1(
        P2_U3088), .C2(n14721), .ZN(P2_U3316) );
  OAI222_X1 U12127 ( .A1(n14302), .A2(n9580), .B1(n14305), .B2(n9579), .C1(
        P1_U3086), .C2(n9578), .ZN(P1_U3344) );
  INV_X1 U12128 ( .A(n12281), .ZN(n12272) );
  OAI222_X1 U12129 ( .A1(P3_U3151), .A2(n12272), .B1(n12694), .B2(n9582), .C1(
        n9581), .C2(n12698), .ZN(P3_U3279) );
  INV_X1 U12130 ( .A(n9583), .ZN(n9584) );
  NOR2_X1 U12131 ( .A1(n9607), .A2(n9604), .ZN(n9603) );
  AND2_X1 U12132 ( .A1(n14609), .A2(n9588), .ZN(n9589) );
  INV_X1 U12133 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13862) );
  OAI22_X1 U12134 ( .A1(n13741), .A2(n10312), .B1(n9595), .B2(n13862), .ZN(
        n9593) );
  AOI21_X1 U12135 ( .B1(n13860), .B2(n10343), .A(n9593), .ZN(n9599) );
  OR2_X1 U12136 ( .A1(n10404), .A2(n13741), .ZN(n9598) );
  OAI22_X1 U12137 ( .A1(n13739), .A2(n10312), .B1(n9595), .B2(n9594), .ZN(
        n9596) );
  INV_X1 U12138 ( .A(n9596), .ZN(n9597) );
  NAND2_X1 U12139 ( .A1(n9598), .A2(n9597), .ZN(n9694) );
  AOI22_X1 U12140 ( .A1(n14464), .A2(n13875), .B1(n14457), .B2(n13859), .ZN(
        n9612) );
  AND2_X1 U12141 ( .A1(n9602), .A2(n9601), .ZN(n10311) );
  NAND2_X1 U12142 ( .A1(n9603), .A2(n10311), .ZN(n9605) );
  NAND2_X1 U12143 ( .A1(n9607), .A2(n9606), .ZN(n9610) );
  INV_X1 U12144 ( .A(n9608), .ZN(n9609) );
  NAND2_X1 U12145 ( .A1(n9610), .A2(n9609), .ZN(n9958) );
  OR2_X1 U12146 ( .A1(n9958), .A2(P1_U3086), .ZN(n9708) );
  AOI22_X1 U12147 ( .A1(n14481), .A2(n10400), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n9708), .ZN(n9611) );
  NAND2_X1 U12148 ( .A1(n9612), .A2(n9611), .ZN(P1_U3232) );
  AOI21_X1 U12149 ( .B1(n11112), .B2(n9716), .A(n9613), .ZN(n9634) );
  MUX2_X1 U12150 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11202), .S(n9760), .Z(
        n9633) );
  NAND2_X1 U12151 ( .A1(n9634), .A2(n9633), .ZN(n9632) );
  NAND2_X1 U12152 ( .A1(n9760), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9614) );
  MUX2_X1 U12153 ( .A(n11303), .B(P1_REG2_REG_14__SCAN_IN), .S(n10823), .Z(
        n9615) );
  AOI21_X1 U12154 ( .B1(n9632), .B2(n9614), .A(n9615), .ZN(n10816) );
  INV_X1 U12155 ( .A(n9632), .ZN(n9617) );
  NAND2_X1 U12156 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  OAI21_X1 U12157 ( .B1(n9617), .B2(n9616), .A(n14563), .ZN(n9627) );
  NAND2_X1 U12158 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14437)
         );
  OAI21_X1 U12159 ( .B1(n14575), .B2(n15294), .A(n14437), .ZN(n9618) );
  AOI21_X1 U12160 ( .B1(n10823), .B2(n13963), .A(n9618), .ZN(n9626) );
  MUX2_X1 U12161 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n8014), .S(n10823), .Z(
        n9623) );
  NAND2_X1 U12162 ( .A1(n9716), .A2(n7947), .ZN(n9619) );
  NAND2_X1 U12163 ( .A1(n9620), .A2(n9619), .ZN(n9629) );
  INV_X1 U12164 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14503) );
  MUX2_X1 U12165 ( .A(n14503), .B(P1_REG1_REG_13__SCAN_IN), .S(n9760), .Z(
        n9628) );
  NAND2_X1 U12166 ( .A1(n9760), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U12167 ( .A1(n9622), .A2(n9623), .ZN(n10825) );
  OAI21_X1 U12168 ( .B1(n9623), .B2(n9622), .A(n10825), .ZN(n9624) );
  NAND2_X1 U12169 ( .A1(n9624), .A2(n14566), .ZN(n9625) );
  OAI211_X1 U12170 ( .C1(n10816), .C2(n9627), .A(n9626), .B(n9625), .ZN(
        P1_U3257) );
  INV_X1 U12171 ( .A(n9760), .ZN(n9639) );
  AOI21_X1 U12172 ( .B1(n9629), .B2(n9628), .A(n14557), .ZN(n9631) );
  NAND2_X1 U12173 ( .A1(n9631), .A2(n9630), .ZN(n9638) );
  NAND2_X1 U12174 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13798)
         );
  OAI211_X1 U12175 ( .C1(n9634), .C2(n9633), .A(n14563), .B(n9632), .ZN(n9635)
         );
  NAND2_X1 U12176 ( .A1(n13798), .A2(n9635), .ZN(n9636) );
  AOI21_X1 U12177 ( .B1(n14544), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9636), .ZN(
        n9637) );
  OAI211_X1 U12178 ( .C1(n14571), .C2(n9639), .A(n9638), .B(n9637), .ZN(
        P1_U3256) );
  OR2_X1 U12179 ( .A1(n6521), .A2(n9641), .ZN(n9642) );
  NAND2_X1 U12180 ( .A1(n13073), .A2(n9459), .ZN(n9736) );
  XNOR2_X1 U12181 ( .A(n9737), .B(n9736), .ZN(n9739) );
  INV_X1 U12182 ( .A(n9644), .ZN(n9645) );
  XOR2_X1 U12183 ( .A(n9739), .B(n9740), .Z(n9660) );
  NAND2_X1 U12184 ( .A1(n12958), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9654) );
  NAND2_X1 U12185 ( .A1(n12941), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9653) );
  AND2_X1 U12186 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9749) );
  NOR2_X1 U12187 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9648) );
  NOR2_X1 U12188 ( .A1(n9749), .A2(n9648), .ZN(n9920) );
  NAND2_X1 U12189 ( .A1(n12004), .A2(n9920), .ZN(n9652) );
  NAND2_X1 U12190 ( .A1(n12959), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U12191 ( .A1(n13072), .A2(n13407), .ZN(n9656) );
  NAND2_X1 U12192 ( .A1(n13074), .A2(n13405), .ZN(n9655) );
  NAND2_X1 U12193 ( .A1(n9656), .A2(n9655), .ZN(n9881) );
  NOR2_X1 U12194 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9535), .ZN(n14679) );
  AOI21_X1 U12195 ( .B1(n12783), .B2(n9881), .A(n14679), .ZN(n9658) );
  NAND2_X1 U12196 ( .A1(n14657), .A2(n12820), .ZN(n9657) );
  OAI211_X1 U12197 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n14660), .A(n9658), .B(
        n9657), .ZN(n9659) );
  AOI21_X1 U12198 ( .B1(n9660), .B2(n14644), .A(n9659), .ZN(n9661) );
  INV_X1 U12199 ( .A(n9661), .ZN(P2_U3190) );
  NAND2_X1 U12200 ( .A1(n9662), .A2(n9034), .ZN(n9663) );
  NAND2_X1 U12201 ( .A1(n9664), .A2(n9663), .ZN(n9675) );
  INV_X1 U12202 ( .A(n9665), .ZN(n9687) );
  NAND2_X1 U12203 ( .A1(n9687), .A2(n9666), .ZN(n9667) );
  AOI21_X1 U12204 ( .B1(n9732), .B2(n9667), .A(n14873), .ZN(n9674) );
  OAI21_X1 U12205 ( .B1(n9669), .B2(P3_REG1_REG_1__SCAN_IN), .A(n9668), .ZN(
        n9670) );
  NAND2_X1 U12206 ( .A1(n12362), .A2(n9670), .ZN(n9672) );
  NAND2_X1 U12207 ( .A1(n14862), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n9671) );
  OAI211_X1 U12208 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n9998), .A(n9672), .B(
        n9671), .ZN(n9673) );
  AOI211_X1 U12209 ( .C1(n12307), .C2(n9675), .A(n9674), .B(n9673), .ZN(n9676)
         );
  OAI21_X1 U12210 ( .B1(n9677), .B2(n14885), .A(n9676), .ZN(P3_U3183) );
  NOR3_X1 U12211 ( .A1(n12307), .A2(n12362), .A3(n14893), .ZN(n9688) );
  AND2_X1 U12212 ( .A1(n12307), .A2(n9678), .ZN(n9681) );
  OAI22_X1 U12213 ( .A1(n14883), .A2(n9679), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10253), .ZN(n9680) );
  AOI211_X1 U12214 ( .C1(n9682), .C2(n12362), .A(n9681), .B(n9680), .ZN(n9686)
         );
  NAND2_X1 U12215 ( .A1(n9683), .A2(n14893), .ZN(n9684) );
  MUX2_X1 U12216 ( .A(n9684), .B(n14885), .S(P3_IR_REG_0__SCAN_IN), .Z(n9685)
         );
  OAI211_X1 U12217 ( .C1(n9688), .C2(n9687), .A(n9686), .B(n9685), .ZN(
        P3_U3182) );
  INV_X1 U12218 ( .A(n14481), .ZN(n14461) );
  NOR2_X2 U12219 ( .A1(n13808), .A2(n14136), .ZN(n14459) );
  INV_X1 U12220 ( .A(n14459), .ZN(n14470) );
  OAI22_X1 U12221 ( .A1(n10404), .A2(n14470), .B1(n14471), .B2(n10405), .ZN(
        n9689) );
  AOI21_X1 U12222 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n9708), .A(n9689), .ZN(
        n9699) );
  XNOR2_X1 U12223 ( .A(n9690), .B(n13705), .ZN(n9692) );
  NOR2_X1 U12224 ( .A1(n9692), .A2(n9691), .ZN(n9701) );
  NAND2_X1 U12225 ( .A1(n9697), .A2(n14464), .ZN(n9698) );
  OAI211_X1 U12226 ( .C1(n7725), .C2(n14461), .A(n9699), .B(n9698), .ZN(
        P1_U3222) );
  OAI22_X1 U12227 ( .A1(n10405), .A2(n13740), .B1(n14585), .B2(n13741), .ZN(
        n9950) );
  OAI22_X1 U12228 ( .A1(n10405), .A2(n13741), .B1(n14585), .B2(n13739), .ZN(
        n9700) );
  XNOR2_X1 U12229 ( .A(n9700), .B(n13705), .ZN(n9951) );
  XOR2_X1 U12230 ( .A(n9950), .B(n9951), .Z(n9705) );
  INV_X1 U12231 ( .A(n9701), .ZN(n9702) );
  NAND2_X1 U12232 ( .A1(n9703), .A2(n9702), .ZN(n9704) );
  NAND2_X1 U12233 ( .A1(n9704), .A2(n9705), .ZN(n9953) );
  OAI21_X1 U12234 ( .B1(n9705), .B2(n9704), .A(n9953), .ZN(n9706) );
  NAND2_X1 U12235 ( .A1(n9706), .A2(n14464), .ZN(n9710) );
  AOI21_X1 U12236 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n9708), .A(n9707), .ZN(
        n9709) );
  OAI211_X1 U12237 ( .C1(n14585), .C2(n14461), .A(n9710), .B(n9709), .ZN(
        P1_U3237) );
  INV_X1 U12238 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n15218) );
  NAND2_X1 U12239 ( .A1(n12445), .A2(P3_U3897), .ZN(n9711) );
  OAI21_X1 U12240 ( .B1(P3_U3897), .B2(n15218), .A(n9711), .ZN(P3_U3515) );
  OAI21_X1 U12241 ( .B1(n9712), .B2(P2_IR_REG_11__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9713) );
  XNOR2_X1 U12242 ( .A(n9713), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10887) );
  INV_X1 U12243 ( .A(n10887), .ZN(n14739) );
  INV_X1 U12244 ( .A(n10885), .ZN(n9715) );
  INV_X1 U12245 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n15119) );
  OAI222_X1 U12246 ( .A1(P2_U3088), .A2(n14739), .B1(n13578), .B2(n9715), .C1(
        n15119), .C2(n13580), .ZN(P2_U3315) );
  OAI222_X1 U12247 ( .A1(P1_U3086), .A2(n9716), .B1(n14305), .B2(n9715), .C1(
        n9714), .C2(n14302), .ZN(P1_U3343) );
  OAI21_X1 U12248 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9729) );
  OAI21_X1 U12249 ( .B1(n9722), .B2(n9721), .A(n9720), .ZN(n9723) );
  NAND2_X1 U12250 ( .A1(n12362), .A2(n9723), .ZN(n9725) );
  NAND2_X1 U12251 ( .A1(n14862), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n9724) );
  OAI211_X1 U12252 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n14925), .A(n9725), .B(
        n9724), .ZN(n9728) );
  NOR2_X1 U12253 ( .A1(n14885), .A2(n9726), .ZN(n9727) );
  AOI211_X1 U12254 ( .C1(n12307), .C2(n9729), .A(n9728), .B(n9727), .ZN(n9735)
         );
  AND3_X1 U12255 ( .A1(n9732), .A2(n9731), .A3(n9730), .ZN(n9733) );
  OAI21_X1 U12256 ( .B1(n9763), .B2(n9733), .A(n14893), .ZN(n9734) );
  NAND2_X1 U12257 ( .A1(n9735), .A2(n9734), .ZN(P3_U3184) );
  INV_X1 U12258 ( .A(n9736), .ZN(n9738) );
  AND2_X1 U12259 ( .A1(n13072), .A2(n9459), .ZN(n9746) );
  NAND2_X1 U12260 ( .A1(n9741), .A2(n6524), .ZN(n9743) );
  INV_X2 U12261 ( .A(n6521), .ZN(n11862) );
  AOI22_X1 U12262 ( .A1(n11862), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n11861), 
        .B2(n13098), .ZN(n9742) );
  NAND2_X1 U12263 ( .A1(n9743), .A2(n9742), .ZN(n12824) );
  INV_X2 U12264 ( .A(n9744), .ZN(n11976) );
  XNOR2_X1 U12265 ( .A(n12824), .B(n11976), .ZN(n9745) );
  NOR2_X1 U12266 ( .A1(n9745), .A2(n9746), .ZN(n9851) );
  AOI21_X1 U12267 ( .B1(n9746), .B2(n9745), .A(n9851), .ZN(n9747) );
  NAND2_X1 U12268 ( .A1(n9748), .A2(n9747), .ZN(n9853) );
  OAI21_X1 U12269 ( .B1(n9748), .B2(n9747), .A(n9853), .ZN(n9757) );
  INV_X1 U12270 ( .A(n12824), .ZN(n10260) );
  INV_X1 U12271 ( .A(n13073), .ZN(n10118) );
  NAND2_X1 U12272 ( .A1(n12958), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9753) );
  NAND2_X1 U12273 ( .A1(n12941), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U12274 ( .A1(n9749), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9858) );
  OAI21_X1 U12275 ( .B1(n9749), .B2(P2_REG3_REG_5__SCAN_IN), .A(n9858), .ZN(
        n10218) );
  INV_X1 U12276 ( .A(n10218), .ZN(n9867) );
  NAND2_X1 U12277 ( .A1(n12004), .A2(n9867), .ZN(n9751) );
  NAND2_X1 U12278 ( .A1(n12959), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9750) );
  NAND4_X1 U12279 ( .A1(n9753), .A2(n9752), .A3(n9751), .A4(n9750), .ZN(n13071) );
  INV_X1 U12280 ( .A(n13071), .ZN(n10180) );
  INV_X1 U12281 ( .A(n13407), .ZN(n14799) );
  OAI22_X1 U12282 ( .A1(n10118), .A2(n13318), .B1(n10180), .B2(n14799), .ZN(
        n9912) );
  AOI22_X1 U12283 ( .A1(n9912), .A2(n12783), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3088), .ZN(n9755) );
  NAND2_X1 U12284 ( .A1(n12800), .A2(n9920), .ZN(n9754) );
  OAI211_X1 U12285 ( .C1(n10260), .C2(n14415), .A(n9755), .B(n9754), .ZN(n9756) );
  AOI21_X1 U12286 ( .B1(n9757), .B2(n14644), .A(n9756), .ZN(n9758) );
  INV_X1 U12287 ( .A(n9758), .ZN(P2_U3202) );
  INV_X1 U12288 ( .A(n11207), .ZN(n9823) );
  AOI22_X1 U12289 ( .A1(n9760), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9759), .ZN(n9761) );
  OAI21_X1 U12290 ( .B1(n9823), .B2(n14305), .A(n9761), .ZN(P1_U3342) );
  INV_X1 U12291 ( .A(n9826), .ZN(n9765) );
  NOR3_X1 U12292 ( .A1(n9763), .A2(n9762), .A3(n7548), .ZN(n9764) );
  OAI21_X1 U12293 ( .B1(n9765), .B2(n9764), .A(n14893), .ZN(n9773) );
  OAI21_X1 U12294 ( .B1(n9766), .B2(P3_REG2_REG_3__SCAN_IN), .A(n9837), .ZN(
        n9771) );
  AOI21_X1 U12295 ( .B1(n9044), .B2(n9767), .A(n9831), .ZN(n9769) );
  INV_X1 U12296 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10429) );
  NOR2_X1 U12297 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10429), .ZN(n10235) );
  AOI21_X1 U12298 ( .B1(n14862), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10235), .ZN(
        n9768) );
  OAI21_X1 U12299 ( .B1(n14897), .B2(n9769), .A(n9768), .ZN(n9770) );
  AOI21_X1 U12300 ( .B1(n12307), .B2(n9771), .A(n9770), .ZN(n9772) );
  OAI211_X1 U12301 ( .C1(n14885), .C2(n9774), .A(n9773), .B(n9772), .ZN(
        P3_U3185) );
  INV_X1 U12302 ( .A(n9775), .ZN(n9776) );
  OAI222_X1 U12303 ( .A1(P3_U3151), .A2(n12323), .B1(n12698), .B2(n9777), .C1(
        n12694), .C2(n9776), .ZN(P3_U3278) );
  INV_X1 U12304 ( .A(n9788), .ZN(n9784) );
  AND3_X1 U12305 ( .A1(n9780), .A2(n9779), .A3(n9778), .ZN(n9783) );
  INV_X1 U12306 ( .A(n9789), .ZN(n9781) );
  OR2_X1 U12307 ( .A1(n9798), .A2(n9781), .ZN(n9782) );
  OAI211_X1 U12308 ( .C1(n9793), .C2(n9784), .A(n9783), .B(n9782), .ZN(n9785)
         );
  NAND2_X1 U12309 ( .A1(n9785), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9787) );
  OR2_X1 U12310 ( .A1(n9798), .A2(n11835), .ZN(n9786) );
  NOR2_X1 U12311 ( .A1(n12195), .A2(P3_U3151), .ZN(n10108) );
  NAND3_X1 U12312 ( .A1(n9793), .A2(n9788), .A3(n15013), .ZN(n9791) );
  NAND2_X1 U12313 ( .A1(n9798), .A2(n9789), .ZN(n9790) );
  NAND2_X1 U12314 ( .A1(n9791), .A2(n9790), .ZN(n9792) );
  NAND2_X1 U12315 ( .A1(n8921), .A2(n9894), .ZN(n11628) );
  AND2_X1 U12316 ( .A1(n14943), .A2(n11628), .ZN(n11787) );
  INV_X1 U12317 ( .A(n11787), .ZN(n9801) );
  NAND3_X1 U12318 ( .A1(n9793), .A2(n14980), .A3(n9794), .ZN(n9796) );
  NOR2_X1 U12319 ( .A1(n14951), .A2(n15013), .ZN(n9795) );
  INV_X1 U12320 ( .A(n14341), .ZN(n12198) );
  INV_X1 U12321 ( .A(n11835), .ZN(n9797) );
  NAND2_X1 U12322 ( .A1(n9798), .A2(n9797), .ZN(n9994) );
  INV_X1 U12323 ( .A(n9993), .ZN(n9799) );
  OAI22_X1 U12324 ( .A1(n9894), .A2(n12198), .B1(n8522), .B2(n12192), .ZN(
        n9800) );
  AOI21_X1 U12325 ( .B1(n14343), .B2(n9801), .A(n9800), .ZN(n9802) );
  OAI21_X1 U12326 ( .B1(n10108), .B2(n10253), .A(n9802), .ZN(P3_U3172) );
  INV_X1 U12327 ( .A(n9803), .ZN(n9806) );
  NOR3_X1 U12328 ( .A1(n9828), .A2(n9804), .A3(n7547), .ZN(n9805) );
  OAI21_X1 U12329 ( .B1(n9806), .B2(n9805), .A(n14893), .ZN(n9818) );
  OAI21_X1 U12330 ( .B1(n9808), .B2(P3_REG2_REG_5__SCAN_IN), .A(n9807), .ZN(
        n9816) );
  AND2_X1 U12331 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n10539) );
  INV_X1 U12332 ( .A(n10539), .ZN(n9809) );
  OAI21_X1 U12333 ( .B1(n14883), .B2(n7562), .A(n9809), .ZN(n9815) );
  AOI21_X1 U12334 ( .B1(n9053), .B2(n9811), .A(n9810), .ZN(n9812) );
  OAI22_X1 U12335 ( .A1(n9813), .A2(n14885), .B1(n9812), .B2(n14897), .ZN(
        n9814) );
  AOI211_X1 U12336 ( .C1(n12307), .C2(n9816), .A(n9815), .B(n9814), .ZN(n9817)
         );
  NAND2_X1 U12337 ( .A1(n9818), .A2(n9817), .ZN(P3_U3187) );
  NAND2_X1 U12338 ( .A1(n9819), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9820) );
  MUX2_X1 U12339 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9820), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9821) );
  AND2_X1 U12340 ( .A1(n9821), .A2(n10076), .ZN(n14751) );
  INV_X1 U12341 ( .A(n14751), .ZN(n10092) );
  OAI222_X1 U12342 ( .A1(P2_U3088), .A2(n10092), .B1(n13578), .B2(n9823), .C1(
        n9822), .C2(n13580), .ZN(P2_U3314) );
  AND3_X1 U12343 ( .A1(n9826), .A2(n9825), .A3(n9824), .ZN(n9827) );
  OAI21_X1 U12344 ( .B1(n9828), .B2(n9827), .A(n14893), .ZN(n9844) );
  OR3_X1 U12345 ( .A1(n9831), .A2(n9830), .A3(n9829), .ZN(n9832) );
  AOI21_X1 U12346 ( .B1(n9833), .B2(n9832), .A(n14897), .ZN(n9842) );
  INV_X1 U12347 ( .A(n9834), .ZN(n9836) );
  NAND3_X1 U12348 ( .A1(n9837), .A2(n9836), .A3(n9835), .ZN(n9838) );
  AOI21_X1 U12349 ( .B1(n9839), .B2(n9838), .A(n14903), .ZN(n9841) );
  NOR2_X1 U12350 ( .A1(n14883), .A2(n15082), .ZN(n9840) );
  AND2_X1 U12351 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10334) );
  NOR4_X1 U12352 ( .A1(n9842), .A2(n9841), .A3(n9840), .A4(n10334), .ZN(n9843)
         );
  OAI211_X1 U12353 ( .C1(n14885), .C2(n7060), .A(n9844), .B(n9843), .ZN(
        P3_U3186) );
  AND2_X1 U12354 ( .A1(n13071), .A2(n6520), .ZN(n9850) );
  OR2_X1 U12355 ( .A1(n9845), .A2(n11375), .ZN(n9848) );
  AOI22_X1 U12356 ( .A1(n11862), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n11861), 
        .B2(n9846), .ZN(n9847) );
  NAND2_X1 U12357 ( .A1(n9848), .A2(n9847), .ZN(n12834) );
  XNOR2_X1 U12358 ( .A(n12834), .B(n11976), .ZN(n9849) );
  NOR2_X1 U12359 ( .A1(n9849), .A2(n9850), .ZN(n9964) );
  AOI21_X1 U12360 ( .B1(n9850), .B2(n9849), .A(n9964), .ZN(n9855) );
  INV_X1 U12361 ( .A(n9851), .ZN(n9852) );
  NAND2_X1 U12362 ( .A1(n9853), .A2(n9852), .ZN(n9854) );
  OAI21_X1 U12363 ( .B1(n9855), .B2(n9854), .A(n9966), .ZN(n9856) );
  NAND2_X1 U12364 ( .A1(n9856), .A2(n14644), .ZN(n9869) );
  NAND2_X1 U12365 ( .A1(n12958), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U12366 ( .A1(n12941), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9862) );
  AND2_X1 U12367 ( .A1(n9858), .A2(n9857), .ZN(n9859) );
  NOR2_X1 U12368 ( .A1(n9971), .A2(n9859), .ZN(n10184) );
  NAND2_X1 U12369 ( .A1(n12004), .A2(n10184), .ZN(n9861) );
  NAND2_X1 U12370 ( .A1(n12959), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9860) );
  NAND4_X1 U12371 ( .A1(n9863), .A2(n9862), .A3(n9861), .A4(n9860), .ZN(n13070) );
  INV_X1 U12372 ( .A(n13070), .ZN(n10522) );
  OAI21_X1 U12373 ( .B1(n14419), .B2(n10522), .A(n9864), .ZN(n9866) );
  INV_X1 U12374 ( .A(n13072), .ZN(n10206) );
  OAI22_X1 U12375 ( .A1(n7205), .A2(n14415), .B1(n14418), .B2(n10206), .ZN(
        n9865) );
  AOI211_X1 U12376 ( .C1(n9867), .C2(n12800), .A(n9866), .B(n9865), .ZN(n9868)
         );
  NAND2_X1 U12377 ( .A1(n9869), .A2(n9868), .ZN(P2_U3199) );
  NAND2_X1 U12378 ( .A1(n13075), .A2(n9348), .ZN(n9870) );
  INV_X1 U12379 ( .A(n9871), .ZN(n9938) );
  NAND2_X1 U12380 ( .A1(n14800), .A2(n9348), .ZN(n9872) );
  INV_X1 U12381 ( .A(n13006), .ZN(n10114) );
  INV_X1 U12382 ( .A(n13074), .ZN(n9934) );
  INV_X1 U12383 ( .A(n6534), .ZN(n14829) );
  NAND2_X1 U12384 ( .A1(n9934), .A2(n14829), .ZN(n9873) );
  NAND2_X1 U12385 ( .A1(n10113), .A2(n9873), .ZN(n9874) );
  NAND2_X1 U12386 ( .A1(n9874), .A2(n13008), .ZN(n9899) );
  OAI21_X1 U12387 ( .B1(n9874), .B2(n13008), .A(n9899), .ZN(n10166) );
  INV_X1 U12388 ( .A(n10166), .ZN(n9884) );
  OR2_X1 U12389 ( .A1(n9333), .A2(n13412), .ZN(n14802) );
  INV_X1 U12390 ( .A(n14802), .ZN(n9876) );
  NAND2_X1 U12391 ( .A1(n9876), .A2(n12968), .ZN(n14822) );
  INV_X1 U12392 ( .A(n13005), .ZN(n9933) );
  NAND2_X1 U12393 ( .A1(n9932), .A2(n9877), .ZN(n10116) );
  NAND2_X1 U12394 ( .A1(n10116), .A2(n13006), .ZN(n10117) );
  NAND2_X1 U12395 ( .A1(n9934), .A2(n6534), .ZN(n9878) );
  NAND2_X1 U12396 ( .A1(n10117), .A2(n9878), .ZN(n9909) );
  XNOR2_X1 U12397 ( .A(n9909), .B(n9908), .ZN(n9882) );
  NAND2_X1 U12398 ( .A1(n13048), .A2(n9333), .ZN(n9880) );
  OR2_X1 U12399 ( .A1(n13412), .A2(n12968), .ZN(n9879) );
  NAND2_X2 U12400 ( .A1(n9880), .A2(n9879), .ZN(n14798) );
  AOI21_X1 U12401 ( .B1(n9882), .B2(n14798), .A(n9881), .ZN(n10161) );
  OR2_X1 U12402 ( .A1(n9381), .A2(n9883), .ZN(n10122) );
  OAI211_X1 U12403 ( .C1(n10125), .C2(n6522), .A(n10803), .B(n9915), .ZN(
        n10164) );
  OAI211_X1 U12404 ( .C1(n9884), .C2(n13529), .A(n10161), .B(n10164), .ZN(
        n10270) );
  INV_X1 U12405 ( .A(n14817), .ZN(n14820) );
  OR2_X1 U12406 ( .A1(n9885), .A2(n14820), .ZN(n14818) );
  NAND3_X1 U12407 ( .A1(n9887), .A2(n9886), .A3(n9903), .ZN(n9888) );
  INV_X1 U12408 ( .A(n14816), .ZN(n9889) );
  NAND2_X1 U12409 ( .A1(n14861), .A2(n14843), .ZN(n13502) );
  OAI22_X1 U12410 ( .A1(n13502), .A2(n6522), .B1(n14861), .B2(n9231), .ZN(
        n9890) );
  AOI21_X1 U12411 ( .B1(n10270), .B2(n14861), .A(n9890), .ZN(n9891) );
  INV_X1 U12412 ( .A(n9891), .ZN(P2_U3502) );
  NOR3_X1 U12413 ( .A1(n11787), .A2(n14980), .A3(n9892), .ZN(n9893) );
  AOI21_X1 U12414 ( .B1(n14944), .B2(n6823), .A(n9893), .ZN(n10257) );
  OAI22_X1 U12415 ( .A1(n12612), .A2(n9894), .B1(n15031), .B2(n8523), .ZN(
        n9895) );
  INV_X1 U12416 ( .A(n9895), .ZN(n9896) );
  OAI21_X1 U12417 ( .B1(n10257), .B2(n15029), .A(n9896), .ZN(P3_U3459) );
  INV_X1 U12418 ( .A(n12669), .ZN(n12664) );
  AOI22_X1 U12419 ( .A1(n12664), .A2(n10255), .B1(n15018), .B2(
        P3_REG0_REG_0__SCAN_IN), .ZN(n9897) );
  OAI21_X1 U12420 ( .B1(n10257), .B2(n15018), .A(n9897), .ZN(P3_U3390) );
  NAND2_X1 U12421 ( .A1(n10118), .A2(n6522), .ZN(n9898) );
  NAND2_X1 U12422 ( .A1(n9899), .A2(n9898), .ZN(n9901) );
  XNOR2_X1 U12423 ( .A(n13072), .B(n12824), .ZN(n13010) );
  INV_X1 U12424 ( .A(n13010), .ZN(n9900) );
  NAND2_X1 U12425 ( .A1(n9901), .A2(n9900), .ZN(n10179) );
  OAI21_X1 U12426 ( .B1(n9901), .B2(n9900), .A(n10179), .ZN(n9902) );
  INV_X1 U12427 ( .A(n9902), .ZN(n10001) );
  AND3_X1 U12428 ( .A1(n14817), .A2(n9904), .A3(n9903), .ZN(n9905) );
  NAND2_X1 U12429 ( .A1(n14816), .A2(n9905), .ZN(n9917) );
  INV_X1 U12430 ( .A(n12807), .ZN(n9906) );
  NAND2_X1 U12431 ( .A1(n9906), .A2(n10205), .ZN(n9907) );
  NAND2_X1 U12432 ( .A1(n9909), .A2(n9908), .ZN(n9911) );
  NAND2_X1 U12433 ( .A1(n10118), .A2(n12820), .ZN(n9910) );
  AOI21_X1 U12434 ( .B1(n9913), .B2(n14798), .A(n9912), .ZN(n10000) );
  MUX2_X1 U12435 ( .A(n9914), .B(n10000), .S(n14809), .Z(n9925) );
  AOI21_X1 U12436 ( .B1(n9915), .B2(n12824), .A(n9459), .ZN(n9916) );
  NAND2_X1 U12437 ( .A1(n9916), .A2(n10215), .ZN(n9999) );
  INV_X1 U12438 ( .A(n9999), .ZN(n9923) );
  INV_X1 U12439 ( .A(n13412), .ZN(n13052) );
  INV_X1 U12440 ( .A(n9918), .ZN(n9919) );
  INV_X1 U12441 ( .A(n9920), .ZN(n9921) );
  OAI22_X1 U12442 ( .A1(n13390), .A2(n10260), .B1(n14803), .B2(n9921), .ZN(
        n9922) );
  AOI21_X1 U12443 ( .B1(n9923), .B2(n13425), .A(n9922), .ZN(n9924) );
  OAI211_X1 U12444 ( .C1(n10001), .C2(n13396), .A(n9925), .B(n9924), .ZN(
        P2_U3261) );
  INV_X1 U12445 ( .A(n12347), .ZN(n9929) );
  INV_X1 U12446 ( .A(n9926), .ZN(n9927) );
  OAI222_X1 U12447 ( .A1(P3_U3151), .A2(n9929), .B1(n12698), .B2(n9928), .C1(
        n12694), .C2(n9927), .ZN(P3_U3277) );
  OAI222_X1 U12448 ( .A1(P3_U3151), .A2(n6525), .B1(n12694), .B2(n9931), .C1(
        n9930), .C2(n12698), .ZN(P3_U3276) );
  OAI21_X1 U12449 ( .B1(n13007), .B2(n9933), .A(n9932), .ZN(n9941) );
  OAI22_X1 U12450 ( .A1(n9935), .A2(n13318), .B1(n9934), .B2(n14799), .ZN(
        n9940) );
  INV_X1 U12451 ( .A(n9936), .ZN(n9937) );
  AOI21_X1 U12452 ( .B1(n13007), .B2(n9938), .A(n9937), .ZN(n10006) );
  NOR2_X1 U12453 ( .A1(n10006), .A2(n10205), .ZN(n9939) );
  AOI211_X1 U12454 ( .C1(n14798), .C2(n9941), .A(n9940), .B(n9939), .ZN(n10005) );
  INV_X2 U12455 ( .A(n14809), .ZN(n14811) );
  OAI211_X1 U12456 ( .C1(n9348), .C2(n14797), .A(n10803), .B(n10122), .ZN(
        n10004) );
  INV_X1 U12457 ( .A(n10004), .ZN(n9942) );
  INV_X1 U12458 ( .A(n14803), .ZN(n14783) );
  AOI22_X1 U12459 ( .A1(n9942), .A2(n13425), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n14783), .ZN(n9943) );
  OAI21_X1 U12460 ( .B1(n13083), .B2(n14809), .A(n9943), .ZN(n9945) );
  NAND2_X1 U12461 ( .A1(n14809), .A2(n12807), .ZN(n14805) );
  NOR2_X1 U12462 ( .A1(n10006), .A2(n14805), .ZN(n9944) );
  AOI211_X1 U12463 ( .C1(n14785), .C2(n9381), .A(n9945), .B(n9944), .ZN(n9946)
         );
  OAI21_X1 U12464 ( .B1(n10005), .B2(n14811), .A(n9946), .ZN(P2_U3264) );
  NAND2_X1 U12465 ( .A1(n13857), .A2(n10605), .ZN(n9948) );
  INV_X2 U12466 ( .A(n13739), .ZN(n13702) );
  NAND2_X1 U12467 ( .A1(n13702), .A2(n10388), .ZN(n9947) );
  NAND2_X1 U12468 ( .A1(n9948), .A2(n9947), .ZN(n9949) );
  XNOR2_X1 U12469 ( .A(n9949), .B(n13705), .ZN(n10192) );
  INV_X1 U12470 ( .A(n10388), .ZN(n14591) );
  OAI22_X1 U12471 ( .A1(n10365), .A2(n13740), .B1(n14591), .B2(n13741), .ZN(
        n10191) );
  XNOR2_X1 U12472 ( .A(n10192), .B(n10191), .ZN(n9957) );
  INV_X1 U12473 ( .A(n10194), .ZN(n9955) );
  AOI211_X1 U12474 ( .C1(n9957), .C2(n9956), .A(n14476), .B(n9955), .ZN(n9963)
         );
  INV_X1 U12475 ( .A(n14485), .ZN(n13835) );
  AOI22_X1 U12476 ( .A1(n9959), .A2(n13835), .B1(n14481), .B2(n10388), .ZN(
        n9961) );
  INV_X1 U12477 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9959) );
  NOR2_X1 U12478 ( .A1(n9959), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13901) );
  AOI21_X1 U12479 ( .B1(n14457), .B2(n13855), .A(n13901), .ZN(n9960) );
  OAI211_X1 U12480 ( .C1(n10405), .C2(n14470), .A(n9961), .B(n9960), .ZN(n9962) );
  OR2_X1 U12481 ( .A1(n9963), .A2(n9962), .ZN(P1_U3218) );
  INV_X1 U12482 ( .A(n9964), .ZN(n9965) );
  NAND2_X1 U12483 ( .A1(n13070), .A2(n6520), .ZN(n10056) );
  OR2_X1 U12484 ( .A1(n9967), .A2(n11375), .ZN(n9969) );
  AOI22_X1 U12485 ( .A1(n11862), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n11861), 
        .B2(n14690), .ZN(n9968) );
  NAND2_X1 U12486 ( .A1(n9969), .A2(n9968), .ZN(n14835) );
  XNOR2_X1 U12487 ( .A(n14835), .B(n11976), .ZN(n10055) );
  XOR2_X1 U12488 ( .A(n10056), .B(n10055), .Z(n10058) );
  XNOR2_X1 U12489 ( .A(n10059), .B(n10058), .ZN(n9980) );
  NAND2_X1 U12490 ( .A1(n12958), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U12491 ( .A1(n12941), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9975) );
  NAND2_X1 U12492 ( .A1(n9971), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10064) );
  OR2_X1 U12493 ( .A1(n9971), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9972) );
  AND2_X1 U12494 ( .A1(n10064), .A2(n9972), .ZN(n14784) );
  NAND2_X1 U12495 ( .A1(n12004), .A2(n14784), .ZN(n9974) );
  NAND2_X1 U12496 ( .A1(n12959), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9973) );
  NAND4_X1 U12497 ( .A1(n9976), .A2(n9975), .A3(n9974), .A4(n9973), .ZN(n13069) );
  INV_X1 U12498 ( .A(n13069), .ZN(n10649) );
  AOI22_X1 U12499 ( .A1(n12801), .A2(n13071), .B1(n12800), .B2(n10184), .ZN(
        n9977) );
  NAND2_X1 U12500 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14699) );
  OAI211_X1 U12501 ( .C1(n10649), .C2(n14419), .A(n9977), .B(n14699), .ZN(
        n9978) );
  AOI21_X1 U12502 ( .B1(n14835), .B2(n14657), .A(n9978), .ZN(n9979) );
  OAI21_X1 U12503 ( .B1(n9980), .B2(n14652), .A(n9979), .ZN(P2_U3211) );
  NAND2_X1 U12504 ( .A1(n12199), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n9981) );
  OAI21_X1 U12505 ( .B1(n11782), .B2(n12199), .A(n9981), .ZN(P3_U3521) );
  NAND2_X1 U12506 ( .A1(n12199), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n9982) );
  OAI21_X1 U12507 ( .B1(n12370), .B2(n12199), .A(n9982), .ZN(P3_U3520) );
  INV_X1 U12508 ( .A(n11819), .ZN(n9984) );
  NAND2_X1 U12509 ( .A1(n12674), .A2(n9984), .ZN(n9986) );
  MUX2_X1 U12510 ( .A(n9983), .B(n8923), .S(n12095), .Z(n9991) );
  INV_X1 U12511 ( .A(n9990), .ZN(n14942) );
  AOI21_X1 U12512 ( .B1(n9987), .B2(n12095), .A(n14942), .ZN(n9988) );
  NAND2_X1 U12513 ( .A1(n9991), .A2(n9988), .ZN(n10101) );
  NAND3_X1 U12514 ( .A1(n9983), .A2(n14943), .A3(n12095), .ZN(n9989) );
  OAI211_X1 U12515 ( .C1(n9991), .C2(n9990), .A(n10101), .B(n9989), .ZN(n9992)
         );
  NAND2_X1 U12516 ( .A1(n9992), .A2(n14343), .ZN(n9997) );
  OR2_X1 U12517 ( .A1(n9994), .A2(n9993), .ZN(n14336) );
  INV_X1 U12518 ( .A(n14336), .ZN(n12190) );
  OAI22_X1 U12519 ( .A1(n14941), .A2(n12198), .B1(n10425), .B2(n12192), .ZN(
        n9995) );
  AOI21_X1 U12520 ( .B1(n12190), .B2(n8921), .A(n9995), .ZN(n9996) );
  OAI211_X1 U12521 ( .C1(n10108), .C2(n9998), .A(n9997), .B(n9996), .ZN(
        P3_U3162) );
  OAI211_X1 U12522 ( .C1(n10001), .C2(n13529), .A(n10000), .B(n9999), .ZN(
        n10262) );
  OAI22_X1 U12523 ( .A1(n13502), .A2(n10260), .B1(n14861), .B2(n9232), .ZN(
        n10002) );
  AOI21_X1 U12524 ( .B1(n10262), .B2(n14861), .A(n10002), .ZN(n10003) );
  INV_X1 U12525 ( .A(n10003), .ZN(P2_U3503) );
  OAI211_X1 U12526 ( .C1(n10006), .C2(n14822), .A(n10005), .B(n10004), .ZN(
        n10266) );
  OAI22_X1 U12527 ( .A1(n13502), .A2(n9348), .B1(n14861), .B2(n9227), .ZN(
        n10007) );
  AOI21_X1 U12528 ( .B1(n10266), .B2(n14861), .A(n10007), .ZN(n10008) );
  INV_X1 U12529 ( .A(n10008), .ZN(P2_U3500) );
  NAND2_X1 U12530 ( .A1(n10011), .A2(n10010), .ZN(n10358) );
  NAND2_X1 U12531 ( .A1(n10405), .A2(n14585), .ZN(n10013) );
  NAND2_X1 U12532 ( .A1(n10014), .A2(n10013), .ZN(n10377) );
  INV_X1 U12533 ( .A(n10379), .ZN(n10015) );
  NAND2_X1 U12534 ( .A1(n10365), .A2(n14591), .ZN(n10016) );
  NAND2_X1 U12535 ( .A1(n10017), .A2(n10016), .ZN(n10446) );
  XOR2_X1 U12536 ( .A(n10446), .B(n10023), .Z(n10399) );
  INV_X1 U12537 ( .A(n10018), .ZN(n10019) );
  NAND2_X1 U12538 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  NAND2_X1 U12539 ( .A1(n10365), .A2(n10388), .ZN(n10022) );
  NAND2_X1 U12540 ( .A1(n10378), .A2(n10022), .ZN(n10455) );
  XOR2_X1 U12541 ( .A(n10023), .B(n10455), .Z(n10024) );
  AOI222_X1 U12542 ( .A1(n14264), .A2(n10024), .B1(n13854), .B2(n14152), .C1(
        n13857), .C2(n14154), .ZN(n10391) );
  OR2_X1 U12543 ( .A1(n10415), .A2(n10400), .ZN(n10402) );
  NAND2_X1 U12544 ( .A1(n10456), .A2(n10385), .ZN(n10025) );
  AND2_X1 U12545 ( .A1(n10575), .A2(n10025), .ZN(n10393) );
  INV_X1 U12546 ( .A(n9590), .ZN(n14618) );
  AOI22_X1 U12547 ( .A1(n10393), .A2(n14618), .B1(n14617), .B2(n10456), .ZN(
        n10026) );
  OAI211_X1 U12548 ( .C1(n14623), .C2(n10399), .A(n10391), .B(n10026), .ZN(
        n10028) );
  NAND2_X1 U12549 ( .A1(n10028), .A2(n14636), .ZN(n10027) );
  OAI21_X1 U12550 ( .B1(n14636), .B2(n9418), .A(n10027), .ZN(P1_U3532) );
  INV_X1 U12551 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10030) );
  NAND2_X1 U12552 ( .A1(n10028), .A2(n14627), .ZN(n10029) );
  OAI21_X1 U12553 ( .B1(n14627), .B2(n10030), .A(n10029), .ZN(P1_U3471) );
  AOI21_X1 U12554 ( .B1(n10034), .B2(n10032), .A(n10132), .ZN(n10054) );
  INV_X1 U12555 ( .A(n10033), .ZN(n10040) );
  MUX2_X1 U12556 ( .A(n10035), .B(n10034), .S(n12691), .Z(n10036) );
  NAND2_X1 U12557 ( .A1(n10036), .A2(n10147), .ZN(n10143) );
  INV_X1 U12558 ( .A(n10036), .ZN(n10037) );
  NAND2_X1 U12559 ( .A1(n10037), .A2(n10049), .ZN(n10038) );
  AND2_X1 U12560 ( .A1(n10143), .A2(n10038), .ZN(n10039) );
  OAI21_X1 U12561 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(n10144) );
  INV_X1 U12562 ( .A(n10144), .ZN(n10043) );
  NOR3_X1 U12563 ( .A1(n10041), .A2(n10040), .A3(n10039), .ZN(n10042) );
  OAI21_X1 U12564 ( .B1(n10043), .B2(n10042), .A(n14893), .ZN(n10053) );
  AOI21_X1 U12565 ( .B1(n10035), .B2(n10046), .A(n10148), .ZN(n10047) );
  INV_X1 U12566 ( .A(n10047), .ZN(n10051) );
  AND2_X1 U12567 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10861) );
  AOI21_X1 U12568 ( .B1(n14862), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n10861), .ZN(
        n10048) );
  OAI21_X1 U12569 ( .B1(n14885), .B2(n10049), .A(n10048), .ZN(n10050) );
  AOI21_X1 U12570 ( .B1(n10051), .B2(n12307), .A(n10050), .ZN(n10052) );
  OAI211_X1 U12571 ( .C1(n10054), .C2(n14897), .A(n10053), .B(n10052), .ZN(
        P3_U3189) );
  INV_X1 U12572 ( .A(n10055), .ZN(n10057) );
  OR2_X1 U12573 ( .A1(n10060), .A2(n11375), .ZN(n10063) );
  AOI22_X1 U12574 ( .A1(n11862), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11861), 
        .B2(n10061), .ZN(n10062) );
  NAND2_X1 U12575 ( .A1(n10063), .A2(n10062), .ZN(n14786) );
  XNOR2_X1 U12576 ( .A(n14786), .B(n11976), .ZN(n10280) );
  NAND2_X1 U12577 ( .A1(n13069), .A2(n6520), .ZN(n10279) );
  XNOR2_X1 U12578 ( .A(n10280), .B(n10279), .ZN(n10282) );
  XNOR2_X1 U12579 ( .A(n10283), .B(n10282), .ZN(n10075) );
  INV_X1 U12580 ( .A(n14784), .ZN(n10072) );
  NAND2_X1 U12581 ( .A1(n12958), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U12582 ( .A1(n12941), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10068) );
  NAND2_X1 U12583 ( .A1(n10064), .A2(n10296), .ZN(n10065) );
  AND2_X1 U12584 ( .A1(n10290), .A2(n10065), .ZN(n10693) );
  NAND2_X1 U12585 ( .A1(n12004), .A2(n10693), .ZN(n10067) );
  NAND2_X1 U12586 ( .A1(n12959), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n10066) );
  NAND4_X1 U12587 ( .A1(n10069), .A2(n10068), .A3(n10067), .A4(n10066), .ZN(
        n13068) );
  INV_X1 U12588 ( .A(n13068), .ZN(n10770) );
  OAI22_X1 U12589 ( .A1(n10522), .A2(n13318), .B1(n10770), .B2(n14799), .ZN(
        n10525) );
  NAND2_X1 U12590 ( .A1(n10525), .A2(n12783), .ZN(n10071) );
  OAI211_X1 U12591 ( .C1(n14660), .C2(n10072), .A(n10071), .B(n10070), .ZN(
        n10073) );
  AOI21_X1 U12592 ( .B1(n14786), .B2(n14657), .A(n10073), .ZN(n10074) );
  OAI21_X1 U12593 ( .B1(n10075), .B2(n14652), .A(n10074), .ZN(P2_U3185) );
  INV_X1 U12594 ( .A(n10823), .ZN(n10818) );
  OAI222_X1 U12595 ( .A1(P1_U3086), .A2(n10818), .B1(n14305), .B2(n11376), 
        .C1(n15126), .C2(n14302), .ZN(P1_U3341) );
  NAND2_X1 U12596 ( .A1(n10076), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10077) );
  XNOR2_X1 U12597 ( .A(n10077), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11377) );
  INV_X1 U12598 ( .A(n11377), .ZN(n10931) );
  OAI222_X1 U12599 ( .A1(n13580), .A2(n10078), .B1(n13574), .B2(n11376), .C1(
        n10931), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U12600 ( .A(n11516), .ZN(n10082) );
  NAND2_X1 U12601 ( .A1(n10302), .A2(n10079), .ZN(n10241) );
  NAND2_X1 U12602 ( .A1(n10241), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10080) );
  XNOR2_X1 U12603 ( .A(n10080), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11517) );
  INV_X1 U12604 ( .A(n11517), .ZN(n11179) );
  OAI222_X1 U12605 ( .A1(n13580), .A2(n10081), .B1(n13574), .B2(n10082), .C1(
        n11179), .C2(P2_U3088), .ZN(P2_U3311) );
  OAI222_X1 U12606 ( .A1(P1_U3086), .A2(n10822), .B1(n14305), .B2(n10082), 
        .C1(n15244), .C2(n14302), .ZN(P1_U3339) );
  INV_X1 U12607 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15206) );
  AOI22_X1 U12608 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n14739), .B1(n10887), 
        .B2(n15206), .ZN(n14734) );
  INV_X1 U12609 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15083) );
  OAI21_X1 U12610 ( .B1(n9293), .B2(n10086), .A(n10083), .ZN(n14726) );
  MUX2_X1 U12611 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n15083), .S(n10748), .Z(
        n14725) );
  NAND2_X1 U12612 ( .A1(n14726), .A2(n14725), .ZN(n14724) );
  OAI21_X1 U12613 ( .B1(n15083), .B2(n14721), .A(n14724), .ZN(n14735) );
  NOR2_X1 U12614 ( .A1(n14734), .A2(n14735), .ZN(n14733) );
  INV_X1 U12615 ( .A(n14733), .ZN(n10084) );
  OAI21_X1 U12616 ( .B1(n10887), .B2(P2_REG1_REG_12__SCAN_IN), .A(n10084), 
        .ZN(n14748) );
  XNOR2_X1 U12617 ( .A(n14751), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n14749) );
  NOR2_X1 U12618 ( .A1(n14748), .A2(n14749), .ZN(n14746) );
  AOI21_X1 U12619 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n14751), .A(n14746), 
        .ZN(n10934) );
  XNOR2_X1 U12620 ( .A(n11377), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n10933) );
  XNOR2_X1 U12621 ( .A(n10934), .B(n10933), .ZN(n10098) );
  NAND2_X1 U12622 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14424)
         );
  NOR2_X1 U12623 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n10887), .ZN(n10089) );
  INV_X1 U12624 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10087) );
  OAI21_X1 U12625 ( .B1(n9300), .B2(n10086), .A(n10085), .ZN(n14719) );
  MUX2_X1 U12626 ( .A(n10087), .B(P2_REG2_REG_11__SCAN_IN), .S(n10748), .Z(
        n14718) );
  NOR2_X1 U12627 ( .A1(n14719), .A2(n14718), .ZN(n14717) );
  AOI21_X1 U12628 ( .B1(n10087), .B2(n14721), .A(n14717), .ZN(n14732) );
  INV_X1 U12629 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10088) );
  AOI22_X1 U12630 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n14739), .B1(n10887), 
        .B2(n10088), .ZN(n14731) );
  NOR2_X1 U12631 ( .A1(n14732), .A2(n14731), .ZN(n14730) );
  NOR2_X1 U12632 ( .A1(n14753), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10093) );
  INV_X1 U12633 ( .A(n14753), .ZN(n10091) );
  INV_X1 U12634 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10090) );
  OAI22_X1 U12635 ( .A1(n10093), .A2(n10092), .B1(n10091), .B2(n10090), .ZN(
        n10924) );
  XNOR2_X1 U12636 ( .A(n10931), .B(n10924), .ZN(n10094) );
  NAND2_X1 U12637 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10094), .ZN(n10925) );
  OAI211_X1 U12638 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n10094), .A(n14776), 
        .B(n10925), .ZN(n10095) );
  AND2_X1 U12639 ( .A1(n14424), .A2(n10095), .ZN(n10097) );
  AOI22_X1 U12640 ( .A1(n14768), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(n14770), 
        .B2(n11377), .ZN(n10096) );
  OAI211_X1 U12641 ( .C1(n10098), .C2(n14747), .A(n10097), .B(n10096), .ZN(
        P2_U3228) );
  INV_X2 U12642 ( .A(n12095), .ZN(n12046) );
  XNOR2_X1 U12643 ( .A(n14924), .B(n12046), .ZN(n10230) );
  XNOR2_X1 U12644 ( .A(n10230), .B(n14945), .ZN(n10103) );
  XNOR2_X1 U12645 ( .A(n14941), .B(n12046), .ZN(n10099) );
  NAND2_X1 U12646 ( .A1(n8522), .A2(n10099), .ZN(n10100) );
  NAND2_X1 U12647 ( .A1(n10101), .A2(n10100), .ZN(n10102) );
  NAND2_X1 U12648 ( .A1(n10104), .A2(n14343), .ZN(n10107) );
  INV_X1 U12649 ( .A(n14911), .ZN(n14931) );
  OAI22_X1 U12650 ( .A1(n12198), .A2(n14924), .B1(n14931), .B2(n12192), .ZN(
        n10105) );
  AOI21_X1 U12651 ( .B1(n12190), .B2(n6823), .A(n10105), .ZN(n10106) );
  OAI211_X1 U12652 ( .C1(n10108), .C2(n14925), .A(n10107), .B(n10106), .ZN(
        P3_U3177) );
  INV_X1 U12653 ( .A(n10109), .ZN(n10111) );
  OAI222_X1 U12654 ( .A1(n12698), .A2(n10112), .B1(n12694), .B2(n10111), .C1(
        n10110), .C2(P3_U3151), .ZN(P3_U3275) );
  OAI21_X1 U12655 ( .B1(n10115), .B2(n10114), .A(n10113), .ZN(n14832) );
  INV_X1 U12656 ( .A(n14832), .ZN(n10130) );
  OAI21_X1 U12657 ( .B1(n10116), .B2(n13006), .A(n10117), .ZN(n10120) );
  OAI22_X1 U12658 ( .A1(n14800), .A2(n13318), .B1(n10118), .B2(n14799), .ZN(
        n10119) );
  AOI21_X1 U12659 ( .B1(n10120), .B2(n14798), .A(n10119), .ZN(n10121) );
  OAI21_X1 U12660 ( .B1(n10130), .B2(n10205), .A(n10121), .ZN(n14830) );
  NAND2_X1 U12661 ( .A1(n14830), .A2(n14809), .ZN(n10129) );
  NAND2_X1 U12662 ( .A1(n10122), .A2(n6534), .ZN(n10123) );
  NAND2_X1 U12663 ( .A1(n10123), .A2(n10803), .ZN(n10124) );
  OR2_X1 U12664 ( .A1(n10125), .A2(n10124), .ZN(n14828) );
  AOI22_X1 U12665 ( .A1(n14811), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n14783), .ZN(n10126) );
  OAI21_X1 U12666 ( .B1(n14789), .B2(n14828), .A(n10126), .ZN(n10127) );
  AOI21_X1 U12667 ( .B1(n14785), .B2(n6534), .A(n10127), .ZN(n10128) );
  OAI211_X1 U12668 ( .C1(n10130), .C2(n14805), .A(n10129), .B(n10128), .ZN(
        P2_U3263) );
  NAND2_X1 U12669 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10487), .ZN(n10133) );
  OAI21_X1 U12670 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10487), .A(n10133), .ZN(
        n10134) );
  AOI21_X1 U12671 ( .B1(n10135), .B2(n10134), .A(n10486), .ZN(n10160) );
  MUX2_X1 U12672 ( .A(n10137), .B(n10136), .S(n12691), .Z(n10139) );
  INV_X1 U12673 ( .A(n10487), .ZN(n10138) );
  NAND2_X1 U12674 ( .A1(n10139), .A2(n10138), .ZN(n10471) );
  INV_X1 U12675 ( .A(n10139), .ZN(n10140) );
  NAND2_X1 U12676 ( .A1(n10140), .A2(n10487), .ZN(n10141) );
  NAND2_X1 U12677 ( .A1(n10471), .A2(n10141), .ZN(n10142) );
  AOI21_X1 U12678 ( .B1(n10144), .B2(n10143), .A(n10142), .ZN(n10479) );
  AND3_X1 U12679 ( .A1(n10144), .A2(n10143), .A3(n10142), .ZN(n10145) );
  OAI21_X1 U12680 ( .B1(n10479), .B2(n10145), .A(n14893), .ZN(n10159) );
  NOR2_X1 U12681 ( .A1(n10147), .A2(n10146), .ZN(n10149) );
  NAND2_X1 U12682 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10487), .ZN(n10150) );
  OAI21_X1 U12683 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10487), .A(n10150), .ZN(
        n10151) );
  AOI21_X1 U12684 ( .B1(n10152), .B2(n10151), .A(n10484), .ZN(n10153) );
  INV_X1 U12685 ( .A(n10153), .ZN(n10157) );
  NOR2_X1 U12686 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10154), .ZN(n11037) );
  AOI21_X1 U12687 ( .B1(n14862), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11037), .ZN(
        n10155) );
  OAI21_X1 U12688 ( .B1(n14885), .B2(n10487), .A(n10155), .ZN(n10156) );
  AOI21_X1 U12689 ( .B1(n10157), .B2(n12307), .A(n10156), .ZN(n10158) );
  OAI211_X1 U12690 ( .C1(n10160), .C2(n14897), .A(n10159), .B(n10158), .ZN(
        P3_U3190) );
  MUX2_X1 U12691 ( .A(n10162), .B(n10161), .S(n14809), .Z(n10168) );
  AOI22_X1 U12692 ( .A1(n14785), .A2(n12820), .B1(n9535), .B2(n14783), .ZN(
        n10163) );
  OAI21_X1 U12693 ( .B1(n14789), .B2(n10164), .A(n10163), .ZN(n10165) );
  AOI21_X1 U12694 ( .B1(n10166), .B2(n14792), .A(n10165), .ZN(n10167) );
  NAND2_X1 U12695 ( .A1(n10168), .A2(n10167), .ZN(P2_U3262) );
  NAND2_X1 U12696 ( .A1(n10206), .A2(n12824), .ZN(n10207) );
  NAND2_X1 U12697 ( .A1(n10209), .A2(n10207), .ZN(n10169) );
  XNOR2_X1 U12698 ( .A(n12834), .B(n13071), .ZN(n13011) );
  NAND2_X1 U12699 ( .A1(n10169), .A2(n13011), .ZN(n10171) );
  NAND2_X1 U12700 ( .A1(n12834), .A2(n10180), .ZN(n10172) );
  NAND2_X1 U12701 ( .A1(n10171), .A2(n10172), .ZN(n10170) );
  XNOR2_X1 U12702 ( .A(n14835), .B(n13070), .ZN(n13012) );
  INV_X1 U12703 ( .A(n13012), .ZN(n10517) );
  NAND3_X1 U12704 ( .A1(n10171), .A2(n10517), .A3(n10172), .ZN(n10173) );
  NAND2_X1 U12705 ( .A1(n10524), .A2(n10173), .ZN(n10174) );
  NAND2_X1 U12706 ( .A1(n10174), .A2(n14798), .ZN(n10176) );
  AOI22_X1 U12707 ( .A1(n13405), .A2(n13071), .B1(n13069), .B2(n13407), .ZN(
        n10175) );
  AND2_X1 U12708 ( .A1(n10176), .A2(n10175), .ZN(n14841) );
  MUX2_X1 U12709 ( .A(n10177), .B(n14841), .S(n14809), .Z(n10188) );
  NAND2_X1 U12710 ( .A1(n10260), .A2(n10206), .ZN(n10178) );
  NAND2_X1 U12711 ( .A1(n10179), .A2(n10178), .ZN(n10204) );
  INV_X1 U12712 ( .A(n13011), .ZN(n10208) );
  NAND2_X1 U12713 ( .A1(n10204), .A2(n10208), .ZN(n10203) );
  NAND2_X1 U12714 ( .A1(n7205), .A2(n10180), .ZN(n10181) );
  XNOR2_X1 U12715 ( .A(n10518), .B(n10517), .ZN(n14834) );
  NAND2_X1 U12716 ( .A1(n10217), .A2(n14835), .ZN(n10182) );
  NAND2_X1 U12717 ( .A1(n10182), .A2(n10803), .ZN(n10183) );
  OR2_X1 U12718 ( .A1(n10183), .A2(n10527), .ZN(n14836) );
  AOI22_X1 U12719 ( .A1(n14835), .A2(n14785), .B1(n14783), .B2(n10184), .ZN(
        n10185) );
  OAI21_X1 U12720 ( .B1(n14836), .B2(n14789), .A(n10185), .ZN(n10186) );
  AOI21_X1 U12721 ( .B1(n14834), .B2(n14792), .A(n10186), .ZN(n10187) );
  NAND2_X1 U12722 ( .A1(n10188), .A2(n10187), .ZN(P2_U3259) );
  INV_X1 U12723 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n15108) );
  INV_X1 U12724 ( .A(n12387), .ZN(n10189) );
  NAND2_X1 U12725 ( .A1(n10189), .A2(P3_U3897), .ZN(n10190) );
  OAI21_X1 U12726 ( .B1(P3_U3897), .B2(n15108), .A(n10190), .ZN(P3_U3519) );
  OR2_X1 U12727 ( .A1(n13740), .A2(n10585), .ZN(n10196) );
  OR2_X1 U12728 ( .A1(n10453), .A2(n13741), .ZN(n10195) );
  NAND2_X1 U12729 ( .A1(n10196), .A2(n10195), .ZN(n10337) );
  OR2_X1 U12730 ( .A1(n10453), .A2(n13739), .ZN(n10197) );
  OAI21_X1 U12731 ( .B1(n10585), .B2(n13741), .A(n10197), .ZN(n10198) );
  XNOR2_X1 U12732 ( .A(n10198), .B(n13705), .ZN(n10338) );
  XNOR2_X1 U12733 ( .A(n10339), .B(n10338), .ZN(n10202) );
  INV_X1 U12734 ( .A(n13854), .ZN(n10459) );
  NAND2_X1 U12735 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13906) );
  OAI21_X1 U12736 ( .B1(n14471), .B2(n10459), .A(n13906), .ZN(n10200) );
  OAI22_X1 U12737 ( .A1(n14461), .A2(n10453), .B1(n10395), .B2(n14485), .ZN(
        n10199) );
  AOI211_X1 U12738 ( .C1(n14459), .C2(n13857), .A(n10200), .B(n10199), .ZN(
        n10201) );
  OAI21_X1 U12739 ( .B1(n10202), .B2(n14476), .A(n10201), .ZN(P1_U3230) );
  OAI21_X1 U12740 ( .B1(n10204), .B2(n10208), .A(n10203), .ZN(n10213) );
  INV_X1 U12741 ( .A(n10213), .ZN(n10225) );
  INV_X1 U12742 ( .A(n10205), .ZN(n14847) );
  OAI22_X1 U12743 ( .A1(n10206), .A2(n13318), .B1(n10522), .B2(n14799), .ZN(
        n10212) );
  NAND3_X1 U12744 ( .A1(n10209), .A2(n10208), .A3(n10207), .ZN(n10210) );
  INV_X1 U12745 ( .A(n14798), .ZN(n13369) );
  AOI21_X1 U12746 ( .B1(n10171), .B2(n10210), .A(n13369), .ZN(n10211) );
  AOI211_X1 U12747 ( .C1(n14847), .C2(n10213), .A(n10212), .B(n10211), .ZN(
        n10224) );
  MUX2_X1 U12748 ( .A(n10214), .B(n10224), .S(n14809), .Z(n10221) );
  AOI21_X1 U12749 ( .B1(n10215), .B2(n12834), .A(n9459), .ZN(n10216) );
  AND2_X1 U12750 ( .A1(n10217), .A2(n10216), .ZN(n10222) );
  OAI22_X1 U12751 ( .A1(n7205), .A2(n13390), .B1(n14803), .B2(n10218), .ZN(
        n10219) );
  AOI21_X1 U12752 ( .B1(n10222), .B2(n13425), .A(n10219), .ZN(n10220) );
  OAI211_X1 U12753 ( .C1(n10225), .C2(n14805), .A(n10221), .B(n10220), .ZN(
        P2_U3260) );
  INV_X1 U12754 ( .A(n10222), .ZN(n10223) );
  OAI211_X1 U12755 ( .C1(n10225), .C2(n14822), .A(n10224), .B(n10223), .ZN(
        n10274) );
  OAI22_X1 U12756 ( .A1(n13502), .A2(n7205), .B1(n14861), .B2(n10226), .ZN(
        n10227) );
  AOI21_X1 U12757 ( .B1(n10274), .B2(n14861), .A(n10227), .ZN(n10228) );
  INV_X1 U12758 ( .A(n10228), .ZN(P2_U3504) );
  XNOR2_X1 U12759 ( .A(n10320), .B(n14911), .ZN(n10232) );
  NAND2_X1 U12760 ( .A1(n10425), .A2(n10230), .ZN(n10233) );
  AND2_X1 U12761 ( .A1(n10232), .A2(n10233), .ZN(n10231) );
  INV_X1 U12762 ( .A(n10330), .ZN(n10326) );
  NOR3_X1 U12763 ( .A1(n10326), .A2(n10234), .A3(n12174), .ZN(n10239) );
  INV_X1 U12764 ( .A(n12192), .ZN(n14333) );
  AOI22_X1 U12765 ( .A1(n12190), .A2(n14945), .B1(n14333), .B2(n12206), .ZN(
        n10237) );
  AOI21_X1 U12766 ( .B1(n14341), .B2(n14971), .A(n10235), .ZN(n10236) );
  OAI211_X1 U12767 ( .C1(n14347), .C2(P3_REG3_REG_3__SCAN_IN), .A(n10237), .B(
        n10236), .ZN(n10238) );
  OR2_X1 U12768 ( .A1(n10239), .A2(n10238), .ZN(P3_U3158) );
  INV_X1 U12769 ( .A(n11547), .ZN(n10245) );
  INV_X1 U12770 ( .A(n11273), .ZN(n11282) );
  OAI222_X1 U12771 ( .A1(n14302), .A2(n10240), .B1(n14305), .B2(n10245), .C1(
        P1_U3086), .C2(n11282), .ZN(P1_U3338) );
  OAI21_X1 U12772 ( .B1(n10241), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10242) );
  MUX2_X1 U12773 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10242), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n10243) );
  AND2_X1 U12774 ( .A1(n10243), .A2(n10637), .ZN(n14769) );
  INV_X1 U12775 ( .A(n14769), .ZN(n11175) );
  OAI222_X1 U12776 ( .A1(P2_U3088), .A2(n11175), .B1(n13574), .B2(n10245), 
        .C1(n10244), .C2(n13580), .ZN(P2_U3310) );
  NAND2_X1 U12777 ( .A1(n12672), .A2(n10246), .ZN(n10247) );
  OAI21_X1 U12778 ( .B1(n12672), .B2(n10248), .A(n10247), .ZN(n10249) );
  INV_X1 U12779 ( .A(n10249), .ZN(n10250) );
  NAND2_X1 U12780 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  INV_X1 U12781 ( .A(n14951), .ZN(n14927) );
  OR2_X1 U12782 ( .A1(n10252), .A2(n14927), .ZN(n11053) );
  OAI22_X1 U12783 ( .A1(n14955), .A2(n15155), .B1(n10253), .B2(n14926), .ZN(
        n10254) );
  AOI21_X1 U12784 ( .B1(n14919), .B2(n10255), .A(n10254), .ZN(n10256) );
  OAI21_X1 U12785 ( .B1(n10257), .B2(n14957), .A(n10256), .ZN(P3_U3233) );
  AND2_X2 U12786 ( .A1(n10258), .A2(n14816), .ZN(n14855) );
  NAND2_X1 U12787 ( .A1(n14855), .A2(n14843), .ZN(n13556) );
  INV_X1 U12788 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10259) );
  OAI22_X1 U12789 ( .A1(n13556), .A2(n10260), .B1(n14855), .B2(n10259), .ZN(
        n10261) );
  AOI21_X1 U12790 ( .B1(n10262), .B2(n14855), .A(n10261), .ZN(n10263) );
  INV_X1 U12791 ( .A(n10263), .ZN(P2_U3442) );
  INV_X1 U12792 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10264) );
  OAI22_X1 U12793 ( .A1(n13556), .A2(n9348), .B1(n14855), .B2(n10264), .ZN(
        n10265) );
  AOI21_X1 U12794 ( .B1(n10266), .B2(n14855), .A(n10265), .ZN(n10267) );
  INV_X1 U12795 ( .A(n10267), .ZN(P2_U3433) );
  INV_X1 U12796 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10268) );
  OAI22_X1 U12797 ( .A1(n13556), .A2(n6522), .B1(n14855), .B2(n10268), .ZN(
        n10269) );
  AOI21_X1 U12798 ( .B1(n10270), .B2(n14855), .A(n10269), .ZN(n10271) );
  INV_X1 U12799 ( .A(n10271), .ZN(P2_U3439) );
  INV_X1 U12800 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10272) );
  OAI22_X1 U12801 ( .A1(n13556), .A2(n7205), .B1(n14855), .B2(n10272), .ZN(
        n10273) );
  AOI21_X1 U12802 ( .B1(n10274), .B2(n14855), .A(n10273), .ZN(n10275) );
  INV_X1 U12803 ( .A(n10275), .ZN(P2_U3445) );
  OR2_X1 U12804 ( .A1(n10276), .A2(n11375), .ZN(n10278) );
  AOI22_X1 U12805 ( .A1(n11862), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n11861), 
        .B2(n13114), .ZN(n10277) );
  NAND2_X1 U12806 ( .A1(n10278), .A2(n10277), .ZN(n12857) );
  INV_X1 U12807 ( .A(n12857), .ZN(n10655) );
  INV_X1 U12808 ( .A(n10279), .ZN(n10281) );
  AND2_X1 U12809 ( .A1(n13068), .A2(n6520), .ZN(n10285) );
  XNOR2_X1 U12810 ( .A(n12857), .B(n11976), .ZN(n10284) );
  NOR2_X1 U12811 ( .A1(n10284), .A2(n10285), .ZN(n10502) );
  AOI21_X1 U12812 ( .B1(n10285), .B2(n10284), .A(n10502), .ZN(n10286) );
  NAND2_X1 U12813 ( .A1(n10287), .A2(n10286), .ZN(n10504) );
  OAI21_X1 U12814 ( .B1(n10287), .B2(n10286), .A(n10504), .ZN(n10288) );
  NAND2_X1 U12815 ( .A1(n10288), .A2(n14644), .ZN(n10299) );
  NAND2_X1 U12816 ( .A1(n11977), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10295) );
  NAND2_X1 U12817 ( .A1(n12958), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10294) );
  INV_X1 U12818 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10289) );
  AND2_X1 U12819 ( .A1(n10290), .A2(n10289), .ZN(n10291) );
  NOR2_X1 U12820 ( .A1(n10508), .A2(n10291), .ZN(n13420) );
  NAND2_X1 U12821 ( .A1(n12004), .A2(n13420), .ZN(n10293) );
  NAND2_X1 U12822 ( .A1(n12959), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n10292) );
  NAND4_X1 U12823 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n13067) );
  AOI22_X1 U12824 ( .A1(n13405), .A2(n13069), .B1(n13067), .B2(n13407), .ZN(
        n10651) );
  INV_X1 U12825 ( .A(n12783), .ZN(n14649) );
  OAI22_X1 U12826 ( .A1(n10651), .A2(n14649), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10296), .ZN(n10297) );
  AOI21_X1 U12827 ( .B1(n10693), .B2(n12800), .A(n10297), .ZN(n10298) );
  OAI211_X1 U12828 ( .C1(n10655), .C2(n14415), .A(n10299), .B(n10298), .ZN(
        P2_U3193) );
  INV_X1 U12829 ( .A(n11383), .ZN(n10304) );
  OAI222_X1 U12830 ( .A1(n14554), .A2(P1_U3086), .B1(n14305), .B2(n10304), 
        .C1(n10300), .C2(n14302), .ZN(P1_U3340) );
  OR2_X1 U12831 ( .A1(n10302), .A2(n10301), .ZN(n10303) );
  XNOR2_X1 U12832 ( .A(n10303), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14759) );
  INV_X1 U12833 ( .A(n14759), .ZN(n10936) );
  OAI222_X1 U12834 ( .A1(n13580), .A2(n10305), .B1(n13574), .B2(n10304), .C1(
        P2_U3088), .C2(n10936), .ZN(P2_U3312) );
  INV_X2 U12835 ( .A(n14076), .ZN(n14159) );
  OAI22_X1 U12836 ( .A1(n14159), .A2(n10310), .B1(n10309), .B2(n14106), .ZN(
        n10314) );
  NOR2_X2 U12837 ( .A1(n13989), .A2(n6669), .ZN(n14167) );
  AOI21_X1 U12838 ( .B1(n14112), .B2(n14161), .A(n10312), .ZN(n10313) );
  AOI211_X1 U12839 ( .C1(n14159), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10314), .B(
        n10313), .ZN(n10319) );
  NAND2_X1 U12840 ( .A1(n14076), .A2(n14264), .ZN(n14116) );
  INV_X1 U12841 ( .A(n14116), .ZN(n11484) );
  INV_X1 U12842 ( .A(n10315), .ZN(n10316) );
  OAI21_X1 U12843 ( .B1(n11484), .B2(n14114), .A(n10317), .ZN(n10318) );
  NAND2_X1 U12844 ( .A1(n10319), .A2(n10318), .ZN(P1_U3293) );
  INV_X1 U12845 ( .A(n10320), .ZN(n10321) );
  AND2_X1 U12846 ( .A1(n10321), .A2(n14911), .ZN(n10327) );
  INV_X1 U12847 ( .A(n12206), .ZN(n10424) );
  XNOR2_X1 U12848 ( .A(n10322), .B(n12046), .ZN(n10323) );
  NAND2_X1 U12849 ( .A1(n10424), .A2(n10323), .ZN(n10535) );
  INV_X1 U12850 ( .A(n10323), .ZN(n10324) );
  NAND2_X1 U12851 ( .A1(n10324), .A2(n12206), .ZN(n10325) );
  NAND2_X1 U12852 ( .A1(n10535), .A2(n10325), .ZN(n10328) );
  OAI21_X1 U12853 ( .B1(n10326), .B2(n10327), .A(n10328), .ZN(n10331) );
  NOR2_X1 U12854 ( .A1(n10328), .A2(n10327), .ZN(n10329) );
  NAND2_X1 U12855 ( .A1(n10330), .A2(n10329), .ZN(n10536) );
  AOI21_X1 U12856 ( .B1(n10331), .B2(n10536), .A(n12174), .ZN(n10332) );
  INV_X1 U12857 ( .A(n10332), .ZN(n10336) );
  INV_X1 U12858 ( .A(n14910), .ZN(n10909) );
  OAI22_X1 U12859 ( .A1(n14931), .A2(n14336), .B1(n10909), .B2(n12192), .ZN(
        n10333) );
  AOI211_X1 U12860 ( .C1(n14973), .C2(n14341), .A(n10334), .B(n10333), .ZN(
        n10335) );
  OAI211_X1 U12861 ( .C1(n14921), .C2(n14347), .A(n10336), .B(n10335), .ZN(
        P3_U3170) );
  NAND2_X1 U12862 ( .A1(n10579), .A2(n13702), .ZN(n10341) );
  NAND2_X1 U12863 ( .A1(n13854), .A2(n13697), .ZN(n10340) );
  NAND2_X1 U12864 ( .A1(n10341), .A2(n10340), .ZN(n10342) );
  XNOR2_X1 U12865 ( .A(n10342), .B(n13705), .ZN(n10347) );
  NAND2_X1 U12866 ( .A1(n10579), .A2(n13697), .ZN(n10345) );
  NAND2_X1 U12867 ( .A1(n10343), .A2(n13854), .ZN(n10344) );
  NAND2_X1 U12868 ( .A1(n10345), .A2(n10344), .ZN(n10346) );
  NOR2_X1 U12869 ( .A1(n10347), .A2(n10346), .ZN(n10601) );
  INV_X1 U12870 ( .A(n10601), .ZN(n10348) );
  NAND2_X1 U12871 ( .A1(n10347), .A2(n10346), .ZN(n10600) );
  NAND2_X1 U12872 ( .A1(n10348), .A2(n10600), .ZN(n10349) );
  XNOR2_X1 U12873 ( .A(n10602), .B(n10349), .ZN(n10354) );
  INV_X1 U12874 ( .A(n13853), .ZN(n10606) );
  OAI21_X1 U12875 ( .B1(n14471), .B2(n10606), .A(n10350), .ZN(n10351) );
  AOI21_X1 U12876 ( .B1(n14459), .B2(n13855), .A(n10351), .ZN(n10353) );
  AOI22_X1 U12877 ( .A1(n13835), .A2(n10578), .B1(n14481), .B2(n10579), .ZN(
        n10352) );
  OAI211_X1 U12878 ( .C1(n10354), .C2(n14476), .A(n10353), .B(n10352), .ZN(
        P1_U3227) );
  INV_X1 U12879 ( .A(n10355), .ZN(n10357) );
  OAI222_X1 U12880 ( .A1(n12694), .A2(n10357), .B1(n12698), .B2(n10356), .C1(
        P3_U3151), .C2(n10418), .ZN(P3_U3274) );
  CLKBUF_X1 U12881 ( .A(n10358), .Z(n10359) );
  XNOR2_X1 U12882 ( .A(n10359), .B(n10364), .ZN(n14584) );
  INV_X1 U12883 ( .A(n10360), .ZN(n10361) );
  NAND2_X1 U12884 ( .A1(n14076), .A2(n10361), .ZN(n14019) );
  OAI21_X1 U12885 ( .B1(n10364), .B2(n10363), .A(n10362), .ZN(n10367) );
  AOI21_X1 U12886 ( .B1(n10367), .B2(n14264), .A(n10366), .ZN(n10368) );
  OAI21_X1 U12887 ( .B1(n14584), .B2(n14010), .A(n10368), .ZN(n14587) );
  NAND2_X1 U12888 ( .A1(n14587), .A2(n14076), .ZN(n10376) );
  AND2_X1 U12889 ( .A1(n10402), .A2(n10374), .ZN(n10369) );
  OR2_X1 U12890 ( .A1(n10369), .A2(n10386), .ZN(n14586) );
  INV_X1 U12891 ( .A(n14586), .ZN(n10370) );
  NAND2_X1 U12892 ( .A1(n14167), .A2(n10370), .ZN(n10372) );
  INV_X1 U12893 ( .A(n14106), .ZN(n14157) );
  NAND2_X1 U12894 ( .A1(n14157), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n10371) );
  OAI211_X1 U12895 ( .C1(n9394), .C2(n14076), .A(n10372), .B(n10371), .ZN(
        n10373) );
  AOI21_X1 U12896 ( .B1(n14110), .B2(n10374), .A(n10373), .ZN(n10375) );
  OAI211_X1 U12897 ( .C1(n14584), .C2(n14019), .A(n10376), .B(n10375), .ZN(
        P1_U3291) );
  XNOR2_X1 U12898 ( .A(n10377), .B(n10379), .ZN(n14590) );
  OAI21_X1 U12899 ( .B1(n10380), .B2(n10379), .A(n10378), .ZN(n10383) );
  OAI22_X1 U12900 ( .A1(n10585), .A2(n14138), .B1(n10405), .B2(n14136), .ZN(
        n10382) );
  NOR2_X1 U12901 ( .A1(n14590), .A2(n14010), .ZN(n10381) );
  AOI211_X1 U12902 ( .C1(n14264), .C2(n10383), .A(n10382), .B(n10381), .ZN(
        n14593) );
  MUX2_X1 U12903 ( .A(n10384), .B(n14593), .S(n14076), .Z(n10390) );
  OAI21_X1 U12904 ( .B1(n10386), .B2(n14591), .A(n10385), .ZN(n14592) );
  OAI22_X1 U12905 ( .A1(n14112), .A2(n14592), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14106), .ZN(n10387) );
  AOI21_X1 U12906 ( .B1(n14110), .B2(n10388), .A(n10387), .ZN(n10389) );
  OAI211_X1 U12907 ( .C1(n14590), .C2(n14019), .A(n10390), .B(n10389), .ZN(
        P1_U3290) );
  MUX2_X1 U12908 ( .A(n10392), .B(n10391), .S(n14076), .Z(n10398) );
  NAND2_X1 U12909 ( .A1(n14167), .A2(n10393), .ZN(n10394) );
  OAI21_X1 U12910 ( .B1(n14106), .B2(n10395), .A(n10394), .ZN(n10396) );
  AOI21_X1 U12911 ( .B1(n14110), .B2(n10456), .A(n10396), .ZN(n10397) );
  OAI211_X1 U12912 ( .C1(n14164), .C2(n10399), .A(n10398), .B(n10397), .ZN(
        P1_U3289) );
  NAND2_X1 U12913 ( .A1(n10415), .A2(n10400), .ZN(n10401) );
  NAND2_X1 U12914 ( .A1(n10402), .A2(n10401), .ZN(n14579) );
  XNOR2_X1 U12915 ( .A(n13859), .B(n14579), .ZN(n10403) );
  MUX2_X1 U12916 ( .A(n10009), .B(n10403), .S(n10404), .Z(n10409) );
  OAI22_X1 U12917 ( .A1(n10405), .A2(n14138), .B1(n10404), .B2(n14136), .ZN(
        n10408) );
  XOR2_X1 U12918 ( .A(n10009), .B(n10406), .Z(n10414) );
  NOR2_X1 U12919 ( .A1(n10414), .A2(n14010), .ZN(n10407) );
  AOI211_X1 U12920 ( .C1(n14264), .C2(n10409), .A(n10408), .B(n10407), .ZN(
        n14580) );
  INV_X1 U12921 ( .A(n14579), .ZN(n10413) );
  NOR2_X1 U12922 ( .A1(n14106), .A2(n10410), .ZN(n10412) );
  NOR2_X1 U12923 ( .A1(n14076), .A2(n9395), .ZN(n10411) );
  AOI211_X1 U12924 ( .C1(n10413), .C2(n14167), .A(n10412), .B(n10411), .ZN(
        n10417) );
  INV_X1 U12925 ( .A(n14019), .ZN(n14064) );
  INV_X1 U12926 ( .A(n10414), .ZN(n14583) );
  AOI22_X1 U12927 ( .A1(n14064), .A2(n14583), .B1(n14110), .B2(n10415), .ZN(
        n10416) );
  OAI211_X1 U12928 ( .C1(n14580), .C2(n14159), .A(n10417), .B(n10416), .ZN(
        P1_U3292) );
  NOR2_X1 U12929 ( .A1(n14951), .A2(n10418), .ZN(n14939) );
  NAND2_X1 U12930 ( .A1(n14955), .A2(n14939), .ZN(n10971) );
  NAND2_X1 U12931 ( .A1(n14955), .A2(n14978), .ZN(n10419) );
  INV_X1 U12932 ( .A(n14380), .ZN(n11437) );
  XNOR2_X1 U12933 ( .A(n10420), .B(n10421), .ZN(n14966) );
  INV_X1 U12934 ( .A(n10422), .ZN(n10423) );
  NOR2_X1 U12935 ( .A1(n10423), .A2(n11788), .ZN(n14907) );
  AOI211_X1 U12936 ( .C1(n11788), .C2(n10423), .A(n14949), .B(n14907), .ZN(
        n10427) );
  OAI22_X1 U12937 ( .A1(n10425), .A2(n14932), .B1(n10424), .B2(n14930), .ZN(
        n10426) );
  NOR2_X1 U12938 ( .A1(n10427), .A2(n10426), .ZN(n14968) );
  MUX2_X1 U12939 ( .A(n10428), .B(n14968), .S(n14955), .Z(n10431) );
  AOI22_X1 U12940 ( .A1(n14919), .A2(n14971), .B1(n14952), .B2(n10429), .ZN(
        n10430) );
  OAI211_X1 U12941 ( .C1(n11437), .C2(n14966), .A(n10431), .B(n10430), .ZN(
        P3_U3230) );
  XNOR2_X1 U12942 ( .A(n10432), .B(n11793), .ZN(n14979) );
  INV_X1 U12943 ( .A(n14979), .ZN(n10442) );
  OAI21_X1 U12944 ( .B1(n6676), .B2(n10434), .A(n6795), .ZN(n10435) );
  NAND2_X1 U12945 ( .A1(n10435), .A2(n14934), .ZN(n10437) );
  AOI22_X1 U12946 ( .A1(n14946), .A2(n12206), .B1(n12205), .B2(n14944), .ZN(
        n10436) );
  AND2_X1 U12947 ( .A1(n10437), .A2(n10436), .ZN(n14985) );
  MUX2_X1 U12948 ( .A(n14985), .B(n10438), .S(n14957), .Z(n10441) );
  INV_X1 U12949 ( .A(n10542), .ZN(n10439) );
  AOI22_X1 U12950 ( .A1(n14919), .A2(n14981), .B1(n14952), .B2(n10439), .ZN(
        n10440) );
  OAI211_X1 U12951 ( .C1(n11437), .C2(n10442), .A(n10441), .B(n10440), .ZN(
        P3_U3228) );
  INV_X1 U12952 ( .A(n14219), .ZN(n14608) );
  INV_X1 U12953 ( .A(n10443), .ZN(n10444) );
  INV_X1 U12954 ( .A(n10571), .ZN(n10448) );
  NAND2_X1 U12955 ( .A1(n10448), .A2(n10447), .ZN(n10573) );
  INV_X1 U12956 ( .A(n10579), .ZN(n14598) );
  NAND2_X1 U12957 ( .A1(n14598), .A2(n10459), .ZN(n10449) );
  INV_X1 U12958 ( .A(n10546), .ZN(n10450) );
  OAI21_X1 U12959 ( .B1(n10451), .B2(n10450), .A(n10553), .ZN(n10598) );
  INV_X1 U12960 ( .A(n10612), .ZN(n10603) );
  NOR2_X1 U12961 ( .A1(n10574), .A2(n10603), .ZN(n10452) );
  OR2_X1 U12962 ( .A1(n10561), .A2(n10452), .ZN(n10594) );
  OAI22_X1 U12963 ( .A1(n10594), .A2(n9590), .B1(n10603), .B2(n14609), .ZN(
        n10467) );
  NAND2_X1 U12964 ( .A1(n13855), .A2(n10453), .ZN(n10454) );
  NAND2_X1 U12965 ( .A1(n10455), .A2(n10454), .ZN(n10458) );
  NAND2_X1 U12966 ( .A1(n10456), .A2(n10585), .ZN(n10457) );
  NAND2_X1 U12967 ( .A1(n10458), .A2(n10457), .ZN(n10582) );
  NAND2_X1 U12968 ( .A1(n10582), .A2(n10581), .ZN(n10461) );
  NAND2_X1 U12969 ( .A1(n10579), .A2(n10459), .ZN(n10460) );
  NAND2_X1 U12970 ( .A1(n10461), .A2(n10460), .ZN(n10547) );
  XNOR2_X1 U12971 ( .A(n10547), .B(n10546), .ZN(n10462) );
  NAND2_X1 U12972 ( .A1(n10462), .A2(n14264), .ZN(n10466) );
  NAND2_X1 U12973 ( .A1(n13854), .A2(n14154), .ZN(n10464) );
  NAND2_X1 U12974 ( .A1(n13852), .A2(n14152), .ZN(n10463) );
  AND2_X1 U12975 ( .A1(n10464), .A2(n10463), .ZN(n10610) );
  INV_X1 U12976 ( .A(n14010), .ZN(n14057) );
  NAND2_X1 U12977 ( .A1(n10598), .A2(n14057), .ZN(n10465) );
  NAND3_X1 U12978 ( .A1(n10466), .A2(n10610), .A3(n10465), .ZN(n10595) );
  AOI211_X1 U12979 ( .C1(n14608), .C2(n10598), .A(n10467), .B(n10595), .ZN(
        n10469) );
  OR2_X1 U12980 ( .A1(n10469), .A2(n14625), .ZN(n10468) );
  OAI21_X1 U12981 ( .B1(n14627), .B2(n7820), .A(n10468), .ZN(P1_U3477) );
  OR2_X1 U12982 ( .A1(n10469), .A2(n14634), .ZN(n10470) );
  OAI21_X1 U12983 ( .B1(n14636), .B2(n7818), .A(n10470), .ZN(P1_U3534) );
  INV_X1 U12984 ( .A(n10471), .ZN(n10478) );
  MUX2_X1 U12985 ( .A(n10473), .B(n10472), .S(n12691), .Z(n10474) );
  NAND2_X1 U12986 ( .A1(n10474), .A2(n10708), .ZN(n10722) );
  INV_X1 U12987 ( .A(n10474), .ZN(n10475) );
  NAND2_X1 U12988 ( .A1(n10475), .A2(n10488), .ZN(n10476) );
  AND2_X1 U12989 ( .A1(n10722), .A2(n10476), .ZN(n10477) );
  OAI21_X1 U12990 ( .B1(n10479), .B2(n10478), .A(n10477), .ZN(n10723) );
  INV_X1 U12991 ( .A(n10723), .ZN(n10481) );
  NOR3_X1 U12992 ( .A1(n10479), .A2(n10478), .A3(n10477), .ZN(n10480) );
  OAI21_X1 U12993 ( .B1(n10481), .B2(n10480), .A(n14893), .ZN(n10483) );
  AND2_X1 U12994 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n10852) );
  AOI21_X1 U12995 ( .B1(n14862), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10852), .ZN(
        n10482) );
  OAI211_X1 U12996 ( .C1(n14885), .C2(n10488), .A(n10483), .B(n10482), .ZN(
        n10493) );
  AOI21_X1 U12997 ( .B1(n10473), .B2(n10485), .A(n10709), .ZN(n10491) );
  AOI21_X1 U12998 ( .B1(n10472), .B2(n10489), .A(n10702), .ZN(n10490) );
  OAI22_X1 U12999 ( .A1(n10491), .A2(n14903), .B1(n10490), .B2(n14897), .ZN(
        n10492) );
  OR2_X1 U13000 ( .A1(n10493), .A2(n10492), .ZN(P3_U3191) );
  OR2_X1 U13001 ( .A1(n10494), .A2(n11375), .ZN(n10499) );
  OAI22_X1 U13002 ( .A1(n6521), .A2(n10496), .B1(n14705), .B2(n10495), .ZN(
        n10497) );
  INV_X1 U13003 ( .A(n10497), .ZN(n10498) );
  INV_X1 U13004 ( .A(n13424), .ZN(n10812) );
  AND2_X1 U13005 ( .A1(n13067), .A2(n6520), .ZN(n10501) );
  XNOR2_X1 U13006 ( .A(n13424), .B(n11976), .ZN(n10500) );
  NOR2_X1 U13007 ( .A1(n10500), .A2(n10501), .ZN(n10731) );
  AOI21_X1 U13008 ( .B1(n10501), .B2(n10500), .A(n10731), .ZN(n10506) );
  INV_X1 U13009 ( .A(n10502), .ZN(n10503) );
  NAND2_X1 U13010 ( .A1(n10504), .A2(n10503), .ZN(n10505) );
  NAND2_X1 U13011 ( .A1(n10505), .A2(n10506), .ZN(n10733) );
  OAI21_X1 U13012 ( .B1(n10506), .B2(n10505), .A(n10733), .ZN(n10507) );
  NAND2_X1 U13013 ( .A1(n10507), .A2(n14644), .ZN(n10516) );
  NOR2_X1 U13014 ( .A1(n10508), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10509) );
  OR2_X1 U13015 ( .A1(n10741), .A2(n10509), .ZN(n14647) );
  INV_X1 U13016 ( .A(n14647), .ZN(n10778) );
  NAND2_X1 U13017 ( .A1(n12004), .A2(n10778), .ZN(n10513) );
  NAND2_X1 U13018 ( .A1(n12958), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10512) );
  NAND2_X1 U13019 ( .A1(n12959), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U13020 ( .A1(n12941), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10510) );
  NAND4_X1 U13021 ( .A1(n10513), .A2(n10512), .A3(n10511), .A4(n10510), .ZN(
        n13066) );
  AOI22_X1 U13022 ( .A1(n13405), .A2(n13068), .B1(n13066), .B2(n13407), .ZN(
        n10808) );
  NAND2_X1 U13023 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14714) );
  OAI21_X1 U13024 ( .B1(n10808), .B2(n14649), .A(n14714), .ZN(n10514) );
  AOI21_X1 U13025 ( .B1(n13420), .B2(n12800), .A(n10514), .ZN(n10515) );
  OAI211_X1 U13026 ( .C1(n10812), .C2(n14415), .A(n10516), .B(n10515), .ZN(
        P2_U3203) );
  NAND2_X1 U13027 ( .A1(n10518), .A2(n10517), .ZN(n10520) );
  OR2_X1 U13028 ( .A1(n14835), .A2(n13070), .ZN(n10519) );
  NAND2_X1 U13029 ( .A1(n10520), .A2(n10519), .ZN(n10521) );
  XNOR2_X1 U13030 ( .A(n14786), .B(n10649), .ZN(n13015) );
  NAND2_X1 U13031 ( .A1(n10521), .A2(n13015), .ZN(n10642) );
  OAI21_X1 U13032 ( .B1(n10521), .B2(n13015), .A(n10642), .ZN(n14793) );
  INV_X1 U13033 ( .A(n14793), .ZN(n10528) );
  NAND2_X1 U13034 ( .A1(n14835), .A2(n10522), .ZN(n10523) );
  XOR2_X1 U13035 ( .A(n10648), .B(n13015), .Z(n10526) );
  AOI21_X1 U13036 ( .B1(n10526), .B2(n14798), .A(n10525), .ZN(n14795) );
  INV_X1 U13037 ( .A(n14786), .ZN(n10531) );
  INV_X1 U13038 ( .A(n10645), .ZN(n10646) );
  OAI211_X1 U13039 ( .C1(n10531), .C2(n10527), .A(n10646), .B(n10803), .ZN(
        n14790) );
  OAI211_X1 U13040 ( .C1(n13529), .C2(n10528), .A(n14795), .B(n14790), .ZN(
        n10533) );
  OAI22_X1 U13041 ( .A1(n13502), .A2(n10531), .B1(n14861), .B2(n9264), .ZN(
        n10529) );
  AOI21_X1 U13042 ( .B1(n10533), .B2(n14861), .A(n10529), .ZN(n10530) );
  INV_X1 U13043 ( .A(n10530), .ZN(P2_U3506) );
  INV_X1 U13044 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15092) );
  OAI22_X1 U13045 ( .A1(n13556), .A2(n10531), .B1(n14855), .B2(n15092), .ZN(
        n10532) );
  AOI21_X1 U13046 ( .B1(n10533), .B2(n14855), .A(n10532), .ZN(n10534) );
  INV_X1 U13047 ( .A(n10534), .ZN(P2_U3451) );
  XNOR2_X1 U13048 ( .A(n11655), .B(n6517), .ZN(n10835) );
  XNOR2_X1 U13049 ( .A(n10835), .B(n14910), .ZN(n10538) );
  NAND2_X1 U13050 ( .A1(n10536), .A2(n10535), .ZN(n10537) );
  OAI21_X1 U13051 ( .B1(n10538), .B2(n10537), .A(n10858), .ZN(n10544) );
  AOI22_X1 U13052 ( .A1(n12190), .A2(n12206), .B1(n14333), .B2(n12205), .ZN(
        n10541) );
  AOI21_X1 U13053 ( .B1(n14341), .B2(n14981), .A(n10539), .ZN(n10540) );
  OAI211_X1 U13054 ( .C1(n14347), .C2(n10542), .A(n10541), .B(n10540), .ZN(
        n10543) );
  AOI21_X1 U13055 ( .B1(n10544), .B2(n14343), .A(n10543), .ZN(n10545) );
  INV_X1 U13056 ( .A(n10545), .ZN(P3_U3167) );
  NAND2_X1 U13057 ( .A1(n10547), .A2(n10546), .ZN(n10549) );
  NAND2_X1 U13058 ( .A1(n10612), .A2(n10606), .ZN(n10548) );
  INV_X1 U13059 ( .A(n10554), .ZN(n10550) );
  XNOR2_X1 U13060 ( .A(n10622), .B(n10550), .ZN(n10551) );
  NAND2_X1 U13061 ( .A1(n10551), .A2(n14264), .ZN(n10559) );
  AOI22_X1 U13062 ( .A1(n14154), .A2(n13853), .B1(n13851), .B2(n14152), .ZN(
        n10558) );
  OR2_X1 U13063 ( .A1(n10612), .A2(n13853), .ZN(n10552) );
  NAND2_X1 U13064 ( .A1(n10553), .A2(n10552), .ZN(n10555) );
  OR2_X1 U13065 ( .A1(n10555), .A2(n10554), .ZN(n10556) );
  NAND2_X1 U13066 ( .A1(n10556), .A2(n10617), .ZN(n14607) );
  NAND2_X1 U13067 ( .A1(n14607), .A2(n14057), .ZN(n10557) );
  NAND3_X1 U13068 ( .A1(n10559), .A2(n10558), .A3(n10557), .ZN(n14605) );
  MUX2_X1 U13069 ( .A(n14605), .B(P1_REG2_REG_7__SCAN_IN), .S(n14159), .Z(
        n10560) );
  INV_X1 U13070 ( .A(n10560), .ZN(n10567) );
  INV_X1 U13071 ( .A(n10689), .ZN(n14603) );
  NAND2_X1 U13072 ( .A1(n14603), .A2(n10561), .ZN(n10661) );
  OR2_X1 U13073 ( .A1(n10561), .A2(n14603), .ZN(n10562) );
  NAND2_X1 U13074 ( .A1(n10661), .A2(n10562), .ZN(n14604) );
  OAI22_X1 U13075 ( .A1(n14161), .A2(n14603), .B1(n14106), .B2(n10683), .ZN(
        n10563) );
  INV_X1 U13076 ( .A(n10563), .ZN(n10564) );
  OAI21_X1 U13077 ( .B1(n14604), .B2(n14112), .A(n10564), .ZN(n10565) );
  AOI21_X1 U13078 ( .B1(n14607), .B2(n14064), .A(n10565), .ZN(n10566) );
  NAND2_X1 U13079 ( .A1(n10567), .A2(n10566), .ZN(P1_U3286) );
  INV_X1 U13080 ( .A(n10568), .ZN(n10570) );
  OAI22_X1 U13081 ( .A1(n11836), .A2(P3_U3151), .B1(SI_22_), .B2(n12698), .ZN(
        n10569) );
  AOI21_X1 U13082 ( .B1(n10570), .B2(n12680), .A(n10569), .ZN(P3_U3273) );
  NAND2_X1 U13083 ( .A1(n10571), .A2(n10581), .ZN(n10572) );
  NAND2_X1 U13084 ( .A1(n10573), .A2(n10572), .ZN(n14602) );
  INV_X1 U13085 ( .A(n10574), .ZN(n10577) );
  NAND2_X1 U13086 ( .A1(n10575), .A2(n10579), .ZN(n10576) );
  NAND2_X1 U13087 ( .A1(n10577), .A2(n10576), .ZN(n14599) );
  AOI22_X1 U13088 ( .A1(n14110), .A2(n10579), .B1(n14157), .B2(n10578), .ZN(
        n10580) );
  OAI21_X1 U13089 ( .B1(n14112), .B2(n14599), .A(n10580), .ZN(n10590) );
  XNOR2_X1 U13090 ( .A(n10581), .B(n10582), .ZN(n10583) );
  NAND2_X1 U13091 ( .A1(n10583), .A2(n14264), .ZN(n10588) );
  NAND2_X1 U13092 ( .A1(n13853), .A2(n14152), .ZN(n10584) );
  OAI21_X1 U13093 ( .B1(n10585), .B2(n14136), .A(n10584), .ZN(n10586) );
  AOI21_X1 U13094 ( .B1(n14602), .B2(n14057), .A(n10586), .ZN(n10587) );
  NAND2_X1 U13095 ( .A1(n10588), .A2(n10587), .ZN(n14600) );
  MUX2_X1 U13096 ( .A(n14600), .B(P1_REG2_REG_5__SCAN_IN), .S(n14159), .Z(
        n10589) );
  AOI211_X1 U13097 ( .C1(n14064), .C2(n14602), .A(n10590), .B(n10589), .ZN(
        n10591) );
  INV_X1 U13098 ( .A(n10591), .ZN(P1_U3288) );
  INV_X1 U13099 ( .A(n10615), .ZN(n10592) );
  AOI22_X1 U13100 ( .A1(n14110), .A2(n10612), .B1(n10592), .B2(n14157), .ZN(
        n10593) );
  OAI21_X1 U13101 ( .B1(n14112), .B2(n10594), .A(n10593), .ZN(n10597) );
  MUX2_X1 U13102 ( .A(n10595), .B(P1_REG2_REG_6__SCAN_IN), .S(n14159), .Z(
        n10596) );
  AOI211_X1 U13103 ( .C1(n14064), .C2(n10598), .A(n10597), .B(n10596), .ZN(
        n10599) );
  INV_X1 U13104 ( .A(n10599), .ZN(P1_U3287) );
  OAI22_X1 U13105 ( .A1(n10603), .A2(n13739), .B1(n10606), .B2(n13741), .ZN(
        n10604) );
  XNOR2_X1 U13106 ( .A(n10604), .B(n13705), .ZN(n10674) );
  NOR2_X1 U13107 ( .A1(n10606), .A2(n13740), .ZN(n10607) );
  AOI21_X1 U13108 ( .B1(n10612), .B2(n13697), .A(n10607), .ZN(n10677) );
  XNOR2_X1 U13109 ( .A(n10674), .B(n10677), .ZN(n10608) );
  NAND2_X1 U13110 ( .A1(n10609), .A2(n10608), .ZN(n10675) );
  OAI211_X1 U13111 ( .C1(n10609), .C2(n10608), .A(n10675), .B(n14464), .ZN(
        n10614) );
  NAND2_X1 U13112 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n13926) );
  OAI21_X1 U13113 ( .B1(n13808), .B2(n10610), .A(n13926), .ZN(n10611) );
  AOI21_X1 U13114 ( .B1(n14481), .B2(n10612), .A(n10611), .ZN(n10613) );
  OAI211_X1 U13115 ( .C1(n14485), .C2(n10615), .A(n10614), .B(n10613), .ZN(
        P1_U3239) );
  OR2_X1 U13116 ( .A1(n10689), .A2(n13852), .ZN(n10616) );
  OR2_X1 U13117 ( .A1(n11030), .A2(n13851), .ZN(n10618) );
  OAI21_X1 U13118 ( .B1(n10619), .B2(n10627), .A(n10788), .ZN(n10620) );
  INV_X1 U13119 ( .A(n10620), .ZN(n14622) );
  AND2_X1 U13120 ( .A1(n10689), .A2(n10679), .ZN(n10621) );
  OR2_X1 U13121 ( .A1(n10689), .A2(n10679), .ZN(n10623) );
  INV_X1 U13122 ( .A(n10666), .ZN(n10626) );
  NOR2_X1 U13123 ( .A1(n11030), .A2(n10624), .ZN(n10625) );
  INV_X1 U13124 ( .A(n10627), .ZN(n10628) );
  OAI21_X1 U13125 ( .B1(n10629), .B2(n10628), .A(n10785), .ZN(n10630) );
  AOI222_X1 U13126 ( .A1(n14264), .A2(n10630), .B1(n13849), .B2(n14152), .C1(
        n13851), .C2(n14154), .ZN(n14621) );
  MUX2_X1 U13127 ( .A(n10631), .B(n14621), .S(n14076), .Z(n10635) );
  OR2_X1 U13128 ( .A1(n10661), .A2(n11030), .ZN(n10662) );
  AOI21_X1 U13129 ( .B1(n14616), .B2(n10662), .A(n10790), .ZN(n14619) );
  INV_X1 U13130 ( .A(n14616), .ZN(n10632) );
  OAI22_X1 U13131 ( .A1(n10632), .A2(n14161), .B1(n14106), .B2(n11165), .ZN(
        n10633) );
  AOI21_X1 U13132 ( .B1(n14619), .B2(n14167), .A(n10633), .ZN(n10634) );
  OAI211_X1 U13133 ( .C1(n14622), .C2(n14164), .A(n10635), .B(n10634), .ZN(
        P1_U3284) );
  INV_X1 U13134 ( .A(n11848), .ZN(n10639) );
  INV_X1 U13135 ( .A(n11286), .ZN(n14570) );
  OAI222_X1 U13136 ( .A1(n14302), .A2(n10636), .B1(n14305), .B2(n10639), .C1(
        n14570), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13137 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10640) );
  NAND2_X1 U13138 ( .A1(n10637), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10638) );
  XNOR2_X1 U13139 ( .A(n10638), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13128) );
  INV_X1 U13140 ( .A(n13128), .ZN(n11183) );
  OAI222_X1 U13141 ( .A1(n13580), .A2(n10640), .B1(n13574), .B2(n10639), .C1(
        P2_U3088), .C2(n11183), .ZN(P2_U3309) );
  XNOR2_X1 U13142 ( .A(n12857), .B(n13068), .ZN(n13016) );
  OR2_X1 U13143 ( .A1(n14786), .A2(n13069), .ZN(n10641) );
  INV_X1 U13144 ( .A(n10766), .ZN(n10643) );
  AOI21_X1 U13145 ( .B1(n13016), .B2(n10644), .A(n10643), .ZN(n10699) );
  AND2_X2 U13146 ( .A1(n10655), .A2(n10645), .ZN(n10802) );
  AOI211_X1 U13147 ( .C1(n12857), .C2(n10646), .A(n9459), .B(n10802), .ZN(
        n10692) );
  OR2_X1 U13148 ( .A1(n14786), .A2(n10649), .ZN(n10647) );
  OAI211_X1 U13149 ( .C1(n10650), .C2(n13016), .A(n14798), .B(n10772), .ZN(
        n10652) );
  NAND2_X1 U13150 ( .A1(n10652), .A2(n10651), .ZN(n10696) );
  AOI211_X1 U13151 ( .C1(n10699), .C2(n14833), .A(n10692), .B(n10696), .ZN(
        n10658) );
  INV_X1 U13152 ( .A(n13502), .ZN(n10977) );
  AOI22_X1 U13153 ( .A1(n10977), .A2(n12857), .B1(n13449), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n10653) );
  OAI21_X1 U13154 ( .B1(n10658), .B2(n13449), .A(n10653), .ZN(P2_U3507) );
  INV_X1 U13155 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10654) );
  OAI22_X1 U13156 ( .A1(n10655), .A2(n13556), .B1(n14855), .B2(n10654), .ZN(
        n10656) );
  INV_X1 U13157 ( .A(n10656), .ZN(n10657) );
  OAI21_X1 U13158 ( .B1(n10658), .B2(n13539), .A(n10657), .ZN(P2_U3454) );
  OAI21_X1 U13159 ( .B1(n10660), .B2(n10666), .A(n10659), .ZN(n14614) );
  INV_X1 U13160 ( .A(n10661), .ZN(n10663) );
  INV_X1 U13161 ( .A(n11030), .ZN(n14610) );
  OAI21_X1 U13162 ( .B1(n10663), .B2(n14610), .A(n10662), .ZN(n14611) );
  INV_X1 U13163 ( .A(n11028), .ZN(n10664) );
  AOI22_X1 U13164 ( .A1(n14110), .A2(n11030), .B1(n10664), .B2(n14157), .ZN(
        n10665) );
  OAI21_X1 U13165 ( .B1(n14611), .B2(n14112), .A(n10665), .ZN(n10672) );
  XNOR2_X1 U13166 ( .A(n10667), .B(n10666), .ZN(n10668) );
  NAND2_X1 U13167 ( .A1(n10668), .A2(n14264), .ZN(n10670) );
  AOI22_X1 U13168 ( .A1(n14154), .A2(n13852), .B1(n13850), .B2(n14152), .ZN(
        n10669) );
  NAND2_X1 U13169 ( .A1(n10670), .A2(n10669), .ZN(n14612) );
  MUX2_X1 U13170 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n14612), .S(n14076), .Z(
        n10671) );
  AOI211_X1 U13171 ( .C1(n14114), .C2(n14614), .A(n10672), .B(n10671), .ZN(
        n10673) );
  INV_X1 U13172 ( .A(n10673), .ZN(P1_U3285) );
  INV_X1 U13173 ( .A(n10674), .ZN(n10676) );
  OAI21_X1 U13174 ( .B1(n10677), .B2(n10676), .A(n10675), .ZN(n10682) );
  OAI22_X1 U13175 ( .A1(n14603), .A2(n13739), .B1(n10679), .B2(n13741), .ZN(
        n10678) );
  XNOR2_X1 U13176 ( .A(n10678), .B(n13705), .ZN(n11016) );
  NOR2_X1 U13177 ( .A1(n10679), .A2(n13740), .ZN(n10680) );
  AOI21_X1 U13178 ( .B1(n10689), .B2(n13697), .A(n10680), .ZN(n11017) );
  XNOR2_X1 U13179 ( .A(n11016), .B(n11017), .ZN(n10681) );
  NAND2_X1 U13180 ( .A1(n10682), .A2(n10681), .ZN(n11020) );
  OAI211_X1 U13181 ( .C1(n10682), .C2(n10681), .A(n11020), .B(n14464), .ZN(
        n10691) );
  NOR2_X1 U13182 ( .A1(n14485), .A2(n10683), .ZN(n10688) );
  NAND2_X1 U13183 ( .A1(n14459), .A2(n13853), .ZN(n10686) );
  NAND2_X1 U13184 ( .A1(n14457), .A2(n13851), .ZN(n10685) );
  NAND3_X1 U13185 ( .A1(n10686), .A2(n10685), .A3(n10684), .ZN(n10687) );
  AOI211_X1 U13186 ( .C1(n10689), .C2(n14481), .A(n10688), .B(n10687), .ZN(
        n10690) );
  NAND2_X1 U13187 ( .A1(n10691), .A2(n10690), .ZN(P1_U3213) );
  INV_X1 U13188 ( .A(n10692), .ZN(n10695) );
  AOI22_X1 U13189 ( .A1(n12857), .A2(n14785), .B1(n14783), .B2(n10693), .ZN(
        n10694) );
  OAI21_X1 U13190 ( .B1(n10695), .B2(n14789), .A(n10694), .ZN(n10698) );
  MUX2_X1 U13191 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10696), .S(n14809), .Z(
        n10697) );
  AOI211_X1 U13192 ( .C1(n14792), .C2(n10699), .A(n10698), .B(n10697), .ZN(
        n10700) );
  INV_X1 U13193 ( .A(n10700), .ZN(P2_U3257) );
  NOR2_X1 U13194 ( .A1(n10708), .A2(n10701), .ZN(n10703) );
  INV_X1 U13195 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10715) );
  MUX2_X1 U13196 ( .A(n10715), .B(P3_REG1_REG_10__SCAN_IN), .S(n11080), .Z(
        n10705) );
  INV_X1 U13197 ( .A(n11075), .ZN(n10704) );
  AOI21_X1 U13198 ( .B1(n10706), .B2(n10705), .A(n10704), .ZN(n10730) );
  NOR2_X1 U13199 ( .A1(n10708), .A2(n10707), .ZN(n10710) );
  INV_X1 U13200 ( .A(n10712), .ZN(n10714) );
  MUX2_X1 U13201 ( .A(n10716), .B(P3_REG2_REG_10__SCAN_IN), .S(n11080), .Z(
        n10711) );
  INV_X1 U13202 ( .A(n10711), .ZN(n10713) );
  OAI21_X1 U13203 ( .B1(n10714), .B2(n10713), .A(n11082), .ZN(n10728) );
  MUX2_X1 U13204 ( .A(n10716), .B(n10715), .S(n12691), .Z(n10718) );
  INV_X1 U13205 ( .A(n11080), .ZN(n10717) );
  NAND2_X1 U13206 ( .A1(n10718), .A2(n10717), .ZN(n11089) );
  INV_X1 U13207 ( .A(n10718), .ZN(n10719) );
  NAND2_X1 U13208 ( .A1(n10719), .A2(n11080), .ZN(n10720) );
  NAND2_X1 U13209 ( .A1(n11089), .A2(n10720), .ZN(n10721) );
  AOI21_X1 U13210 ( .B1(n10723), .B2(n10722), .A(n10721), .ZN(n11091) );
  AND3_X1 U13211 ( .A1(n10723), .A2(n10722), .A3(n10721), .ZN(n10724) );
  OAI21_X1 U13212 ( .B1(n11091), .B2(n10724), .A(n14893), .ZN(n10726) );
  AND2_X1 U13213 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n12075) );
  AOI21_X1 U13214 ( .B1(n14862), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n12075), 
        .ZN(n10725) );
  OAI211_X1 U13215 ( .C1(n14885), .C2(n11080), .A(n10726), .B(n10725), .ZN(
        n10727) );
  AOI21_X1 U13216 ( .B1(n12307), .B2(n10728), .A(n10727), .ZN(n10729) );
  OAI21_X1 U13217 ( .B1(n10730), .B2(n14897), .A(n10729), .ZN(P3_U3192) );
  INV_X1 U13218 ( .A(n10731), .ZN(n10732) );
  OR2_X1 U13219 ( .A1(n10734), .A2(n11375), .ZN(n10737) );
  AOI22_X1 U13220 ( .A1(n11862), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10735), 
        .B2(n11861), .ZN(n10736) );
  NAND2_X2 U13221 ( .A1(n10737), .A2(n10736), .ZN(n14639) );
  XNOR2_X1 U13222 ( .A(n14639), .B(n11976), .ZN(n10739) );
  NAND2_X1 U13223 ( .A1(n13066), .A2(n6520), .ZN(n10738) );
  XNOR2_X1 U13224 ( .A(n10739), .B(n10738), .ZN(n14637) );
  INV_X1 U13225 ( .A(n10738), .ZN(n10740) );
  NAND2_X1 U13226 ( .A1(n12958), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10746) );
  NAND2_X1 U13227 ( .A1(n12941), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10745) );
  OR2_X1 U13228 ( .A1(n10741), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10742) );
  AND2_X1 U13229 ( .A1(n10752), .A2(n10742), .ZN(n11005) );
  NAND2_X1 U13230 ( .A1(n12004), .A2(n11005), .ZN(n10744) );
  NAND2_X1 U13231 ( .A1(n12959), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10743) );
  NAND4_X1 U13232 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        n13065) );
  NAND2_X1 U13233 ( .A1(n13065), .A2(n6520), .ZN(n10882) );
  NAND2_X1 U13234 ( .A1(n10747), .A2(n12963), .ZN(n10750) );
  AOI22_X1 U13235 ( .A1(n10748), .A2(n11861), .B1(n11862), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n10749) );
  XNOR2_X1 U13236 ( .A(n14844), .B(n11976), .ZN(n10881) );
  XOR2_X1 U13237 ( .A(n10882), .B(n10881), .Z(n10883) );
  XNOR2_X1 U13238 ( .A(n10884), .B(n10883), .ZN(n10764) );
  INV_X1 U13239 ( .A(n11005), .ZN(n10761) );
  NAND2_X1 U13240 ( .A1(n12941), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10757) );
  NAND2_X1 U13241 ( .A1(n12958), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10756) );
  INV_X1 U13242 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10751) );
  NAND2_X1 U13243 ( .A1(n10752), .A2(n10751), .ZN(n10753) );
  AND2_X1 U13244 ( .A1(n10893), .A2(n10753), .ZN(n11144) );
  NAND2_X1 U13245 ( .A1(n12004), .A2(n11144), .ZN(n10755) );
  NAND2_X1 U13246 ( .A1(n12959), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10754) );
  NAND4_X1 U13247 ( .A1(n10757), .A2(n10756), .A3(n10755), .A4(n10754), .ZN(
        n13064) );
  NAND2_X1 U13248 ( .A1(n13064), .A2(n13407), .ZN(n10759) );
  NAND2_X1 U13249 ( .A1(n13066), .A2(n13405), .ZN(n10758) );
  NAND2_X1 U13250 ( .A1(n10759), .A2(n10758), .ZN(n11000) );
  AOI22_X1 U13251 ( .A1(n12783), .A2(n11000), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10760) );
  OAI21_X1 U13252 ( .B1(n10761), .B2(n14660), .A(n10760), .ZN(n10762) );
  AOI21_X1 U13253 ( .B1(n14844), .B2(n14657), .A(n10762), .ZN(n10763) );
  OAI21_X1 U13254 ( .B1(n10764), .B2(n14652), .A(n10763), .ZN(P2_U3208) );
  NAND2_X1 U13255 ( .A1(n12857), .A2(n13068), .ZN(n10765) );
  XNOR2_X1 U13256 ( .A(n13424), .B(n13067), .ZN(n13017) );
  INV_X1 U13257 ( .A(n13017), .ZN(n10767) );
  NAND2_X1 U13258 ( .A1(n13424), .A2(n13067), .ZN(n10768) );
  NAND2_X1 U13259 ( .A1(n10769), .A2(n10768), .ZN(n11009) );
  XNOR2_X1 U13260 ( .A(n14639), .B(n13066), .ZN(n13019) );
  XNOR2_X1 U13261 ( .A(n11009), .B(n13019), .ZN(n10976) );
  INV_X1 U13262 ( .A(n10976), .ZN(n10783) );
  OR2_X1 U13263 ( .A1(n12857), .A2(n10770), .ZN(n10771) );
  INV_X1 U13264 ( .A(n13067), .ZN(n10773) );
  OR2_X1 U13265 ( .A1(n13424), .A2(n10773), .ZN(n10774) );
  OAI211_X1 U13266 ( .C1(n10775), .C2(n13019), .A(n10996), .B(n14798), .ZN(
        n10776) );
  AOI22_X1 U13267 ( .A1(n13405), .A2(n13067), .B1(n13065), .B2(n13407), .ZN(
        n14642) );
  NAND2_X1 U13268 ( .A1(n10776), .A2(n14642), .ZN(n10974) );
  INV_X1 U13269 ( .A(n11002), .ZN(n10777) );
  AOI211_X1 U13270 ( .C1(n14639), .C2(n10805), .A(n9459), .B(n10777), .ZN(
        n10975) );
  NAND2_X1 U13271 ( .A1(n10975), .A2(n13425), .ZN(n10780) );
  AOI22_X1 U13272 ( .A1(n14811), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10778), 
        .B2(n14783), .ZN(n10779) );
  OAI211_X1 U13273 ( .C1(n7239), .C2(n13390), .A(n10780), .B(n10779), .ZN(
        n10781) );
  AOI21_X1 U13274 ( .B1(n10974), .B2(n14809), .A(n10781), .ZN(n10782) );
  OAI21_X1 U13275 ( .B1(n10783), .B2(n13396), .A(n10782), .ZN(P2_U3255) );
  NAND2_X1 U13276 ( .A1(n14616), .A2(n11025), .ZN(n10784) );
  XNOR2_X1 U13277 ( .A(n10946), .B(n10945), .ZN(n10990) );
  OR2_X1 U13278 ( .A1(n14616), .A2(n13850), .ZN(n10787) );
  NAND2_X1 U13279 ( .A1(n10789), .A2(n10945), .ZN(n10951) );
  OAI21_X1 U13280 ( .B1(n10789), .B2(n10945), .A(n10951), .ZN(n10987) );
  INV_X1 U13281 ( .A(n10790), .ZN(n10791) );
  AOI211_X1 U13282 ( .C1(n11345), .C2(n10791), .A(n9590), .B(n7019), .ZN(
        n10986) );
  NAND2_X1 U13283 ( .A1(n13848), .A2(n14152), .ZN(n10984) );
  INV_X1 U13284 ( .A(n10984), .ZN(n10793) );
  NOR2_X1 U13285 ( .A1(n13989), .A2(n10792), .ZN(n14063) );
  OAI21_X1 U13286 ( .B1(n10986), .B2(n10793), .A(n14063), .ZN(n10796) );
  NAND2_X1 U13287 ( .A1(n13850), .A2(n14154), .ZN(n10985) );
  OAI22_X1 U13288 ( .A1(n14159), .A2(n10985), .B1(n11348), .B2(n14106), .ZN(
        n10794) );
  AOI21_X1 U13289 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n14159), .A(n10794), 
        .ZN(n10795) );
  OAI211_X1 U13290 ( .C1(n6948), .C2(n14161), .A(n10796), .B(n10795), .ZN(
        n10797) );
  AOI21_X1 U13291 ( .B1(n14114), .B2(n10987), .A(n10797), .ZN(n10798) );
  OAI21_X1 U13292 ( .B1(n10990), .B2(n14116), .A(n10798), .ZN(P1_U3283) );
  INV_X1 U13293 ( .A(n11860), .ZN(n10800) );
  OAI222_X1 U13294 ( .A1(n11295), .A2(P1_U3086), .B1(n14305), .B2(n10800), 
        .C1(n10799), .C2(n14302), .ZN(P1_U3336) );
  OAI222_X1 U13295 ( .A1(n13580), .A2(n15116), .B1(n13578), .B2(n10800), .C1(
        n13412), .C2(P2_U3088), .ZN(P2_U3308) );
  XNOR2_X1 U13296 ( .A(n10801), .B(n13017), .ZN(n13418) );
  OR2_X1 U13297 ( .A1(n10802), .A2(n10812), .ZN(n10804) );
  AND3_X1 U13298 ( .A1(n10805), .A2(n10804), .A3(n10803), .ZN(n13426) );
  OAI211_X1 U13299 ( .C1(n10807), .C2(n13017), .A(n10806), .B(n14798), .ZN(
        n10809) );
  NAND2_X1 U13300 ( .A1(n10809), .A2(n10808), .ZN(n13419) );
  AOI211_X1 U13301 ( .C1(n14833), .C2(n13418), .A(n13426), .B(n13419), .ZN(
        n10815) );
  AOI22_X1 U13302 ( .A1(n13424), .A2(n10977), .B1(n13449), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10810) );
  OAI21_X1 U13303 ( .B1(n10815), .B2(n13449), .A(n10810), .ZN(P2_U3508) );
  INV_X1 U13304 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10811) );
  OAI22_X1 U13305 ( .A1(n10812), .A2(n13556), .B1(n14855), .B2(n10811), .ZN(
        n10813) );
  INV_X1 U13306 ( .A(n10813), .ZN(n10814) );
  OAI21_X1 U13307 ( .B1(n10815), .B2(n13539), .A(n10814), .ZN(P2_U3457) );
  MUX2_X1 U13308 ( .A(n11479), .B(P1_REG2_REG_17__SCAN_IN), .S(n11273), .Z(
        n11274) );
  INV_X1 U13309 ( .A(n10816), .ZN(n10817) );
  OAI21_X1 U13310 ( .B1(n10818), .B2(n11303), .A(n10817), .ZN(n10819) );
  NOR2_X1 U13311 ( .A1(n10827), .A2(n10819), .ZN(n10820) );
  XNOR2_X1 U13312 ( .A(n10819), .B(n10827), .ZN(n14551) );
  NOR2_X1 U13313 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14551), .ZN(n14550) );
  NOR2_X1 U13314 ( .A1(n10820), .A2(n14550), .ZN(n13969) );
  NAND2_X1 U13315 ( .A1(n10822), .A2(n13964), .ZN(n10821) );
  OAI211_X1 U13316 ( .C1(n10822), .C2(n13964), .A(n13969), .B(n10821), .ZN(
        n13967) );
  OAI21_X1 U13317 ( .B1(n13964), .B2(n10822), .A(n13967), .ZN(n11276) );
  XOR2_X1 U13318 ( .A(n11274), .B(n11276), .Z(n10834) );
  NOR2_X1 U13319 ( .A1(n14571), .A2(n11282), .ZN(n10832) );
  NAND2_X1 U13320 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3086), .ZN(n14466)
         );
  XNOR2_X1 U13321 ( .A(n11273), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11284) );
  OR2_X1 U13322 ( .A1(n10823), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10824) );
  AND2_X1 U13323 ( .A1(n10825), .A2(n10824), .ZN(n10828) );
  XNOR2_X1 U13324 ( .A(n10828), .B(n10827), .ZN(n14549) );
  NOR2_X1 U13325 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14549), .ZN(n14548) );
  INV_X1 U13326 ( .A(n14548), .ZN(n10826) );
  OAI21_X1 U13327 ( .B1(n10828), .B2(n10827), .A(n10826), .ZN(n13959) );
  XNOR2_X1 U13328 ( .A(n13966), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n13960) );
  NOR2_X1 U13329 ( .A1(n13959), .A2(n13960), .ZN(n13958) );
  AOI21_X1 U13330 ( .B1(n13966), .B2(P1_REG1_REG_16__SCAN_IN), .A(n13958), 
        .ZN(n11285) );
  XOR2_X1 U13331 ( .A(n11284), .B(n11285), .Z(n10829) );
  NAND2_X1 U13332 ( .A1(n10829), .A2(n14566), .ZN(n10830) );
  NAND2_X1 U13333 ( .A1(n14466), .A2(n10830), .ZN(n10831) );
  AOI211_X1 U13334 ( .C1(n14544), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n10832), 
        .B(n10831), .ZN(n10833) );
  OAI21_X1 U13335 ( .B1(n10834), .B2(n14552), .A(n10833), .ZN(P1_U3260) );
  XNOR2_X1 U13336 ( .A(n10850), .B(n12095), .ZN(n11117) );
  XNOR2_X1 U13337 ( .A(n11117), .B(n12202), .ZN(n10848) );
  XNOR2_X1 U13338 ( .A(n10871), .B(n12095), .ZN(n11033) );
  XNOR2_X1 U13339 ( .A(n10916), .B(n12095), .ZN(n10859) );
  XNOR2_X1 U13340 ( .A(n11038), .B(n12095), .ZN(n10840) );
  XNOR2_X1 U13341 ( .A(n10840), .B(n12203), .ZN(n10838) );
  NAND2_X1 U13342 ( .A1(n10909), .A2(n10835), .ZN(n10857) );
  OAI211_X1 U13343 ( .C1(n10859), .C2(n12205), .A(n10838), .B(n10857), .ZN(
        n10836) );
  NOR2_X1 U13344 ( .A1(n11033), .A2(n10836), .ZN(n10837) );
  INV_X1 U13345 ( .A(n12204), .ZN(n10908) );
  INV_X1 U13346 ( .A(n10838), .ZN(n11035) );
  OAI21_X1 U13347 ( .B1(n10908), .B2(n11035), .A(n11033), .ZN(n10843) );
  NAND2_X1 U13348 ( .A1(n10859), .A2(n12205), .ZN(n10860) );
  INV_X1 U13349 ( .A(n11033), .ZN(n10839) );
  OAI21_X1 U13350 ( .B1(n11035), .B2(n10860), .A(n10839), .ZN(n10842) );
  INV_X1 U13351 ( .A(n10840), .ZN(n10841) );
  AOI22_X1 U13352 ( .A1(n10843), .A2(n10842), .B1(n10841), .B2(n12203), .ZN(
        n10844) );
  INV_X1 U13353 ( .A(n12071), .ZN(n10846) );
  AOI21_X1 U13354 ( .B1(n10848), .B2(n10847), .A(n10846), .ZN(n10856) );
  INV_X1 U13355 ( .A(n12203), .ZN(n10849) );
  OAI22_X1 U13356 ( .A1(n12198), .A2(n10850), .B1(n10849), .B2(n14336), .ZN(
        n10851) );
  AOI211_X1 U13357 ( .C1(n14333), .C2(n14371), .A(n10852), .B(n10851), .ZN(
        n10855) );
  INV_X1 U13358 ( .A(n11054), .ZN(n10853) );
  NAND2_X1 U13359 ( .A1(n12195), .A2(n10853), .ZN(n10854) );
  OAI211_X1 U13360 ( .C1(n10856), .C2(n12174), .A(n10855), .B(n10854), .ZN(
        P3_U3171) );
  AND2_X1 U13361 ( .A1(n10858), .A2(n10857), .ZN(n12178) );
  XOR2_X1 U13362 ( .A(n10859), .B(n12205), .Z(n12177) );
  NAND2_X1 U13363 ( .A1(n12178), .A2(n12177), .ZN(n12176) );
  NAND2_X1 U13364 ( .A1(n12176), .A2(n10860), .ZN(n11034) );
  XNOR2_X1 U13365 ( .A(n11034), .B(n11033), .ZN(n10866) );
  AOI22_X1 U13366 ( .A1(n14333), .A2(n12203), .B1(n12190), .B2(n12205), .ZN(
        n10864) );
  AOI21_X1 U13367 ( .B1(n14341), .B2(n10862), .A(n10861), .ZN(n10863) );
  OAI211_X1 U13368 ( .C1(n14347), .C2(n10868), .A(n10864), .B(n10863), .ZN(
        n10865) );
  AOI21_X1 U13369 ( .B1(n10866), .B2(n14343), .A(n10865), .ZN(n10867) );
  INV_X1 U13370 ( .A(n10867), .ZN(P3_U3153) );
  INV_X1 U13371 ( .A(n10868), .ZN(n10877) );
  NAND2_X1 U13372 ( .A1(n10906), .A2(n11660), .ZN(n10869) );
  XNOR2_X1 U13373 ( .A(n10869), .B(n11794), .ZN(n14993) );
  NAND2_X1 U13374 ( .A1(n14993), .A2(n14978), .ZN(n10876) );
  OAI211_X1 U13375 ( .C1(n10872), .C2(n10871), .A(n10870), .B(n14934), .ZN(
        n10874) );
  AOI22_X1 U13376 ( .A1(n14944), .A2(n12203), .B1(n12205), .B2(n14946), .ZN(
        n10873) );
  AND2_X1 U13377 ( .A1(n10874), .A2(n10873), .ZN(n10875) );
  NAND2_X1 U13378 ( .A1(n10876), .A2(n10875), .ZN(n14997) );
  AOI21_X1 U13379 ( .B1(n14952), .B2(n10877), .A(n14997), .ZN(n10880) );
  INV_X1 U13380 ( .A(n10971), .ZN(n14953) );
  OAI22_X1 U13381 ( .A1(n14354), .A2(n14994), .B1(n10035), .B2(n14955), .ZN(
        n10878) );
  AOI21_X1 U13382 ( .B1(n14993), .B2(n14953), .A(n10878), .ZN(n10879) );
  OAI21_X1 U13383 ( .B1(n10880), .B2(n14957), .A(n10879), .ZN(P3_U3226) );
  NAND2_X1 U13384 ( .A1(n10885), .A2(n12963), .ZN(n10889) );
  NOR2_X1 U13385 ( .A1(n6521), .A2(n15119), .ZN(n10886) );
  AOI21_X1 U13386 ( .B1(n10887), .B2(n11861), .A(n10886), .ZN(n10888) );
  XNOR2_X1 U13387 ( .A(n12880), .B(n11948), .ZN(n10891) );
  NAND2_X1 U13388 ( .A1(n13064), .A2(n6520), .ZN(n10890) );
  NOR2_X1 U13389 ( .A1(n10891), .A2(n10890), .ZN(n11520) );
  NOR2_X1 U13390 ( .A1(n11520), .A2(n6663), .ZN(n10892) );
  XNOR2_X1 U13391 ( .A(n11521), .B(n10892), .ZN(n10905) );
  INV_X1 U13392 ( .A(n11144), .ZN(n10902) );
  NAND2_X1 U13393 ( .A1(n12941), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U13394 ( .A1(n10893), .A2(n14648), .ZN(n10894) );
  NAND2_X1 U13395 ( .A1(n11388), .A2(n10894), .ZN(n14661) );
  INV_X1 U13396 ( .A(n14661), .ZN(n11223) );
  NAND2_X1 U13397 ( .A1(n12004), .A2(n11223), .ZN(n10897) );
  NAND2_X1 U13398 ( .A1(n12959), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10896) );
  NAND2_X1 U13399 ( .A1(n12958), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10895) );
  NAND4_X1 U13400 ( .A1(n10898), .A2(n10897), .A3(n10896), .A4(n10895), .ZN(
        n13063) );
  NAND2_X1 U13401 ( .A1(n13063), .A2(n13407), .ZN(n10900) );
  NAND2_X1 U13402 ( .A1(n13065), .A2(n13405), .ZN(n10899) );
  NAND2_X1 U13403 ( .A1(n10900), .A2(n10899), .ZN(n11141) );
  AOI22_X1 U13404 ( .A1(n12783), .A2(n11141), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10901) );
  OAI21_X1 U13405 ( .B1(n10902), .B2(n14660), .A(n10901), .ZN(n10903) );
  AOI21_X1 U13406 ( .B1(n12880), .B2(n14657), .A(n10903), .ZN(n10904) );
  OAI21_X1 U13407 ( .B1(n10905), .B2(n14652), .A(n10904), .ZN(P2_U3196) );
  OAI21_X1 U13408 ( .B1(n10907), .B2(n11791), .A(n10906), .ZN(n14990) );
  INV_X1 U13409 ( .A(n14990), .ZN(n10920) );
  OAI22_X1 U13410 ( .A1(n10909), .A2(n14932), .B1(n10908), .B2(n14930), .ZN(
        n10914) );
  INV_X1 U13411 ( .A(n10910), .ZN(n10911) );
  AOI211_X1 U13412 ( .C1(n11791), .C2(n10912), .A(n14949), .B(n10911), .ZN(
        n10913) );
  AOI211_X1 U13413 ( .C1(n14978), .C2(n14990), .A(n10914), .B(n10913), .ZN(
        n14987) );
  MUX2_X1 U13414 ( .A(n10915), .B(n14987), .S(n14955), .Z(n10919) );
  NOR2_X1 U13415 ( .A1(n10916), .A2(n15013), .ZN(n14989) );
  INV_X1 U13416 ( .A(n12181), .ZN(n10917) );
  AOI22_X1 U13417 ( .A1(n14379), .A2(n14989), .B1(n14952), .B2(n10917), .ZN(
        n10918) );
  OAI211_X1 U13418 ( .C1(n10920), .C2(n10971), .A(n10919), .B(n10918), .ZN(
        P3_U3227) );
  NAND2_X1 U13419 ( .A1(n10921), .A2(n12680), .ZN(n10922) );
  OAI211_X1 U13420 ( .C1(n10923), .C2(n12698), .A(n10922), .B(n11839), .ZN(
        P3_U3272) );
  NAND2_X1 U13421 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11538)
         );
  OAI21_X1 U13422 ( .B1(n14740), .B2(n11179), .A(n11538), .ZN(n10943) );
  INV_X1 U13423 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11178) );
  AOI22_X1 U13424 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n11517), .B1(n11179), 
        .B2(n11178), .ZN(n10930) );
  NAND2_X1 U13425 ( .A1(n11377), .A2(n10924), .ZN(n10926) );
  NAND2_X1 U13426 ( .A1(n10926), .A2(n10925), .ZN(n10927) );
  NAND2_X1 U13427 ( .A1(n10927), .A2(n14759), .ZN(n10928) );
  XOR2_X1 U13428 ( .A(n14759), .B(n10927), .Z(n14761) );
  NAND2_X1 U13429 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14761), .ZN(n14760) );
  NAND2_X1 U13430 ( .A1(n10928), .A2(n14760), .ZN(n10929) );
  NAND2_X1 U13431 ( .A1(n10930), .A2(n10929), .ZN(n11177) );
  OAI211_X1 U13432 ( .C1(n10930), .C2(n10929), .A(n14776), .B(n11177), .ZN(
        n10941) );
  INV_X1 U13433 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10932) );
  OAI22_X1 U13434 ( .A1(n10934), .A2(n10933), .B1(n10932), .B2(n10931), .ZN(
        n10935) );
  XNOR2_X1 U13435 ( .A(n10935), .B(n14759), .ZN(n14762) );
  INV_X1 U13436 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15200) );
  INV_X1 U13437 ( .A(n10935), .ZN(n10937) );
  OAI22_X1 U13438 ( .A1(n14762), .A2(n15200), .B1(n10937), .B2(n10936), .ZN(
        n10939) );
  XNOR2_X1 U13439 ( .A(n11179), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n10938) );
  NAND2_X1 U13440 ( .A1(n10938), .A2(n10939), .ZN(n11169) );
  OAI211_X1 U13441 ( .C1(n10939), .C2(n10938), .A(n14774), .B(n11169), .ZN(
        n10940) );
  NAND2_X1 U13442 ( .A1(n10941), .A2(n10940), .ZN(n10942) );
  AOI211_X1 U13443 ( .C1(n14768), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n10943), 
        .B(n10942), .ZN(n10944) );
  INV_X1 U13444 ( .A(n10944), .ZN(P2_U3230) );
  INV_X1 U13445 ( .A(n13849), .ZN(n14469) );
  XNOR2_X1 U13446 ( .A(n11104), .B(n10952), .ZN(n10947) );
  NAND2_X1 U13447 ( .A1(n10947), .A2(n14264), .ZN(n10949) );
  AOI22_X1 U13448 ( .A1(n14154), .A2(n13849), .B1(n13847), .B2(n14152), .ZN(
        n10948) );
  OR2_X1 U13449 ( .A1(n11345), .A2(n13849), .ZN(n10950) );
  NAND2_X1 U13450 ( .A1(n10951), .A2(n10950), .ZN(n10953) );
  OR2_X1 U13451 ( .A1(n10953), .A2(n10952), .ZN(n10954) );
  NAND2_X1 U13452 ( .A1(n6835), .A2(n10954), .ZN(n14507) );
  NAND2_X1 U13453 ( .A1(n14504), .A2(n10955), .ZN(n10956) );
  NAND2_X1 U13454 ( .A1(n11111), .A2(n10956), .ZN(n14505) );
  OAI22_X1 U13455 ( .A1(n14076), .A2(n10957), .B1(n14484), .B2(n14106), .ZN(
        n10958) );
  AOI21_X1 U13456 ( .B1(n14504), .B2(n14110), .A(n10958), .ZN(n10959) );
  OAI21_X1 U13457 ( .B1(n14505), .B2(n14112), .A(n10959), .ZN(n10960) );
  AOI21_X1 U13458 ( .B1(n14507), .B2(n14114), .A(n10960), .ZN(n10961) );
  OAI21_X1 U13459 ( .B1(n14509), .B2(n14159), .A(n10961), .ZN(P1_U3282) );
  XNOR2_X1 U13460 ( .A(n10962), .B(n11789), .ZN(n10964) );
  INV_X1 U13461 ( .A(n10964), .ZN(n15000) );
  XNOR2_X1 U13462 ( .A(n10963), .B(n7478), .ZN(n10967) );
  NAND2_X1 U13463 ( .A1(n10964), .A2(n14978), .ZN(n10966) );
  AOI22_X1 U13464 ( .A1(n14946), .A2(n12204), .B1(n12202), .B2(n14944), .ZN(
        n10965) );
  OAI211_X1 U13465 ( .C1(n10967), .C2(n14949), .A(n10966), .B(n10965), .ZN(
        n15002) );
  NAND2_X1 U13466 ( .A1(n15002), .A2(n14955), .ZN(n10970) );
  NAND2_X1 U13467 ( .A1(n11038), .A2(n14980), .ZN(n14999) );
  OAI22_X1 U13468 ( .A1(n11053), .A2(n14999), .B1(n6573), .B2(n14926), .ZN(
        n10968) );
  AOI21_X1 U13469 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14957), .A(n10968), .ZN(
        n10969) );
  OAI211_X1 U13470 ( .C1(n15000), .C2(n10971), .A(n10970), .B(n10969), .ZN(
        P3_U3225) );
  INV_X1 U13471 ( .A(n11868), .ZN(n11014) );
  OAI222_X1 U13472 ( .A1(P1_U3086), .A2(n10973), .B1(n14305), .B2(n11014), 
        .C1(n10972), .C2(n14302), .ZN(P1_U3335) );
  AOI211_X1 U13473 ( .C1(n14833), .C2(n10976), .A(n10975), .B(n10974), .ZN(
        n10983) );
  AOI22_X1 U13474 ( .A1(n14639), .A2(n10977), .B1(n13449), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n10978) );
  OAI21_X1 U13475 ( .B1(n10983), .B2(n13449), .A(n10978), .ZN(P2_U3509) );
  INV_X1 U13476 ( .A(n13556), .ZN(n10981) );
  INV_X1 U13477 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10979) );
  NOR2_X1 U13478 ( .A1(n14855), .A2(n10979), .ZN(n10980) );
  AOI21_X1 U13479 ( .B1(n14639), .B2(n10981), .A(n10980), .ZN(n10982) );
  OAI21_X1 U13480 ( .B1(n10983), .B2(n13539), .A(n10982), .ZN(P2_U3460) );
  NAND2_X1 U13481 ( .A1(n10985), .A2(n10984), .ZN(n11351) );
  AOI211_X1 U13482 ( .C1(n14617), .C2(n11345), .A(n11351), .B(n10986), .ZN(
        n10989) );
  NAND2_X1 U13483 ( .A1(n10987), .A2(n14615), .ZN(n10988) );
  OAI211_X1 U13484 ( .C1(n10990), .C2(n14275), .A(n10989), .B(n10988), .ZN(
        n10992) );
  NAND2_X1 U13485 ( .A1(n10992), .A2(n14636), .ZN(n10991) );
  OAI21_X1 U13486 ( .B1(n14636), .B2(n9432), .A(n10991), .ZN(P1_U3538) );
  NAND2_X1 U13487 ( .A1(n10992), .A2(n14627), .ZN(n10993) );
  OAI21_X1 U13488 ( .B1(n14627), .B2(n7909), .A(n10993), .ZN(P1_U3489) );
  INV_X1 U13489 ( .A(n13066), .ZN(n10994) );
  OR2_X1 U13490 ( .A1(n14639), .A2(n10994), .ZN(n10995) );
  XNOR2_X1 U13491 ( .A(n14844), .B(n13065), .ZN(n13022) );
  INV_X1 U13492 ( .A(n13022), .ZN(n10997) );
  NAND2_X1 U13493 ( .A1(n10998), .A2(n10997), .ZN(n10999) );
  NAND2_X1 U13494 ( .A1(n11135), .A2(n10999), .ZN(n11001) );
  AOI21_X1 U13495 ( .B1(n11001), .B2(n14798), .A(n11000), .ZN(n14853) );
  NAND2_X1 U13496 ( .A1(n14844), .A2(n11002), .ZN(n11003) );
  NAND2_X1 U13497 ( .A1(n11003), .A2(n10803), .ZN(n11004) );
  OR2_X1 U13498 ( .A1(n11143), .A2(n11004), .ZN(n14846) );
  INV_X1 U13499 ( .A(n14846), .ZN(n11008) );
  AOI22_X1 U13500 ( .A1(n14811), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11005), 
        .B2(n14783), .ZN(n11006) );
  OAI21_X1 U13501 ( .B1(n7241), .B2(n13390), .A(n11006), .ZN(n11007) );
  AOI21_X1 U13502 ( .B1(n11008), .B2(n13425), .A(n11007), .ZN(n11013) );
  NAND2_X1 U13503 ( .A1(n11009), .A2(n7141), .ZN(n11011) );
  NAND2_X1 U13504 ( .A1(n14639), .A2(n13066), .ZN(n11010) );
  XNOR2_X1 U13505 ( .A(n11150), .B(n13022), .ZN(n14849) );
  NAND2_X1 U13506 ( .A1(n14849), .A2(n14792), .ZN(n11012) );
  OAI211_X1 U13507 ( .C1(n14853), .C2(n14811), .A(n11013), .B(n11012), .ZN(
        P2_U3254) );
  OAI222_X1 U13508 ( .A1(n13580), .A2(n11869), .B1(P2_U3088), .B2(n13039), 
        .C1(n13578), .C2(n11014), .ZN(P2_U3307) );
  AOI22_X1 U13509 ( .A1(n11030), .A2(n13702), .B1(n13697), .B2(n13851), .ZN(
        n11015) );
  XNOR2_X1 U13510 ( .A(n11015), .B(n13705), .ZN(n11154) );
  AOI22_X1 U13511 ( .A1(n11030), .A2(n13697), .B1(n10343), .B2(n13851), .ZN(
        n11153) );
  XNOR2_X1 U13512 ( .A(n11154), .B(n11153), .ZN(n11023) );
  AOI21_X1 U13513 ( .B1(n11023), .B2(n11022), .A(n11021), .ZN(n11032) );
  OAI21_X1 U13514 ( .B1(n14471), .B2(n11025), .A(n11024), .ZN(n11026) );
  AOI21_X1 U13515 ( .B1(n14459), .B2(n13852), .A(n11026), .ZN(n11027) );
  OAI21_X1 U13516 ( .B1(n11028), .B2(n14485), .A(n11027), .ZN(n11029) );
  AOI21_X1 U13517 ( .B1(n11030), .B2(n14481), .A(n11029), .ZN(n11031) );
  OAI21_X1 U13518 ( .B1(n11032), .B2(n14476), .A(n11031), .ZN(P1_U3221) );
  MUX2_X1 U13519 ( .A(n11034), .B(n12204), .S(n11033), .Z(n11036) );
  XNOR2_X1 U13520 ( .A(n11036), .B(n11035), .ZN(n11042) );
  AOI22_X1 U13521 ( .A1(n12190), .A2(n12204), .B1(n14333), .B2(n12202), .ZN(
        n11040) );
  AOI21_X1 U13522 ( .B1(n14341), .B2(n11038), .A(n11037), .ZN(n11039) );
  OAI211_X1 U13523 ( .C1(n14347), .C2(n6573), .A(n11040), .B(n11039), .ZN(
        n11041) );
  AOI21_X1 U13524 ( .B1(n11042), .B2(n14343), .A(n11041), .ZN(n11043) );
  INV_X1 U13525 ( .A(n11043), .ZN(P3_U3161) );
  NAND2_X1 U13526 ( .A1(n10963), .A2(n11044), .ZN(n11046) );
  NAND2_X1 U13527 ( .A1(n11046), .A2(n11045), .ZN(n11047) );
  XNOR2_X1 U13528 ( .A(n11047), .B(n11666), .ZN(n11051) );
  XNOR2_X1 U13529 ( .A(n11048), .B(n6819), .ZN(n15004) );
  NAND2_X1 U13530 ( .A1(n15004), .A2(n14978), .ZN(n11050) );
  AOI22_X1 U13531 ( .A1(n14946), .A2(n12203), .B1(n14371), .B2(n14944), .ZN(
        n11049) );
  OAI211_X1 U13532 ( .C1(n11051), .C2(n14949), .A(n11050), .B(n11049), .ZN(
        n15009) );
  INV_X1 U13533 ( .A(n15009), .ZN(n11058) );
  NAND2_X1 U13534 ( .A1(n11052), .A2(n14980), .ZN(n15005) );
  NOR2_X1 U13535 ( .A1(n11053), .A2(n15005), .ZN(n11056) );
  OAI22_X1 U13536 ( .A1(n14955), .A2(n10473), .B1(n11054), .B2(n14926), .ZN(
        n11055) );
  AOI211_X1 U13537 ( .C1(n15004), .C2(n14953), .A(n11056), .B(n11055), .ZN(
        n11057) );
  OAI21_X1 U13538 ( .B1(n11058), .B2(n14957), .A(n11057), .ZN(P3_U3224) );
  NAND2_X1 U13539 ( .A1(n10963), .A2(n11059), .ZN(n11061) );
  NAND2_X1 U13540 ( .A1(n11061), .A2(n11060), .ZN(n11063) );
  XNOR2_X1 U13541 ( .A(n11063), .B(n11062), .ZN(n11064) );
  NAND2_X1 U13542 ( .A1(n11064), .A2(n14934), .ZN(n11066) );
  AOI22_X1 U13543 ( .A1(n14946), .A2(n12202), .B1(n12076), .B2(n14944), .ZN(
        n11065) );
  NAND2_X1 U13544 ( .A1(n11066), .A2(n11065), .ZN(n15015) );
  INV_X1 U13545 ( .A(n15015), .ZN(n11071) );
  XNOR2_X1 U13546 ( .A(n11067), .B(n11677), .ZN(n15012) );
  NOR2_X1 U13547 ( .A1(n14354), .A2(n15014), .ZN(n11069) );
  OAI22_X1 U13548 ( .A1(n14955), .A2(n10716), .B1(n12078), .B2(n14926), .ZN(
        n11068) );
  AOI211_X1 U13549 ( .C1(n15012), .C2(n14380), .A(n11069), .B(n11068), .ZN(
        n11070) );
  OAI21_X1 U13550 ( .B1(n11071), .B2(n14957), .A(n11070), .ZN(P3_U3223) );
  INV_X1 U13551 ( .A(n11888), .ZN(n11188) );
  OAI222_X1 U13552 ( .A1(P1_U3086), .A2(n11073), .B1(n14305), .B2(n11188), 
        .C1(n11072), .C2(n14302), .ZN(P1_U3334) );
  NAND2_X1 U13553 ( .A1(n11080), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11074) );
  NAND2_X1 U13554 ( .A1(n12216), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12207) );
  OAI21_X1 U13555 ( .B1(n12216), .B2(P3_REG1_REG_12__SCAN_IN), .A(n12207), 
        .ZN(n11078) );
  INV_X1 U13556 ( .A(n12208), .ZN(n11077) );
  AOI21_X1 U13557 ( .B1(n11079), .B2(n11078), .A(n11077), .ZN(n11098) );
  NAND2_X1 U13558 ( .A1(n11080), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n11081) );
  NOR2_X1 U13559 ( .A1(n6995), .A2(n11083), .ZN(n11084) );
  NOR2_X1 U13560 ( .A1(n11084), .A2(n14863), .ZN(n12233) );
  NAND2_X1 U13561 ( .A1(n12216), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12234) );
  OAI21_X1 U13562 ( .B1(n12216), .B2(P3_REG2_REG_12__SCAN_IN), .A(n12234), 
        .ZN(n12232) );
  XNOR2_X1 U13563 ( .A(n12233), .B(n12232), .ZN(n11088) );
  INV_X1 U13564 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11085) );
  OR2_X1 U13565 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11085), .ZN(n11247) );
  OAI21_X1 U13566 ( .B1(n14883), .B2(n15285), .A(n11247), .ZN(n11087) );
  NOR2_X1 U13567 ( .A1(n14885), .A2(n12216), .ZN(n11086) );
  AOI211_X1 U13568 ( .C1(n12307), .C2(n11088), .A(n11087), .B(n11086), .ZN(
        n11097) );
  MUX2_X1 U13569 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12691), .Z(n11092) );
  INV_X1 U13570 ( .A(n11092), .ZN(n11093) );
  INV_X1 U13571 ( .A(n11089), .ZN(n11090) );
  NOR2_X1 U13572 ( .A1(n11091), .A2(n11090), .ZN(n14869) );
  XNOR2_X1 U13573 ( .A(n11092), .B(n14866), .ZN(n14868) );
  NOR2_X1 U13574 ( .A1(n14869), .A2(n14868), .ZN(n14867) );
  AOI21_X1 U13575 ( .B1(n6995), .B2(n11093), .A(n14867), .ZN(n11095) );
  MUX2_X1 U13576 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12691), .Z(n12217) );
  XOR2_X1 U13577 ( .A(n12217), .B(n12216), .Z(n11094) );
  NAND2_X1 U13578 ( .A1(n11095), .A2(n11094), .ZN(n14892) );
  OAI211_X1 U13579 ( .C1(n11095), .C2(n11094), .A(n14892), .B(n14893), .ZN(
        n11096) );
  OAI211_X1 U13580 ( .C1(n11098), .C2(n14897), .A(n11097), .B(n11096), .ZN(
        P3_U3194) );
  OR2_X1 U13581 ( .A1(n14504), .A2(n13848), .ZN(n11099) );
  OAI21_X1 U13582 ( .B1(n11102), .B2(n11101), .A(n11197), .ZN(n11253) );
  INV_X1 U13583 ( .A(n13848), .ZN(n13589) );
  OAI22_X1 U13584 ( .A1(n13589), .A2(n14136), .B1(n14427), .B2(n14138), .ZN(
        n11109) );
  OR2_X1 U13585 ( .A1(n14504), .A2(n13589), .ZN(n11105) );
  NAND2_X1 U13586 ( .A1(n11106), .A2(n11105), .ZN(n11190) );
  XNOR2_X1 U13587 ( .A(n11190), .B(n11189), .ZN(n11107) );
  NOR2_X1 U13588 ( .A1(n11107), .A2(n14275), .ZN(n11108) );
  AOI211_X1 U13589 ( .C1(n14057), .C2(n11253), .A(n11109), .B(n11108), .ZN(
        n11256) );
  INV_X1 U13590 ( .A(n11200), .ZN(n11110) );
  AOI21_X1 U13591 ( .B1(n13601), .B2(n11111), .A(n11110), .ZN(n11254) );
  NOR2_X1 U13592 ( .A1(n7016), .A2(n14161), .ZN(n11114) );
  OAI22_X1 U13593 ( .A1(n14076), .A2(n11112), .B1(n13764), .B2(n14106), .ZN(
        n11113) );
  AOI211_X1 U13594 ( .C1(n11254), .C2(n14167), .A(n11114), .B(n11113), .ZN(
        n11116) );
  NAND2_X1 U13595 ( .A1(n11253), .A2(n14064), .ZN(n11115) );
  OAI211_X1 U13596 ( .C1(n11256), .C2(n14159), .A(n11116), .B(n11115), .ZN(
        P1_U3281) );
  XNOR2_X1 U13597 ( .A(n15014), .B(n12046), .ZN(n11121) );
  XNOR2_X1 U13598 ( .A(n11121), .B(n14371), .ZN(n12073) );
  INV_X1 U13599 ( .A(n12202), .ZN(n11119) );
  INV_X1 U13600 ( .A(n11117), .ZN(n11118) );
  NAND2_X1 U13601 ( .A1(n11119), .A2(n11118), .ZN(n12070) );
  AND2_X1 U13602 ( .A1(n12073), .A2(n12070), .ZN(n11120) );
  INV_X1 U13603 ( .A(n11121), .ZN(n11122) );
  NAND2_X1 U13604 ( .A1(n11122), .A2(n14371), .ZN(n11123) );
  XNOR2_X1 U13605 ( .A(n11130), .B(n6517), .ZN(n11124) );
  NAND2_X1 U13606 ( .A1(n11125), .A2(n11124), .ZN(n11241) );
  NAND2_X1 U13607 ( .A1(n11242), .A2(n11241), .ZN(n11126) );
  XNOR2_X1 U13608 ( .A(n11126), .B(n11318), .ZN(n11132) );
  AND2_X1 U13609 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n14877) );
  AOI21_X1 U13610 ( .B1(n14333), .B2(n14372), .A(n14877), .ZN(n11128) );
  NAND2_X1 U13611 ( .A1(n12190), .A2(n14371), .ZN(n11127) );
  OAI211_X1 U13612 ( .C1(n14347), .C2(n14374), .A(n11128), .B(n11127), .ZN(
        n11129) );
  AOI21_X1 U13613 ( .B1(n11130), .B2(n14341), .A(n11129), .ZN(n11131) );
  OAI21_X1 U13614 ( .B1(n11132), .B2(n12174), .A(n11131), .ZN(P3_U3176) );
  INV_X1 U13615 ( .A(n13065), .ZN(n11133) );
  NAND2_X1 U13616 ( .A1(n14844), .A2(n11133), .ZN(n11134) );
  INV_X1 U13617 ( .A(n13064), .ZN(n11136) );
  OR2_X1 U13618 ( .A1(n12880), .A2(n11136), .ZN(n11212) );
  NAND2_X1 U13619 ( .A1(n12880), .A2(n11136), .ZN(n11137) );
  NAND2_X1 U13620 ( .A1(n11212), .A2(n11137), .ZN(n13021) );
  AOI21_X1 U13621 ( .B1(n11138), .B2(n13021), .A(n13369), .ZN(n11142) );
  INV_X1 U13622 ( .A(n13021), .ZN(n11139) );
  AOI21_X1 U13623 ( .B1(n11142), .B2(n11213), .A(n11141), .ZN(n11230) );
  INV_X1 U13624 ( .A(n12880), .ZN(n11231) );
  OAI211_X1 U13625 ( .C1(n11231), .C2(n11143), .A(n10803), .B(n11222), .ZN(
        n11229) );
  INV_X1 U13626 ( .A(n11229), .ZN(n11147) );
  AOI22_X1 U13627 ( .A1(n14811), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11144), 
        .B2(n14783), .ZN(n11145) );
  OAI21_X1 U13628 ( .B1(n11231), .B2(n13390), .A(n11145), .ZN(n11146) );
  AOI21_X1 U13629 ( .B1(n11147), .B2(n13425), .A(n11146), .ZN(n11152) );
  AND2_X1 U13630 ( .A1(n14844), .A2(n13065), .ZN(n11149) );
  OR2_X1 U13631 ( .A1(n14844), .A2(n13065), .ZN(n11148) );
  XNOR2_X1 U13632 ( .A(n11211), .B(n13021), .ZN(n11233) );
  NAND2_X1 U13633 ( .A1(n11233), .A2(n14792), .ZN(n11151) );
  OAI211_X1 U13634 ( .C1(n11230), .C2(n14811), .A(n11152), .B(n11151), .ZN(
        P2_U3253) );
  NAND2_X1 U13635 ( .A1(n11154), .A2(n11153), .ZN(n11155) );
  AOI22_X1 U13636 ( .A1(n14616), .A2(n13697), .B1(n10343), .B2(n13850), .ZN(
        n11338) );
  NAND2_X1 U13637 ( .A1(n14616), .A2(n13702), .ZN(n11158) );
  NAND2_X1 U13638 ( .A1(n13850), .A2(n13697), .ZN(n11157) );
  NAND2_X1 U13639 ( .A1(n11158), .A2(n11157), .ZN(n11159) );
  XNOR2_X1 U13640 ( .A(n11159), .B(n13705), .ZN(n11337) );
  XOR2_X1 U13641 ( .A(n11338), .B(n11337), .Z(n11160) );
  AOI21_X1 U13642 ( .B1(n11161), .B2(n11160), .A(n11340), .ZN(n11168) );
  OAI21_X1 U13643 ( .B1(n14471), .B2(n14469), .A(n11162), .ZN(n11163) );
  AOI21_X1 U13644 ( .B1(n14459), .B2(n13851), .A(n11163), .ZN(n11164) );
  OAI21_X1 U13645 ( .B1(n11165), .B2(n14485), .A(n11164), .ZN(n11166) );
  AOI21_X1 U13646 ( .B1(n14616), .B2(n14481), .A(n11166), .ZN(n11167) );
  OAI21_X1 U13647 ( .B1(n11168), .B2(n14476), .A(n11167), .ZN(P1_U3231) );
  XNOR2_X1 U13648 ( .A(n11175), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14772) );
  INV_X1 U13649 ( .A(n14772), .ZN(n11172) );
  INV_X1 U13650 ( .A(n11169), .ZN(n11170) );
  AOI21_X1 U13651 ( .B1(n11517), .B2(P2_REG1_REG_16__SCAN_IN), .A(n11170), 
        .ZN(n14771) );
  INV_X1 U13652 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11171) );
  OAI22_X1 U13653 ( .A1(n11172), .A2(n14771), .B1(n11175), .B2(n11171), .ZN(
        n13127) );
  XOR2_X1 U13654 ( .A(n13128), .B(n13127), .Z(n11173) );
  NAND2_X1 U13655 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11173), .ZN(n13129) );
  OAI21_X1 U13656 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n11173), .A(n13129), 
        .ZN(n11187) );
  NAND2_X1 U13657 ( .A1(n14769), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11180) );
  INV_X1 U13658 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U13659 ( .A1(n11175), .A2(n11174), .ZN(n11176) );
  AND2_X1 U13660 ( .A1(n11176), .A2(n11180), .ZN(n14778) );
  OAI21_X1 U13661 ( .B1(n11179), .B2(n11178), .A(n11177), .ZN(n14777) );
  NAND2_X1 U13662 ( .A1(n14778), .A2(n14777), .ZN(n14775) );
  NAND2_X1 U13663 ( .A1(n11180), .A2(n14775), .ZN(n13123) );
  XNOR2_X1 U13664 ( .A(n13128), .B(n13123), .ZN(n11181) );
  NOR2_X1 U13665 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11181), .ZN(n13124) );
  AOI21_X1 U13666 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n11181), .A(n13124), 
        .ZN(n11182) );
  INV_X1 U13667 ( .A(n14776), .ZN(n14738) );
  OR2_X1 U13668 ( .A1(n11182), .A2(n14738), .ZN(n11186) );
  AND2_X1 U13669 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n12781) );
  NOR2_X1 U13670 ( .A1(n14740), .A2(n11183), .ZN(n11184) );
  AOI211_X1 U13671 ( .C1(n14768), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n12781), 
        .B(n11184), .ZN(n11185) );
  OAI211_X1 U13672 ( .C1(n11187), .C2(n14747), .A(n11186), .B(n11185), .ZN(
        P2_U3232) );
  NAND2_X1 U13673 ( .A1(n11190), .A2(n11189), .ZN(n11192) );
  INV_X1 U13674 ( .A(n13847), .ZN(n14472) );
  OR2_X1 U13675 ( .A1(n13601), .A2(n14472), .ZN(n11191) );
  NAND2_X1 U13676 ( .A1(n11192), .A2(n11191), .ZN(n11309) );
  XNOR2_X1 U13677 ( .A(n11309), .B(n11308), .ZN(n11195) );
  NAND2_X1 U13678 ( .A1(n13847), .A2(n14154), .ZN(n11193) );
  OAI21_X1 U13679 ( .B1(n13833), .B2(n14138), .A(n11193), .ZN(n11194) );
  AOI21_X1 U13680 ( .B1(n11195), .B2(n14264), .A(n11194), .ZN(n14502) );
  NOR2_X1 U13681 ( .A1(n11198), .A2(n11308), .ZN(n11199) );
  OR2_X1 U13682 ( .A1(n11301), .A2(n11199), .ZN(n14500) );
  INV_X1 U13683 ( .A(n11305), .ZN(n11304) );
  NAND2_X1 U13684 ( .A1(n13610), .A2(n11200), .ZN(n11201) );
  NAND2_X1 U13685 ( .A1(n11304), .A2(n11201), .ZN(n14498) );
  OAI22_X1 U13686 ( .A1(n14076), .A2(n11202), .B1(n13797), .B2(n14106), .ZN(
        n11203) );
  AOI21_X1 U13687 ( .B1(n13610), .B2(n14110), .A(n11203), .ZN(n11204) );
  OAI21_X1 U13688 ( .B1(n14498), .B2(n14112), .A(n11204), .ZN(n11205) );
  AOI21_X1 U13689 ( .B1(n14500), .B2(n14114), .A(n11205), .ZN(n11206) );
  OAI21_X1 U13690 ( .B1(n14502), .B2(n14159), .A(n11206), .ZN(P1_U3280) );
  NAND2_X1 U13691 ( .A1(n11207), .A2(n12963), .ZN(n11209) );
  AOI22_X1 U13692 ( .A1(n11862), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n11861), 
        .B2(n14751), .ZN(n11208) );
  XNOR2_X1 U13693 ( .A(n14658), .B(n13063), .ZN(n13023) );
  NOR2_X1 U13694 ( .A1(n12880), .A2(n13064), .ZN(n11210) );
  XOR2_X1 U13695 ( .A(n13023), .B(n11404), .Z(n13528) );
  OAI211_X1 U13696 ( .C1(n11214), .C2(n13023), .A(n11374), .B(n14798), .ZN(
        n11220) );
  INV_X1 U13697 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11215) );
  XNOR2_X1 U13698 ( .A(n11388), .B(n11215), .ZN(n14426) );
  INV_X1 U13699 ( .A(n14426), .ZN(n11444) );
  NAND2_X1 U13700 ( .A1(n12004), .A2(n11444), .ZN(n11219) );
  NAND2_X1 U13701 ( .A1(n12941), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11218) );
  NAND2_X1 U13702 ( .A1(n12959), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n11217) );
  NAND2_X1 U13703 ( .A1(n12958), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11216) );
  NAND4_X1 U13704 ( .A1(n11219), .A2(n11218), .A3(n11217), .A4(n11216), .ZN(
        n13062) );
  AOI22_X1 U13705 ( .A1(n13405), .A2(n13064), .B1(n13062), .B2(n13407), .ZN(
        n14650) );
  NAND2_X1 U13706 ( .A1(n11220), .A2(n14650), .ZN(n13525) );
  INV_X1 U13707 ( .A(n14658), .ZN(n11226) );
  INV_X1 U13708 ( .A(n11443), .ZN(n11221) );
  AOI211_X1 U13709 ( .C1(n14658), .C2(n11222), .A(n9459), .B(n11221), .ZN(
        n13526) );
  NAND2_X1 U13710 ( .A1(n13526), .A2(n13425), .ZN(n11225) );
  AOI22_X1 U13711 ( .A1(n14811), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11223), 
        .B2(n14783), .ZN(n11224) );
  OAI211_X1 U13712 ( .C1(n11226), .C2(n13390), .A(n11225), .B(n11224), .ZN(
        n11227) );
  AOI21_X1 U13713 ( .B1(n13525), .B2(n14809), .A(n11227), .ZN(n11228) );
  OAI21_X1 U13714 ( .B1(n13528), .B2(n13396), .A(n11228), .ZN(P2_U3252) );
  OAI211_X1 U13715 ( .C1(n11231), .C2(n14837), .A(n11230), .B(n11229), .ZN(
        n11232) );
  AOI21_X1 U13716 ( .B1(n14833), .B2(n11233), .A(n11232), .ZN(n11236) );
  NAND2_X1 U13717 ( .A1(n13539), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n11234) );
  OAI21_X1 U13718 ( .B1(n11236), .B2(n13539), .A(n11234), .ZN(P2_U3466) );
  NAND2_X1 U13719 ( .A1(n13449), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11235) );
  OAI21_X1 U13720 ( .B1(n11236), .B2(n13449), .A(n11235), .ZN(P2_U3511) );
  XNOR2_X1 U13721 ( .A(n14393), .B(n12046), .ZN(n11238) );
  NAND2_X1 U13722 ( .A1(n11238), .A2(n11237), .ZN(n11262) );
  INV_X1 U13723 ( .A(n11238), .ZN(n11239) );
  NAND2_X1 U13724 ( .A1(n11239), .A2(n14372), .ZN(n11240) );
  AND2_X1 U13725 ( .A1(n11262), .A2(n11240), .ZN(n11245) );
  NAND2_X1 U13726 ( .A1(n11241), .A2(n11318), .ZN(n11243) );
  OAI21_X1 U13727 ( .B1(n11245), .B2(n11244), .A(n11263), .ZN(n11246) );
  NAND2_X1 U13728 ( .A1(n11246), .A2(n14343), .ZN(n11252) );
  INV_X1 U13729 ( .A(n11324), .ZN(n11250) );
  NAND2_X1 U13730 ( .A1(n12190), .A2(n12076), .ZN(n11248) );
  OAI211_X1 U13731 ( .C1(n11432), .C2(n12192), .A(n11248), .B(n11247), .ZN(
        n11249) );
  AOI21_X1 U13732 ( .B1(n12195), .B2(n11250), .A(n11249), .ZN(n11251) );
  OAI211_X1 U13733 ( .C1(n12198), .C2(n14393), .A(n11252), .B(n11251), .ZN(
        P3_U3164) );
  INV_X1 U13734 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11259) );
  INV_X1 U13735 ( .A(n11253), .ZN(n11257) );
  AOI22_X1 U13736 ( .A1(n11254), .A2(n14618), .B1(n14617), .B2(n13601), .ZN(
        n11255) );
  OAI211_X1 U13737 ( .C1(n11257), .C2(n14219), .A(n11256), .B(n11255), .ZN(
        n11260) );
  NAND2_X1 U13738 ( .A1(n11260), .A2(n14627), .ZN(n11258) );
  OAI21_X1 U13739 ( .B1(n14627), .B2(n11259), .A(n11258), .ZN(P1_U3495) );
  NAND2_X1 U13740 ( .A1(n11260), .A2(n14636), .ZN(n11261) );
  OAI21_X1 U13741 ( .B1(n14636), .B2(n7947), .A(n11261), .ZN(P1_U3540) );
  XNOR2_X1 U13742 ( .A(n14366), .B(n12095), .ZN(n11264) );
  AND2_X1 U13743 ( .A1(n11264), .A2(n11432), .ZN(n11360) );
  INV_X1 U13744 ( .A(n11360), .ZN(n11266) );
  INV_X1 U13745 ( .A(n11264), .ZN(n11265) );
  NAND2_X1 U13746 ( .A1(n11265), .A2(n12201), .ZN(n11359) );
  NAND2_X1 U13747 ( .A1(n11266), .A2(n11359), .ZN(n11267) );
  XNOR2_X1 U13748 ( .A(n11361), .B(n11267), .ZN(n11272) );
  AND2_X1 U13749 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n14901) );
  NOR2_X1 U13750 ( .A1(n14337), .A2(n12192), .ZN(n11268) );
  AOI211_X1 U13751 ( .C1(n12190), .C2(n14372), .A(n14901), .B(n11268), .ZN(
        n11269) );
  OAI21_X1 U13752 ( .B1(n14362), .B2(n14347), .A(n11269), .ZN(n11270) );
  AOI21_X1 U13753 ( .B1(n14366), .B2(n14341), .A(n11270), .ZN(n11271) );
  OAI21_X1 U13754 ( .B1(n11272), .B2(n12174), .A(n11271), .ZN(P3_U3174) );
  INV_X1 U13755 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n11299) );
  NAND2_X1 U13756 ( .A1(n11273), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11278) );
  INV_X1 U13757 ( .A(n11274), .ZN(n11275) );
  NAND2_X1 U13758 ( .A1(n11276), .A2(n11275), .ZN(n11277) );
  NAND2_X1 U13759 ( .A1(n11278), .A2(n11277), .ZN(n11279) );
  XOR2_X1 U13760 ( .A(n11286), .B(n11279), .Z(n14564) );
  NAND2_X1 U13761 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14564), .ZN(n14562) );
  NAND2_X1 U13762 ( .A1(n11279), .A2(n11286), .ZN(n11280) );
  NAND2_X1 U13763 ( .A1(n14562), .A2(n11280), .ZN(n11281) );
  XOR2_X1 U13764 ( .A(n11281), .B(P1_REG2_REG_19__SCAN_IN), .Z(n11294) );
  INV_X1 U13765 ( .A(n11294), .ZN(n11292) );
  OAI22_X1 U13766 ( .A1(n11285), .A2(n11284), .B1(n11283), .B2(n11282), .ZN(
        n11287) );
  XOR2_X1 U13767 ( .A(n11286), .B(n11287), .Z(n14567) );
  NAND2_X1 U13768 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14567), .ZN(n14565) );
  NAND2_X1 U13769 ( .A1(n11287), .A2(n11286), .ZN(n11288) );
  NAND2_X1 U13770 ( .A1(n14565), .A2(n11288), .ZN(n11290) );
  XNOR2_X1 U13771 ( .A(n11290), .B(n11289), .ZN(n11293) );
  OAI21_X1 U13772 ( .B1(n11293), .B2(n14557), .A(n14571), .ZN(n11291) );
  AOI21_X1 U13773 ( .B1(n14563), .B2(n11292), .A(n11291), .ZN(n11297) );
  AOI22_X1 U13774 ( .A1(n11294), .A2(n14563), .B1(n11293), .B2(n14566), .ZN(
        n11296) );
  MUX2_X1 U13775 ( .A(n11297), .B(n11296), .S(n11295), .Z(n11298) );
  NAND2_X1 U13776 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13729)
         );
  OAI211_X1 U13777 ( .C1(n11299), .C2(n14575), .A(n11298), .B(n13729), .ZN(
        P1_U3262) );
  OAI21_X1 U13778 ( .B1(n11302), .B2(n6959), .A(n11413), .ZN(n14491) );
  OAI22_X1 U13779 ( .A1(n14076), .A2(n11303), .B1(n14439), .B2(n14106), .ZN(
        n11307) );
  INV_X1 U13780 ( .A(n14436), .ZN(n14492) );
  OAI21_X1 U13781 ( .B1(n14492), .B2(n11305), .A(n11420), .ZN(n14493) );
  NOR2_X1 U13782 ( .A1(n14493), .A2(n14112), .ZN(n11306) );
  AOI211_X1 U13783 ( .C1(n14110), .C2(n14436), .A(n11307), .B(n11306), .ZN(
        n11316) );
  NAND2_X1 U13784 ( .A1(n11309), .A2(n7407), .ZN(n11311) );
  OR2_X1 U13785 ( .A1(n13610), .A2(n14427), .ZN(n11310) );
  XNOR2_X1 U13786 ( .A(n11416), .B(n6959), .ZN(n11312) );
  NAND2_X1 U13787 ( .A1(n11312), .A2(n14264), .ZN(n11314) );
  INV_X1 U13788 ( .A(n14441), .ZN(n13845) );
  AOI22_X1 U13789 ( .A1(n13845), .A2(n14152), .B1(n14154), .B2(n13846), .ZN(
        n11313) );
  NAND2_X1 U13790 ( .A1(n11314), .A2(n11313), .ZN(n14494) );
  NAND2_X1 U13791 ( .A1(n14494), .A2(n14076), .ZN(n11315) );
  OAI211_X1 U13792 ( .C1(n14491), .C2(n14164), .A(n11316), .B(n11315), .ZN(
        P1_U3279) );
  AOI21_X1 U13793 ( .B1(n11317), .B2(n11799), .A(n14949), .ZN(n11321) );
  OAI22_X1 U13794 ( .A1(n11318), .A2(n14932), .B1(n11432), .B2(n14930), .ZN(
        n11319) );
  AOI21_X1 U13795 ( .B1(n11321), .B2(n11320), .A(n11319), .ZN(n14394) );
  OAI21_X1 U13796 ( .B1(n11323), .B2(n11799), .A(n11322), .ZN(n14397) );
  NOR2_X1 U13797 ( .A1(n14354), .A2(n14393), .ZN(n11327) );
  OAI22_X1 U13798 ( .A1(n14955), .A2(n11325), .B1(n11324), .B2(n14926), .ZN(
        n11326) );
  AOI211_X1 U13799 ( .C1(n14397), .C2(n14380), .A(n11327), .B(n11326), .ZN(
        n11328) );
  OAI21_X1 U13800 ( .B1(n14957), .B2(n14394), .A(n11328), .ZN(P3_U3221) );
  INV_X1 U13801 ( .A(n11329), .ZN(n11330) );
  OAI222_X1 U13802 ( .A1(P3_U3151), .A2(n11332), .B1(n12698), .B2(n11331), 
        .C1(n12694), .C2(n11330), .ZN(P3_U3271) );
  INV_X1 U13803 ( .A(n11930), .ZN(n11609) );
  OAI222_X1 U13804 ( .A1(n13580), .A2(n11931), .B1(n13578), .B2(n11609), .C1(
        P2_U3088), .C2(n11333), .ZN(P2_U3303) );
  XNOR2_X1 U13805 ( .A(n11335), .B(n11334), .ZN(n11899) );
  INV_X1 U13806 ( .A(n11899), .ZN(n11336) );
  OAI222_X1 U13807 ( .A1(n13580), .A2(n15205), .B1(n13578), .B2(n11336), .C1(
        n12968), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U13808 ( .A(n11337), .ZN(n11339) );
  NAND2_X1 U13809 ( .A1(n11345), .A2(n13702), .ZN(n11342) );
  NAND2_X1 U13810 ( .A1(n13849), .A2(n13697), .ZN(n11341) );
  NAND2_X1 U13811 ( .A1(n11342), .A2(n11341), .ZN(n11343) );
  XNOR2_X1 U13812 ( .A(n11343), .B(n13705), .ZN(n13593) );
  NOR2_X1 U13813 ( .A1(n14469), .A2(n13740), .ZN(n11344) );
  AOI21_X1 U13814 ( .B1(n11345), .B2(n13697), .A(n11344), .ZN(n13591) );
  XNOR2_X1 U13815 ( .A(n13593), .B(n13591), .ZN(n11346) );
  OAI211_X1 U13816 ( .C1(n11347), .C2(n11346), .A(n13595), .B(n14464), .ZN(
        n11353) );
  INV_X1 U13817 ( .A(n13808), .ZN(n13825) );
  NOR2_X1 U13818 ( .A1(n14485), .A2(n11348), .ZN(n11349) );
  AOI211_X1 U13819 ( .C1(n13825), .C2(n11351), .A(n11350), .B(n11349), .ZN(
        n11352) );
  OAI211_X1 U13820 ( .C1(n6948), .C2(n14461), .A(n11353), .B(n11352), .ZN(
        P1_U3217) );
  NAND2_X1 U13821 ( .A1(n11914), .A2(n14296), .ZN(n11355) );
  OAI211_X1 U13822 ( .C1(n11356), .C2(n14302), .A(n11355), .B(n11354), .ZN(
        P1_U3332) );
  NAND2_X1 U13823 ( .A1(n11914), .A2(n13564), .ZN(n11358) );
  OR2_X1 U13824 ( .A1(n11357), .A2(P2_U3088), .ZN(n13046) );
  OAI211_X1 U13825 ( .C1(n11915), .C2(n13580), .A(n11358), .B(n13046), .ZN(
        P2_U3304) );
  XNOR2_X1 U13826 ( .A(n12614), .B(n12095), .ZN(n11486) );
  XNOR2_X1 U13827 ( .A(n11486), .B(n14337), .ZN(n11488) );
  XOR2_X1 U13828 ( .A(n11488), .B(n11489), .Z(n11366) );
  AOI22_X1 U13829 ( .A1(n14333), .A2(n12537), .B1(P3_REG3_REG_14__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11363) );
  NAND2_X1 U13830 ( .A1(n12190), .A2(n12201), .ZN(n11362) );
  OAI211_X1 U13831 ( .C1(n14347), .C2(n11433), .A(n11363), .B(n11362), .ZN(
        n11364) );
  AOI21_X1 U13832 ( .B1(n12614), .B2(n14341), .A(n11364), .ZN(n11365) );
  OAI21_X1 U13833 ( .B1(n11366), .B2(n12174), .A(n11365), .ZN(P3_U3155) );
  INV_X1 U13834 ( .A(n11367), .ZN(n11368) );
  OAI222_X1 U13835 ( .A1(P3_U3151), .A2(n11369), .B1(n12698), .B2(n15275), 
        .C1(n12694), .C2(n11368), .ZN(P3_U3270) );
  INV_X1 U13836 ( .A(n11945), .ZN(n11371) );
  OAI222_X1 U13837 ( .A1(n13580), .A2(n15291), .B1(n13578), .B2(n11371), .C1(
        P2_U3088), .C2(n11370), .ZN(P2_U3302) );
  OAI222_X1 U13838 ( .A1(n11372), .A2(P1_U3086), .B1(n14305), .B2(n11371), 
        .C1(n15151), .C2(n14302), .ZN(P1_U3330) );
  INV_X1 U13839 ( .A(n13063), .ZN(n14417) );
  OR2_X1 U13840 ( .A1(n14658), .A2(n14417), .ZN(n11373) );
  OR2_X1 U13841 ( .A1(n11376), .A2(n11375), .ZN(n11379) );
  AOI22_X1 U13842 ( .A1(n11862), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n11861), 
        .B2(n11377), .ZN(n11378) );
  INV_X1 U13843 ( .A(n13062), .ZN(n11381) );
  NAND2_X1 U13844 ( .A1(n13521), .A2(n11381), .ZN(n11380) );
  OR2_X1 U13845 ( .A1(n13521), .A2(n11381), .ZN(n11382) );
  NAND2_X1 U13846 ( .A1(n11383), .A2(n12963), .ZN(n11385) );
  AOI22_X1 U13847 ( .A1(n11862), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n11861), 
        .B2(n14759), .ZN(n11384) );
  INV_X1 U13848 ( .A(n11388), .ZN(n11386) );
  AOI21_X1 U13849 ( .B1(n11386), .B2(P2_REG3_REG_14__SCAN_IN), .A(
        P2_REG3_REG_15__SCAN_IN), .ZN(n11389) );
  NAND2_X1 U13850 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n11387) );
  NOR2_X1 U13851 ( .A1(n11389), .A2(n11395), .ZN(n12799) );
  NAND2_X1 U13852 ( .A1(n12799), .A2(n12004), .ZN(n11393) );
  NAND2_X1 U13853 ( .A1(n12958), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n11392) );
  NAND2_X1 U13854 ( .A1(n12941), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11391) );
  NAND2_X1 U13855 ( .A1(n12959), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n11390) );
  XNOR2_X1 U13856 ( .A(n11543), .B(n11557), .ZN(n11394) );
  NAND2_X1 U13857 ( .A1(n11394), .A2(n14798), .ZN(n11402) );
  NOR2_X1 U13858 ( .A1(n11395), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11396) );
  OR2_X1 U13859 ( .A1(n11534), .A2(n11396), .ZN(n13402) );
  NAND2_X1 U13860 ( .A1(n12958), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11398) );
  NAND2_X1 U13861 ( .A1(n11977), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11397) );
  AND2_X1 U13862 ( .A1(n11398), .A2(n11397), .ZN(n11400) );
  NAND2_X1 U13863 ( .A1(n12959), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n11399) );
  OAI211_X1 U13864 ( .C1(n13402), .C2(n11887), .A(n11400), .B(n11399), .ZN(
        n13061) );
  AOI22_X1 U13865 ( .A1(n13061), .A2(n13407), .B1(n13062), .B2(n13405), .ZN(
        n11401) );
  AND2_X1 U13866 ( .A1(n11402), .A2(n11401), .ZN(n11504) );
  OR2_X1 U13867 ( .A1(n14658), .A2(n13063), .ZN(n11403) );
  NAND2_X1 U13868 ( .A1(n11404), .A2(n11403), .ZN(n11406) );
  NAND2_X1 U13869 ( .A1(n14658), .A2(n13063), .ZN(n11405) );
  NAND2_X1 U13870 ( .A1(n11406), .A2(n11405), .ZN(n11446) );
  NAND2_X1 U13871 ( .A1(n13521), .A2(n13062), .ZN(n11438) );
  INV_X1 U13872 ( .A(n11438), .ZN(n11407) );
  OR2_X1 U13873 ( .A1(n13521), .A2(n13062), .ZN(n11439) );
  OAI21_X2 U13874 ( .B1(n11446), .B2(n11407), .A(n11439), .ZN(n11558) );
  XNOR2_X1 U13875 ( .A(n11558), .B(n11557), .ZN(n11502) );
  AOI21_X1 U13876 ( .B1(n12897), .B2(n11442), .A(n9459), .ZN(n11408) );
  AND2_X1 U13877 ( .A1(n11408), .A2(n13401), .ZN(n11501) );
  NAND2_X1 U13878 ( .A1(n11501), .A2(n13425), .ZN(n11410) );
  AOI22_X1 U13879 ( .A1(n14811), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12799), 
        .B2(n14783), .ZN(n11409) );
  OAI211_X1 U13880 ( .C1(n6846), .C2(n13390), .A(n11410), .B(n11409), .ZN(
        n11411) );
  AOI21_X1 U13881 ( .B1(n11502), .B2(n14792), .A(n11411), .ZN(n11412) );
  OAI21_X1 U13882 ( .B1(n11504), .B2(n14811), .A(n11412), .ZN(P2_U3250) );
  XNOR2_X1 U13883 ( .A(n11459), .B(n11458), .ZN(n14490) );
  INV_X1 U13884 ( .A(n14490), .ZN(n11427) );
  XNOR2_X1 U13885 ( .A(n11457), .B(n11458), .ZN(n11417) );
  NAND2_X1 U13886 ( .A1(n11417), .A2(n14264), .ZN(n11419) );
  AOI22_X1 U13887 ( .A1(n6793), .A2(n14154), .B1(n14152), .B2(n14458), .ZN(
        n11418) );
  NAND2_X1 U13888 ( .A1(n11419), .A2(n11418), .ZN(n14488) );
  INV_X1 U13889 ( .A(n13622), .ZN(n14486) );
  INV_X1 U13890 ( .A(n11420), .ZN(n11422) );
  NOR2_X1 U13891 ( .A1(n13622), .A2(n11420), .ZN(n11462) );
  INV_X1 U13892 ( .A(n11462), .ZN(n11421) );
  OAI21_X1 U13893 ( .B1(n14486), .B2(n11422), .A(n11421), .ZN(n14487) );
  AOI22_X1 U13894 ( .A1(n14159), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13836), 
        .B2(n14157), .ZN(n11424) );
  NAND2_X1 U13895 ( .A1(n13622), .A2(n14110), .ZN(n11423) );
  OAI211_X1 U13896 ( .C1(n14487), .C2(n14112), .A(n11424), .B(n11423), .ZN(
        n11425) );
  AOI21_X1 U13897 ( .B1(n14488), .B2(n14076), .A(n11425), .ZN(n11426) );
  OAI21_X1 U13898 ( .B1(n11427), .B2(n14164), .A(n11426), .ZN(P1_U3278) );
  INV_X1 U13899 ( .A(n11430), .ZN(n11800) );
  XNOR2_X1 U13900 ( .A(n11428), .B(n11800), .ZN(n12616) );
  XNOR2_X1 U13901 ( .A(n11429), .B(n11430), .ZN(n11431) );
  OAI222_X1 U13902 ( .A1(n14930), .A2(n11490), .B1(n14932), .B2(n11432), .C1(
        n11431), .C2(n14949), .ZN(n12613) );
  NAND2_X1 U13903 ( .A1(n12613), .A2(n14955), .ZN(n11436) );
  OAI22_X1 U13904 ( .A1(n14955), .A2(n12220), .B1(n11433), .B2(n14926), .ZN(
        n11434) );
  AOI21_X1 U13905 ( .B1(n12614), .B2(n14919), .A(n11434), .ZN(n11435) );
  OAI211_X1 U13906 ( .C1(n11437), .C2(n12616), .A(n11436), .B(n11435), .ZN(
        P3_U3219) );
  NAND2_X1 U13907 ( .A1(n11439), .A2(n11438), .ZN(n13025) );
  XOR2_X1 U13908 ( .A(n11440), .B(n13025), .Z(n11441) );
  AOI222_X1 U13909 ( .A1(n14798), .A2(n11441), .B1(n13063), .B2(n13405), .C1(
        n13406), .C2(n13407), .ZN(n13523) );
  AOI211_X1 U13910 ( .C1(n13521), .C2(n11443), .A(n9459), .B(n6847), .ZN(
        n13520) );
  INV_X1 U13911 ( .A(n13521), .ZN(n14416) );
  AOI22_X1 U13912 ( .A1(n14811), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11444), 
        .B2(n14783), .ZN(n11445) );
  OAI21_X1 U13913 ( .B1(n14416), .B2(n13390), .A(n11445), .ZN(n11448) );
  XOR2_X1 U13914 ( .A(n13025), .B(n11446), .Z(n13524) );
  NOR2_X1 U13915 ( .A1(n13524), .A2(n13396), .ZN(n11447) );
  AOI211_X1 U13916 ( .C1(n13520), .C2(n13425), .A(n11448), .B(n11447), .ZN(
        n11449) );
  OAI21_X1 U13917 ( .B1(n14811), .B2(n13523), .A(n11449), .ZN(P2_U3251) );
  INV_X1 U13918 ( .A(n11967), .ZN(n11452) );
  OAI222_X1 U13919 ( .A1(P1_U3086), .A2(n11450), .B1(n14305), .B2(n11452), 
        .C1(n8483), .C2(n14302), .ZN(P1_U3329) );
  OAI222_X1 U13920 ( .A1(P2_U3088), .A2(n11453), .B1(n13578), .B2(n11452), 
        .C1(n15117), .C2(n13580), .ZN(P2_U3301) );
  XNOR2_X1 U13921 ( .A(n11474), .B(n11460), .ZN(n14274) );
  INV_X1 U13922 ( .A(n11460), .ZN(n11473) );
  OAI21_X1 U13923 ( .B1(n11461), .B2(n11473), .A(n11471), .ZN(n14272) );
  NAND2_X1 U13924 ( .A1(n11462), .A2(n13631), .ZN(n11477) );
  OAI21_X1 U13925 ( .B1(n11462), .B2(n13631), .A(n11477), .ZN(n14270) );
  OR2_X1 U13926 ( .A1(n14441), .A2(n14136), .ZN(n11464) );
  NAND2_X1 U13927 ( .A1(n14440), .A2(n14152), .ZN(n11463) );
  NAND2_X1 U13928 ( .A1(n11464), .A2(n11463), .ZN(n14268) );
  INV_X1 U13929 ( .A(n14453), .ZN(n11465) );
  AOI22_X1 U13930 ( .A1(n14076), .A2(n14268), .B1(n11465), .B2(n14157), .ZN(
        n11466) );
  OAI21_X1 U13931 ( .B1(n13964), .B2(n14076), .A(n11466), .ZN(n11467) );
  AOI21_X1 U13932 ( .B1(n14450), .B2(n14110), .A(n11467), .ZN(n11468) );
  OAI21_X1 U13933 ( .B1(n14270), .B2(n14112), .A(n11468), .ZN(n11469) );
  AOI21_X1 U13934 ( .B1(n14272), .B2(n14114), .A(n11469), .ZN(n11470) );
  OAI21_X1 U13935 ( .B1(n14116), .B2(n14274), .A(n11470), .ZN(P1_U3277) );
  XNOR2_X1 U13936 ( .A(n11579), .B(n11472), .ZN(n14267) );
  INV_X1 U13937 ( .A(n11472), .ZN(n11476) );
  AOI21_X1 U13938 ( .B1(n11476), .B2(n11475), .A(n11586), .ZN(n14265) );
  INV_X1 U13939 ( .A(n11477), .ZN(n11478) );
  INV_X1 U13940 ( .A(n14259), .ZN(n14462) );
  OAI21_X1 U13941 ( .B1(n11478), .B2(n14462), .A(n6546), .ZN(n14262) );
  NOR2_X1 U13942 ( .A1(n14076), .A2(n11479), .ZN(n11481) );
  AOI22_X1 U13943 ( .A1(n14456), .A2(n14152), .B1(n14154), .B2(n14458), .ZN(
        n14261) );
  OAI22_X1 U13944 ( .A1(n14159), .A2(n14261), .B1(n14468), .B2(n14106), .ZN(
        n11480) );
  AOI211_X1 U13945 ( .C1(n14259), .C2(n14110), .A(n11481), .B(n11480), .ZN(
        n11482) );
  OAI21_X1 U13946 ( .B1(n14262), .B2(n14112), .A(n11482), .ZN(n11483) );
  AOI21_X1 U13947 ( .B1(n14265), .B2(n11484), .A(n11483), .ZN(n11485) );
  OAI21_X1 U13948 ( .B1(n14164), .B2(n14267), .A(n11485), .ZN(P1_U3276) );
  NAND2_X1 U13949 ( .A1(n11486), .A2(n14337), .ZN(n11487) );
  XNOR2_X1 U13950 ( .A(n14342), .B(n12095), .ZN(n11491) );
  XNOR2_X1 U13951 ( .A(n11491), .B(n12537), .ZN(n14339) );
  NAND2_X1 U13952 ( .A1(n11491), .A2(n11490), .ZN(n11492) );
  XNOR2_X1 U13953 ( .A(n12547), .B(n12095), .ZN(n12017) );
  XNOR2_X1 U13954 ( .A(n12017), .B(n14332), .ZN(n11494) );
  AOI21_X1 U13955 ( .B1(n11495), .B2(n11494), .A(n12174), .ZN(n11496) );
  NAND2_X1 U13956 ( .A1(n11496), .A2(n12019), .ZN(n11500) );
  NAND2_X1 U13957 ( .A1(n12190), .A2(n12537), .ZN(n11497) );
  NAND2_X1 U13958 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12274)
         );
  OAI211_X1 U13959 ( .C1(n12020), .C2(n12192), .A(n11497), .B(n12274), .ZN(
        n11498) );
  AOI21_X1 U13960 ( .B1(n12195), .B2(n12545), .A(n11498), .ZN(n11499) );
  OAI211_X1 U13961 ( .C1(n12547), .C2(n12198), .A(n11500), .B(n11499), .ZN(
        P3_U3166) );
  INV_X1 U13962 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11505) );
  AOI21_X1 U13963 ( .B1(n11502), .B2(n14833), .A(n11501), .ZN(n11503) );
  AND2_X1 U13964 ( .A1(n11504), .A2(n11503), .ZN(n11507) );
  MUX2_X1 U13965 ( .A(n11505), .B(n11507), .S(n14855), .Z(n11506) );
  OAI21_X1 U13966 ( .B1(n6846), .B2(n13556), .A(n11506), .ZN(P2_U3475) );
  MUX2_X1 U13967 ( .A(n15200), .B(n11507), .S(n14861), .Z(n11508) );
  OAI21_X1 U13968 ( .B1(n6846), .B2(n13502), .A(n11508), .ZN(P2_U3514) );
  XOR2_X1 U13969 ( .A(n11509), .B(n11802), .Z(n11510) );
  OAI222_X1 U13970 ( .A1(n14930), .A2(n12131), .B1(n14932), .B2(n14337), .C1(
        n11510), .C2(n14949), .ZN(n12608) );
  INV_X1 U13971 ( .A(n12608), .ZN(n11515) );
  XNOR2_X1 U13972 ( .A(n11511), .B(n11802), .ZN(n12609) );
  INV_X1 U13973 ( .A(n14342), .ZN(n12670) );
  NOR2_X1 U13974 ( .A1(n12670), .A2(n14354), .ZN(n11513) );
  OAI22_X1 U13975 ( .A1(n14955), .A2(n15185), .B1(n14348), .B2(n14926), .ZN(
        n11512) );
  AOI211_X1 U13976 ( .C1(n12609), .C2(n14380), .A(n11513), .B(n11512), .ZN(
        n11514) );
  OAI21_X1 U13977 ( .B1(n11515), .B2(n14957), .A(n11514), .ZN(P3_U3218) );
  NAND2_X1 U13978 ( .A1(n13061), .A2(n6520), .ZN(n11841) );
  NAND2_X1 U13979 ( .A1(n11516), .A2(n12963), .ZN(n11519) );
  AOI22_X1 U13980 ( .A1(n11862), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n11861), 
        .B2(n11517), .ZN(n11518) );
  XNOR2_X1 U13981 ( .A(n13514), .B(n11976), .ZN(n11843) );
  XOR2_X1 U13982 ( .A(n11841), .B(n11843), .Z(n11533) );
  NAND2_X1 U13983 ( .A1(n13062), .A2(n6520), .ZN(n11525) );
  INV_X1 U13984 ( .A(n11525), .ZN(n11527) );
  XNOR2_X1 U13985 ( .A(n13521), .B(n11976), .ZN(n11526) );
  AND2_X1 U13986 ( .A1(n13063), .A2(n6520), .ZN(n11522) );
  NAND2_X1 U13987 ( .A1(n11523), .A2(n11522), .ZN(n11524) );
  OAI21_X1 U13988 ( .B1(n11523), .B2(n11522), .A(n11524), .ZN(n14653) );
  XNOR2_X1 U13989 ( .A(n11526), .B(n11525), .ZN(n14413) );
  NAND2_X1 U13990 ( .A1(n14414), .A2(n14413), .ZN(n14412) );
  OAI21_X1 U13991 ( .B1(n11527), .B2(n11526), .A(n14412), .ZN(n11530) );
  XNOR2_X1 U13992 ( .A(n12897), .B(n11976), .ZN(n11528) );
  XNOR2_X1 U13993 ( .A(n11530), .B(n11528), .ZN(n12797) );
  NOR2_X1 U13994 ( .A1(n14420), .A2(n10803), .ZN(n12796) );
  NAND2_X1 U13995 ( .A1(n12797), .A2(n12796), .ZN(n12795) );
  INV_X1 U13996 ( .A(n11528), .ZN(n11529) );
  OR2_X1 U13997 ( .A1(n11530), .A2(n11529), .ZN(n11531) );
  AOI21_X1 U13998 ( .B1(n11533), .B2(n11532), .A(n12742), .ZN(n11542) );
  NOR2_X1 U13999 ( .A1(n11534), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11535) );
  OR2_X1 U14000 ( .A1(n11550), .A2(n11535), .ZN(n12744) );
  AOI22_X1 U14001 ( .A1(n12941), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n12959), 
        .B2(P2_REG0_REG_17__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U14002 ( .A1(n12958), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n11536) );
  OAI211_X1 U14003 ( .C1(n12744), .C2(n11887), .A(n11537), .B(n11536), .ZN(
        n13408) );
  INV_X1 U14004 ( .A(n13408), .ZN(n12902) );
  OAI21_X1 U14005 ( .B1(n14419), .B2(n12902), .A(n11538), .ZN(n11540) );
  OAI22_X1 U14006 ( .A1(n14418), .A2(n14420), .B1(n14660), .B2(n13402), .ZN(
        n11539) );
  AOI211_X1 U14007 ( .C1(n13514), .C2(n14657), .A(n11540), .B(n11539), .ZN(
        n11541) );
  OAI21_X1 U14008 ( .B1(n11542), .B2(n14652), .A(n11541), .ZN(P2_U3198) );
  OR2_X1 U14009 ( .A1(n12897), .A2(n14420), .ZN(n11544) );
  INV_X1 U14010 ( .A(n13061), .ZN(n11545) );
  XNOR2_X1 U14011 ( .A(n13514), .B(n11545), .ZN(n13403) );
  INV_X1 U14012 ( .A(n13403), .ZN(n13413) );
  OR2_X1 U14013 ( .A1(n13514), .A2(n11545), .ZN(n11546) );
  NAND2_X1 U14014 ( .A1(n11547), .A2(n12963), .ZN(n11549) );
  AOI22_X1 U14015 ( .A1(n11862), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n11861), 
        .B2(n14769), .ZN(n11548) );
  XNOR2_X1 U14016 ( .A(n13509), .B(n13408), .ZN(n13028) );
  XNOR2_X1 U14017 ( .A(n13177), .B(n11560), .ZN(n11556) );
  OR2_X1 U14018 ( .A1(n11550), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U14019 ( .A1(n11874), .A2(n11551), .ZN(n13387) );
  AOI22_X1 U14020 ( .A1(n12941), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n12959), 
        .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n11553) );
  NAND2_X1 U14021 ( .A1(n12958), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n11552) );
  OAI211_X1 U14022 ( .C1(n13387), .C2(n11887), .A(n11553), .B(n11552), .ZN(
        n13155) );
  AND2_X1 U14023 ( .A1(n13061), .A2(n13405), .ZN(n11554) );
  AOI21_X1 U14024 ( .B1(n13155), .B2(n13407), .A(n11554), .ZN(n12746) );
  INV_X1 U14025 ( .A(n12746), .ZN(n11555) );
  AOI21_X1 U14026 ( .B1(n11556), .B2(n14798), .A(n11555), .ZN(n13511) );
  OR2_X1 U14027 ( .A1(n12897), .A2(n13406), .ZN(n11559) );
  NAND2_X1 U14028 ( .A1(n11561), .A2(n11560), .ZN(n13154) );
  OAI21_X1 U14029 ( .B1(n11561), .B2(n11560), .A(n13154), .ZN(n13512) );
  OAI22_X1 U14030 ( .A1(n14809), .A2(n11174), .B1(n12744), .B2(n14803), .ZN(
        n11562) );
  AOI21_X1 U14031 ( .B1(n13509), .B2(n14785), .A(n11562), .ZN(n11565) );
  INV_X1 U14032 ( .A(n13509), .ZN(n12751) );
  OR2_X1 U14033 ( .A1(n13400), .A2(n12751), .ZN(n11563) );
  AND3_X1 U14034 ( .A1(n13386), .A2(n10803), .A3(n11563), .ZN(n13508) );
  NAND2_X1 U14035 ( .A1(n13508), .A2(n13425), .ZN(n11564) );
  OAI211_X1 U14036 ( .C1(n13512), .C2(n13396), .A(n11565), .B(n11564), .ZN(
        n11566) );
  INV_X1 U14037 ( .A(n11566), .ZN(n11567) );
  OAI21_X1 U14038 ( .B1(n14811), .B2(n13511), .A(n11567), .ZN(P2_U3248) );
  INV_X1 U14039 ( .A(n11987), .ZN(n13575) );
  OAI222_X1 U14040 ( .A1(n13873), .A2(P1_U3086), .B1(n14305), .B2(n13575), 
        .C1(n11568), .C2(n14302), .ZN(P1_U3327) );
  INV_X1 U14041 ( .A(n12964), .ZN(n13567) );
  OAI222_X1 U14042 ( .A1(n14305), .A2(n13567), .B1(n11569), .B2(P1_U3086), 
        .C1(n11771), .C2(n14302), .ZN(P1_U3325) );
  INV_X1 U14043 ( .A(n11570), .ZN(n11574) );
  AOI22_X1 U14044 ( .A1(n14352), .A2(n14952), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n14957), .ZN(n11571) );
  OAI21_X1 U14045 ( .B1(n11572), .B2(n14354), .A(n11571), .ZN(n11573) );
  AOI21_X1 U14046 ( .B1(n11574), .B2(n14380), .A(n11573), .ZN(n11575) );
  OAI21_X1 U14047 ( .B1(n11576), .B2(n14957), .A(n11575), .ZN(P3_U3204) );
  INV_X1 U14048 ( .A(n13840), .ZN(n13582) );
  NAND2_X1 U14049 ( .A1(n11599), .A2(n14135), .ZN(n11580) );
  NAND2_X1 U14050 ( .A1(n14127), .A2(n14126), .ZN(n14125) );
  NAND2_X1 U14051 ( .A1(n14088), .A2(n14087), .ZN(n14086) );
  OAI21_X1 U14052 ( .B1(n14228), .B2(n14105), .A(n14086), .ZN(n14081) );
  INV_X1 U14053 ( .A(n14068), .ZN(n14082) );
  INV_X1 U14054 ( .A(n14022), .ZN(n14020) );
  INV_X1 U14055 ( .A(n11596), .ZN(n11582) );
  NAND2_X1 U14056 ( .A1(n11583), .A2(n11582), .ZN(n13996) );
  OAI21_X1 U14057 ( .B1(n11583), .B2(n11582), .A(n13996), .ZN(n14187) );
  INV_X1 U14058 ( .A(n13839), .ZN(n11597) );
  INV_X1 U14059 ( .A(n13842), .ZN(n13773) );
  INV_X1 U14060 ( .A(n11587), .ZN(n11588) );
  INV_X1 U14061 ( .A(n14126), .ZN(n14118) );
  INV_X1 U14062 ( .A(n14236), .ZN(n14100) );
  AOI22_X1 U14063 ( .A1(n14096), .A2(n14097), .B1(n14100), .B2(n13844), .ZN(
        n14085) );
  INV_X1 U14064 ( .A(n14087), .ZN(n11591) );
  INV_X1 U14065 ( .A(n14105), .ZN(n13718) );
  AOI21_X1 U14066 ( .B1(n14085), .B2(n11591), .A(n11590), .ZN(n14069) );
  INV_X1 U14067 ( .A(n13843), .ZN(n11592) );
  INV_X1 U14068 ( .A(n14047), .ZN(n14036) );
  NOR2_X1 U14069 ( .A1(n14201), .A2(n13772), .ZN(n11595) );
  NAND2_X1 U14070 ( .A1(n14188), .A2(n14076), .ZN(n11604) );
  OAI22_X1 U14071 ( .A1(n14076), .A2(n11598), .B1(n13748), .B2(n14106), .ZN(
        n11602) );
  NAND2_X1 U14072 ( .A1(n14101), .A2(n14100), .ZN(n14099) );
  OAI21_X1 U14073 ( .B1(n14011), .B2(n14189), .A(n13984), .ZN(n14190) );
  NOR2_X1 U14074 ( .A1(n14190), .A2(n14112), .ZN(n11601) );
  AOI211_X1 U14075 ( .C1(n14110), .C2(n13982), .A(n11602), .B(n11601), .ZN(
        n11603) );
  OAI211_X1 U14076 ( .C1(n14164), .C2(n14187), .A(n11604), .B(n11603), .ZN(
        P1_U3265) );
  INV_X1 U14077 ( .A(n11605), .ZN(n11607) );
  OAI222_X1 U14078 ( .A1(n12694), .A2(n11607), .B1(n12698), .B2(n11606), .C1(
        P3_U3151), .C2(n11833), .ZN(P3_U3267) );
  OAI222_X1 U14079 ( .A1(n11610), .A2(P1_U3086), .B1(n14305), .B2(n11609), 
        .C1(n11608), .C2(n14302), .ZN(P1_U3331) );
  MUX2_X1 U14080 ( .A(n11613), .B(n11612), .S(n11736), .Z(n11745) );
  INV_X1 U14081 ( .A(n12396), .ZN(n12400) );
  MUX2_X1 U14082 ( .A(n12395), .B(n11614), .S(n11736), .Z(n11743) );
  NAND2_X1 U14083 ( .A1(n11616), .A2(n11615), .ZN(n11617) );
  NAND2_X1 U14084 ( .A1(n11617), .A2(n12418), .ZN(n11618) );
  MUX2_X1 U14085 ( .A(n11618), .B(n12418), .S(n11736), .Z(n11741) );
  INV_X1 U14086 ( .A(n11619), .ZN(n11621) );
  MUX2_X1 U14087 ( .A(n11621), .B(n11620), .S(n11736), .Z(n11735) );
  NAND3_X1 U14088 ( .A1(n12112), .A2(n12458), .A3(n11736), .ZN(n11732) );
  INV_X1 U14089 ( .A(n11622), .ZN(n11624) );
  MUX2_X1 U14090 ( .A(n11626), .B(n11625), .S(n11755), .Z(n11729) );
  MUX2_X1 U14091 ( .A(n8923), .B(n11629), .S(n11755), .Z(n11635) );
  NAND2_X1 U14092 ( .A1(n11628), .A2(n11633), .ZN(n11627) );
  NAND2_X1 U14093 ( .A1(n11627), .A2(n11755), .ZN(n11631) );
  NAND3_X1 U14094 ( .A1(n11629), .A2(n11628), .A3(n11836), .ZN(n11630) );
  NAND2_X1 U14095 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  OAI211_X1 U14096 ( .C1(n11633), .C2(n14943), .A(n11632), .B(n8923), .ZN(
        n11634) );
  NAND3_X1 U14097 ( .A1(n11635), .A2(n14922), .A3(n11634), .ZN(n11644) );
  NAND2_X1 U14098 ( .A1(n11641), .A2(n11636), .ZN(n11639) );
  NAND2_X1 U14099 ( .A1(n11646), .A2(n11637), .ZN(n11638) );
  MUX2_X1 U14100 ( .A(n11639), .B(n11638), .S(n11736), .Z(n11640) );
  INV_X1 U14101 ( .A(n11640), .ZN(n11643) );
  OAI21_X1 U14102 ( .B1(n11641), .B2(n11755), .A(n14908), .ZN(n11642) );
  AOI21_X1 U14103 ( .B1(n11644), .B2(n11643), .A(n11642), .ZN(n11648) );
  NOR2_X1 U14104 ( .A1(n11645), .A2(n11755), .ZN(n11647) );
  OAI22_X1 U14105 ( .A1(n11648), .A2(n11647), .B1(n11736), .B2(n11646), .ZN(
        n11649) );
  OAI211_X1 U14106 ( .C1(n11736), .C2(n11650), .A(n11649), .B(n11793), .ZN(
        n11654) );
  NAND2_X1 U14107 ( .A1(n11660), .A2(n11651), .ZN(n11652) );
  NAND2_X1 U14108 ( .A1(n11652), .A2(n11736), .ZN(n11653) );
  NAND2_X1 U14109 ( .A1(n11654), .A2(n11653), .ZN(n11659) );
  NAND2_X1 U14110 ( .A1(n14910), .A2(n11655), .ZN(n11656) );
  AOI21_X1 U14111 ( .B1(n11658), .B2(n11656), .A(n11736), .ZN(n11657) );
  AOI21_X1 U14112 ( .B1(n11659), .B2(n11658), .A(n11657), .ZN(n11665) );
  OAI21_X1 U14113 ( .B1(n11736), .B2(n11660), .A(n11794), .ZN(n11664) );
  NAND2_X1 U14114 ( .A1(n12204), .A2(n14994), .ZN(n11662) );
  MUX2_X1 U14115 ( .A(n11662), .B(n11661), .S(n11736), .Z(n11663) );
  OAI211_X1 U14116 ( .C1(n11665), .C2(n11664), .A(n11789), .B(n11663), .ZN(
        n11671) );
  NOR2_X1 U14117 ( .A1(n11677), .A2(n11666), .ZN(n11795) );
  NAND2_X1 U14118 ( .A1(n12203), .A2(n11667), .ZN(n11668) );
  MUX2_X1 U14119 ( .A(n11669), .B(n11668), .S(n11736), .Z(n11670) );
  NAND3_X1 U14120 ( .A1(n11671), .A2(n11795), .A3(n11670), .ZN(n11681) );
  MUX2_X1 U14121 ( .A(n11673), .B(n11672), .S(n11755), .Z(n11678) );
  MUX2_X1 U14122 ( .A(n11675), .B(n11674), .S(n11736), .Z(n11676) );
  OAI21_X1 U14123 ( .B1(n11678), .B2(n11677), .A(n11676), .ZN(n11679) );
  NOR2_X1 U14124 ( .A1(n11679), .A2(n14376), .ZN(n11680) );
  NAND2_X1 U14125 ( .A1(n11681), .A2(n11680), .ZN(n11685) );
  NAND2_X1 U14126 ( .A1(n11691), .A2(n11682), .ZN(n11683) );
  NAND2_X1 U14127 ( .A1(n11683), .A2(n11755), .ZN(n11684) );
  NAND2_X1 U14128 ( .A1(n11685), .A2(n11684), .ZN(n11689) );
  AOI21_X1 U14129 ( .B1(n11688), .B2(n11686), .A(n11755), .ZN(n11687) );
  AOI21_X1 U14130 ( .B1(n11689), .B2(n11688), .A(n11687), .ZN(n11696) );
  INV_X1 U14131 ( .A(n11690), .ZN(n11692) );
  OAI21_X1 U14132 ( .B1(n11691), .B2(n11755), .A(n14364), .ZN(n11695) );
  MUX2_X1 U14133 ( .A(n11693), .B(n11692), .S(n11755), .Z(n11694) );
  OAI21_X1 U14134 ( .B1(n11696), .B2(n11695), .A(n11694), .ZN(n11697) );
  NAND2_X1 U14135 ( .A1(n11697), .A2(n11800), .ZN(n11701) );
  MUX2_X1 U14136 ( .A(n11699), .B(n11698), .S(n11736), .Z(n11700) );
  NAND3_X1 U14137 ( .A1(n11701), .A2(n11802), .A3(n11700), .ZN(n11706) );
  NAND2_X1 U14138 ( .A1(n11709), .A2(n11702), .ZN(n11703) );
  NAND2_X1 U14139 ( .A1(n11703), .A2(n11755), .ZN(n11705) );
  INV_X1 U14140 ( .A(n11708), .ZN(n11704) );
  AOI21_X1 U14141 ( .B1(n11706), .B2(n11705), .A(n11704), .ZN(n11711) );
  AOI21_X1 U14142 ( .B1(n11708), .B2(n11707), .A(n11755), .ZN(n11710) );
  OAI22_X1 U14143 ( .A1(n11711), .A2(n11710), .B1(n11709), .B2(n11755), .ZN(
        n11718) );
  INV_X1 U14144 ( .A(n11712), .ZN(n11717) );
  NAND2_X1 U14145 ( .A1(n11714), .A2(n11713), .ZN(n11715) );
  NAND2_X1 U14146 ( .A1(n11715), .A2(n11719), .ZN(n11716) );
  NAND3_X1 U14147 ( .A1(n11725), .A2(n11716), .A3(n11736), .ZN(n11721) );
  AOI22_X1 U14148 ( .A1(n11718), .A2(n12531), .B1(n11717), .B2(n11721), .ZN(
        n11723) );
  NAND3_X1 U14149 ( .A1(n11724), .A2(n11719), .A3(n11755), .ZN(n11720) );
  NAND2_X1 U14150 ( .A1(n11721), .A2(n11720), .ZN(n11722) );
  OAI21_X1 U14151 ( .B1(n11723), .B2(n12517), .A(n11722), .ZN(n11727) );
  MUX2_X1 U14152 ( .A(n11725), .B(n11724), .S(n11736), .Z(n11726) );
  NAND3_X1 U14153 ( .A1(n11727), .A2(n8936), .A3(n11726), .ZN(n11728) );
  NAND3_X1 U14154 ( .A1(n12472), .A2(n11729), .A3(n11728), .ZN(n11731) );
  OR3_X1 U14155 ( .A1(n12112), .A2(n12458), .A3(n11736), .ZN(n11730) );
  NAND4_X1 U14156 ( .A1(n12461), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n11734) );
  NAND3_X1 U14157 ( .A1(n11735), .A2(n11734), .A3(n11733), .ZN(n11738) );
  NAND3_X1 U14158 ( .A1(n12449), .A2(n12162), .A3(n11736), .ZN(n11737) );
  NAND2_X1 U14159 ( .A1(n11738), .A2(n11737), .ZN(n11739) );
  NAND2_X1 U14160 ( .A1(n12430), .A2(n11739), .ZN(n11740) );
  NAND3_X1 U14161 ( .A1(n12421), .A2(n11741), .A3(n11740), .ZN(n11742) );
  NAND3_X1 U14162 ( .A1(n12400), .A2(n11743), .A3(n11742), .ZN(n11744) );
  NAND2_X1 U14163 ( .A1(n11745), .A2(n11744), .ZN(n11746) );
  AND2_X1 U14164 ( .A1(n11746), .A2(n12382), .ZN(n11747) );
  NAND2_X1 U14165 ( .A1(n7038), .A2(n11747), .ZN(n11752) );
  NAND2_X1 U14166 ( .A1(n11748), .A2(n11751), .ZN(n11749) );
  AND2_X1 U14167 ( .A1(n11752), .A2(n11749), .ZN(n11757) );
  INV_X1 U14168 ( .A(n11750), .ZN(n11754) );
  OAI211_X1 U14169 ( .C1(n11754), .C2(n11753), .A(n11752), .B(n11751), .ZN(
        n11756) );
  INV_X1 U14170 ( .A(n11758), .ZN(n11823) );
  INV_X1 U14171 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14293) );
  AOI22_X1 U14172 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n11760), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n14293), .ZN(n11761) );
  XOR2_X1 U14173 ( .A(n11762), .B(n11761), .Z(n12681) );
  INV_X1 U14174 ( .A(SI_31_), .ZN(n12676) );
  NOR2_X1 U14175 ( .A1(n6529), .A2(n12676), .ZN(n11763) );
  INV_X1 U14176 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n14353) );
  NAND2_X1 U14177 ( .A1(n6532), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11766) );
  INV_X1 U14178 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n15181) );
  OR2_X1 U14179 ( .A1(n8563), .A2(n15181), .ZN(n11765) );
  OAI211_X1 U14180 ( .C1(n14353), .C2(n11767), .A(n11766), .B(n11765), .ZN(
        n11768) );
  INV_X1 U14181 ( .A(n11768), .ZN(n11769) );
  NAND2_X1 U14182 ( .A1(n11770), .A2(n11769), .ZN(n14351) );
  NAND2_X1 U14183 ( .A1(n14383), .A2(n14351), .ZN(n11784) );
  AOI22_X1 U14184 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n13566), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n11771), .ZN(n11772) );
  XNOR2_X1 U14185 ( .A(n11773), .B(n11772), .ZN(n12683) );
  NAND2_X1 U14186 ( .A1(n12683), .A2(n11774), .ZN(n11777) );
  INV_X1 U14187 ( .A(SI_30_), .ZN(n12684) );
  OR2_X1 U14188 ( .A1(n11775), .A2(n12684), .ZN(n11776) );
  NAND2_X1 U14189 ( .A1(n14387), .A2(n11782), .ZN(n11778) );
  NAND2_X1 U14190 ( .A1(n11784), .A2(n11778), .ZN(n11816) );
  INV_X1 U14191 ( .A(n11779), .ZN(n11780) );
  NOR2_X1 U14192 ( .A1(n11816), .A2(n11780), .ZN(n11821) );
  OR2_X1 U14193 ( .A1(n14387), .A2(n11782), .ZN(n11783) );
  NAND2_X1 U14194 ( .A1(n11815), .A2(n11784), .ZN(n11785) );
  AND2_X2 U14195 ( .A1(n11786), .A2(n11785), .ZN(n11832) );
  AND4_X1 U14196 ( .A1(n14922), .A2(n11788), .A3(n14908), .A4(n11787), .ZN(
        n11792) );
  INV_X1 U14197 ( .A(n9983), .ZN(n11790) );
  NAND4_X1 U14198 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(
        n11797) );
  NAND3_X1 U14199 ( .A1(n11795), .A2(n11794), .A3(n11793), .ZN(n11796) );
  NOR3_X1 U14200 ( .A1(n11797), .A2(n11796), .A3(n14376), .ZN(n11798) );
  AND4_X1 U14201 ( .A1(n11800), .A2(n11799), .A3(n14364), .A4(n11798), .ZN(
        n11801) );
  NAND3_X1 U14202 ( .A1(n12541), .A2(n11802), .A3(n11801), .ZN(n11803) );
  NOR2_X1 U14203 ( .A1(n11804), .A2(n11803), .ZN(n11805) );
  NAND2_X1 U14204 ( .A1(n11806), .A2(n11805), .ZN(n11807) );
  NOR2_X1 U14205 ( .A1(n12503), .A2(n11807), .ZN(n11808) );
  NAND3_X1 U14206 ( .A1(n12472), .A2(n8936), .A3(n11808), .ZN(n11809) );
  NOR2_X1 U14207 ( .A1(n12442), .A2(n11809), .ZN(n11810) );
  NAND4_X1 U14208 ( .A1(n12421), .A2(n12430), .A3(n12461), .A4(n11810), .ZN(
        n11811) );
  NOR2_X1 U14209 ( .A1(n12396), .A2(n11811), .ZN(n11812) );
  NAND3_X1 U14210 ( .A1(n7038), .A2(n12382), .A3(n11812), .ZN(n11813) );
  XNOR2_X1 U14211 ( .A(n11818), .B(n11817), .ZN(n11820) );
  OAI22_X1 U14212 ( .A1(n11820), .A2(n11819), .B1(n11832), .B2(n14951), .ZN(
        n11831) );
  INV_X1 U14213 ( .A(n14387), .ZN(n11822) );
  OAI21_X1 U14214 ( .B1(n11822), .B2(n14351), .A(n11821), .ZN(n11827) );
  NOR2_X1 U14215 ( .A1(n11824), .A2(n11823), .ZN(n11826) );
  OAI22_X1 U14216 ( .A1(n11827), .A2(n11826), .B1(n14383), .B2(n11825), .ZN(
        n11828) );
  XNOR2_X1 U14217 ( .A(n11828), .B(n6525), .ZN(n11830) );
  NOR3_X1 U14218 ( .A1(n11835), .A2(n11834), .A3(n11833), .ZN(n11838) );
  OAI21_X1 U14219 ( .B1(n11839), .B2(n11836), .A(P3_B_REG_SCAN_IN), .ZN(n11837) );
  OAI22_X1 U14220 ( .A1(n11840), .A2(n11839), .B1(n11838), .B2(n11837), .ZN(
        P3_U3296) );
  INV_X1 U14221 ( .A(n11841), .ZN(n11842) );
  NOR2_X1 U14222 ( .A1(n11843), .A2(n11842), .ZN(n12741) );
  NAND2_X1 U14223 ( .A1(n13408), .A2(n6520), .ZN(n11845) );
  XNOR2_X1 U14224 ( .A(n11844), .B(n11845), .ZN(n12740) );
  INV_X1 U14225 ( .A(n11844), .ZN(n11846) );
  NAND2_X1 U14226 ( .A1(n11846), .A2(n11845), .ZN(n11847) );
  NAND2_X1 U14227 ( .A1(n11848), .A2(n12963), .ZN(n11850) );
  AOI22_X1 U14228 ( .A1(n11862), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n11861), 
        .B2(n13128), .ZN(n11849) );
  XNOR2_X1 U14229 ( .A(n13504), .B(n11948), .ZN(n11852) );
  NAND2_X1 U14230 ( .A1(n13155), .A2(n6520), .ZN(n11851) );
  NOR2_X1 U14231 ( .A1(n11852), .A2(n11851), .ZN(n11853) );
  AOI21_X1 U14232 ( .B1(n11852), .B2(n11851), .A(n11853), .ZN(n12779) );
  INV_X1 U14233 ( .A(n11853), .ZN(n11854) );
  XNOR2_X1 U14234 ( .A(n11874), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n13376) );
  NAND2_X1 U14235 ( .A1(n13376), .A2(n12004), .ZN(n11859) );
  INV_X1 U14236 ( .A(n12958), .ZN(n11923) );
  INV_X1 U14237 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13500) );
  NAND2_X1 U14238 ( .A1(n12959), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n11856) );
  NAND2_X1 U14239 ( .A1(n12941), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n11855) );
  OAI211_X1 U14240 ( .C1(n11923), .C2(n13500), .A(n11856), .B(n11855), .ZN(
        n11857) );
  INV_X1 U14241 ( .A(n11857), .ZN(n11858) );
  NAND2_X1 U14242 ( .A1(n11859), .A2(n11858), .ZN(n13158) );
  NAND2_X1 U14243 ( .A1(n13158), .A2(n6520), .ZN(n11866) );
  NAND2_X1 U14244 ( .A1(n11860), .A2(n12963), .ZN(n11864) );
  AOI22_X1 U14245 ( .A1(n11862), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11861), 
        .B2(n13052), .ZN(n11863) );
  XNOR2_X1 U14246 ( .A(n13375), .B(n11976), .ZN(n11865) );
  XOR2_X1 U14247 ( .A(n11866), .B(n11865), .Z(n12716) );
  INV_X1 U14248 ( .A(n11865), .ZN(n11867) );
  NAND2_X1 U14249 ( .A1(n11867), .A2(n11866), .ZN(n12763) );
  NAND2_X1 U14250 ( .A1(n11868), .A2(n12963), .ZN(n11871) );
  OR2_X1 U14251 ( .A1(n6521), .A2(n11869), .ZN(n11870) );
  INV_X1 U14252 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n12717) );
  INV_X1 U14253 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n11872) );
  OAI21_X1 U14254 ( .B1(n11874), .B2(n12717), .A(n11872), .ZN(n11875) );
  NAND2_X1 U14255 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n11873) );
  AND2_X1 U14256 ( .A1(n11875), .A2(n11881), .ZN(n13360) );
  NAND2_X1 U14257 ( .A1(n13360), .A2(n12004), .ZN(n11880) );
  INV_X1 U14258 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n15302) );
  NAND2_X1 U14259 ( .A1(n11977), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n11877) );
  NAND2_X1 U14260 ( .A1(n12958), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n11876) );
  OAI211_X1 U14261 ( .C1(n9650), .C2(n15302), .A(n11877), .B(n11876), .ZN(
        n11878) );
  INV_X1 U14262 ( .A(n11878), .ZN(n11879) );
  NAND2_X1 U14263 ( .A1(n11880), .A2(n11879), .ZN(n13160) );
  NAND2_X1 U14264 ( .A1(n13160), .A2(n6520), .ZN(n11892) );
  XNOR2_X1 U14265 ( .A(n11891), .B(n11892), .ZN(n12762) );
  INV_X1 U14266 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12729) );
  AND2_X1 U14267 ( .A1(n11881), .A2(n12729), .ZN(n11882) );
  OR2_X1 U14268 ( .A1(n11882), .A2(n11902), .ZN(n12728) );
  INV_X1 U14269 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n15295) );
  NAND2_X1 U14270 ( .A1(n12941), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n11884) );
  NAND2_X1 U14271 ( .A1(n12959), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n11883) );
  OAI211_X1 U14272 ( .C1(n15295), .C2(n11923), .A(n11884), .B(n11883), .ZN(
        n11885) );
  INV_X1 U14273 ( .A(n11885), .ZN(n11886) );
  OAI21_X1 U14274 ( .B1(n12728), .B2(n11887), .A(n11886), .ZN(n13162) );
  NAND2_X1 U14275 ( .A1(n13162), .A2(n6520), .ZN(n11895) );
  NAND2_X1 U14276 ( .A1(n11888), .A2(n12963), .ZN(n11890) );
  OR2_X1 U14277 ( .A1(n6521), .A2(n15216), .ZN(n11889) );
  XNOR2_X1 U14278 ( .A(n13488), .B(n11976), .ZN(n11897) );
  XOR2_X1 U14279 ( .A(n11895), .B(n11897), .Z(n12724) );
  INV_X1 U14280 ( .A(n12724), .ZN(n11894) );
  INV_X1 U14281 ( .A(n11891), .ZN(n11893) );
  NAND2_X1 U14282 ( .A1(n11893), .A2(n11892), .ZN(n12723) );
  INV_X1 U14283 ( .A(n11895), .ZN(n11896) );
  NAND2_X1 U14284 ( .A1(n11897), .A2(n11896), .ZN(n11898) );
  NAND2_X1 U14285 ( .A1(n11899), .A2(n12963), .ZN(n11901) );
  OR2_X1 U14286 ( .A1(n6521), .A2(n15205), .ZN(n11900) );
  XNOR2_X1 U14287 ( .A(n13482), .B(n11948), .ZN(n11910) );
  XNOR2_X1 U14288 ( .A(n11912), .B(n11910), .ZN(n12772) );
  NOR2_X1 U14289 ( .A1(n11902), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n11903) );
  OR2_X1 U14290 ( .A1(n11918), .A2(n11903), .ZN(n13329) );
  INV_X1 U14291 ( .A(n13329), .ZN(n12773) );
  NAND2_X1 U14292 ( .A1(n12773), .A2(n12004), .ZN(n11909) );
  INV_X1 U14293 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n11906) );
  NAND2_X1 U14294 ( .A1(n12959), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n11905) );
  NAND2_X1 U14295 ( .A1(n12941), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n11904) );
  OAI211_X1 U14296 ( .C1(n11923), .C2(n11906), .A(n11905), .B(n11904), .ZN(
        n11907) );
  INV_X1 U14297 ( .A(n11907), .ZN(n11908) );
  NOR2_X1 U14298 ( .A1(n13310), .A2(n10803), .ZN(n12771) );
  INV_X1 U14299 ( .A(n11910), .ZN(n11911) );
  NAND2_X1 U14300 ( .A1(n11912), .A2(n11911), .ZN(n11913) );
  NAND2_X1 U14301 ( .A1(n11914), .A2(n12963), .ZN(n11917) );
  OR2_X1 U14302 ( .A1(n6521), .A2(n11915), .ZN(n11916) );
  XNOR2_X1 U14303 ( .A(n13476), .B(n11948), .ZN(n11928) );
  OR2_X1 U14304 ( .A1(n11918), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n11919) );
  NAND2_X1 U14305 ( .A1(n11918), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n11935) );
  AND2_X1 U14306 ( .A1(n11919), .A2(n11935), .ZN(n13304) );
  NAND2_X1 U14307 ( .A1(n13304), .A2(n12004), .ZN(n11926) );
  INV_X1 U14308 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n11922) );
  NAND2_X1 U14309 ( .A1(n12959), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n11921) );
  NAND2_X1 U14310 ( .A1(n12941), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n11920) );
  OAI211_X1 U14311 ( .C1(n11923), .C2(n11922), .A(n11921), .B(n11920), .ZN(
        n11924) );
  INV_X1 U14312 ( .A(n11924), .ZN(n11925) );
  NAND2_X1 U14313 ( .A1(n11926), .A2(n11925), .ZN(n13286) );
  NAND2_X1 U14314 ( .A1(n13286), .A2(n9459), .ZN(n12707) );
  NAND2_X1 U14315 ( .A1(n11930), .A2(n12963), .ZN(n11933) );
  OR2_X1 U14316 ( .A1(n6521), .A2(n11931), .ZN(n11932) );
  XNOR2_X1 U14317 ( .A(n13470), .B(n11976), .ZN(n11943) );
  NAND2_X1 U14318 ( .A1(n12941), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U14319 ( .A1(n12958), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n11940) );
  INV_X1 U14320 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n11934) );
  NAND2_X1 U14321 ( .A1(n11934), .A2(n11935), .ZN(n11937) );
  INV_X1 U14322 ( .A(n11935), .ZN(n11936) );
  NAND2_X1 U14323 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n11936), .ZN(n11950) );
  AND2_X1 U14324 ( .A1(n11937), .A2(n11950), .ZN(n13292) );
  NAND2_X1 U14325 ( .A1(n12004), .A2(n13292), .ZN(n11939) );
  NAND2_X1 U14326 ( .A1(n12959), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n11938) );
  NAND4_X1 U14327 ( .A1(n11941), .A2(n11940), .A3(n11939), .A4(n11938), .ZN(
        n13311) );
  AND2_X1 U14328 ( .A1(n13311), .A2(n6520), .ZN(n11942) );
  NAND2_X1 U14329 ( .A1(n11943), .A2(n11942), .ZN(n11944) );
  OAI21_X1 U14330 ( .B1(n11943), .B2(n11942), .A(n11944), .ZN(n12753) );
  NAND2_X1 U14331 ( .A1(n12754), .A2(n11944), .ZN(n12733) );
  NAND2_X1 U14332 ( .A1(n11945), .A2(n12963), .ZN(n11947) );
  OR2_X1 U14333 ( .A1(n6521), .A2(n15291), .ZN(n11946) );
  XNOR2_X1 U14334 ( .A(n13276), .B(n11948), .ZN(n11957) );
  NAND2_X1 U14335 ( .A1(n12958), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U14336 ( .A1(n12941), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n11954) );
  INV_X1 U14337 ( .A(n11950), .ZN(n11949) );
  NAND2_X1 U14338 ( .A1(n11949), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n11961) );
  INV_X1 U14339 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n15141) );
  NAND2_X1 U14340 ( .A1(n15141), .A2(n11950), .ZN(n11951) );
  AND2_X1 U14341 ( .A1(n11961), .A2(n11951), .ZN(n13277) );
  NAND2_X1 U14342 ( .A1(n12004), .A2(n13277), .ZN(n11953) );
  NAND2_X1 U14343 ( .A1(n12959), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n11952) );
  NAND4_X1 U14344 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n13287) );
  NAND2_X1 U14345 ( .A1(n13287), .A2(n9459), .ZN(n11956) );
  NOR2_X1 U14346 ( .A1(n11957), .A2(n11956), .ZN(n11958) );
  AOI21_X1 U14347 ( .B1(n11957), .B2(n11956), .A(n11958), .ZN(n12735) );
  INV_X1 U14348 ( .A(n11958), .ZN(n11959) );
  NAND2_X1 U14349 ( .A1(n12958), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n11966) );
  NAND2_X1 U14350 ( .A1(n12941), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n11965) );
  INV_X1 U14351 ( .A(n11961), .ZN(n11960) );
  NAND2_X1 U14352 ( .A1(n11960), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n11994) );
  INV_X1 U14353 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n15231) );
  NAND2_X1 U14354 ( .A1(n11961), .A2(n15231), .ZN(n11962) );
  AND2_X1 U14355 ( .A1(n11994), .A2(n11962), .ZN(n12790) );
  NAND2_X1 U14356 ( .A1(n12004), .A2(n12790), .ZN(n11964) );
  NAND2_X1 U14357 ( .A1(n12959), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n11963) );
  NAND4_X1 U14358 ( .A1(n11966), .A2(n11965), .A3(n11964), .A4(n11963), .ZN(
        n13238) );
  NAND2_X1 U14359 ( .A1(n13238), .A2(n9459), .ZN(n11970) );
  NAND2_X1 U14360 ( .A1(n11967), .A2(n12963), .ZN(n11969) );
  OR2_X1 U14361 ( .A1(n6521), .A2(n15117), .ZN(n11968) );
  XOR2_X1 U14362 ( .A(n11970), .B(n11972), .Z(n12789) );
  INV_X1 U14363 ( .A(n11970), .ZN(n11971) );
  NAND2_X1 U14364 ( .A1(n13576), .A2(n12963), .ZN(n11975) );
  OR2_X1 U14365 ( .A1(n6521), .A2(n13579), .ZN(n11974) );
  XNOR2_X1 U14366 ( .A(n13454), .B(n11976), .ZN(n11983) );
  NAND2_X1 U14367 ( .A1(n12958), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n11981) );
  NAND2_X1 U14368 ( .A1(n11977), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n11980) );
  XNOR2_X1 U14369 ( .A(n11994), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13243) );
  NAND2_X1 U14370 ( .A1(n12004), .A2(n13243), .ZN(n11979) );
  NAND2_X1 U14371 ( .A1(n12959), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n11978) );
  NAND4_X1 U14372 ( .A1(n11981), .A2(n11980), .A3(n11979), .A4(n11978), .ZN(
        n13252) );
  AND2_X1 U14373 ( .A1(n13252), .A2(n9459), .ZN(n11982) );
  NAND2_X1 U14374 ( .A1(n11983), .A2(n11982), .ZN(n11986) );
  OAI21_X1 U14375 ( .B1(n11983), .B2(n11982), .A(n11986), .ZN(n12700) );
  NAND2_X1 U14376 ( .A1(n11987), .A2(n12963), .ZN(n11990) );
  OR2_X1 U14377 ( .A1(n6521), .A2(n11988), .ZN(n11989) );
  NAND2_X1 U14378 ( .A1(n12941), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n11999) );
  NAND2_X1 U14379 ( .A1(n12959), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n11998) );
  INV_X1 U14380 ( .A(n11994), .ZN(n11992) );
  AND2_X1 U14381 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n11991) );
  NAND2_X1 U14382 ( .A1(n11992), .A2(n11991), .ZN(n12003) );
  INV_X1 U14383 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12701) );
  INV_X1 U14384 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n11993) );
  OAI21_X1 U14385 ( .B1(n11994), .B2(n12701), .A(n11993), .ZN(n11995) );
  AND2_X1 U14386 ( .A1(n12003), .A2(n11995), .ZN(n12002) );
  NAND2_X1 U14387 ( .A1(n12004), .A2(n12002), .ZN(n11997) );
  NAND2_X1 U14388 ( .A1(n12958), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n11996) );
  NAND4_X1 U14389 ( .A1(n11999), .A2(n11998), .A3(n11997), .A4(n11996), .ZN(
        n13237) );
  NAND2_X1 U14390 ( .A1(n13237), .A2(n6520), .ZN(n12000) );
  INV_X1 U14391 ( .A(n12002), .ZN(n13225) );
  NAND2_X1 U14392 ( .A1(n12958), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n12008) );
  NAND2_X1 U14393 ( .A1(n11977), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n12007) );
  INV_X1 U14394 ( .A(n12003), .ZN(n13210) );
  NAND2_X1 U14395 ( .A1(n12004), .A2(n13210), .ZN(n12006) );
  NAND2_X1 U14396 ( .A1(n12959), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n12005) );
  NAND4_X1 U14397 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(
        n13060) );
  NAND2_X1 U14398 ( .A1(n13060), .A2(n13407), .ZN(n12010) );
  NAND2_X1 U14399 ( .A1(n13252), .A2(n13405), .ZN(n12009) );
  NAND2_X1 U14400 ( .A1(n12010), .A2(n12009), .ZN(n13219) );
  AOI22_X1 U14401 ( .A1(n12783), .A2(n13219), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12011) );
  OAI21_X1 U14402 ( .B1(n13225), .B2(n14660), .A(n12011), .ZN(n12012) );
  AOI21_X1 U14403 ( .B1(n13228), .B2(n14657), .A(n12012), .ZN(n12013) );
  XNOR2_X1 U14404 ( .A(n12014), .B(n12046), .ZN(n12015) );
  INV_X1 U14405 ( .A(n12193), .ZN(n12403) );
  NOR2_X1 U14406 ( .A1(n12015), .A2(n12403), .ZN(n12092) );
  AOI21_X1 U14407 ( .B1(n12015), .B2(n12403), .A(n12092), .ZN(n12052) );
  XNOR2_X1 U14408 ( .A(n12639), .B(n12046), .ZN(n12039) );
  INV_X1 U14409 ( .A(n12039), .ZN(n12061) );
  XNOR2_X1 U14410 ( .A(n12635), .B(n12046), .ZN(n12016) );
  NAND2_X1 U14411 ( .A1(n12016), .A2(n12066), .ZN(n12040) );
  OAI21_X1 U14412 ( .B1(n12016), .B2(n12066), .A(n12040), .ZN(n12139) );
  NAND2_X1 U14413 ( .A1(n12017), .A2(n14332), .ZN(n12018) );
  XNOR2_X1 U14414 ( .A(n12659), .B(n12095), .ZN(n12021) );
  XNOR2_X1 U14415 ( .A(n12021), .B(n12538), .ZN(n12126) );
  NAND2_X1 U14416 ( .A1(n12021), .A2(n12020), .ZN(n12022) );
  XNOR2_X1 U14417 ( .A(n12511), .B(n12095), .ZN(n12166) );
  AND2_X1 U14418 ( .A1(n12166), .A2(n12494), .ZN(n12023) );
  XNOR2_X1 U14419 ( .A(n12655), .B(n12095), .ZN(n12024) );
  XNOR2_X1 U14420 ( .A(n12024), .B(n12169), .ZN(n12083) );
  NAND2_X1 U14421 ( .A1(n12084), .A2(n12083), .ZN(n12026) );
  NAND2_X1 U14422 ( .A1(n12024), .A2(n12509), .ZN(n12025) );
  NAND2_X1 U14423 ( .A1(n12026), .A2(n12025), .ZN(n12151) );
  XNOR2_X1 U14424 ( .A(n12650), .B(n12095), .ZN(n12027) );
  XNOR2_X1 U14425 ( .A(n12027), .B(n12200), .ZN(n12150) );
  NAND2_X1 U14426 ( .A1(n12151), .A2(n12150), .ZN(n12030) );
  INV_X1 U14427 ( .A(n12027), .ZN(n12028) );
  NAND2_X1 U14428 ( .A1(n12028), .A2(n12200), .ZN(n12029) );
  XNOR2_X1 U14429 ( .A(n12112), .B(n12095), .ZN(n12031) );
  NAND2_X1 U14430 ( .A1(n12031), .A2(n12458), .ZN(n12034) );
  INV_X1 U14431 ( .A(n12031), .ZN(n12032) );
  NAND2_X1 U14432 ( .A1(n12032), .A2(n12480), .ZN(n12033) );
  NAND2_X1 U14433 ( .A1(n12034), .A2(n12033), .ZN(n12108) );
  XNOR2_X1 U14434 ( .A(n12642), .B(n12095), .ZN(n12035) );
  NAND2_X1 U14435 ( .A1(n12036), .A2(n12035), .ZN(n12038) );
  NAND2_X1 U14436 ( .A1(n12038), .A2(n12037), .ZN(n12159) );
  INV_X1 U14437 ( .A(n12040), .ZN(n12118) );
  XNOR2_X1 U14438 ( .A(n12041), .B(n12095), .ZN(n12042) );
  NAND2_X1 U14439 ( .A1(n12042), .A2(n12145), .ZN(n12045) );
  INV_X1 U14440 ( .A(n12042), .ZN(n12043) );
  INV_X1 U14441 ( .A(n12145), .ZN(n12429) );
  NAND2_X1 U14442 ( .A1(n12043), .A2(n12429), .ZN(n12044) );
  AND2_X1 U14443 ( .A1(n12045), .A2(n12044), .ZN(n12117) );
  NAND2_X1 U14444 ( .A1(n12116), .A2(n12045), .ZN(n12187) );
  XNOR2_X1 U14445 ( .A(n12047), .B(n6517), .ZN(n12048) );
  NOR2_X1 U14446 ( .A1(n12048), .A2(n12415), .ZN(n12049) );
  AOI21_X1 U14447 ( .B1(n12048), .B2(n12415), .A(n12049), .ZN(n12188) );
  NAND2_X1 U14448 ( .A1(n12187), .A2(n12188), .ZN(n12186) );
  INV_X1 U14449 ( .A(n12049), .ZN(n12050) );
  NAND2_X1 U14450 ( .A1(n12186), .A2(n12050), .ZN(n12051) );
  NAND2_X1 U14451 ( .A1(n12051), .A2(n12052), .ZN(n12094) );
  OAI21_X1 U14452 ( .B1(n12052), .B2(n12051), .A(n12094), .ZN(n12053) );
  NAND2_X1 U14453 ( .A1(n12053), .A2(n14343), .ZN(n12059) );
  NAND2_X1 U14454 ( .A1(n12415), .A2(n12190), .ZN(n12054) );
  OAI21_X1 U14455 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n12055), .A(n12054), .ZN(
        n12057) );
  NOR2_X1 U14456 ( .A1(n12387), .A2(n12192), .ZN(n12056) );
  AOI211_X1 U14457 ( .C1(n12390), .C2(n12195), .A(n12057), .B(n12056), .ZN(
        n12058) );
  OAI211_X1 U14458 ( .C1(n12624), .C2(n12198), .A(n12059), .B(n12058), .ZN(
        P3_U3154) );
  INV_X1 U14459 ( .A(n12060), .ZN(n12062) );
  NOR2_X1 U14460 ( .A1(n12062), .A2(n12061), .ZN(n12137) );
  AOI21_X1 U14461 ( .B1(n12062), .B2(n12061), .A(n12137), .ZN(n12063) );
  NAND2_X1 U14462 ( .A1(n12063), .A2(n12162), .ZN(n12140) );
  OAI21_X1 U14463 ( .B1(n12162), .B2(n12063), .A(n12140), .ZN(n12064) );
  NAND2_X1 U14464 ( .A1(n12064), .A2(n14343), .ZN(n12069) );
  AOI22_X1 U14465 ( .A1(n12444), .A2(n12190), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12065) );
  OAI21_X1 U14466 ( .B1(n12066), .B2(n12192), .A(n12065), .ZN(n12067) );
  AOI21_X1 U14467 ( .B1(n12448), .B2(n12195), .A(n12067), .ZN(n12068) );
  OAI211_X1 U14468 ( .C1(n12639), .C2(n12198), .A(n12069), .B(n12068), .ZN(
        P3_U3156) );
  AND2_X1 U14469 ( .A1(n12071), .A2(n12070), .ZN(n12074) );
  OAI211_X1 U14470 ( .C1(n12074), .C2(n12073), .A(n14343), .B(n12072), .ZN(
        n12082) );
  AOI21_X1 U14471 ( .B1(n14333), .B2(n12076), .A(n12075), .ZN(n12081) );
  AOI22_X1 U14472 ( .A1(n12190), .A2(n12202), .B1(n14341), .B2(n12077), .ZN(
        n12080) );
  OR2_X1 U14473 ( .A1(n14347), .A2(n12078), .ZN(n12079) );
  NAND4_X1 U14474 ( .A1(n12082), .A2(n12081), .A3(n12080), .A4(n12079), .ZN(
        P3_U3157) );
  XOR2_X1 U14475 ( .A(n12084), .B(n12083), .Z(n12085) );
  NAND2_X1 U14476 ( .A1(n12085), .A2(n14343), .ZN(n12091) );
  INV_X1 U14477 ( .A(n12086), .ZN(n12499) );
  NOR2_X1 U14478 ( .A1(n14347), .A2(n12499), .ZN(n12089) );
  NAND2_X1 U14479 ( .A1(n12525), .A2(n12190), .ZN(n12087) );
  NAND2_X1 U14480 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12353)
         );
  OAI211_X1 U14481 ( .C1(n12495), .C2(n12192), .A(n12087), .B(n12353), .ZN(
        n12088) );
  NOR2_X1 U14482 ( .A1(n12089), .A2(n12088), .ZN(n12090) );
  OAI211_X1 U14483 ( .C1(n12198), .C2(n12655), .A(n12091), .B(n12090), .ZN(
        P3_U3159) );
  INV_X1 U14484 ( .A(n12092), .ZN(n12093) );
  NAND2_X1 U14485 ( .A1(n12094), .A2(n12093), .ZN(n12097) );
  XNOR2_X1 U14486 ( .A(n12373), .B(n12095), .ZN(n12096) );
  XNOR2_X1 U14487 ( .A(n12097), .B(n12096), .ZN(n12104) );
  OAI22_X1 U14488 ( .A1(n12193), .A2(n14336), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12098), .ZN(n12101) );
  INV_X1 U14489 ( .A(n12375), .ZN(n12099) );
  OAI22_X1 U14490 ( .A1(n12370), .A2(n12192), .B1(n12099), .B2(n14347), .ZN(
        n12100) );
  AOI211_X1 U14491 ( .C1(n12102), .C2(n14341), .A(n12101), .B(n12100), .ZN(
        n12103) );
  OAI21_X1 U14492 ( .B1(n12104), .B2(n12174), .A(n12103), .ZN(P3_U3160) );
  INV_X1 U14493 ( .A(n12105), .ZN(n12106) );
  AOI21_X1 U14494 ( .B1(n12108), .B2(n12107), .A(n12106), .ZN(n12115) );
  OAI22_X1 U14495 ( .A1(n12495), .A2(n14336), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12109), .ZN(n12111) );
  NOR2_X1 U14496 ( .A1(n12470), .A2(n12192), .ZN(n12110) );
  AOI211_X1 U14497 ( .C1(n12473), .C2(n12195), .A(n12111), .B(n12110), .ZN(
        n12114) );
  NAND2_X1 U14498 ( .A1(n12112), .A2(n14341), .ZN(n12113) );
  OAI211_X1 U14499 ( .C1(n12115), .C2(n12174), .A(n12114), .B(n12113), .ZN(
        P3_U3163) );
  INV_X1 U14500 ( .A(n12116), .ZN(n12120) );
  NOR3_X1 U14501 ( .A1(n12141), .A2(n12118), .A3(n12117), .ZN(n12119) );
  OAI21_X1 U14502 ( .B1(n12120), .B2(n12119), .A(n14343), .ZN(n12124) );
  AOI22_X1 U14503 ( .A1(n12445), .A2(n12190), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12121) );
  OAI21_X1 U14504 ( .B1(n12386), .B2(n12192), .A(n12121), .ZN(n12122) );
  AOI21_X1 U14505 ( .B1(n12423), .B2(n12195), .A(n12122), .ZN(n12123) );
  OAI211_X1 U14506 ( .C1(n12631), .C2(n12198), .A(n12124), .B(n12123), .ZN(
        P3_U3165) );
  INV_X1 U14507 ( .A(n12659), .ZN(n12136) );
  OAI21_X1 U14508 ( .B1(n12127), .B2(n12126), .A(n12125), .ZN(n12128) );
  NAND2_X1 U14509 ( .A1(n12128), .A2(n14343), .ZN(n12135) );
  NOR2_X1 U14510 ( .A1(n12129), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12296) );
  AOI21_X1 U14511 ( .B1(n12525), .B2(n14333), .A(n12296), .ZN(n12130) );
  OAI21_X1 U14512 ( .B1(n12131), .B2(n14336), .A(n12130), .ZN(n12132) );
  AOI21_X1 U14513 ( .B1(n12133), .B2(n12195), .A(n12132), .ZN(n12134) );
  OAI211_X1 U14514 ( .C1(n12136), .C2(n12198), .A(n12135), .B(n12134), .ZN(
        P3_U3168) );
  INV_X1 U14515 ( .A(n12137), .ZN(n12138) );
  AND3_X1 U14516 ( .A1(n12140), .A2(n12139), .A3(n12138), .ZN(n12142) );
  OAI21_X1 U14517 ( .B1(n12142), .B2(n12141), .A(n14343), .ZN(n12149) );
  INV_X1 U14518 ( .A(n12435), .ZN(n12143) );
  NOR2_X1 U14519 ( .A1(n12143), .A2(n14347), .ZN(n12147) );
  INV_X1 U14520 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12144) );
  OAI22_X1 U14521 ( .A1(n12145), .A2(n12192), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12144), .ZN(n12146) );
  AOI211_X1 U14522 ( .C1(n12190), .C2(n12456), .A(n12147), .B(n12146), .ZN(
        n12148) );
  OAI211_X1 U14523 ( .C1(n12635), .C2(n12198), .A(n12149), .B(n12148), .ZN(
        P3_U3169) );
  XNOR2_X1 U14524 ( .A(n12151), .B(n12150), .ZN(n12156) );
  NAND2_X1 U14525 ( .A1(n12195), .A2(n12487), .ZN(n12153) );
  AOI22_X1 U14526 ( .A1(n12480), .A2(n14333), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12152) );
  OAI211_X1 U14527 ( .C1(n12169), .C2(n14336), .A(n12153), .B(n12152), .ZN(
        n12154) );
  AOI21_X1 U14528 ( .B1(n12650), .B2(n14341), .A(n12154), .ZN(n12155) );
  OAI21_X1 U14529 ( .B1(n12156), .B2(n12174), .A(n12155), .ZN(P3_U3173) );
  INV_X1 U14530 ( .A(n12157), .ZN(n12158) );
  AOI21_X1 U14531 ( .B1(n12444), .B2(n12159), .A(n12158), .ZN(n12165) );
  NAND2_X1 U14532 ( .A1(n12195), .A2(n12463), .ZN(n12161) );
  AOI22_X1 U14533 ( .A1(n12480), .A2(n12190), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12160) );
  OAI211_X1 U14534 ( .C1(n12162), .C2(n12192), .A(n12161), .B(n12160), .ZN(
        n12163) );
  AOI21_X1 U14535 ( .B1(n12642), .B2(n14341), .A(n12163), .ZN(n12164) );
  OAI21_X1 U14536 ( .B1(n12165), .B2(n12174), .A(n12164), .ZN(P3_U3175) );
  XNOR2_X1 U14537 ( .A(n12166), .B(n12494), .ZN(n12167) );
  XNOR2_X1 U14538 ( .A(n12168), .B(n12167), .ZN(n12175) );
  NAND2_X1 U14539 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12320)
         );
  OAI21_X1 U14540 ( .B1(n12169), .B2(n12192), .A(n12320), .ZN(n12170) );
  AOI21_X1 U14541 ( .B1(n12190), .B2(n12538), .A(n12170), .ZN(n12171) );
  OAI21_X1 U14542 ( .B1(n12512), .B2(n14347), .A(n12171), .ZN(n12172) );
  AOI21_X1 U14543 ( .B1(n12511), .B2(n14341), .A(n12172), .ZN(n12173) );
  OAI21_X1 U14544 ( .B1(n12175), .B2(n12174), .A(n12173), .ZN(P3_U3178) );
  OAI211_X1 U14545 ( .C1(n12178), .C2(n12177), .A(n12176), .B(n14343), .ZN(
        n12185) );
  AOI21_X1 U14546 ( .B1(n14341), .B2(n12180), .A(n12179), .ZN(n12184) );
  AOI22_X1 U14547 ( .A1(n12190), .A2(n14910), .B1(n14333), .B2(n12204), .ZN(
        n12183) );
  OR2_X1 U14548 ( .A1(n14347), .A2(n12181), .ZN(n12182) );
  NAND4_X1 U14549 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        P3_U3179) );
  OAI21_X1 U14550 ( .B1(n12188), .B2(n12187), .A(n12186), .ZN(n12189) );
  NAND2_X1 U14551 ( .A1(n12189), .A2(n14343), .ZN(n12197) );
  AOI22_X1 U14552 ( .A1(n12429), .A2(n12190), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12191) );
  OAI21_X1 U14553 ( .B1(n12193), .B2(n12192), .A(n12191), .ZN(n12194) );
  AOI21_X1 U14554 ( .B1(n12407), .B2(n12195), .A(n12194), .ZN(n12196) );
  OAI211_X1 U14555 ( .C1(n12627), .C2(n12198), .A(n12197), .B(n12196), .ZN(
        P3_U3180) );
  MUX2_X1 U14556 ( .A(n14351), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12199), .Z(
        P3_U3522) );
  MUX2_X1 U14557 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12403), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14558 ( .A(n12415), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12199), .Z(
        P3_U3517) );
  MUX2_X1 U14559 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12429), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14560 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12456), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14561 ( .A(n12444), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12199), .Z(
        P3_U3513) );
  MUX2_X1 U14562 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12480), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14563 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12200), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14564 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12509), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14565 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12525), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14566 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12538), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14567 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n14332), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14568 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12537), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14569 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n14360), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14570 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12201), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14571 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n14372), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14572 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n14371), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14573 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12202), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14574 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12203), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14575 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12204), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14576 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12205), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14577 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n14910), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14578 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12206), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14579 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n14911), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14580 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n6823), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14581 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n8921), .S(P3_U3897), .Z(
        P3_U3491) );
  NOR2_X1 U14582 ( .A1(n14882), .A2(n12209), .ZN(n12210) );
  INV_X1 U14583 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14888) );
  INV_X1 U14584 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12211) );
  OR2_X1 U14585 ( .A1(n12231), .A2(n12211), .ZN(n12246) );
  NAND2_X1 U14586 ( .A1(n12231), .A2(n12211), .ZN(n12212) );
  NAND2_X1 U14587 ( .A1(n12246), .A2(n12212), .ZN(n12222) );
  AOI21_X1 U14588 ( .B1(n12213), .B2(n12222), .A(n12243), .ZN(n12242) );
  INV_X1 U14589 ( .A(n14885), .ZN(n12330) );
  INV_X1 U14590 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n12215) );
  NAND2_X1 U14591 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n12214)
         );
  OAI21_X1 U14592 ( .B1(n14883), .B2(n12215), .A(n12214), .ZN(n12230) );
  NAND2_X1 U14593 ( .A1(n12217), .A2(n12216), .ZN(n14891) );
  MUX2_X1 U14594 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12691), .Z(n12218) );
  XNOR2_X1 U14595 ( .A(n12218), .B(n14882), .ZN(n14890) );
  NAND3_X1 U14596 ( .A1(n14892), .A2(n14891), .A3(n14890), .ZN(n14889) );
  INV_X1 U14597 ( .A(n12218), .ZN(n12219) );
  NAND2_X1 U14598 ( .A1(n12219), .A2(n14882), .ZN(n12226) );
  OR2_X1 U14599 ( .A1(n12231), .A2(n12220), .ZN(n12256) );
  NAND2_X1 U14600 ( .A1(n12231), .A2(n12220), .ZN(n12221) );
  NAND2_X1 U14601 ( .A1(n12256), .A2(n12221), .ZN(n12237) );
  INV_X1 U14602 ( .A(n12237), .ZN(n12224) );
  INV_X1 U14603 ( .A(n12222), .ZN(n12223) );
  MUX2_X1 U14604 ( .A(n12224), .B(n12223), .S(n12691), .Z(n12225) );
  NAND3_X1 U14605 ( .A1(n14889), .A2(n12226), .A3(n12225), .ZN(n12248) );
  INV_X1 U14606 ( .A(n12248), .ZN(n12228) );
  AOI21_X1 U14607 ( .B1(n14889), .B2(n12226), .A(n12225), .ZN(n12227) );
  NOR3_X1 U14608 ( .A1(n12228), .A2(n12227), .A3(n14873), .ZN(n12229) );
  AOI211_X1 U14609 ( .C1(n12330), .C2(n12231), .A(n12230), .B(n12229), .ZN(
        n12241) );
  AOI21_X1 U14610 ( .B1(n12238), .B2(n12237), .A(n12254), .ZN(n12239) );
  OR2_X1 U14611 ( .A1(n12239), .A2(n14903), .ZN(n12240) );
  OAI211_X1 U14612 ( .C1(n12242), .C2(n14897), .A(n12241), .B(n12240), .ZN(
        P3_U3196) );
  AOI21_X1 U14613 ( .B1(n12610), .B2(n12244), .A(n12263), .ZN(n12261) );
  INV_X1 U14614 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12245) );
  NAND2_X1 U14615 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14334)
         );
  OAI21_X1 U14616 ( .B1(n14883), .B2(n12245), .A(n14334), .ZN(n12253) );
  MUX2_X1 U14617 ( .A(n12256), .B(n12246), .S(n12691), .Z(n12247) );
  NAND2_X1 U14618 ( .A1(n12248), .A2(n12247), .ZN(n12266) );
  XNOR2_X1 U14619 ( .A(n12266), .B(n12277), .ZN(n12250) );
  MUX2_X1 U14620 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12691), .Z(n12249) );
  NOR2_X1 U14621 ( .A1(n12250), .A2(n12249), .ZN(n12267) );
  AOI21_X1 U14622 ( .B1(n12250), .B2(n12249), .A(n12267), .ZN(n12251) );
  NOR2_X1 U14623 ( .A1(n12251), .A2(n14873), .ZN(n12252) );
  AOI211_X1 U14624 ( .C1(n12330), .C2(n12268), .A(n12253), .B(n12252), .ZN(
        n12260) );
  INV_X1 U14625 ( .A(n12254), .ZN(n12255) );
  AOI21_X1 U14626 ( .B1(n15185), .B2(n12257), .A(n12278), .ZN(n12258) );
  OR2_X1 U14627 ( .A1(n12258), .A2(n14903), .ZN(n12259) );
  OAI211_X1 U14628 ( .C1(n12261), .C2(n14897), .A(n12260), .B(n12259), .ZN(
        P3_U3197) );
  NAND2_X1 U14629 ( .A1(n12272), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12308) );
  NAND2_X1 U14630 ( .A1(n12281), .A2(n12270), .ZN(n12264) );
  NAND2_X1 U14631 ( .A1(n12308), .A2(n12264), .ZN(n12265) );
  AOI21_X1 U14632 ( .B1(n6649), .B2(n12265), .A(n6558), .ZN(n12290) );
  INV_X1 U14633 ( .A(n12266), .ZN(n12269) );
  AOI21_X1 U14634 ( .B1(n12269), .B2(n12268), .A(n12267), .ZN(n12301) );
  MUX2_X1 U14635 ( .A(n12280), .B(n12270), .S(n12691), .Z(n12271) );
  NAND2_X1 U14636 ( .A1(n12271), .A2(n12281), .ZN(n12299) );
  NAND2_X1 U14637 ( .A1(n12272), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12291) );
  MUX2_X1 U14638 ( .A(n12291), .B(n12308), .S(n12691), .Z(n12298) );
  NAND2_X1 U14639 ( .A1(n12299), .A2(n12298), .ZN(n12273) );
  XNOR2_X1 U14640 ( .A(n12301), .B(n12273), .ZN(n12288) );
  NAND2_X1 U14641 ( .A1(n12330), .A2(n12281), .ZN(n12275) );
  OAI211_X1 U14642 ( .C1(n15271), .C2(n14883), .A(n12275), .B(n12274), .ZN(
        n12287) );
  AND2_X1 U14643 ( .A1(n12277), .A2(n12276), .ZN(n12279) );
  NAND2_X1 U14644 ( .A1(n12281), .A2(n12280), .ZN(n12282) );
  NAND2_X1 U14645 ( .A1(n12291), .A2(n12282), .ZN(n12283) );
  NAND2_X1 U14646 ( .A1(n12284), .A2(n12283), .ZN(n12285) );
  AOI21_X1 U14647 ( .B1(n12292), .B2(n12285), .A(n14903), .ZN(n12286) );
  AOI211_X1 U14648 ( .C1(n14893), .C2(n12288), .A(n12287), .B(n12286), .ZN(
        n12289) );
  OAI21_X1 U14649 ( .B1(n12290), .B2(n14897), .A(n12289), .ZN(P3_U3198) );
  INV_X1 U14650 ( .A(n12293), .ZN(n12294) );
  OAI21_X1 U14651 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n12295), .A(n12318), 
        .ZN(n12306) );
  AOI21_X1 U14652 ( .B1(n14862), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12296), 
        .ZN(n12297) );
  OAI21_X1 U14653 ( .B1(n14885), .B2(n12323), .A(n12297), .ZN(n12305) );
  MUX2_X1 U14654 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12691), .Z(n12324) );
  XNOR2_X1 U14655 ( .A(n12324), .B(n12323), .ZN(n12303) );
  INV_X1 U14656 ( .A(n12298), .ZN(n12300) );
  OAI21_X1 U14657 ( .B1(n12301), .B2(n12300), .A(n12299), .ZN(n12302) );
  NOR2_X1 U14658 ( .A1(n12302), .A2(n12303), .ZN(n12322) );
  AOI211_X1 U14659 ( .C1(n12303), .C2(n12302), .A(n14873), .B(n12322), .ZN(
        n12304) );
  AOI211_X1 U14660 ( .C1(n12307), .C2(n12306), .A(n12305), .B(n12304), .ZN(
        n12315) );
  INV_X1 U14661 ( .A(n12309), .ZN(n12311) );
  NAND2_X1 U14662 ( .A1(n12312), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n12336) );
  OAI21_X1 U14663 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n12312), .A(n12336), 
        .ZN(n12313) );
  NAND2_X1 U14664 ( .A1(n12313), .A2(n12362), .ZN(n12314) );
  NAND2_X1 U14665 ( .A1(n12315), .A2(n12314), .ZN(P3_U3199) );
  OR2_X1 U14666 ( .A1(n12347), .A2(n12513), .ZN(n12341) );
  NAND2_X1 U14667 ( .A1(n12347), .A2(n12513), .ZN(n12316) );
  NAND2_X1 U14668 ( .A1(n12341), .A2(n12316), .ZN(n12317) );
  AOI21_X1 U14669 ( .B1(n12318), .B2(n6591), .A(n12317), .ZN(n12343) );
  AND3_X1 U14670 ( .A1(n12318), .A2(n6591), .A3(n12317), .ZN(n12319) );
  NOR2_X1 U14671 ( .A1(n12343), .A2(n12319), .ZN(n12340) );
  OAI21_X1 U14672 ( .B1(n14883), .B2(n12321), .A(n12320), .ZN(n12329) );
  MUX2_X1 U14673 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12691), .Z(n12326) );
  AOI21_X1 U14674 ( .B1(n12324), .B2(n12323), .A(n12322), .ZN(n12348) );
  XNOR2_X1 U14675 ( .A(n12348), .B(n12347), .ZN(n12325) );
  NOR2_X1 U14676 ( .A1(n12325), .A2(n12326), .ZN(n12346) );
  AOI21_X1 U14677 ( .B1(n12326), .B2(n12325), .A(n12346), .ZN(n12327) );
  NOR2_X1 U14678 ( .A1(n12327), .A2(n14873), .ZN(n12328) );
  AOI211_X1 U14679 ( .C1(n12330), .C2(n12347), .A(n12329), .B(n12328), .ZN(
        n12339) );
  INV_X1 U14680 ( .A(n12331), .ZN(n12335) );
  INV_X1 U14681 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12332) );
  OR2_X1 U14682 ( .A1(n12347), .A2(n12332), .ZN(n12357) );
  NAND2_X1 U14683 ( .A1(n12347), .A2(n12332), .ZN(n12333) );
  NAND2_X1 U14684 ( .A1(n12357), .A2(n12333), .ZN(n12334) );
  AND3_X1 U14685 ( .A1(n12336), .A2(n12335), .A3(n12334), .ZN(n12337) );
  OAI21_X1 U14686 ( .B1(n12359), .B2(n12337), .A(n12362), .ZN(n12338) );
  OAI211_X1 U14687 ( .C1(n12340), .C2(n14903), .A(n12339), .B(n12338), .ZN(
        P3_U3200) );
  INV_X1 U14688 ( .A(n12341), .ZN(n12342) );
  NOR2_X1 U14689 ( .A1(n12343), .A2(n12342), .ZN(n12345) );
  XNOR2_X1 U14690 ( .A(n6525), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12349) );
  INV_X1 U14691 ( .A(n12349), .ZN(n12344) );
  XNOR2_X1 U14692 ( .A(n12345), .B(n12344), .ZN(n12366) );
  AOI21_X1 U14693 ( .B1(n12348), .B2(n12347), .A(n12346), .ZN(n12351) );
  XNOR2_X1 U14694 ( .A(n6525), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12360) );
  MUX2_X1 U14695 ( .A(n12349), .B(n12360), .S(n12691), .Z(n12350) );
  XNOR2_X1 U14696 ( .A(n12351), .B(n12350), .ZN(n12356) );
  NAND2_X1 U14697 ( .A1(n14862), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12352) );
  OAI211_X1 U14698 ( .C1(n14885), .C2(n6525), .A(n12353), .B(n12352), .ZN(
        n12355) );
  AOI21_X1 U14699 ( .B1(n12356), .B2(n14893), .A(n12355), .ZN(n12365) );
  INV_X1 U14700 ( .A(n12357), .ZN(n12358) );
  NOR2_X1 U14701 ( .A1(n12359), .A2(n12358), .ZN(n12361) );
  XNOR2_X1 U14702 ( .A(n12361), .B(n12360), .ZN(n12363) );
  NAND2_X1 U14703 ( .A1(n12363), .A2(n12362), .ZN(n12364) );
  OAI211_X1 U14704 ( .C1(n12366), .C2(n14903), .A(n12365), .B(n12364), .ZN(
        P3_U3201) );
  NAND2_X1 U14705 ( .A1(n12403), .A2(n14946), .ZN(n12368) );
  OAI211_X1 U14706 ( .C1(n12370), .C2(n14930), .A(n12369), .B(n12368), .ZN(
        n12550) );
  INV_X1 U14707 ( .A(n12550), .ZN(n12379) );
  INV_X1 U14708 ( .A(n12371), .ZN(n12372) );
  NOR2_X1 U14709 ( .A1(n6589), .A2(n12372), .ZN(n12374) );
  XNOR2_X1 U14710 ( .A(n12374), .B(n12373), .ZN(n12551) );
  AOI22_X1 U14711 ( .A1(n12375), .A2(n14952), .B1(n14957), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12376) );
  OAI21_X1 U14712 ( .B1(n12620), .B2(n14354), .A(n12376), .ZN(n12377) );
  AOI21_X1 U14713 ( .B1(n12551), .B2(n14380), .A(n12377), .ZN(n12378) );
  OAI21_X1 U14714 ( .B1(n12379), .B2(n14957), .A(n12378), .ZN(P3_U3205) );
  AND2_X1 U14715 ( .A1(n12384), .A2(n12383), .ZN(n12385) );
  OAI22_X1 U14716 ( .A1(n12387), .A2(n14930), .B1(n12386), .B2(n14932), .ZN(
        n12388) );
  AOI21_X1 U14717 ( .B1(n12555), .B2(n14978), .A(n12388), .ZN(n12389) );
  INV_X1 U14718 ( .A(n12554), .ZN(n12394) );
  AOI22_X1 U14719 ( .A1(n12390), .A2(n14952), .B1(n14957), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12391) );
  OAI21_X1 U14720 ( .B1(n12624), .B2(n14354), .A(n12391), .ZN(n12392) );
  AOI21_X1 U14721 ( .B1(n12555), .B2(n14953), .A(n12392), .ZN(n12393) );
  OAI21_X1 U14722 ( .B1(n12394), .B2(n14957), .A(n12393), .ZN(P3_U3206) );
  NAND2_X1 U14723 ( .A1(n12420), .A2(n12395), .ZN(n12397) );
  NAND2_X1 U14724 ( .A1(n12397), .A2(n12396), .ZN(n12399) );
  NAND2_X1 U14725 ( .A1(n12399), .A2(n12398), .ZN(n12406) );
  XNOR2_X1 U14726 ( .A(n12401), .B(n12400), .ZN(n12402) );
  NAND2_X1 U14727 ( .A1(n12402), .A2(n14934), .ZN(n12405) );
  AOI22_X1 U14728 ( .A1(n12403), .A2(n14944), .B1(n14946), .B2(n12429), .ZN(
        n12404) );
  OAI211_X1 U14729 ( .C1(n14967), .C2(n12406), .A(n12405), .B(n12404), .ZN(
        n12557) );
  INV_X1 U14730 ( .A(n12557), .ZN(n12411) );
  INV_X1 U14731 ( .A(n12406), .ZN(n12558) );
  AOI22_X1 U14732 ( .A1(n12407), .A2(n14952), .B1(n14957), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12408) );
  OAI21_X1 U14733 ( .B1(n12627), .B2(n14354), .A(n12408), .ZN(n12409) );
  AOI21_X1 U14734 ( .B1(n12558), .B2(n14953), .A(n12409), .ZN(n12410) );
  OAI21_X1 U14735 ( .B1(n12411), .B2(n14957), .A(n12410), .ZN(P3_U3207) );
  OAI211_X1 U14736 ( .C1(n12414), .C2(n12413), .A(n12412), .B(n14934), .ZN(
        n12417) );
  AOI22_X1 U14737 ( .A1(n12415), .A2(n14944), .B1(n14946), .B2(n12445), .ZN(
        n12416) );
  NAND2_X1 U14738 ( .A1(n12417), .A2(n12416), .ZN(n12561) );
  INV_X1 U14739 ( .A(n12561), .ZN(n12427) );
  NAND2_X1 U14740 ( .A1(n12431), .A2(n12430), .ZN(n12419) );
  NAND2_X1 U14741 ( .A1(n12419), .A2(n12418), .ZN(n12422) );
  OAI21_X1 U14742 ( .B1(n12422), .B2(n12421), .A(n12420), .ZN(n12562) );
  AOI22_X1 U14743 ( .A1(n12423), .A2(n14952), .B1(n14957), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12424) );
  OAI21_X1 U14744 ( .B1(n12631), .B2(n14354), .A(n12424), .ZN(n12425) );
  AOI21_X1 U14745 ( .B1(n12562), .B2(n14380), .A(n12425), .ZN(n12426) );
  OAI21_X1 U14746 ( .B1(n12427), .B2(n14957), .A(n12426), .ZN(P3_U3208) );
  AOI21_X1 U14747 ( .B1(n12430), .B2(n12428), .A(n6863), .ZN(n12434) );
  AOI22_X1 U14748 ( .A1(n12429), .A2(n14944), .B1(n14946), .B2(n12456), .ZN(
        n12433) );
  XNOR2_X1 U14749 ( .A(n12431), .B(n12430), .ZN(n12566) );
  NAND2_X1 U14750 ( .A1(n12566), .A2(n14978), .ZN(n12432) );
  OAI211_X1 U14751 ( .C1(n12434), .C2(n14949), .A(n12433), .B(n12432), .ZN(
        n12565) );
  INV_X1 U14752 ( .A(n12565), .ZN(n12439) );
  AOI22_X1 U14753 ( .A1(n14952), .A2(n12435), .B1(n14957), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12436) );
  OAI21_X1 U14754 ( .B1(n12635), .B2(n14354), .A(n12436), .ZN(n12437) );
  AOI21_X1 U14755 ( .B1(n12566), .B2(n14953), .A(n12437), .ZN(n12438) );
  OAI21_X1 U14756 ( .B1(n12439), .B2(n14957), .A(n12438), .ZN(P3_U3209) );
  XNOR2_X1 U14757 ( .A(n12440), .B(n12442), .ZN(n12569) );
  OAI211_X1 U14758 ( .C1(n12443), .C2(n12442), .A(n12441), .B(n14934), .ZN(
        n12447) );
  AOI22_X1 U14759 ( .A1(n12445), .A2(n14944), .B1(n14946), .B2(n12444), .ZN(
        n12446) );
  AND2_X1 U14760 ( .A1(n12447), .A2(n12446), .ZN(n12571) );
  AOI22_X1 U14761 ( .A1(n14957), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12448), 
        .B2(n14952), .ZN(n12451) );
  NAND2_X1 U14762 ( .A1(n12449), .A2(n14919), .ZN(n12450) );
  OAI211_X1 U14763 ( .C1(n12571), .C2(n14957), .A(n12451), .B(n12450), .ZN(
        n12452) );
  AOI21_X1 U14764 ( .B1(n14380), .B2(n12569), .A(n12452), .ZN(n12453) );
  INV_X1 U14765 ( .A(n12453), .ZN(P3_U3210) );
  INV_X1 U14766 ( .A(n12461), .ZN(n12454) );
  XNOR2_X1 U14767 ( .A(n12455), .B(n12454), .ZN(n12460) );
  NAND2_X1 U14768 ( .A1(n12456), .A2(n14944), .ZN(n12457) );
  OAI21_X1 U14769 ( .B1(n12458), .B2(n14932), .A(n12457), .ZN(n12459) );
  AOI21_X1 U14770 ( .B1(n12460), .B2(n14934), .A(n12459), .ZN(n12576) );
  XNOR2_X1 U14771 ( .A(n12462), .B(n12461), .ZN(n12574) );
  INV_X1 U14772 ( .A(n12642), .ZN(n12465) );
  AOI22_X1 U14773 ( .A1(n14957), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n14952), 
        .B2(n12463), .ZN(n12464) );
  OAI21_X1 U14774 ( .B1(n12465), .B2(n14354), .A(n12464), .ZN(n12466) );
  AOI21_X1 U14775 ( .B1(n12574), .B2(n14380), .A(n12466), .ZN(n12467) );
  OAI21_X1 U14776 ( .B1(n12576), .B2(n14957), .A(n12467), .ZN(P3_U3211) );
  XOR2_X1 U14777 ( .A(n12472), .B(n12468), .Z(n12469) );
  OAI222_X1 U14778 ( .A1(n14930), .A2(n12470), .B1(n14932), .B2(n12495), .C1(
        n14949), .C2(n12469), .ZN(n12579) );
  INV_X1 U14779 ( .A(n12579), .ZN(n12477) );
  XOR2_X1 U14780 ( .A(n12472), .B(n12471), .Z(n12580) );
  AOI22_X1 U14781 ( .A1(n14957), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12473), 
        .B2(n14952), .ZN(n12474) );
  OAI21_X1 U14782 ( .B1(n12647), .B2(n14354), .A(n12474), .ZN(n12475) );
  AOI21_X1 U14783 ( .B1(n12580), .B2(n14380), .A(n12475), .ZN(n12476) );
  OAI21_X1 U14784 ( .B1(n12477), .B2(n14957), .A(n12476), .ZN(P3_U3212) );
  OAI211_X1 U14785 ( .C1(n12483), .C2(n12479), .A(n12478), .B(n14934), .ZN(
        n12482) );
  AOI22_X1 U14786 ( .A1(n12480), .A2(n14944), .B1(n14946), .B2(n12509), .ZN(
        n12481) );
  AND2_X1 U14787 ( .A1(n12482), .A2(n12481), .ZN(n12585) );
  NAND2_X1 U14788 ( .A1(n12484), .A2(n12483), .ZN(n12485) );
  AND2_X1 U14789 ( .A1(n12486), .A2(n12485), .ZN(n12583) );
  INV_X1 U14790 ( .A(n12650), .ZN(n12489) );
  AOI22_X1 U14791 ( .A1(n14957), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n14952), 
        .B2(n12487), .ZN(n12488) );
  OAI21_X1 U14792 ( .B1(n12489), .B2(n14354), .A(n12488), .ZN(n12490) );
  AOI21_X1 U14793 ( .B1(n12583), .B2(n14380), .A(n12490), .ZN(n12491) );
  OAI21_X1 U14794 ( .B1(n12585), .B2(n14957), .A(n12491), .ZN(P3_U3213) );
  OAI211_X1 U14795 ( .C1(n12493), .C2(n12503), .A(n12492), .B(n14934), .ZN(
        n12498) );
  OAI22_X1 U14796 ( .A1(n12495), .A2(n14930), .B1(n12494), .B2(n14932), .ZN(
        n12496) );
  INV_X1 U14797 ( .A(n12496), .ZN(n12497) );
  AND2_X1 U14798 ( .A1(n12498), .A2(n12497), .ZN(n12590) );
  INV_X1 U14799 ( .A(n12655), .ZN(n12502) );
  OAI22_X1 U14800 ( .A1(n14955), .A2(n12500), .B1(n12499), .B2(n14926), .ZN(
        n12501) );
  AOI21_X1 U14801 ( .B1(n12502), .B2(n14919), .A(n12501), .ZN(n12506) );
  XNOR2_X1 U14802 ( .A(n12504), .B(n12503), .ZN(n12588) );
  NAND2_X1 U14803 ( .A1(n12588), .A2(n14380), .ZN(n12505) );
  OAI211_X1 U14804 ( .C1(n12590), .C2(n14957), .A(n12506), .B(n12505), .ZN(
        P3_U3214) );
  OAI21_X1 U14805 ( .B1(n6656), .B2(n12517), .A(n12508), .ZN(n12510) );
  AOI222_X1 U14806 ( .A1(n14934), .A2(n12510), .B1(n12509), .B2(n14944), .C1(
        n12538), .C2(n14946), .ZN(n12596) );
  NAND2_X1 U14807 ( .A1(n12511), .A2(n14980), .ZN(n12594) );
  INV_X1 U14808 ( .A(n12594), .ZN(n12515) );
  OAI22_X1 U14809 ( .A1(n14955), .A2(n12513), .B1(n12512), .B2(n14926), .ZN(
        n12514) );
  AOI21_X1 U14810 ( .B1(n12515), .B2(n14379), .A(n12514), .ZN(n12520) );
  NAND2_X1 U14811 ( .A1(n12518), .A2(n12517), .ZN(n12593) );
  NAND3_X1 U14812 ( .A1(n12516), .A2(n12593), .A3(n14380), .ZN(n12519) );
  OAI211_X1 U14813 ( .C1(n12596), .C2(n14957), .A(n12520), .B(n12519), .ZN(
        P3_U3215) );
  NAND3_X1 U14814 ( .A1(n12521), .A2(n12531), .A3(n12522), .ZN(n12523) );
  NAND3_X1 U14815 ( .A1(n12524), .A2(n14934), .A3(n12523), .ZN(n12527) );
  AOI22_X1 U14816 ( .A1(n12525), .A2(n14944), .B1(n14946), .B2(n14332), .ZN(
        n12526) );
  OAI22_X1 U14817 ( .A1(n14955), .A2(n12529), .B1(n12528), .B2(n14926), .ZN(
        n12530) );
  AOI21_X1 U14818 ( .B1(n12659), .B2(n14919), .A(n12530), .ZN(n12534) );
  XNOR2_X1 U14819 ( .A(n12532), .B(n12531), .ZN(n12597) );
  NAND2_X1 U14820 ( .A1(n12597), .A2(n14380), .ZN(n12533) );
  OAI211_X1 U14821 ( .C1(n12599), .C2(n14957), .A(n12534), .B(n12533), .ZN(
        P3_U3216) );
  NAND2_X1 U14822 ( .A1(n12535), .A2(n12541), .ZN(n12536) );
  NAND3_X1 U14823 ( .A1(n12521), .A2(n14934), .A3(n12536), .ZN(n12540) );
  AOI22_X1 U14824 ( .A1(n12538), .A2(n14944), .B1(n14946), .B2(n12537), .ZN(
        n12539) );
  AND2_X1 U14825 ( .A1(n12540), .A2(n12539), .ZN(n12604) );
  OR2_X1 U14826 ( .A1(n12542), .A2(n12541), .ZN(n12543) );
  NAND2_X1 U14827 ( .A1(n12544), .A2(n12543), .ZN(n12602) );
  AOI22_X1 U14828 ( .A1(n14957), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n14952), 
        .B2(n12545), .ZN(n12546) );
  OAI21_X1 U14829 ( .B1(n12547), .B2(n14354), .A(n12546), .ZN(n12548) );
  AOI21_X1 U14830 ( .B1(n12602), .B2(n14380), .A(n12548), .ZN(n12549) );
  OAI21_X1 U14831 ( .B1(n12604), .B2(n14957), .A(n12549), .ZN(P3_U3217) );
  INV_X1 U14832 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12552) );
  OAI21_X1 U14833 ( .B1(n12620), .B2(n12612), .A(n12553), .ZN(P3_U3487) );
  INV_X1 U14834 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12556) );
  INV_X1 U14835 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12559) );
  AOI21_X1 U14836 ( .B1(n14992), .B2(n12558), .A(n12557), .ZN(n12625) );
  MUX2_X1 U14837 ( .A(n12559), .B(n12625), .S(n15031), .Z(n12560) );
  OAI21_X1 U14838 ( .B1(n12627), .B2(n12612), .A(n12560), .ZN(P3_U3485) );
  INV_X1 U14839 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12563) );
  AOI21_X1 U14840 ( .B1(n15011), .B2(n12562), .A(n12561), .ZN(n12628) );
  MUX2_X1 U14841 ( .A(n12563), .B(n12628), .S(n15031), .Z(n12564) );
  OAI21_X1 U14842 ( .B1(n12631), .B2(n12612), .A(n12564), .ZN(P3_U3484) );
  INV_X1 U14843 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12567) );
  AOI21_X1 U14844 ( .B1(n14992), .B2(n12566), .A(n12565), .ZN(n12632) );
  MUX2_X1 U14845 ( .A(n12567), .B(n12632), .S(n15031), .Z(n12568) );
  OAI21_X1 U14846 ( .B1(n12635), .B2(n12612), .A(n12568), .ZN(P3_U3483) );
  NAND2_X1 U14847 ( .A1(n12569), .A2(n15011), .ZN(n12570) );
  NAND2_X1 U14848 ( .A1(n12571), .A2(n12570), .ZN(n12636) );
  MUX2_X1 U14849 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12636), .S(n15031), .Z(
        n12572) );
  INV_X1 U14850 ( .A(n12572), .ZN(n12573) );
  OAI21_X1 U14851 ( .B1(n12639), .B2(n12612), .A(n12573), .ZN(P3_U3482) );
  INV_X1 U14852 ( .A(n12612), .ZN(n12606) );
  NAND2_X1 U14853 ( .A1(n12574), .A2(n15011), .ZN(n12575) );
  NAND2_X1 U14854 ( .A1(n12576), .A2(n12575), .ZN(n12640) );
  MUX2_X1 U14855 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n12640), .S(n15031), .Z(
        n12577) );
  AOI21_X1 U14856 ( .B1(n12606), .B2(n12642), .A(n12577), .ZN(n12578) );
  INV_X1 U14857 ( .A(n12578), .ZN(P3_U3481) );
  INV_X1 U14858 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12581) );
  AOI21_X1 U14859 ( .B1(n12580), .B2(n15011), .A(n12579), .ZN(n12644) );
  MUX2_X1 U14860 ( .A(n12581), .B(n12644), .S(n15031), .Z(n12582) );
  OAI21_X1 U14861 ( .B1(n12647), .B2(n12612), .A(n12582), .ZN(P3_U3480) );
  NAND2_X1 U14862 ( .A1(n12583), .A2(n15011), .ZN(n12584) );
  NAND2_X1 U14863 ( .A1(n12585), .A2(n12584), .ZN(n12648) );
  MUX2_X1 U14864 ( .A(n12648), .B(P3_REG1_REG_20__SCAN_IN), .S(n15029), .Z(
        n12586) );
  AOI21_X1 U14865 ( .B1(n12606), .B2(n12650), .A(n12586), .ZN(n12587) );
  INV_X1 U14866 ( .A(n12587), .ZN(P3_U3479) );
  NAND2_X1 U14867 ( .A1(n12588), .A2(n15011), .ZN(n12589) );
  AND2_X1 U14868 ( .A1(n12590), .A2(n12589), .ZN(n12653) );
  MUX2_X1 U14869 ( .A(n12591), .B(n12653), .S(n15031), .Z(n12592) );
  OAI21_X1 U14870 ( .B1(n12612), .B2(n12655), .A(n12592), .ZN(P3_U3478) );
  NAND3_X1 U14871 ( .A1(n12516), .A2(n12593), .A3(n15011), .ZN(n12595) );
  NAND3_X1 U14872 ( .A1(n12596), .A2(n12595), .A3(n12594), .ZN(n12656) );
  MUX2_X1 U14873 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12656), .S(n15031), .Z(
        P3_U3477) );
  NAND2_X1 U14874 ( .A1(n12597), .A2(n15011), .ZN(n12598) );
  NAND2_X1 U14875 ( .A1(n12599), .A2(n12598), .ZN(n12657) );
  MUX2_X1 U14876 ( .A(n12657), .B(P3_REG1_REG_17__SCAN_IN), .S(n15029), .Z(
        n12600) );
  AOI21_X1 U14877 ( .B1(n12606), .B2(n12659), .A(n12600), .ZN(n12601) );
  INV_X1 U14878 ( .A(n12601), .ZN(P3_U3476) );
  NAND2_X1 U14879 ( .A1(n12602), .A2(n15011), .ZN(n12603) );
  NAND2_X1 U14880 ( .A1(n12604), .A2(n12603), .ZN(n12661) );
  MUX2_X1 U14881 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12661), .S(n15031), .Z(
        n12605) );
  AOI21_X1 U14882 ( .B1(n12606), .B2(n12663), .A(n12605), .ZN(n12607) );
  INV_X1 U14883 ( .A(n12607), .ZN(P3_U3475) );
  AOI21_X1 U14884 ( .B1(n12609), .B2(n15011), .A(n12608), .ZN(n12666) );
  MUX2_X1 U14885 ( .A(n12610), .B(n12666), .S(n15031), .Z(n12611) );
  OAI21_X1 U14886 ( .B1(n12670), .B2(n12612), .A(n12611), .ZN(P3_U3474) );
  AOI21_X1 U14887 ( .B1(n14980), .B2(n12614), .A(n12613), .ZN(n12615) );
  OAI21_X1 U14888 ( .B1(n12617), .B2(n12616), .A(n12615), .ZN(n12671) );
  MUX2_X1 U14889 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n12671), .S(n15031), .Z(
        P3_U3473) );
  INV_X1 U14890 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12618) );
  OAI21_X1 U14891 ( .B1(n12620), .B2(n12669), .A(n12619), .ZN(P3_U3455) );
  INV_X1 U14892 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12622) );
  MUX2_X1 U14893 ( .A(n12622), .B(n12621), .S(n15019), .Z(n12623) );
  OAI21_X1 U14894 ( .B1(n12624), .B2(n12669), .A(n12623), .ZN(P3_U3454) );
  MUX2_X1 U14895 ( .A(n15165), .B(n12625), .S(n15019), .Z(n12626) );
  OAI21_X1 U14896 ( .B1(n12627), .B2(n12669), .A(n12626), .ZN(P3_U3453) );
  INV_X1 U14897 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12629) );
  MUX2_X1 U14898 ( .A(n12629), .B(n12628), .S(n15019), .Z(n12630) );
  OAI21_X1 U14899 ( .B1(n12631), .B2(n12669), .A(n12630), .ZN(P3_U3452) );
  INV_X1 U14900 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12633) );
  MUX2_X1 U14901 ( .A(n12633), .B(n12632), .S(n15019), .Z(n12634) );
  OAI21_X1 U14902 ( .B1(n12635), .B2(n12669), .A(n12634), .ZN(P3_U3451) );
  MUX2_X1 U14903 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n12636), .S(n15019), .Z(
        n12637) );
  INV_X1 U14904 ( .A(n12637), .ZN(n12638) );
  OAI21_X1 U14905 ( .B1(n12639), .B2(n12669), .A(n12638), .ZN(P3_U3450) );
  MUX2_X1 U14906 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n12640), .S(n15019), .Z(
        n12641) );
  AOI21_X1 U14907 ( .B1(n12664), .B2(n12642), .A(n12641), .ZN(n12643) );
  INV_X1 U14908 ( .A(n12643), .ZN(P3_U3449) );
  INV_X1 U14909 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12645) );
  MUX2_X1 U14910 ( .A(n12645), .B(n12644), .S(n15019), .Z(n12646) );
  OAI21_X1 U14911 ( .B1(n12647), .B2(n12669), .A(n12646), .ZN(P3_U3448) );
  MUX2_X1 U14912 ( .A(n12648), .B(P3_REG0_REG_20__SCAN_IN), .S(n15018), .Z(
        n12649) );
  AOI21_X1 U14913 ( .B1(n12664), .B2(n12650), .A(n12649), .ZN(n12651) );
  INV_X1 U14914 ( .A(n12651), .ZN(P3_U3447) );
  MUX2_X1 U14915 ( .A(n12653), .B(n12652), .S(n15018), .Z(n12654) );
  OAI21_X1 U14916 ( .B1(n12669), .B2(n12655), .A(n12654), .ZN(P3_U3446) );
  MUX2_X1 U14917 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n12656), .S(n15019), .Z(
        P3_U3444) );
  MUX2_X1 U14918 ( .A(n12657), .B(P3_REG0_REG_17__SCAN_IN), .S(n15018), .Z(
        n12658) );
  AOI21_X1 U14919 ( .B1(n12664), .B2(n12659), .A(n12658), .ZN(n12660) );
  INV_X1 U14920 ( .A(n12660), .ZN(P3_U3441) );
  MUX2_X1 U14921 ( .A(n12661), .B(P3_REG0_REG_16__SCAN_IN), .S(n15018), .Z(
        n12662) );
  AOI21_X1 U14922 ( .B1(n12664), .B2(n12663), .A(n12662), .ZN(n12665) );
  INV_X1 U14923 ( .A(n12665), .ZN(P3_U3438) );
  INV_X1 U14924 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12667) );
  MUX2_X1 U14925 ( .A(n12667), .B(n12666), .S(n15019), .Z(n12668) );
  OAI21_X1 U14926 ( .B1(n12670), .B2(n12669), .A(n12668), .ZN(P3_U3435) );
  MUX2_X1 U14927 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n12671), .S(n15019), .Z(
        P3_U3432) );
  MUX2_X1 U14928 ( .A(P3_D_REG_1__SCAN_IN), .B(n12672), .S(n12673), .Z(
        P3_U3377) );
  MUX2_X1 U14929 ( .A(P3_D_REG_0__SCAN_IN), .B(n12674), .S(n12673), .Z(
        P3_U3376) );
  NAND3_X1 U14930 ( .A1(n12675), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12677) );
  OAI22_X1 U14931 ( .A1(n12678), .A2(n12677), .B1(n12676), .B2(n12698), .ZN(
        n12679) );
  AOI21_X1 U14932 ( .B1(n12681), .B2(n12680), .A(n12679), .ZN(n12682) );
  INV_X1 U14933 ( .A(n12682), .ZN(P3_U3264) );
  INV_X1 U14934 ( .A(n12683), .ZN(n12685) );
  OAI222_X1 U14935 ( .A1(P3_U3151), .A2(n12686), .B1(n12694), .B2(n12685), 
        .C1(n12684), .C2(n12698), .ZN(P3_U3265) );
  INV_X1 U14936 ( .A(n12687), .ZN(n12688) );
  INV_X1 U14937 ( .A(n12690), .ZN(n12693) );
  OAI222_X1 U14938 ( .A1(n12694), .A2(n12693), .B1(n12698), .B2(n12692), .C1(
        P3_U3151), .C2(n12691), .ZN(P3_U3268) );
  INV_X1 U14939 ( .A(n12695), .ZN(n12696) );
  OAI222_X1 U14940 ( .A1(P3_U3151), .A2(n12699), .B1(n12698), .B2(n12697), 
        .C1(n12694), .C2(n12696), .ZN(P3_U3269) );
  NOR2_X1 U14941 ( .A1(n14418), .A2(n13274), .ZN(n12703) );
  INV_X1 U14942 ( .A(n13237), .ZN(n13204) );
  OAI22_X1 U14943 ( .A1(n14419), .A2(n13204), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12701), .ZN(n12702) );
  AOI211_X1 U14944 ( .C1(n12800), .C2(n13243), .A(n12703), .B(n12702), .ZN(
        n12704) );
  OAI211_X1 U14945 ( .C1(n13240), .C2(n14415), .A(n12705), .B(n12704), .ZN(
        P2_U3186) );
  XOR2_X1 U14946 ( .A(n12707), .B(n12706), .Z(n12713) );
  INV_X1 U14947 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12708) );
  OAI22_X1 U14948 ( .A1(n14419), .A2(n13273), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12708), .ZN(n12711) );
  INV_X1 U14949 ( .A(n13304), .ZN(n12709) );
  OAI22_X1 U14950 ( .A1(n13310), .A2(n14418), .B1(n12709), .B2(n14660), .ZN(
        n12710) );
  AOI211_X1 U14951 ( .C1(n13476), .C2(n14657), .A(n12711), .B(n12710), .ZN(
        n12712) );
  OAI21_X1 U14952 ( .B1(n12713), .B2(n14652), .A(n12712), .ZN(P2_U3188) );
  INV_X1 U14953 ( .A(n12765), .ZN(n12714) );
  AOI21_X1 U14954 ( .B1(n12716), .B2(n12715), .A(n12714), .ZN(n12721) );
  AOI22_X1 U14955 ( .A1(n13160), .A2(n13407), .B1(n13405), .B2(n13155), .ZN(
        n13368) );
  OAI22_X1 U14956 ( .A1(n13368), .A2(n14649), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12717), .ZN(n12718) );
  AOI21_X1 U14957 ( .B1(n13376), .B2(n12800), .A(n12718), .ZN(n12720) );
  NAND2_X1 U14958 ( .A1(n13375), .A2(n14657), .ZN(n12719) );
  OAI211_X1 U14959 ( .C1(n12721), .C2(n14652), .A(n12720), .B(n12719), .ZN(
        P2_U3191) );
  INV_X1 U14960 ( .A(n13488), .ZN(n13347) );
  NAND2_X1 U14961 ( .A1(n12722), .A2(n12723), .ZN(n12725) );
  AOI21_X1 U14962 ( .B1(n12725), .B2(n12724), .A(n14652), .ZN(n12727) );
  NAND2_X1 U14963 ( .A1(n12727), .A2(n12726), .ZN(n12732) );
  INV_X1 U14964 ( .A(n12728), .ZN(n13344) );
  INV_X1 U14965 ( .A(n13310), .ZN(n13164) );
  AOI22_X1 U14966 ( .A1(n13164), .A2(n13407), .B1(n13405), .B2(n13160), .ZN(
        n13339) );
  OAI22_X1 U14967 ( .A1(n13339), .A2(n14649), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12729), .ZN(n12730) );
  AOI21_X1 U14968 ( .B1(n13344), .B2(n12800), .A(n12730), .ZN(n12731) );
  OAI211_X1 U14969 ( .C1(n13347), .C2(n14415), .A(n12732), .B(n12731), .ZN(
        P2_U3195) );
  INV_X1 U14970 ( .A(n13276), .ZN(n13548) );
  OAI211_X1 U14971 ( .C1(n12733), .C2(n12735), .A(n12734), .B(n14644), .ZN(
        n12739) );
  NOR2_X1 U14972 ( .A1(n14418), .A2(n13273), .ZN(n12737) );
  OAI22_X1 U14973 ( .A1(n14419), .A2(n13274), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15141), .ZN(n12736) );
  AOI211_X1 U14974 ( .C1(n12800), .C2(n13277), .A(n12737), .B(n12736), .ZN(
        n12738) );
  OAI211_X1 U14975 ( .C1(n13548), .C2(n14415), .A(n12739), .B(n12738), .ZN(
        P2_U3197) );
  NOR3_X1 U14976 ( .A1(n12742), .A2(n12741), .A3(n12740), .ZN(n12743) );
  OAI21_X1 U14977 ( .B1(n6658), .B2(n12743), .A(n14644), .ZN(n12750) );
  INV_X1 U14978 ( .A(n12744), .ZN(n12748) );
  INV_X1 U14979 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12745) );
  OAI22_X1 U14980 ( .A1(n12746), .A2(n14649), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12745), .ZN(n12747) );
  AOI21_X1 U14981 ( .B1(n12748), .B2(n12800), .A(n12747), .ZN(n12749) );
  OAI211_X1 U14982 ( .C1(n12751), .C2(n14415), .A(n12750), .B(n12749), .ZN(
        P2_U3200) );
  AOI21_X1 U14983 ( .B1(n12752), .B2(n12753), .A(n14652), .ZN(n12755) );
  NAND2_X1 U14984 ( .A1(n12755), .A2(n12754), .ZN(n12759) );
  AOI22_X1 U14985 ( .A1(n12798), .A2(n13287), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12758) );
  AOI22_X1 U14986 ( .A1(n13286), .A2(n12801), .B1(n13292), .B2(n12800), .ZN(
        n12757) );
  NAND2_X1 U14987 ( .A1(n13470), .A2(n14657), .ZN(n12756) );
  NAND4_X1 U14988 ( .A1(n12759), .A2(n12758), .A3(n12757), .A4(n12756), .ZN(
        P2_U3201) );
  INV_X1 U14989 ( .A(n13360), .ZN(n12761) );
  INV_X1 U14990 ( .A(n13162), .ZN(n13319) );
  INV_X1 U14991 ( .A(n13158), .ZN(n13183) );
  OAI22_X1 U14992 ( .A1(n13319), .A2(n14799), .B1(n13183), .B2(n13318), .ZN(
        n13355) );
  AOI22_X1 U14993 ( .A1(n13355), .A2(n12783), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12760) );
  OAI21_X1 U14994 ( .B1(n12761), .B2(n14660), .A(n12760), .ZN(n12768) );
  INV_X1 U14995 ( .A(n12762), .ZN(n12764) );
  NAND3_X1 U14996 ( .A1(n12765), .A2(n12764), .A3(n12763), .ZN(n12766) );
  AOI21_X1 U14997 ( .B1(n12722), .B2(n12766), .A(n14652), .ZN(n12767) );
  AOI211_X1 U14998 ( .C1(n13493), .C2(n14657), .A(n12768), .B(n12767), .ZN(
        n12769) );
  INV_X1 U14999 ( .A(n12769), .ZN(P2_U3205) );
  OAI211_X1 U15000 ( .C1(n12772), .C2(n12771), .A(n12770), .B(n14644), .ZN(
        n12777) );
  AOI22_X1 U15001 ( .A1(n13286), .A2(n12798), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12776) );
  AOI22_X1 U15002 ( .A1(n12800), .A2(n12773), .B1(n13162), .B2(n12801), .ZN(
        n12775) );
  NAND2_X1 U15003 ( .A1(n13482), .A2(n14657), .ZN(n12774) );
  NAND4_X1 U15004 ( .A1(n12777), .A2(n12776), .A3(n12775), .A4(n12774), .ZN(
        P2_U3207) );
  INV_X1 U15005 ( .A(n13504), .ZN(n13391) );
  OAI211_X1 U15006 ( .C1(n12780), .C2(n12779), .A(n12778), .B(n14644), .ZN(
        n12785) );
  OAI22_X1 U15007 ( .A1(n13183), .A2(n14799), .B1(n12902), .B2(n13318), .ZN(
        n13383) );
  NOR2_X1 U15008 ( .A1(n14660), .A2(n13387), .ZN(n12782) );
  AOI211_X1 U15009 ( .C1(n13383), .C2(n12783), .A(n12782), .B(n12781), .ZN(
        n12784) );
  OAI211_X1 U15010 ( .C1(n13391), .C2(n14415), .A(n12785), .B(n12784), .ZN(
        P2_U3210) );
  INV_X1 U15011 ( .A(n12786), .ZN(n12787) );
  AOI21_X1 U15012 ( .B1(n12789), .B2(n12788), .A(n12787), .ZN(n12794) );
  INV_X1 U15013 ( .A(n13252), .ZN(n13198) );
  OAI22_X1 U15014 ( .A1(n14419), .A2(n13198), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15231), .ZN(n12792) );
  INV_X1 U15015 ( .A(n13287), .ZN(n13195) );
  INV_X1 U15016 ( .A(n12790), .ZN(n13256) );
  OAI22_X1 U15017 ( .A1(n14418), .A2(n13195), .B1(n14660), .B2(n13256), .ZN(
        n12791) );
  AOI211_X1 U15018 ( .C1(n13460), .C2(n14657), .A(n12792), .B(n12791), .ZN(
        n12793) );
  OAI21_X1 U15019 ( .B1(n12794), .B2(n14652), .A(n12793), .ZN(P2_U3212) );
  OAI211_X1 U15020 ( .C1(n12797), .C2(n12796), .A(n12795), .B(n14644), .ZN(
        n12805) );
  AOI22_X1 U15021 ( .A1(n12798), .A2(n13061), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12804) );
  AOI22_X1 U15022 ( .A1(n12801), .A2(n13062), .B1(n12800), .B2(n12799), .ZN(
        n12803) );
  NAND2_X1 U15023 ( .A1(n12897), .A2(n14657), .ZN(n12802) );
  NAND4_X1 U15024 ( .A1(n12805), .A2(n12804), .A3(n12803), .A4(n12802), .ZN(
        P2_U3213) );
  INV_X1 U15025 ( .A(n6571), .ZN(n12806) );
  NAND2_X1 U15026 ( .A1(n13004), .A2(n12806), .ZN(n12809) );
  NAND3_X1 U15027 ( .A1(n13005), .A2(n12809), .A3(n12886), .ZN(n12808) );
  MUX2_X1 U15028 ( .A(n13075), .B(n9381), .S(n12833), .Z(n12811) );
  MUX2_X1 U15029 ( .A(n13075), .B(n9381), .S(n12886), .Z(n12810) );
  INV_X1 U15030 ( .A(n12811), .ZN(n12812) );
  MUX2_X1 U15031 ( .A(n13074), .B(n6534), .S(n12886), .Z(n12816) );
  MUX2_X1 U15032 ( .A(n6534), .B(n13074), .S(n12886), .Z(n12814) );
  NAND2_X1 U15033 ( .A1(n12815), .A2(n12814), .ZN(n12819) );
  MUX2_X1 U15034 ( .A(n13073), .B(n12820), .S(n12886), .Z(n12821) );
  INV_X1 U15035 ( .A(n12822), .ZN(n12823) );
  MUX2_X1 U15036 ( .A(n13072), .B(n12824), .S(n12886), .Z(n12828) );
  NAND2_X1 U15037 ( .A1(n12827), .A2(n12828), .ZN(n12826) );
  MUX2_X1 U15038 ( .A(n12824), .B(n13072), .S(n12886), .Z(n12825) );
  NAND2_X1 U15039 ( .A1(n12826), .A2(n12825), .ZN(n12832) );
  INV_X1 U15040 ( .A(n12827), .ZN(n12830) );
  INV_X1 U15041 ( .A(n12828), .ZN(n12829) );
  NAND2_X1 U15042 ( .A1(n12830), .A2(n12829), .ZN(n12831) );
  NAND2_X1 U15043 ( .A1(n12832), .A2(n12831), .ZN(n12837) );
  MUX2_X1 U15044 ( .A(n12834), .B(n13071), .S(n12886), .Z(n12838) );
  NAND2_X1 U15045 ( .A1(n12837), .A2(n12838), .ZN(n12836) );
  MUX2_X1 U15046 ( .A(n12834), .B(n13071), .S(n12973), .Z(n12835) );
  NAND2_X1 U15047 ( .A1(n12836), .A2(n12835), .ZN(n12842) );
  INV_X1 U15048 ( .A(n12837), .ZN(n12840) );
  INV_X1 U15049 ( .A(n12838), .ZN(n12839) );
  NAND2_X1 U15050 ( .A1(n12840), .A2(n12839), .ZN(n12841) );
  NAND2_X1 U15051 ( .A1(n12842), .A2(n12841), .ZN(n12845) );
  MUX2_X1 U15052 ( .A(n14835), .B(n13070), .S(n12973), .Z(n12846) );
  NAND2_X1 U15053 ( .A1(n12845), .A2(n12846), .ZN(n12844) );
  MUX2_X1 U15054 ( .A(n14835), .B(n13070), .S(n12997), .Z(n12843) );
  NAND2_X1 U15055 ( .A1(n12844), .A2(n12843), .ZN(n12850) );
  INV_X1 U15056 ( .A(n12845), .ZN(n12848) );
  INV_X1 U15057 ( .A(n12846), .ZN(n12847) );
  NAND2_X1 U15058 ( .A1(n12848), .A2(n12847), .ZN(n12849) );
  NAND2_X1 U15059 ( .A1(n12850), .A2(n12849), .ZN(n12854) );
  MUX2_X1 U15060 ( .A(n13069), .B(n14786), .S(n12973), .Z(n12853) );
  NAND2_X1 U15061 ( .A1(n12854), .A2(n12853), .ZN(n12852) );
  MUX2_X1 U15062 ( .A(n14786), .B(n13069), .S(n12973), .Z(n12851) );
  NAND2_X1 U15063 ( .A1(n12852), .A2(n12851), .ZN(n12856) );
  OR2_X1 U15064 ( .A1(n12854), .A2(n12853), .ZN(n12855) );
  MUX2_X1 U15065 ( .A(n13068), .B(n12857), .S(n12997), .Z(n12861) );
  NAND2_X1 U15066 ( .A1(n12860), .A2(n12861), .ZN(n12859) );
  MUX2_X1 U15067 ( .A(n13068), .B(n12857), .S(n12973), .Z(n12858) );
  NAND2_X1 U15068 ( .A1(n12859), .A2(n12858), .ZN(n12865) );
  INV_X1 U15069 ( .A(n12860), .ZN(n12863) );
  INV_X1 U15070 ( .A(n12861), .ZN(n12862) );
  NAND2_X1 U15071 ( .A1(n12863), .A2(n12862), .ZN(n12864) );
  MUX2_X1 U15072 ( .A(n13067), .B(n13424), .S(n12973), .Z(n12867) );
  MUX2_X1 U15073 ( .A(n13067), .B(n13424), .S(n12997), .Z(n12866) );
  INV_X1 U15074 ( .A(n12867), .ZN(n12868) );
  MUX2_X1 U15075 ( .A(n13066), .B(n14639), .S(n12997), .Z(n12872) );
  NAND2_X1 U15076 ( .A1(n12871), .A2(n12872), .ZN(n12870) );
  MUX2_X1 U15077 ( .A(n13066), .B(n14639), .S(n12973), .Z(n12869) );
  NAND2_X1 U15078 ( .A1(n12870), .A2(n12869), .ZN(n12876) );
  INV_X1 U15079 ( .A(n12871), .ZN(n12874) );
  INV_X1 U15080 ( .A(n12872), .ZN(n12873) );
  NAND2_X1 U15081 ( .A1(n12874), .A2(n12873), .ZN(n12875) );
  NAND2_X1 U15082 ( .A1(n12876), .A2(n12875), .ZN(n12879) );
  MUX2_X1 U15083 ( .A(n13065), .B(n14844), .S(n12973), .Z(n12878) );
  MUX2_X1 U15084 ( .A(n13065), .B(n14844), .S(n12997), .Z(n12877) );
  MUX2_X1 U15085 ( .A(n13064), .B(n12880), .S(n12997), .Z(n12883) );
  MUX2_X1 U15086 ( .A(n13064), .B(n12880), .S(n12973), .Z(n12881) );
  NAND2_X1 U15087 ( .A1(n12882), .A2(n12881), .ZN(n12885) );
  NAND2_X1 U15088 ( .A1(n12885), .A2(n12884), .ZN(n12888) );
  MUX2_X1 U15089 ( .A(n13063), .B(n14658), .S(n12973), .Z(n12889) );
  MUX2_X1 U15090 ( .A(n13063), .B(n14658), .S(n12997), .Z(n12887) );
  INV_X1 U15091 ( .A(n12889), .ZN(n12890) );
  MUX2_X1 U15092 ( .A(n13062), .B(n13521), .S(n12997), .Z(n12893) );
  MUX2_X1 U15093 ( .A(n13062), .B(n13521), .S(n12973), .Z(n12891) );
  NAND2_X1 U15094 ( .A1(n12892), .A2(n12891), .ZN(n12896) );
  INV_X1 U15095 ( .A(n12893), .ZN(n12894) );
  MUX2_X1 U15096 ( .A(n13406), .B(n12897), .S(n12973), .Z(n12899) );
  MUX2_X1 U15097 ( .A(n13406), .B(n12897), .S(n12997), .Z(n12898) );
  MUX2_X1 U15098 ( .A(n13061), .B(n13514), .S(n12997), .Z(n12903) );
  MUX2_X1 U15099 ( .A(n13061), .B(n13514), .S(n12973), .Z(n12900) );
  INV_X1 U15100 ( .A(n12900), .ZN(n12901) );
  NAND2_X1 U15101 ( .A1(n13509), .A2(n12902), .ZN(n13178) );
  OR2_X1 U15102 ( .A1(n13509), .A2(n12902), .ZN(n13175) );
  MUX2_X1 U15103 ( .A(n13178), .B(n13175), .S(n12973), .Z(n12906) );
  NAND2_X1 U15104 ( .A1(n12904), .A2(n12903), .ZN(n12905) );
  NAND3_X1 U15105 ( .A1(n12907), .A2(n12906), .A3(n12905), .ZN(n12909) );
  MUX2_X1 U15106 ( .A(n13178), .B(n13175), .S(n12997), .Z(n12908) );
  NAND2_X1 U15107 ( .A1(n12909), .A2(n12908), .ZN(n12912) );
  INV_X1 U15108 ( .A(n13155), .ZN(n13180) );
  MUX2_X1 U15109 ( .A(n13180), .B(n13391), .S(n12997), .Z(n12911) );
  MUX2_X1 U15110 ( .A(n13155), .B(n13504), .S(n12973), .Z(n12910) );
  NAND2_X1 U15111 ( .A1(n12912), .A2(n12911), .ZN(n12913) );
  MUX2_X1 U15112 ( .A(n13375), .B(n13158), .S(n12997), .Z(n12916) );
  MUX2_X1 U15113 ( .A(n13158), .B(n13375), .S(n12997), .Z(n12915) );
  MUX2_X1 U15114 ( .A(n13160), .B(n13493), .S(n12997), .Z(n12919) );
  NAND2_X1 U15115 ( .A1(n12920), .A2(n12919), .ZN(n12918) );
  MUX2_X1 U15116 ( .A(n13160), .B(n13493), .S(n12973), .Z(n12917) );
  NAND2_X1 U15117 ( .A1(n12918), .A2(n12917), .ZN(n12922) );
  NAND2_X1 U15118 ( .A1(n12922), .A2(n12921), .ZN(n12925) );
  MUX2_X1 U15119 ( .A(n13162), .B(n13488), .S(n12973), .Z(n12924) );
  MUX2_X1 U15120 ( .A(n13162), .B(n13488), .S(n12997), .Z(n12923) );
  MUX2_X1 U15121 ( .A(n13164), .B(n13482), .S(n12997), .Z(n12928) );
  MUX2_X1 U15122 ( .A(n13164), .B(n13482), .S(n12973), .Z(n12926) );
  NAND2_X1 U15123 ( .A1(n12927), .A2(n12926), .ZN(n12930) );
  NAND2_X1 U15124 ( .A1(n12930), .A2(n12929), .ZN(n12933) );
  MUX2_X1 U15125 ( .A(n13286), .B(n13476), .S(n12973), .Z(n12932) );
  MUX2_X1 U15126 ( .A(n13286), .B(n13476), .S(n12997), .Z(n12931) );
  MUX2_X1 U15127 ( .A(n13311), .B(n13470), .S(n12997), .Z(n12936) );
  MUX2_X1 U15128 ( .A(n13311), .B(n13470), .S(n12973), .Z(n12934) );
  NAND2_X1 U15129 ( .A1(n12935), .A2(n12934), .ZN(n12939) );
  OR2_X1 U15130 ( .A1(n6521), .A2(n11760), .ZN(n12940) );
  NAND2_X1 U15131 ( .A1(n12958), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12944) );
  NAND2_X1 U15132 ( .A1(n12941), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n12943) );
  NAND2_X1 U15133 ( .A1(n12959), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n12942) );
  XNOR2_X1 U15134 ( .A(n13141), .B(n13145), .ZN(n13036) );
  MUX2_X1 U15135 ( .A(n13204), .B(n13542), .S(n12997), .Z(n12980) );
  MUX2_X1 U15136 ( .A(n13237), .B(n13228), .S(n12973), .Z(n12978) );
  INV_X1 U15137 ( .A(n13060), .ZN(n13001) );
  OAI21_X1 U15138 ( .B1(n12980), .B2(n12978), .A(n12979), .ZN(n12945) );
  MUX2_X1 U15139 ( .A(n13198), .B(n13240), .S(n12973), .Z(n12955) );
  MUX2_X1 U15140 ( .A(n13252), .B(n13454), .S(n12997), .Z(n12954) );
  INV_X1 U15141 ( .A(n13460), .ZN(n13259) );
  MUX2_X1 U15142 ( .A(n13274), .B(n13259), .S(n12973), .Z(n12988) );
  MUX2_X1 U15143 ( .A(n13238), .B(n13460), .S(n12997), .Z(n12987) );
  AND2_X1 U15144 ( .A1(n12988), .A2(n12987), .ZN(n12946) );
  NOR2_X1 U15145 ( .A1(n12989), .A2(n12946), .ZN(n12949) );
  MUX2_X1 U15146 ( .A(n13548), .B(n13195), .S(n12997), .Z(n12951) );
  MUX2_X1 U15147 ( .A(n13287), .B(n13276), .S(n12997), .Z(n12950) );
  NAND2_X1 U15148 ( .A1(n12951), .A2(n12950), .ZN(n12947) );
  INV_X1 U15149 ( .A(n12949), .ZN(n12993) );
  INV_X1 U15150 ( .A(n12950), .ZN(n12953) );
  INV_X1 U15151 ( .A(n12951), .ZN(n12952) );
  NAND2_X1 U15152 ( .A1(n12953), .A2(n12952), .ZN(n12992) );
  INV_X1 U15153 ( .A(n12954), .ZN(n12957) );
  INV_X1 U15154 ( .A(n12955), .ZN(n12956) );
  NAND2_X1 U15155 ( .A1(n12957), .A2(n12956), .ZN(n12984) );
  INV_X1 U15156 ( .A(n13145), .ZN(n13058) );
  NAND2_X1 U15157 ( .A1(n13058), .A2(n12997), .ZN(n12971) );
  MUX2_X1 U15158 ( .A(n12971), .B(n13058), .S(n13141), .Z(n12977) );
  NAND2_X1 U15159 ( .A1(n12958), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n12962) );
  NAND2_X1 U15160 ( .A1(n12941), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n12961) );
  NAND2_X1 U15161 ( .A1(n12959), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n12960) );
  NAND3_X1 U15162 ( .A1(n12962), .A2(n12961), .A3(n12960), .ZN(n13059) );
  NAND2_X1 U15163 ( .A1(n12964), .A2(n12963), .ZN(n12967) );
  OR2_X1 U15164 ( .A1(n6521), .A2(n13566), .ZN(n12966) );
  MUX2_X1 U15165 ( .A(n13059), .B(n13140), .S(n12997), .Z(n12996) );
  OAI211_X1 U15166 ( .C1(n14802), .C2(n12968), .A(n13048), .B(n13042), .ZN(
        n12969) );
  INV_X1 U15167 ( .A(n12969), .ZN(n12970) );
  INV_X1 U15168 ( .A(n13059), .ZN(n13206) );
  AOI21_X1 U15169 ( .B1(n12971), .B2(n12970), .A(n13206), .ZN(n12972) );
  AOI21_X1 U15170 ( .B1(n13140), .B2(n12973), .A(n12972), .ZN(n12995) );
  OAI22_X1 U15171 ( .A1(n12996), .A2(n12995), .B1(n12975), .B2(n12974), .ZN(
        n12976) );
  NAND2_X1 U15172 ( .A1(n12977), .A2(n12976), .ZN(n12983) );
  INV_X1 U15173 ( .A(n13036), .ZN(n12981) );
  NAND4_X1 U15174 ( .A1(n12981), .A2(n12980), .A3(n12979), .A4(n12978), .ZN(
        n12982) );
  OAI211_X1 U15175 ( .C1(n12985), .C2(n12984), .A(n12983), .B(n12982), .ZN(
        n12986) );
  INV_X1 U15176 ( .A(n12986), .ZN(n12991) );
  OAI211_X1 U15177 ( .C1(n12993), .C2(n12992), .A(n12991), .B(n12990), .ZN(
        n12994) );
  NAND2_X1 U15178 ( .A1(n12996), .A2(n12995), .ZN(n13000) );
  NAND3_X1 U15179 ( .A1(n13141), .A2(n13145), .A3(n12997), .ZN(n12999) );
  OR3_X1 U15180 ( .A1(n13141), .A2(n13145), .A3(n12997), .ZN(n12998) );
  INV_X1 U15181 ( .A(n13046), .ZN(n13051) );
  XNOR2_X1 U15182 ( .A(n13140), .B(n13206), .ZN(n13035) );
  NAND2_X1 U15183 ( .A1(n13228), .A2(n13237), .ZN(n13173) );
  OR2_X1 U15184 ( .A1(n13228), .A2(n13237), .ZN(n13002) );
  NAND2_X1 U15185 ( .A1(n13173), .A2(n13002), .ZN(n13172) );
  XNOR2_X1 U15186 ( .A(n13460), .B(n13274), .ZN(n13254) );
  XNOR2_X1 U15187 ( .A(n13276), .B(n13195), .ZN(n13269) );
  XNOR2_X1 U15188 ( .A(n13470), .B(n13273), .ZN(n13290) );
  XNOR2_X1 U15189 ( .A(n13482), .B(n13310), .ZN(n13326) );
  NAND2_X1 U15190 ( .A1(n13488), .A2(n13319), .ZN(n13189) );
  OR2_X1 U15191 ( .A1(n13488), .A2(n13319), .ZN(n13003) );
  NAND2_X1 U15192 ( .A1(n13189), .A2(n13003), .ZN(n13188) );
  INV_X1 U15193 ( .A(n13160), .ZN(n13185) );
  XNOR2_X1 U15194 ( .A(n13493), .B(n13185), .ZN(n13351) );
  XNOR2_X1 U15195 ( .A(n13375), .B(n13183), .ZN(n13371) );
  XNOR2_X1 U15196 ( .A(n13504), .B(n13155), .ZN(n13395) );
  AND2_X1 U15197 ( .A1(n13005), .A2(n13004), .ZN(n14823) );
  NAND4_X1 U15198 ( .A1(n13007), .A2(n14823), .A3(n9333), .A4(n13006), .ZN(
        n13009) );
  NOR2_X1 U15199 ( .A1(n13009), .A2(n13008), .ZN(n13013) );
  NAND4_X1 U15200 ( .A1(n13013), .A2(n13012), .A3(n13011), .A4(n13010), .ZN(
        n13014) );
  NOR2_X1 U15201 ( .A1(n13015), .A2(n13014), .ZN(n13018) );
  NAND4_X1 U15202 ( .A1(n13019), .A2(n13018), .A3(n13017), .A4(n13016), .ZN(
        n13020) );
  NOR2_X1 U15203 ( .A1(n13021), .A2(n13020), .ZN(n13024) );
  NAND4_X1 U15204 ( .A1(n13025), .A2(n13024), .A3(n13023), .A4(n13022), .ZN(
        n13026) );
  NOR2_X1 U15205 ( .A1(n13403), .A2(n13026), .ZN(n13029) );
  NAND4_X1 U15206 ( .A1(n13395), .A2(n13029), .A3(n13028), .A4(n13027), .ZN(
        n13030) );
  OR4_X1 U15207 ( .A1(n13188), .A2(n13351), .A3(n13371), .A4(n13030), .ZN(
        n13031) );
  OR4_X1 U15208 ( .A1(n13269), .A2(n13290), .A3(n13326), .A4(n13031), .ZN(
        n13032) );
  NOR2_X1 U15209 ( .A1(n13254), .A2(n13032), .ZN(n13033) );
  XNOR2_X1 U15210 ( .A(n13476), .B(n13286), .ZN(n13307) );
  NAND4_X1 U15211 ( .A1(n13172), .A2(n13033), .A3(n13247), .A4(n13307), .ZN(
        n13034) );
  XNOR2_X1 U15212 ( .A(n13037), .B(n13052), .ZN(n13038) );
  OAI21_X1 U15213 ( .B1(n13048), .B2(n13039), .A(n13412), .ZN(n13040) );
  OAI21_X1 U15214 ( .B1(n13049), .B2(n6571), .A(n13040), .ZN(n13041) );
  NAND3_X1 U15215 ( .A1(n13047), .A2(n13051), .A3(n13041), .ZN(n13056) );
  INV_X1 U15216 ( .A(n13042), .ZN(n13043) );
  NAND4_X1 U15217 ( .A1(n14817), .A2(n13044), .A3(n13043), .A4(n13405), .ZN(
        n13045) );
  OAI211_X1 U15218 ( .C1(n13049), .C2(n13046), .A(n13045), .B(P2_B_REG_SCAN_IN), .ZN(n13055) );
  MUX2_X1 U15219 ( .A(n13049), .B(n13048), .S(n9333), .Z(n13050) );
  NAND4_X1 U15220 ( .A1(n13053), .A2(n13052), .A3(n13051), .A4(n13050), .ZN(
        n13054) );
  NAND4_X1 U15221 ( .A1(n13057), .A2(n13056), .A3(n13055), .A4(n13054), .ZN(
        P2_U3328) );
  MUX2_X1 U15222 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13058), .S(n6523), .Z(
        P2_U3562) );
  MUX2_X1 U15223 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13059), .S(n6523), .Z(
        P2_U3561) );
  MUX2_X1 U15224 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13060), .S(n6523), .Z(
        P2_U3560) );
  MUX2_X1 U15225 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13237), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15226 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13252), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15227 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13238), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15228 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13287), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15229 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13311), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15230 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13286), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15231 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13164), .S(n6523), .Z(
        P2_U3553) );
  MUX2_X1 U15232 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13162), .S(n6523), .Z(
        P2_U3552) );
  MUX2_X1 U15233 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13160), .S(n6523), .Z(
        P2_U3551) );
  MUX2_X1 U15234 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13158), .S(n6523), .Z(
        P2_U3550) );
  MUX2_X1 U15235 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13155), .S(n6523), .Z(
        P2_U3549) );
  MUX2_X1 U15236 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13408), .S(n6523), .Z(
        P2_U3548) );
  MUX2_X1 U15237 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13061), .S(n6523), .Z(
        P2_U3547) );
  MUX2_X1 U15238 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13406), .S(n6523), .Z(
        P2_U3546) );
  MUX2_X1 U15239 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13062), .S(n6523), .Z(
        P2_U3545) );
  MUX2_X1 U15240 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13063), .S(n6523), .Z(
        P2_U3544) );
  MUX2_X1 U15241 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13064), .S(n6523), .Z(
        P2_U3543) );
  MUX2_X1 U15242 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13065), .S(n6523), .Z(
        P2_U3542) );
  MUX2_X1 U15243 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13066), .S(n6523), .Z(
        P2_U3541) );
  MUX2_X1 U15244 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13067), .S(n6523), .Z(
        P2_U3540) );
  MUX2_X1 U15245 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13068), .S(n6523), .Z(
        P2_U3539) );
  MUX2_X1 U15246 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13069), .S(n6523), .Z(
        P2_U3538) );
  MUX2_X1 U15247 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13070), .S(n6523), .Z(
        P2_U3537) );
  MUX2_X1 U15248 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13071), .S(n6523), .Z(
        P2_U3536) );
  MUX2_X1 U15249 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13072), .S(n6523), .Z(
        P2_U3535) );
  MUX2_X1 U15250 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13073), .S(n6523), .Z(
        P2_U3534) );
  MUX2_X1 U15251 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13074), .S(n6523), .Z(
        P2_U3533) );
  MUX2_X1 U15252 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13075), .S(n6523), .Z(
        P2_U3532) );
  MUX2_X1 U15253 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9385), .S(n6523), .Z(
        P2_U3531) );
  INV_X1 U15254 ( .A(n13082), .ZN(n13078) );
  INV_X1 U15255 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13076) );
  OAI22_X1 U15256 ( .A1(n14744), .A2(n7617), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13076), .ZN(n13077) );
  AOI21_X1 U15257 ( .B1(n13078), .B2(n14770), .A(n13077), .ZN(n13090) );
  INV_X1 U15258 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14856) );
  INV_X1 U15259 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n13085) );
  MUX2_X1 U15260 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9227), .S(n13082), .Z(
        n13079) );
  OAI21_X1 U15261 ( .B1(n14856), .B2(n13085), .A(n13079), .ZN(n13080) );
  NAND3_X1 U15262 ( .A1(n14774), .A2(n13081), .A3(n13080), .ZN(n13089) );
  INV_X1 U15263 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n14808) );
  MUX2_X1 U15264 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n13083), .S(n13082), .Z(
        n13084) );
  OAI21_X1 U15265 ( .B1(n14808), .B2(n13085), .A(n13084), .ZN(n13086) );
  NAND3_X1 U15266 ( .A1(n14776), .A2(n13087), .A3(n13086), .ZN(n13088) );
  NAND3_X1 U15267 ( .A1(n13090), .A2(n13089), .A3(n13088), .ZN(P2_U3215) );
  NAND2_X1 U15268 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n13091) );
  OAI21_X1 U15269 ( .B1(n14740), .B2(n13092), .A(n13091), .ZN(n13093) );
  AOI21_X1 U15270 ( .B1(n14768), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n13093), .ZN(
        n13105) );
  MUX2_X1 U15271 ( .A(n9914), .B(P2_REG2_REG_4__SCAN_IN), .S(n13098), .Z(
        n13094) );
  NAND3_X1 U15272 ( .A1(n14683), .A2(n13095), .A3(n13094), .ZN(n13096) );
  NAND3_X1 U15273 ( .A1(n14776), .A2(n13097), .A3(n13096), .ZN(n13104) );
  MUX2_X1 U15274 ( .A(n9232), .B(P2_REG1_REG_4__SCAN_IN), .S(n13098), .Z(
        n13099) );
  NAND3_X1 U15275 ( .A1(n14680), .A2(n13100), .A3(n13099), .ZN(n13101) );
  NAND3_X1 U15276 ( .A1(n14774), .A2(n13102), .A3(n13101), .ZN(n13103) );
  NAND3_X1 U15277 ( .A1(n13105), .A2(n13104), .A3(n13103), .ZN(P2_U3218) );
  NAND2_X1 U15278 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n13106) );
  OAI21_X1 U15279 ( .B1(n14740), .B2(n13107), .A(n13106), .ZN(n13108) );
  AOI21_X1 U15280 ( .B1(n14768), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n13108), .ZN(
        n13122) );
  MUX2_X1 U15281 ( .A(n9296), .B(P2_REG2_REG_8__SCAN_IN), .S(n13114), .Z(
        n13109) );
  NAND3_X1 U15282 ( .A1(n13111), .A2(n13110), .A3(n13109), .ZN(n13112) );
  NAND3_X1 U15283 ( .A1(n13113), .A2(n14776), .A3(n13112), .ZN(n13121) );
  INV_X1 U15284 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15262) );
  MUX2_X1 U15285 ( .A(n15262), .B(P2_REG1_REG_8__SCAN_IN), .S(n13114), .Z(
        n13115) );
  NAND3_X1 U15286 ( .A1(n13117), .A2(n13116), .A3(n13115), .ZN(n13118) );
  NAND3_X1 U15287 ( .A1(n13119), .A2(n14774), .A3(n13118), .ZN(n13120) );
  NAND3_X1 U15288 ( .A1(n13122), .A2(n13121), .A3(n13120), .ZN(P2_U3222) );
  INV_X1 U15289 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n15214) );
  NOR2_X1 U15290 ( .A1(n13128), .A2(n13123), .ZN(n13125) );
  NOR2_X1 U15291 ( .A1(n13125), .A2(n13124), .ZN(n13126) );
  XOR2_X1 U15292 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13126), .Z(n13135) );
  INV_X1 U15293 ( .A(n13135), .ZN(n13133) );
  NAND2_X1 U15294 ( .A1(n13128), .A2(n13127), .ZN(n13130) );
  NAND2_X1 U15295 ( .A1(n13130), .A2(n13129), .ZN(n13131) );
  XNOR2_X1 U15296 ( .A(n13500), .B(n13131), .ZN(n13134) );
  NOR2_X1 U15297 ( .A1(n13134), .A2(n14747), .ZN(n13132) );
  AOI211_X1 U15298 ( .C1(n13133), .C2(n14776), .A(n14770), .B(n13132), .ZN(
        n13137) );
  AOI22_X1 U15299 ( .A1(n13135), .A2(n14776), .B1(n14774), .B2(n13134), .ZN(
        n13136) );
  MUX2_X1 U15300 ( .A(n13137), .B(n13136), .S(n13412), .Z(n13139) );
  NAND2_X1 U15301 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3088), .ZN(n13138)
         );
  OAI211_X1 U15302 ( .C1(n15214), .C2(n14744), .A(n13139), .B(n13138), .ZN(
        P2_U3233) );
  NAND2_X1 U15303 ( .A1(n13359), .A2(n13347), .ZN(n13343) );
  AND2_X2 U15304 ( .A1(n13275), .A2(n13259), .ZN(n13260) );
  AND2_X2 U15305 ( .A1(n13260), .A2(n13240), .ZN(n13242) );
  XNOR2_X1 U15306 ( .A(n13149), .B(n13141), .ZN(n13142) );
  NOR2_X1 U15307 ( .A1(n13142), .A2(n9459), .ZN(n13432) );
  NAND2_X1 U15308 ( .A1(n13432), .A2(n13425), .ZN(n13147) );
  INV_X1 U15309 ( .A(P2_B_REG_SCAN_IN), .ZN(n13143) );
  OR2_X1 U15310 ( .A1(n13577), .A2(n13143), .ZN(n13144) );
  NAND2_X1 U15311 ( .A1(n13407), .A2(n13144), .ZN(n13205) );
  NOR2_X1 U15312 ( .A1(n13145), .A2(n13205), .ZN(n13431) );
  INV_X1 U15313 ( .A(n13431), .ZN(n13435) );
  NOR2_X1 U15314 ( .A1(n13435), .A2(n14811), .ZN(n13151) );
  AOI21_X1 U15315 ( .B1(n14811), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13151), 
        .ZN(n13146) );
  OAI211_X1 U15316 ( .C1(n13533), .C2(n13390), .A(n13147), .B(n13146), .ZN(
        P2_U3234) );
  OR2_X1 U15317 ( .A1(n13209), .A2(n13537), .ZN(n13148) );
  NAND3_X1 U15318 ( .A1(n13149), .A2(n13148), .A3(n10803), .ZN(n13436) );
  NOR2_X1 U15319 ( .A1(n13537), .A2(n13390), .ZN(n13150) );
  AOI211_X1 U15320 ( .C1(n14811), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13151), 
        .B(n13150), .ZN(n13152) );
  OAI21_X1 U15321 ( .B1(n14789), .B2(n13436), .A(n13152), .ZN(P2_U3235) );
  NAND2_X1 U15322 ( .A1(n13509), .A2(n13408), .ZN(n13153) );
  NAND2_X1 U15323 ( .A1(n13154), .A2(n13153), .ZN(n13394) );
  OR2_X2 U15324 ( .A1(n13394), .A2(n13395), .ZN(n13392) );
  OR2_X1 U15325 ( .A1(n13504), .A2(n13155), .ZN(n13156) );
  NOR2_X1 U15326 ( .A1(n13375), .A2(n13158), .ZN(n13157) );
  NAND2_X1 U15327 ( .A1(n13375), .A2(n13158), .ZN(n13159) );
  AND2_X1 U15328 ( .A1(n13493), .A2(n13160), .ZN(n13161) );
  NOR2_X1 U15329 ( .A1(n13488), .A2(n13162), .ZN(n13163) );
  NAND2_X1 U15330 ( .A1(n13327), .A2(n13326), .ZN(n13480) );
  NAND2_X1 U15331 ( .A1(n13482), .A2(n13164), .ZN(n13165) );
  OR2_X1 U15332 ( .A1(n13476), .A2(n13286), .ZN(n13166) );
  INV_X1 U15333 ( .A(n13290), .ZN(n13284) );
  NAND2_X1 U15334 ( .A1(n13470), .A2(n13311), .ZN(n13167) );
  OR2_X1 U15335 ( .A1(n13276), .A2(n13287), .ZN(n13168) );
  NAND2_X1 U15336 ( .A1(n13267), .A2(n13168), .ZN(n13170) );
  NAND2_X1 U15337 ( .A1(n13276), .A2(n13287), .ZN(n13169) );
  AND2_X1 U15338 ( .A1(n13460), .A2(n13238), .ZN(n13171) );
  NAND2_X1 U15339 ( .A1(n13224), .A2(n13223), .ZN(n13222) );
  NAND2_X1 U15340 ( .A1(n13222), .A2(n13173), .ZN(n13174) );
  INV_X1 U15341 ( .A(n13175), .ZN(n13176) );
  OR2_X2 U15342 ( .A1(n13177), .A2(n13176), .ZN(n13179) );
  AND2_X1 U15343 ( .A1(n13504), .A2(n13180), .ZN(n13182) );
  NOR2_X1 U15344 ( .A1(n13375), .A2(n13183), .ZN(n13184) );
  INV_X1 U15345 ( .A(n13351), .ZN(n13353) );
  NAND2_X1 U15346 ( .A1(n13493), .A2(n13185), .ZN(n13186) );
  OR2_X1 U15347 ( .A1(n13482), .A2(n13310), .ZN(n13190) );
  INV_X1 U15348 ( .A(n13286), .ZN(n13320) );
  NAND2_X1 U15349 ( .A1(n13476), .A2(n13320), .ZN(n13191) );
  OR2_X1 U15350 ( .A1(n13476), .A2(n13320), .ZN(n13192) );
  NAND2_X1 U15351 ( .A1(n13470), .A2(n13273), .ZN(n13268) );
  INV_X1 U15352 ( .A(n13269), .ZN(n13266) );
  NAND2_X1 U15353 ( .A1(n13276), .A2(n13195), .ZN(n13196) );
  OR2_X1 U15354 ( .A1(n13460), .A2(n13274), .ZN(n13197) );
  NAND2_X1 U15355 ( .A1(n13454), .A2(n13198), .ZN(n13199) );
  NAND2_X1 U15356 ( .A1(n13200), .A2(n13199), .ZN(n13216) );
  INV_X1 U15357 ( .A(n13216), .ZN(n13201) );
  OAI21_X1 U15358 ( .B1(n13204), .B2(n13228), .A(n13218), .ZN(n13203) );
  NOR2_X1 U15359 ( .A1(n13206), .A2(n13205), .ZN(n13207) );
  AOI21_X1 U15360 ( .B1(n13237), .B2(n13405), .A(n13207), .ZN(n13208) );
  NAND2_X1 U15361 ( .A1(n13442), .A2(n14809), .ZN(n13215) );
  AOI211_X1 U15362 ( .C1(n13439), .C2(n13231), .A(n9459), .B(n13209), .ZN(
        n13441) );
  AOI22_X1 U15363 ( .A1(n14811), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n13210), 
        .B2(n14783), .ZN(n13211) );
  OAI21_X1 U15364 ( .B1(n13212), .B2(n13390), .A(n13211), .ZN(n13213) );
  AOI21_X1 U15365 ( .B1(n13441), .B2(n13425), .A(n13213), .ZN(n13214) );
  OAI211_X1 U15366 ( .C1(n13444), .C2(n13396), .A(n13215), .B(n13214), .ZN(
        P2_U3236) );
  NAND2_X1 U15367 ( .A1(n13216), .A2(n13223), .ZN(n13217) );
  NAND3_X1 U15368 ( .A1(n13218), .A2(n14798), .A3(n13217), .ZN(n13221) );
  INV_X1 U15369 ( .A(n13219), .ZN(n13220) );
  NAND2_X1 U15370 ( .A1(n13221), .A2(n13220), .ZN(n13447) );
  OAI21_X1 U15371 ( .B1(n13224), .B2(n13223), .A(n13222), .ZN(n13445) );
  INV_X1 U15372 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13226) );
  OAI22_X1 U15373 ( .A1(n14809), .A2(n13226), .B1(n13225), .B2(n14803), .ZN(
        n13227) );
  AOI21_X1 U15374 ( .B1(n13228), .B2(n14785), .A(n13227), .ZN(n13233) );
  INV_X1 U15375 ( .A(n13242), .ZN(n13229) );
  AOI21_X1 U15376 ( .B1(n13229), .B2(n13228), .A(n9459), .ZN(n13230) );
  AND2_X1 U15377 ( .A1(n13231), .A2(n13230), .ZN(n13446) );
  NAND2_X1 U15378 ( .A1(n13446), .A2(n13425), .ZN(n13232) );
  OAI211_X1 U15379 ( .C1(n13445), .C2(n13396), .A(n13233), .B(n13232), .ZN(
        n13234) );
  AOI21_X1 U15380 ( .B1(n13447), .B2(n14809), .A(n13234), .ZN(n13235) );
  INV_X1 U15381 ( .A(n13235), .ZN(P2_U3237) );
  XNOR2_X1 U15382 ( .A(n13236), .B(n13247), .ZN(n13239) );
  OAI21_X1 U15383 ( .B1(n13260), .B2(n13240), .A(n10803), .ZN(n13241) );
  AOI22_X1 U15384 ( .A1(n14811), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13243), 
        .B2(n14783), .ZN(n13245) );
  NAND2_X1 U15385 ( .A1(n13454), .A2(n14785), .ZN(n13244) );
  OAI211_X1 U15386 ( .C1(n13457), .C2(n14789), .A(n13245), .B(n13244), .ZN(
        n13246) );
  INV_X1 U15387 ( .A(n13246), .ZN(n13250) );
  NAND2_X1 U15388 ( .A1(n13248), .A2(n13247), .ZN(n13452) );
  NAND3_X1 U15389 ( .A1(n13453), .A2(n13452), .A3(n14792), .ZN(n13249) );
  OAI211_X1 U15390 ( .C1(n13458), .C2(n14811), .A(n13250), .B(n13249), .ZN(
        P2_U3238) );
  XOR2_X1 U15391 ( .A(n13254), .B(n13251), .Z(n13253) );
  AOI222_X1 U15392 ( .A1(n14798), .A2(n13253), .B1(n13252), .B2(n13407), .C1(
        n13287), .C2(n13405), .ZN(n13462) );
  XNOR2_X1 U15393 ( .A(n13255), .B(n13254), .ZN(n13463) );
  INV_X1 U15394 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13257) );
  OAI22_X1 U15395 ( .A1(n14809), .A2(n13257), .B1(n13256), .B2(n14803), .ZN(
        n13258) );
  AOI21_X1 U15396 ( .B1(n13460), .B2(n14785), .A(n13258), .ZN(n13263) );
  OAI21_X1 U15397 ( .B1(n13275), .B2(n13259), .A(n10803), .ZN(n13261) );
  NOR2_X1 U15398 ( .A1(n13261), .A2(n13260), .ZN(n13459) );
  NAND2_X1 U15399 ( .A1(n13459), .A2(n13425), .ZN(n13262) );
  OAI211_X1 U15400 ( .C1(n13463), .C2(n13396), .A(n13263), .B(n13262), .ZN(
        n13264) );
  INV_X1 U15401 ( .A(n13264), .ZN(n13265) );
  OAI21_X1 U15402 ( .B1(n13462), .B2(n14811), .A(n13265), .ZN(P2_U3239) );
  XNOR2_X1 U15403 ( .A(n13267), .B(n13266), .ZN(n13466) );
  INV_X1 U15404 ( .A(n13466), .ZN(n13282) );
  NAND3_X1 U15405 ( .A1(n13283), .A2(n13269), .A3(n13268), .ZN(n13270) );
  AND2_X1 U15406 ( .A1(n13271), .A2(n13270), .ZN(n13272) );
  OAI222_X1 U15407 ( .A1(n14799), .A2(n13274), .B1(n13318), .B2(n13273), .C1(
        n13369), .C2(n13272), .ZN(n13464) );
  AOI211_X1 U15408 ( .C1(n13276), .C2(n6569), .A(n9459), .B(n13275), .ZN(
        n13465) );
  NAND2_X1 U15409 ( .A1(n13465), .A2(n13425), .ZN(n13279) );
  AOI22_X1 U15410 ( .A1(n14811), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13277), 
        .B2(n14783), .ZN(n13278) );
  OAI211_X1 U15411 ( .C1(n13548), .C2(n13390), .A(n13279), .B(n13278), .ZN(
        n13280) );
  AOI21_X1 U15412 ( .B1(n13464), .B2(n14809), .A(n13280), .ZN(n13281) );
  OAI21_X1 U15413 ( .B1(n13282), .B2(n13396), .A(n13281), .ZN(P2_U3240) );
  OAI21_X1 U15414 ( .B1(n13285), .B2(n13284), .A(n13283), .ZN(n13288) );
  AOI222_X1 U15415 ( .A1(n14798), .A2(n13288), .B1(n13287), .B2(n13407), .C1(
        n13286), .C2(n13405), .ZN(n13472) );
  OAI21_X1 U15416 ( .B1(n13290), .B2(n6622), .A(n13289), .ZN(n13473) );
  INV_X1 U15417 ( .A(n13473), .ZN(n13297) );
  INV_X1 U15418 ( .A(n13470), .ZN(n13295) );
  AOI21_X1 U15419 ( .B1(n13302), .B2(n13470), .A(n9459), .ZN(n13291) );
  AND2_X1 U15420 ( .A1(n13291), .A2(n6569), .ZN(n13469) );
  NAND2_X1 U15421 ( .A1(n13469), .A2(n13425), .ZN(n13294) );
  AOI22_X1 U15422 ( .A1(n14811), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13292), 
        .B2(n14783), .ZN(n13293) );
  OAI211_X1 U15423 ( .C1(n13295), .C2(n13390), .A(n13294), .B(n13293), .ZN(
        n13296) );
  AOI21_X1 U15424 ( .B1(n13297), .B2(n14792), .A(n13296), .ZN(n13298) );
  OAI21_X1 U15425 ( .B1(n13472), .B2(n14811), .A(n13298), .ZN(P2_U3241) );
  INV_X1 U15426 ( .A(n13299), .ZN(n13300) );
  AOI21_X1 U15427 ( .B1(n13307), .B2(n13301), .A(n13300), .ZN(n13479) );
  INV_X1 U15428 ( .A(n13302), .ZN(n13303) );
  AOI211_X1 U15429 ( .C1(n13476), .C2(n13324), .A(n9459), .B(n13303), .ZN(
        n13474) );
  AOI22_X1 U15430 ( .A1(n13304), .A2(n14783), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14811), .ZN(n13305) );
  OAI21_X1 U15431 ( .B1(n7229), .B2(n13390), .A(n13305), .ZN(n13306) );
  AOI21_X1 U15432 ( .B1(n13474), .B2(n13425), .A(n13306), .ZN(n13316) );
  XOR2_X1 U15433 ( .A(n13308), .B(n13307), .Z(n13309) );
  NAND2_X1 U15434 ( .A1(n13309), .A2(n14798), .ZN(n13477) );
  INV_X1 U15435 ( .A(n13477), .ZN(n13314) );
  OR2_X1 U15436 ( .A1(n13310), .A2(n13318), .ZN(n13313) );
  NAND2_X1 U15437 ( .A1(n13311), .A2(n13407), .ZN(n13312) );
  NAND2_X1 U15438 ( .A1(n13313), .A2(n13312), .ZN(n13475) );
  OAI21_X1 U15439 ( .B1(n13314), .B2(n13475), .A(n14809), .ZN(n13315) );
  OAI211_X1 U15440 ( .C1(n13479), .C2(n13396), .A(n13316), .B(n13315), .ZN(
        P2_U3242) );
  AOI21_X1 U15441 ( .B1(n13317), .B2(n13326), .A(n13369), .ZN(n13323) );
  OAI22_X1 U15442 ( .A1(n13320), .A2(n14799), .B1(n13319), .B2(n13318), .ZN(
        n13321) );
  AOI21_X1 U15443 ( .B1(n13323), .B2(n13322), .A(n13321), .ZN(n13485) );
  AOI21_X1 U15444 ( .B1(n13482), .B2(n13343), .A(n9459), .ZN(n13325) );
  NAND2_X1 U15445 ( .A1(n13325), .A2(n13324), .ZN(n13483) );
  OR2_X1 U15446 ( .A1(n13327), .A2(n13326), .ZN(n13481) );
  NAND3_X1 U15447 ( .A1(n13481), .A2(n13480), .A3(n14792), .ZN(n13332) );
  INV_X1 U15448 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13328) );
  OAI22_X1 U15449 ( .A1(n13329), .A2(n14803), .B1(n13328), .B2(n14809), .ZN(
        n13330) );
  AOI21_X1 U15450 ( .B1(n13482), .B2(n14785), .A(n13330), .ZN(n13331) );
  OAI211_X1 U15451 ( .C1(n13483), .C2(n14789), .A(n13332), .B(n13331), .ZN(
        n13333) );
  INV_X1 U15452 ( .A(n13333), .ZN(n13334) );
  OAI21_X1 U15453 ( .B1(n14811), .B2(n13485), .A(n13334), .ZN(P2_U3243) );
  XNOR2_X1 U15454 ( .A(n13335), .B(n13338), .ZN(n13491) );
  OAI21_X1 U15455 ( .B1(n13338), .B2(n13337), .A(n13336), .ZN(n13341) );
  INV_X1 U15456 ( .A(n13339), .ZN(n13340) );
  AOI21_X1 U15457 ( .B1(n13341), .B2(n14798), .A(n13340), .ZN(n13490) );
  INV_X1 U15458 ( .A(n13490), .ZN(n13349) );
  OR2_X1 U15459 ( .A1(n13359), .A2(n13347), .ZN(n13342) );
  AND3_X1 U15460 ( .A1(n13343), .A2(n10803), .A3(n13342), .ZN(n13487) );
  NAND2_X1 U15461 ( .A1(n13487), .A2(n13425), .ZN(n13346) );
  AOI22_X1 U15462 ( .A1(n13344), .A2(n14783), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n14811), .ZN(n13345) );
  OAI211_X1 U15463 ( .C1(n13347), .C2(n13390), .A(n13346), .B(n13345), .ZN(
        n13348) );
  AOI21_X1 U15464 ( .B1(n13349), .B2(n14809), .A(n13348), .ZN(n13350) );
  OAI21_X1 U15465 ( .B1(n13491), .B2(n13396), .A(n13350), .ZN(P2_U3244) );
  XNOR2_X1 U15466 ( .A(n13352), .B(n13351), .ZN(n13496) );
  XNOR2_X1 U15467 ( .A(n13354), .B(n13353), .ZN(n13356) );
  AOI21_X1 U15468 ( .B1(n13356), .B2(n14798), .A(n13355), .ZN(n13495) );
  INV_X1 U15469 ( .A(n13495), .ZN(n13365) );
  INV_X1 U15470 ( .A(n13493), .ZN(n13363) );
  NAND2_X1 U15471 ( .A1(n13373), .A2(n13493), .ZN(n13357) );
  NAND2_X1 U15472 ( .A1(n13357), .A2(n10803), .ZN(n13358) );
  NOR2_X1 U15473 ( .A1(n13359), .A2(n13358), .ZN(n13492) );
  NAND2_X1 U15474 ( .A1(n13492), .A2(n13425), .ZN(n13362) );
  AOI22_X1 U15475 ( .A1(n13360), .A2(n14783), .B1(n14811), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n13361) );
  OAI211_X1 U15476 ( .C1(n13363), .C2(n13390), .A(n13362), .B(n13361), .ZN(
        n13364) );
  AOI21_X1 U15477 ( .B1(n13365), .B2(n14809), .A(n13364), .ZN(n13366) );
  OAI21_X1 U15478 ( .B1(n13496), .B2(n13396), .A(n13366), .ZN(P2_U3245) );
  XOR2_X1 U15479 ( .A(n13371), .B(n13367), .Z(n13370) );
  OAI21_X1 U15480 ( .B1(n13370), .B2(n13369), .A(n13368), .ZN(n13497) );
  INV_X1 U15481 ( .A(n13497), .ZN(n13381) );
  XNOR2_X1 U15482 ( .A(n13372), .B(n13371), .ZN(n13499) );
  INV_X1 U15483 ( .A(n13373), .ZN(n13374) );
  AOI211_X1 U15484 ( .C1(n13375), .C2(n13385), .A(n9459), .B(n13374), .ZN(
        n13498) );
  NAND2_X1 U15485 ( .A1(n13498), .A2(n13425), .ZN(n13378) );
  AOI22_X1 U15486 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(n14811), .B1(n13376), 
        .B2(n14783), .ZN(n13377) );
  OAI211_X1 U15487 ( .C1(n7237), .C2(n13390), .A(n13378), .B(n13377), .ZN(
        n13379) );
  AOI21_X1 U15488 ( .B1(n13499), .B2(n14792), .A(n13379), .ZN(n13380) );
  OAI21_X1 U15489 ( .B1(n13381), .B2(n14811), .A(n13380), .ZN(P2_U3246) );
  XNOR2_X1 U15490 ( .A(n13382), .B(n13395), .ZN(n13384) );
  AOI21_X1 U15491 ( .B1(n13384), .B2(n14798), .A(n13383), .ZN(n13506) );
  AOI211_X1 U15492 ( .C1(n13504), .C2(n13386), .A(n9459), .B(n7238), .ZN(
        n13503) );
  INV_X1 U15493 ( .A(n13387), .ZN(n13388) );
  AOI22_X1 U15494 ( .A1(n14811), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13388), 
        .B2(n14783), .ZN(n13389) );
  OAI21_X1 U15495 ( .B1(n13391), .B2(n13390), .A(n13389), .ZN(n13398) );
  INV_X1 U15496 ( .A(n13392), .ZN(n13393) );
  AOI21_X1 U15497 ( .B1(n13395), .B2(n13394), .A(n13393), .ZN(n13507) );
  NOR2_X1 U15498 ( .A1(n13507), .A2(n13396), .ZN(n13397) );
  AOI211_X1 U15499 ( .C1(n13503), .C2(n13425), .A(n13398), .B(n13397), .ZN(
        n13399) );
  OAI21_X1 U15500 ( .B1(n14811), .B2(n13506), .A(n13399), .ZN(P2_U3247) );
  AOI211_X1 U15501 ( .C1(n13514), .C2(n13401), .A(n9459), .B(n13400), .ZN(
        n13513) );
  NOR2_X1 U15502 ( .A1(n13402), .A2(n14803), .ZN(n13411) );
  XNOR2_X1 U15503 ( .A(n13404), .B(n13403), .ZN(n13409) );
  AOI222_X1 U15504 ( .A1(n14798), .A2(n13409), .B1(n13408), .B2(n13407), .C1(
        n13406), .C2(n13405), .ZN(n13519) );
  INV_X1 U15505 ( .A(n13519), .ZN(n13410) );
  AOI211_X1 U15506 ( .C1(n13513), .C2(n13412), .A(n13411), .B(n13410), .ZN(
        n13417) );
  AOI22_X1 U15507 ( .A1(n13514), .A2(n14785), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n14811), .ZN(n13416) );
  NAND2_X1 U15508 ( .A1(n13414), .A2(n13413), .ZN(n13515) );
  NAND3_X1 U15509 ( .A1(n13516), .A2(n13515), .A3(n14792), .ZN(n13415) );
  OAI211_X1 U15510 ( .C1(n13417), .C2(n14811), .A(n13416), .B(n13415), .ZN(
        P2_U3249) );
  NAND2_X1 U15511 ( .A1(n13418), .A2(n14792), .ZN(n13430) );
  NAND2_X1 U15512 ( .A1(n13419), .A2(n14809), .ZN(n13429) );
  INV_X1 U15513 ( .A(n13420), .ZN(n13421) );
  OAI22_X1 U15514 ( .A1(n14809), .A2(n13422), .B1(n13421), .B2(n14803), .ZN(
        n13423) );
  AOI21_X1 U15515 ( .B1(n13424), .B2(n14785), .A(n13423), .ZN(n13428) );
  NAND2_X1 U15516 ( .A1(n13426), .A2(n13425), .ZN(n13427) );
  NAND4_X1 U15517 ( .A1(n13430), .A2(n13429), .A3(n13428), .A4(n13427), .ZN(
        P2_U3256) );
  INV_X1 U15518 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13433) );
  NOR2_X1 U15519 ( .A1(n13432), .A2(n13431), .ZN(n13530) );
  MUX2_X1 U15520 ( .A(n13433), .B(n13530), .S(n14861), .Z(n13434) );
  OAI21_X1 U15521 ( .B1(n13533), .B2(n13502), .A(n13434), .ZN(P2_U3530) );
  NAND2_X1 U15522 ( .A1(n13436), .A2(n13435), .ZN(n13534) );
  MUX2_X1 U15523 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13534), .S(n14861), .Z(
        n13437) );
  INV_X1 U15524 ( .A(n13437), .ZN(n13438) );
  OAI21_X1 U15525 ( .B1(n13537), .B2(n13502), .A(n13438), .ZN(P2_U3529) );
  OAI21_X1 U15526 ( .B1(n13444), .B2(n13529), .A(n13443), .ZN(n13538) );
  MUX2_X1 U15527 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13538), .S(n14861), .Z(
        P2_U3528) );
  NOR2_X1 U15528 ( .A1(n13447), .A2(n13446), .ZN(n13448) );
  OR2_X1 U15529 ( .A1(n13540), .A2(n13449), .ZN(n13450) );
  NAND2_X1 U15530 ( .A1(n13450), .A2(n7538), .ZN(n13451) );
  OAI21_X1 U15531 ( .B1(n13542), .B2(n13502), .A(n13451), .ZN(P2_U3527) );
  NAND3_X1 U15532 ( .A1(n13453), .A2(n14833), .A3(n13452), .ZN(n13456) );
  NAND2_X1 U15533 ( .A1(n13454), .A2(n14843), .ZN(n13455) );
  MUX2_X1 U15534 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13543), .S(n14861), .Z(
        P2_U3526) );
  AOI21_X1 U15535 ( .B1(n14843), .B2(n13460), .A(n13459), .ZN(n13461) );
  OAI211_X1 U15536 ( .C1(n13529), .C2(n13463), .A(n13462), .B(n13461), .ZN(
        n13544) );
  MUX2_X1 U15537 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13544), .S(n14861), .Z(
        P2_U3525) );
  INV_X1 U15538 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13467) );
  AOI211_X1 U15539 ( .C1(n14833), .C2(n13466), .A(n13465), .B(n13464), .ZN(
        n13545) );
  MUX2_X1 U15540 ( .A(n13467), .B(n13545), .S(n14861), .Z(n13468) );
  OAI21_X1 U15541 ( .B1(n13548), .B2(n13502), .A(n13468), .ZN(P2_U3524) );
  AOI21_X1 U15542 ( .B1(n14843), .B2(n13470), .A(n13469), .ZN(n13471) );
  OAI211_X1 U15543 ( .C1(n13529), .C2(n13473), .A(n13472), .B(n13471), .ZN(
        n13549) );
  MUX2_X1 U15544 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13549), .S(n14861), .Z(
        P2_U3523) );
  AOI211_X1 U15545 ( .C1(n14843), .C2(n13476), .A(n13475), .B(n13474), .ZN(
        n13478) );
  OAI211_X1 U15546 ( .C1(n13479), .C2(n13529), .A(n13478), .B(n13477), .ZN(
        n13550) );
  MUX2_X1 U15547 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13550), .S(n14861), .Z(
        P2_U3522) );
  NAND3_X1 U15548 ( .A1(n13481), .A2(n14833), .A3(n13480), .ZN(n13486) );
  NAND2_X1 U15549 ( .A1(n13482), .A2(n14843), .ZN(n13484) );
  NAND4_X1 U15550 ( .A1(n13486), .A2(n13485), .A3(n13484), .A4(n13483), .ZN(
        n13551) );
  MUX2_X1 U15551 ( .A(n13551), .B(P2_REG1_REG_22__SCAN_IN), .S(n13449), .Z(
        P2_U3521) );
  AOI21_X1 U15552 ( .B1(n14843), .B2(n13488), .A(n13487), .ZN(n13489) );
  OAI211_X1 U15553 ( .C1(n13491), .C2(n13529), .A(n13490), .B(n13489), .ZN(
        n13552) );
  MUX2_X1 U15554 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13552), .S(n14861), .Z(
        P2_U3520) );
  AOI21_X1 U15555 ( .B1(n14843), .B2(n13493), .A(n13492), .ZN(n13494) );
  OAI211_X1 U15556 ( .C1(n13496), .C2(n13529), .A(n13495), .B(n13494), .ZN(
        n13553) );
  MUX2_X1 U15557 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13553), .S(n14861), .Z(
        P2_U3519) );
  AOI211_X1 U15558 ( .C1(n13499), .C2(n14833), .A(n13498), .B(n13497), .ZN(
        n13554) );
  MUX2_X1 U15559 ( .A(n13500), .B(n13554), .S(n14861), .Z(n13501) );
  OAI21_X1 U15560 ( .B1(n7237), .B2(n13502), .A(n13501), .ZN(P2_U3518) );
  AOI21_X1 U15561 ( .B1(n14843), .B2(n13504), .A(n13503), .ZN(n13505) );
  OAI211_X1 U15562 ( .C1(n13507), .C2(n13529), .A(n13506), .B(n13505), .ZN(
        n13557) );
  MUX2_X1 U15563 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13557), .S(n14861), .Z(
        P2_U3517) );
  AOI21_X1 U15564 ( .B1(n14843), .B2(n13509), .A(n13508), .ZN(n13510) );
  OAI211_X1 U15565 ( .C1(n13512), .C2(n13529), .A(n13511), .B(n13510), .ZN(
        n13558) );
  MUX2_X1 U15566 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13558), .S(n14861), .Z(
        P2_U3516) );
  AOI21_X1 U15567 ( .B1(n14843), .B2(n13514), .A(n13513), .ZN(n13518) );
  NAND3_X1 U15568 ( .A1(n13516), .A2(n14833), .A3(n13515), .ZN(n13517) );
  NAND3_X1 U15569 ( .A1(n13519), .A2(n13518), .A3(n13517), .ZN(n13559) );
  MUX2_X1 U15570 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13559), .S(n14861), .Z(
        P2_U3515) );
  AOI21_X1 U15571 ( .B1(n14843), .B2(n13521), .A(n13520), .ZN(n13522) );
  OAI211_X1 U15572 ( .C1(n13529), .C2(n13524), .A(n13523), .B(n13522), .ZN(
        n13560) );
  MUX2_X1 U15573 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13560), .S(n14861), .Z(
        P2_U3513) );
  AOI211_X1 U15574 ( .C1(n14843), .C2(n14658), .A(n13526), .B(n13525), .ZN(
        n13527) );
  OAI21_X1 U15575 ( .B1(n13529), .B2(n13528), .A(n13527), .ZN(n13561) );
  MUX2_X1 U15576 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13561), .S(n14861), .Z(
        P2_U3512) );
  INV_X1 U15577 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13531) );
  MUX2_X1 U15578 ( .A(n13531), .B(n13530), .S(n14855), .Z(n13532) );
  OAI21_X1 U15579 ( .B1(n13533), .B2(n13556), .A(n13532), .ZN(P2_U3498) );
  MUX2_X1 U15580 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13534), .S(n14855), .Z(
        n13535) );
  INV_X1 U15581 ( .A(n13535), .ZN(n13536) );
  OAI21_X1 U15582 ( .B1(n13537), .B2(n13556), .A(n13536), .ZN(P2_U3497) );
  MUX2_X1 U15583 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13538), .S(n14855), .Z(
        P2_U3496) );
  OAI21_X1 U15584 ( .B1(n13542), .B2(n13556), .A(n13541), .ZN(P2_U3495) );
  MUX2_X1 U15585 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13543), .S(n14855), .Z(
        P2_U3494) );
  MUX2_X1 U15586 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13544), .S(n14855), .Z(
        P2_U3493) );
  INV_X1 U15587 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13546) );
  MUX2_X1 U15588 ( .A(n13546), .B(n13545), .S(n14855), .Z(n13547) );
  OAI21_X1 U15589 ( .B1(n13548), .B2(n13556), .A(n13547), .ZN(P2_U3492) );
  MUX2_X1 U15590 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13549), .S(n14855), .Z(
        P2_U3491) );
  MUX2_X1 U15591 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13550), .S(n14855), .Z(
        P2_U3490) );
  MUX2_X1 U15592 ( .A(n13551), .B(P2_REG0_REG_22__SCAN_IN), .S(n13539), .Z(
        P2_U3489) );
  MUX2_X1 U15593 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13552), .S(n14855), .Z(
        P2_U3488) );
  MUX2_X1 U15594 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13553), .S(n14855), .Z(
        P2_U3487) );
  INV_X1 U15595 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n15225) );
  MUX2_X1 U15596 ( .A(n15225), .B(n13554), .S(n14855), .Z(n13555) );
  OAI21_X1 U15597 ( .B1(n7237), .B2(n13556), .A(n13555), .ZN(P2_U3486) );
  MUX2_X1 U15598 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13557), .S(n14855), .Z(
        P2_U3484) );
  MUX2_X1 U15599 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13558), .S(n14855), .Z(
        P2_U3481) );
  MUX2_X1 U15600 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13559), .S(n14855), .Z(
        P2_U3478) );
  MUX2_X1 U15601 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13560), .S(n14855), .Z(
        P2_U3472) );
  MUX2_X1 U15602 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13561), .S(n14855), .Z(
        P2_U3469) );
  NAND3_X1 U15603 ( .A1(n9320), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13562) );
  OAI22_X1 U15604 ( .A1(n6545), .A2(n13562), .B1(n11760), .B2(n13580), .ZN(
        n13563) );
  AOI21_X1 U15605 ( .B1(n14297), .B2(n13564), .A(n13563), .ZN(n13565) );
  INV_X1 U15606 ( .A(n13565), .ZN(P2_U3296) );
  OAI222_X1 U15607 ( .A1(n13578), .A2(n13567), .B1(P2_U3088), .B2(n9324), .C1(
        n13566), .C2(n13580), .ZN(P2_U3297) );
  INV_X1 U15608 ( .A(n13568), .ZN(n14300) );
  OAI222_X1 U15609 ( .A1(n13580), .A2(n13570), .B1(n13578), .B2(n14300), .C1(
        n13569), .C2(P2_U3088), .ZN(P2_U3298) );
  AOI21_X1 U15610 ( .B1(n13572), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13571), 
        .ZN(n13573) );
  OAI21_X1 U15611 ( .B1(n13575), .B2(n13574), .A(n13573), .ZN(P2_U3299) );
  INV_X1 U15612 ( .A(n13576), .ZN(n14304) );
  OAI222_X1 U15613 ( .A1(n13580), .A2(n13579), .B1(n13578), .B2(n14304), .C1(
        n13577), .C2(P2_U3088), .ZN(P2_U3300) );
  MUX2_X1 U15614 ( .A(n13581), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI22_X1 U15615 ( .A1(n14012), .A2(n13741), .B1(n13582), .B2(n13740), .ZN(
        n13734) );
  NAND2_X1 U15616 ( .A1(n14195), .A2(n13702), .ZN(n13584) );
  NAND2_X1 U15617 ( .A1(n13840), .A2(n13697), .ZN(n13583) );
  NAND2_X1 U15618 ( .A1(n13584), .A2(n13583), .ZN(n13585) );
  XNOR2_X1 U15619 ( .A(n13585), .B(n13705), .ZN(n13733) );
  XOR2_X1 U15620 ( .A(n13734), .B(n13733), .Z(n13737) );
  NAND2_X1 U15621 ( .A1(n14504), .A2(n13702), .ZN(n13587) );
  NAND2_X1 U15622 ( .A1(n13848), .A2(n13697), .ZN(n13586) );
  NAND2_X1 U15623 ( .A1(n13587), .A2(n13586), .ZN(n13588) );
  XNOR2_X1 U15624 ( .A(n13588), .B(n13705), .ZN(n13598) );
  NOR2_X1 U15625 ( .A1(n13589), .A2(n13740), .ZN(n13590) );
  AOI21_X1 U15626 ( .B1(n14504), .B2(n13697), .A(n13590), .ZN(n13596) );
  XNOR2_X1 U15627 ( .A(n13598), .B(n13596), .ZN(n14473) );
  INV_X1 U15628 ( .A(n13591), .ZN(n13592) );
  NAND2_X1 U15629 ( .A1(n13593), .A2(n13592), .ZN(n14474) );
  AND2_X1 U15630 ( .A1(n14473), .A2(n14474), .ZN(n13594) );
  INV_X1 U15631 ( .A(n13596), .ZN(n13597) );
  NOR2_X1 U15632 ( .A1(n14472), .A2(n13740), .ZN(n13600) );
  AOI21_X1 U15633 ( .B1(n13601), .B2(n13697), .A(n13600), .ZN(n13606) );
  NAND2_X1 U15634 ( .A1(n13601), .A2(n13702), .ZN(n13603) );
  NAND2_X1 U15635 ( .A1(n13847), .A2(n13697), .ZN(n13602) );
  NAND2_X1 U15636 ( .A1(n13603), .A2(n13602), .ZN(n13604) );
  XNOR2_X1 U15637 ( .A(n13604), .B(n13705), .ZN(n13605) );
  XOR2_X1 U15638 ( .A(n13606), .B(n13605), .Z(n13760) );
  OAI22_X1 U15639 ( .A1(n14497), .A2(n13739), .B1(n14427), .B2(n13741), .ZN(
        n13608) );
  XNOR2_X1 U15640 ( .A(n13608), .B(n13705), .ZN(n13615) );
  NOR2_X1 U15641 ( .A1(n14427), .A2(n13740), .ZN(n13609) );
  AOI21_X1 U15642 ( .B1(n13610), .B2(n13697), .A(n13609), .ZN(n13616) );
  XNOR2_X1 U15643 ( .A(n13615), .B(n13616), .ZN(n13795) );
  NAND2_X1 U15644 ( .A1(n14436), .A2(n13702), .ZN(n13612) );
  OR2_X1 U15645 ( .A1(n13833), .A2(n13741), .ZN(n13611) );
  NAND2_X1 U15646 ( .A1(n13612), .A2(n13611), .ZN(n13613) );
  XNOR2_X1 U15647 ( .A(n13613), .B(n13705), .ZN(n13619) );
  NOR2_X1 U15648 ( .A1(n13833), .A2(n13740), .ZN(n13614) );
  AOI21_X1 U15649 ( .B1(n14436), .B2(n13697), .A(n13614), .ZN(n13620) );
  XNOR2_X1 U15650 ( .A(n13619), .B(n13620), .ZN(n14428) );
  INV_X1 U15651 ( .A(n13615), .ZN(n13617) );
  OR2_X1 U15652 ( .A1(n13617), .A2(n13616), .ZN(n14429) );
  INV_X1 U15653 ( .A(n13619), .ZN(n13621) );
  NAND2_X1 U15654 ( .A1(n13622), .A2(n13702), .ZN(n13624) );
  OR2_X1 U15655 ( .A1(n14441), .A2(n13741), .ZN(n13623) );
  NAND2_X1 U15656 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  XNOR2_X1 U15657 ( .A(n13625), .B(n13705), .ZN(n13626) );
  OAI22_X1 U15658 ( .A1(n14486), .A2(n13741), .B1(n14441), .B2(n13740), .ZN(
        n13830) );
  INV_X1 U15659 ( .A(n13626), .ZN(n13627) );
  NOR2_X1 U15660 ( .A1(n13628), .A2(n13627), .ZN(n14444) );
  OAI22_X1 U15661 ( .A1(n13631), .A2(n13739), .B1(n13629), .B2(n13741), .ZN(
        n13630) );
  XNOR2_X1 U15662 ( .A(n13630), .B(n13705), .ZN(n13635) );
  OR2_X1 U15663 ( .A1(n13631), .A2(n13741), .ZN(n13633) );
  NAND2_X1 U15664 ( .A1(n10343), .A2(n14458), .ZN(n13632) );
  NAND2_X1 U15665 ( .A1(n13633), .A2(n13632), .ZN(n13636) );
  XNOR2_X1 U15666 ( .A(n13635), .B(n13636), .ZN(n14443) );
  NOR2_X1 U15667 ( .A1(n14444), .A2(n14443), .ZN(n13634) );
  INV_X1 U15668 ( .A(n13635), .ZN(n13638) );
  INV_X1 U15669 ( .A(n13636), .ZN(n13637) );
  NAND2_X1 U15670 ( .A1(n13638), .A2(n13637), .ZN(n13639) );
  NAND2_X1 U15671 ( .A1(n14259), .A2(n13702), .ZN(n13641) );
  NAND2_X1 U15672 ( .A1(n14440), .A2(n13697), .ZN(n13640) );
  NAND2_X1 U15673 ( .A1(n13641), .A2(n13640), .ZN(n13642) );
  XNOR2_X1 U15674 ( .A(n13642), .B(n13705), .ZN(n13643) );
  AOI22_X1 U15675 ( .A1(n14259), .A2(n13697), .B1(n10343), .B2(n14440), .ZN(
        n13644) );
  XNOR2_X1 U15676 ( .A(n13643), .B(n13644), .ZN(n14454) );
  INV_X1 U15677 ( .A(n13643), .ZN(n13645) );
  NAND2_X1 U15678 ( .A1(n13645), .A2(n13644), .ZN(n13646) );
  NAND2_X1 U15679 ( .A1(n13647), .A2(n13646), .ZN(n13814) );
  OAI22_X1 U15680 ( .A1(n11599), .A2(n13741), .B1(n14135), .B2(n13740), .ZN(
        n13652) );
  NAND2_X1 U15681 ( .A1(n14254), .A2(n13702), .ZN(n13649) );
  NAND2_X1 U15682 ( .A1(n14456), .A2(n13697), .ZN(n13648) );
  NAND2_X1 U15683 ( .A1(n13649), .A2(n13648), .ZN(n13650) );
  XNOR2_X1 U15684 ( .A(n13650), .B(n13705), .ZN(n13651) );
  XOR2_X1 U15685 ( .A(n13652), .B(n13651), .Z(n13813) );
  INV_X1 U15686 ( .A(n13651), .ZN(n13654) );
  INV_X1 U15687 ( .A(n13652), .ZN(n13653) );
  NAND2_X1 U15688 ( .A1(n13654), .A2(n13653), .ZN(n13655) );
  OAI22_X1 U15689 ( .A1(n14143), .A2(n13739), .B1(n13816), .B2(n13741), .ZN(
        n13656) );
  XNOR2_X1 U15690 ( .A(n13656), .B(n13705), .ZN(n13659) );
  OAI22_X1 U15691 ( .A1(n14143), .A2(n13741), .B1(n13816), .B2(n13740), .ZN(
        n13658) );
  XNOR2_X1 U15692 ( .A(n13659), .B(n13658), .ZN(n13724) );
  NAND2_X1 U15693 ( .A1(n13659), .A2(n13658), .ZN(n13660) );
  NAND2_X1 U15694 ( .A1(n13726), .A2(n13660), .ZN(n13788) );
  OAI22_X1 U15695 ( .A1(n14124), .A2(n13739), .B1(n14137), .B2(n13741), .ZN(
        n13661) );
  XNOR2_X1 U15696 ( .A(n13661), .B(n13705), .ZN(n13665) );
  AND2_X1 U15697 ( .A1(n14103), .A2(n10343), .ZN(n13662) );
  AOI21_X1 U15698 ( .B1(n14244), .B2(n13697), .A(n13662), .ZN(n13663) );
  XNOR2_X1 U15699 ( .A(n13665), .B(n13663), .ZN(n13787) );
  NAND2_X1 U15700 ( .A1(n13788), .A2(n13787), .ZN(n13786) );
  INV_X1 U15701 ( .A(n13663), .ZN(n13664) );
  NAND2_X1 U15702 ( .A1(n13665), .A2(n13664), .ZN(n13666) );
  AOI22_X1 U15703 ( .A1(n14236), .A2(n13702), .B1(n13697), .B2(n13844), .ZN(
        n13667) );
  XNOR2_X1 U15704 ( .A(n13667), .B(n13705), .ZN(n13670) );
  AOI22_X1 U15705 ( .A1(n14236), .A2(n13697), .B1(n10343), .B2(n13844), .ZN(
        n13669) );
  XNOR2_X1 U15706 ( .A(n13670), .B(n13669), .ZN(n13754) );
  INV_X1 U15707 ( .A(n13754), .ZN(n13668) );
  NAND2_X1 U15708 ( .A1(n13670), .A2(n13669), .ZN(n13671) );
  OAI22_X1 U15709 ( .A1(n14090), .A2(n13741), .B1(n13718), .B2(n13740), .ZN(
        n13676) );
  NAND2_X1 U15710 ( .A1(n14228), .A2(n13702), .ZN(n13673) );
  NAND2_X1 U15711 ( .A1(n14105), .A2(n13697), .ZN(n13672) );
  NAND2_X1 U15712 ( .A1(n13673), .A2(n13672), .ZN(n13674) );
  XNOR2_X1 U15713 ( .A(n13674), .B(n13705), .ZN(n13675) );
  XOR2_X1 U15714 ( .A(n13676), .B(n13675), .Z(n13805) );
  INV_X1 U15715 ( .A(n13675), .ZN(n13678) );
  INV_X1 U15716 ( .A(n13676), .ZN(n13677) );
  NAND2_X1 U15717 ( .A1(n13678), .A2(n13677), .ZN(n13679) );
  NAND2_X1 U15718 ( .A1(n14074), .A2(n13702), .ZN(n13681) );
  NAND2_X1 U15719 ( .A1(n13843), .A2(n13697), .ZN(n13680) );
  NAND2_X1 U15720 ( .A1(n13681), .A2(n13680), .ZN(n13682) );
  XNOR2_X1 U15721 ( .A(n13682), .B(n13705), .ZN(n13683) );
  AOI22_X1 U15722 ( .A1(n14074), .A2(n13697), .B1(n10343), .B2(n13843), .ZN(
        n13684) );
  XNOR2_X1 U15723 ( .A(n13683), .B(n13684), .ZN(n13717) );
  INV_X1 U15724 ( .A(n13683), .ZN(n13685) );
  NAND2_X1 U15725 ( .A1(n14216), .A2(n13702), .ZN(n13687) );
  NAND2_X1 U15726 ( .A1(n13842), .A2(n13697), .ZN(n13686) );
  NAND2_X1 U15727 ( .A1(n13687), .A2(n13686), .ZN(n13688) );
  XNOR2_X1 U15728 ( .A(n13688), .B(n13705), .ZN(n13689) );
  AOI22_X1 U15729 ( .A1(n14216), .A2(n13697), .B1(n10343), .B2(n13842), .ZN(
        n13690) );
  XNOR2_X1 U15730 ( .A(n13689), .B(n13690), .ZN(n13779) );
  NAND2_X1 U15731 ( .A1(n13778), .A2(n13779), .ZN(n13693) );
  INV_X1 U15732 ( .A(n13689), .ZN(n13691) );
  NAND2_X1 U15733 ( .A1(n13691), .A2(n13690), .ZN(n13692) );
  NAND2_X1 U15734 ( .A1(n13693), .A2(n13692), .ZN(n13770) );
  NAND2_X1 U15735 ( .A1(n14209), .A2(n13702), .ZN(n13695) );
  NAND2_X1 U15736 ( .A1(n13841), .A2(n13697), .ZN(n13694) );
  NAND2_X1 U15737 ( .A1(n13695), .A2(n13694), .ZN(n13696) );
  XNOR2_X1 U15738 ( .A(n13696), .B(n13705), .ZN(n13698) );
  AOI22_X1 U15739 ( .A1(n14209), .A2(n13697), .B1(n10343), .B2(n13841), .ZN(
        n13699) );
  XNOR2_X1 U15740 ( .A(n13698), .B(n13699), .ZN(n13771) );
  INV_X1 U15741 ( .A(n13698), .ZN(n13700) );
  NAND2_X1 U15742 ( .A1(n13700), .A2(n13699), .ZN(n13701) );
  OAI22_X1 U15743 ( .A1(n14031), .A2(n13741), .B1(n13772), .B2(n13740), .ZN(
        n13708) );
  NAND2_X1 U15744 ( .A1(n14201), .A2(n13702), .ZN(n13704) );
  NAND2_X1 U15745 ( .A1(n14004), .A2(n13697), .ZN(n13703) );
  NAND2_X1 U15746 ( .A1(n13704), .A2(n13703), .ZN(n13706) );
  XNOR2_X1 U15747 ( .A(n13706), .B(n13705), .ZN(n13707) );
  XOR2_X1 U15748 ( .A(n13708), .B(n13707), .Z(n13822) );
  INV_X1 U15749 ( .A(n13707), .ZN(n13710) );
  INV_X1 U15750 ( .A(n13708), .ZN(n13709) );
  XOR2_X1 U15751 ( .A(n13737), .B(n13738), .Z(n13715) );
  AOI22_X1 U15752 ( .A1(n14459), .A2(n14004), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13712) );
  NAND2_X1 U15753 ( .A1(n14457), .A2(n14003), .ZN(n13711) );
  OAI211_X1 U15754 ( .C1(n14485), .C2(n14013), .A(n13712), .B(n13711), .ZN(
        n13713) );
  AOI21_X1 U15755 ( .B1(n14195), .B2(n14481), .A(n13713), .ZN(n13714) );
  OAI21_X1 U15756 ( .B1(n13715), .B2(n14476), .A(n13714), .ZN(P1_U3214) );
  XOR2_X1 U15757 ( .A(n13717), .B(n13716), .Z(n13723) );
  INV_X1 U15758 ( .A(n14075), .ZN(n13720) );
  OAI22_X1 U15759 ( .A1(n13718), .A2(n14136), .B1(n13773), .B2(n14138), .ZN(
        n14221) );
  AOI22_X1 U15760 ( .A1(n14221), .A2(n13825), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13719) );
  OAI21_X1 U15761 ( .B1(n13720), .B2(n14485), .A(n13719), .ZN(n13721) );
  AOI21_X1 U15762 ( .B1(n14074), .B2(n14481), .A(n13721), .ZN(n13722) );
  OAI21_X1 U15763 ( .B1(n13723), .B2(n14476), .A(n13722), .ZN(P1_U3216) );
  AOI21_X1 U15764 ( .B1(n13725), .B2(n13724), .A(n14476), .ZN(n13727) );
  NAND2_X1 U15765 ( .A1(n13727), .A2(n13726), .ZN(n13732) );
  NAND2_X1 U15766 ( .A1(n14459), .A2(n14456), .ZN(n13728) );
  OAI211_X1 U15767 ( .C1(n14471), .C2(n14137), .A(n13729), .B(n13728), .ZN(
        n13730) );
  AOI21_X1 U15768 ( .B1(n14141), .B2(n13835), .A(n13730), .ZN(n13731) );
  OAI211_X1 U15769 ( .C1(n14143), .C2(n14461), .A(n13732), .B(n13731), .ZN(
        P1_U3219) );
  INV_X1 U15770 ( .A(n13733), .ZN(n13736) );
  INV_X1 U15771 ( .A(n13734), .ZN(n13735) );
  INV_X1 U15772 ( .A(n14003), .ZN(n13994) );
  OAI22_X1 U15773 ( .A1(n14189), .A2(n13739), .B1(n13994), .B2(n13741), .ZN(
        n13744) );
  OAI22_X1 U15774 ( .A1(n14189), .A2(n13741), .B1(n13994), .B2(n13740), .ZN(
        n13742) );
  XNOR2_X1 U15775 ( .A(n13742), .B(n13705), .ZN(n13743) );
  XOR2_X1 U15776 ( .A(n13744), .B(n13743), .Z(n13745) );
  AOI22_X1 U15777 ( .A1(n14459), .A2(n13840), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13747) );
  NAND2_X1 U15778 ( .A1(n14457), .A2(n13839), .ZN(n13746) );
  OAI211_X1 U15779 ( .C1(n14485), .C2(n13748), .A(n13747), .B(n13746), .ZN(
        n13749) );
  AOI21_X1 U15780 ( .B1(n13982), .B2(n14481), .A(n13749), .ZN(n13750) );
  INV_X1 U15781 ( .A(n13751), .ZN(n13752) );
  AOI21_X1 U15782 ( .B1(n13754), .B2(n13753), .A(n13752), .ZN(n13759) );
  AOI22_X1 U15783 ( .A1(n14457), .A2(n14105), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13756) );
  NAND2_X1 U15784 ( .A1(n14459), .A2(n14103), .ZN(n13755) );
  OAI211_X1 U15785 ( .C1(n14485), .C2(n14107), .A(n13756), .B(n13755), .ZN(
        n13757) );
  AOI21_X1 U15786 ( .B1(n14236), .B2(n14481), .A(n13757), .ZN(n13758) );
  OAI21_X1 U15787 ( .B1(n13759), .B2(n14476), .A(n13758), .ZN(P1_U3223) );
  AOI21_X1 U15788 ( .B1(n13761), .B2(n13760), .A(n14476), .ZN(n13763) );
  NAND2_X1 U15789 ( .A1(n13763), .A2(n13762), .ZN(n13769) );
  NOR2_X1 U15790 ( .A1(n14485), .A2(n13764), .ZN(n13767) );
  OAI22_X1 U15791 ( .A1(n14471), .A2(n14427), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13765), .ZN(n13766) );
  AOI211_X1 U15792 ( .C1(n14459), .C2(n13848), .A(n13767), .B(n13766), .ZN(
        n13768) );
  OAI211_X1 U15793 ( .C1(n7016), .C2(n14461), .A(n13769), .B(n13768), .ZN(
        P1_U3224) );
  XOR2_X1 U15794 ( .A(n13771), .B(n13770), .Z(n13777) );
  OAI22_X1 U15795 ( .A1(n13773), .A2(n14136), .B1(n13772), .B2(n14138), .ZN(
        n14208) );
  AOI22_X1 U15796 ( .A1(n13825), .A2(n14208), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13774) );
  OAI21_X1 U15797 ( .B1(n14038), .B2(n14485), .A(n13774), .ZN(n13775) );
  AOI21_X1 U15798 ( .B1(n14209), .B2(n14481), .A(n13775), .ZN(n13776) );
  OAI21_X1 U15799 ( .B1(n13777), .B2(n14476), .A(n13776), .ZN(P1_U3225) );
  XOR2_X1 U15800 ( .A(n13779), .B(n13778), .Z(n13785) );
  NAND2_X1 U15801 ( .A1(n13843), .A2(n14154), .ZN(n13781) );
  NAND2_X1 U15802 ( .A1(n13841), .A2(n14152), .ZN(n13780) );
  NAND2_X1 U15803 ( .A1(n13781), .A2(n13780), .ZN(n14056) );
  AOI22_X1 U15804 ( .A1(n14056), .A2(n13825), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13782) );
  OAI21_X1 U15805 ( .B1(n14059), .B2(n14485), .A(n13782), .ZN(n13783) );
  AOI21_X1 U15806 ( .B1(n14216), .B2(n14481), .A(n13783), .ZN(n13784) );
  OAI21_X1 U15807 ( .B1(n13785), .B2(n14476), .A(n13784), .ZN(P1_U3229) );
  OAI211_X1 U15808 ( .C1(n13788), .C2(n13787), .A(n13786), .B(n14464), .ZN(
        n13794) );
  NAND2_X1 U15809 ( .A1(n13844), .A2(n14152), .ZN(n13790) );
  OR2_X1 U15810 ( .A1(n13816), .A2(n14136), .ZN(n13789) );
  AND2_X1 U15811 ( .A1(n13790), .A2(n13789), .ZN(n14120) );
  OAI22_X1 U15812 ( .A1(n14120), .A2(n13808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13791), .ZN(n13792) );
  AOI21_X1 U15813 ( .B1(n14122), .B2(n13835), .A(n13792), .ZN(n13793) );
  OAI211_X1 U15814 ( .C1(n14124), .C2(n14461), .A(n13794), .B(n13793), .ZN(
        P1_U3233) );
  OAI211_X1 U15815 ( .C1(n13796), .C2(n13795), .A(n14430), .B(n14464), .ZN(
        n13802) );
  NOR2_X1 U15816 ( .A1(n14485), .A2(n13797), .ZN(n13800) );
  OAI21_X1 U15817 ( .B1(n14471), .B2(n13833), .A(n13798), .ZN(n13799) );
  AOI211_X1 U15818 ( .C1(n14459), .C2(n13847), .A(n13800), .B(n13799), .ZN(
        n13801) );
  OAI211_X1 U15819 ( .C1(n14497), .C2(n14461), .A(n13802), .B(n13801), .ZN(
        P1_U3234) );
  OAI21_X1 U15820 ( .B1(n13805), .B2(n13804), .A(n13803), .ZN(n13806) );
  NAND2_X1 U15821 ( .A1(n13806), .A2(n14464), .ZN(n13812) );
  INV_X1 U15822 ( .A(n14089), .ZN(n13810) );
  AND2_X1 U15823 ( .A1(n13844), .A2(n14154), .ZN(n13807) );
  AOI21_X1 U15824 ( .B1(n13843), .B2(n14152), .A(n13807), .ZN(n14230) );
  INV_X1 U15825 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15230) );
  OAI22_X1 U15826 ( .A1(n14230), .A2(n13808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15230), .ZN(n13809) );
  AOI21_X1 U15827 ( .B1(n13810), .B2(n13835), .A(n13809), .ZN(n13811) );
  OAI211_X1 U15828 ( .C1(n14461), .C2(n14090), .A(n13812), .B(n13811), .ZN(
        P1_U3235) );
  XOR2_X1 U15829 ( .A(n13814), .B(n13813), .Z(n13820) );
  NOR2_X1 U15830 ( .A1(n14485), .A2(n14156), .ZN(n13818) );
  NAND2_X1 U15831 ( .A1(n14459), .A2(n14440), .ZN(n13815) );
  NAND2_X1 U15832 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14573)
         );
  OAI211_X1 U15833 ( .C1(n14471), .C2(n13816), .A(n13815), .B(n14573), .ZN(
        n13817) );
  AOI211_X1 U15834 ( .C1(n14254), .C2(n14481), .A(n13818), .B(n13817), .ZN(
        n13819) );
  OAI21_X1 U15835 ( .B1(n13820), .B2(n14476), .A(n13819), .ZN(P1_U3238) );
  XOR2_X1 U15836 ( .A(n13822), .B(n13821), .Z(n13829) );
  NAND2_X1 U15837 ( .A1(n13841), .A2(n14154), .ZN(n13824) );
  NAND2_X1 U15838 ( .A1(n13840), .A2(n14152), .ZN(n13823) );
  NAND2_X1 U15839 ( .A1(n13824), .A2(n13823), .ZN(n14024) );
  AOI22_X1 U15840 ( .A1(n13825), .A2(n14024), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13826) );
  OAI21_X1 U15841 ( .B1(n14026), .B2(n14485), .A(n13826), .ZN(n13827) );
  AOI21_X1 U15842 ( .B1(n14201), .B2(n14481), .A(n13827), .ZN(n13828) );
  OAI21_X1 U15843 ( .B1(n13829), .B2(n14476), .A(n13828), .ZN(P1_U3240) );
  OAI211_X1 U15844 ( .C1(n13831), .C2(n13830), .A(n14442), .B(n14464), .ZN(
        n13838) );
  AOI22_X1 U15845 ( .A1(n14457), .A2(n14458), .B1(P1_REG3_REG_15__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13832) );
  OAI21_X1 U15846 ( .B1(n13833), .B2(n14470), .A(n13832), .ZN(n13834) );
  AOI21_X1 U15847 ( .B1(n13836), .B2(n13835), .A(n13834), .ZN(n13837) );
  OAI211_X1 U15848 ( .C1(n14486), .C2(n14461), .A(n13838), .B(n13837), .ZN(
        P1_U3241) );
  MUX2_X1 U15849 ( .A(n13987), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13856), .Z(
        P1_U3590) );
  MUX2_X1 U15850 ( .A(n13839), .B(P1_DATAO_REG_29__SCAN_IN), .S(n13856), .Z(
        P1_U3589) );
  MUX2_X1 U15851 ( .A(n14003), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13856), .Z(
        P1_U3588) );
  MUX2_X1 U15852 ( .A(n13840), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13856), .Z(
        P1_U3587) );
  MUX2_X1 U15853 ( .A(n14004), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13856), .Z(
        P1_U3586) );
  MUX2_X1 U15854 ( .A(n13841), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13856), .Z(
        P1_U3585) );
  MUX2_X1 U15855 ( .A(n13842), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13856), .Z(
        P1_U3584) );
  MUX2_X1 U15856 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13843), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15857 ( .A(n14105), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13856), .Z(
        P1_U3582) );
  MUX2_X1 U15858 ( .A(n13844), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13856), .Z(
        P1_U3581) );
  MUX2_X1 U15859 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14103), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15860 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14153), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15861 ( .A(n14456), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13856), .Z(
        P1_U3578) );
  MUX2_X1 U15862 ( .A(n14440), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13856), .Z(
        P1_U3577) );
  MUX2_X1 U15863 ( .A(n14458), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13856), .Z(
        P1_U3576) );
  MUX2_X1 U15864 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13845), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15865 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n6793), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15866 ( .A(n13846), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13856), .Z(
        P1_U3573) );
  MUX2_X1 U15867 ( .A(n13847), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13856), .Z(
        P1_U3572) );
  MUX2_X1 U15868 ( .A(n13848), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13856), .Z(
        P1_U3571) );
  MUX2_X1 U15869 ( .A(n13849), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13856), .Z(
        P1_U3570) );
  MUX2_X1 U15870 ( .A(n13850), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13856), .Z(
        P1_U3569) );
  MUX2_X1 U15871 ( .A(n13851), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13856), .Z(
        P1_U3568) );
  MUX2_X1 U15872 ( .A(n13852), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13856), .Z(
        P1_U3567) );
  MUX2_X1 U15873 ( .A(n13853), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13856), .Z(
        P1_U3566) );
  MUX2_X1 U15874 ( .A(n13854), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13856), .Z(
        P1_U3565) );
  MUX2_X1 U15875 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13855), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15876 ( .A(n13857), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13856), .Z(
        P1_U3563) );
  MUX2_X1 U15877 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13858), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15878 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13859), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15879 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13860), .S(P1_U4016), .Z(
        P1_U3560) );
  MUX2_X1 U15880 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n15154), .S(n13867), .Z(
        n13861) );
  OAI21_X1 U15881 ( .B1(n9594), .B2(n13862), .A(n13861), .ZN(n13863) );
  NAND3_X1 U15882 ( .A1(n14566), .A2(n13864), .A3(n13863), .ZN(n13872) );
  OAI211_X1 U15883 ( .C1(n13877), .C2(n13866), .A(n14563), .B(n13865), .ZN(
        n13871) );
  INV_X1 U15884 ( .A(n13867), .ZN(n13868) );
  NAND2_X1 U15885 ( .A1(n13963), .A2(n13868), .ZN(n13870) );
  AOI22_X1 U15886 ( .A1(n14544), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13869) );
  NAND4_X1 U15887 ( .A1(n13872), .A2(n13871), .A3(n13870), .A4(n13869), .ZN(
        P1_U3244) );
  NOR2_X1 U15888 ( .A1(n6530), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13874) );
  NOR2_X1 U15889 ( .A1(n13874), .A2(n13873), .ZN(n14541) );
  INV_X1 U15890 ( .A(n13875), .ZN(n13876) );
  MUX2_X1 U15891 ( .A(n13877), .B(n13876), .S(n6530), .Z(n13879) );
  NAND2_X1 U15892 ( .A1(n13879), .A2(n13878), .ZN(n13880) );
  OAI211_X1 U15893 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14541), .A(n13880), .B(
        P1_U4016), .ZN(n13925) );
  AOI22_X1 U15894 ( .A1(n14544), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13891) );
  OAI21_X1 U15895 ( .B1(n13882), .B2(n13881), .A(n13899), .ZN(n13883) );
  OAI22_X1 U15896 ( .A1(n13884), .A2(n14571), .B1(n14552), .B2(n13883), .ZN(
        n13885) );
  INV_X1 U15897 ( .A(n13885), .ZN(n13890) );
  OAI21_X1 U15898 ( .B1(n13887), .B2(n13886), .A(n13894), .ZN(n13888) );
  OR2_X1 U15899 ( .A1(n14557), .A2(n13888), .ZN(n13889) );
  NAND4_X1 U15900 ( .A1(n13925), .A2(n13891), .A3(n13890), .A4(n13889), .ZN(
        P1_U3245) );
  MUX2_X1 U15901 ( .A(n9415), .B(P1_REG1_REG_3__SCAN_IN), .S(n13896), .Z(
        n13892) );
  NAND3_X1 U15902 ( .A1(n13894), .A2(n13893), .A3(n13892), .ZN(n13895) );
  NAND3_X1 U15903 ( .A1(n14566), .A2(n13910), .A3(n13895), .ZN(n13905) );
  NAND2_X1 U15904 ( .A1(n13963), .A2(n13896), .ZN(n13904) );
  MUX2_X1 U15905 ( .A(n10384), .B(P1_REG2_REG_3__SCAN_IN), .S(n13896), .Z(
        n13897) );
  NAND3_X1 U15906 ( .A1(n13899), .A2(n13898), .A3(n13897), .ZN(n13900) );
  NAND3_X1 U15907 ( .A1(n14563), .A2(n13919), .A3(n13900), .ZN(n13903) );
  AOI21_X1 U15908 ( .B1(n14544), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n13901), .ZN(
        n13902) );
  NAND4_X1 U15909 ( .A1(n13905), .A2(n13904), .A3(n13903), .A4(n13902), .ZN(
        P1_U3246) );
  INV_X1 U15910 ( .A(n13906), .ZN(n13907) );
  AOI21_X1 U15911 ( .B1(n14544), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n13907), .ZN(
        n13924) );
  MUX2_X1 U15912 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9418), .S(n13914), .Z(
        n13908) );
  NAND3_X1 U15913 ( .A1(n13910), .A2(n13909), .A3(n13908), .ZN(n13911) );
  NAND2_X1 U15914 ( .A1(n13912), .A2(n13911), .ZN(n13913) );
  OAI22_X1 U15915 ( .A1(n13914), .A2(n14571), .B1(n14557), .B2(n13913), .ZN(
        n13915) );
  INV_X1 U15916 ( .A(n13915), .ZN(n13923) );
  INV_X1 U15917 ( .A(n13916), .ZN(n13921) );
  NAND3_X1 U15918 ( .A1(n13919), .A2(n13918), .A3(n13917), .ZN(n13920) );
  NAND3_X1 U15919 ( .A1(n14563), .A2(n13921), .A3(n13920), .ZN(n13922) );
  NAND4_X1 U15920 ( .A1(n13925), .A2(n13924), .A3(n13923), .A4(n13922), .ZN(
        P1_U3247) );
  OAI21_X1 U15921 ( .B1(n14575), .B2(n13927), .A(n13926), .ZN(n13928) );
  AOI21_X1 U15922 ( .B1(n13929), .B2(n13963), .A(n13928), .ZN(n13942) );
  NAND2_X1 U15923 ( .A1(n13931), .A2(n13930), .ZN(n13932) );
  NAND3_X1 U15924 ( .A1(n14566), .A2(n13933), .A3(n13932), .ZN(n13941) );
  INV_X1 U15925 ( .A(n13934), .ZN(n13939) );
  NAND3_X1 U15926 ( .A1(n13937), .A2(n13936), .A3(n13935), .ZN(n13938) );
  NAND3_X1 U15927 ( .A1(n14563), .A2(n13939), .A3(n13938), .ZN(n13940) );
  NAND3_X1 U15928 ( .A1(n13942), .A2(n13941), .A3(n13940), .ZN(P1_U3249) );
  OR3_X1 U15929 ( .A1(n13945), .A2(n13944), .A3(n13943), .ZN(n13946) );
  NAND3_X1 U15930 ( .A1(n13947), .A2(n14563), .A3(n13946), .ZN(n13957) );
  INV_X1 U15931 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n13948) );
  NAND2_X1 U15932 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14482)
         );
  OAI21_X1 U15933 ( .B1(n14575), .B2(n13948), .A(n14482), .ZN(n13949) );
  AOI21_X1 U15934 ( .B1(n13963), .B2(n13950), .A(n13949), .ZN(n13956) );
  OAI21_X1 U15935 ( .B1(n13953), .B2(n13952), .A(n13951), .ZN(n13954) );
  NAND2_X1 U15936 ( .A1(n13954), .A2(n14566), .ZN(n13955) );
  NAND3_X1 U15937 ( .A1(n13957), .A2(n13956), .A3(n13955), .ZN(P1_U3254) );
  NAND2_X1 U15938 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14451)
         );
  AOI211_X1 U15939 ( .C1(n13960), .C2(n13959), .A(n14557), .B(n13958), .ZN(
        n13961) );
  INV_X1 U15940 ( .A(n13961), .ZN(n13962) );
  AND2_X1 U15941 ( .A1(n14451), .A2(n13962), .ZN(n13972) );
  AOI22_X1 U15942 ( .A1(n13963), .A2(n13966), .B1(n14544), .B2(
        P1_ADDR_REG_16__SCAN_IN), .ZN(n13971) );
  NAND2_X1 U15943 ( .A1(n13966), .A2(n13964), .ZN(n13965) );
  OAI21_X1 U15944 ( .B1(n13966), .B2(n13964), .A(n13965), .ZN(n13968) );
  OAI211_X1 U15945 ( .C1(n13969), .C2(n13968), .A(n13967), .B(n14563), .ZN(
        n13970) );
  NAND3_X1 U15946 ( .A1(n13972), .A2(n13971), .A3(n13970), .ZN(P1_U3259) );
  NAND2_X1 U15947 ( .A1(n14169), .A2(n14167), .ZN(n13977) );
  INV_X1 U15948 ( .A(P1_B_REG_SCAN_IN), .ZN(n13973) );
  NOR2_X1 U15949 ( .A1(n6530), .A2(n13973), .ZN(n13974) );
  NOR2_X1 U15950 ( .A1(n14138), .A2(n13974), .ZN(n13986) );
  NAND2_X1 U15951 ( .A1(n13975), .A2(n13986), .ZN(n14173) );
  NOR2_X1 U15952 ( .A1(n14159), .A2(n14173), .ZN(n13979) );
  AOI21_X1 U15953 ( .B1(n14159), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13979), 
        .ZN(n13976) );
  OAI211_X1 U15954 ( .C1(n14171), .C2(n14161), .A(n13977), .B(n13976), .ZN(
        P1_U3263) );
  XNOR2_X1 U15955 ( .A(n13983), .B(n13978), .ZN(n14172) );
  NAND2_X1 U15956 ( .A1(n14172), .A2(n14167), .ZN(n13981) );
  AOI21_X1 U15957 ( .B1(n14159), .B2(P1_REG2_REG_30__SCAN_IN), .A(n13979), 
        .ZN(n13980) );
  OAI211_X1 U15958 ( .C1(n14175), .C2(n14161), .A(n13981), .B(n13980), .ZN(
        P1_U3264) );
  AOI21_X1 U15959 ( .B1(n13985), .B2(n13984), .A(n13983), .ZN(n14181) );
  INV_X1 U15960 ( .A(n13985), .ZN(n14179) );
  NAND2_X1 U15961 ( .A1(n13987), .A2(n13986), .ZN(n14178) );
  OAI22_X1 U15962 ( .A1(n13989), .A2(n14178), .B1(n13988), .B2(n14106), .ZN(
        n13991) );
  NAND2_X1 U15963 ( .A1(n14003), .A2(n14154), .ZN(n14177) );
  NOR2_X1 U15964 ( .A1(n14159), .A2(n14177), .ZN(n13990) );
  AOI211_X1 U15965 ( .C1(n14159), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13991), 
        .B(n13990), .ZN(n13992) );
  OAI21_X1 U15966 ( .B1(n14179), .B2(n14161), .A(n13992), .ZN(n13993) );
  AOI21_X1 U15967 ( .B1(n14181), .B2(n14167), .A(n13993), .ZN(n14000) );
  NAND2_X1 U15968 ( .A1(n13996), .A2(n13995), .ZN(n13998) );
  XNOR2_X1 U15969 ( .A(n13998), .B(n13997), .ZN(n14176) );
  NAND2_X1 U15970 ( .A1(n14176), .A2(n14114), .ZN(n13999) );
  OAI211_X1 U15971 ( .C1(n14183), .C2(n14116), .A(n14000), .B(n13999), .ZN(
        P1_U3356) );
  AOI21_X1 U15972 ( .B1(n14005), .B2(n14002), .A(n14001), .ZN(n14198) );
  AOI22_X1 U15973 ( .A1(n14154), .A2(n14004), .B1(n14003), .B2(n14152), .ZN(
        n14009) );
  XNOR2_X1 U15974 ( .A(n14006), .B(n14005), .ZN(n14007) );
  NAND2_X1 U15975 ( .A1(n14007), .A2(n14264), .ZN(n14008) );
  OAI211_X1 U15976 ( .C1(n14198), .C2(n14010), .A(n14009), .B(n14008), .ZN(
        n14200) );
  NAND2_X1 U15977 ( .A1(n14200), .A2(n14076), .ZN(n14018) );
  AOI21_X1 U15978 ( .B1(n14195), .B2(n14029), .A(n14011), .ZN(n14196) );
  NOR2_X1 U15979 ( .A1(n14012), .A2(n14161), .ZN(n14016) );
  OAI22_X1 U15980 ( .A1(n14076), .A2(n14014), .B1(n14013), .B2(n14106), .ZN(
        n14015) );
  AOI211_X1 U15981 ( .C1(n14196), .C2(n14167), .A(n14016), .B(n14015), .ZN(
        n14017) );
  OAI211_X1 U15982 ( .C1(n14198), .C2(n14019), .A(n14018), .B(n14017), .ZN(
        P1_U3266) );
  XNOR2_X1 U15983 ( .A(n14021), .B(n14020), .ZN(n14205) );
  XNOR2_X1 U15984 ( .A(n14023), .B(n14022), .ZN(n14025) );
  AOI21_X1 U15985 ( .B1(n14025), .B2(n14264), .A(n14024), .ZN(n14204) );
  OAI21_X1 U15986 ( .B1(n14026), .B2(n14106), .A(n14204), .ZN(n14027) );
  NAND2_X1 U15987 ( .A1(n14027), .A2(n14076), .ZN(n14034) );
  NAND2_X1 U15988 ( .A1(n14037), .A2(n14201), .ZN(n14028) );
  AND2_X1 U15989 ( .A1(n14029), .A2(n14028), .ZN(n14202) );
  INV_X1 U15990 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14030) );
  OAI22_X1 U15991 ( .A1(n14031), .A2(n14161), .B1(n14030), .B2(n14076), .ZN(
        n14032) );
  AOI21_X1 U15992 ( .B1(n14202), .B2(n14167), .A(n14032), .ZN(n14033) );
  OAI211_X1 U15993 ( .C1(n14205), .C2(n14164), .A(n14034), .B(n14033), .ZN(
        P1_U3267) );
  AOI21_X1 U15994 ( .B1(n14036), .B2(n14035), .A(n6615), .ZN(n14213) );
  OAI21_X1 U15995 ( .B1(n6547), .B2(n14042), .A(n14037), .ZN(n14206) );
  INV_X1 U15996 ( .A(n14206), .ZN(n14044) );
  INV_X1 U15997 ( .A(n14208), .ZN(n14039) );
  OAI22_X1 U15998 ( .A1(n14159), .A2(n14039), .B1(n14038), .B2(n14106), .ZN(
        n14040) );
  AOI21_X1 U15999 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n14159), .A(n14040), 
        .ZN(n14041) );
  OAI21_X1 U16000 ( .B1(n14042), .B2(n14161), .A(n14041), .ZN(n14043) );
  AOI21_X1 U16001 ( .B1(n14044), .B2(n14167), .A(n14043), .ZN(n14049) );
  AOI21_X1 U16002 ( .B1(n14047), .B2(n14046), .A(n14045), .ZN(n14210) );
  NAND2_X1 U16003 ( .A1(n14210), .A2(n14114), .ZN(n14048) );
  OAI211_X1 U16004 ( .C1(n14213), .C2(n14116), .A(n14049), .B(n14048), .ZN(
        P1_U3268) );
  OAI21_X1 U16005 ( .B1(n14051), .B2(n6727), .A(n6836), .ZN(n14214) );
  OAI211_X1 U16006 ( .C1(n6651), .C2(n14053), .A(n14052), .B(n14264), .ZN(
        n14054) );
  INV_X1 U16007 ( .A(n14054), .ZN(n14055) );
  AOI211_X1 U16008 ( .C1(n14057), .C2(n14214), .A(n14056), .B(n14055), .ZN(
        n14218) );
  AOI211_X1 U16009 ( .C1(n14216), .C2(n14071), .A(n9590), .B(n6547), .ZN(
        n14215) );
  INV_X1 U16010 ( .A(n14216), .ZN(n14058) );
  NOR2_X1 U16011 ( .A1(n14058), .A2(n14161), .ZN(n14062) );
  OAI22_X1 U16012 ( .A1(n14076), .A2(n14060), .B1(n14059), .B2(n14106), .ZN(
        n14061) );
  AOI211_X1 U16013 ( .C1(n14215), .C2(n14063), .A(n14062), .B(n14061), .ZN(
        n14066) );
  NAND2_X1 U16014 ( .A1(n14214), .A2(n14064), .ZN(n14065) );
  OAI211_X1 U16015 ( .C1(n14218), .C2(n14159), .A(n14066), .B(n14065), .ZN(
        P1_U3269) );
  AOI21_X1 U16016 ( .B1(n14069), .B2(n14068), .A(n14067), .ZN(n14227) );
  INV_X1 U16017 ( .A(n14070), .ZN(n14073) );
  INV_X1 U16018 ( .A(n14071), .ZN(n14072) );
  AOI21_X1 U16019 ( .B1(n14074), .B2(n14073), .A(n14072), .ZN(n14223) );
  AOI22_X1 U16020 ( .A1(n14221), .A2(n14076), .B1(n14075), .B2(n14157), .ZN(
        n14078) );
  NAND2_X1 U16021 ( .A1(n14159), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14077) );
  OAI211_X1 U16022 ( .C1(n11600), .C2(n14161), .A(n14078), .B(n14077), .ZN(
        n14079) );
  AOI21_X1 U16023 ( .B1(n14223), .B2(n14167), .A(n14079), .ZN(n14084) );
  AOI21_X1 U16024 ( .B1(n14082), .B2(n14081), .A(n14080), .ZN(n14224) );
  NAND2_X1 U16025 ( .A1(n14224), .A2(n14114), .ZN(n14083) );
  OAI211_X1 U16026 ( .C1(n14227), .C2(n14116), .A(n14084), .B(n14083), .ZN(
        P1_U3270) );
  XNOR2_X1 U16027 ( .A(n14085), .B(n14087), .ZN(n14235) );
  OAI21_X1 U16028 ( .B1(n14088), .B2(n14087), .A(n14086), .ZN(n14233) );
  XNOR2_X1 U16029 ( .A(n14228), .B(n14099), .ZN(n14231) );
  OAI22_X1 U16030 ( .A1(n14230), .A2(n14159), .B1(n14089), .B2(n14106), .ZN(
        n14092) );
  NOR2_X1 U16031 ( .A1(n14090), .A2(n14161), .ZN(n14091) );
  AOI211_X1 U16032 ( .C1(n14159), .C2(P1_REG2_REG_22__SCAN_IN), .A(n14092), 
        .B(n14091), .ZN(n14093) );
  OAI21_X1 U16033 ( .B1(n14231), .B2(n14112), .A(n14093), .ZN(n14094) );
  AOI21_X1 U16034 ( .B1(n14233), .B2(n14114), .A(n14094), .ZN(n14095) );
  OAI21_X1 U16035 ( .B1(n14235), .B2(n14116), .A(n14095), .ZN(P1_U3271) );
  XNOR2_X1 U16036 ( .A(n14096), .B(n14097), .ZN(n14243) );
  XNOR2_X1 U16037 ( .A(n14098), .B(n14097), .ZN(n14241) );
  OAI21_X1 U16038 ( .B1(n14101), .B2(n14100), .A(n14099), .ZN(n14239) );
  NOR2_X1 U16039 ( .A1(n14076), .A2(n14102), .ZN(n14109) );
  AND2_X1 U16040 ( .A1(n14103), .A2(n14154), .ZN(n14104) );
  AOI21_X1 U16041 ( .B1(n14105), .B2(n14152), .A(n14104), .ZN(n14238) );
  OAI22_X1 U16042 ( .A1(n14238), .A2(n14159), .B1(n14107), .B2(n14106), .ZN(
        n14108) );
  AOI211_X1 U16043 ( .C1(n14236), .C2(n14110), .A(n14109), .B(n14108), .ZN(
        n14111) );
  OAI21_X1 U16044 ( .B1(n14239), .B2(n14112), .A(n14111), .ZN(n14113) );
  AOI21_X1 U16045 ( .B1(n14241), .B2(n14114), .A(n14113), .ZN(n14115) );
  OAI21_X1 U16046 ( .B1(n14243), .B2(n14116), .A(n14115), .ZN(P1_U3272) );
  OAI211_X1 U16047 ( .C1(n14119), .C2(n14118), .A(n14117), .B(n14264), .ZN(
        n14121) );
  XNOR2_X1 U16048 ( .A(n14124), .B(n14140), .ZN(n14245) );
  AOI22_X1 U16049 ( .A1(n14159), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14122), 
        .B2(n14157), .ZN(n14123) );
  OAI21_X1 U16050 ( .B1(n14124), .B2(n14161), .A(n14123), .ZN(n14129) );
  OAI21_X1 U16051 ( .B1(n14127), .B2(n14126), .A(n14125), .ZN(n14248) );
  NOR2_X1 U16052 ( .A1(n14248), .A2(n14164), .ZN(n14128) );
  AOI211_X1 U16053 ( .C1(n14245), .C2(n14167), .A(n14129), .B(n14128), .ZN(
        n14130) );
  OAI21_X1 U16054 ( .B1(n14159), .B2(n14247), .A(n14130), .ZN(P1_U3273) );
  AOI21_X1 U16055 ( .B1(n14133), .B2(n14132), .A(n14131), .ZN(n14134) );
  OAI222_X1 U16056 ( .A1(n14138), .A2(n14137), .B1(n14136), .B2(n14135), .C1(
        n14275), .C2(n14134), .ZN(n14139) );
  INV_X1 U16057 ( .A(n14139), .ZN(n14252) );
  AOI21_X1 U16058 ( .B1(n14249), .B2(n14155), .A(n7009), .ZN(n14250) );
  AOI22_X1 U16059 ( .A1(n14159), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14141), 
        .B2(n14157), .ZN(n14142) );
  OAI21_X1 U16060 ( .B1(n14143), .B2(n14161), .A(n14142), .ZN(n14147) );
  XNOR2_X1 U16061 ( .A(n14145), .B(n14144), .ZN(n14253) );
  NOR2_X1 U16062 ( .A1(n14253), .A2(n14164), .ZN(n14146) );
  AOI211_X1 U16063 ( .C1(n14250), .C2(n14167), .A(n14147), .B(n14146), .ZN(
        n14148) );
  OAI21_X1 U16064 ( .B1(n14252), .B2(n14159), .A(n14148), .ZN(P1_U3274) );
  XNOR2_X1 U16065 ( .A(n14150), .B(n14149), .ZN(n14151) );
  AOI222_X1 U16066 ( .A1(n14440), .A2(n14154), .B1(n14153), .B2(n14152), .C1(
        n14264), .C2(n14151), .ZN(n14257) );
  AOI21_X1 U16067 ( .B1(n14254), .B2(n6546), .A(n7010), .ZN(n14255) );
  INV_X1 U16068 ( .A(n14156), .ZN(n14158) );
  AOI22_X1 U16069 ( .A1(n14159), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14158), 
        .B2(n14157), .ZN(n14160) );
  OAI21_X1 U16070 ( .B1(n11599), .B2(n14161), .A(n14160), .ZN(n14166) );
  XNOR2_X1 U16071 ( .A(n14163), .B(n14162), .ZN(n14258) );
  NOR2_X1 U16072 ( .A1(n14258), .A2(n14164), .ZN(n14165) );
  AOI211_X1 U16073 ( .C1(n14255), .C2(n14167), .A(n14166), .B(n14165), .ZN(
        n14168) );
  OAI21_X1 U16074 ( .B1(n14257), .B2(n14159), .A(n14168), .ZN(P1_U3275) );
  NAND2_X1 U16075 ( .A1(n14169), .A2(n14618), .ZN(n14170) );
  OAI211_X1 U16076 ( .C1(n14171), .C2(n14609), .A(n14170), .B(n14173), .ZN(
        n14276) );
  MUX2_X1 U16077 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14276), .S(n14636), .Z(
        P1_U3559) );
  NAND2_X1 U16078 ( .A1(n14172), .A2(n14618), .ZN(n14174) );
  OAI211_X1 U16079 ( .C1(n14175), .C2(n14609), .A(n14174), .B(n14173), .ZN(
        n14277) );
  MUX2_X1 U16080 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14277), .S(n14636), .Z(
        P1_U3558) );
  NAND2_X1 U16081 ( .A1(n14176), .A2(n14615), .ZN(n14186) );
  OAI211_X1 U16082 ( .C1(n14179), .C2(n14609), .A(n14178), .B(n14177), .ZN(
        n14180) );
  AOI21_X1 U16083 ( .B1(n14181), .B2(n14618), .A(n14180), .ZN(n14182) );
  OAI21_X1 U16084 ( .B1(n14183), .B2(n14275), .A(n14182), .ZN(n14184) );
  INV_X1 U16085 ( .A(n14184), .ZN(n14185) );
  NAND2_X1 U16086 ( .A1(n14186), .A2(n14185), .ZN(n14278) );
  MUX2_X1 U16087 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14278), .S(n14636), .Z(
        P1_U3557) );
  INV_X1 U16088 ( .A(n14188), .ZN(n14193) );
  OAI22_X1 U16089 ( .A1(n14190), .A2(n9590), .B1(n14189), .B2(n14609), .ZN(
        n14191) );
  INV_X1 U16090 ( .A(n14191), .ZN(n14192) );
  NAND3_X1 U16091 ( .A1(n14194), .A2(n14193), .A3(n14192), .ZN(n14279) );
  MUX2_X1 U16092 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14279), .S(n14636), .Z(
        P1_U3556) );
  AOI22_X1 U16093 ( .A1(n14196), .A2(n14618), .B1(n14617), .B2(n14195), .ZN(
        n14197) );
  OAI21_X1 U16094 ( .B1(n14198), .B2(n14219), .A(n14197), .ZN(n14199) );
  AOI22_X1 U16095 ( .A1(n14202), .A2(n14618), .B1(n14617), .B2(n14201), .ZN(
        n14203) );
  OAI211_X1 U16096 ( .C1(n14623), .C2(n14205), .A(n14204), .B(n14203), .ZN(
        n14280) );
  MUX2_X1 U16097 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14280), .S(n14636), .Z(
        P1_U3554) );
  NOR2_X1 U16098 ( .A1(n14206), .A2(n9590), .ZN(n14207) );
  AOI211_X1 U16099 ( .C1(n14617), .C2(n14209), .A(n14208), .B(n14207), .ZN(
        n14212) );
  NAND2_X1 U16100 ( .A1(n14210), .A2(n14615), .ZN(n14211) );
  OAI211_X1 U16101 ( .C1(n14213), .C2(n14275), .A(n14212), .B(n14211), .ZN(
        n14281) );
  MUX2_X1 U16102 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14281), .S(n14636), .Z(
        P1_U3553) );
  INV_X1 U16103 ( .A(n14214), .ZN(n14220) );
  AOI21_X1 U16104 ( .B1(n14617), .B2(n14216), .A(n14215), .ZN(n14217) );
  OAI211_X1 U16105 ( .C1(n14220), .C2(n14219), .A(n14218), .B(n14217), .ZN(
        n14282) );
  MUX2_X1 U16106 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14282), .S(n14636), .Z(
        P1_U3552) );
  NOR2_X1 U16107 ( .A1(n11600), .A2(n14609), .ZN(n14222) );
  AOI211_X1 U16108 ( .C1(n14223), .C2(n14618), .A(n14222), .B(n14221), .ZN(
        n14226) );
  NAND2_X1 U16109 ( .A1(n14224), .A2(n14615), .ZN(n14225) );
  OAI211_X1 U16110 ( .C1(n14227), .C2(n14275), .A(n14226), .B(n14225), .ZN(
        n14283) );
  MUX2_X1 U16111 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14283), .S(n14636), .Z(
        P1_U3551) );
  NAND2_X1 U16112 ( .A1(n14228), .A2(n14617), .ZN(n14229) );
  OAI211_X1 U16113 ( .C1(n14231), .C2(n9590), .A(n14230), .B(n14229), .ZN(
        n14232) );
  AOI21_X1 U16114 ( .B1(n14233), .B2(n14615), .A(n14232), .ZN(n14234) );
  OAI21_X1 U16115 ( .B1(n14235), .B2(n14275), .A(n14234), .ZN(n14284) );
  MUX2_X1 U16116 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14284), .S(n14636), .Z(
        P1_U3550) );
  NAND2_X1 U16117 ( .A1(n14236), .A2(n14617), .ZN(n14237) );
  OAI211_X1 U16118 ( .C1(n14239), .C2(n9590), .A(n14238), .B(n14237), .ZN(
        n14240) );
  AOI21_X1 U16119 ( .B1(n14241), .B2(n14615), .A(n14240), .ZN(n14242) );
  OAI21_X1 U16120 ( .B1(n14243), .B2(n14275), .A(n14242), .ZN(n14285) );
  MUX2_X1 U16121 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14285), .S(n14636), .Z(
        P1_U3549) );
  AOI22_X1 U16122 ( .A1(n14245), .A2(n14618), .B1(n14617), .B2(n14244), .ZN(
        n14246) );
  OAI211_X1 U16123 ( .C1(n14623), .C2(n14248), .A(n14247), .B(n14246), .ZN(
        n14286) );
  MUX2_X1 U16124 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14286), .S(n14636), .Z(
        P1_U3548) );
  AOI22_X1 U16125 ( .A1(n14250), .A2(n14618), .B1(n14617), .B2(n14249), .ZN(
        n14251) );
  OAI211_X1 U16126 ( .C1(n14623), .C2(n14253), .A(n14252), .B(n14251), .ZN(
        n14287) );
  MUX2_X1 U16127 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14287), .S(n14636), .Z(
        P1_U3547) );
  AOI22_X1 U16128 ( .A1(n14255), .A2(n14618), .B1(n14617), .B2(n14254), .ZN(
        n14256) );
  OAI211_X1 U16129 ( .C1(n14623), .C2(n14258), .A(n14257), .B(n14256), .ZN(
        n14288) );
  MUX2_X1 U16130 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14288), .S(n14636), .Z(
        P1_U3546) );
  NAND2_X1 U16131 ( .A1(n14259), .A2(n14617), .ZN(n14260) );
  OAI211_X1 U16132 ( .C1(n14262), .C2(n9590), .A(n14261), .B(n14260), .ZN(
        n14263) );
  AOI21_X1 U16133 ( .B1(n14265), .B2(n14264), .A(n14263), .ZN(n14266) );
  OAI21_X1 U16134 ( .B1(n14623), .B2(n14267), .A(n14266), .ZN(n14289) );
  MUX2_X1 U16135 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14289), .S(n14636), .Z(
        P1_U3545) );
  AOI21_X1 U16136 ( .B1(n14450), .B2(n14617), .A(n14268), .ZN(n14269) );
  OAI21_X1 U16137 ( .B1(n14270), .B2(n9590), .A(n14269), .ZN(n14271) );
  AOI21_X1 U16138 ( .B1(n14272), .B2(n14615), .A(n14271), .ZN(n14273) );
  OAI21_X1 U16139 ( .B1(n14275), .B2(n14274), .A(n14273), .ZN(n14290) );
  MUX2_X1 U16140 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14290), .S(n14636), .Z(
        P1_U3544) );
  MUX2_X1 U16141 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14276), .S(n14627), .Z(
        P1_U3527) );
  MUX2_X1 U16142 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14277), .S(n14627), .Z(
        P1_U3526) );
  MUX2_X1 U16143 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14278), .S(n14627), .Z(
        P1_U3525) );
  MUX2_X1 U16144 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14279), .S(n14627), .Z(
        P1_U3524) );
  MUX2_X1 U16145 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14280), .S(n14627), .Z(
        P1_U3522) );
  MUX2_X1 U16146 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14281), .S(n14627), .Z(
        P1_U3521) );
  MUX2_X1 U16147 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14282), .S(n14627), .Z(
        P1_U3520) );
  MUX2_X1 U16148 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14283), .S(n14627), .Z(
        P1_U3519) );
  MUX2_X1 U16149 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14284), .S(n14627), .Z(
        P1_U3518) );
  MUX2_X1 U16150 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14285), .S(n14627), .Z(
        P1_U3517) );
  MUX2_X1 U16151 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14286), .S(n14627), .Z(
        P1_U3516) );
  MUX2_X1 U16152 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14287), .S(n14627), .Z(
        P1_U3515) );
  MUX2_X1 U16153 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14288), .S(n14627), .Z(
        P1_U3513) );
  MUX2_X1 U16154 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14289), .S(n14627), .Z(
        P1_U3510) );
  MUX2_X1 U16155 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14290), .S(n14627), .Z(
        P1_U3507) );
  NAND3_X1 U16156 ( .A1(n14292), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14294) );
  OAI22_X1 U16157 ( .A1(n14291), .A2(n14294), .B1(n14293), .B2(n14302), .ZN(
        n14295) );
  AOI21_X1 U16158 ( .B1(n14297), .B2(n14296), .A(n14295), .ZN(n14298) );
  INV_X1 U16159 ( .A(n14298), .ZN(P1_U3324) );
  OAI222_X1 U16160 ( .A1(n14302), .A2(n14301), .B1(n14305), .B2(n14300), .C1(
        P1_U3086), .C2(n14299), .ZN(P1_U3326) );
  OAI222_X1 U16161 ( .A1(P1_U3086), .A2(n6530), .B1(n14305), .B2(n14304), .C1(
        n14303), .C2(n14302), .ZN(P1_U3328) );
  MUX2_X1 U16162 ( .A(n8348), .B(n14307), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16163 ( .A(n14308), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U16164 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14312) );
  OAI21_X1 U16165 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14312), 
        .ZN(U28) );
  OAI21_X1 U16166 ( .B1(n14315), .B2(n14314), .A(n14313), .ZN(n14316) );
  XNOR2_X1 U16167 ( .A(n14316), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16168 ( .B1(n14319), .B2(n14318), .A(n14317), .ZN(SUB_1596_U57) );
  OAI21_X1 U16169 ( .B1(n14321), .B2(n15086), .A(n14320), .ZN(SUB_1596_U55) );
  OAI21_X1 U16170 ( .B1(n14324), .B2(n14323), .A(n14322), .ZN(n14325) );
  XNOR2_X1 U16171 ( .A(n14325), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  OAI21_X1 U16172 ( .B1(n14328), .B2(n14327), .A(n14326), .ZN(n14329) );
  XNOR2_X1 U16173 ( .A(n14329), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI21_X1 U16174 ( .B1(n14331), .B2(n15226), .A(n14330), .ZN(SUB_1596_U63) );
  NAND2_X1 U16175 ( .A1(n14333), .A2(n14332), .ZN(n14335) );
  OAI211_X1 U16176 ( .C1(n14337), .C2(n14336), .A(n14335), .B(n14334), .ZN(
        n14338) );
  INV_X1 U16177 ( .A(n14338), .ZN(n14346) );
  XNOR2_X1 U16178 ( .A(n14340), .B(n14339), .ZN(n14344) );
  AOI22_X1 U16179 ( .A1(n14344), .A2(n14343), .B1(n14342), .B2(n14341), .ZN(
        n14345) );
  OAI211_X1 U16180 ( .C1(n14348), .C2(n14347), .A(n14346), .B(n14345), .ZN(
        P3_U3181) );
  INV_X1 U16181 ( .A(n14349), .ZN(n14350) );
  AOI22_X1 U16182 ( .A1(n14352), .A2(n14952), .B1(n14386), .B2(n14955), .ZN(
        n14358) );
  OAI22_X1 U16183 ( .A1(n14383), .A2(n14354), .B1(n14353), .B2(n14955), .ZN(
        n14355) );
  INV_X1 U16184 ( .A(n14355), .ZN(n14356) );
  NAND2_X1 U16185 ( .A1(n14358), .A2(n14356), .ZN(P3_U3202) );
  AOI22_X1 U16186 ( .A1(n14387), .A2(n14919), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n14957), .ZN(n14357) );
  NAND2_X1 U16187 ( .A1(n14358), .A2(n14357), .ZN(P3_U3203) );
  XNOR2_X1 U16188 ( .A(n14359), .B(n14364), .ZN(n14361) );
  AOI222_X1 U16189 ( .A1(n14934), .A2(n14361), .B1(n14360), .B2(n14944), .C1(
        n14372), .C2(n14946), .ZN(n14389) );
  INV_X1 U16190 ( .A(n14362), .ZN(n14363) );
  AOI22_X1 U16191 ( .A1(P3_REG2_REG_13__SCAN_IN), .A2(n14957), .B1(n14952), 
        .B2(n14363), .ZN(n14369) );
  XNOR2_X1 U16192 ( .A(n14365), .B(n14364), .ZN(n14392) );
  INV_X1 U16193 ( .A(n14366), .ZN(n14367) );
  NOR2_X1 U16194 ( .A1(n14367), .A2(n15013), .ZN(n14391) );
  AOI22_X1 U16195 ( .A1(n14392), .A2(n14380), .B1(n14391), .B2(n14379), .ZN(
        n14368) );
  OAI211_X1 U16196 ( .C1(n14957), .C2(n14389), .A(n14369), .B(n14368), .ZN(
        P3_U3220) );
  XOR2_X1 U16197 ( .A(n14370), .B(n14376), .Z(n14373) );
  AOI222_X1 U16198 ( .A1(n14934), .A2(n14373), .B1(n14372), .B2(n14944), .C1(
        n14371), .C2(n14946), .ZN(n14399) );
  OAI22_X1 U16199 ( .A1(n14955), .A2(n8686), .B1(n14926), .B2(n14374), .ZN(
        n14375) );
  INV_X1 U16200 ( .A(n14375), .ZN(n14382) );
  XNOR2_X1 U16201 ( .A(n14377), .B(n14376), .ZN(n14402) );
  NOR2_X1 U16202 ( .A1(n14378), .A2(n15013), .ZN(n14401) );
  AOI22_X1 U16203 ( .A1(n14402), .A2(n14380), .B1(n14401), .B2(n14379), .ZN(
        n14381) );
  OAI211_X1 U16204 ( .C1(n14957), .C2(n14399), .A(n14382), .B(n14381), .ZN(
        P3_U3222) );
  OR2_X1 U16205 ( .A1(n14383), .A2(n15013), .ZN(n14385) );
  INV_X1 U16206 ( .A(n14386), .ZN(n14384) );
  AOI22_X1 U16207 ( .A1(n15031), .A2(n14404), .B1(n15181), .B2(n15029), .ZN(
        P3_U3490) );
  AOI21_X1 U16208 ( .B1(n14387), .B2(n14980), .A(n14386), .ZN(n14406) );
  INV_X1 U16209 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U16210 ( .A1(n15031), .A2(n14406), .B1(n14388), .B2(n15029), .ZN(
        P3_U3489) );
  INV_X1 U16211 ( .A(n14389), .ZN(n14390) );
  AOI211_X1 U16212 ( .C1(n14392), .C2(n15011), .A(n14391), .B(n14390), .ZN(
        n14407) );
  AOI22_X1 U16213 ( .A1(n15031), .A2(n14407), .B1(n14888), .B2(n15029), .ZN(
        P3_U3472) );
  NOR2_X1 U16214 ( .A1(n14393), .A2(n15013), .ZN(n14396) );
  INV_X1 U16215 ( .A(n14394), .ZN(n14395) );
  AOI211_X1 U16216 ( .C1(n15011), .C2(n14397), .A(n14396), .B(n14395), .ZN(
        n14409) );
  AOI22_X1 U16217 ( .A1(n15031), .A2(n14409), .B1(n14398), .B2(n15029), .ZN(
        P3_U3471) );
  INV_X1 U16218 ( .A(n14399), .ZN(n14400) );
  AOI211_X1 U16219 ( .C1(n15011), .C2(n14402), .A(n14401), .B(n14400), .ZN(
        n14411) );
  AOI22_X1 U16220 ( .A1(n15031), .A2(n14411), .B1(n8687), .B2(n15029), .ZN(
        P3_U3470) );
  INV_X1 U16221 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14403) );
  AOI22_X1 U16222 ( .A1(n15019), .A2(n14404), .B1(n14403), .B2(n15018), .ZN(
        P3_U3458) );
  AOI22_X1 U16223 ( .A1(n15019), .A2(n14406), .B1(n14405), .B2(n15018), .ZN(
        P3_U3457) );
  AOI22_X1 U16224 ( .A1(n15019), .A2(n14407), .B1(n8717), .B2(n15018), .ZN(
        P3_U3429) );
  INV_X1 U16225 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U16226 ( .A1(n15019), .A2(n14409), .B1(n14408), .B2(n15018), .ZN(
        P3_U3426) );
  INV_X1 U16227 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14410) );
  AOI22_X1 U16228 ( .A1(n15019), .A2(n14411), .B1(n14410), .B2(n15018), .ZN(
        P3_U3423) );
  OAI21_X1 U16229 ( .B1(n14414), .B2(n14413), .A(n14412), .ZN(n14423) );
  NOR2_X1 U16230 ( .A1(n14416), .A2(n14415), .ZN(n14422) );
  OAI22_X1 U16231 ( .A1(n14420), .A2(n14419), .B1(n14418), .B2(n14417), .ZN(
        n14421) );
  AOI211_X1 U16232 ( .C1(n14423), .C2(n14644), .A(n14422), .B(n14421), .ZN(
        n14425) );
  OAI211_X1 U16233 ( .C1(n14660), .C2(n14426), .A(n14425), .B(n14424), .ZN(
        P2_U3187) );
  OAI22_X1 U16234 ( .A1(n14427), .A2(n14470), .B1(n14471), .B2(n14441), .ZN(
        n14435) );
  AOI21_X1 U16235 ( .B1(n14430), .B2(n14429), .A(n14428), .ZN(n14431) );
  INV_X1 U16236 ( .A(n14431), .ZN(n14433) );
  AOI21_X1 U16237 ( .B1(n14433), .B2(n14432), .A(n14476), .ZN(n14434) );
  AOI211_X1 U16238 ( .C1(n14436), .C2(n14481), .A(n14435), .B(n14434), .ZN(
        n14438) );
  OAI211_X1 U16239 ( .C1(n14485), .C2(n14439), .A(n14438), .B(n14437), .ZN(
        P1_U3215) );
  OAI22_X1 U16240 ( .A1(n14441), .A2(n14470), .B1(n14471), .B2(n11584), .ZN(
        n14449) );
  INV_X1 U16241 ( .A(n14442), .ZN(n14445) );
  OAI21_X1 U16242 ( .B1(n14445), .B2(n14444), .A(n14443), .ZN(n14447) );
  AOI21_X1 U16243 ( .B1(n14447), .B2(n14446), .A(n14476), .ZN(n14448) );
  AOI211_X1 U16244 ( .C1(n14450), .C2(n14481), .A(n14449), .B(n14448), .ZN(
        n14452) );
  OAI211_X1 U16245 ( .C1(n14485), .C2(n14453), .A(n14452), .B(n14451), .ZN(
        P1_U3226) );
  XNOR2_X1 U16246 ( .A(n14455), .B(n14454), .ZN(n14465) );
  AOI22_X1 U16247 ( .A1(n14459), .A2(n14458), .B1(n14457), .B2(n14456), .ZN(
        n14460) );
  OAI21_X1 U16248 ( .B1(n14462), .B2(n14461), .A(n14460), .ZN(n14463) );
  AOI21_X1 U16249 ( .B1(n14465), .B2(n14464), .A(n14463), .ZN(n14467) );
  OAI211_X1 U16250 ( .C1(n14485), .C2(n14468), .A(n14467), .B(n14466), .ZN(
        P1_U3228) );
  OAI22_X1 U16251 ( .A1(n14472), .A2(n14471), .B1(n14470), .B2(n14469), .ZN(
        n14480) );
  AOI21_X1 U16252 ( .B1(n13595), .B2(n14474), .A(n14473), .ZN(n14475) );
  INV_X1 U16253 ( .A(n14475), .ZN(n14478) );
  AOI21_X1 U16254 ( .B1(n14478), .B2(n14477), .A(n14476), .ZN(n14479) );
  AOI211_X1 U16255 ( .C1(n14504), .C2(n14481), .A(n14480), .B(n14479), .ZN(
        n14483) );
  OAI211_X1 U16256 ( .C1(n14485), .C2(n14484), .A(n14483), .B(n14482), .ZN(
        P1_U3236) );
  OAI22_X1 U16257 ( .A1(n14487), .A2(n9590), .B1(n14486), .B2(n14609), .ZN(
        n14489) );
  AOI211_X1 U16258 ( .C1(n14490), .C2(n14615), .A(n14489), .B(n14488), .ZN(
        n14510) );
  AOI22_X1 U16259 ( .A1(n14636), .A2(n14510), .B1(n8032), .B2(n14634), .ZN(
        P1_U3543) );
  INV_X1 U16260 ( .A(n14491), .ZN(n14496) );
  OAI22_X1 U16261 ( .A1(n14493), .A2(n9590), .B1(n14492), .B2(n14609), .ZN(
        n14495) );
  AOI211_X1 U16262 ( .C1(n14496), .C2(n14615), .A(n14495), .B(n14494), .ZN(
        n14512) );
  AOI22_X1 U16263 ( .A1(n14636), .A2(n14512), .B1(n8014), .B2(n14634), .ZN(
        P1_U3542) );
  OAI22_X1 U16264 ( .A1(n14498), .A2(n9590), .B1(n14497), .B2(n14609), .ZN(
        n14499) );
  AOI21_X1 U16265 ( .B1(n14500), .B2(n14615), .A(n14499), .ZN(n14501) );
  AND2_X1 U16266 ( .A1(n14502), .A2(n14501), .ZN(n14513) );
  AOI22_X1 U16267 ( .A1(n14636), .A2(n14513), .B1(n14503), .B2(n14634), .ZN(
        P1_U3541) );
  OAI22_X1 U16268 ( .A1(n14505), .A2(n9590), .B1(n7018), .B2(n14609), .ZN(
        n14506) );
  AOI21_X1 U16269 ( .B1(n14507), .B2(n14615), .A(n14506), .ZN(n14508) );
  AOI22_X1 U16270 ( .A1(n14636), .A2(n14515), .B1(n7929), .B2(n14634), .ZN(
        P1_U3539) );
  AOI22_X1 U16271 ( .A1(n14627), .A2(n14510), .B1(n8033), .B2(n14625), .ZN(
        P1_U3504) );
  INV_X1 U16272 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14511) );
  AOI22_X1 U16273 ( .A1(n14627), .A2(n14512), .B1(n14511), .B2(n14625), .ZN(
        P1_U3501) );
  AOI22_X1 U16274 ( .A1(n14627), .A2(n14513), .B1(n7972), .B2(n14625), .ZN(
        P1_U3498) );
  INV_X1 U16275 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14514) );
  AOI22_X1 U16276 ( .A1(n14627), .A2(n14515), .B1(n14514), .B2(n14625), .ZN(
        P1_U3492) );
  OAI21_X1 U16277 ( .B1(n14518), .B2(n14517), .A(n14516), .ZN(n14519) );
  XNOR2_X1 U16278 ( .A(n14519), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI222_X1 U16279 ( .A1(n14745), .A2(n14522), .B1(n14745), .B2(n6787), .C1(
        n14521), .C2(n14520), .ZN(SUB_1596_U68) );
  OAI222_X1 U16280 ( .A1(n14527), .A2(n14526), .B1(n14527), .B2(n14525), .C1(
        n14524), .C2(n14523), .ZN(SUB_1596_U67) );
  OAI222_X1 U16281 ( .A1(n14532), .A2(n14531), .B1(n14532), .B2(n14530), .C1(
        n14529), .C2(n14528), .ZN(SUB_1596_U66) );
  OAI21_X1 U16282 ( .B1(n14535), .B2(n14534), .A(n14533), .ZN(n14536) );
  XNOR2_X1 U16283 ( .A(n14536), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  OAI21_X1 U16284 ( .B1(n14539), .B2(n14538), .A(n14537), .ZN(n14540) );
  XNOR2_X1 U16285 ( .A(n14540), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  OAI21_X1 U16286 ( .B1(n14542), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14541), .ZN(
        n14543) );
  XOR2_X1 U16287 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14543), .Z(n14547) );
  AOI22_X1 U16288 ( .A1(n14544), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14545) );
  OAI21_X1 U16289 ( .B1(n14547), .B2(n14546), .A(n14545), .ZN(P1_U3243) );
  AOI21_X1 U16290 ( .B1(n14549), .B2(P1_REG1_REG_15__SCAN_IN), .A(n14548), 
        .ZN(n14558) );
  AOI21_X1 U16291 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14551), .A(n14550), 
        .ZN(n14553) );
  OR2_X1 U16292 ( .A1(n14553), .A2(n14552), .ZN(n14556) );
  OR2_X1 U16293 ( .A1(n14571), .A2(n14554), .ZN(n14555) );
  OAI211_X1 U16294 ( .C1(n14558), .C2(n14557), .A(n14556), .B(n14555), .ZN(
        n14559) );
  INV_X1 U16295 ( .A(n14559), .ZN(n14561) );
  NAND2_X1 U16296 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14560)
         );
  OAI211_X1 U16297 ( .C1(n15085), .C2(n14575), .A(n14561), .B(n14560), .ZN(
        P1_U3258) );
  OAI211_X1 U16298 ( .C1(n14564), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14563), 
        .B(n14562), .ZN(n14569) );
  OAI211_X1 U16299 ( .C1(n14567), .C2(P1_REG1_REG_18__SCAN_IN), .A(n14566), 
        .B(n14565), .ZN(n14568) );
  OAI211_X1 U16300 ( .C1(n14571), .C2(n14570), .A(n14569), .B(n14568), .ZN(
        n14572) );
  INV_X1 U16301 ( .A(n14572), .ZN(n14574) );
  OAI211_X1 U16302 ( .C1(n14576), .C2(n14575), .A(n14574), .B(n14573), .ZN(
        P1_U3261) );
  AND2_X1 U16303 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14578), .ZN(P1_U3294) );
  AND2_X1 U16304 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14578), .ZN(P1_U3295) );
  AND2_X1 U16305 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14578), .ZN(P1_U3296) );
  AND2_X1 U16306 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14578), .ZN(P1_U3297) );
  AND2_X1 U16307 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14578), .ZN(P1_U3298) );
  AND2_X1 U16308 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14578), .ZN(P1_U3299) );
  AND2_X1 U16309 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14578), .ZN(P1_U3300) );
  INV_X1 U16310 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15272) );
  NOR2_X1 U16311 ( .A1(n14577), .A2(n15272), .ZN(P1_U3301) );
  AND2_X1 U16312 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14578), .ZN(P1_U3302) );
  INV_X1 U16313 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15246) );
  NOR2_X1 U16314 ( .A1(n14577), .A2(n15246), .ZN(P1_U3303) );
  AND2_X1 U16315 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14578), .ZN(P1_U3304) );
  AND2_X1 U16316 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14578), .ZN(P1_U3305) );
  AND2_X1 U16317 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14578), .ZN(P1_U3306) );
  AND2_X1 U16318 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14578), .ZN(P1_U3307) );
  AND2_X1 U16319 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14578), .ZN(P1_U3308) );
  AND2_X1 U16320 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14578), .ZN(P1_U3309) );
  AND2_X1 U16321 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14578), .ZN(P1_U3310) );
  AND2_X1 U16322 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14578), .ZN(P1_U3311) );
  INV_X1 U16323 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15240) );
  NOR2_X1 U16324 ( .A1(n14577), .A2(n15240), .ZN(P1_U3312) );
  AND2_X1 U16325 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14578), .ZN(P1_U3313) );
  AND2_X1 U16326 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14578), .ZN(P1_U3314) );
  AND2_X1 U16327 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14578), .ZN(P1_U3315) );
  AND2_X1 U16328 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14578), .ZN(P1_U3316) );
  AND2_X1 U16329 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14578), .ZN(P1_U3317) );
  AND2_X1 U16330 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14578), .ZN(P1_U3318) );
  INV_X1 U16331 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15164) );
  NOR2_X1 U16332 ( .A1(n14577), .A2(n15164), .ZN(P1_U3319) );
  AND2_X1 U16333 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14578), .ZN(P1_U3320) );
  INV_X1 U16334 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15199) );
  NOR2_X1 U16335 ( .A1(n14577), .A2(n15199), .ZN(P1_U3321) );
  AND2_X1 U16336 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14578), .ZN(P1_U3322) );
  AND2_X1 U16337 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14578), .ZN(P1_U3323) );
  OAI22_X1 U16338 ( .A1(n14579), .A2(n9590), .B1(n7725), .B2(n14609), .ZN(
        n14582) );
  INV_X1 U16339 ( .A(n14580), .ZN(n14581) );
  AOI211_X1 U16340 ( .C1(n14608), .C2(n14583), .A(n14582), .B(n14581), .ZN(
        n14628) );
  AOI22_X1 U16341 ( .A1(n14627), .A2(n14628), .B1(n7679), .B2(n14625), .ZN(
        P1_U3462) );
  INV_X1 U16342 ( .A(n14584), .ZN(n14589) );
  OAI22_X1 U16343 ( .A1(n14586), .A2(n9590), .B1(n14585), .B2(n14609), .ZN(
        n14588) );
  AOI211_X1 U16344 ( .C1(n14608), .C2(n14589), .A(n14588), .B(n14587), .ZN(
        n14629) );
  AOI22_X1 U16345 ( .A1(n14627), .A2(n14629), .B1(n7732), .B2(n14625), .ZN(
        P1_U3465) );
  INV_X1 U16346 ( .A(n14590), .ZN(n14596) );
  OAI22_X1 U16347 ( .A1(n14592), .A2(n9590), .B1(n14591), .B2(n14609), .ZN(
        n14595) );
  INV_X1 U16348 ( .A(n14593), .ZN(n14594) );
  AOI211_X1 U16349 ( .C1(n14608), .C2(n14596), .A(n14595), .B(n14594), .ZN(
        n14630) );
  INV_X1 U16350 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14597) );
  AOI22_X1 U16351 ( .A1(n14627), .A2(n14630), .B1(n14597), .B2(n14625), .ZN(
        P1_U3468) );
  OAI22_X1 U16352 ( .A1(n14599), .A2(n9590), .B1(n14598), .B2(n14609), .ZN(
        n14601) );
  AOI211_X1 U16353 ( .C1(n14608), .C2(n14602), .A(n14601), .B(n14600), .ZN(
        n14631) );
  AOI22_X1 U16354 ( .A1(n14627), .A2(n14631), .B1(n7807), .B2(n14625), .ZN(
        P1_U3474) );
  OAI22_X1 U16355 ( .A1(n14604), .A2(n9590), .B1(n14603), .B2(n14609), .ZN(
        n14606) );
  AOI211_X1 U16356 ( .C1(n14608), .C2(n14607), .A(n14606), .B(n14605), .ZN(
        n14632) );
  AOI22_X1 U16357 ( .A1(n14627), .A2(n14632), .B1(n7842), .B2(n14625), .ZN(
        P1_U3480) );
  OAI22_X1 U16358 ( .A1(n14611), .A2(n9590), .B1(n14610), .B2(n14609), .ZN(
        n14613) );
  AOI211_X1 U16359 ( .C1(n14615), .C2(n14614), .A(n14613), .B(n14612), .ZN(
        n14633) );
  AOI22_X1 U16360 ( .A1(n14627), .A2(n14633), .B1(n7866), .B2(n14625), .ZN(
        P1_U3483) );
  AOI22_X1 U16361 ( .A1(n14619), .A2(n14618), .B1(n14617), .B2(n14616), .ZN(
        n14620) );
  OAI211_X1 U16362 ( .C1(n14623), .C2(n14622), .A(n14621), .B(n14620), .ZN(
        n14624) );
  INV_X1 U16363 ( .A(n14624), .ZN(n14635) );
  INV_X1 U16364 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14626) );
  AOI22_X1 U16365 ( .A1(n14627), .A2(n14635), .B1(n14626), .B2(n14625), .ZN(
        P1_U3486) );
  AOI22_X1 U16366 ( .A1(n14636), .A2(n14628), .B1(n15154), .B2(n14634), .ZN(
        P1_U3529) );
  AOI22_X1 U16367 ( .A1(n14636), .A2(n14629), .B1(n9412), .B2(n14634), .ZN(
        P1_U3530) );
  AOI22_X1 U16368 ( .A1(n14636), .A2(n14630), .B1(n9415), .B2(n14634), .ZN(
        P1_U3531) );
  AOI22_X1 U16369 ( .A1(n14636), .A2(n14631), .B1(n7806), .B2(n14634), .ZN(
        P1_U3533) );
  AOI22_X1 U16370 ( .A1(n14636), .A2(n14632), .B1(n9426), .B2(n14634), .ZN(
        P1_U3535) );
  AOI22_X1 U16371 ( .A1(n14636), .A2(n14633), .B1(n9428), .B2(n14634), .ZN(
        P1_U3536) );
  AOI22_X1 U16372 ( .A1(n14636), .A2(n14635), .B1(n7885), .B2(n14634), .ZN(
        P1_U3537) );
  NOR2_X1 U16373 ( .A1(n14768), .A2(P2_U3947), .ZN(P2_U3087) );
  XOR2_X1 U16374 ( .A(n14638), .B(n14637), .Z(n14645) );
  NAND2_X1 U16375 ( .A1(n14639), .A2(n14657), .ZN(n14641) );
  OAI211_X1 U16376 ( .C1(n14642), .C2(n14649), .A(n14641), .B(n14640), .ZN(
        n14643) );
  AOI21_X1 U16377 ( .B1(n14645), .B2(n14644), .A(n14643), .ZN(n14646) );
  OAI21_X1 U16378 ( .B1(n14647), .B2(n14660), .A(n14646), .ZN(P2_U3189) );
  OAI22_X1 U16379 ( .A1(n14650), .A2(n14649), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14648), .ZN(n14656) );
  AOI211_X1 U16380 ( .C1(n14654), .C2(n14653), .A(n14652), .B(n14651), .ZN(
        n14655) );
  AOI211_X1 U16381 ( .C1(n14658), .C2(n14657), .A(n14656), .B(n14655), .ZN(
        n14659) );
  OAI21_X1 U16382 ( .B1(n14661), .B2(n14660), .A(n14659), .ZN(P2_U3206) );
  AOI22_X1 U16383 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n14774), .B1(n14776), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n14665) );
  AOI22_X1 U16384 ( .A1(n14768), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14664) );
  OAI22_X1 U16385 ( .A1(n14738), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14747), .ZN(n14662) );
  OAI21_X1 U16386 ( .B1(n14770), .B2(n14662), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14663) );
  OAI211_X1 U16387 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14665), .A(n14664), .B(
        n14663), .ZN(P2_U3214) );
  INV_X1 U16388 ( .A(n14666), .ZN(n14667) );
  AOI22_X1 U16389 ( .A1(n14768), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n14770), 
        .B2(n14667), .ZN(n14677) );
  OAI211_X1 U16390 ( .C1(n14670), .C2(n14669), .A(n14776), .B(n14668), .ZN(
        n14676) );
  OAI211_X1 U16391 ( .C1(n14673), .C2(n14672), .A(n14774), .B(n14671), .ZN(
        n14675) );
  NAND2_X1 U16392 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(P2_U3088), .ZN(n14674) );
  NAND4_X1 U16393 ( .A1(n14677), .A2(n14676), .A3(n14675), .A4(n14674), .ZN(
        P2_U3216) );
  AOI22_X1 U16394 ( .A1(n14768), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(n14770), 
        .B2(n14678), .ZN(n14689) );
  INV_X1 U16395 ( .A(n14679), .ZN(n14688) );
  OAI211_X1 U16396 ( .C1(n14682), .C2(n14681), .A(n14774), .B(n14680), .ZN(
        n14687) );
  OAI211_X1 U16397 ( .C1(n14685), .C2(n14684), .A(n14776), .B(n14683), .ZN(
        n14686) );
  NAND4_X1 U16398 ( .A1(n14689), .A2(n14688), .A3(n14687), .A4(n14686), .ZN(
        P2_U3217) );
  AOI22_X1 U16399 ( .A1(n14768), .A2(P2_ADDR_REG_6__SCAN_IN), .B1(n14770), 
        .B2(n14690), .ZN(n14700) );
  OAI211_X1 U16400 ( .C1(n14693), .C2(n14692), .A(n14774), .B(n14691), .ZN(
        n14698) );
  OAI211_X1 U16401 ( .C1(n14696), .C2(n14695), .A(n14776), .B(n14694), .ZN(
        n14697) );
  NAND4_X1 U16402 ( .A1(n14700), .A2(n14699), .A3(n14698), .A4(n14697), .ZN(
        P2_U3220) );
  INV_X1 U16403 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14716) );
  NOR2_X1 U16404 ( .A1(n14702), .A2(n14701), .ZN(n14703) );
  OAI21_X1 U16405 ( .B1(n14704), .B2(n14703), .A(n14776), .ZN(n14713) );
  INV_X1 U16406 ( .A(n14705), .ZN(n14706) );
  NAND2_X1 U16407 ( .A1(n14770), .A2(n14706), .ZN(n14712) );
  AND2_X1 U16408 ( .A1(n14708), .A2(n14707), .ZN(n14709) );
  OAI21_X1 U16409 ( .B1(n14710), .B2(n14709), .A(n14774), .ZN(n14711) );
  AND3_X1 U16410 ( .A1(n14713), .A2(n14712), .A3(n14711), .ZN(n14715) );
  OAI211_X1 U16411 ( .C1(n14716), .C2(n14744), .A(n14715), .B(n14714), .ZN(
        P2_U3223) );
  AOI21_X1 U16412 ( .B1(n14719), .B2(n14718), .A(n14717), .ZN(n14729) );
  INV_X1 U16413 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n14720) );
  NOR2_X1 U16414 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14720), .ZN(n14723) );
  NOR2_X1 U16415 ( .A1(n14740), .A2(n14721), .ZN(n14722) );
  AOI211_X1 U16416 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n14768), .A(n14723), 
        .B(n14722), .ZN(n14728) );
  OAI211_X1 U16417 ( .C1(n14726), .C2(n14725), .A(n14724), .B(n14774), .ZN(
        n14727) );
  OAI211_X1 U16418 ( .C1(n14729), .C2(n14738), .A(n14728), .B(n14727), .ZN(
        P2_U3225) );
  AOI21_X1 U16419 ( .B1(n14732), .B2(n14731), .A(n14730), .ZN(n14737) );
  AOI21_X1 U16420 ( .B1(n14735), .B2(n14734), .A(n14733), .ZN(n14736) );
  OAI222_X1 U16421 ( .A1(n14740), .A2(n14739), .B1(n14738), .B2(n14737), .C1(
        n14747), .C2(n14736), .ZN(n14741) );
  INV_X1 U16422 ( .A(n14741), .ZN(n14743) );
  NAND2_X1 U16423 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14742)
         );
  OAI211_X1 U16424 ( .C1(n14745), .C2(n14744), .A(n14743), .B(n14742), .ZN(
        P2_U3226) );
  AOI22_X1 U16425 ( .A1(n14768), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14758) );
  NAND2_X1 U16426 ( .A1(n14770), .A2(n14751), .ZN(n14757) );
  AOI211_X1 U16427 ( .C1(n14749), .C2(n14748), .A(n14747), .B(n14746), .ZN(
        n14750) );
  INV_X1 U16428 ( .A(n14750), .ZN(n14756) );
  MUX2_X1 U16429 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n10090), .S(n14751), .Z(
        n14754) );
  NAND2_X1 U16430 ( .A1(n14753), .A2(n14754), .ZN(n14752) );
  OAI211_X1 U16431 ( .C1(n14754), .C2(n14753), .A(n14776), .B(n14752), .ZN(
        n14755) );
  NAND4_X1 U16432 ( .A1(n14758), .A2(n14757), .A3(n14756), .A4(n14755), .ZN(
        P2_U3227) );
  AOI22_X1 U16433 ( .A1(n14768), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14767) );
  NAND2_X1 U16434 ( .A1(n14770), .A2(n14759), .ZN(n14766) );
  OAI211_X1 U16435 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14761), .A(n14776), 
        .B(n14760), .ZN(n14765) );
  XNOR2_X1 U16436 ( .A(n14762), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n14763) );
  NAND2_X1 U16437 ( .A1(n14763), .A2(n14774), .ZN(n14764) );
  NAND4_X1 U16438 ( .A1(n14767), .A2(n14766), .A3(n14765), .A4(n14764), .ZN(
        P2_U3229) );
  AOI22_X1 U16439 ( .A1(n14768), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n14782) );
  NAND2_X1 U16440 ( .A1(n14770), .A2(n14769), .ZN(n14781) );
  XNOR2_X1 U16441 ( .A(n14772), .B(n14771), .ZN(n14773) );
  NAND2_X1 U16442 ( .A1(n14774), .A2(n14773), .ZN(n14780) );
  OAI211_X1 U16443 ( .C1(n14778), .C2(n14777), .A(n14776), .B(n14775), .ZN(
        n14779) );
  NAND4_X1 U16444 ( .A1(n14782), .A2(n14781), .A3(n14780), .A4(n14779), .ZN(
        P2_U3231) );
  AOI22_X1 U16445 ( .A1(n14811), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14784), 
        .B2(n14783), .ZN(n14788) );
  NAND2_X1 U16446 ( .A1(n14786), .A2(n14785), .ZN(n14787) );
  OAI211_X1 U16447 ( .C1(n14790), .C2(n14789), .A(n14788), .B(n14787), .ZN(
        n14791) );
  AOI21_X1 U16448 ( .B1(n14793), .B2(n14792), .A(n14791), .ZN(n14794) );
  OAI21_X1 U16449 ( .B1(n14811), .B2(n14795), .A(n14794), .ZN(P2_U3258) );
  NOR2_X1 U16450 ( .A1(n14797), .A2(n14796), .ZN(n14825) );
  NOR2_X1 U16451 ( .A1(n14847), .A2(n14798), .ZN(n14801) );
  OAI22_X1 U16452 ( .A1(n14823), .A2(n14801), .B1(n14800), .B2(n14799), .ZN(
        n14824) );
  AOI21_X1 U16453 ( .B1(n14825), .B2(n14802), .A(n14824), .ZN(n14810) );
  INV_X1 U16454 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n14804) );
  OAI22_X1 U16455 ( .A1(n14823), .A2(n14805), .B1(n14804), .B2(n14803), .ZN(
        n14806) );
  INV_X1 U16456 ( .A(n14806), .ZN(n14807) );
  OAI221_X1 U16457 ( .B1(n14811), .B2(n14810), .C1(n14809), .C2(n14808), .A(
        n14807), .ZN(P2_U3265) );
  INV_X1 U16458 ( .A(n14813), .ZN(n14814) );
  AND2_X1 U16459 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14814), .ZN(P2_U3266) );
  AND2_X1 U16460 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14814), .ZN(P2_U3267) );
  INV_X1 U16461 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15239) );
  NOR2_X1 U16462 ( .A1(n14813), .A2(n15239), .ZN(P2_U3268) );
  INV_X1 U16463 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15183) );
  NOR2_X1 U16464 ( .A1(n14813), .A2(n15183), .ZN(P2_U3269) );
  AND2_X1 U16465 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14814), .ZN(P2_U3270) );
  AND2_X1 U16466 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14814), .ZN(P2_U3271) );
  AND2_X1 U16467 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14814), .ZN(P2_U3272) );
  AND2_X1 U16468 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14814), .ZN(P2_U3273) );
  AND2_X1 U16469 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14814), .ZN(P2_U3274) );
  AND2_X1 U16470 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14814), .ZN(P2_U3275) );
  AND2_X1 U16471 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14814), .ZN(P2_U3276) );
  AND2_X1 U16472 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14814), .ZN(P2_U3277) );
  AND2_X1 U16473 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14814), .ZN(P2_U3278) );
  AND2_X1 U16474 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14814), .ZN(P2_U3279) );
  AND2_X1 U16475 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14814), .ZN(P2_U3280) );
  AND2_X1 U16476 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14814), .ZN(P2_U3281) );
  AND2_X1 U16477 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14814), .ZN(P2_U3282) );
  AND2_X1 U16478 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14814), .ZN(P2_U3283) );
  AND2_X1 U16479 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14814), .ZN(P2_U3284) );
  AND2_X1 U16480 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14814), .ZN(P2_U3285) );
  AND2_X1 U16481 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14814), .ZN(P2_U3286) );
  INV_X1 U16482 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15274) );
  NOR2_X1 U16483 ( .A1(n14813), .A2(n15274), .ZN(P2_U3287) );
  AND2_X1 U16484 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14814), .ZN(P2_U3288) );
  AND2_X1 U16485 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14814), .ZN(P2_U3289) );
  AND2_X1 U16486 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14814), .ZN(P2_U3290) );
  AND2_X1 U16487 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14814), .ZN(P2_U3291) );
  INV_X1 U16488 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15167) );
  NOR2_X1 U16489 ( .A1(n14813), .A2(n15167), .ZN(P2_U3292) );
  INV_X1 U16490 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15305) );
  NOR2_X1 U16491 ( .A1(n14813), .A2(n15305), .ZN(P2_U3293) );
  AND2_X1 U16492 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14814), .ZN(P2_U3294) );
  AND2_X1 U16493 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14814), .ZN(P2_U3295) );
  AOI22_X1 U16494 ( .A1(n14817), .A2(n14816), .B1(n14815), .B2(n14820), .ZN(
        P2_U3416) );
  INV_X1 U16495 ( .A(n14818), .ZN(n14819) );
  AOI21_X1 U16496 ( .B1(n14821), .B2(n14820), .A(n14819), .ZN(P2_U3417) );
  INV_X1 U16497 ( .A(n14822), .ZN(n14848) );
  INV_X1 U16498 ( .A(n14823), .ZN(n14826) );
  AOI211_X1 U16499 ( .C1(n14848), .C2(n14826), .A(n14825), .B(n14824), .ZN(
        n14857) );
  INV_X1 U16500 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14827) );
  AOI22_X1 U16501 ( .A1(n14855), .A2(n14857), .B1(n14827), .B2(n13539), .ZN(
        P2_U3430) );
  OAI21_X1 U16502 ( .B1(n14829), .B2(n14837), .A(n14828), .ZN(n14831) );
  AOI211_X1 U16503 ( .C1(n14848), .C2(n14832), .A(n14831), .B(n14830), .ZN(
        n14858) );
  INV_X1 U16504 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15153) );
  AOI22_X1 U16505 ( .A1(n14855), .A2(n14858), .B1(n15153), .B2(n13539), .ZN(
        P2_U3436) );
  NAND2_X1 U16506 ( .A1(n14834), .A2(n14833), .ZN(n14842) );
  INV_X1 U16507 ( .A(n14835), .ZN(n14838) );
  OAI21_X1 U16508 ( .B1(n14838), .B2(n14837), .A(n14836), .ZN(n14839) );
  INV_X1 U16509 ( .A(n14839), .ZN(n14840) );
  INV_X1 U16510 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15136) );
  AOI22_X1 U16511 ( .A1(n14855), .A2(n14859), .B1(n15136), .B2(n13539), .ZN(
        P2_U3448) );
  NAND2_X1 U16512 ( .A1(n14844), .A2(n14843), .ZN(n14845) );
  AND2_X1 U16513 ( .A1(n14846), .A2(n14845), .ZN(n14852) );
  NAND2_X1 U16514 ( .A1(n14849), .A2(n14847), .ZN(n14851) );
  NAND2_X1 U16515 ( .A1(n14849), .A2(n14848), .ZN(n14850) );
  INV_X1 U16516 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14854) );
  AOI22_X1 U16517 ( .A1(n14855), .A2(n14860), .B1(n14854), .B2(n13539), .ZN(
        P2_U3463) );
  AOI22_X1 U16518 ( .A1(n14861), .A2(n14857), .B1(n14856), .B2(n13449), .ZN(
        P2_U3499) );
  AOI22_X1 U16519 ( .A1(n14861), .A2(n14858), .B1(n9226), .B2(n13449), .ZN(
        P2_U3501) );
  AOI22_X1 U16520 ( .A1(n14861), .A2(n14859), .B1(n9263), .B2(n13449), .ZN(
        P2_U3505) );
  AOI22_X1 U16521 ( .A1(n14861), .A2(n14860), .B1(n15083), .B2(n13449), .ZN(
        P2_U3510) );
  NOR2_X1 U16522 ( .A1(P3_U3897), .A2(n14862), .ZN(P3_U3150) );
  AOI21_X1 U16523 ( .B1(n8686), .B2(n14864), .A(n14863), .ZN(n14879) );
  OAI22_X1 U16524 ( .A1(n14885), .A2(n14866), .B1(n14865), .B2(n14883), .ZN(
        n14876) );
  AOI21_X1 U16525 ( .B1(n14869), .B2(n14868), .A(n14867), .ZN(n14874) );
  AOI21_X1 U16526 ( .B1(n8687), .B2(n14871), .A(n14870), .ZN(n14872) );
  OAI22_X1 U16527 ( .A1(n14874), .A2(n14873), .B1(n14872), .B2(n14897), .ZN(
        n14875) );
  NOR3_X1 U16528 ( .A1(n14877), .A2(n14876), .A3(n14875), .ZN(n14878) );
  OAI21_X1 U16529 ( .B1(n14879), .B2(n14903), .A(n14878), .ZN(P3_U3193) );
  AOI21_X1 U16530 ( .B1(n8716), .B2(n14881), .A(n14880), .ZN(n14904) );
  OAI22_X1 U16531 ( .A1(n14885), .A2(n6828), .B1(n14884), .B2(n14883), .ZN(
        n14900) );
  AOI21_X1 U16532 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n14898) );
  INV_X1 U16533 ( .A(n14889), .ZN(n14895) );
  AOI21_X1 U16534 ( .B1(n14892), .B2(n14891), .A(n14890), .ZN(n14894) );
  OAI21_X1 U16535 ( .B1(n14895), .B2(n14894), .A(n14893), .ZN(n14896) );
  OAI21_X1 U16536 ( .B1(n14898), .B2(n14897), .A(n14896), .ZN(n14899) );
  NOR3_X1 U16537 ( .A1(n14901), .A2(n14900), .A3(n14899), .ZN(n14902) );
  OAI21_X1 U16538 ( .B1(n14904), .B2(n14903), .A(n14902), .ZN(P3_U3195) );
  INV_X1 U16539 ( .A(n14939), .ZN(n14916) );
  XNOR2_X1 U16540 ( .A(n14905), .B(n14908), .ZN(n14974) );
  INV_X1 U16541 ( .A(n14974), .ZN(n14915) );
  NOR2_X1 U16542 ( .A1(n14907), .A2(n14906), .ZN(n14909) );
  XNOR2_X1 U16543 ( .A(n14909), .B(n14908), .ZN(n14913) );
  AOI22_X1 U16544 ( .A1(n14946), .A2(n14911), .B1(n14910), .B2(n14944), .ZN(
        n14912) );
  OAI21_X1 U16545 ( .B1(n14913), .B2(n14949), .A(n14912), .ZN(n14914) );
  AOI21_X1 U16546 ( .B1(n14974), .B2(n14978), .A(n14914), .ZN(n14976) );
  OAI21_X1 U16547 ( .B1(n14916), .B2(n14915), .A(n14976), .ZN(n14917) );
  MUX2_X1 U16548 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n14917), .S(n14955), .Z(
        n14918) );
  AOI21_X1 U16549 ( .B1(n14919), .B2(n14973), .A(n14918), .ZN(n14920) );
  OAI21_X1 U16550 ( .B1(n14921), .B2(n14926), .A(n14920), .ZN(P3_U3229) );
  XNOR2_X1 U16551 ( .A(n14923), .B(n8924), .ZN(n14937) );
  INV_X1 U16552 ( .A(n14937), .ZN(n14964) );
  NOR2_X1 U16553 ( .A1(n14924), .A2(n15013), .ZN(n14963) );
  INV_X1 U16554 ( .A(n14963), .ZN(n14928) );
  OAI22_X1 U16555 ( .A1(n14928), .A2(n14927), .B1(n14926), .B2(n14925), .ZN(
        n14938) );
  XNOR2_X1 U16556 ( .A(n14929), .B(n8924), .ZN(n14935) );
  OAI22_X1 U16557 ( .A1(n8522), .A2(n14932), .B1(n14931), .B2(n14930), .ZN(
        n14933) );
  AOI21_X1 U16558 ( .B1(n14935), .B2(n14934), .A(n14933), .ZN(n14936) );
  OAI21_X1 U16559 ( .B1(n14937), .B2(n14967), .A(n14936), .ZN(n14962) );
  AOI211_X1 U16560 ( .C1(n14939), .C2(n14964), .A(n14938), .B(n14962), .ZN(
        n14940) );
  AOI22_X1 U16561 ( .A1(n14957), .A2(n9086), .B1(n14940), .B2(n14955), .ZN(
        P3_U3231) );
  NOR2_X1 U16562 ( .A1(n14941), .A2(n15013), .ZN(n14959) );
  XNOR2_X1 U16563 ( .A(n9983), .B(n14942), .ZN(n14950) );
  XNOR2_X1 U16564 ( .A(n9983), .B(n14943), .ZN(n14960) );
  NAND2_X1 U16565 ( .A1(n14960), .A2(n14978), .ZN(n14948) );
  AOI22_X1 U16566 ( .A1(n14946), .A2(n8921), .B1(n14945), .B2(n14944), .ZN(
        n14947) );
  OAI211_X1 U16567 ( .C1(n14950), .C2(n14949), .A(n14948), .B(n14947), .ZN(
        n14958) );
  AOI21_X1 U16568 ( .B1(n14959), .B2(n14951), .A(n14958), .ZN(n14956) );
  AOI22_X1 U16569 ( .A1(n14960), .A2(n14953), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n14952), .ZN(n14954) );
  OAI221_X1 U16570 ( .B1(n14957), .B2(n14956), .C1(n14955), .C2(n9034), .A(
        n14954), .ZN(P3_U3232) );
  AOI211_X1 U16571 ( .C1(n14992), .C2(n14960), .A(n14959), .B(n14958), .ZN(
        n15020) );
  INV_X1 U16572 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n14961) );
  AOI22_X1 U16573 ( .A1(n15019), .A2(n15020), .B1(n14961), .B2(n15018), .ZN(
        P3_U3393) );
  AOI211_X1 U16574 ( .C1(n14964), .C2(n14992), .A(n14963), .B(n14962), .ZN(
        n15021) );
  INV_X1 U16575 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n14965) );
  AOI22_X1 U16576 ( .A1(n15019), .A2(n15021), .B1(n14965), .B2(n15018), .ZN(
        P3_U3396) );
  AOI21_X1 U16577 ( .B1(n14967), .B2(n15006), .A(n14966), .ZN(n14970) );
  INV_X1 U16578 ( .A(n14968), .ZN(n14969) );
  AOI211_X1 U16579 ( .C1(n14980), .C2(n14971), .A(n14970), .B(n14969), .ZN(
        n15022) );
  INV_X1 U16580 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U16581 ( .A1(n15019), .A2(n15022), .B1(n14972), .B2(n15018), .ZN(
        P3_U3399) );
  AOI22_X1 U16582 ( .A1(n14974), .A2(n14992), .B1(n14980), .B2(n14973), .ZN(
        n14975) );
  AND2_X1 U16583 ( .A1(n14976), .A2(n14975), .ZN(n15023) );
  INV_X1 U16584 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n14977) );
  AOI22_X1 U16585 ( .A1(n15019), .A2(n15023), .B1(n14977), .B2(n15018), .ZN(
        P3_U3402) );
  NAND2_X1 U16586 ( .A1(n14979), .A2(n14992), .ZN(n14984) );
  NAND2_X1 U16587 ( .A1(n14979), .A2(n14978), .ZN(n14983) );
  NAND2_X1 U16588 ( .A1(n14981), .A2(n14980), .ZN(n14982) );
  INV_X1 U16589 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n14986) );
  AOI22_X1 U16590 ( .A1(n15019), .A2(n15024), .B1(n14986), .B2(n15018), .ZN(
        P3_U3405) );
  INV_X1 U16591 ( .A(n14987), .ZN(n14988) );
  AOI211_X1 U16592 ( .C1(n14992), .C2(n14990), .A(n14989), .B(n14988), .ZN(
        n15025) );
  INV_X1 U16593 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n14991) );
  AOI22_X1 U16594 ( .A1(n15019), .A2(n15025), .B1(n14991), .B2(n15018), .ZN(
        P3_U3408) );
  AND2_X1 U16595 ( .A1(n14993), .A2(n14992), .ZN(n14996) );
  NOR2_X1 U16596 ( .A1(n14994), .A2(n15013), .ZN(n14995) );
  NOR3_X1 U16597 ( .A1(n14997), .A2(n14996), .A3(n14995), .ZN(n15026) );
  INV_X1 U16598 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n14998) );
  AOI22_X1 U16599 ( .A1(n15019), .A2(n15026), .B1(n14998), .B2(n15018), .ZN(
        P3_U3411) );
  OAI21_X1 U16600 ( .B1(n15000), .B2(n15006), .A(n14999), .ZN(n15001) );
  NOR2_X1 U16601 ( .A1(n15002), .A2(n15001), .ZN(n15027) );
  INV_X1 U16602 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15003) );
  AOI22_X1 U16603 ( .A1(n15019), .A2(n15027), .B1(n15003), .B2(n15018), .ZN(
        P3_U3414) );
  INV_X1 U16604 ( .A(n15004), .ZN(n15007) );
  OAI21_X1 U16605 ( .B1(n15007), .B2(n15006), .A(n15005), .ZN(n15008) );
  NOR2_X1 U16606 ( .A1(n15009), .A2(n15008), .ZN(n15028) );
  INV_X1 U16607 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15010) );
  AOI22_X1 U16608 ( .A1(n15019), .A2(n15028), .B1(n15010), .B2(n15018), .ZN(
        P3_U3417) );
  AND2_X1 U16609 ( .A1(n15012), .A2(n15011), .ZN(n15017) );
  NOR2_X1 U16610 ( .A1(n15014), .A2(n15013), .ZN(n15016) );
  NOR3_X1 U16611 ( .A1(n15017), .A2(n15016), .A3(n15015), .ZN(n15030) );
  AOI22_X1 U16612 ( .A1(n15019), .A2(n15030), .B1(n8657), .B2(n15018), .ZN(
        P3_U3420) );
  AOI22_X1 U16613 ( .A1(n15031), .A2(n15020), .B1(n9033), .B2(n15029), .ZN(
        P3_U3460) );
  AOI22_X1 U16614 ( .A1(n15031), .A2(n15021), .B1(n9070), .B2(n15029), .ZN(
        P3_U3461) );
  AOI22_X1 U16615 ( .A1(n15031), .A2(n15022), .B1(n9044), .B2(n15029), .ZN(
        P3_U3462) );
  AOI22_X1 U16616 ( .A1(n15031), .A2(n15023), .B1(n9073), .B2(n15029), .ZN(
        P3_U3463) );
  AOI22_X1 U16617 ( .A1(n15031), .A2(n15024), .B1(n9053), .B2(n15029), .ZN(
        P3_U3464) );
  AOI22_X1 U16618 ( .A1(n15031), .A2(n15025), .B1(n9057), .B2(n15029), .ZN(
        P3_U3465) );
  AOI22_X1 U16619 ( .A1(n15031), .A2(n15026), .B1(n10034), .B2(n15029), .ZN(
        P3_U3466) );
  AOI22_X1 U16620 ( .A1(n15031), .A2(n15027), .B1(n10136), .B2(n15029), .ZN(
        P3_U3467) );
  AOI22_X1 U16621 ( .A1(n15031), .A2(n15028), .B1(n10472), .B2(n15029), .ZN(
        P3_U3468) );
  AOI22_X1 U16622 ( .A1(n15031), .A2(n15030), .B1(n10715), .B2(n15029), .ZN(
        P3_U3469) );
  NOR2_X1 U16623 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n15205), .ZN(n15042) );
  NOR2_X1 U16624 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n15151), .ZN(n15033) );
  NAND4_X1 U16625 ( .A1(n15033), .A2(n15032), .A3(P3_ADDR_REG_7__SCAN_IN), 
        .A4(n15108), .ZN(n15039) );
  NOR4_X1 U16626 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .A3(P3_D_REG_12__SCAN_IN), .A4(P3_DATAO_REG_11__SCAN_IN), .ZN(n15037)
         );
  NOR4_X1 U16627 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_DATAO_REG_16__SCAN_IN), 
        .A3(P3_REG1_REG_31__SCAN_IN), .A4(P3_ADDR_REG_10__SCAN_IN), .ZN(n15036) );
  NOR4_X1 U16628 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(P2_REG1_REG_8__SCAN_IN), 
        .A3(P2_REG0_REG_6__SCAN_IN), .A4(P2_REG0_REG_2__SCAN_IN), .ZN(n15035)
         );
  NOR4_X1 U16629 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(SI_4_), .A3(
        P3_IR_REG_5__SCAN_IN), .A4(P3_REG2_REG_10__SCAN_IN), .ZN(n15034) );
  NAND4_X1 U16630 ( .A1(n15037), .A2(n15036), .A3(n15035), .A4(n15034), .ZN(
        n15038) );
  NOR4_X1 U16631 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(P3_ADDR_REG_4__SCAN_IN), 
        .A3(n15039), .A4(n15038), .ZN(n15040) );
  NAND4_X1 U16632 ( .A1(n15041), .A2(n15042), .A3(n15043), .A4(n15040), .ZN(
        n15075) );
  NOR4_X1 U16633 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(P3_IR_REG_30__SCAN_IN), 
        .A3(P3_REG0_REG_14__SCAN_IN), .A4(P3_REG1_REG_22__SCAN_IN), .ZN(n15047) );
  NOR4_X1 U16634 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .A3(P1_DATAO_REG_12__SCAN_IN), .A4(P2_REG2_REG_26__SCAN_IN), .ZN(
        n15046) );
  NOR4_X1 U16635 ( .A1(SI_8_), .A2(P3_REG3_REG_22__SCAN_IN), .A3(
        P3_ADDR_REG_16__SCAN_IN), .A4(P1_U3086), .ZN(n15045) );
  NOR4_X1 U16636 ( .A1(SI_12_), .A2(P3_REG2_REG_13__SCAN_IN), .A3(
        P3_REG2_REG_12__SCAN_IN), .A4(P3_REG2_REG_11__SCAN_IN), .ZN(n15044) );
  NAND4_X1 U16637 ( .A1(n15047), .A2(n15046), .A3(n15045), .A4(n15044), .ZN(
        n15074) );
  NOR4_X1 U16638 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_REG2_REG_21__SCAN_IN), 
        .A3(P1_REG1_REG_20__SCAN_IN), .A4(P1_REG1_REG_19__SCAN_IN), .ZN(n15051) );
  NOR4_X1 U16639 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(P1_REG1_REG_26__SCAN_IN), 
        .A3(P1_REG0_REG_23__SCAN_IN), .A4(P1_REG1_REG_22__SCAN_IN), .ZN(n15050) );
  NOR4_X1 U16640 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(P1_REG0_REG_6__SCAN_IN), 
        .A3(P1_REG1_REG_1__SCAN_IN), .A4(P1_ADDR_REG_14__SCAN_IN), .ZN(n15049)
         );
  NOR4_X1 U16641 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_1__SCAN_IN), .ZN(n15048) );
  NAND4_X1 U16642 ( .A1(n15051), .A2(n15050), .A3(n15049), .A4(n15048), .ZN(
        n15073) );
  NAND4_X1 U16643 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_REG1_REG_22__SCAN_IN), 
        .A3(P2_REG1_REG_21__SCAN_IN), .A4(P2_REG2_REG_29__SCAN_IN), .ZN(n15055) );
  NAND4_X1 U16644 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), 
        .A3(P3_REG0_REG_0__SCAN_IN), .A4(P3_REG2_REG_0__SCAN_IN), .ZN(n15054)
         );
  NAND4_X1 U16645 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_DATAO_REG_2__SCAN_IN), .A4(P2_REG0_REG_7__SCAN_IN), .ZN(n15053) );
  NAND4_X1 U16646 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .A3(P2_REG0_REG_20__SCAN_IN), .A4(P2_REG0_REG_19__SCAN_IN), .ZN(n15052) );
  NOR4_X1 U16647 ( .A1(n15055), .A2(n15054), .A3(n15053), .A4(n15052), .ZN(
        n15071) );
  NAND4_X1 U16648 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P1_B_REG_SCAN_IN), .A3(
        P1_REG3_REG_18__SCAN_IN), .A4(P3_DATAO_REG_2__SCAN_IN), .ZN(n15059) );
  NAND4_X1 U16649 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(P3_DATAO_REG_24__SCAN_IN), .A3(n15214), .A4(n15086), .ZN(n15058) );
  NAND4_X1 U16650 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(P1_DATAO_REG_6__SCAN_IN), 
        .A3(P3_IR_REG_8__SCAN_IN), .A4(P3_IR_REG_26__SCAN_IN), .ZN(n15057) );
  NAND4_X1 U16651 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), 
        .A3(P3_REG0_REG_26__SCAN_IN), .A4(P1_REG3_REG_15__SCAN_IN), .ZN(n15056) );
  NOR4_X1 U16652 ( .A1(n15059), .A2(n15058), .A3(n15057), .A4(n15056), .ZN(
        n15070) );
  NAND4_X1 U16653 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .A3(P3_ADDR_REG_12__SCAN_IN), .A4(P3_ADDR_REG_9__SCAN_IN), .ZN(n15063)
         );
  NAND4_X1 U16654 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), 
        .A3(P1_REG2_REG_9__SCAN_IN), .A4(P1_REG1_REG_7__SCAN_IN), .ZN(n15062)
         );
  NAND4_X1 U16655 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG1_REG_15__SCAN_IN), 
        .A3(P2_REG2_REG_14__SCAN_IN), .A4(P3_REG0_REG_13__SCAN_IN), .ZN(n15061) );
  NAND4_X1 U16656 ( .A1(SI_25_), .A2(P2_REG2_REG_15__SCAN_IN), .A3(
        P1_REG3_REG_22__SCAN_IN), .A4(P1_REG0_REG_17__SCAN_IN), .ZN(n15060) );
  NOR4_X1 U16657 ( .A1(n15063), .A2(n15062), .A3(n15061), .A4(n15060), .ZN(
        n15069) );
  NAND4_X1 U16658 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .A3(P1_REG3_REG_3__SCAN_IN), .A4(P1_REG1_REG_31__SCAN_IN), .ZN(n15067)
         );
  NAND4_X1 U16659 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(P2_REG1_REG_9__SCAN_IN), 
        .A3(P2_REG1_REG_2__SCAN_IN), .A4(P1_REG0_REG_25__SCAN_IN), .ZN(n15066)
         );
  NAND4_X1 U16660 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(P3_REG3_REG_23__SCAN_IN), .A3(P3_REG0_REG_23__SCAN_IN), .A4(P3_REG2_REG_15__SCAN_IN), .ZN(n15065) );
  NAND4_X1 U16661 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(
        P2_DATAO_REG_14__SCAN_IN), .A3(SI_31_), .A4(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n15064) );
  NOR4_X1 U16662 ( .A1(n15067), .A2(n15066), .A3(n15065), .A4(n15064), .ZN(
        n15068) );
  NAND4_X1 U16663 ( .A1(n15071), .A2(n15070), .A3(n15069), .A4(n15068), .ZN(
        n15072) );
  NOR4_X1 U16664 ( .A1(n15075), .A2(n15074), .A3(n15073), .A4(n15072), .ZN(
        n15325) );
  AOI221_X1 U16665 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n7702), .C2(n15076), .A(P3_RD_REG_SCAN_IN), .ZN(n15323) );
  AOI22_X1 U16666 ( .A1(n15079), .A2(keyinput68), .B1(keyinput78), .B2(n15078), 
        .ZN(n15077) );
  OAI221_X1 U16667 ( .B1(n15079), .B2(keyinput68), .C1(n15078), .C2(keyinput78), .A(n15077), .ZN(n15090) );
  AOI22_X1 U16668 ( .A1(P1_U3086), .A2(keyinput73), .B1(keyinput29), .B2(
        n13973), .ZN(n15080) );
  OAI221_X1 U16669 ( .B1(P1_U3086), .B2(keyinput73), .C1(n13973), .C2(
        keyinput29), .A(n15080), .ZN(n15089) );
  AOI22_X1 U16670 ( .A1(n15083), .A2(keyinput24), .B1(keyinput89), .B2(n15082), 
        .ZN(n15081) );
  OAI221_X1 U16671 ( .B1(n15083), .B2(keyinput24), .C1(n15082), .C2(keyinput89), .A(n15081), .ZN(n15088) );
  AOI22_X1 U16672 ( .A1(n15086), .A2(keyinput7), .B1(n15085), .B2(keyinput120), 
        .ZN(n15084) );
  OAI221_X1 U16673 ( .B1(n15086), .B2(keyinput7), .C1(n15085), .C2(keyinput120), .A(n15084), .ZN(n15087) );
  NOR4_X1 U16674 ( .A1(n15090), .A2(n15089), .A3(n15088), .A4(n15087), .ZN(
        n15134) );
  AOI22_X1 U16675 ( .A1(n8524), .A2(keyinput98), .B1(n15092), .B2(keyinput32), 
        .ZN(n15091) );
  OAI221_X1 U16676 ( .B1(n8524), .B2(keyinput98), .C1(n15092), .C2(keyinput32), 
        .A(n15091), .ZN(n15102) );
  XNOR2_X1 U16677 ( .A(n15093), .B(keyinput1), .ZN(n15101) );
  XNOR2_X1 U16678 ( .A(n15094), .B(keyinput2), .ZN(n15100) );
  XNOR2_X1 U16679 ( .A(P3_IR_REG_25__SCAN_IN), .B(keyinput93), .ZN(n15098) );
  XNOR2_X1 U16680 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput19), .ZN(n15097) );
  XNOR2_X1 U16681 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput77), .ZN(n15096) );
  XNOR2_X1 U16682 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput17), .ZN(n15095) );
  NAND4_X1 U16683 ( .A1(n15098), .A2(n15097), .A3(n15096), .A4(n15095), .ZN(
        n15099) );
  NOR4_X1 U16684 ( .A1(n15102), .A2(n15101), .A3(n15100), .A4(n15099), .ZN(
        n15133) );
  AOI22_X1 U16685 ( .A1(n15104), .A2(keyinput30), .B1(n8686), .B2(keyinput67), 
        .ZN(n15103) );
  OAI221_X1 U16686 ( .B1(n15104), .B2(keyinput30), .C1(n8686), .C2(keyinput67), 
        .A(n15103), .ZN(n15114) );
  AOI22_X1 U16687 ( .A1(n9426), .A2(keyinput64), .B1(n15106), .B2(keyinput45), 
        .ZN(n15105) );
  OAI221_X1 U16688 ( .B1(n9426), .B2(keyinput64), .C1(n15106), .C2(keyinput45), 
        .A(n15105), .ZN(n15113) );
  AOI22_X1 U16689 ( .A1(n8717), .A2(keyinput126), .B1(keyinput100), .B2(n15108), .ZN(n15107) );
  OAI221_X1 U16690 ( .B1(n8717), .B2(keyinput126), .C1(n15108), .C2(
        keyinput100), .A(n15107), .ZN(n15112) );
  XNOR2_X1 U16691 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput124), .ZN(n15110)
         );
  XNOR2_X1 U16692 ( .A(SI_4_), .B(keyinput113), .ZN(n15109) );
  NAND2_X1 U16693 ( .A1(n15110), .A2(n15109), .ZN(n15111) );
  NOR4_X1 U16694 ( .A1(n15114), .A2(n15113), .A3(n15112), .A4(n15111), .ZN(
        n15132) );
  AOI22_X1 U16695 ( .A1(n15117), .A2(keyinput50), .B1(keyinput119), .B2(n15116), .ZN(n15115) );
  OAI221_X1 U16696 ( .B1(n15117), .B2(keyinput50), .C1(n15116), .C2(
        keyinput119), .A(n15115), .ZN(n15130) );
  INV_X1 U16697 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U16698 ( .A1(n15120), .A2(keyinput86), .B1(n15119), .B2(keyinput80), 
        .ZN(n15118) );
  OAI221_X1 U16699 ( .B1(n15120), .B2(keyinput86), .C1(n15119), .C2(keyinput80), .A(n15118), .ZN(n15129) );
  AOI22_X1 U16700 ( .A1(n15123), .A2(keyinput87), .B1(n15122), .B2(keyinput22), 
        .ZN(n15121) );
  OAI221_X1 U16701 ( .B1(n15123), .B2(keyinput87), .C1(n15122), .C2(keyinput22), .A(n15121), .ZN(n15128) );
  AOI22_X1 U16702 ( .A1(n15126), .A2(keyinput47), .B1(keyinput54), .B2(n15125), 
        .ZN(n15124) );
  OAI221_X1 U16703 ( .B1(n15126), .B2(keyinput47), .C1(n15125), .C2(keyinput54), .A(n15124), .ZN(n15127) );
  NOR4_X1 U16704 ( .A1(n15130), .A2(n15129), .A3(n15128), .A4(n15127), .ZN(
        n15131) );
  NAND4_X1 U16705 ( .A1(n15134), .A2(n15133), .A3(n15132), .A4(n15131), .ZN(
        n15321) );
  AOI22_X1 U16706 ( .A1(n14102), .A2(keyinput102), .B1(n15136), .B2(keyinput38), .ZN(n15135) );
  OAI221_X1 U16707 ( .B1(n14102), .B2(keyinput102), .C1(n15136), .C2(
        keyinput38), .A(n15135), .ZN(n15149) );
  AOI22_X1 U16708 ( .A1(n15139), .A2(keyinput123), .B1(keyinput16), .B2(n15138), .ZN(n15137) );
  OAI221_X1 U16709 ( .B1(n15139), .B2(keyinput123), .C1(n15138), .C2(
        keyinput16), .A(n15137), .ZN(n15148) );
  INV_X1 U16710 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U16711 ( .A1(n15142), .A2(keyinput0), .B1(n15141), .B2(keyinput114), 
        .ZN(n15140) );
  OAI221_X1 U16712 ( .B1(n15142), .B2(keyinput0), .C1(n15141), .C2(keyinput114), .A(n15140), .ZN(n15147) );
  INV_X1 U16713 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n15143) );
  XOR2_X1 U16714 ( .A(n15143), .B(keyinput118), .Z(n15145) );
  XNOR2_X1 U16715 ( .A(P3_IR_REG_26__SCAN_IN), .B(keyinput55), .ZN(n15144) );
  NAND2_X1 U16716 ( .A1(n15145), .A2(n15144), .ZN(n15146) );
  NOR4_X1 U16717 ( .A1(n15149), .A2(n15148), .A3(n15147), .A4(n15146), .ZN(
        n15197) );
  AOI22_X1 U16718 ( .A1(n15151), .A2(keyinput110), .B1(keyinput76), .B2(n8546), 
        .ZN(n15150) );
  OAI221_X1 U16719 ( .B1(n15151), .B2(keyinput110), .C1(n8546), .C2(keyinput76), .A(n15150), .ZN(n15162) );
  AOI22_X1 U16720 ( .A1(n15154), .A2(keyinput28), .B1(n15153), .B2(keyinput66), 
        .ZN(n15152) );
  OAI221_X1 U16721 ( .B1(n15154), .B2(keyinput28), .C1(n15153), .C2(keyinput66), .A(n15152), .ZN(n15161) );
  XOR2_X1 U16722 ( .A(n15155), .B(keyinput101), .Z(n15159) );
  XNOR2_X1 U16723 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput72), .ZN(n15158)
         );
  XNOR2_X1 U16724 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput74), .ZN(n15157)
         );
  XNOR2_X1 U16725 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput13), .ZN(n15156)
         );
  NAND4_X1 U16726 ( .A1(n15159), .A2(n15158), .A3(n15157), .A4(n15156), .ZN(
        n15160) );
  NOR3_X1 U16727 ( .A1(n15162), .A2(n15161), .A3(n15160), .ZN(n15196) );
  AOI22_X1 U16728 ( .A1(n15165), .A2(keyinput8), .B1(keyinput96), .B2(n15164), 
        .ZN(n15163) );
  OAI221_X1 U16729 ( .B1(n15165), .B2(keyinput8), .C1(n15164), .C2(keyinput96), 
        .A(n15163), .ZN(n15178) );
  AOI22_X1 U16730 ( .A1(n15168), .A2(keyinput4), .B1(n15167), .B2(keyinput53), 
        .ZN(n15166) );
  OAI221_X1 U16731 ( .B1(n15168), .B2(keyinput4), .C1(n15167), .C2(keyinput53), 
        .A(n15166), .ZN(n15177) );
  AOI22_X1 U16732 ( .A1(n15171), .A2(keyinput71), .B1(keyinput12), .B2(n15170), 
        .ZN(n15169) );
  OAI221_X1 U16733 ( .B1(n15171), .B2(keyinput71), .C1(n15170), .C2(keyinput12), .A(n15169), .ZN(n15176) );
  INV_X1 U16734 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15173) );
  AOI22_X1 U16735 ( .A1(n15174), .A2(keyinput92), .B1(keyinput88), .B2(n15173), 
        .ZN(n15172) );
  OAI221_X1 U16736 ( .B1(n15174), .B2(keyinput92), .C1(n15173), .C2(keyinput88), .A(n15172), .ZN(n15175) );
  NOR4_X1 U16737 ( .A1(n15178), .A2(n15177), .A3(n15176), .A4(n15175), .ZN(
        n15195) );
  INV_X1 U16738 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n15180) );
  AOI22_X1 U16739 ( .A1(n15181), .A2(keyinput14), .B1(n15180), .B2(keyinput6), 
        .ZN(n15179) );
  OAI221_X1 U16740 ( .B1(n15181), .B2(keyinput14), .C1(n15180), .C2(keyinput6), 
        .A(n15179), .ZN(n15193) );
  AOI22_X1 U16741 ( .A1(n15183), .A2(keyinput112), .B1(keyinput97), .B2(n9959), 
        .ZN(n15182) );
  OAI221_X1 U16742 ( .B1(n15183), .B2(keyinput112), .C1(n9959), .C2(keyinput97), .A(n15182), .ZN(n15192) );
  INV_X1 U16743 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U16744 ( .A1(n15186), .A2(keyinput85), .B1(n15185), .B2(keyinput109), .ZN(n15184) );
  OAI221_X1 U16745 ( .B1(n15186), .B2(keyinput85), .C1(n15185), .C2(
        keyinput109), .A(n15184), .ZN(n15191) );
  INV_X1 U16746 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n15189) );
  AOI22_X1 U16747 ( .A1(n15189), .A2(keyinput37), .B1(keyinput103), .B2(n15188), .ZN(n15187) );
  OAI221_X1 U16748 ( .B1(n15189), .B2(keyinput37), .C1(n15188), .C2(
        keyinput103), .A(n15187), .ZN(n15190) );
  NOR4_X1 U16749 ( .A1(n15193), .A2(n15192), .A3(n15191), .A4(n15190), .ZN(
        n15194) );
  NAND4_X1 U16750 ( .A1(n15197), .A2(n15196), .A3(n15195), .A4(n15194), .ZN(
        n15320) );
  AOI22_X1 U16751 ( .A1(n15200), .A2(keyinput11), .B1(keyinput69), .B2(n15199), 
        .ZN(n15198) );
  OAI221_X1 U16752 ( .B1(n15200), .B2(keyinput11), .C1(n15199), .C2(keyinput69), .A(n15198), .ZN(n15212) );
  INV_X1 U16753 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n15202) );
  AOI22_X1 U16754 ( .A1(n15203), .A2(keyinput90), .B1(keyinput79), .B2(n15202), 
        .ZN(n15201) );
  OAI221_X1 U16755 ( .B1(n15203), .B2(keyinput90), .C1(n15202), .C2(keyinput79), .A(n15201), .ZN(n15211) );
  AOI22_X1 U16756 ( .A1(n15206), .A2(keyinput105), .B1(n15205), .B2(keyinput18), .ZN(n15204) );
  OAI221_X1 U16757 ( .B1(n15206), .B2(keyinput105), .C1(n15205), .C2(
        keyinput18), .A(n15204), .ZN(n15210) );
  XNOR2_X1 U16758 ( .A(P3_REG2_REG_12__SCAN_IN), .B(keyinput81), .ZN(n15208)
         );
  XNOR2_X1 U16759 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput21), .ZN(n15207) );
  NAND2_X1 U16760 ( .A1(n15208), .A2(n15207), .ZN(n15209) );
  NOR4_X1 U16761 ( .A1(n15212), .A2(n15211), .A3(n15210), .A4(n15209), .ZN(
        n15254) );
  AOI22_X1 U16762 ( .A1(n15214), .A2(keyinput65), .B1(keyinput20), .B2(n10631), 
        .ZN(n15213) );
  OAI221_X1 U16763 ( .B1(n15214), .B2(keyinput65), .C1(n10631), .C2(keyinput20), .A(n15213), .ZN(n15223) );
  AOI22_X1 U16764 ( .A1(n15216), .A2(keyinput60), .B1(keyinput56), .B2(n10716), 
        .ZN(n15215) );
  OAI221_X1 U16765 ( .B1(n15216), .B2(keyinput60), .C1(n10716), .C2(keyinput56), .A(n15215), .ZN(n15222) );
  AOI22_X1 U16766 ( .A1(n15218), .A2(keyinput27), .B1(n12675), .B2(keyinput106), .ZN(n15217) );
  OAI221_X1 U16767 ( .B1(n15218), .B2(keyinput27), .C1(n12675), .C2(
        keyinput106), .A(n15217), .ZN(n15221) );
  AOI22_X1 U16768 ( .A1(n8093), .A2(keyinput70), .B1(n9226), .B2(keyinput58), 
        .ZN(n15219) );
  OAI221_X1 U16769 ( .B1(n8093), .B2(keyinput70), .C1(n9226), .C2(keyinput58), 
        .A(n15219), .ZN(n15220) );
  NOR4_X1 U16770 ( .A1(n15223), .A2(n15222), .A3(n15221), .A4(n15220), .ZN(
        n15253) );
  AOI22_X1 U16771 ( .A1(n15226), .A2(keyinput48), .B1(n15225), .B2(keyinput116), .ZN(n15224) );
  OAI221_X1 U16772 ( .B1(n15226), .B2(keyinput48), .C1(n15225), .C2(
        keyinput116), .A(n15224), .ZN(n15237) );
  AOI22_X1 U16773 ( .A1(n15228), .A2(keyinput63), .B1(n9164), .B2(keyinput26), 
        .ZN(n15227) );
  OAI221_X1 U16774 ( .B1(n15228), .B2(keyinput63), .C1(n9164), .C2(keyinput26), 
        .A(n15227), .ZN(n15236) );
  AOI22_X1 U16775 ( .A1(n15231), .A2(keyinput15), .B1(keyinput95), .B2(n15230), 
        .ZN(n15229) );
  OAI221_X1 U16776 ( .B1(n15231), .B2(keyinput15), .C1(n15230), .C2(keyinput95), .A(n15229), .ZN(n15235) );
  XOR2_X1 U16777 ( .A(n7820), .B(keyinput82), .Z(n15233) );
  XNOR2_X1 U16778 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput36), .ZN(n15232)
         );
  NAND2_X1 U16779 ( .A1(n15233), .A2(n15232), .ZN(n15234) );
  NOR4_X1 U16780 ( .A1(n15237), .A2(n15236), .A3(n15235), .A4(n15234), .ZN(
        n15252) );
  AOI22_X1 U16781 ( .A1(n15240), .A2(keyinput108), .B1(n15239), .B2(keyinput9), 
        .ZN(n15238) );
  OAI221_X1 U16782 ( .B1(n15240), .B2(keyinput108), .C1(n15239), .C2(keyinput9), .A(n15238), .ZN(n15250) );
  AOI22_X1 U16783 ( .A1(n8500), .A2(keyinput84), .B1(keyinput42), .B2(n10384), 
        .ZN(n15241) );
  OAI221_X1 U16784 ( .B1(n8500), .B2(keyinput84), .C1(n10384), .C2(keyinput42), 
        .A(n15241), .ZN(n15249) );
  AOI22_X1 U16785 ( .A1(n15244), .A2(keyinput62), .B1(keyinput40), .B2(n15243), 
        .ZN(n15242) );
  OAI221_X1 U16786 ( .B1(n15244), .B2(keyinput62), .C1(n15243), .C2(keyinput40), .A(n15242), .ZN(n15248) );
  AOI22_X1 U16787 ( .A1(n15246), .A2(keyinput49), .B1(n12676), .B2(keyinput111), .ZN(n15245) );
  OAI221_X1 U16788 ( .B1(n15246), .B2(keyinput49), .C1(n12676), .C2(
        keyinput111), .A(n15245), .ZN(n15247) );
  NOR4_X1 U16789 ( .A1(n15250), .A2(n15249), .A3(n15248), .A4(n15247), .ZN(
        n15251) );
  NAND4_X1 U16790 ( .A1(n15254), .A2(n15253), .A3(n15252), .A4(n15251), .ZN(
        n15319) );
  INV_X1 U16791 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n15256) );
  AOI22_X1 U16792 ( .A1(n15256), .A2(keyinput57), .B1(keyinput94), .B2(n13257), 
        .ZN(n15255) );
  OAI221_X1 U16793 ( .B1(n15256), .B2(keyinput57), .C1(n13257), .C2(keyinput94), .A(n15255), .ZN(n15260) );
  XOR2_X1 U16794 ( .A(P3_IR_REG_5__SCAN_IN), .B(keyinput23), .Z(n15259) );
  XNOR2_X1 U16795 ( .A(n15257), .B(keyinput43), .ZN(n15258) );
  OR3_X1 U16796 ( .A1(n15260), .A2(n15259), .A3(n15258), .ZN(n15269) );
  AOI22_X1 U16797 ( .A1(n15263), .A2(keyinput107), .B1(n15262), .B2(keyinput91), .ZN(n15261) );
  OAI221_X1 U16798 ( .B1(n15263), .B2(keyinput107), .C1(n15262), .C2(
        keyinput91), .A(n15261), .ZN(n15268) );
  AOI22_X1 U16799 ( .A1(n15266), .A2(keyinput34), .B1(keyinput117), .B2(n15265), .ZN(n15264) );
  OAI221_X1 U16800 ( .B1(n15266), .B2(keyinput34), .C1(n15265), .C2(
        keyinput117), .A(n15264), .ZN(n15267) );
  NOR3_X1 U16801 ( .A1(n15269), .A2(n15268), .A3(n15267), .ZN(n15317) );
  AOI22_X1 U16802 ( .A1(n15272), .A2(keyinput10), .B1(keyinput5), .B2(n15271), 
        .ZN(n15270) );
  OAI221_X1 U16803 ( .B1(n15272), .B2(keyinput10), .C1(n15271), .C2(keyinput5), 
        .A(n15270), .ZN(n15282) );
  AOI22_X1 U16804 ( .A1(n15275), .A2(keyinput3), .B1(n15274), .B2(keyinput127), 
        .ZN(n15273) );
  OAI221_X1 U16805 ( .B1(n15275), .B2(keyinput3), .C1(n15274), .C2(keyinput127), .A(n15273), .ZN(n15281) );
  XOR2_X1 U16806 ( .A(n7947), .B(keyinput75), .Z(n15279) );
  XNOR2_X1 U16807 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput33), .ZN(n15278)
         );
  XNOR2_X1 U16808 ( .A(P2_REG1_REG_22__SCAN_IN), .B(keyinput25), .ZN(n15277)
         );
  XNOR2_X1 U16809 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput52), .ZN(n15276) );
  NAND4_X1 U16810 ( .A1(n15279), .A2(n15278), .A3(n15277), .A4(n15276), .ZN(
        n15280) );
  NOR3_X1 U16811 ( .A1(n15282), .A2(n15281), .A3(n15280), .ZN(n15316) );
  INV_X1 U16812 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15284) );
  AOI22_X1 U16813 ( .A1(n15285), .A2(keyinput61), .B1(keyinput44), .B2(n15284), 
        .ZN(n15283) );
  OAI221_X1 U16814 ( .B1(n15285), .B2(keyinput61), .C1(n15284), .C2(keyinput44), .A(n15283), .ZN(n15288) );
  INV_X1 U16815 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n15286) );
  XNOR2_X1 U16816 ( .A(n15286), .B(keyinput31), .ZN(n15287) );
  NOR2_X1 U16817 ( .A1(n15288), .A2(n15287), .ZN(n15300) );
  AOI22_X1 U16818 ( .A1(n15291), .A2(keyinput122), .B1(keyinput115), .B2(
        n15290), .ZN(n15289) );
  OAI221_X1 U16819 ( .B1(n15291), .B2(keyinput122), .C1(n15290), .C2(
        keyinput115), .A(n15289), .ZN(n15292) );
  INV_X1 U16820 ( .A(n15292), .ZN(n15299) );
  AOI22_X1 U16821 ( .A1(n15295), .A2(keyinput41), .B1(keyinput59), .B2(n15294), 
        .ZN(n15293) );
  OAI221_X1 U16822 ( .B1(n15295), .B2(keyinput41), .C1(n15294), .C2(keyinput59), .A(n15293), .ZN(n15296) );
  INV_X1 U16823 ( .A(n15296), .ZN(n15298) );
  XNOR2_X1 U16824 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput51), .ZN(n15297) );
  AND4_X1 U16825 ( .A1(n15300), .A2(n15299), .A3(n15298), .A4(n15297), .ZN(
        n15315) );
  AOI22_X1 U16826 ( .A1(n15302), .A2(keyinput99), .B1(keyinput104), .B2(n8716), 
        .ZN(n15301) );
  OAI221_X1 U16827 ( .B1(n15302), .B2(keyinput99), .C1(n8716), .C2(keyinput104), .A(n15301), .ZN(n15313) );
  AOI22_X1 U16828 ( .A1(n15305), .A2(keyinput35), .B1(keyinput46), .B2(n15304), 
        .ZN(n15303) );
  OAI221_X1 U16829 ( .B1(n15305), .B2(keyinput35), .C1(n15304), .C2(keyinput46), .A(n15303), .ZN(n15312) );
  AOI22_X1 U16830 ( .A1(n15307), .A2(keyinput39), .B1(n9176), .B2(keyinput83), 
        .ZN(n15306) );
  OAI221_X1 U16831 ( .B1(n15307), .B2(keyinput39), .C1(n9176), .C2(keyinput83), 
        .A(n15306), .ZN(n15311) );
  XNOR2_X1 U16832 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput121), .ZN(n15309) );
  XNOR2_X1 U16833 ( .A(P1_REG1_REG_19__SCAN_IN), .B(keyinput125), .ZN(n15308)
         );
  NAND2_X1 U16834 ( .A1(n15309), .A2(n15308), .ZN(n15310) );
  NOR4_X1 U16835 ( .A1(n15313), .A2(n15312), .A3(n15311), .A4(n15310), .ZN(
        n15314) );
  NAND4_X1 U16836 ( .A1(n15317), .A2(n15316), .A3(n15315), .A4(n15314), .ZN(
        n15318) );
  NOR4_X1 U16837 ( .A1(n15321), .A2(n15320), .A3(n15319), .A4(n15318), .ZN(
        n15322) );
  XOR2_X1 U16838 ( .A(n15323), .B(n15322), .Z(n15324) );
  XNOR2_X1 U16839 ( .A(n15325), .B(n15324), .ZN(U29) );
  OAI21_X1 U16840 ( .B1(n15328), .B2(n15327), .A(n15326), .ZN(SUB_1596_U58) );
  AOI21_X1 U16841 ( .B1(n15331), .B2(n15330), .A(n15329), .ZN(SUB_1596_U59) );
  XOR2_X1 U16842 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15332), .Z(SUB_1596_U53) );
  AOI21_X1 U16843 ( .B1(n15335), .B2(n15334), .A(n15333), .ZN(SUB_1596_U56) );
  INV_X1 U16844 ( .A(n15338), .ZN(n15337) );
  OAI222_X1 U16845 ( .A1(n15340), .A2(n15339), .B1(n15340), .B2(n15338), .C1(
        n15337), .C2(n15336), .ZN(SUB_1596_U60) );
  AOI21_X1 U16846 ( .B1(n15343), .B2(n15342), .A(n15341), .ZN(SUB_1596_U5) );
  OR2_X1 U10666 ( .A1(n8430), .A2(n8429), .ZN(n8432) );
  CLKBUF_X1 U7272 ( .A(n9346), .Z(n10495) );
  INV_X2 U7284 ( .A(n13740), .ZN(n10343) );
  CLKBUF_X1 U7289 ( .A(n8540), .Z(n6538) );
  NAND2_X1 U7301 ( .A1(n6516), .A2(n7041), .ZN(n8490) );
  CLKBUF_X1 U7308 ( .A(n7865), .Z(n8277) );
  NAND2_X2 U7347 ( .A1(n13873), .A2(n14306), .ZN(n7759) );
  INV_X1 U8418 ( .A(n6967), .ZN(n9343) );
  CLKBUF_X1 U9419 ( .A(n12354), .Z(n6525) );
  CLKBUF_X2 U9915 ( .A(n7678), .Z(n11569) );
endmodule

