

module b21_C_AntiSAT_k_128_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192;

  INV_X4 U4822 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U4823 ( .A1(n8403), .A2(n8281), .ZN(n8287) );
  XNOR2_X1 U4824 ( .A(n5525), .B(n5524), .ZN(n7879) );
  XNOR2_X1 U4825 ( .A(n5463), .B(n5462), .ZN(n7796) );
  INV_X2 U4826 ( .A(n4322), .ZN(n8300) );
  NAND2_X1 U4827 ( .A1(n6206), .A2(n9883), .ZN(n8143) );
  CLKBUF_X2 U4828 ( .A(n6741), .Z(n7937) );
  CLKBUF_X2 U4829 ( .A(n5923), .Z(n4319) );
  INV_X1 U4830 ( .A(n5366), .ZN(n5466) );
  OR3_X1 U4831 ( .A1(n6171), .A2(n4863), .A3(P2_IR_REG_29__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U4832 ( .A1(n6159), .A2(n6158), .ZN(n6171) );
  INV_X1 U4833 ( .A(n5923), .ZN(n5808) );
  INV_X1 U4834 ( .A(n7832), .ZN(n7641) );
  INV_X2 U4835 ( .A(n5808), .ZN(n8199) );
  NAND2_X1 U4836 ( .A1(n9253), .A2(n4603), .ZN(n9215) );
  NAND2_X1 U4837 ( .A1(n7004), .A2(n7003), .ZN(n7072) );
  NAND2_X1 U4838 ( .A1(n7832), .A2(n6173), .ZN(n7977) );
  BUF_X1 U4839 ( .A(n5836), .Z(n6006) );
  INV_X1 U4840 ( .A(n5367), .ZN(n5332) );
  AND3_X1 U4841 ( .A1(n5323), .A2(n5322), .A3(n5321), .ZN(n9697) );
  INV_X1 U4842 ( .A(n6876), .ZN(n6797) );
  INV_X1 U4843 ( .A(n6172), .ZN(n6286) );
  INV_X1 U4845 ( .A(n7144), .ZN(n4531) );
  XOR2_X1 U4846 ( .A(n8752), .B(n4322), .Z(n4318) );
  AOI21_X4 U4847 ( .B1(n9215), .B2(n9216), .A(n9222), .ZN(n9219) );
  NAND2_X2 U4848 ( .A1(n5108), .A2(n5076), .ZN(n5366) );
  OAI21_X2 U4849 ( .B1(n8963), .B2(n4700), .A(n4697), .ZN(n8898) );
  NAND2_X2 U4850 ( .A1(n5963), .A2(n8837), .ZN(n8963) );
  NOR2_X2 U4851 ( .A1(n6084), .A2(n6083), .ZN(n4488) );
  OAI211_X2 U4852 ( .C1(n6748), .C2(n7977), .A(n6747), .B(n6746), .ZN(n7048)
         );
  NAND2_X2 U4853 ( .A1(n4411), .A2(n4410), .ZN(n6172) );
  AOI21_X2 U4854 ( .B1(n7606), .B2(n7605), .A(n7604), .ZN(n7738) );
  XNOR2_X2 U4855 ( .A(n4627), .B(n5073), .ZN(n5076) );
  NAND2_X2 U4856 ( .A1(n4628), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4627) );
  AOI22_X2 U4857 ( .A1(n8357), .A2(n8355), .B1(n8295), .B2(n8354), .ZN(n8428)
         );
  AND2_X1 U4858 ( .A1(n5801), .A2(n6150), .ZN(n5923) );
  OAI21_X4 U4859 ( .B1(n6202), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6197) );
  NAND2_X2 U4860 ( .A1(n5560), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U4861 ( .A1(n8292), .A2(n8291), .ZN(n8294) );
  NAND2_X1 U4862 ( .A1(n5981), .A2(n8900), .ZN(n8940) );
  MUX2_X1 U4863 ( .A(n8088), .B(n8087), .S(n8126), .Z(n8098) );
  NAND2_X1 U4864 ( .A1(n8014), .A2(n8012), .ZN(n8149) );
  NAND2_X1 U4865 ( .A1(n8447), .A2(n9894), .ZN(n8006) );
  OR2_X1 U4866 ( .A1(n6897), .A2(n6896), .ZN(n6894) );
  AND2_X1 U4867 ( .A1(n5358), .A2(n5704), .ZN(n7167) );
  INV_X2 U4868 ( .A(n5815), .ZN(n6037) );
  NAND2_X2 U4869 ( .A1(n5809), .A2(n8192), .ZN(n5815) );
  INV_X2 U4870 ( .A(n7040), .ZN(n9894) );
  OR2_X1 U4871 ( .A1(n6725), .A2(n6724), .ZN(n6726) );
  NAND2_X2 U4872 ( .A1(n5805), .A2(n6150), .ZN(n6035) );
  INV_X1 U4873 ( .A(n9820), .ZN(n6928) );
  INV_X1 U4874 ( .A(n7048), .ZN(n6933) );
  INV_X1 U4875 ( .A(n5823), .ZN(n5347) );
  INV_X2 U4876 ( .A(n6206), .ZN(n6883) );
  NAND4_X1 U4877 ( .A1(n5441), .A2(n5440), .A3(n5439), .A4(n5438), .ZN(n8985)
         );
  INV_X1 U4878 ( .A(n5357), .ZN(n8236) );
  INV_X8 U4879 ( .A(n8306), .ZN(n8301) );
  NOR2_X1 U4880 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6080) );
  INV_X1 U4881 ( .A(n8294), .ZN(n8357) );
  OAI21_X1 U4882 ( .B1(n8224), .B2(n7953), .A(n8120), .ZN(n7954) );
  AOI21_X1 U4883 ( .B1(n8500), .B2(n8501), .A(n8113), .ZN(n8226) );
  NOR2_X1 U4884 ( .A1(n9173), .A2(n9174), .ZN(n9172) );
  OR2_X1 U4885 ( .A1(n9143), .A2(n9412), .ZN(n4526) );
  NAND2_X1 U4886 ( .A1(n4651), .A2(n4650), .ZN(n8576) );
  CLKBUF_X1 U4887 ( .A(n8366), .Z(n4405) );
  NAND2_X2 U4888 ( .A1(n5527), .A2(n5526), .ZN(n9225) );
  NAND2_X1 U4889 ( .A1(n8256), .A2(n8255), .ZN(n8366) );
  NAND2_X1 U4890 ( .A1(n9266), .A2(n9249), .ZN(n9244) );
  NAND2_X1 U4891 ( .A1(n7858), .A2(n7857), .ZN(n8759) );
  AOI21_X1 U4892 ( .B1(n4561), .B2(n4560), .A(n4559), .ZN(n5638) );
  NAND2_X1 U4893 ( .A1(n7676), .A2(n7675), .ZN(n8707) );
  OAI21_X1 U4894 ( .B1(n8047), .B2(n8046), .A(n8045), .ZN(n8050) );
  NAND2_X1 U4895 ( .A1(n4600), .A2(n4598), .ZN(n9494) );
  NAND2_X1 U4896 ( .A1(n7824), .A2(n7823), .ZN(n8777) );
  AND2_X1 U4897 ( .A1(n4587), .A2(n7230), .ZN(n7717) );
  NAND2_X1 U4898 ( .A1(n9502), .A2(n5768), .ZN(n9503) );
  NAND2_X1 U4899 ( .A1(n7225), .A2(n8022), .ZN(n7357) );
  NAND2_X1 U4900 ( .A1(n4655), .A2(n4654), .ZN(n7225) );
  NAND2_X1 U4901 ( .A1(n5213), .A2(n5212), .ZN(n9387) );
  NAND2_X1 U4902 ( .A1(n7190), .A2(n4656), .ZN(n4655) );
  NAND2_X1 U4903 ( .A1(n7508), .A2(n7507), .ZN(n8803) );
  OR2_X1 U4904 ( .A1(n8016), .A2(n4492), .ZN(n4489) );
  NAND2_X1 U4905 ( .A1(n4409), .A2(n5273), .ZN(n9561) );
  NAND2_X1 U4906 ( .A1(n7060), .A2(n7059), .ZN(n7350) );
  NAND2_X1 U4907 ( .A1(n9815), .A2(n4741), .ZN(n9814) );
  NAND2_X1 U4908 ( .A1(n5589), .A2(n5706), .ZN(n7524) );
  AOI21_X1 U4909 ( .B1(n6886), .B2(n4852), .A(n4851), .ZN(n4850) );
  NAND2_X1 U4910 ( .A1(n7014), .A2(n7013), .ZN(n7282) );
  NAND2_X1 U4911 ( .A1(n6194), .A2(n8144), .ZN(n6805) );
  INV_X2 U4912 ( .A(n5836), .ZN(n8195) );
  CLKBUF_X1 U4913 ( .A(n5769), .Z(n6687) );
  NAND2_X1 U4914 ( .A1(n6883), .A2(n6998), .ZN(n6236) );
  NAND4_X2 U4915 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n8987)
         );
  NAND4_X1 U4916 ( .A1(n6166), .A2(n6165), .A3(n6164), .A4(n6163), .ZN(n9820)
         );
  AND3_X1 U4917 ( .A1(n6189), .A2(n6188), .A3(n6187), .ZN(n6899) );
  AND2_X1 U4918 ( .A1(n6178), .A2(n6177), .ZN(n6181) );
  INV_X1 U4919 ( .A(n6998), .ZN(n9883) );
  NOR2_X1 U4920 ( .A1(n6998), .A2(n6990), .ZN(n6989) );
  OAI211_X1 U4921 ( .C1(n6736), .C2(n7977), .A(n6735), .B(n6734), .ZN(n9825)
         );
  CLKBUF_X3 U4922 ( .A(n5344), .Z(n4320) );
  INV_X1 U4923 ( .A(n8308), .ZN(n4321) );
  CLKBUF_X3 U4924 ( .A(n8308), .Z(n4322) );
  AOI21_X1 U4925 ( .B1(n4805), .B2(n4980), .A(n4801), .ZN(n4800) );
  NAND2_X1 U4926 ( .A1(n6162), .A2(n4667), .ZN(n4666) );
  XNOR2_X1 U4927 ( .A(n5699), .B(n5698), .ZN(n7164) );
  NAND2_X1 U4928 ( .A1(n6721), .A2(n6720), .ZN(n8308) );
  NAND2_X1 U4929 ( .A1(n5559), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5699) );
  AND2_X2 U4930 ( .A1(n5076), .A2(n8244), .ZN(n5350) );
  INV_X1 U4931 ( .A(n6907), .ZN(n6839) );
  NAND2_X4 U4932 ( .A1(n7832), .A2(n6304), .ZN(n6907) );
  AND2_X1 U4933 ( .A1(n4676), .A2(n4674), .ZN(n5786) );
  NAND2_X1 U4934 ( .A1(n6161), .A2(n4323), .ZN(n8833) );
  XNOR2_X1 U4935 ( .A(n5074), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U4936 ( .A1(n5495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5558) );
  AND2_X1 U4937 ( .A1(n7128), .A2(n7982), .ZN(n8178) );
  MUX2_X1 U4938 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6169), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n6170) );
  XNOR2_X1 U4939 ( .A(n4506), .B(n6199), .ZN(n7260) );
  NAND2_X2 U4940 ( .A1(n6286), .A2(P2_U3152), .ZN(n8830) );
  INV_X2 U4941 ( .A(n6286), .ZN(n5052) );
  INV_X4 U4942 ( .A(n6286), .ZN(n6304) );
  NOR2_X1 U4943 ( .A1(n6200), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6085) );
  OAI21_X1 U4944 ( .B1(n4911), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n4808), .ZN(
        n6173) );
  NOR2_X1 U4945 ( .A1(n4856), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4855) );
  NAND2_X1 U4946 ( .A1(n5060), .A2(n4844), .ZN(n4843) );
  NAND2_X1 U4947 ( .A1(n6100), .A2(n4857), .ZN(n4856) );
  NOR2_X1 U4948 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5056) );
  NOR2_X1 U4949 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4838) );
  NOR2_X1 U4950 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5057) );
  NOR2_X1 U4951 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4620) );
  INV_X1 U4952 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4844) );
  NOR2_X1 U4953 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4578) );
  NOR2_X1 U4954 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5744) );
  INV_X1 U4955 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6335) );
  INV_X1 U4956 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5060) );
  INV_X1 U4957 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4522) );
  INV_X4 U4958 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4959 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6100) );
  NOR2_X2 U4960 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5361) );
  INV_X1 U4961 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5428) );
  INV_X1 U4962 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4518) );
  AOI211_X2 U4963 ( .C1(n7377), .C2(n7376), .A(n5606), .B(n5605), .ZN(n5612)
         );
  AOI21_X2 U4964 ( .B1(n8548), .B2(n8528), .A(n8520), .ZN(n8531) );
  NAND2_X2 U4965 ( .A1(n7951), .A2(n8540), .ZN(n8548) );
  OAI22_X2 U4966 ( .A1(n8248), .A2(n4846), .B1(n8246), .B2(n4845), .ZN(n8365)
         );
  NOR3_X2 U4967 ( .A1(n8631), .A2(n8759), .A3(n4594), .ZN(n4592) );
  NAND2_X1 U4968 ( .A1(n5356), .A2(n6286), .ZN(n5344) );
  NOR2_X2 U4969 ( .A1(n8531), .A2(n7952), .ZN(n8510) );
  XNOR2_X2 U4970 ( .A(n6197), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6234) );
  INV_X4 U4971 ( .A(n6035), .ZN(n8192) );
  NAND2_X1 U4972 ( .A1(n4760), .A2(n4759), .ZN(n5091) );
  AOI21_X1 U4973 ( .B1(n4762), .B2(n4764), .A(n4400), .ZN(n4759) );
  NAND2_X1 U4974 ( .A1(n5129), .A2(n4762), .ZN(n4760) );
  NOR2_X1 U4975 ( .A1(n4960), .A2(n4773), .ZN(n4772) );
  INV_X1 U4976 ( .A(n5252), .ZN(n4960) );
  NAND2_X1 U4977 ( .A1(n4497), .A2(n7128), .ZN(n4496) );
  AOI21_X1 U4978 ( .B1(n4477), .B2(n4476), .A(n4366), .ZN(n4475) );
  INV_X1 U4979 ( .A(n4481), .ZN(n4476) );
  AND2_X1 U4980 ( .A1(n4872), .A2(n4871), .ZN(n4327) );
  INV_X1 U4981 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4872) );
  INV_X1 U4982 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4871) );
  NOR2_X2 U4983 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6174) );
  INV_X1 U4984 ( .A(n4423), .ZN(n4422) );
  OR2_X1 U4985 ( .A1(n9320), .A2(n9321), .ZN(n9299) );
  NAND2_X1 U4986 ( .A1(n5035), .A2(n5034), .ZN(n5129) );
  NAND2_X1 U4987 ( .A1(n4789), .A2(n4787), .ZN(n5035) );
  AOI21_X1 U4988 ( .B1(n4790), .B2(n4383), .A(n4788), .ZN(n4787) );
  AND2_X1 U4989 ( .A1(n4985), .A2(n4984), .ZN(n5177) );
  NAND2_X1 U4990 ( .A1(n4965), .A2(n4964), .ZN(n5234) );
  XNOR2_X1 U4991 ( .A(n4958), .B(SI_11_), .ZN(n5252) );
  NAND2_X1 U4992 ( .A1(n4952), .A2(n4951), .ZN(n5268) );
  INV_X1 U4993 ( .A(n4666), .ZN(n6741) );
  INV_X1 U4994 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6079) );
  INV_X1 U4995 ( .A(n7977), .ZN(n7969) );
  NAND2_X1 U4996 ( .A1(n4373), .A2(n4328), .ZN(n4480) );
  NAND2_X1 U4997 ( .A1(n8530), .A2(n4485), .ZN(n4483) );
  AOI21_X1 U4998 ( .B1(n4423), .B2(n4421), .A(n4420), .ZN(n4419) );
  INV_X1 U4999 ( .A(n4424), .ZN(n4421) );
  INV_X1 U5000 ( .A(n9096), .ZN(n4420) );
  AND2_X1 U5001 ( .A1(n8647), .A2(n8062), .ZN(n4505) );
  INV_X1 U5002 ( .A(n7502), .ZN(n4900) );
  INV_X1 U5003 ( .A(n7260), .ZN(n8173) );
  AOI21_X1 U5004 ( .B1(n4736), .B2(n4734), .A(n4364), .ZN(n4733) );
  INV_X1 U5005 ( .A(n4738), .ZN(n4734) );
  INV_X1 U5006 ( .A(n4736), .ZN(n4735) );
  OR2_X1 U5007 ( .A1(n8797), .A2(n7800), .ZN(n8051) );
  NAND2_X1 U5008 ( .A1(n4642), .A2(n4640), .ZN(n7676) );
  NOR2_X1 U5009 ( .A1(n4643), .A2(n4641), .ZN(n4640) );
  AND2_X1 U5010 ( .A1(n8040), .A2(n7987), .ZN(n8042) );
  INV_X1 U5011 ( .A(n7569), .ZN(n4591) );
  NOR2_X1 U5012 ( .A1(n7191), .A2(n4657), .ZN(n4656) );
  INV_X1 U5013 ( .A(n8014), .ZN(n4657) );
  INV_X1 U5014 ( .A(n8987), .ZN(n5814) );
  NAND2_X1 U5015 ( .A1(n5953), .A2(n7705), .ZN(n5959) );
  NAND2_X1 U5016 ( .A1(n8186), .A2(n5771), .ZN(n5682) );
  NOR2_X1 U5017 ( .A1(n9434), .A2(n4542), .ZN(n4541) );
  OR2_X1 U5018 ( .A1(n9434), .A2(n9100), .ZN(n9131) );
  OR2_X1 U5019 ( .A1(n9225), .A2(n9239), .ZN(n9096) );
  OR2_X1 U5020 ( .A1(n5471), .A2(n5457), .ZN(n5517) );
  OR2_X1 U5021 ( .A1(n9467), .A2(n9472), .ZN(n4536) );
  NOR2_X1 U5022 ( .A1(n9089), .A2(n4832), .ZN(n4831) );
  NOR2_X1 U5023 ( .A1(n9338), .A2(n9323), .ZN(n9089) );
  INV_X1 U5024 ( .A(n9086), .ZN(n4832) );
  NAND2_X1 U5025 ( .A1(n6684), .A2(n5806), .ZN(n5836) );
  OR2_X1 U5026 ( .A1(n8980), .A2(n9703), .ZN(n7605) );
  OR2_X1 U5027 ( .A1(n8985), .A2(n5848), .ZN(n5706) );
  AND2_X1 U5028 ( .A1(n7267), .A2(n7266), .ZN(n4837) );
  INV_X1 U5029 ( .A(n7274), .ZN(n7267) );
  AND2_X1 U5030 ( .A1(n8987), .A2(n7144), .ZN(n6683) );
  INV_X1 U5031 ( .A(n4791), .ZN(n4790) );
  OAI21_X1 U5032 ( .B1(n4794), .B2(n4383), .A(n5029), .ZN(n4791) );
  AND2_X1 U5033 ( .A1(n5005), .A2(n5004), .ZN(n5475) );
  XNOR2_X1 U5034 ( .A(n4988), .B(SI_17_), .ZN(n5160) );
  OAI21_X1 U5035 ( .B1(n4557), .B2(n4553), .A(n4945), .ZN(n4552) );
  NAND2_X1 U5036 ( .A1(n4558), .A2(n4347), .ZN(n4553) );
  XNOR2_X1 U5037 ( .A(n4321), .B(n9825), .ZN(n4870) );
  NOR2_X1 U5038 ( .A1(n4878), .A2(n4343), .ZN(n4877) );
  NAND2_X1 U5039 ( .A1(n4849), .A2(n4847), .ZN(n6905) );
  AOI21_X1 U5040 ( .B1(n4850), .B2(n4853), .A(n4848), .ZN(n4847) );
  INV_X1 U5041 ( .A(n6861), .ZN(n4848) );
  OR2_X1 U5042 ( .A1(n8135), .A2(n7985), .ZN(n4639) );
  OR2_X1 U5043 ( .A1(n8491), .A2(n7979), .ZN(n8131) );
  NAND2_X1 U5044 ( .A1(n4494), .A2(n4402), .ZN(n4493) );
  INV_X1 U5045 ( .A(n9584), .ZN(n8491) );
  OR2_X1 U5046 ( .A1(n8224), .A2(n4648), .ZN(n7968) );
  NAND2_X1 U5047 ( .A1(n8121), .A2(n4649), .ZN(n4648) );
  NAND2_X1 U5048 ( .A1(n7939), .A2(n7938), .ZN(n8719) );
  NAND2_X1 U5049 ( .A1(n8108), .A2(n7915), .ZN(n8509) );
  INV_X1 U5050 ( .A(n4750), .ZN(n8521) );
  AOI21_X1 U5051 ( .B1(n4753), .B2(n8164), .A(n7891), .ZN(n4751) );
  INV_X1 U5052 ( .A(n4753), .ZN(n4752) );
  NAND2_X1 U5053 ( .A1(n7950), .A2(n4652), .ZN(n4651) );
  NOR2_X1 U5054 ( .A1(n8594), .A2(n4653), .ZN(n4652) );
  INV_X1 U5055 ( .A(n8079), .ZN(n4653) );
  OR2_X1 U5056 ( .A1(n8769), .A2(n8349), .ZN(n8079) );
  NAND2_X1 U5057 ( .A1(n8618), .A2(n7845), .ZN(n7846) );
  OR2_X1 U5058 ( .A1(n8773), .A2(n8638), .ZN(n7845) );
  OR2_X1 U5059 ( .A1(n8784), .A2(n8663), .ZN(n8063) );
  NAND2_X1 U5060 ( .A1(n8674), .A2(n8658), .ZN(n8652) );
  OR2_X1 U5061 ( .A1(n8797), .A2(n8692), .ZN(n4463) );
  NAND2_X1 U5062 ( .A1(n7556), .A2(n4644), .ZN(n4642) );
  AND2_X1 U5063 ( .A1(n8033), .A2(n8032), .ZN(n4644) );
  AOI21_X1 U5064 ( .B1(n4468), .B2(n4756), .A(n4467), .ZN(n4465) );
  OR2_X1 U5065 ( .A1(n7569), .A2(n7558), .ZN(n8032) );
  NAND2_X1 U5066 ( .A1(n4662), .A2(n4487), .ZN(n6168) );
  NOR2_X1 U5067 ( .A1(n4663), .A2(n6298), .ZN(n4662) );
  NAND2_X1 U5068 ( .A1(n4327), .A2(n4855), .ZN(n4663) );
  AND3_X1 U5069 ( .A1(n4664), .A2(n4665), .A3(n4488), .ZN(n6099) );
  AND2_X1 U5070 ( .A1(n4350), .A2(n4327), .ZN(n4664) );
  AND2_X1 U5071 ( .A1(n4665), .A2(n4516), .ZN(n4515) );
  NOR2_X1 U5072 ( .A1(n4517), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n4516) );
  NAND2_X1 U5073 ( .A1(n4522), .A2(n4518), .ZN(n4517) );
  NAND2_X1 U5074 ( .A1(n4342), .A2(n4520), .ZN(n6978) );
  INV_X1 U5075 ( .A(n4521), .ZN(n4520) );
  NAND2_X1 U5076 ( .A1(n8937), .A2(n4713), .ZN(n4712) );
  AND2_X1 U5077 ( .A1(n5995), .A2(n5994), .ZN(n8860) );
  NAND2_X1 U5078 ( .A1(n4711), .A2(n8938), .ZN(n4710) );
  INV_X1 U5079 ( .A(n8937), .ZN(n4711) );
  AND3_X1 U5080 ( .A1(n5474), .A2(n5473), .A3(n5472), .ZN(n8920) );
  CLKBUF_X2 U5081 ( .A(n5365), .Z(n5437) );
  CLKBUF_X2 U5082 ( .A(n5367), .Z(n5500) );
  AOI21_X1 U5083 ( .B1(n4821), .B2(n9107), .A(n4332), .ZN(n4818) );
  NAND2_X1 U5084 ( .A1(n5093), .A2(n5092), .ZN(n9417) );
  NOR2_X1 U5085 ( .A1(n9159), .A2(n4822), .ZN(n4821) );
  OR2_X1 U5086 ( .A1(n9243), .A2(n4422), .ZN(n4414) );
  AND2_X1 U5087 ( .A1(n4377), .A2(n4416), .ZN(n4415) );
  NAND2_X1 U5088 ( .A1(n4419), .A2(n4422), .ZN(n4416) );
  NOR2_X1 U5089 ( .A1(n9236), .A2(n4604), .ZN(n4603) );
  INV_X1 U5090 ( .A(n9127), .ZN(n4604) );
  NAND2_X1 U5091 ( .A1(n9269), .A2(n9270), .ZN(n9268) );
  NAND2_X1 U5092 ( .A1(n9294), .A2(n4432), .ZN(n4428) );
  NOR2_X1 U5093 ( .A1(n9285), .A2(n5646), .ZN(n4612) );
  INV_X1 U5094 ( .A(n9294), .ZN(n4434) );
  NAND2_X1 U5095 ( .A1(n9481), .A2(n9085), .ZN(n9086) );
  NAND2_X1 U5096 ( .A1(n9347), .A2(n9354), .ZN(n9348) );
  AOI21_X1 U5097 ( .B1(n9365), .B2(n4389), .A(n4449), .ZN(n9087) );
  NOR2_X1 U5098 ( .A1(n9372), .A2(n9084), .ZN(n4449) );
  INV_X1 U5099 ( .A(n4320), .ZN(n5496) );
  NOR2_X1 U5100 ( .A1(n4783), .A2(n5054), .ZN(n4782) );
  AND2_X1 U5101 ( .A1(n4842), .A2(n5059), .ZN(n4839) );
  NOR2_X1 U5102 ( .A1(n4344), .A2(n4843), .ZN(n4842) );
  INV_X1 U5103 ( .A(n4798), .ZN(n5178) );
  AOI21_X1 U5104 ( .B1(n4807), .B2(n4799), .A(n4802), .ZN(n4798) );
  OAI21_X1 U5105 ( .B1(n5268), .B2(n4771), .A(n4770), .ZN(n5235) );
  INV_X1 U5106 ( .A(n4769), .ZN(n5253) );
  AOI21_X1 U5107 ( .B1(n5268), .B2(n4907), .A(n4773), .ZN(n4769) );
  XNOR2_X1 U5108 ( .A(n5268), .B(n4907), .ZN(n7076) );
  NAND2_X1 U5109 ( .A1(n5401), .A2(n5400), .ZN(n4937) );
  NAND2_X1 U5110 ( .A1(n7918), .A2(n7917), .ZN(n8730) );
  NAND2_X1 U5111 ( .A1(n7916), .A2(n7969), .ZN(n7918) );
  XNOR2_X1 U5112 ( .A(n6737), .B(n4870), .ZN(n6925) );
  NAND2_X1 U5113 ( .A1(n7072), .A2(n7071), .ZN(n7106) );
  NOR2_X1 U5114 ( .A1(n7981), .A2(n4639), .ZN(n4629) );
  NAND2_X1 U5115 ( .A1(n7924), .A2(n7923), .ZN(n8438) );
  NAND2_X1 U5116 ( .A1(n8020), .A2(n8152), .ZN(n4492) );
  INV_X1 U5117 ( .A(n4492), .ZN(n4491) );
  NAND2_X1 U5118 ( .A1(n4641), .A2(n8126), .ZN(n4510) );
  INV_X1 U5119 ( .A(n4505), .ZN(n4504) );
  AND2_X1 U5120 ( .A1(n4502), .A2(n8069), .ZN(n4501) );
  NAND2_X1 U5121 ( .A1(n4505), .A2(n4503), .ZN(n4502) );
  NAND2_X1 U5122 ( .A1(n4335), .A2(n5639), .ZN(n4572) );
  NOR2_X1 U5123 ( .A1(n4403), .A2(n4571), .ZN(n4570) );
  AND2_X1 U5124 ( .A1(n5640), .A2(n9125), .ZN(n4571) );
  NOR2_X1 U5125 ( .A1(n5651), .A2(n5650), .ZN(n5654) );
  NAND2_X1 U5126 ( .A1(n4566), .A2(n4565), .ZN(n5651) );
  INV_X1 U5127 ( .A(n4892), .ZN(n4891) );
  OAI21_X1 U5128 ( .B1(n4894), .B2(n4893), .A(n8344), .ZN(n4892) );
  INV_X1 U5129 ( .A(n8274), .ZN(n4893) );
  AND2_X1 U5130 ( .A1(n9189), .A2(n9103), .ZN(n9134) );
  NAND2_X1 U5131 ( .A1(n4806), .A2(n4974), .ZN(n4805) );
  INV_X1 U5132 ( .A(n5191), .ZN(n4806) );
  NOR2_X1 U5133 ( .A1(n4975), .A2(n4804), .ZN(n4803) );
  INV_X1 U5134 ( .A(n4970), .ZN(n4804) );
  INV_X1 U5135 ( .A(n5207), .ZN(n4975) );
  NAND2_X1 U5136 ( .A1(n4413), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4810) );
  INV_X1 U5137 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4413) );
  NOR2_X2 U5138 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .ZN(
        n4911) );
  AND2_X1 U5139 ( .A1(n8491), .A2(n7979), .ZN(n8125) );
  INV_X1 U5140 ( .A(n8833), .ZN(n6162) );
  OR2_X1 U5141 ( .A1(n8719), .A2(n8313), .ZN(n8127) );
  OR2_X1 U5142 ( .A1(n8741), .A2(n8390), .ZN(n8107) );
  OR2_X1 U5143 ( .A1(n8745), .A2(n8562), .ZN(n7890) );
  AOI21_X1 U5144 ( .B1(n4724), .B2(n4729), .A(n8877), .ZN(n4722) );
  INV_X1 U5145 ( .A(n4724), .ZN(n4723) );
  INV_X1 U5146 ( .A(n8876), .ZN(n4720) );
  AND2_X1 U5147 ( .A1(n8868), .A2(n4694), .ZN(n4693) );
  INV_X1 U5148 ( .A(n4910), .ZN(n4694) );
  XNOR2_X1 U5149 ( .A(n5868), .B(n6006), .ZN(n7319) );
  OR2_X1 U5150 ( .A1(n9424), .A2(n8951), .ZN(n5673) );
  OR2_X1 U5151 ( .A1(n9420), .A2(n9176), .ZN(n5676) );
  NOR2_X1 U5152 ( .A1(n9424), .A2(n9106), .ZN(n4822) );
  NOR2_X1 U5153 ( .A1(n4611), .A2(n9134), .ZN(n4608) );
  OR2_X1 U5154 ( .A1(n5542), .A2(n8883), .ZN(n5544) );
  INV_X1 U5155 ( .A(n9134), .ZN(n5727) );
  OR2_X1 U5156 ( .A1(n9225), .A2(n9446), .ZN(n4542) );
  INV_X1 U5157 ( .A(n5501), .ZN(n5101) );
  OR2_X1 U5158 ( .A1(n9461), .A2(n4536), .ZN(n4535) );
  NOR2_X1 U5159 ( .A1(n9387), .A2(n9612), .ZN(n4534) );
  OR2_X1 U5160 ( .A1(n9080), .A2(n4387), .ZN(n4444) );
  NOR2_X1 U5161 ( .A1(n4444), .A2(n4441), .ZN(n4442) );
  OR2_X1 U5162 ( .A1(n9561), .A2(n8978), .ZN(n7731) );
  NAND2_X1 U5163 ( .A1(n4574), .A2(n4573), .ZN(n7737) );
  AND2_X1 U5164 ( .A1(n8979), .A2(n4346), .ZN(n4573) );
  NOR2_X1 U5165 ( .A1(n6314), .A2(n6286), .ZN(n4528) );
  NAND2_X1 U5166 ( .A1(n8236), .A2(n5823), .ZN(n5704) );
  NAND2_X1 U5167 ( .A1(n4448), .A2(n9075), .ZN(n4446) );
  AND2_X1 U5168 ( .A1(n5034), .A2(n5033), .ZN(n5137) );
  INV_X1 U5169 ( .A(n5024), .ZN(n4792) );
  NOR2_X1 U5170 ( .A1(n5025), .A2(n4795), .ZN(n4794) );
  INV_X1 U5171 ( .A(n5020), .ZN(n4795) );
  XNOR2_X1 U5172 ( .A(n4993), .B(SI_18_), .ZN(n5148) );
  OAI21_X1 U5173 ( .B1(n5161), .B2(n4991), .A(n4990), .ZN(n5149) );
  INV_X1 U5174 ( .A(n5160), .ZN(n4991) );
  AOI21_X1 U5175 ( .B1(n5268), .B2(n4352), .A(n4766), .ZN(n4765) );
  NAND2_X1 U5176 ( .A1(n4767), .A2(n4965), .ZN(n4766) );
  NAND2_X1 U5177 ( .A1(n4947), .A2(n4946), .ZN(n4951) );
  OAI21_X1 U5178 ( .B1(n4558), .B2(n4936), .A(n4940), .ZN(n4557) );
  NAND2_X1 U5179 ( .A1(n6912), .A2(n6911), .ZN(n7199) );
  INV_X1 U5180 ( .A(n4884), .ZN(n4883) );
  OAI21_X1 U5181 ( .B1(n4886), .B2(n4885), .A(n8412), .ZN(n4884) );
  INV_X1 U5182 ( .A(n8260), .ZN(n4885) );
  INV_X1 U5183 ( .A(n8365), .ZN(n8256) );
  NAND2_X1 U5184 ( .A1(n6371), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7896) );
  INV_X1 U5185 ( .A(n8338), .ZN(n8269) );
  NAND2_X1 U5186 ( .A1(n7473), .A2(n7472), .ZN(n7503) );
  INV_X1 U5187 ( .A(n7239), .ZN(n4874) );
  INV_X1 U5188 ( .A(n6859), .ZN(n4851) );
  INV_X1 U5189 ( .A(n6848), .ZN(n4852) );
  INV_X1 U5190 ( .A(n6886), .ZN(n4853) );
  AND2_X1 U5191 ( .A1(n7638), .A2(n4897), .ZN(n4896) );
  NAND2_X1 U5192 ( .A1(n4898), .A2(n7475), .ZN(n4897) );
  INV_X1 U5193 ( .A(n6738), .ZN(n7875) );
  OR2_X1 U5194 ( .A1(n6318), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U5195 ( .A1(n4477), .A2(n8225), .ZN(n4474) );
  OAI21_X1 U5196 ( .B1(n4475), .B2(n4472), .A(n4370), .ZN(n4471) );
  AND2_X1 U5197 ( .A1(n7931), .A2(n7930), .ZN(n8314) );
  AND2_X1 U5198 ( .A1(n4328), .A2(n4485), .ZN(n4481) );
  NAND2_X1 U5199 ( .A1(n4486), .A2(n8390), .ZN(n4485) );
  AND2_X1 U5200 ( .A1(n8107), .A2(n8094), .ZN(n8530) );
  OR2_X1 U5201 ( .A1(n8571), .A2(n8392), .ZN(n4902) );
  NOR2_X1 U5202 ( .A1(n8540), .A2(n4754), .ZN(n4753) );
  INV_X1 U5203 ( .A(n4902), .ZN(n4754) );
  AOI21_X1 U5204 ( .B1(n8575), .B2(n8162), .A(n4452), .ZN(n8565) );
  NOR2_X1 U5205 ( .A1(n8759), .A2(n8596), .ZN(n4452) );
  INV_X1 U5206 ( .A(n7850), .ZN(n6369) );
  AND2_X1 U5207 ( .A1(n8080), .A2(n8578), .ZN(n4650) );
  NOR2_X1 U5208 ( .A1(n7855), .A2(n4739), .ZN(n4738) );
  INV_X1 U5209 ( .A(n4903), .ZN(n4739) );
  NAND2_X1 U5210 ( .A1(n4737), .A2(n4740), .ZN(n4736) );
  INV_X1 U5211 ( .A(n8603), .ZN(n4737) );
  OR2_X1 U5212 ( .A1(n4597), .A2(n8607), .ZN(n4903) );
  NOR2_X1 U5213 ( .A1(n8649), .A2(n8777), .ZN(n7829) );
  AND2_X1 U5214 ( .A1(n4338), .A2(n8063), .ZN(n4661) );
  NAND2_X1 U5215 ( .A1(n7948), .A2(n7947), .ZN(n8648) );
  NOR2_X1 U5216 ( .A1(n4362), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U5217 ( .A1(n8648), .A2(n8647), .ZN(n8646) );
  NOR2_X1 U5218 ( .A1(n7807), .A2(n8647), .ZN(n4747) );
  AOI21_X1 U5219 ( .B1(n8684), .B2(n4461), .A(n4359), .ZN(n4460) );
  OR2_X1 U5220 ( .A1(n8667), .A2(n8666), .ZN(n4749) );
  NAND2_X1 U5221 ( .A1(n4743), .A2(n4329), .ZN(n4464) );
  AOI21_X1 U5222 ( .B1(n4324), .B2(n8042), .A(n4358), .ZN(n4742) );
  OR2_X1 U5223 ( .A1(n7714), .A2(n8042), .ZN(n4744) );
  AND2_X1 U5224 ( .A1(n8048), .A2(n8706), .ZN(n8045) );
  INV_X1 U5225 ( .A(n8045), .ZN(n7669) );
  NAND2_X1 U5226 ( .A1(n7358), .A2(n8029), .ZN(n7556) );
  INV_X1 U5227 ( .A(n8442), .ZN(n7558) );
  INV_X1 U5228 ( .A(n8440), .ZN(n7678) );
  INV_X1 U5229 ( .A(n8441), .ZN(n7555) );
  NAND2_X1 U5230 ( .A1(n7357), .A2(n8027), .ZN(n7358) );
  AND2_X1 U5231 ( .A1(n8032), .A2(n8031), .ZN(n8154) );
  NAND2_X1 U5232 ( .A1(n7222), .A2(n7226), .ZN(n7352) );
  NAND2_X1 U5233 ( .A1(n7217), .A2(n8150), .ZN(n7216) );
  NAND2_X1 U5234 ( .A1(n6942), .A2(n6941), .ZN(n7190) );
  INV_X1 U5235 ( .A(n9819), .ZN(n7033) );
  INV_X1 U5236 ( .A(n8446), .ZN(n7182) );
  AND2_X1 U5237 ( .A1(n6276), .A2(n6205), .ZN(n9818) );
  INV_X1 U5238 ( .A(n9873), .ZN(n6597) );
  AND2_X1 U5239 ( .A1(n6262), .A2(n6227), .ZN(n6763) );
  NAND2_X1 U5240 ( .A1(n4469), .A2(n4475), .ZN(n8218) );
  OR2_X1 U5241 ( .A1(n8521), .A2(n4478), .ZN(n4469) );
  NAND2_X1 U5242 ( .A1(n7906), .A2(n7905), .ZN(n8737) );
  NAND2_X1 U5243 ( .A1(n7628), .A2(n7627), .ZN(n8797) );
  AOI22_X1 U5244 ( .A1(n6171), .A2(n4862), .B1(n4860), .B2(n4859), .ZN(n4858)
         );
  NAND2_X1 U5245 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4861), .ZN(n4860) );
  NAND2_X1 U5246 ( .A1(n6099), .A2(n4854), .ZN(n6167) );
  INV_X1 U5247 ( .A(n4856), .ZN(n4854) );
  NOR2_X1 U5248 ( .A1(n4521), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n4519) );
  INV_X1 U5249 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6078) );
  NOR2_X1 U5250 ( .A1(n6319), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U5251 ( .A1(n5099), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5186) );
  INV_X1 U5252 ( .A(n5200), .ZN(n5099) );
  INV_X1 U5253 ( .A(n4703), .ZN(n4701) );
  OR2_X1 U5254 ( .A1(n8960), .A2(n8961), .ZN(n4704) );
  NAND2_X1 U5255 ( .A1(n6068), .A2(n6070), .ZN(n6069) );
  NOR2_X1 U5256 ( .A1(n5817), .A2(n5816), .ZN(n6130) );
  INV_X1 U5257 ( .A(n4710), .ZN(n4709) );
  AND2_X1 U5258 ( .A1(n8860), .A2(n4707), .ZN(n4706) );
  NAND2_X1 U5259 ( .A1(n4710), .A2(n4708), .ZN(n4707) );
  INV_X1 U5260 ( .A(n4688), .ZN(n4687) );
  OAI21_X1 U5261 ( .B1(n5928), .B2(n4689), .A(n5939), .ZN(n4688) );
  INV_X1 U5262 ( .A(n5934), .ZN(n4689) );
  AOI21_X1 U5263 ( .B1(n4683), .B2(n4684), .A(n4682), .ZN(n4681) );
  XNOR2_X1 U5264 ( .A(n5826), .B(n8195), .ZN(n5830) );
  XNOR2_X1 U5265 ( .A(n5837), .B(n6006), .ZN(n5843) );
  OR2_X1 U5266 ( .A1(n6125), .A2(n5792), .ZN(n7139) );
  NAND2_X1 U5267 ( .A1(n5962), .A2(n5961), .ZN(n8837) );
  AND2_X1 U5268 ( .A1(n5694), .A2(n5739), .ZN(n4757) );
  OR2_X1 U5269 ( .A1(n8186), .A2(n5771), .ZN(n5739) );
  INV_X1 U5270 ( .A(n5350), .ZN(n5484) );
  OR2_X1 U5271 ( .A1(n5484), .A2(n5417), .ZN(n5424) );
  NAND2_X1 U5272 ( .A1(n5466), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5354) );
  INV_X1 U5273 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5237) );
  OR2_X1 U5274 ( .A1(n5269), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5271) );
  AOI21_X1 U5275 ( .B1(n7415), .B2(n5214), .A(n7414), .ZN(n7578) );
  INV_X1 U5276 ( .A(n4782), .ZN(n4777) );
  AND2_X1 U5277 ( .A1(n5676), .A2(n9136), .ZN(n9159) );
  OR2_X1 U5278 ( .A1(n9166), .A2(n9107), .ZN(n4823) );
  INV_X1 U5279 ( .A(n4822), .ZN(n4820) );
  NAND2_X1 U5280 ( .A1(n9219), .A2(n9130), .ZN(n4609) );
  AND2_X1 U5281 ( .A1(n9131), .A2(n9130), .ZN(n9205) );
  OR2_X1 U5282 ( .A1(n9446), .A2(n8933), .ZN(n9216) );
  AND2_X1 U5283 ( .A1(n9096), .A2(n9097), .ZN(n9222) );
  AND2_X1 U5284 ( .A1(n4325), .A2(n9095), .ZN(n4424) );
  NAND2_X1 U5285 ( .A1(n4371), .A2(n4325), .ZN(n4423) );
  AND3_X1 U5286 ( .A1(n5461), .A2(n5460), .A3(n5459), .ZN(n9273) );
  NAND2_X1 U5287 ( .A1(n9268), .A2(n9126), .ZN(n9253) );
  NAND2_X1 U5288 ( .A1(n9261), .A2(n9093), .ZN(n9243) );
  OR2_X1 U5289 ( .A1(n5503), .A2(n5479), .ZN(n5481) );
  NAND2_X1 U5290 ( .A1(n4432), .A2(n9091), .ZN(n4431) );
  NAND2_X1 U5291 ( .A1(n4428), .A2(n4427), .ZN(n9261) );
  NOR2_X1 U5292 ( .A1(n4430), .A2(n9270), .ZN(n4427) );
  NAND2_X1 U5293 ( .A1(n9299), .A2(n9123), .ZN(n9302) );
  OR2_X1 U5294 ( .A1(n4333), .A2(n4386), .ZN(n4825) );
  NAND2_X1 U5295 ( .A1(n9087), .A2(n4826), .ZN(n4824) );
  NOR2_X1 U5296 ( .A1(n4827), .A2(n4386), .ZN(n4826) );
  AOI21_X1 U5297 ( .B1(n4833), .B2(n4831), .A(n4830), .ZN(n4829) );
  NOR2_X1 U5298 ( .A1(n9476), .A2(n9088), .ZN(n4830) );
  NAND2_X1 U5299 ( .A1(n9087), .A2(n4831), .ZN(n4828) );
  AOI21_X1 U5300 ( .B1(n4617), .B2(n4616), .A(n4615), .ZN(n4614) );
  INV_X1 U5301 ( .A(n9355), .ZN(n4833) );
  AOI21_X1 U5302 ( .B1(n9378), .B2(n9380), .A(n9082), .ZN(n9365) );
  NAND2_X1 U5303 ( .A1(n9116), .A2(n9115), .ZN(n9362) );
  AND2_X1 U5304 ( .A1(n5619), .A2(n9379), .ZN(n9399) );
  NAND2_X1 U5305 ( .A1(n5097), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5246) );
  NOR2_X2 U5306 ( .A1(n7609), .A2(n9561), .ZN(n9562) );
  INV_X1 U5307 ( .A(n4599), .ZN(n4598) );
  OAI21_X1 U5308 ( .B1(n7739), .B2(n5600), .A(n7740), .ZN(n4599) );
  INV_X1 U5309 ( .A(n9304), .ZN(n9552) );
  INV_X1 U5310 ( .A(n4836), .ZN(n4835) );
  AOI21_X1 U5311 ( .B1(n4836), .B2(n7393), .A(n4349), .ZN(n4834) );
  AND2_X1 U5312 ( .A1(n7397), .A2(n7390), .ZN(n4836) );
  NAND2_X1 U5313 ( .A1(n7345), .A2(n7344), .ZN(n7391) );
  INV_X1 U5314 ( .A(n9641), .ZN(n7384) );
  AND2_X1 U5315 ( .A1(n7341), .A2(n7340), .ZN(n7375) );
  AND2_X1 U5316 ( .A1(n7262), .A2(n7261), .ZN(n7274) );
  NAND2_X1 U5317 ( .A1(n7265), .A2(n7272), .ZN(n7523) );
  AND3_X1 U5318 ( .A1(n5435), .A2(n5434), .A3(n5433), .ZN(n5848) );
  AND2_X1 U5319 ( .A1(n7149), .A2(n7148), .ZN(n7166) );
  XNOR2_X1 U5320 ( .A(n5838), .B(n9670), .ZN(n7168) );
  INV_X1 U5321 ( .A(n9556), .ZN(n9306) );
  INV_X1 U5322 ( .A(n4451), .ZN(n4450) );
  OAI21_X1 U5323 ( .B1(n9415), .B2(n9704), .A(n4621), .ZN(n4451) );
  NAND2_X1 U5324 ( .A1(n9417), .A2(n9712), .ZN(n4621) );
  NAND2_X1 U5325 ( .A1(n5139), .A2(n5138), .ZN(n9430) );
  OR2_X1 U5326 ( .A1(n4320), .A2(n7724), .ZN(n5540) );
  NAND2_X1 U5327 ( .A1(n5498), .A2(n5497), .ZN(n9467) );
  AND3_X1 U5328 ( .A1(n5304), .A2(n5303), .A3(n5302), .ZN(n9703) );
  NAND2_X1 U5329 ( .A1(n9497), .A2(n9718), .ZN(n9708) );
  AOI21_X1 U5330 ( .B1(n4782), .B2(n5080), .A(n4399), .ZN(n4781) );
  NAND2_X1 U5331 ( .A1(n4785), .A2(n5054), .ZN(n4784) );
  INV_X1 U5332 ( .A(n5080), .ZN(n4785) );
  OR2_X1 U5333 ( .A1(n5091), .A2(n5088), .ZN(n5045) );
  XNOR2_X1 U5334 ( .A(n5081), .B(n5080), .ZN(n8216) );
  XNOR2_X1 U5335 ( .A(n5116), .B(n5115), .ZN(n7925) );
  NAND2_X1 U5336 ( .A1(n4761), .A2(n5040), .ZN(n5116) );
  NAND2_X1 U5337 ( .A1(n5129), .A2(n5128), .ZN(n4761) );
  NOR2_X1 U5338 ( .A1(n5064), .A2(n4675), .ZN(n4674) );
  OR2_X1 U5339 ( .A1(n5756), .A2(n4677), .ZN(n4676) );
  NOR2_X1 U5340 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4675) );
  OAI21_X1 U5341 ( .B1(n5454), .B2(n5453), .A(n5014), .ZN(n5513) );
  NAND2_X1 U5342 ( .A1(n5597), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5598) );
  INV_X1 U5343 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5741) );
  INV_X1 U5344 ( .A(n4714), .ZN(n4619) );
  INV_X1 U5345 ( .A(n5318), .ZN(n4558) );
  INV_X1 U5346 ( .A(n4557), .ZN(n4556) );
  NAND2_X1 U5347 ( .A1(n4933), .A2(n4932), .ZN(n5401) );
  OR2_X1 U5348 ( .A1(n5361), .A2(n9535), .ZN(n5429) );
  NAND2_X1 U5349 ( .A1(n7081), .A2(n7080), .ZN(n7569) );
  NAND2_X1 U5350 ( .A1(n7458), .A2(n7457), .ZN(n7718) );
  NAND2_X1 U5351 ( .A1(n7812), .A2(n7811), .ZN(n8784) );
  NAND2_X1 U5352 ( .A1(n4866), .A2(n4865), .ZN(n4864) );
  NAND2_X1 U5353 ( .A1(n4868), .A2(n6733), .ZN(n4869) );
  NAND2_X1 U5354 ( .A1(n7073), .A2(n4406), .ZN(n7105) );
  INV_X1 U5355 ( .A(n7101), .ZN(n4406) );
  NAND2_X1 U5356 ( .A1(n7849), .A2(n7848), .ZN(n8769) );
  INV_X1 U5357 ( .A(n7001), .ZN(n7004) );
  NAND2_X1 U5358 ( .A1(n7246), .A2(n7245), .ZN(n8041) );
  NAND2_X1 U5359 ( .A1(n6894), .A2(n6727), .ZN(n6878) );
  NAND2_X1 U5360 ( .A1(n6769), .A2(n7366), .ZN(n8421) );
  OR2_X1 U5361 ( .A1(n6768), .A2(n6759), .ZN(n8423) );
  OAI21_X1 U5362 ( .B1(n8168), .B2(n4639), .A(n4638), .ZN(n4637) );
  NAND2_X1 U5363 ( .A1(n8135), .A2(n7985), .ZN(n4638) );
  INV_X1 U5364 ( .A(n7968), .ZN(n7976) );
  AND2_X1 U5365 ( .A1(n8177), .A2(n4635), .ZN(n4634) );
  NAND2_X1 U5366 ( .A1(n8301), .A2(n7983), .ZN(n8177) );
  AOI21_X1 U5367 ( .B1(n8176), .B2(n4635), .A(n4631), .ZN(n4630) );
  INV_X1 U5368 ( .A(n8182), .ZN(n4631) );
  OR2_X1 U5369 ( .A1(n8227), .A2(n4672), .ZN(n4671) );
  NAND2_X1 U5370 ( .A1(n4388), .A2(n4673), .ZN(n4672) );
  INV_X1 U5371 ( .A(n8496), .ZN(n8221) );
  NOR2_X1 U5372 ( .A1(n8723), .A2(n8718), .ZN(n4669) );
  OR2_X1 U5373 ( .A1(n9840), .A2(n6545), .ZN(n7366) );
  NAND3_X2 U5374 ( .A1(n6183), .A2(n6184), .A3(n4454), .ZN(n6998) );
  NAND2_X1 U5375 ( .A1(n7832), .A2(n4455), .ZN(n4454) );
  OR2_X1 U5376 ( .A1(n8722), .A2(n9877), .ZN(n4458) );
  NAND2_X1 U5377 ( .A1(n8720), .A2(n9827), .ZN(n4586) );
  NAND2_X1 U5378 ( .A1(n5184), .A2(n5183), .ZN(n9481) );
  INV_X1 U5379 ( .A(n9338), .ZN(n9476) );
  NAND2_X1 U5380 ( .A1(n5456), .A2(n5455), .ZN(n9452) );
  INV_X1 U5381 ( .A(n9074), .ZN(n9507) );
  NAND2_X1 U5382 ( .A1(n5197), .A2(n5196), .ZN(n9488) );
  NAND2_X1 U5383 ( .A1(n5536), .A2(n5535), .ZN(n9239) );
  NAND4_X1 U5384 ( .A1(n5331), .A2(n5330), .A3(n5329), .A4(n5328), .ZN(n8981)
         );
  AND2_X1 U5385 ( .A1(n9003), .A2(n4408), .ZN(n6592) );
  NAND2_X1 U5386 ( .A1(n9002), .A2(n10108), .ZN(n4408) );
  NAND2_X1 U5387 ( .A1(n4818), .A2(n4817), .ZN(n4816) );
  OAI21_X1 U5388 ( .B1(n9109), .B2(n4818), .A(n4814), .ZN(n4813) );
  NAND2_X1 U5389 ( .A1(n4624), .A2(n9142), .ZN(n9416) );
  NAND2_X1 U5390 ( .A1(n4625), .A2(n9501), .ZN(n4624) );
  XNOR2_X1 U5391 ( .A(n9139), .B(n4817), .ZN(n4625) );
  NOR2_X1 U5392 ( .A1(n5071), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n4626) );
  AOI21_X1 U5393 ( .B1(n4334), .B2(n4491), .A(n4369), .ZN(n4490) );
  AND2_X1 U5394 ( .A1(n8708), .A2(n8049), .ZN(n4508) );
  INV_X1 U5395 ( .A(n8666), .ZN(n4503) );
  NAND2_X1 U5396 ( .A1(n5625), .A2(n5644), .ZN(n4563) );
  NOR2_X1 U5397 ( .A1(n5622), .A2(n5621), .ZN(n4564) );
  NOR2_X1 U5398 ( .A1(n5631), .A2(n9355), .ZN(n4560) );
  NAND2_X1 U5399 ( .A1(n4500), .A2(n4499), .ZN(n8071) );
  AOI21_X1 U5400 ( .B1(n4501), .B2(n4504), .A(n4659), .ZN(n4499) );
  NOR2_X1 U5401 ( .A1(n4568), .A2(n5642), .ZN(n4567) );
  OAI21_X1 U5402 ( .B1(n5647), .B2(n4572), .A(n4570), .ZN(n4569) );
  NAND2_X1 U5403 ( .A1(n5641), .A2(n5644), .ZN(n4568) );
  NAND2_X1 U5404 ( .A1(n5664), .A2(n5665), .ZN(n4404) );
  AOI21_X1 U5405 ( .B1(n5641), .B2(n5490), .A(n4403), .ZN(n5491) );
  NAND2_X1 U5406 ( .A1(n5679), .A2(n5681), .ZN(n5688) );
  INV_X1 U5407 ( .A(n4763), .ZN(n4762) );
  OAI21_X1 U5408 ( .B1(n5128), .B2(n4764), .A(n5115), .ZN(n4763) );
  INV_X1 U5409 ( .A(n5040), .ZN(n4764) );
  INV_X1 U5410 ( .A(n5137), .ZN(n4788) );
  NAND2_X1 U5411 ( .A1(n4997), .A2(n4996), .ZN(n5000) );
  AND2_X1 U5412 ( .A1(n4803), .A2(n4980), .ZN(n4797) );
  INV_X1 U5413 ( .A(n5177), .ZN(n4801) );
  INV_X1 U5414 ( .A(n5234), .ZN(n4768) );
  AOI21_X1 U5415 ( .B1(n4891), .B2(n4893), .A(n4355), .ZN(n4889) );
  NOR2_X1 U5416 ( .A1(n6757), .A2(n6756), .ZN(n6760) );
  AND2_X1 U5417 ( .A1(n8283), .A2(n8385), .ZN(n8289) );
  OR2_X1 U5418 ( .A1(n8737), .A2(n8109), .ZN(n8108) );
  OR2_X1 U5419 ( .A1(n8759), .A2(n8347), .ZN(n8085) );
  NAND2_X1 U5420 ( .A1(n4595), .A2(n8593), .ZN(n4594) );
  INV_X1 U5421 ( .A(n4596), .ZN(n4595) );
  NAND2_X1 U5422 ( .A1(n8615), .A2(n4597), .ZN(n4596) );
  OR2_X1 U5423 ( .A1(n7838), .A2(n6368), .ZN(n7850) );
  INV_X1 U5424 ( .A(n8054), .ZN(n4646) );
  INV_X1 U5425 ( .A(n4463), .ZN(n4461) );
  OR2_X1 U5426 ( .A1(n7510), .A2(n7509), .ZN(n7645) );
  NAND2_X1 U5427 ( .A1(n6365), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7510) );
  INV_X1 U5428 ( .A(n7476), .ZN(n6365) );
  OR2_X1 U5429 ( .A1(n7718), .A2(n7678), .ZN(n8040) );
  OR2_X1 U5430 ( .A1(n7248), .A2(n7247), .ZN(n7476) );
  INV_X1 U5431 ( .A(n8156), .ZN(n4467) );
  NAND2_X1 U5432 ( .A1(n6364), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7248) );
  INV_X1 U5433 ( .A(n7090), .ZN(n6364) );
  OR2_X1 U5434 ( .A1(n7083), .A2(n7082), .ZN(n7090) );
  OR2_X1 U5435 ( .A1(n7350), .A2(n7356), .ZN(n8027) );
  NAND2_X1 U5436 ( .A1(n6771), .A2(n9830), .ZN(n8007) );
  NAND2_X1 U5437 ( .A1(n6928), .A2(n6876), .ZN(n7999) );
  INV_X1 U5438 ( .A(n8144), .ZN(n6238) );
  NAND2_X1 U5439 ( .A1(n4863), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4861) );
  NAND2_X1 U5440 ( .A1(n8826), .A2(n4863), .ZN(n4859) );
  NOR2_X1 U5441 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(n8826), .ZN(n4862) );
  INV_X1 U5442 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U5443 ( .A1(n4810), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4808) );
  OR2_X1 U5444 ( .A1(n5880), .A2(n7297), .ZN(n5899) );
  INV_X1 U5445 ( .A(n4712), .ZN(n4708) );
  AOI21_X1 U5446 ( .B1(n4678), .B2(n5913), .A(n4679), .ZN(n4683) );
  INV_X1 U5447 ( .A(n6106), .ZN(n4679) );
  INV_X1 U5448 ( .A(n6070), .ZN(n4678) );
  INV_X1 U5449 ( .A(n6105), .ZN(n4682) );
  OR2_X1 U5450 ( .A1(n6687), .A2(n9274), .ZN(n5689) );
  INV_X1 U5451 ( .A(n4821), .ZN(n4819) );
  NAND2_X1 U5452 ( .A1(n5103), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5529) );
  INV_X1 U5453 ( .A(n4831), .ZN(n4827) );
  NOR2_X1 U5454 ( .A1(n9355), .A2(n5629), .ZN(n4617) );
  OR2_X1 U5455 ( .A1(n7610), .A2(n9711), .ZN(n7609) );
  NOR2_X1 U5456 ( .A1(n4602), .A2(n5600), .ZN(n4601) );
  INV_X1 U5457 ( .A(n7737), .ZN(n4602) );
  AND2_X1 U5458 ( .A1(n5385), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5384) );
  OR2_X1 U5459 ( .A1(n8981), .A2(n9697), .ZN(n7395) );
  AND2_X1 U5460 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5385) );
  NAND2_X1 U5461 ( .A1(n6140), .A2(n6642), .ZN(n4575) );
  NAND2_X1 U5462 ( .A1(n4576), .A2(n5539), .ZN(n4574) );
  NAND2_X1 U5463 ( .A1(n4530), .A2(n9670), .ZN(n7173) );
  INV_X1 U5464 ( .A(n7172), .ZN(n4530) );
  INV_X1 U5465 ( .A(n5051), .ZN(n4783) );
  NAND2_X1 U5466 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n4677) );
  NAND2_X1 U5467 ( .A1(n5236), .A2(n4840), .ZN(n4715) );
  INV_X1 U5468 ( .A(n4843), .ZN(n4841) );
  INV_X1 U5469 ( .A(n4805), .ZN(n4799) );
  NAND2_X1 U5470 ( .A1(n5058), .A2(n4716), .ZN(n4714) );
  NOR2_X1 U5471 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4716) );
  NAND2_X1 U5472 ( .A1(n4980), .A2(n4979), .ZN(n5191) );
  XNOR2_X1 U5473 ( .A(n4972), .B(SI_14_), .ZN(n5207) );
  NAND2_X1 U5474 ( .A1(n4967), .A2(n4966), .ZN(n4970) );
  NAND2_X1 U5475 ( .A1(n5220), .A2(n4901), .ZN(n4971) );
  INV_X1 U5476 ( .A(n4772), .ZN(n4771) );
  AOI21_X1 U5477 ( .B1(n4772), .B2(n4774), .A(n4368), .ZN(n4770) );
  INV_X1 U5478 ( .A(n4957), .ZN(n4773) );
  NOR2_X2 U5479 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5055) );
  NAND2_X1 U5480 ( .A1(n4911), .A2(n4809), .ZN(n4410) );
  INV_X1 U5481 ( .A(n4810), .ZN(n4412) );
  NOR2_X1 U5482 ( .A1(n8397), .A2(n4895), .ZN(n4894) );
  INV_X1 U5483 ( .A(n8271), .ZN(n4895) );
  OR2_X1 U5484 ( .A1(n8273), .A2(n8272), .ZN(n8274) );
  INV_X1 U5485 ( .A(n4870), .ZN(n4866) );
  INV_X1 U5486 ( .A(n6737), .ZN(n4865) );
  NOR2_X1 U5487 ( .A1(n8374), .A2(n4887), .ZN(n4886) );
  INV_X1 U5488 ( .A(n8257), .ZN(n4887) );
  AND2_X1 U5489 ( .A1(n6760), .A2(n8180), .ZN(n6770) );
  NAND2_X1 U5490 ( .A1(n4496), .A2(n8175), .ZN(n4495) );
  INV_X1 U5491 ( .A(n8183), .ZN(n4635) );
  OR3_X1 U5492 ( .A1(n6356), .A2(P2_IR_REG_10__SCAN_IN), .A3(
        P2_IR_REG_11__SCAN_IN), .ZN(n6380) );
  NOR2_X1 U5493 ( .A1(n8219), .A2(n8719), .ZN(n8490) );
  NAND2_X1 U5494 ( .A1(n8438), .A2(n9821), .ZN(n4673) );
  NAND2_X1 U5495 ( .A1(n8496), .A2(n8223), .ZN(n8219) );
  NAND2_X1 U5496 ( .A1(n8541), .A2(n4486), .ZN(n8522) );
  INV_X1 U5497 ( .A(n8530), .ZN(n8520) );
  OR2_X1 U5498 ( .A1(n7859), .A2(n6370), .ZN(n7870) );
  NAND2_X1 U5499 ( .A1(n4453), .A2(n4731), .ZN(n8575) );
  AOI21_X1 U5500 ( .B1(n4733), .B2(n4735), .A(n4336), .ZN(n4731) );
  NAND2_X1 U5501 ( .A1(n7846), .A2(n4733), .ZN(n4453) );
  NOR2_X1 U5502 ( .A1(n8631), .A2(n4596), .ZN(n8609) );
  OAI21_X1 U5503 ( .B1(n8648), .B2(n4660), .A(n4658), .ZN(n8623) );
  INV_X1 U5504 ( .A(n4661), .ZN(n4660) );
  AOI21_X1 U5505 ( .B1(n4661), .B2(n8644), .A(n4659), .ZN(n4658) );
  NOR2_X1 U5506 ( .A1(n8631), .A2(n8773), .ZN(n8619) );
  AND2_X1 U5507 ( .A1(n8078), .A2(n8602), .ZN(n8624) );
  AOI21_X1 U5508 ( .B1(n4747), .B2(n8666), .A(n4392), .ZN(n4746) );
  NAND2_X1 U5509 ( .A1(n6366), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7814) );
  INV_X1 U5510 ( .A(n7653), .ZN(n6366) );
  NAND2_X1 U5511 ( .A1(n6367), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7838) );
  INV_X1 U5512 ( .A(n7814), .ZN(n6367) );
  AOI21_X1 U5513 ( .B1(n8707), .B2(n7946), .A(n7945), .ZN(n8691) );
  NAND2_X1 U5514 ( .A1(n4582), .A2(n4581), .ZN(n8687) );
  NOR2_X1 U5515 ( .A1(n4589), .A2(n7718), .ZN(n4587) );
  NAND2_X1 U5516 ( .A1(n7230), .A2(n4345), .ZN(n7559) );
  NAND2_X1 U5517 ( .A1(n7230), .A2(n9906), .ZN(n7363) );
  NAND2_X1 U5518 ( .A1(n4655), .A2(n8019), .ZN(n7192) );
  AND2_X1 U5519 ( .A1(n8152), .A2(n8019), .ZN(n4654) );
  NAND2_X1 U5520 ( .A1(n6798), .A2(n4741), .ZN(n6801) );
  NOR2_X1 U5521 ( .A1(n9831), .A2(n7048), .ZN(n7037) );
  INV_X1 U5522 ( .A(n9825), .ZN(n9830) );
  OR2_X1 U5523 ( .A1(n9826), .A2(n9825), .ZN(n9831) );
  NAND2_X1 U5524 ( .A1(n6989), .A2(n6797), .ZN(n9826) );
  OR2_X1 U5525 ( .A1(n9915), .A2(n7982), .ZN(n6545) );
  NOR2_X1 U5526 ( .A1(n6314), .A2(n4456), .ZN(n4455) );
  INV_X1 U5527 ( .A(n6173), .ZN(n4456) );
  NAND2_X1 U5528 ( .A1(n8719), .A2(n8804), .ZN(n4585) );
  INV_X1 U5529 ( .A(n9914), .ZN(n8804) );
  OR2_X1 U5530 ( .A1(n6722), .A2(n8178), .ZN(n9914) );
  NOR2_X1 U5531 ( .A1(n6757), .A2(n6230), .ZN(n6546) );
  NAND2_X1 U5532 ( .A1(n6087), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6104) );
  INV_X1 U5533 ( .A(n6085), .ZN(n6202) );
  AND2_X1 U5534 ( .A1(n6340), .A2(n6337), .ZN(n6488) );
  INV_X1 U5535 ( .A(n4665), .ZN(n6298) );
  NOR2_X1 U5536 ( .A1(n6298), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6300) );
  INV_X1 U5537 ( .A(n6037), .ZN(n8197) );
  INV_X1 U5538 ( .A(n5805), .ZN(n5801) );
  AOI21_X1 U5539 ( .B1(n4722), .B2(n4723), .A(n4720), .ZN(n4719) );
  INV_X1 U5540 ( .A(n4722), .ZN(n4721) );
  NAND2_X1 U5541 ( .A1(n8960), .A2(n8961), .ZN(n4703) );
  NOR2_X1 U5542 ( .A1(n8908), .A2(n4725), .ZN(n4724) );
  INV_X1 U5543 ( .A(n4728), .ZN(n4725) );
  NAND2_X1 U5544 ( .A1(n8848), .A2(n4730), .ZN(n4728) );
  NAND2_X1 U5545 ( .A1(n8850), .A2(n4727), .ZN(n4726) );
  INV_X1 U5546 ( .A(n6249), .ZN(n5860) );
  AOI21_X1 U5547 ( .B1(n4693), .B2(n8917), .A(n4692), .ZN(n4691) );
  INV_X1 U5548 ( .A(n4909), .ZN(n4692) );
  NAND2_X1 U5549 ( .A1(n6128), .A2(n5822), .ZN(n6676) );
  INV_X1 U5550 ( .A(n5186), .ZN(n5100) );
  OR2_X1 U5551 ( .A1(n5171), .A2(n5154), .ZN(n5501) );
  OR2_X1 U5552 ( .A1(n5228), .A2(n5098), .ZN(n5200) );
  AOI21_X1 U5553 ( .B1(n9169), .B2(n5335), .A(n5135), .ZN(n8951) );
  AND2_X1 U5554 ( .A1(n5551), .A2(n5550), .ZN(n9100) );
  AND4_X1 U5555 ( .A1(n5159), .A2(n5158), .A3(n5157), .A4(n5156), .ZN(n8902)
         );
  AND4_X1 U5556 ( .A1(n5176), .A2(n5175), .A3(n5174), .A4(n5173), .ZN(n9323)
         );
  AOI21_X1 U5557 ( .B1(n8989), .B2(n8988), .A(n8990), .ZN(n8992) );
  NOR2_X1 U5558 ( .A1(n6515), .A2(n6623), .ZN(n6556) );
  AND2_X1 U5559 ( .A1(n6567), .A2(n6566), .ZN(n10159) );
  NOR2_X1 U5560 ( .A1(n4819), .A2(n4817), .ZN(n4812) );
  NAND2_X1 U5561 ( .A1(n4818), .A2(n4815), .ZN(n4814) );
  NAND2_X1 U5562 ( .A1(n4819), .A2(n4817), .ZN(n4815) );
  NAND2_X1 U5563 ( .A1(n9154), .A2(n9144), .ZN(n9143) );
  AOI21_X1 U5564 ( .B1(n4608), .B2(n9132), .A(n4606), .ZN(n4605) );
  INV_X1 U5565 ( .A(n4608), .ZN(n4607) );
  INV_X1 U5566 ( .A(n9133), .ZN(n4606) );
  AND2_X1 U5567 ( .A1(n5141), .A2(n5140), .ZN(n9187) );
  NAND2_X1 U5568 ( .A1(n4541), .A2(n9189), .ZN(n4540) );
  NOR2_X1 U5569 ( .A1(n9244), .A2(n4539), .ZN(n9199) );
  INV_X1 U5570 ( .A(n4541), .ZN(n4539) );
  NOR2_X1 U5571 ( .A1(n9244), .A2(n4542), .ZN(n9212) );
  INV_X1 U5572 ( .A(n5481), .ZN(n5102) );
  NOR2_X1 U5573 ( .A1(n9333), .A2(n4535), .ZN(n9280) );
  NOR2_X1 U5574 ( .A1(n9333), .A2(n4536), .ZN(n9295) );
  NAND2_X1 U5575 ( .A1(n9372), .A2(n4534), .ZN(n4533) );
  AND4_X1 U5576 ( .A1(n5190), .A2(n5189), .A3(n5188), .A4(n5187), .ZN(n9363)
         );
  AND4_X1 U5577 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n9364)
         );
  INV_X1 U5578 ( .A(n4534), .ZN(n4532) );
  INV_X1 U5579 ( .A(n4439), .ZN(n4438) );
  OAI21_X1 U5580 ( .B1(n4326), .B2(n4444), .A(n9079), .ZN(n4439) );
  OR2_X1 U5581 ( .A1(n5246), .A2(n5226), .ZN(n5228) );
  AND2_X1 U5582 ( .A1(n9562), .A2(n9507), .ZN(n9502) );
  NAND2_X1 U5583 ( .A1(n9548), .A2(n7739), .ZN(n7743) );
  NAND2_X1 U5584 ( .A1(n7738), .A2(n7737), .ZN(n9548) );
  OR2_X1 U5585 ( .A1(n6125), .A2(n6139), .ZN(n9556) );
  NOR2_X1 U5586 ( .A1(n7380), .A2(n7389), .ZN(n7400) );
  NAND2_X1 U5587 ( .A1(n5384), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5395) );
  AND3_X1 U5588 ( .A1(n5407), .A2(n5406), .A3(n5405), .ZN(n9641) );
  OR2_X1 U5589 ( .A1(n7379), .A2(n7384), .ZN(n7380) );
  AND2_X1 U5590 ( .A1(n5603), .A2(n5604), .ZN(n7376) );
  INV_X1 U5591 ( .A(n7376), .ZN(n7342) );
  NAND2_X1 U5592 ( .A1(n7375), .A2(n7342), .ZN(n7374) );
  OR2_X1 U5593 ( .A1(n7531), .A2(n7339), .ZN(n7379) );
  NAND2_X1 U5594 ( .A1(n5706), .A2(n5586), .ZN(n7153) );
  AND2_X1 U5595 ( .A1(n5346), .A2(n4527), .ZN(n4529) );
  NAND2_X1 U5596 ( .A1(n8236), .A2(n4531), .ZN(n7172) );
  AND2_X1 U5597 ( .A1(n6048), .A2(n6139), .ZN(n9304) );
  INV_X1 U5598 ( .A(n5793), .ZN(n7152) );
  INV_X1 U5599 ( .A(n6654), .ZN(n6650) );
  NAND2_X1 U5600 ( .A1(n5083), .A2(n5082), .ZN(n9412) );
  NAND2_X1 U5601 ( .A1(n5131), .A2(n5130), .ZN(n9424) );
  INV_X1 U5602 ( .A(n4443), .ZN(n9398) );
  AOI21_X1 U5603 ( .B1(n4447), .B2(n4326), .A(n4387), .ZN(n4443) );
  NAND2_X1 U5604 ( .A1(n9076), .A2(n4448), .ZN(n4447) );
  OR2_X1 U5605 ( .A1(n9076), .A2(n9075), .ZN(n4445) );
  NAND2_X1 U5606 ( .A1(n4574), .A2(n4346), .ZN(n9711) );
  NAND2_X1 U5607 ( .A1(n7521), .A2(n7266), .ZN(n7269) );
  INV_X1 U5608 ( .A(n9712), .ZN(n9702) );
  XNOR2_X1 U5609 ( .A(n5091), .B(n5090), .ZN(n8241) );
  XNOR2_X1 U5610 ( .A(n5129), .B(n5128), .ZN(n7916) );
  NAND2_X1 U5611 ( .A1(n4786), .A2(n4790), .ZN(n5136) );
  OR2_X1 U5612 ( .A1(n5021), .A2(n4383), .ZN(n4786) );
  XNOR2_X1 U5613 ( .A(n5538), .B(n5537), .ZN(n7892) );
  NAND2_X1 U5614 ( .A1(n4793), .A2(n5024), .ZN(n5538) );
  NAND2_X1 U5615 ( .A1(n4951), .A2(n4949), .ZN(n5292) );
  NAND2_X1 U5616 ( .A1(n4556), .A2(n4347), .ZN(n4555) );
  INV_X1 U5617 ( .A(n4552), .ZN(n4551) );
  AND2_X1 U5618 ( .A1(n5300), .A2(n5238), .ZN(n5290) );
  NAND2_X1 U5619 ( .A1(n6905), .A2(n6904), .ZN(n7001) );
  NAND2_X1 U5620 ( .A1(n7503), .A2(n4898), .ZN(n7693) );
  NAND2_X1 U5621 ( .A1(n7869), .A2(n7868), .ZN(n8752) );
  AOI21_X1 U5622 ( .B1(n4883), .B2(n4885), .A(n4354), .ZN(n4881) );
  AND2_X1 U5623 ( .A1(n6186), .A2(n6185), .ZN(n6189) );
  NAND2_X1 U5624 ( .A1(n4890), .A2(n8274), .ZN(n8345) );
  NAND2_X1 U5625 ( .A1(n8336), .A2(n4894), .ZN(n4890) );
  OAI211_X1 U5626 ( .C1(n4879), .C2(n4343), .A(n7464), .B(n4873), .ZN(n7470)
         );
  INV_X1 U5627 ( .A(n8247), .ZN(n4845) );
  NOR2_X1 U5628 ( .A1(n8249), .A2(n8247), .ZN(n4846) );
  NAND2_X1 U5629 ( .A1(n7806), .A2(n7805), .ZN(n8788) );
  NAND2_X1 U5630 ( .A1(n6849), .A2(n6848), .ZN(n6885) );
  NAND2_X1 U5631 ( .A1(n6885), .A2(n6886), .ZN(n6884) );
  NAND2_X1 U5632 ( .A1(n4405), .A2(n8257), .ZN(n8375) );
  NAND2_X1 U5633 ( .A1(n7881), .A2(n7880), .ZN(n8745) );
  NAND2_X1 U5634 ( .A1(n8336), .A2(n8271), .ZN(n8398) );
  INV_X1 U5635 ( .A(n8692), .ZN(n7800) );
  INV_X1 U5636 ( .A(n4879), .ZN(n4876) );
  AOI21_X1 U5637 ( .B1(n4879), .B2(n4878), .A(n4343), .ZN(n4875) );
  NAND2_X1 U5638 ( .A1(n4882), .A2(n8260), .ZN(n8413) );
  NAND2_X1 U5639 ( .A1(n4405), .A2(n4886), .ZN(n4882) );
  OAI21_X1 U5640 ( .B1(n6849), .B2(n4853), .A(n4850), .ZN(n6860) );
  INV_X1 U5641 ( .A(n8423), .ZN(n8425) );
  NAND2_X1 U5642 ( .A1(n7694), .A2(n7639), .ZN(n8248) );
  OAI21_X1 U5643 ( .B1(n8429), .B2(n4666), .A(n7914), .ZN(n8502) );
  AND2_X1 U5644 ( .A1(n6322), .A2(n6321), .ZN(n6471) );
  AND2_X1 U5645 ( .A1(n6618), .A2(n6436), .ZN(n7626) );
  INV_X1 U5646 ( .A(n9736), .ZN(n9797) );
  AND2_X1 U5647 ( .A1(n7972), .A2(n7971), .ZN(n9584) );
  AND2_X1 U5648 ( .A1(n4473), .A2(n4470), .ZN(n7940) );
  INV_X1 U5649 ( .A(n4471), .ZN(n4470) );
  OR2_X1 U5650 ( .A1(n8521), .A2(n4474), .ZN(n4473) );
  INV_X1 U5651 ( .A(n7962), .ZN(n7963) );
  NAND2_X1 U5652 ( .A1(n4479), .A2(n4480), .ZN(n8495) );
  NAND2_X1 U5653 ( .A1(n8521), .A2(n4481), .ZN(n4479) );
  NAND2_X1 U5654 ( .A1(n4482), .A2(n4485), .ZN(n8508) );
  OR2_X1 U5655 ( .A1(n8521), .A2(n8530), .ZN(n4482) );
  AND2_X1 U5656 ( .A1(n8750), .A2(n4753), .ZN(n8538) );
  NAND2_X1 U5657 ( .A1(n8565), .A2(n8564), .ZN(n8750) );
  AND2_X1 U5658 ( .A1(n4651), .A2(n8080), .ZN(n8577) );
  NAND2_X1 U5659 ( .A1(n7950), .A2(n8079), .ZN(n8595) );
  NAND2_X1 U5660 ( .A1(n4732), .A2(n4736), .ZN(n8588) );
  NAND2_X1 U5661 ( .A1(n7846), .A2(n4738), .ZN(n4732) );
  NAND2_X1 U5662 ( .A1(n7846), .A2(n4903), .ZN(n8601) );
  NAND2_X1 U5663 ( .A1(n8646), .A2(n4661), .ZN(n8636) );
  NAND2_X1 U5664 ( .A1(n4749), .A2(n4747), .ZN(n8643) );
  NAND2_X1 U5665 ( .A1(n8685), .A2(n8684), .ZN(n8683) );
  NAND2_X1 U5666 ( .A1(n4464), .A2(n4463), .ZN(n8685) );
  NAND2_X1 U5667 ( .A1(n4743), .A2(n4742), .ZN(n8699) );
  NAND2_X1 U5668 ( .A1(n4744), .A2(n4324), .ZN(n7799) );
  NAND2_X1 U5669 ( .A1(n4744), .A2(n7668), .ZN(n7670) );
  AND2_X1 U5670 ( .A1(n4642), .A2(n8025), .ZN(n7715) );
  NAND2_X1 U5671 ( .A1(n7556), .A2(n8032), .ZN(n7672) );
  NAND2_X1 U5672 ( .A1(n7352), .A2(n4755), .ZN(n7554) );
  NAND2_X1 U5673 ( .A1(n7352), .A2(n7351), .ZN(n7354) );
  NAND2_X1 U5674 ( .A1(n7216), .A2(n7185), .ZN(n7188) );
  NAND2_X1 U5675 ( .A1(n7190), .A2(n8014), .ZN(n7208) );
  NAND2_X1 U5676 ( .A1(n9838), .A2(n9824), .ZN(n8718) );
  INV_X1 U5677 ( .A(n4671), .ZN(n8727) );
  INV_X1 U5678 ( .A(n4667), .ZN(n8239) );
  NAND3_X1 U5679 ( .A1(n4580), .A2(n6168), .A3(n4579), .ZN(n7955) );
  NAND2_X1 U5680 ( .A1(n6157), .A2(n8826), .ZN(n4579) );
  NAND2_X1 U5681 ( .A1(n6167), .A2(n4360), .ZN(n4580) );
  OR2_X1 U5682 ( .A1(n6085), .A2(n8826), .ZN(n4506) );
  NAND2_X1 U5683 ( .A1(n4665), .A2(n4342), .ZN(n6095) );
  INV_X1 U5684 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6437) );
  INV_X1 U5685 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9967) );
  INV_X1 U5686 ( .A(n6663), .ZN(n7505) );
  INV_X1 U5687 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10117) );
  INV_X1 U5688 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7078) );
  INV_X1 U5689 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7057) );
  INV_X1 U5690 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7011) );
  INV_X1 U5691 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6909) );
  INV_X1 U5692 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10140) );
  NAND2_X1 U5693 ( .A1(n5515), .A2(n5514), .ZN(n9446) );
  INV_X1 U5694 ( .A(n9073), .ZN(n9555) );
  NAND2_X1 U5695 ( .A1(n6069), .A2(n5913), .ZN(n6108) );
  NAND2_X1 U5696 ( .A1(n4705), .A2(n4710), .ZN(n8859) );
  NAND2_X1 U5697 ( .A1(n8940), .A2(n4712), .ZN(n4705) );
  NAND2_X1 U5698 ( .A1(n5118), .A2(n5117), .ZN(n9420) );
  AOI21_X1 U5699 ( .B1(n4696), .B2(n4910), .A(n4695), .ZN(n8867) );
  INV_X1 U5700 ( .A(n8916), .ZN(n4696) );
  NAND2_X1 U5701 ( .A1(n4702), .A2(n4703), .ZN(n8891) );
  NAND2_X1 U5702 ( .A1(n8963), .A2(n4704), .ZN(n4702) );
  AOI21_X1 U5703 ( .B1(n4699), .B2(n4698), .A(n4398), .ZN(n4697) );
  INV_X1 U5704 ( .A(n4704), .ZN(n4698) );
  NAND2_X1 U5705 ( .A1(n4726), .A2(n4728), .ZN(n8907) );
  AND4_X1 U5706 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n7746)
         );
  NAND2_X1 U5707 ( .A1(n5478), .A2(n5477), .ZN(n9461) );
  AOI21_X1 U5708 ( .B1(n4687), .B2(n4689), .A(n4367), .ZN(n4685) );
  NAND2_X1 U5709 ( .A1(n5225), .A2(n5224), .ZN(n9612) );
  AND4_X1 U5710 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n8977)
         );
  NAND2_X1 U5711 ( .A1(n5152), .A2(n5151), .ZN(n9472) );
  NAND2_X1 U5712 ( .A1(n9642), .A2(n9712), .ZN(n8959) );
  AND2_X1 U5713 ( .A1(n6059), .A2(n6651), .ZN(n9633) );
  NAND2_X1 U5714 ( .A1(n6056), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9648) );
  OR3_X1 U5715 ( .A1(n6057), .A2(n6048), .A3(n9712), .ZN(n8972) );
  INV_X1 U5716 ( .A(n4758), .ZN(n4547) );
  AOI21_X1 U5717 ( .B1(n5697), .B2(n9274), .A(n7164), .ZN(n4758) );
  INV_X1 U5718 ( .A(n9100), .ZN(n8975) );
  INV_X1 U5719 ( .A(n8920), .ZN(n9255) );
  NAND4_X1 U5720 ( .A1(n5399), .A2(n5398), .A3(n5397), .A4(n5396), .ZN(n8982)
         );
  OR2_X1 U5721 ( .A1(n5548), .A2(n5391), .ZN(n5398) );
  NAND4_X1 U5722 ( .A1(n5390), .A2(n5389), .A3(n5388), .A4(n5387), .ZN(n8983)
         );
  OR2_X1 U5723 ( .A1(n5548), .A2(n6589), .ZN(n5389) );
  NAND4_X1 U5724 ( .A1(n5425), .A2(n5424), .A3(n5423), .A4(n5422), .ZN(n8984)
         );
  OR2_X1 U5725 ( .A1(n5366), .A2(n5436), .ZN(n5439) );
  AND3_X1 U5726 ( .A1(n5369), .A2(n4905), .A3(n5368), .ZN(n5370) );
  NAND2_X1 U5727 ( .A1(n5335), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5336) );
  OR2_X1 U5728 ( .A1(n5365), .A2(n5349), .ZN(n5352) );
  NAND2_X1 U5729 ( .A1(n6592), .A2(n4407), .ZN(n6590) );
  INV_X1 U5730 ( .A(n6514), .ZN(n4407) );
  NOR2_X1 U5731 ( .A1(n6564), .A2(n6563), .ZN(n6636) );
  AOI21_X1 U5732 ( .B1(n6568), .B2(n10164), .A(n10158), .ZN(n6570) );
  NOR2_X1 U5733 ( .A1(n6703), .A2(n6702), .ZN(n6706) );
  AND2_X1 U5734 ( .A1(n7581), .A2(n7580), .ZN(n9018) );
  OAI22_X1 U5735 ( .A1(n9018), .A2(n9017), .B1(n7582), .B2(n9023), .ZN(n9033)
         );
  OAI211_X1 U5736 ( .C1(n5081), .C2(n4778), .A(n5069), .B(n4776), .ZN(n8186)
         );
  NAND2_X1 U5737 ( .A1(n4396), .A2(n4784), .ZN(n4778) );
  XOR2_X1 U5738 ( .A(n8186), .B(n9409), .Z(n8188) );
  INV_X1 U5739 ( .A(n4526), .ZN(n9409) );
  NAND2_X1 U5740 ( .A1(n9143), .A2(n4622), .ZN(n9415) );
  OR2_X1 U5741 ( .A1(n9154), .A2(n9144), .ZN(n4622) );
  NAND2_X1 U5742 ( .A1(n9151), .A2(n9153), .ZN(n9423) );
  NAND2_X1 U5743 ( .A1(n4823), .A2(n4820), .ZN(n9152) );
  AOI21_X1 U5744 ( .B1(n9193), .B2(n9501), .A(n9192), .ZN(n9432) );
  NAND2_X1 U5745 ( .A1(n4609), .A2(n4610), .ZN(n9191) );
  INV_X1 U5746 ( .A(n9430), .ZN(n9189) );
  NOR2_X1 U5747 ( .A1(n9219), .A2(n9129), .ZN(n9204) );
  NAND2_X1 U5748 ( .A1(n4414), .A2(n4419), .ZN(n9098) );
  NAND2_X1 U5749 ( .A1(n4418), .A2(n4423), .ZN(n9223) );
  NAND2_X1 U5750 ( .A1(n9243), .A2(n4424), .ZN(n4418) );
  OR2_X1 U5751 ( .A1(n4320), .A2(n7619), .ZN(n5526) );
  NAND2_X1 U5752 ( .A1(n9253), .A2(n9127), .ZN(n9235) );
  AND2_X1 U5753 ( .A1(n4425), .A2(n4426), .ZN(n9229) );
  NAND2_X1 U5754 ( .A1(n9243), .A2(n9095), .ZN(n4425) );
  INV_X1 U5755 ( .A(n9452), .ZN(n9249) );
  AND2_X1 U5756 ( .A1(n4428), .A2(n4429), .ZN(n9263) );
  NAND2_X1 U5757 ( .A1(n9302), .A2(n9124), .ZN(n9286) );
  NAND2_X1 U5758 ( .A1(n4433), .A2(n4435), .ZN(n9279) );
  NAND2_X1 U5759 ( .A1(n4434), .A2(n4437), .ZN(n4433) );
  NAND2_X1 U5760 ( .A1(n4828), .A2(n4829), .ZN(n9312) );
  AND2_X1 U5761 ( .A1(n5167), .A2(n5166), .ZN(n9338) );
  OAI21_X1 U5762 ( .B1(n9087), .B2(n4833), .A(n9086), .ZN(n9331) );
  NAND2_X1 U5763 ( .A1(n4618), .A2(n9118), .ZN(n9356) );
  NAND2_X1 U5764 ( .A1(n9362), .A2(n9117), .ZN(n4618) );
  INV_X1 U5765 ( .A(n9087), .ZN(n9346) );
  INV_X1 U5766 ( .A(n9488), .ZN(n9372) );
  NAND2_X1 U5767 ( .A1(n5242), .A2(n5241), .ZN(n9596) );
  NAND2_X1 U5768 ( .A1(n5256), .A2(n5255), .ZN(n9074) );
  NAND2_X1 U5769 ( .A1(n7076), .A2(n5539), .ZN(n4409) );
  INV_X1 U5770 ( .A(n9711), .ZN(n7730) );
  AND2_X1 U5771 ( .A1(n7391), .A2(n7390), .ZN(n7392) );
  INV_X1 U5772 ( .A(n9697), .ZN(n7389) );
  AND3_X1 U5773 ( .A1(n5383), .A2(n5382), .A3(n5381), .ZN(n7494) );
  AND3_X1 U5774 ( .A1(n5416), .A2(n5415), .A3(n5414), .ZN(n7535) );
  INV_X1 U5775 ( .A(n9594), .ZN(n9559) );
  AND2_X1 U5776 ( .A1(n6050), .A2(n6650), .ZN(n9594) );
  AND2_X1 U5777 ( .A1(n7140), .A2(n7152), .ZN(n6050) );
  NOR2_X1 U5778 ( .A1(n5775), .A2(n5774), .ZN(n9578) );
  NAND2_X1 U5779 ( .A1(n5773), .A2(n5772), .ZN(n5774) );
  NOR2_X1 U5780 ( .A1(n8188), .A2(n9704), .ZN(n5775) );
  NAND2_X1 U5781 ( .A1(n8186), .A2(n9712), .ZN(n5773) );
  INV_X1 U5782 ( .A(n4523), .ZN(n9514) );
  OAI21_X1 U5783 ( .B1(n9410), .B2(n4525), .A(n4524), .ZN(n4523) );
  AOI21_X1 U5784 ( .B1(n9412), .B2(n9712), .A(n9411), .ZN(n4524) );
  NAND2_X1 U5785 ( .A1(n4526), .A2(n9713), .ZN(n4525) );
  NAND2_X1 U5786 ( .A1(n4623), .A2(n4357), .ZN(n9517) );
  INV_X1 U5787 ( .A(n9416), .ZN(n4623) );
  INV_X2 U5788 ( .A(n9722), .ZN(n9724) );
  NAND2_X1 U5789 ( .A1(n7140), .A2(n6329), .ZN(n9666) );
  OR2_X1 U5790 ( .A1(n5081), .A2(n4784), .ZN(n4780) );
  CLKBUF_X1 U5791 ( .A(n5753), .Z(n5754) );
  INV_X1 U5792 ( .A(n5786), .ZN(n7725) );
  INV_X1 U5793 ( .A(n5756), .ZN(n5760) );
  XNOR2_X1 U5794 ( .A(n5513), .B(n5512), .ZN(n7867) );
  INV_X1 U5795 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6381) );
  INV_X1 U5796 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10104) );
  INV_X1 U5797 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6342) );
  INV_X1 U5798 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6325) );
  INV_X1 U5799 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6323) );
  OAI21_X1 U5800 ( .B1(n4937), .B2(n4558), .A(n4556), .ZN(n5299) );
  INV_X1 U5801 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U5802 ( .A1(n4937), .A2(n4936), .ZN(n5319) );
  INV_X1 U5803 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6309) );
  INV_X1 U5804 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6317) );
  INV_X1 U5805 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6308) );
  XNOR2_X1 U5806 ( .A(n5432), .B(n5431), .ZN(n6529) );
  NOR2_X1 U5807 ( .A1(n7445), .A2(n10182), .ZN(n9962) );
  NAND2_X1 U5808 ( .A1(n7106), .A2(n7075), .ZN(n7240) );
  NAND2_X1 U5809 ( .A1(n6877), .A2(n6733), .ZN(n6926) );
  INV_X1 U5810 ( .A(n4634), .ZN(n4633) );
  NAND2_X1 U5811 ( .A1(n4670), .A2(n4668), .ZN(P2_U3268) );
  AOI211_X1 U5812 ( .C1(n8725), .C2(n8716), .A(n4669), .B(n8228), .ZN(n4668)
         );
  NAND2_X1 U5813 ( .A1(n4671), .A2(n9838), .ZN(n4670) );
  NAND2_X1 U5814 ( .A1(n4584), .A2(n4583), .ZN(P2_U3549) );
  NAND2_X1 U5815 ( .A1(n9931), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4583) );
  NAND2_X1 U5816 ( .A1(n8809), .A2(n9934), .ZN(n4584) );
  NAND2_X1 U5817 ( .A1(n4457), .A2(n4397), .ZN(P2_U3517) );
  NAND2_X1 U5818 ( .A1(n8809), .A2(n9923), .ZN(n4457) );
  OR2_X1 U5819 ( .A1(n6171), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4323) );
  NAND4_X1 U5820 ( .A1(n6210), .A2(n6209), .A3(n6208), .A4(n6207), .ZN(n6771)
         );
  AND2_X1 U5821 ( .A1(n7669), .A2(n7668), .ZN(n4324) );
  OR2_X1 U5822 ( .A1(n5377), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5379) );
  OR2_X1 U5823 ( .A1(n9446), .A2(n9256), .ZN(n4325) );
  AND2_X1 U5824 ( .A1(n4446), .A2(n9495), .ZN(n4326) );
  NAND2_X1 U5825 ( .A1(n4331), .A2(n4431), .ZN(n4430) );
  NAND2_X1 U5826 ( .A1(n8517), .A2(n8109), .ZN(n4328) );
  AND2_X1 U5827 ( .A1(n4742), .A2(n8698), .ZN(n4329) );
  INV_X1 U5828 ( .A(n4756), .ZN(n4755) );
  NAND2_X1 U5829 ( .A1(n7353), .A2(n7351), .ZN(n4756) );
  AND3_X1 U5830 ( .A1(n8168), .A2(n7985), .A3(n4634), .ZN(n4330) );
  INV_X1 U5831 ( .A(n8917), .ZN(n4695) );
  INV_X1 U5832 ( .A(n8070), .ZN(n4659) );
  INV_X1 U5833 ( .A(n8120), .ZN(n4649) );
  NAND2_X1 U5834 ( .A1(n8121), .A2(n8122), .ZN(n8225) );
  INV_X1 U5835 ( .A(n8225), .ZN(n4472) );
  NAND2_X1 U5836 ( .A1(n7894), .A2(n7893), .ZN(n8741) );
  INV_X1 U5837 ( .A(n8741), .ZN(n4486) );
  OR2_X1 U5838 ( .A1(n9461), .A2(n9307), .ZN(n4331) );
  NAND2_X1 U5839 ( .A1(n7798), .A2(n7797), .ZN(n8762) );
  AND2_X1 U5840 ( .A1(n9118), .A2(n5628), .ZN(n9117) );
  INV_X1 U5841 ( .A(n9117), .ZN(n4616) );
  NAND2_X1 U5842 ( .A1(n8007), .A2(n6940), .ZN(n9813) );
  INV_X1 U5843 ( .A(n9813), .ZN(n4741) );
  AND2_X1 U5844 ( .A1(n9420), .A2(n9108), .ZN(n4332) );
  AND2_X1 U5845 ( .A1(n4829), .A2(n9321), .ZN(n4333) );
  OR2_X1 U5846 ( .A1(n8015), .A2(n8150), .ZN(n4334) );
  AND2_X1 U5847 ( .A1(n9125), .A2(n5562), .ZN(n4335) );
  INV_X1 U5848 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4717) );
  XNOR2_X1 U5849 ( .A(n5598), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5769) );
  AND2_X1 U5850 ( .A1(n8593), .A2(n8608), .ZN(n4336) );
  OR2_X1 U5851 ( .A1(n9458), .A2(n8920), .ZN(n5641) );
  INV_X1 U5852 ( .A(n8041), .ZN(n4590) );
  AND2_X1 U5853 ( .A1(n9461), .A2(n9307), .ZN(n4337) );
  AND2_X1 U5854 ( .A1(n8076), .A2(n8070), .ZN(n4338) );
  AND2_X1 U5855 ( .A1(n8027), .A2(n8023), .ZN(n8153) );
  INV_X1 U5856 ( .A(n9461), .ZN(n9284) );
  INV_X1 U5857 ( .A(n4700), .ZN(n4699) );
  OR2_X1 U5858 ( .A1(n8889), .A2(n4701), .ZN(n4700) );
  INV_X1 U5859 ( .A(n8324), .ZN(n4484) );
  OR2_X1 U5860 ( .A1(n9503), .A2(n4532), .ZN(n4339) );
  INV_X1 U5861 ( .A(n9091), .ZN(n4437) );
  NAND2_X1 U5862 ( .A1(n4681), .A2(n4680), .ZN(n6115) );
  OAI21_X1 U5863 ( .B1(n7072), .B2(n4876), .A(n4875), .ZN(n7465) );
  NAND2_X1 U5864 ( .A1(n4665), .A2(n4522), .ZN(n4521) );
  AND2_X1 U5865 ( .A1(n6014), .A2(n6013), .ZN(n4340) );
  AND2_X1 U5866 ( .A1(n8833), .A2(n4667), .ZN(n4341) );
  INV_X1 U5867 ( .A(n9109), .ZN(n4817) );
  AND2_X1 U5868 ( .A1(n4488), .A2(n4327), .ZN(n4342) );
  NOR2_X1 U5869 ( .A1(n7238), .A2(n7237), .ZN(n4343) );
  NAND2_X1 U5870 ( .A1(n5371), .A2(n5370), .ZN(n5838) );
  NOR2_X1 U5871 ( .A1(n4715), .A2(n4714), .ZN(n5150) );
  NAND2_X1 U5872 ( .A1(n4417), .A2(n4415), .ZN(n9182) );
  XNOR2_X1 U5873 ( .A(n8730), .B(n8438), .ZN(n8501) );
  INV_X1 U5874 ( .A(n8938), .ZN(n4713) );
  INV_X1 U5875 ( .A(n4341), .ZN(n7912) );
  NAND4_X1 U5876 ( .A1(n5744), .A2(n5063), .A3(n5062), .A4(n5061), .ZN(n4344)
         );
  NAND2_X1 U5877 ( .A1(n7927), .A2(n7926), .ZN(n8724) );
  OR2_X1 U5878 ( .A1(n9561), .A2(n7746), .ZN(n7741) );
  AND2_X1 U5879 ( .A1(n9906), .A2(n4591), .ZN(n4345) );
  AND2_X1 U5880 ( .A1(n5294), .A2(n4575), .ZN(n4346) );
  NAND2_X1 U5881 ( .A1(n4480), .A2(n8166), .ZN(n4478) );
  AND2_X1 U5882 ( .A1(n4945), .A2(n4944), .ZN(n4347) );
  AND2_X1 U5883 ( .A1(n9446), .A2(n9256), .ZN(n4348) );
  NOR2_X1 U5884 ( .A1(n9507), .A2(n9555), .ZN(n4441) );
  NAND2_X1 U5885 ( .A1(n7836), .A2(n7835), .ZN(n8773) );
  INV_X1 U5886 ( .A(n8773), .ZN(n4597) );
  AND2_X1 U5887 ( .A1(n8980), .A2(n7600), .ZN(n4349) );
  AND4_X1 U5888 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n4350)
         );
  INV_X1 U5889 ( .A(n5585), .ZN(n4403) );
  INV_X1 U5890 ( .A(n7987), .ZN(n4641) );
  NAND2_X1 U5891 ( .A1(n9098), .A2(n9097), .ZN(n9197) );
  AND2_X1 U5892 ( .A1(n4726), .A2(n4724), .ZN(n4351) );
  AND2_X1 U5893 ( .A1(n4770), .A2(n4768), .ZN(n4352) );
  OR2_X1 U5894 ( .A1(n9387), .A2(n9364), .ZN(n9115) );
  INV_X1 U5895 ( .A(n5913), .ZN(n4684) );
  AND2_X1 U5896 ( .A1(n4548), .A2(n4546), .ZN(n4353) );
  NAND2_X1 U5897 ( .A1(n4578), .A2(n6174), .ZN(n6295) );
  AND2_X1 U5898 ( .A1(n8263), .A2(n8262), .ZN(n4354) );
  AND2_X1 U5899 ( .A1(n8277), .A2(n8276), .ZN(n4355) );
  INV_X1 U5900 ( .A(n4907), .ZN(n4774) );
  AND2_X1 U5901 ( .A1(n8021), .A2(n8022), .ZN(n8152) );
  NAND3_X1 U5902 ( .A1(n5338), .A2(n5337), .A3(n5336), .ZN(n5823) );
  INV_X1 U5903 ( .A(n4729), .ZN(n4727) );
  NOR2_X1 U5904 ( .A1(n8848), .A2(n4730), .ZN(n4729) );
  AND2_X1 U5905 ( .A1(n8051), .A2(n8052), .ZN(n8708) );
  INV_X1 U5906 ( .A(n4577), .ZN(n8513) );
  NOR2_X1 U5907 ( .A1(n8522), .A2(n8737), .ZN(n4577) );
  NOR2_X1 U5908 ( .A1(n9244), .A2(n4540), .ZN(n4538) );
  AND2_X1 U5909 ( .A1(n5639), .A2(n5643), .ZN(n9313) );
  INV_X1 U5910 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9535) );
  AND2_X1 U5911 ( .A1(n5673), .A2(n5672), .ZN(n9107) );
  AND2_X1 U5912 ( .A1(n7569), .A2(n8442), .ZN(n4356) );
  INV_X1 U5913 ( .A(n4611), .ZN(n4610) );
  OAI21_X1 U5914 ( .B1(n9132), .B2(n5658), .A(n9131), .ZN(n4611) );
  AND2_X1 U5915 ( .A1(n9418), .A2(n4450), .ZN(n4357) );
  AND2_X1 U5916 ( .A1(n8803), .A2(n8711), .ZN(n4358) );
  INV_X1 U5917 ( .A(n5356), .ZN(n6140) );
  INV_X1 U5918 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4863) );
  NOR2_X1 U5919 ( .A1(n8792), .A2(n8710), .ZN(n4359) );
  AND2_X1 U5920 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4360) );
  INV_X1 U5921 ( .A(n4543), .ZN(n9230) );
  NOR2_X1 U5922 ( .A1(n9244), .A2(n9446), .ZN(n4543) );
  OR2_X1 U5923 ( .A1(n9472), .A2(n8902), .ZN(n5639) );
  INV_X1 U5924 ( .A(n7855), .ZN(n4740) );
  NOR2_X1 U5925 ( .A1(n5900), .A2(n5899), .ZN(n4361) );
  INV_X1 U5926 ( .A(n4589), .ZN(n4588) );
  NAND2_X1 U5927 ( .A1(n4345), .A2(n4590), .ZN(n4589) );
  INV_X1 U5928 ( .A(n4436), .ZN(n4435) );
  NOR2_X1 U5929 ( .A1(n9298), .A2(n9322), .ZN(n4436) );
  AND2_X1 U5930 ( .A1(n8788), .A2(n8059), .ZN(n4362) );
  INV_X1 U5931 ( .A(n7807), .ZN(n4748) );
  AND2_X1 U5932 ( .A1(n8788), .A2(n8693), .ZN(n7807) );
  NOR2_X1 U5933 ( .A1(n8593), .A2(n8608), .ZN(n4364) );
  NAND2_X1 U5934 ( .A1(n4519), .A2(n4342), .ZN(n4365) );
  NOR2_X1 U5935 ( .A1(n8730), .A2(n8438), .ZN(n4366) );
  INV_X1 U5936 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5761) );
  AND2_X1 U5937 ( .A1(n5941), .A2(n7777), .ZN(n4367) );
  INV_X1 U5938 ( .A(n4899), .ZN(n4898) );
  OR2_X1 U5939 ( .A1(n7623), .A2(n4900), .ZN(n4899) );
  AND2_X1 U5940 ( .A1(n4959), .A2(SI_11_), .ZN(n4368) );
  NAND2_X1 U5941 ( .A1(n8024), .A2(n8023), .ZN(n4369) );
  OR2_X1 U5942 ( .A1(n8724), .A2(n4484), .ZN(n4370) );
  NAND2_X1 U5943 ( .A1(n4942), .A2(n4941), .ZN(n4945) );
  OR2_X1 U5944 ( .A1(n8724), .A2(n8324), .ZN(n8121) );
  INV_X1 U5945 ( .A(n4478), .ZN(n4477) );
  OR2_X1 U5946 ( .A1(n9094), .A2(n4348), .ZN(n4371) );
  NAND2_X1 U5947 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n4372) );
  NAND2_X1 U5948 ( .A1(n8509), .A2(n4483), .ZN(n4373) );
  NAND2_X1 U5949 ( .A1(n4823), .A2(n4821), .ZN(n9151) );
  INV_X1 U5950 ( .A(n8684), .ZN(n4462) );
  INV_X1 U5951 ( .A(n4980), .ZN(n4802) );
  AND2_X1 U5952 ( .A1(n4617), .A2(n9115), .ZN(n4374) );
  AND2_X1 U5953 ( .A1(n8721), .A2(n4585), .ZN(n4375) );
  AND2_X1 U5954 ( .A1(n4462), .A2(n8053), .ZN(n4376) );
  AND2_X1 U5955 ( .A1(n9099), .A2(n9097), .ZN(n4377) );
  AND2_X1 U5956 ( .A1(n5362), .A2(n5364), .ZN(n4378) );
  AND2_X1 U5957 ( .A1(n8917), .A2(n8868), .ZN(n4379) );
  AND2_X1 U5958 ( .A1(n7187), .A2(n7185), .ZN(n4380) );
  AND2_X1 U5959 ( .A1(n4372), .A2(n5065), .ZN(n4381) );
  OR2_X1 U5960 ( .A1(n8041), .A2(n7555), .ZN(n8033) );
  NAND2_X1 U5961 ( .A1(n4329), .A2(n8684), .ZN(n4382) );
  INV_X1 U5962 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4809) );
  OR2_X2 U5963 ( .A1(n7986), .A2(n6234), .ZN(n8137) );
  NAND2_X1 U5964 ( .A1(n8189), .A2(n7260), .ZN(n6722) );
  OR2_X1 U5965 ( .A1(n5537), .A2(n4792), .ZN(n4383) );
  NAND2_X1 U5966 ( .A1(n8270), .A2(n8269), .ZN(n8336) );
  NOR2_X1 U5967 ( .A1(n9503), .A2(n4533), .ZN(n9347) );
  NAND2_X1 U5968 ( .A1(n5179), .A2(n5060), .ZN(n5162) );
  NOR2_X1 U5969 ( .A1(n9503), .A2(n9612), .ZN(n4384) );
  NAND3_X1 U5970 ( .A1(n5236), .A2(n5058), .A3(n4717), .ZN(n4385) );
  AND2_X1 U5971 ( .A1(n9472), .A2(n9305), .ZN(n4386) );
  NAND2_X1 U5972 ( .A1(n7503), .A2(n7502), .ZN(n7624) );
  NAND2_X1 U5973 ( .A1(n6116), .A2(n5934), .ZN(n7776) );
  AND2_X1 U5974 ( .A1(n9596), .A2(n9077), .ZN(n4387) );
  NAND2_X1 U5975 ( .A1(n5164), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U5976 ( .A1(n4647), .A2(n8054), .ZN(n8661) );
  NAND2_X1 U5977 ( .A1(n4445), .A2(n4448), .ZN(n9492) );
  OR2_X1 U5978 ( .A1(n8313), .A2(n8662), .ZN(n4388) );
  INV_X1 U5979 ( .A(n9119), .ZN(n4615) );
  NAND2_X1 U5980 ( .A1(n5929), .A2(n5928), .ZN(n6116) );
  OR2_X1 U5981 ( .A1(n9488), .A2(n9083), .ZN(n4389) );
  NAND2_X1 U5982 ( .A1(n5236), .A2(n5058), .ZN(n5221) );
  INV_X1 U5983 ( .A(n8596), .ZN(n8347) );
  AND2_X1 U5984 ( .A1(n8646), .A2(n8063), .ZN(n4390) );
  NOR2_X1 U5985 ( .A1(n4337), .A2(n4436), .ZN(n4432) );
  INV_X1 U5986 ( .A(n4537), .ZN(n9315) );
  NOR2_X1 U5987 ( .A1(n9333), .A2(n9472), .ZN(n4537) );
  AND2_X1 U5988 ( .A1(n4828), .A2(n4333), .ZN(n4391) );
  NOR2_X1 U5989 ( .A1(n8784), .A2(n8637), .ZN(n4392) );
  INV_X1 U5990 ( .A(n4593), .ZN(n8589) );
  NOR2_X1 U5991 ( .A1(n8631), .A2(n4594), .ZN(n4593) );
  AND2_X1 U5992 ( .A1(n5150), .A2(n4904), .ZN(n5748) );
  AND2_X1 U5993 ( .A1(n5462), .A2(n5005), .ZN(n4393) );
  AND2_X1 U5994 ( .A1(n4749), .A2(n4748), .ZN(n4394) );
  INV_X1 U5995 ( .A(n9094), .ZN(n4426) );
  INV_X1 U5996 ( .A(n4430), .ZN(n4429) );
  INV_X2 U5997 ( .A(n5341), .ZN(n5539) );
  OAI21_X1 U5998 ( .B1(n7345), .B2(n4835), .A(n4834), .ZN(n7736) );
  NAND2_X1 U5999 ( .A1(n6099), .A2(n6100), .ZN(n6097) );
  NAND2_X1 U6000 ( .A1(n7230), .A2(n4588), .ZN(n4395) );
  AOI21_X1 U6001 ( .B1(n4755), .B2(n8153), .A(n4356), .ZN(n4468) );
  AND2_X1 U6002 ( .A1(n4781), .A2(n5539), .ZN(n4396) );
  OR2_X1 U6003 ( .A1(n9923), .A2(n6377), .ZN(n4397) );
  OAI21_X1 U6004 ( .B1(n7222), .B2(n4756), .A(n4468), .ZN(n7665) );
  NAND2_X1 U6005 ( .A1(n5374), .A2(n5373), .ZN(n5588) );
  NAND2_X1 U6006 ( .A1(n7644), .A2(n7643), .ZN(n8792) );
  INV_X1 U6007 ( .A(n8792), .ZN(n4581) );
  NAND2_X1 U6008 ( .A1(n7391), .A2(n4836), .ZN(n7601) );
  AND2_X1 U6009 ( .A1(n5977), .A2(n5976), .ZN(n4398) );
  AND2_X1 U6010 ( .A1(n4783), .A2(n5054), .ZN(n4399) );
  INV_X1 U6011 ( .A(n4582), .ZN(n8700) );
  NOR2_X1 U6012 ( .A1(n8701), .A2(n8797), .ZN(n4582) );
  AND2_X1 U6013 ( .A1(n7075), .A2(n4874), .ZN(n4879) );
  AND2_X1 U6014 ( .A1(n5043), .A2(n5042), .ZN(n4400) );
  INV_X1 U6015 ( .A(n8025), .ZN(n4643) );
  AND2_X1 U6016 ( .A1(n4396), .A2(n4777), .ZN(n4401) );
  OR2_X1 U6017 ( .A1(n6654), .A2(n6688), .ZN(n9704) );
  INV_X1 U6018 ( .A(n9704), .ZN(n9713) );
  AND2_X1 U6019 ( .A1(n6690), .A2(n6689), .ZN(n9553) );
  INV_X1 U6020 ( .A(n9553), .ZN(n9501) );
  NAND2_X1 U6021 ( .A1(n6878), .A2(n6879), .ZN(n6877) );
  OAI211_X1 U6022 ( .C1(n6878), .C2(n4869), .A(n4867), .B(n4864), .ZN(n6751)
         );
  AND2_X1 U6023 ( .A1(n6722), .A2(n8171), .ZN(n4402) );
  INV_X1 U6024 ( .A(n7985), .ZN(n7982) );
  MUX2_X1 U6025 ( .A(n5686), .B(n5685), .S(n5689), .Z(n5695) );
  NAND2_X1 U6026 ( .A1(n5718), .A2(n5689), .ZN(n4565) );
  OAI21_X1 U6027 ( .B1(n5627), .B2(n5626), .A(n5689), .ZN(n4562) );
  OAI21_X1 U6028 ( .B1(n8510), .B2(n8509), .A(n8108), .ZN(n8500) );
  AND2_X1 U6029 ( .A1(n8000), .A2(n7999), .ZN(n8144) );
  AND2_X1 U6030 ( .A1(n5648), .A2(n5511), .ZN(n5718) );
  NAND2_X1 U6031 ( .A1(n4986), .A2(n4985), .ZN(n5161) );
  OAI21_X1 U6032 ( .B1(n5493), .B2(n5492), .A(n5000), .ZN(n5476) );
  NOR2_X2 U6033 ( .A1(n5688), .A2(n5687), .ZN(n5684) );
  OR2_X2 U6034 ( .A1(n5671), .A2(n4404), .ZN(n5669) );
  INV_X2 U6035 ( .A(n5755), .ZN(n5064) );
  NOR4_X1 U6036 ( .A1(n5647), .A2(n5646), .A3(n5645), .A4(n5644), .ZN(n5649)
         );
  OAI21_X2 U6037 ( .B1(n5592), .B2(n5591), .A(n7262), .ZN(n5602) );
  NAND2_X1 U6038 ( .A1(n5695), .A2(n4757), .ZN(n4550) );
  NOR4_X2 U6039 ( .A1(n5617), .A2(n5616), .A3(n7742), .A4(n5615), .ZN(n5624)
         );
  OAI211_X1 U6040 ( .C1(n4564), .C2(n4563), .A(n4562), .B(n9117), .ZN(n4561)
         );
  OAI21_X1 U6041 ( .B1(n4549), .B2(n5582), .A(n9061), .ZN(n4548) );
  AND2_X1 U6042 ( .A1(n7069), .A2(n7103), .ZN(n7073) );
  NAND2_X1 U6043 ( .A1(n4498), .A2(n4501), .ZN(n8077) );
  NAND2_X1 U6044 ( .A1(n4412), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4411) );
  INV_X1 U6045 ( .A(n4496), .ZN(n4494) );
  NAND2_X1 U6046 ( .A1(n4495), .A2(n4493), .ZN(n8176) );
  NAND2_X1 U6047 ( .A1(n8141), .A2(n8140), .ZN(n4497) );
  AOI21_X1 U6048 ( .B1(n8030), .B2(n8029), .A(n8028), .ZN(n8035) );
  OAI211_X1 U6049 ( .C1(n4636), .C2(n4633), .A(n4632), .B(n4630), .ZN(P2_U3244) );
  NOR2_X1 U6050 ( .A1(n8948), .A2(n8947), .ZN(n8946) );
  NAND2_X1 U6051 ( .A1(n4995), .A2(n4994), .ZN(n5493) );
  NAND2_X1 U6052 ( .A1(n4545), .A2(n4920), .ZN(n5427) );
  NAND2_X1 U6053 ( .A1(n4544), .A2(n4924), .ZN(n5411) );
  NAND2_X1 U6054 ( .A1(n5476), .A2(n5475), .ZN(n4775) );
  NAND2_X1 U6055 ( .A1(n4796), .A2(n4800), .ZN(n4986) );
  NAND2_X1 U6056 ( .A1(n5293), .A2(n4950), .ZN(n4952) );
  NAND2_X1 U6057 ( .A1(n9243), .A2(n4419), .ZN(n4417) );
  NAND2_X1 U6058 ( .A1(n9076), .A2(n4442), .ZN(n4440) );
  NAND2_X1 U6059 ( .A1(n4440), .A2(n4438), .ZN(n9378) );
  INV_X1 U6060 ( .A(n4441), .ZN(n4448) );
  AND3_X2 U6061 ( .A1(n6174), .A2(n6078), .A3(n4578), .ZN(n4665) );
  NAND3_X1 U6062 ( .A1(n4458), .A2(n4375), .A3(n4586), .ZN(n8809) );
  INV_X1 U6063 ( .A(n4743), .ZN(n4459) );
  OAI21_X1 U6064 ( .B1(n4459), .B2(n4382), .A(n4460), .ZN(n8667) );
  NAND2_X1 U6065 ( .A1(n7222), .A2(n4468), .ZN(n4466) );
  NAND2_X1 U6066 ( .A1(n4466), .A2(n4465), .ZN(n7667) );
  NAND2_X1 U6067 ( .A1(n6300), .A2(n4488), .ZN(n6646) );
  AND2_X1 U6068 ( .A1(n4350), .A2(n4488), .ZN(n4487) );
  OAI21_X1 U6069 ( .B1(n8017), .B2(n4489), .A(n4490), .ZN(n8030) );
  OR2_X1 U6070 ( .A1(n8058), .A2(n4504), .ZN(n4498) );
  NAND2_X1 U6071 ( .A1(n8058), .A2(n4501), .ZN(n4500) );
  NAND2_X1 U6072 ( .A1(n4507), .A2(n4376), .ZN(n8057) );
  NAND2_X1 U6073 ( .A1(n4509), .A2(n4508), .ZN(n4507) );
  NAND3_X1 U6074 ( .A1(n4514), .A2(n4511), .A3(n4510), .ZN(n4509) );
  NAND2_X1 U6075 ( .A1(n4513), .A2(n4512), .ZN(n4511) );
  NOR2_X1 U6076 ( .A1(n4641), .A2(n8126), .ZN(n4512) );
  NAND2_X1 U6077 ( .A1(n8038), .A2(n8040), .ZN(n4513) );
  INV_X1 U6078 ( .A(n8050), .ZN(n4514) );
  NAND2_X1 U6079 ( .A1(n4342), .A2(n4515), .ZN(n6200) );
  NAND2_X1 U6080 ( .A1(n4839), .A2(n5193), .ZN(n5755) );
  AND2_X2 U6081 ( .A1(n4619), .A2(n5236), .ZN(n5193) );
  AND2_X1 U6082 ( .A1(n5193), .A2(n5059), .ZN(n5179) );
  NAND2_X1 U6083 ( .A1(n5356), .A2(n6304), .ZN(n5341) );
  NAND2_X2 U6084 ( .A1(n5753), .A2(n7789), .ZN(n5356) );
  NAND2_X1 U6085 ( .A1(n5356), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U6086 ( .A1(n5345), .A2(n4529), .ZN(n5357) );
  INV_X1 U6087 ( .A(n9670), .ZN(n7177) );
  NOR2_X2 U6088 ( .A1(n7173), .A2(n9626), .ZN(n7530) );
  AND2_X2 U6089 ( .A1(n5363), .A2(n4378), .ZN(n9670) );
  NOR3_X4 U6090 ( .A1(n9333), .A2(n9458), .A3(n4535), .ZN(n9266) );
  INV_X1 U6091 ( .A(n4538), .ZN(n9185) );
  NAND2_X1 U6092 ( .A1(n5427), .A2(n5426), .ZN(n4544) );
  NAND2_X1 U6093 ( .A1(n5360), .A2(n5359), .ZN(n4545) );
  AOI21_X1 U6094 ( .B1(n4550), .B2(n5701), .A(n4547), .ZN(n4546) );
  NOR2_X1 U6095 ( .A1(n6125), .A2(n4550), .ZN(n4549) );
  INV_X1 U6096 ( .A(n4937), .ZN(n4554) );
  OAI21_X1 U6097 ( .B1(n4555), .B2(n4554), .A(n4551), .ZN(n5293) );
  OR2_X1 U6098 ( .A1(n5633), .A2(n5634), .ZN(n4559) );
  NAND2_X1 U6099 ( .A1(n4569), .A2(n4567), .ZN(n4566) );
  INV_X1 U6100 ( .A(n7056), .ZN(n4576) );
  NOR2_X2 U6101 ( .A1(n8730), .A2(n8513), .ZN(n8496) );
  NOR2_X2 U6102 ( .A1(n8687), .A2(n8788), .ZN(n8674) );
  INV_X1 U6103 ( .A(n4592), .ZN(n8581) );
  NAND2_X1 U6104 ( .A1(n7738), .A2(n4601), .ZN(n4600) );
  OAI21_X1 U6105 ( .B1(n9219), .B2(n4607), .A(n4605), .ZN(n9173) );
  NAND2_X1 U6106 ( .A1(n9302), .A2(n4612), .ZN(n9288) );
  NAND2_X1 U6107 ( .A1(n9116), .A2(n4374), .ZN(n4613) );
  NAND2_X1 U6108 ( .A1(n4613), .A2(n4614), .ZN(n9340) );
  AND4_X2 U6109 ( .A1(n5361), .A2(n5055), .A3(n5428), .A4(n4838), .ZN(n5236)
         );
  AND3_X2 U6110 ( .A1(n4620), .A2(n5057), .A3(n5056), .ZN(n5058) );
  NAND2_X1 U6111 ( .A1(n5064), .A2(n5761), .ZN(n5072) );
  NAND2_X1 U6112 ( .A1(n5064), .A2(n4626), .ZN(n4628) );
  NOR2_X1 U6113 ( .A1(n4629), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U6114 ( .A1(n7981), .A2(n4330), .ZN(n4632) );
  NAND2_X1 U6115 ( .A1(n8691), .A2(n8055), .ZN(n4647) );
  NAND2_X1 U6116 ( .A1(n4647), .A2(n4645), .ZN(n7948) );
  NOR2_X2 U6117 ( .A1(n8226), .A2(n8225), .ZN(n8224) );
  NAND2_X1 U6118 ( .A1(n4363), .A2(n4858), .ZN(n4667) );
  NAND2_X2 U6119 ( .A1(n6236), .A2(n6982), .ZN(n8145) );
  NAND2_X1 U6120 ( .A1(n6068), .A2(n4683), .ZN(n4680) );
  NAND2_X1 U6121 ( .A1(n5929), .A2(n4687), .ZN(n4686) );
  NAND2_X2 U6122 ( .A1(n4686), .A2(n4685), .ZN(n7709) );
  NAND2_X1 U6123 ( .A1(n8916), .A2(n4379), .ZN(n4690) );
  NAND2_X1 U6124 ( .A1(n4690), .A2(n4691), .ZN(n8926) );
  NAND2_X1 U6125 ( .A1(n8898), .A2(n8899), .ZN(n5981) );
  OAI21_X2 U6126 ( .B1(n8940), .B2(n4709), .A(n4706), .ZN(n8858) );
  INV_X1 U6127 ( .A(n8850), .ZN(n4718) );
  OAI21_X1 U6128 ( .B1(n4718), .B2(n4721), .A(n4719), .ZN(n8875) );
  INV_X1 U6129 ( .A(n8847), .ZN(n4730) );
  NAND2_X1 U6130 ( .A1(n7714), .A2(n4324), .ZN(n4743) );
  NAND2_X1 U6131 ( .A1(n8667), .A2(n4747), .ZN(n4745) );
  NAND2_X1 U6132 ( .A1(n4745), .A2(n4746), .ZN(n8630) );
  INV_X1 U6133 ( .A(n4749), .ZN(n8669) );
  OAI21_X1 U6134 ( .B1(n8565), .B2(n4752), .A(n4751), .ZN(n4750) );
  NAND2_X1 U6135 ( .A1(n8750), .A2(n4902), .ZN(n8539) );
  NAND2_X1 U6136 ( .A1(n7216), .A2(n4380), .ZN(n7221) );
  INV_X1 U6137 ( .A(n4765), .ZN(n5220) );
  NAND3_X1 U6138 ( .A1(n4770), .A2(n4771), .A3(n4768), .ZN(n4767) );
  NAND2_X1 U6139 ( .A1(n4775), .A2(n5005), .ZN(n5463) );
  NAND2_X1 U6140 ( .A1(n4775), .A2(n4393), .ZN(n5009) );
  NAND2_X1 U6141 ( .A1(n5081), .A2(n4782), .ZN(n4779) );
  NAND2_X1 U6142 ( .A1(n5081), .A2(n4401), .ZN(n4776) );
  NAND3_X1 U6143 ( .A1(n4780), .A2(n4781), .A3(n4779), .ZN(n9540) );
  NAND2_X1 U6144 ( .A1(n5021), .A2(n4790), .ZN(n4789) );
  NAND2_X1 U6145 ( .A1(n5021), .A2(n4794), .ZN(n4793) );
  NAND2_X1 U6146 ( .A1(n5021), .A2(n5020), .ZN(n5525) );
  NAND2_X1 U6147 ( .A1(n4971), .A2(n4803), .ZN(n4807) );
  NAND2_X1 U6148 ( .A1(n4971), .A2(n4797), .ZN(n4796) );
  NAND2_X1 U6149 ( .A1(n4971), .A2(n4970), .ZN(n5208) );
  NAND2_X1 U6150 ( .A1(n4807), .A2(n4974), .ZN(n5192) );
  OAI211_X1 U6151 ( .C1(n9166), .C2(n4816), .A(n4813), .B(n4811), .ZN(n9414)
         );
  NAND2_X1 U6152 ( .A1(n9166), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U6153 ( .A1(n4824), .A2(n4825), .ZN(n9294) );
  NAND2_X1 U6154 ( .A1(n9182), .A2(n9102), .ZN(n9105) );
  NAND2_X1 U6155 ( .A1(n4837), .A2(n7521), .ZN(n7341) );
  NAND3_X1 U6156 ( .A1(n5055), .A2(n5361), .A3(n5428), .ZN(n5377) );
  AND2_X1 U6157 ( .A1(n4841), .A2(n5059), .ZN(n4840) );
  NAND2_X1 U6158 ( .A1(n5067), .A2(n4381), .ZN(n5075) );
  NAND2_X1 U6159 ( .A1(n5067), .A2(n5065), .ZN(n5074) );
  NAND2_X2 U6160 ( .A1(n5072), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6161 ( .A1(n6849), .A2(n4850), .ZN(n4849) );
  INV_X1 U6162 ( .A(n6168), .ZN(n6159) );
  OR2_X1 U6163 ( .A1(n4869), .A2(n6879), .ZN(n4867) );
  INV_X1 U6164 ( .A(n6925), .ZN(n4868) );
  NAND2_X1 U6165 ( .A1(n7072), .A2(n4877), .ZN(n4873) );
  INV_X1 U6166 ( .A(n7071), .ZN(n4878) );
  NAND2_X1 U6167 ( .A1(n8366), .A2(n4883), .ZN(n4880) );
  NAND2_X1 U6168 ( .A1(n4880), .A2(n4881), .ZN(n8339) );
  NAND2_X1 U6169 ( .A1(n8336), .A2(n4891), .ZN(n4888) );
  NAND2_X1 U6170 ( .A1(n4888), .A2(n4889), .ZN(n8278) );
  OAI21_X2 U6171 ( .B1(n7473), .B2(n4899), .A(n4896), .ZN(n7694) );
  NAND2_X1 U6172 ( .A1(n8950), .A2(n8949), .ZN(n8958) );
  OR2_X1 U6173 ( .A1(n8723), .A2(n9877), .ZN(n8729) );
  OR2_X1 U6174 ( .A1(n5888), .A2(n5898), .ZN(n5889) );
  AND2_X1 U6175 ( .A1(n8727), .A2(n8726), .ZN(n8728) );
  INV_X1 U6176 ( .A(n5959), .ZN(n5962) );
  INV_X1 U6177 ( .A(n5076), .ZN(n5107) );
  AND2_X1 U6178 ( .A1(n7554), .A2(n7355), .ZN(n7568) );
  INV_X1 U6179 ( .A(n5769), .ZN(n5804) );
  NAND2_X1 U6180 ( .A1(n5804), .A2(n5805), .ZN(n6684) );
  NAND2_X1 U6181 ( .A1(n5357), .A2(n8192), .ZN(n5824) );
  INV_X1 U6182 ( .A(n9331), .ZN(n9332) );
  NAND2_X1 U6183 ( .A1(n8286), .A2(n8285), .ZN(n8292) );
  NOR2_X1 U6184 ( .A1(n5815), .A2(n5814), .ZN(n5816) );
  INV_X1 U6185 ( .A(n8946), .ZN(n8950) );
  OAI211_X2 U6186 ( .C1(n6305), .C2(n7977), .A(n6176), .B(n6175), .ZN(n6876)
         );
  XNOR2_X1 U6187 ( .A(n5874), .B(n6006), .ZN(n5879) );
  AOI21_X1 U6188 ( .B1(n8948), .B2(n8947), .A(n8972), .ZN(n8949) );
  NOR2_X1 U6189 ( .A1(n8287), .A2(n4318), .ZN(n8382) );
  XNOR2_X1 U6190 ( .A(n8287), .B(n4318), .ZN(n8330) );
  NAND2_X1 U6191 ( .A1(n6171), .A2(n6170), .ZN(n6205) );
  OAI222_X1 U6192 ( .A1(n8245), .A2(n8834), .B1(P1_U3084), .B2(n8244), .C1(
        n8243), .C2(n8242), .ZN(P1_U3324) );
  INV_X1 U6193 ( .A(n8244), .ZN(n5108) );
  NAND2_X1 U6194 ( .A1(n8244), .A2(n5107), .ZN(n5367) );
  AND2_X1 U6195 ( .A1(n4970), .A2(n4969), .ZN(n4901) );
  AND4_X1 U6196 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n5741), .ZN(n4904)
         );
  OR2_X1 U6197 ( .A1(n5366), .A2(n6142), .ZN(n4905) );
  AND2_X1 U6198 ( .A1(n9969), .A2(n5070), .ZN(n4906) );
  AND2_X1 U6199 ( .A1(n4957), .A2(n4956), .ZN(n4907) );
  OR2_X1 U6200 ( .A1(n6757), .A2(n6599), .ZN(n9931) );
  NAND2_X1 U6201 ( .A1(n6546), .A2(n6596), .ZN(n9921) );
  AND2_X1 U6202 ( .A1(n9722), .A2(n5799), .ZN(n4908) );
  INV_X1 U6203 ( .A(n9377), .ZN(n9327) );
  NAND2_X1 U6204 ( .A1(n6012), .A2(n6011), .ZN(n4909) );
  NAND2_X1 U6205 ( .A1(n6000), .A2(n6001), .ZN(n4910) );
  AND2_X1 U6206 ( .A1(n7888), .A2(n7887), .ZN(n8358) );
  INV_X1 U6207 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U6208 ( .A1(n7177), .A2(n8192), .ZN(n5834) );
  INV_X1 U6209 ( .A(n9176), .ZN(n9108) );
  INV_X1 U6210 ( .A(n7603), .ZN(n7604) );
  OR2_X1 U6211 ( .A1(n8278), .A2(n8280), .ZN(n8281) );
  INV_X1 U6212 ( .A(n7870), .ZN(n6371) );
  INV_X1 U6213 ( .A(n8502), .ZN(n8109) );
  AOI22_X1 U6214 ( .A1(n4484), .A2(n9821), .B1(n8486), .B2(n8437), .ZN(n7962)
         );
  INV_X1 U6215 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U6216 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  NAND2_X1 U6217 ( .A1(n5835), .A2(n5834), .ZN(n5837) );
  INV_X1 U6218 ( .A(n5517), .ZN(n5103) );
  INV_X1 U6219 ( .A(n9205), .ZN(n9099) );
  INV_X1 U6220 ( .A(n9236), .ZN(n9128) );
  INV_X1 U6221 ( .A(n5260), .ZN(n5097) );
  INV_X1 U6222 ( .A(n7494), .ZN(n7339) );
  NAND2_X1 U6223 ( .A1(n4906), .A2(n5066), .ZN(n5071) );
  INV_X1 U6224 ( .A(n5148), .ZN(n4992) );
  INV_X1 U6225 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5059) );
  INV_X1 U6226 ( .A(n5292), .ZN(n4950) );
  INV_X1 U6227 ( .A(n7002), .ZN(n7003) );
  AOI21_X1 U6228 ( .B1(n8382), .B2(n8290), .A(n8289), .ZN(n8291) );
  NAND2_X1 U6229 ( .A1(n6725), .A2(n6724), .ZN(n6727) );
  OAI22_X1 U6230 ( .A1(n7976), .A2(n7975), .B1(n7974), .B2(n8131), .ZN(n7981)
         );
  OR2_X1 U6231 ( .A1(n7896), .A2(n6372), .ZN(n7907) );
  NAND2_X1 U6232 ( .A1(n6369), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7859) );
  OR2_X1 U6233 ( .A1(n7645), .A2(n7659), .ZN(n7653) );
  INV_X1 U6234 ( .A(n8154), .ZN(n7353) );
  INV_X1 U6235 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6434) );
  INV_X1 U6236 ( .A(n5284), .ZN(n5096) );
  NAND2_X1 U6237 ( .A1(n5100), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5171) );
  INV_X1 U6238 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5282) );
  INV_X1 U6239 ( .A(n5960), .ZN(n5961) );
  OR2_X1 U6240 ( .A1(n5544), .A2(n8954), .ZN(n5141) );
  NAND2_X1 U6241 ( .A1(n5101), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5503) );
  INV_X1 U6242 ( .A(n9417), .ZN(n9144) );
  NAND2_X1 U6243 ( .A1(n5102), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5471) );
  AOI21_X1 U6244 ( .B1(n7330), .B2(n7329), .A(n7328), .ZN(n7394) );
  NAND2_X1 U6245 ( .A1(n4977), .A2(n4976), .ZN(n4980) );
  NAND2_X1 U6246 ( .A1(n4962), .A2(n4961), .ZN(n4965) );
  XNOR2_X1 U6247 ( .A(n8745), .B(n8300), .ZN(n8386) );
  OR2_X1 U6248 ( .A1(n8259), .A2(n8258), .ZN(n8260) );
  NAND2_X1 U6249 ( .A1(n8407), .A2(n9818), .ZN(n8415) );
  OR2_X1 U6250 ( .A1(n7907), .A2(n9968), .ZN(n7929) );
  AND2_X1 U6251 ( .A1(n8769), .A2(n8625), .ZN(n7855) );
  INV_X1 U6252 ( .A(n8443), .ZN(n7356) );
  AND2_X1 U6253 ( .A1(n6234), .A2(n8173), .ZN(n6276) );
  NAND2_X1 U6254 ( .A1(n6839), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6183) );
  OR2_X1 U6255 ( .A1(n6722), .A2(n8172), .ZN(n9915) );
  OAI21_X1 U6256 ( .B1(n8946), .B2(n6041), .A(n6040), .ZN(n6042) );
  NAND2_X1 U6257 ( .A1(n5096), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5277) );
  OR2_X1 U6258 ( .A1(n5308), .A2(n5282), .ZN(n5284) );
  OR2_X1 U6259 ( .A1(n5277), .A2(n5258), .ZN(n5260) );
  AND3_X1 U6260 ( .A1(n5079), .A2(n5078), .A3(n5077), .ZN(n5771) );
  OR2_X1 U6261 ( .A1(n9022), .A2(n9021), .ZN(n9019) );
  AND2_X1 U6262 ( .A1(n6045), .A2(n6330), .ZN(n7141) );
  INV_X1 U6263 ( .A(n9411), .ZN(n5772) );
  AND2_X1 U6264 ( .A1(n5040), .A2(n5039), .ZN(n5128) );
  AND2_X1 U6265 ( .A1(n5020), .A2(n5019), .ZN(n5512) );
  INV_X1 U6266 ( .A(n8416), .ZN(n8433) );
  INV_X1 U6267 ( .A(n6770), .ZN(n6768) );
  INV_X1 U6268 ( .A(n7958), .ZN(n7934) );
  AND2_X1 U6269 ( .A1(n6272), .A2(n6271), .ZN(n9804) );
  INV_X1 U6270 ( .A(n9734), .ZN(n9802) );
  AND2_X1 U6271 ( .A1(n7799), .A2(n7671), .ZN(n8802) );
  AND2_X1 U6272 ( .A1(n6276), .A2(n6260), .ZN(n9821) );
  AND2_X1 U6273 ( .A1(n6226), .A2(n9841), .ZN(n6757) );
  INV_X1 U6274 ( .A(n9915), .ZN(n9827) );
  OR2_X1 U6275 ( .A1(n8669), .A2(n8668), .ZN(n8791) );
  AND2_X1 U6276 ( .A1(n8670), .A2(n9905), .ZN(n9877) );
  AND2_X1 U6277 ( .A1(n6545), .A2(n6754), .ZN(n6596) );
  AND2_X1 U6278 ( .A1(n6225), .A2(n6224), .ZN(n9841) );
  OAI21_X1 U6279 ( .B1(n9171), .B2(n8959), .A(n6063), .ZN(n6064) );
  AND2_X1 U6280 ( .A1(n6034), .A2(n6033), .ZN(n6041) );
  INV_X1 U6281 ( .A(n8972), .ZN(n9643) );
  INV_X1 U6282 ( .A(n8959), .ZN(n8970) );
  AND2_X1 U6283 ( .A1(n5126), .A2(n5125), .ZN(n9176) );
  OR2_X1 U6284 ( .A1(n9056), .A2(n5754), .ZN(n10154) );
  INV_X1 U6285 ( .A(n9274), .ZN(n9061) );
  INV_X1 U6286 ( .A(n9107), .ZN(n9174) );
  INV_X1 U6287 ( .A(n5633), .ZN(n9339) );
  INV_X1 U6288 ( .A(n5848), .ZN(n9626) );
  INV_X1 U6289 ( .A(n9389), .ZN(n9566) );
  NAND2_X1 U6290 ( .A1(n5804), .A2(n7293), .ZN(n6654) );
  INV_X1 U6291 ( .A(n9708), .ZN(n9485) );
  NAND2_X1 U6292 ( .A1(n5790), .A2(n5789), .ZN(n6329) );
  AND2_X1 U6293 ( .A1(n5272), .A2(n5271), .ZN(n6575) );
  XNOR2_X1 U6294 ( .A(n4938), .B(SI_7_), .ZN(n5318) );
  INV_X1 U6295 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7426) );
  OR3_X1 U6296 ( .A1(n7622), .A2(n7771), .A3(n7728), .ZN(n6262) );
  NAND2_X1 U6297 ( .A1(n6766), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8416) );
  INV_X1 U6298 ( .A(n8358), .ZN(n8562) );
  INV_X1 U6299 ( .A(n9804), .ZN(n8475) );
  INV_X1 U6300 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U6301 ( .A1(n9838), .A2(n6241), .ZN(n8704) );
  NAND2_X1 U6302 ( .A1(n6235), .A2(n7366), .ZN(n9838) );
  NOR2_X1 U6303 ( .A1(n9841), .A2(n9840), .ZN(n9854) );
  CLKBUF_X1 U6304 ( .A(n9854), .Z(n9874) );
  XNOR2_X1 U6305 ( .A(n6090), .B(n6089), .ZN(n7622) );
  INV_X1 U6306 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7803) );
  INV_X1 U6307 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7243) );
  INV_X1 U6308 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6297) );
  INV_X1 U6309 ( .A(n6064), .ZN(n6065) );
  INV_X1 U6310 ( .A(n9434), .ZN(n9203) );
  NAND2_X1 U6311 ( .A1(n5147), .A2(n5146), .ZN(n9103) );
  OR2_X1 U6312 ( .A1(n9056), .A2(n6139), .ZN(n10163) );
  OR2_X1 U6313 ( .A1(n6348), .A2(n6350), .ZN(n10162) );
  OR2_X1 U6314 ( .A1(P1_U3083), .A2(n6151), .ZN(n10167) );
  OR2_X1 U6315 ( .A1(n9605), .A2(n7347), .ZN(n9392) );
  AND2_X1 U6316 ( .A1(n9559), .A2(n7143), .ZN(n9377) );
  INV_X1 U6317 ( .A(n9595), .ZN(n9401) );
  OR2_X1 U6318 ( .A1(n6696), .A2(n7138), .ZN(n9731) );
  INV_X2 U6319 ( .A(n9731), .ZN(n9733) );
  OR2_X1 U6320 ( .A1(n6696), .A2(n6046), .ZN(n9722) );
  AND2_X1 U6321 ( .A1(n6150), .A2(n5764), .ZN(n7140) );
  XNOR2_X1 U6322 ( .A(n5762), .B(n5761), .ZN(n7759) );
  INV_X1 U6323 ( .A(n5800), .ZN(n7293) );
  INV_X1 U6324 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6438) );
  INV_X1 U6325 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6338) );
  NOR2_X1 U6326 ( .A1(n9962), .A2(n9961), .ZN(n9960) );
  AOI21_X1 U6327 ( .B1(n9578), .B2(n9724), .A(n4908), .ZN(P1_U3522) );
  INV_X1 U6328 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6289) );
  INV_X1 U6329 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6306) );
  MUX2_X1 U6330 ( .A(n6289), .B(n6306), .S(n6172), .Z(n4918) );
  XNOR2_X1 U6331 ( .A(n4918), .B(SI_2_), .ZN(n5359) );
  NAND3_X1 U6332 ( .A1(n6172), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n4913) );
  AND2_X1 U6333 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4912) );
  NAND2_X1 U6334 ( .A1(n6173), .A2(n4912), .ZN(n6192) );
  NAND2_X1 U6335 ( .A1(n4913), .A2(n6192), .ZN(n4915) );
  INV_X1 U6336 ( .A(SI_1_), .ZN(n4914) );
  XNOR2_X1 U6337 ( .A(n4915), .B(n4914), .ZN(n5340) );
  MUX2_X1 U6338 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6172), .Z(n5339) );
  NAND2_X1 U6339 ( .A1(n5340), .A2(n5339), .ZN(n4917) );
  NAND2_X1 U6340 ( .A1(n4915), .A2(SI_1_), .ZN(n4916) );
  NAND2_X1 U6341 ( .A1(n4917), .A2(n4916), .ZN(n5360) );
  INV_X1 U6342 ( .A(n4918), .ZN(n4919) );
  NAND2_X1 U6343 ( .A1(n4919), .A2(SI_2_), .ZN(n4920) );
  INV_X1 U6344 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4921) );
  INV_X1 U6345 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6307) );
  MUX2_X1 U6346 ( .A(n4921), .B(n6307), .S(n6172), .Z(n4922) );
  XNOR2_X1 U6347 ( .A(n4922), .B(SI_3_), .ZN(n5426) );
  INV_X1 U6348 ( .A(n4922), .ZN(n4923) );
  NAND2_X1 U6349 ( .A1(n4923), .A2(SI_3_), .ZN(n4924) );
  MUX2_X1 U6350 ( .A(n6297), .B(n6308), .S(n5052), .Z(n4925) );
  XNOR2_X1 U6351 ( .A(n4925), .B(SI_4_), .ZN(n5410) );
  NAND2_X1 U6352 ( .A1(n5411), .A2(n5410), .ZN(n4928) );
  INV_X1 U6353 ( .A(n4925), .ZN(n4926) );
  NAND2_X1 U6354 ( .A1(n4926), .A2(SI_4_), .ZN(n4927) );
  NAND2_X1 U6355 ( .A1(n4928), .A2(n4927), .ZN(n5376) );
  INV_X1 U6356 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4929) );
  MUX2_X1 U6357 ( .A(n4929), .B(n6317), .S(n6304), .Z(n4930) );
  XNOR2_X1 U6358 ( .A(n4930), .B(SI_5_), .ZN(n5375) );
  NAND2_X1 U6359 ( .A1(n5376), .A2(n5375), .ZN(n4933) );
  INV_X1 U6360 ( .A(n4930), .ZN(n4931) );
  NAND2_X1 U6361 ( .A1(n4931), .A2(SI_5_), .ZN(n4932) );
  MUX2_X1 U6362 ( .A(n10140), .B(n6309), .S(n6304), .Z(n4934) );
  XNOR2_X1 U6363 ( .A(n4934), .B(SI_6_), .ZN(n5400) );
  INV_X1 U6364 ( .A(n4934), .ZN(n4935) );
  NAND2_X1 U6365 ( .A1(n4935), .A2(SI_6_), .ZN(n4936) );
  MUX2_X1 U6366 ( .A(n6909), .B(n6316), .S(n6304), .Z(n4938) );
  INV_X1 U6367 ( .A(n4938), .ZN(n4939) );
  NAND2_X1 U6368 ( .A1(n4939), .A2(SI_7_), .ZN(n4940) );
  MUX2_X1 U6369 ( .A(n7011), .B(n6323), .S(n6304), .Z(n4942) );
  INV_X1 U6370 ( .A(SI_8_), .ZN(n4941) );
  INV_X1 U6371 ( .A(n4942), .ZN(n4943) );
  NAND2_X1 U6372 ( .A1(n4943), .A2(SI_8_), .ZN(n4944) );
  MUX2_X1 U6373 ( .A(n7057), .B(n6325), .S(n6304), .Z(n4947) );
  INV_X1 U6374 ( .A(SI_9_), .ZN(n4946) );
  INV_X1 U6375 ( .A(n4947), .ZN(n4948) );
  NAND2_X1 U6376 ( .A1(n4948), .A2(SI_9_), .ZN(n4949) );
  MUX2_X1 U6377 ( .A(n7078), .B(n6338), .S(n5052), .Z(n4954) );
  INV_X1 U6378 ( .A(SI_10_), .ZN(n4953) );
  NAND2_X1 U6379 ( .A1(n4954), .A2(n4953), .ZN(n4957) );
  INV_X1 U6380 ( .A(n4954), .ZN(n4955) );
  NAND2_X1 U6381 ( .A1(n4955), .A2(SI_10_), .ZN(n4956) );
  MUX2_X1 U6382 ( .A(n7243), .B(n6342), .S(n5052), .Z(n4958) );
  INV_X1 U6383 ( .A(n4958), .ZN(n4959) );
  MUX2_X1 U6384 ( .A(n10117), .B(n10104), .S(n6304), .Z(n4962) );
  INV_X1 U6385 ( .A(SI_12_), .ZN(n4961) );
  INV_X1 U6386 ( .A(n4962), .ZN(n4963) );
  NAND2_X1 U6387 ( .A1(n4963), .A2(SI_12_), .ZN(n4964) );
  MUX2_X1 U6388 ( .A(n9967), .B(n6381), .S(n5052), .Z(n4967) );
  INV_X1 U6389 ( .A(SI_13_), .ZN(n4966) );
  INV_X1 U6390 ( .A(n4967), .ZN(n4968) );
  NAND2_X1 U6391 ( .A1(n4968), .A2(SI_13_), .ZN(n4969) );
  MUX2_X1 U6392 ( .A(n6437), .B(n6438), .S(n5052), .Z(n4972) );
  INV_X1 U6393 ( .A(n4972), .ZN(n4973) );
  NAND2_X1 U6394 ( .A1(n4973), .A2(SI_14_), .ZN(n4974) );
  INV_X1 U6395 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6620) );
  INV_X1 U6396 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6621) );
  MUX2_X1 U6397 ( .A(n6620), .B(n6621), .S(n6304), .Z(n4977) );
  INV_X1 U6398 ( .A(SI_15_), .ZN(n4976) );
  INV_X1 U6399 ( .A(n4977), .ZN(n4978) );
  NAND2_X1 U6400 ( .A1(n4978), .A2(SI_15_), .ZN(n4979) );
  INV_X1 U6401 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6649) );
  MUX2_X1 U6402 ( .A(n7803), .B(n6649), .S(n5052), .Z(n4982) );
  INV_X1 U6403 ( .A(SI_16_), .ZN(n4981) );
  NAND2_X1 U6404 ( .A1(n4982), .A2(n4981), .ZN(n4985) );
  INV_X1 U6405 ( .A(n4982), .ZN(n4983) );
  NAND2_X1 U6406 ( .A1(n4983), .A2(SI_16_), .ZN(n4984) );
  INV_X1 U6407 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7809) );
  INV_X1 U6408 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4987) );
  MUX2_X1 U6409 ( .A(n7809), .B(n4987), .S(n5052), .Z(n4988) );
  INV_X1 U6410 ( .A(n4988), .ZN(n4989) );
  NAND2_X1 U6411 ( .A1(n4989), .A2(SI_17_), .ZN(n4990) );
  MUX2_X1 U6412 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6304), .Z(n4993) );
  NAND2_X1 U6413 ( .A1(n5149), .A2(n4992), .ZN(n4995) );
  NAND2_X1 U6414 ( .A1(n4993), .A2(SI_18_), .ZN(n4994) );
  INV_X1 U6415 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7833) );
  INV_X1 U6416 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7027) );
  MUX2_X1 U6417 ( .A(n7833), .B(n7027), .S(n6304), .Z(n4997) );
  INV_X1 U6418 ( .A(SI_19_), .ZN(n4996) );
  INV_X1 U6419 ( .A(n4997), .ZN(n4998) );
  NAND2_X1 U6420 ( .A1(n4998), .A2(SI_19_), .ZN(n4999) );
  NAND2_X1 U6421 ( .A1(n5000), .A2(n4999), .ZN(n5492) );
  INV_X1 U6422 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7127) );
  INV_X1 U6423 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7162) );
  MUX2_X1 U6424 ( .A(n7127), .B(n7162), .S(n6304), .Z(n5002) );
  INV_X1 U6425 ( .A(SI_20_), .ZN(n5001) );
  NAND2_X1 U6426 ( .A1(n5002), .A2(n5001), .ZN(n5005) );
  INV_X1 U6427 ( .A(n5002), .ZN(n5003) );
  NAND2_X1 U6428 ( .A1(n5003), .A2(SI_20_), .ZN(n5004) );
  INV_X1 U6429 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7259) );
  INV_X1 U6430 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7291) );
  MUX2_X1 U6431 ( .A(n7259), .B(n7291), .S(n6304), .Z(n5006) );
  XNOR2_X1 U6432 ( .A(n5006), .B(SI_21_), .ZN(n5462) );
  INV_X1 U6433 ( .A(n5006), .ZN(n5007) );
  NAND2_X1 U6434 ( .A1(n5007), .A2(SI_21_), .ZN(n5008) );
  NAND2_X1 U6435 ( .A1(n5009), .A2(n5008), .ZN(n5454) );
  INV_X1 U6436 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8191) );
  INV_X1 U6437 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7373) );
  MUX2_X1 U6438 ( .A(n8191), .B(n7373), .S(n5052), .Z(n5011) );
  INV_X1 U6439 ( .A(SI_22_), .ZN(n5010) );
  NAND2_X1 U6440 ( .A1(n5011), .A2(n5010), .ZN(n5014) );
  INV_X1 U6441 ( .A(n5011), .ZN(n5012) );
  NAND2_X1 U6442 ( .A1(n5012), .A2(SI_22_), .ZN(n5013) );
  NAND2_X1 U6443 ( .A1(n5014), .A2(n5013), .ZN(n5453) );
  INV_X1 U6444 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5015) );
  INV_X1 U6445 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7501) );
  MUX2_X1 U6446 ( .A(n5015), .B(n7501), .S(n6304), .Z(n5017) );
  INV_X1 U6447 ( .A(SI_23_), .ZN(n5016) );
  NAND2_X1 U6448 ( .A1(n5017), .A2(n5016), .ZN(n5020) );
  INV_X1 U6449 ( .A(n5017), .ZN(n5018) );
  NAND2_X1 U6450 ( .A1(n5018), .A2(SI_23_), .ZN(n5019) );
  NAND2_X1 U6451 ( .A1(n5513), .A2(n5512), .ZN(n5021) );
  INV_X1 U6452 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7621) );
  INV_X1 U6453 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7619) );
  MUX2_X1 U6454 ( .A(n7621), .B(n7619), .S(n6304), .Z(n5022) );
  XNOR2_X1 U6455 ( .A(n5022), .B(SI_24_), .ZN(n5524) );
  INV_X1 U6456 ( .A(n5524), .ZN(n5025) );
  INV_X1 U6457 ( .A(n5022), .ZN(n5023) );
  NAND2_X1 U6458 ( .A1(n5023), .A2(SI_24_), .ZN(n5024) );
  INV_X1 U6459 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7726) );
  INV_X1 U6460 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7724) );
  MUX2_X1 U6461 ( .A(n7726), .B(n7724), .S(n6304), .Z(n5026) );
  INV_X1 U6462 ( .A(SI_25_), .ZN(n10003) );
  NAND2_X1 U6463 ( .A1(n5026), .A2(n10003), .ZN(n5029) );
  INV_X1 U6464 ( .A(n5026), .ZN(n5027) );
  NAND2_X1 U6465 ( .A1(n5027), .A2(SI_25_), .ZN(n5028) );
  NAND2_X1 U6466 ( .A1(n5029), .A2(n5028), .ZN(n5537) );
  INV_X1 U6467 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7770) );
  INV_X1 U6468 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7758) );
  MUX2_X1 U6469 ( .A(n7770), .B(n7758), .S(n6304), .Z(n5031) );
  INV_X1 U6470 ( .A(SI_26_), .ZN(n5030) );
  NAND2_X1 U6471 ( .A1(n5031), .A2(n5030), .ZN(n5034) );
  INV_X1 U6472 ( .A(n5031), .ZN(n5032) );
  NAND2_X1 U6473 ( .A1(n5032), .A2(SI_26_), .ZN(n5033) );
  INV_X1 U6474 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7784) );
  INV_X1 U6475 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7787) );
  MUX2_X1 U6476 ( .A(n7784), .B(n7787), .S(n6304), .Z(n5037) );
  INV_X1 U6477 ( .A(SI_27_), .ZN(n5036) );
  NAND2_X1 U6478 ( .A1(n5037), .A2(n5036), .ZN(n5040) );
  INV_X1 U6479 ( .A(n5037), .ZN(n5038) );
  NAND2_X1 U6480 ( .A1(n5038), .A2(SI_27_), .ZN(n5039) );
  INV_X1 U6481 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5041) );
  INV_X1 U6482 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8238) );
  MUX2_X1 U6483 ( .A(n5041), .B(n8238), .S(n6304), .Z(n5043) );
  XNOR2_X1 U6484 ( .A(n5043), .B(SI_28_), .ZN(n5115) );
  INV_X1 U6485 ( .A(SI_28_), .ZN(n5042) );
  INV_X1 U6486 ( .A(SI_29_), .ZN(n5088) );
  NAND2_X1 U6487 ( .A1(n5091), .A2(n5088), .ZN(n5044) );
  MUX2_X1 U6488 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6304), .Z(n5089) );
  NAND2_X1 U6489 ( .A1(n5044), .A2(n5089), .ZN(n5046) );
  NAND2_X1 U6490 ( .A1(n5046), .A2(n5045), .ZN(n5081) );
  INV_X1 U6491 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10137) );
  INV_X1 U6492 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8217) );
  MUX2_X1 U6493 ( .A(n10137), .B(n8217), .S(n6304), .Z(n5048) );
  INV_X1 U6494 ( .A(SI_30_), .ZN(n5047) );
  NAND2_X1 U6495 ( .A1(n5048), .A2(n5047), .ZN(n5051) );
  INV_X1 U6496 ( .A(n5048), .ZN(n5049) );
  NAND2_X1 U6497 ( .A1(n5049), .A2(SI_30_), .ZN(n5050) );
  NAND2_X1 U6498 ( .A1(n5051), .A2(n5050), .ZN(n5080) );
  MUX2_X1 U6499 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n5052), .Z(n5053) );
  XNOR2_X1 U6500 ( .A(n5053), .B(SI_31_), .ZN(n5054) );
  NOR2_X1 U6501 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5063) );
  NOR2_X1 U6502 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5062) );
  NOR2_X1 U6503 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5061) );
  NAND2_X1 U6504 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5065) );
  INV_X1 U6505 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5066) );
  XNOR2_X2 U6506 ( .A(n5067), .B(n5066), .ZN(n7789) );
  INV_X1 U6507 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5068) );
  OR2_X1 U6508 ( .A1(n4320), .A2(n5068), .ZN(n5069) );
  INV_X1 U6509 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9969) );
  INV_X1 U6510 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5070) );
  INV_X1 U6511 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5073) );
  XNOR2_X2 U6512 ( .A(n5075), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U6513 ( .A1(n5350), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5079) );
  INV_X1 U6514 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8184) );
  OR2_X1 U6515 ( .A1(n5500), .A2(n8184), .ZN(n5078) );
  INV_X1 U6516 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9577) );
  OR2_X1 U6517 ( .A1(n5548), .A2(n9577), .ZN(n5077) );
  NAND2_X1 U6518 ( .A1(n8216), .A2(n5539), .ZN(n5083) );
  OR2_X1 U6519 ( .A1(n4320), .A2(n8217), .ZN(n5082) );
  INV_X1 U6520 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6521 ( .A1(n5332), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U6522 ( .A1(n5350), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5084) );
  OAI211_X1 U6523 ( .C1(n5548), .C2(n5086), .A(n5085), .B(n5084), .ZN(n9140)
         );
  INV_X1 U6524 ( .A(n9140), .ZN(n5579) );
  OR2_X1 U6525 ( .A1(n9412), .A2(n5579), .ZN(n5087) );
  NAND2_X1 U6526 ( .A1(n5682), .A2(n5087), .ZN(n5738) );
  NAND2_X1 U6527 ( .A1(n5738), .A2(n8186), .ZN(n5679) );
  XNOR2_X1 U6528 ( .A(n5089), .B(n5088), .ZN(n5090) );
  NAND2_X1 U6529 ( .A1(n8241), .A2(n5539), .ZN(n5093) );
  INV_X1 U6530 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8243) );
  OR2_X1 U6531 ( .A1(n4320), .A2(n8243), .ZN(n5092) );
  INV_X1 U6532 ( .A(n5395), .ZN(n5094) );
  NAND2_X1 U6533 ( .A1(n5094), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5326) );
  INV_X1 U6534 ( .A(n5326), .ZN(n5095) );
  NAND2_X1 U6535 ( .A1(n5095), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5308) );
  INV_X1 U6536 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5258) );
  INV_X1 U6537 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6538 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_REG3_REG_15__SCAN_IN), 
        .ZN(n5098) );
  INV_X1 U6539 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5154) );
  INV_X1 U6540 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5479) );
  INV_X1 U6541 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5457) );
  INV_X1 U6542 ( .A(n5529), .ZN(n5104) );
  NAND2_X1 U6543 ( .A1(n5104), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5542) );
  INV_X1 U6544 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8883) );
  INV_X1 U6545 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8954) );
  INV_X1 U6546 ( .A(n5141), .ZN(n5106) );
  AND2_X1 U6547 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5105) );
  NAND2_X1 U6548 ( .A1(n5106), .A2(n5105), .ZN(n5121) );
  INV_X1 U6549 ( .A(n5121), .ZN(n9145) );
  NAND2_X2 U6550 ( .A1(n5108), .A2(n5107), .ZN(n5365) );
  NAND2_X1 U6551 ( .A1(n9145), .A2(n5335), .ZN(n5114) );
  INV_X1 U6552 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6553 ( .A1(n5466), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6554 ( .A1(n5332), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5109) );
  OAI211_X1 U6555 ( .C1(n5484), .C2(n5111), .A(n5110), .B(n5109), .ZN(n5112)
         );
  INV_X1 U6556 ( .A(n5112), .ZN(n5113) );
  NAND2_X1 U6557 ( .A1(n5114), .A2(n5113), .ZN(n8974) );
  INV_X1 U6558 ( .A(n8974), .ZN(n5690) );
  OR2_X1 U6559 ( .A1(n9417), .A2(n5690), .ZN(n5127) );
  NAND2_X1 U6560 ( .A1(n7925), .A2(n5539), .ZN(n5118) );
  OR2_X1 U6561 ( .A1(n4320), .A2(n8238), .ZN(n5117) );
  INV_X1 U6562 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6060) );
  INV_X1 U6563 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5119) );
  OAI21_X1 U6564 ( .B1(n5141), .B2(n6060), .A(n5119), .ZN(n5120) );
  NAND2_X1 U6565 ( .A1(n5121), .A2(n5120), .ZN(n8205) );
  OR2_X1 U6566 ( .A1(n8205), .A2(n5365), .ZN(n5126) );
  INV_X1 U6567 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10126) );
  NAND2_X1 U6568 ( .A1(n5466), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6569 ( .A1(n5332), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5122) );
  OAI211_X1 U6570 ( .C1(n5484), .C2(n10126), .A(n5123), .B(n5122), .ZN(n5124)
         );
  INV_X1 U6571 ( .A(n5124), .ZN(n5125) );
  AND2_X1 U6572 ( .A1(n5127), .A2(n5676), .ZN(n5556) );
  INV_X1 U6573 ( .A(n5556), .ZN(n5731) );
  NAND2_X1 U6574 ( .A1(n7916), .A2(n5539), .ZN(n5131) );
  OR2_X1 U6575 ( .A1(n4320), .A2(n7787), .ZN(n5130) );
  XNOR2_X1 U6576 ( .A(n5141), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9169) );
  INV_X1 U6577 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6578 ( .A1(n5332), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6579 ( .A1(n5350), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5132) );
  OAI211_X1 U6580 ( .C1(n5548), .C2(n5134), .A(n5133), .B(n5132), .ZN(n5135)
         );
  XNOR2_X1 U6581 ( .A(n5136), .B(n5137), .ZN(n7904) );
  NAND2_X1 U6582 ( .A1(n7904), .A2(n5539), .ZN(n5139) );
  OR2_X1 U6583 ( .A1(n4320), .A2(n7758), .ZN(n5138) );
  NAND2_X1 U6584 ( .A1(n5544), .A2(n8954), .ZN(n5140) );
  NAND2_X1 U6585 ( .A1(n9187), .A2(n5335), .ZN(n5147) );
  INV_X1 U6586 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6587 ( .A1(n5332), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6588 ( .A1(n5350), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5142) );
  OAI211_X1 U6589 ( .C1(n5548), .C2(n5144), .A(n5143), .B(n5142), .ZN(n5145)
         );
  INV_X1 U6590 ( .A(n5145), .ZN(n5146) );
  XNOR2_X1 U6591 ( .A(n5149), .B(n5148), .ZN(n7820) );
  NAND2_X1 U6592 ( .A1(n7820), .A2(n5539), .ZN(n5152) );
  INV_X1 U6593 ( .A(n5150), .ZN(n5164) );
  XNOR2_X1 U6594 ( .A(n5494), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9051) );
  AOI22_X1 U6595 ( .A1(n5496), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6140), .B2(
        n9051), .ZN(n5151) );
  NAND2_X1 U6596 ( .A1(n5466), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5159) );
  INV_X1 U6597 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5153) );
  OR2_X1 U6598 ( .A1(n5484), .A2(n5153), .ZN(n5158) );
  NAND2_X1 U6599 ( .A1(n5171), .A2(n5154), .ZN(n5155) );
  NAND2_X1 U6600 ( .A1(n5501), .A2(n5155), .ZN(n9326) );
  OR2_X1 U6601 ( .A1(n5437), .A2(n9326), .ZN(n5157) );
  INV_X1 U6602 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9316) );
  OR2_X1 U6603 ( .A1(n5500), .A2(n9316), .ZN(n5156) );
  NAND2_X1 U6604 ( .A1(n9472), .A2(n8902), .ZN(n5643) );
  XNOR2_X1 U6605 ( .A(n5161), .B(n5160), .ZN(n7808) );
  NAND2_X1 U6606 ( .A1(n7808), .A2(n5539), .ZN(n5167) );
  NAND2_X1 U6607 ( .A1(n5162), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5163) );
  MUX2_X1 U6608 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5163), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n5165) );
  AND2_X1 U6609 ( .A1(n5165), .A2(n5164), .ZN(n9031) );
  AOI22_X1 U6610 ( .A1(n5496), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6140), .B2(
        n9031), .ZN(n5166) );
  NAND2_X1 U6611 ( .A1(n5466), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5176) );
  INV_X1 U6612 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n5168) );
  OR2_X1 U6613 ( .A1(n5484), .A2(n5168), .ZN(n5175) );
  INV_X1 U6614 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6615 ( .A1(n5186), .A2(n5169), .ZN(n5170) );
  NAND2_X1 U6616 ( .A1(n5171), .A2(n5170), .ZN(n9335) );
  OR2_X1 U6617 ( .A1(n5437), .A2(n9335), .ZN(n5174) );
  INV_X1 U6618 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5172) );
  OR2_X1 U6619 ( .A1(n5500), .A2(n5172), .ZN(n5173) );
  NAND2_X1 U6620 ( .A1(n9476), .A2(n9323), .ZN(n9121) );
  NAND2_X1 U6621 ( .A1(n5643), .A2(n9121), .ZN(n5636) );
  XNOR2_X1 U6622 ( .A(n5178), .B(n5177), .ZN(n7801) );
  NAND2_X1 U6623 ( .A1(n7801), .A2(n5539), .ZN(n5184) );
  NOR2_X1 U6624 ( .A1(n5179), .A2(n9535), .ZN(n5180) );
  MUX2_X1 U6625 ( .A(n9535), .B(n5180), .S(P1_IR_REG_16__SCAN_IN), .Z(n5182)
         );
  INV_X1 U6626 ( .A(n5162), .ZN(n5181) );
  OR2_X1 U6627 ( .A1(n5182), .A2(n5181), .ZN(n9023) );
  INV_X1 U6628 ( .A(n9023), .ZN(n7592) );
  AOI22_X1 U6629 ( .A1(n5496), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6140), .B2(
        n7592), .ZN(n5183) );
  NAND2_X1 U6630 ( .A1(n5350), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5190) );
  INV_X1 U6631 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7582) );
  OR2_X1 U6632 ( .A1(n5548), .A2(n7582), .ZN(n5189) );
  INV_X1 U6633 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U6634 ( .A1(n5200), .A2(n9964), .ZN(n5185) );
  NAND2_X1 U6635 ( .A1(n5186), .A2(n5185), .ZN(n9351) );
  OR2_X1 U6636 ( .A1(n5437), .A2(n9351), .ZN(n5188) );
  INV_X1 U6637 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7591) );
  OR2_X1 U6638 ( .A1(n5500), .A2(n7591), .ZN(n5187) );
  NAND2_X1 U6639 ( .A1(n9481), .A2(n9363), .ZN(n9119) );
  NOR2_X1 U6640 ( .A1(n5636), .A2(n4615), .ZN(n5447) );
  OR2_X1 U6641 ( .A1(n9481), .A2(n9363), .ZN(n5563) );
  XNOR2_X1 U6642 ( .A(n5192), .B(n5191), .ZN(n7640) );
  NAND2_X1 U6643 ( .A1(n7640), .A2(n5539), .ZN(n5197) );
  NOR2_X1 U6644 ( .A1(n5193), .A2(n9535), .ZN(n5194) );
  MUX2_X1 U6645 ( .A(n9535), .B(n5194), .S(P1_IR_REG_15__SCAN_IN), .Z(n5195)
         );
  OR2_X1 U6646 ( .A1(n5195), .A2(n5179), .ZN(n7587) );
  INV_X1 U6647 ( .A(n7587), .ZN(n7579) );
  AOI22_X1 U6648 ( .A1(n5496), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6140), .B2(
        n7579), .ZN(n5196) );
  NAND2_X1 U6649 ( .A1(n5350), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5206) );
  INV_X1 U6650 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5198) );
  OR2_X1 U6651 ( .A1(n5548), .A2(n5198), .ZN(n5205) );
  INV_X1 U6652 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5215) );
  INV_X1 U6653 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5199) );
  OAI21_X1 U6654 ( .B1(n5228), .B2(n5215), .A(n5199), .ZN(n5201) );
  NAND2_X1 U6655 ( .A1(n5201), .A2(n5200), .ZN(n9369) );
  OR2_X1 U6656 ( .A1(n5437), .A2(n9369), .ZN(n5204) );
  INV_X1 U6657 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5202) );
  OR2_X1 U6658 ( .A1(n5500), .A2(n5202), .ZN(n5203) );
  NAND4_X1 U6659 ( .A1(n5206), .A2(n5205), .A3(n5204), .A4(n5203), .ZN(n9083)
         );
  INV_X1 U6660 ( .A(n9083), .ZN(n9084) );
  OR2_X1 U6661 ( .A1(n9488), .A2(n9084), .ZN(n9118) );
  XNOR2_X1 U6662 ( .A(n5208), .B(n5207), .ZN(n7625) );
  NAND2_X1 U6663 ( .A1(n7625), .A2(n5539), .ZN(n5213) );
  NAND2_X1 U6664 ( .A1(n4385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5209) );
  MUX2_X1 U6665 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5209), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5211) );
  INV_X1 U6666 ( .A(n5193), .ZN(n5210) );
  AND2_X1 U6667 ( .A1(n5211), .A2(n5210), .ZN(n7124) );
  AOI22_X1 U6668 ( .A1(n5496), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6140), .B2(
        n7124), .ZN(n5212) );
  NAND2_X1 U6669 ( .A1(n5350), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5219) );
  INV_X1 U6670 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5214) );
  OR2_X1 U6671 ( .A1(n5548), .A2(n5214), .ZN(n5218) );
  XNOR2_X1 U6672 ( .A(n5228), .B(n5215), .ZN(n9384) );
  OR2_X1 U6673 ( .A1(n5437), .A2(n9384), .ZN(n5217) );
  INV_X1 U6674 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9385) );
  OR2_X1 U6675 ( .A1(n5500), .A2(n9385), .ZN(n5216) );
  XNOR2_X1 U6676 ( .A(n5220), .B(n4901), .ZN(n7504) );
  NAND2_X1 U6677 ( .A1(n7504), .A2(n5539), .ZN(n5225) );
  NAND2_X1 U6678 ( .A1(n5221), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5222) );
  MUX2_X1 U6679 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5222), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n5223) );
  AND2_X1 U6680 ( .A1(n5223), .A2(n4385), .ZN(n7120) );
  AOI22_X1 U6681 ( .A1(n5496), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6140), .B2(
        n7120), .ZN(n5224) );
  NAND2_X1 U6682 ( .A1(n5350), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5232) );
  INV_X1 U6683 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6704) );
  OR2_X1 U6684 ( .A1(n5548), .A2(n6704), .ZN(n5231) );
  NAND2_X1 U6685 ( .A1(n5246), .A2(n5226), .ZN(n5227) );
  NAND2_X1 U6686 ( .A1(n5228), .A2(n5227), .ZN(n9403) );
  OR2_X1 U6687 ( .A1(n5437), .A2(n9403), .ZN(n5230) );
  INV_X1 U6688 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9404) );
  OR2_X1 U6689 ( .A1(n5500), .A2(n9404), .ZN(n5229) );
  NAND4_X1 U6690 ( .A1(n5232), .A2(n5231), .A3(n5230), .A4(n5229), .ZN(n9078)
         );
  INV_X1 U6691 ( .A(n9078), .ZN(n5266) );
  NAND2_X1 U6692 ( .A1(n9612), .A2(n5266), .ZN(n9379) );
  INV_X1 U6693 ( .A(n9379), .ZN(n9113) );
  NAND2_X1 U6694 ( .A1(n9115), .A2(n9113), .ZN(n5233) );
  NAND2_X1 U6695 ( .A1(n9387), .A2(n9364), .ZN(n5564) );
  AND2_X1 U6696 ( .A1(n5233), .A2(n5564), .ZN(n5625) );
  NAND2_X1 U6697 ( .A1(n9488), .A2(n9084), .ZN(n5628) );
  XNOR2_X1 U6698 ( .A(n5235), .B(n5234), .ZN(n7454) );
  NAND2_X1 U6699 ( .A1(n7454), .A2(n5539), .ZN(n5242) );
  AND2_X1 U6700 ( .A1(n5236), .A2(n5237), .ZN(n5300) );
  INV_X1 U6701 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5238) );
  INV_X1 U6702 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6703 ( .A1(n5290), .A2(n5239), .ZN(n5269) );
  OAI21_X1 U6704 ( .B1(n5271), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5240) );
  XNOR2_X1 U6705 ( .A(n5240), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6709) );
  AOI22_X1 U6706 ( .A1(n5496), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6140), .B2(
        n6709), .ZN(n5241) );
  NAND2_X1 U6707 ( .A1(n5350), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5251) );
  INV_X1 U6708 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5243) );
  OR2_X1 U6709 ( .A1(n5548), .A2(n5243), .ZN(n5250) );
  INV_X1 U6710 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U6711 ( .A1(n5260), .A2(n5244), .ZN(n5245) );
  NAND2_X1 U6712 ( .A1(n5246), .A2(n5245), .ZN(n9592) );
  OR2_X1 U6713 ( .A1(n5437), .A2(n9592), .ZN(n5249) );
  INV_X1 U6714 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5247) );
  OR2_X1 U6715 ( .A1(n5500), .A2(n5247), .ZN(n5248) );
  NAND2_X1 U6716 ( .A1(n9596), .A2(n8977), .ZN(n9111) );
  INV_X1 U6717 ( .A(n9111), .ZN(n5267) );
  OR2_X1 U6718 ( .A1(n9596), .A2(n8977), .ZN(n5618) );
  XNOR2_X1 U6719 ( .A(n5253), .B(n5252), .ZN(n7241) );
  NAND2_X1 U6720 ( .A1(n7241), .A2(n5539), .ZN(n5256) );
  NAND2_X1 U6721 ( .A1(n5271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5254) );
  XNOR2_X1 U6722 ( .A(n5254), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6610) );
  AOI22_X1 U6723 ( .A1(n5496), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6140), .B2(
        n6610), .ZN(n5255) );
  NAND2_X1 U6724 ( .A1(n5350), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5265) );
  INV_X1 U6725 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5257) );
  OR2_X1 U6726 ( .A1(n5548), .A2(n5257), .ZN(n5264) );
  NAND2_X1 U6727 ( .A1(n5277), .A2(n5258), .ZN(n5259) );
  NAND2_X1 U6728 ( .A1(n5260), .A2(n5259), .ZN(n7752) );
  OR2_X1 U6729 ( .A1(n5437), .A2(n7752), .ZN(n5263) );
  INV_X1 U6730 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5261) );
  OR2_X1 U6731 ( .A1(n5500), .A2(n5261), .ZN(n5262) );
  NAND4_X1 U6732 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n9073)
         );
  OR2_X1 U6733 ( .A1(n9074), .A2(n9555), .ZN(n9493) );
  AND2_X1 U6734 ( .A1(n5618), .A2(n9493), .ZN(n9110) );
  OR2_X1 U6735 ( .A1(n9612), .A2(n5266), .ZN(n5619) );
  OAI211_X1 U6736 ( .C1(n5267), .C2(n9110), .A(n9115), .B(n5619), .ZN(n5623)
         );
  NAND3_X1 U6737 ( .A1(n5625), .A2(n5628), .A3(n5623), .ZN(n5316) );
  NAND2_X1 U6738 ( .A1(n5269), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5270) );
  MUX2_X1 U6739 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5270), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5272) );
  AOI22_X1 U6740 ( .A1(n5496), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6140), .B2(
        n6575), .ZN(n5273) );
  NAND2_X1 U6741 ( .A1(n5350), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5281) );
  INV_X1 U6742 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5274) );
  OR2_X1 U6743 ( .A1(n5500), .A2(n5274), .ZN(n5280) );
  INV_X1 U6744 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6745 ( .A1(n5284), .A2(n5275), .ZN(n5276) );
  NAND2_X1 U6746 ( .A1(n5277), .A2(n5276), .ZN(n9558) );
  OR2_X1 U6747 ( .A1(n5437), .A2(n9558), .ZN(n5279) );
  INV_X1 U6748 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6568) );
  OR2_X1 U6749 ( .A1(n5548), .A2(n6568), .ZN(n5278) );
  INV_X1 U6750 ( .A(n7741), .ZN(n5600) );
  NAND2_X1 U6751 ( .A1(n9561), .A2(n7746), .ZN(n5607) );
  NAND2_X1 U6752 ( .A1(n5350), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6753 ( .A1(n5308), .A2(n5282), .ZN(n5283) );
  NAND2_X1 U6754 ( .A1(n5284), .A2(n5283), .ZN(n7611) );
  OR2_X1 U6755 ( .A1(n5437), .A2(n7611), .ZN(n5288) );
  INV_X1 U6756 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5285) );
  OR2_X1 U6757 ( .A1(n5500), .A2(n5285), .ZN(n5287) );
  INV_X1 U6758 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6565) );
  OR2_X1 U6759 ( .A1(n5548), .A2(n6565), .ZN(n5286) );
  NAND4_X1 U6760 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .ZN(n8979)
         );
  INV_X1 U6761 ( .A(n8979), .ZN(n9551) );
  OR2_X1 U6762 ( .A1(n5290), .A2(n9535), .ZN(n5291) );
  XNOR2_X1 U6763 ( .A(n5291), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6642) );
  INV_X1 U6764 ( .A(n6642), .ZN(n6326) );
  XNOR2_X1 U6765 ( .A(n5293), .B(n5292), .ZN(n7056) );
  OR2_X1 U6766 ( .A1(n4320), .A2(n6325), .ZN(n5294) );
  NAND2_X1 U6767 ( .A1(n9551), .A2(n9711), .ZN(n9547) );
  AND2_X1 U6768 ( .A1(n5607), .A2(n9547), .ZN(n7739) );
  NAND2_X1 U6769 ( .A1(n9074), .A2(n9555), .ZN(n7740) );
  NAND2_X1 U6770 ( .A1(n9111), .A2(n7740), .ZN(n5620) );
  INV_X1 U6771 ( .A(n5620), .ZN(n5295) );
  OAI211_X1 U6772 ( .C1(n5600), .C2(n7739), .A(n9379), .B(n5295), .ZN(n5296)
         );
  INV_X1 U6773 ( .A(n5296), .ZN(n5297) );
  AND2_X1 U6774 ( .A1(n5297), .A2(n5564), .ZN(n5298) );
  NAND2_X1 U6775 ( .A1(n5628), .A2(n5298), .ZN(n5449) );
  XNOR2_X1 U6776 ( .A(n5299), .B(n4347), .ZN(n7009) );
  OR2_X1 U6777 ( .A1(n5341), .A2(n7009), .ZN(n5304) );
  OR2_X1 U6778 ( .A1(n4320), .A2(n6323), .ZN(n5303) );
  OR2_X1 U6779 ( .A1(n5300), .A2(n9535), .ZN(n5301) );
  XNOR2_X1 U6780 ( .A(n5301), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6573) );
  INV_X1 U6781 ( .A(n6573), .ZN(n6518) );
  OR2_X1 U6782 ( .A1(n5356), .A2(n6518), .ZN(n5302) );
  NAND2_X1 U6783 ( .A1(n5350), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5313) );
  INV_X1 U6784 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5305) );
  OR2_X1 U6785 ( .A1(n5548), .A2(n5305), .ZN(n5312) );
  INV_X1 U6786 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6787 ( .A1(n5326), .A2(n5306), .ZN(n5307) );
  NAND2_X1 U6788 ( .A1(n5308), .A2(n5307), .ZN(n7312) );
  OR2_X1 U6789 ( .A1(n5437), .A2(n7312), .ZN(n5311) );
  INV_X1 U6790 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5309) );
  OR2_X1 U6791 ( .A1(n5500), .A2(n5309), .ZN(n5310) );
  NAND4_X1 U6792 ( .A1(n5313), .A2(n5312), .A3(n5311), .A4(n5310), .ZN(n8980)
         );
  NAND2_X1 U6793 ( .A1(n9703), .A2(n8980), .ZN(n7603) );
  AND2_X1 U6794 ( .A1(n7737), .A2(n7603), .ZN(n5613) );
  AND2_X1 U6795 ( .A1(n5613), .A2(n7741), .ZN(n5314) );
  OR2_X1 U6796 ( .A1(n5449), .A2(n5314), .ZN(n5315) );
  NAND4_X1 U6797 ( .A1(n5563), .A2(n9118), .A3(n5316), .A4(n5315), .ZN(n5317)
         );
  OR2_X1 U6798 ( .A1(n9476), .A2(n9323), .ZN(n9120) );
  NAND2_X1 U6799 ( .A1(n5639), .A2(n9120), .ZN(n5635) );
  AND2_X1 U6800 ( .A1(n5635), .A2(n5643), .ZN(n9301) );
  AOI21_X1 U6801 ( .B1(n5447), .B2(n5317), .A(n9301), .ZN(n5717) );
  XNOR2_X1 U6802 ( .A(n5319), .B(n5318), .ZN(n6906) );
  OR2_X1 U6803 ( .A1(n5341), .A2(n6906), .ZN(n5323) );
  OR2_X1 U6804 ( .A1(n4320), .A2(n6316), .ZN(n5322) );
  OR2_X1 U6805 ( .A1(n5236), .A2(n9535), .ZN(n5320) );
  XNOR2_X1 U6806 ( .A(n5320), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6533) );
  INV_X1 U6807 ( .A(n6533), .ZN(n6558) );
  OR2_X1 U6808 ( .A1(n5356), .A2(n6558), .ZN(n5321) );
  NAND2_X1 U6809 ( .A1(n5350), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5331) );
  INV_X1 U6810 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6516) );
  OR2_X1 U6811 ( .A1(n5548), .A2(n6516), .ZN(n5330) );
  INV_X1 U6812 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6813 ( .A1(n5395), .A2(n5324), .ZN(n5325) );
  NAND2_X1 U6814 ( .A1(n5326), .A2(n5325), .ZN(n7333) );
  OR2_X1 U6815 ( .A1(n5437), .A2(n7333), .ZN(n5329) );
  INV_X1 U6816 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5327) );
  OR2_X1 U6817 ( .A1(n5500), .A2(n5327), .ZN(n5328) );
  NAND2_X1 U6818 ( .A1(n9697), .A2(n8981), .ZN(n5711) );
  INV_X1 U6819 ( .A(n5711), .ZN(n5606) );
  NAND2_X1 U6820 ( .A1(n5332), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6821 ( .A1(n5350), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5333) );
  AND2_X1 U6822 ( .A1(n5334), .A2(n5333), .ZN(n5338) );
  NAND2_X1 U6823 ( .A1(n5466), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5337) );
  INV_X1 U6824 ( .A(n5365), .ZN(n5335) );
  XNOR2_X1 U6825 ( .A(n5340), .B(n5339), .ZN(n6314) );
  INV_X1 U6826 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5343) );
  CLKBUF_X2 U6827 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n9541) );
  NAND2_X1 U6828 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9541), .ZN(n5342) );
  XNOR2_X1 U6829 ( .A(n5343), .B(n5342), .ZN(n9655) );
  OR2_X1 U6830 ( .A1(n5356), .A2(n9655), .ZN(n5346) );
  INV_X1 U6831 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6315) );
  OR2_X1 U6832 ( .A1(n5344), .A2(n6315), .ZN(n5345) );
  NAND2_X1 U6833 ( .A1(n5347), .A2(n5357), .ZN(n5565) );
  INV_X1 U6834 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5348) );
  OR2_X1 U6835 ( .A1(n5367), .A2(n5348), .ZN(n5353) );
  INV_X1 U6836 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6837 ( .A1(n5350), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U6838 ( .A1(n6304), .A2(SI_0_), .ZN(n5355) );
  XNOR2_X1 U6839 ( .A(n5355), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9542) );
  MUX2_X1 U6840 ( .A(n9541), .B(n9542), .S(n5356), .Z(n7144) );
  OR2_X1 U6841 ( .A1(n8987), .A2(n4531), .ZN(n6686) );
  NAND2_X1 U6842 ( .A1(n5565), .A2(n6686), .ZN(n5358) );
  XNOR2_X1 U6843 ( .A(n5360), .B(n5359), .ZN(n6305) );
  OR2_X1 U6844 ( .A1(n5341), .A2(n6305), .ZN(n5364) );
  OR2_X1 U6845 ( .A1(n4320), .A2(n6306), .ZN(n5363) );
  XNOR2_X1 U6846 ( .A(n5429), .B(n5428), .ZN(n6527) );
  OR2_X1 U6847 ( .A1(n5356), .A2(n6527), .ZN(n5362) );
  NAND2_X1 U6848 ( .A1(n5350), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5371) );
  INV_X1 U6849 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6152) );
  OR2_X1 U6850 ( .A1(n5365), .A2(n6152), .ZN(n5369) );
  INV_X1 U6851 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6142) );
  INV_X1 U6852 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6526) );
  OR2_X1 U6853 ( .A1(n5367), .A2(n6526), .ZN(n5368) );
  NAND2_X1 U6854 ( .A1(n9670), .A2(n5838), .ZN(n5703) );
  NAND2_X1 U6855 ( .A1(n7167), .A2(n5703), .ZN(n5374) );
  INV_X1 U6856 ( .A(n5838), .ZN(n5372) );
  NAND2_X1 U6857 ( .A1(n5372), .A2(n7177), .ZN(n5373) );
  XNOR2_X1 U6858 ( .A(n5376), .B(n5375), .ZN(n6853) );
  OR2_X1 U6859 ( .A1(n5341), .A2(n6853), .ZN(n5383) );
  OR2_X1 U6860 ( .A1(n4320), .A2(n6317), .ZN(n5382) );
  NAND2_X1 U6861 ( .A1(n5377), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5378) );
  MUX2_X1 U6862 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5378), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5380) );
  NAND2_X1 U6863 ( .A1(n5380), .A2(n5379), .ZN(n6595) );
  OR2_X1 U6864 ( .A1(n5356), .A2(n6595), .ZN(n5381) );
  NAND2_X1 U6865 ( .A1(n5350), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5390) );
  INV_X1 U6866 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6589) );
  INV_X1 U6867 ( .A(n5384), .ZN(n5393) );
  INV_X1 U6868 ( .A(n5385), .ZN(n5421) );
  INV_X1 U6869 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10094) );
  NAND2_X1 U6870 ( .A1(n5421), .A2(n10094), .ZN(n5386) );
  NAND2_X1 U6871 ( .A1(n5393), .A2(n5386), .ZN(n7490) );
  OR2_X1 U6872 ( .A1(n5437), .A2(n7490), .ZN(n5388) );
  INV_X1 U6873 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6530) );
  OR2_X1 U6874 ( .A1(n5500), .A2(n6530), .ZN(n5387) );
  NAND2_X1 U6875 ( .A1(n7494), .A2(n8983), .ZN(n7261) );
  INV_X1 U6876 ( .A(n7261), .ZN(n5408) );
  NAND2_X1 U6877 ( .A1(n5350), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5399) );
  INV_X1 U6878 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5391) );
  INV_X1 U6879 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7382) );
  OR2_X1 U6880 ( .A1(n5500), .A2(n7382), .ZN(n5397) );
  INV_X1 U6881 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U6882 ( .A1(n5393), .A2(n5392), .ZN(n5394) );
  NAND2_X1 U6883 ( .A1(n5395), .A2(n5394), .ZN(n9647) );
  OR2_X1 U6884 ( .A1(n5437), .A2(n9647), .ZN(n5396) );
  XNOR2_X1 U6885 ( .A(n5401), .B(n5400), .ZN(n6842) );
  OR2_X1 U6886 ( .A1(n5341), .A2(n6842), .ZN(n5407) );
  OR2_X1 U6887 ( .A1(n4320), .A2(n6309), .ZN(n5406) );
  NAND2_X1 U6888 ( .A1(n5379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5402) );
  MUX2_X1 U6889 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5402), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5403) );
  INV_X1 U6890 ( .A(n5403), .ZN(n5404) );
  NOR2_X1 U6891 ( .A1(n5404), .A2(n5236), .ZN(n6630) );
  INV_X1 U6892 ( .A(n6630), .ZN(n6512) );
  OR2_X1 U6893 ( .A1(n5356), .A2(n6512), .ZN(n5405) );
  OR2_X1 U6894 ( .A1(n8982), .A2(n9641), .ZN(n5603) );
  NAND2_X1 U6895 ( .A1(n5408), .A2(n5603), .ZN(n5409) );
  NAND2_X1 U6896 ( .A1(n9641), .A2(n8982), .ZN(n5604) );
  NAND2_X1 U6897 ( .A1(n5409), .A2(n5604), .ZN(n7328) );
  XNOR2_X1 U6898 ( .A(n5411), .B(n5410), .ZN(n6748) );
  OR2_X1 U6899 ( .A1(n5341), .A2(n6748), .ZN(n5416) );
  OR2_X1 U6900 ( .A1(n4320), .A2(n6308), .ZN(n5415) );
  OAI21_X1 U6901 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6902 ( .A1(n5429), .A2(n5412), .ZN(n5413) );
  XNOR2_X1 U6903 ( .A(n5413), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9002) );
  OR2_X1 U6904 ( .A1(n5356), .A2(n9002), .ZN(n5414) );
  NAND2_X1 U6905 ( .A1(n5466), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5425) );
  INV_X1 U6906 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5417) );
  INV_X1 U6907 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5419) );
  INV_X1 U6908 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6909 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  NAND2_X1 U6910 ( .A1(n5421), .A2(n5420), .ZN(n7534) );
  OR2_X1 U6911 ( .A1(n5437), .A2(n7534), .ZN(n5423) );
  INV_X1 U6912 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7529) );
  OR2_X1 U6913 ( .A1(n5500), .A2(n7529), .ZN(n5422) );
  NAND2_X1 U6914 ( .A1(n7535), .A2(n8984), .ZN(n7272) );
  XNOR2_X1 U6915 ( .A(n5427), .B(n5426), .ZN(n6736) );
  OR2_X1 U6916 ( .A1(n5341), .A2(n6736), .ZN(n5435) );
  OR2_X1 U6917 ( .A1(n4320), .A2(n6307), .ZN(n5434) );
  NAND2_X1 U6918 ( .A1(n5429), .A2(n5428), .ZN(n5430) );
  NAND2_X1 U6919 ( .A1(n5430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5432) );
  INV_X1 U6920 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5431) );
  OR2_X1 U6921 ( .A1(n5356), .A2(n6529), .ZN(n5433) );
  NAND2_X1 U6922 ( .A1(n5350), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5441) );
  INV_X1 U6923 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6528) );
  OR2_X1 U6924 ( .A1(n5500), .A2(n6528), .ZN(n5440) );
  INV_X1 U6925 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5436) );
  OR2_X1 U6926 ( .A1(n5437), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U6927 ( .A1(n5848), .A2(n8985), .ZN(n5586) );
  AND2_X1 U6928 ( .A1(n7272), .A2(n5586), .ZN(n5708) );
  INV_X1 U6929 ( .A(n5708), .ZN(n5442) );
  NOR2_X1 U6930 ( .A1(n7328), .A2(n5442), .ZN(n5446) );
  NAND2_X1 U6931 ( .A1(n7272), .A2(n7261), .ZN(n5591) );
  INV_X1 U6932 ( .A(n5591), .ZN(n5444) );
  OR2_X1 U6933 ( .A1(n8984), .A2(n7535), .ZN(n7265) );
  NAND2_X1 U6934 ( .A1(n7265), .A2(n5706), .ZN(n5443) );
  NAND2_X1 U6935 ( .A1(n5444), .A2(n5443), .ZN(n5445) );
  OR2_X1 U6936 ( .A1(n8983), .A2(n7494), .ZN(n7262) );
  AND2_X1 U6937 ( .A1(n5603), .A2(n7262), .ZN(n7329) );
  NAND2_X1 U6938 ( .A1(n5445), .A2(n7329), .ZN(n5568) );
  AOI22_X1 U6939 ( .A1(n5588), .A2(n5446), .B1(n5568), .B2(n5604), .ZN(n5452)
         );
  INV_X1 U6940 ( .A(n5447), .ZN(n5451) );
  INV_X1 U6941 ( .A(n7605), .ZN(n5448) );
  OR2_X1 U6942 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  NOR2_X1 U6943 ( .A1(n5451), .A2(n5450), .ZN(n5715) );
  OAI211_X1 U6944 ( .C1(n5606), .C2(n5452), .A(n5715), .B(n7395), .ZN(n5510)
         );
  XNOR2_X1 U6945 ( .A(n5454), .B(n5453), .ZN(n7856) );
  NAND2_X1 U6946 ( .A1(n7856), .A2(n5539), .ZN(n5456) );
  OR2_X1 U6947 ( .A1(n4320), .A2(n7373), .ZN(n5455) );
  NAND2_X1 U6948 ( .A1(n5471), .A2(n5457), .ZN(n5458) );
  AND2_X1 U6949 ( .A1(n5517), .A2(n5458), .ZN(n9247) );
  NAND2_X1 U6950 ( .A1(n9247), .A2(n5335), .ZN(n5461) );
  AOI22_X1 U6951 ( .A1(n5466), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n5350), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6952 ( .A1(n5332), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U6953 ( .A1(n9452), .A2(n9273), .ZN(n9127) );
  NAND2_X1 U6954 ( .A1(n7796), .A2(n5539), .ZN(n5465) );
  OR2_X1 U6955 ( .A1(n4320), .A2(n7291), .ZN(n5464) );
  NAND2_X2 U6956 ( .A1(n5465), .A2(n5464), .ZN(n9458) );
  NAND2_X1 U6957 ( .A1(n5350), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6958 ( .A1(n5466), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5467) );
  AND2_X1 U6959 ( .A1(n5468), .A2(n5467), .ZN(n5474) );
  INV_X1 U6960 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6961 ( .A1(n5481), .A2(n5469), .ZN(n5470) );
  NAND2_X1 U6962 ( .A1(n5471), .A2(n5470), .ZN(n9264) );
  OR2_X1 U6963 ( .A1(n9264), .A2(n5365), .ZN(n5473) );
  NAND2_X1 U6964 ( .A1(n5332), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5472) );
  XNOR2_X1 U6965 ( .A(n5476), .B(n5475), .ZN(n7847) );
  NAND2_X1 U6966 ( .A1(n7847), .A2(n5539), .ZN(n5478) );
  OR2_X1 U6967 ( .A1(n4320), .A2(n7162), .ZN(n5477) );
  NAND2_X1 U6968 ( .A1(n5503), .A2(n5479), .ZN(n5480) );
  AND2_X1 U6969 ( .A1(n5481), .A2(n5480), .ZN(n9282) );
  NAND2_X1 U6970 ( .A1(n5335), .A2(n9282), .ZN(n5489) );
  INV_X1 U6971 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5482) );
  OR2_X1 U6972 ( .A1(n5548), .A2(n5482), .ZN(n5488) );
  INV_X1 U6973 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n5483) );
  OR2_X1 U6974 ( .A1(n5484), .A2(n5483), .ZN(n5487) );
  INV_X1 U6975 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5485) );
  OR2_X1 U6976 ( .A1(n5500), .A2(n5485), .ZN(n5486) );
  NAND4_X1 U6977 ( .A1(n5489), .A2(n5488), .A3(n5487), .A4(n5486), .ZN(n9307)
         );
  INV_X1 U6978 ( .A(n9307), .ZN(n9092) );
  NAND2_X1 U6979 ( .A1(n9461), .A2(n9092), .ZN(n5584) );
  INV_X1 U6980 ( .A(n5584), .ZN(n5490) );
  NAND2_X1 U6981 ( .A1(n9458), .A2(n8920), .ZN(n5585) );
  AND2_X1 U6982 ( .A1(n9127), .A2(n5491), .ZN(n5648) );
  INV_X1 U6983 ( .A(n5648), .ZN(n5509) );
  XNOR2_X1 U6984 ( .A(n5493), .B(n5492), .ZN(n7831) );
  NAND2_X1 U6985 ( .A1(n7831), .A2(n5539), .ZN(n5498) );
  INV_X1 U6986 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U6987 ( .A1(n5494), .A2(n5743), .ZN(n5495) );
  XNOR2_X1 U6988 ( .A(n5558), .B(n5741), .ZN(n9274) );
  AOI22_X1 U6989 ( .A1(n5496), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9061), .B2(
        n6140), .ZN(n5497) );
  NAND2_X1 U6990 ( .A1(n5350), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5508) );
  INV_X1 U6991 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5499) );
  OR2_X1 U6992 ( .A1(n5500), .A2(n5499), .ZN(n5507) );
  INV_X1 U6993 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U6994 ( .A1(n5501), .A2(n10120), .ZN(n5502) );
  NAND2_X1 U6995 ( .A1(n5503), .A2(n5502), .ZN(n8862) );
  OR2_X1 U6996 ( .A1(n5437), .A2(n8862), .ZN(n5506) );
  INV_X1 U6997 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5504) );
  OR2_X1 U6998 ( .A1(n5548), .A2(n5504), .ZN(n5505) );
  NAND4_X1 U6999 ( .A1(n5508), .A2(n5507), .A3(n5506), .A4(n5505), .ZN(n9090)
         );
  INV_X1 U7000 ( .A(n9090), .ZN(n9322) );
  NAND2_X1 U7001 ( .A1(n9467), .A2(n9322), .ZN(n9124) );
  INV_X1 U7002 ( .A(n9124), .ZN(n5646) );
  OR2_X1 U7003 ( .A1(n5509), .A2(n5646), .ZN(n5722) );
  AOI21_X1 U7004 ( .B1(n5717), .B2(n5510), .A(n5722), .ZN(n5522) );
  OR2_X1 U7005 ( .A1(n9461), .A2(n9092), .ZN(n9125) );
  OR2_X1 U7006 ( .A1(n9467), .A2(n9322), .ZN(n5562) );
  NAND2_X1 U7007 ( .A1(n5641), .A2(n4335), .ZN(n5511) );
  NAND2_X1 U7008 ( .A1(n7867), .A2(n5539), .ZN(n5515) );
  OR2_X1 U7009 ( .A1(n4320), .A2(n7501), .ZN(n5514) );
  INV_X1 U7010 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5521) );
  INV_X1 U7011 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7012 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  NAND2_X1 U7013 ( .A1(n5529), .A2(n5518), .ZN(n8851) );
  OR2_X1 U7014 ( .A1(n8851), .A2(n5365), .ZN(n5520) );
  AOI22_X1 U7015 ( .A1(n5332), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n5350), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n5519) );
  OAI211_X1 U7016 ( .C1(n5548), .C2(n5521), .A(n5520), .B(n5519), .ZN(n9256)
         );
  INV_X1 U7017 ( .A(n9256), .ZN(n8933) );
  INV_X1 U7018 ( .A(n9216), .ZN(n5652) );
  OR2_X1 U7019 ( .A1(n9452), .A2(n9273), .ZN(n5720) );
  INV_X1 U7020 ( .A(n5720), .ZN(n5642) );
  NOR4_X1 U7021 ( .A1(n5522), .A2(n5718), .A3(n5652), .A4(n5642), .ZN(n5523)
         );
  NAND2_X1 U7022 ( .A1(n9446), .A2(n8933), .ZN(n5723) );
  INV_X1 U7023 ( .A(n5723), .ZN(n5653) );
  NOR2_X1 U7024 ( .A1(n5523), .A2(n5653), .ZN(n5552) );
  NAND2_X1 U7025 ( .A1(n7879), .A2(n5539), .ZN(n5527) );
  INV_X1 U7026 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U7027 ( .A1(n5529), .A2(n5528), .ZN(n5530) );
  NAND2_X1 U7028 ( .A1(n5542), .A2(n5530), .ZN(n9214) );
  OR2_X1 U7029 ( .A1(n9214), .A2(n5365), .ZN(n5536) );
  INV_X1 U7030 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7031 ( .A1(n5350), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7032 ( .A1(n5332), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5531) );
  OAI211_X1 U7033 ( .C1(n5533), .C2(n5548), .A(n5532), .B(n5531), .ZN(n5534)
         );
  INV_X1 U7034 ( .A(n5534), .ZN(n5535) );
  INV_X1 U7035 ( .A(n9239), .ZN(n8854) );
  NOR2_X1 U7036 ( .A1(n9225), .A2(n8854), .ZN(n9129) );
  NAND2_X1 U7037 ( .A1(n7892), .A2(n5539), .ZN(n5541) );
  NAND2_X2 U7038 ( .A1(n5541), .A2(n5540), .ZN(n9434) );
  NAND2_X1 U7039 ( .A1(n5542), .A2(n8883), .ZN(n5543) );
  NAND2_X1 U7040 ( .A1(n5544), .A2(n5543), .ZN(n8880) );
  OR2_X1 U7041 ( .A1(n8880), .A2(n5365), .ZN(n5551) );
  INV_X1 U7042 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7043 ( .A1(n5332), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7044 ( .A1(n5350), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5545) );
  OAI211_X1 U7045 ( .C1(n5548), .C2(n5547), .A(n5546), .B(n5545), .ZN(n5549)
         );
  INV_X1 U7046 ( .A(n5549), .ZN(n5550) );
  NAND2_X1 U7047 ( .A1(n9434), .A2(n9100), .ZN(n9130) );
  NAND2_X1 U7048 ( .A1(n9225), .A2(n8854), .ZN(n5657) );
  AND2_X1 U7049 ( .A1(n9130), .A2(n5657), .ZN(n5702) );
  OAI21_X1 U7050 ( .B1(n5552), .B2(n9129), .A(n5702), .ZN(n5553) );
  NAND4_X1 U7051 ( .A1(n5673), .A2(n5727), .A3(n5553), .A4(n9131), .ZN(n5557)
         );
  INV_X1 U7052 ( .A(n5673), .ZN(n9158) );
  INV_X1 U7053 ( .A(n9103), .ZN(n9175) );
  NAND2_X1 U7054 ( .A1(n9430), .A2(n9175), .ZN(n9133) );
  NAND2_X1 U7055 ( .A1(n9420), .A2(n9176), .ZN(n9136) );
  NAND2_X1 U7056 ( .A1(n9424), .A2(n8951), .ZN(n5672) );
  OAI211_X1 U7057 ( .C1(n9158), .C2(n9133), .A(n9136), .B(n5672), .ZN(n5555)
         );
  AND2_X1 U7058 ( .A1(n9417), .A2(n5690), .ZN(n5554) );
  AOI21_X1 U7059 ( .B1(n5556), .B2(n5555), .A(n5554), .ZN(n5734) );
  OAI21_X1 U7060 ( .B1(n5579), .B2(n5771), .A(n9412), .ZN(n5681) );
  OAI211_X1 U7061 ( .C1(n5731), .C2(n5557), .A(n5734), .B(n5681), .ZN(n5561)
         );
  NAND2_X1 U7062 ( .A1(n5558), .A2(n5741), .ZN(n5559) );
  INV_X1 U7063 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7064 ( .A1(n5699), .A2(n5698), .ZN(n5560) );
  XNOR2_X2 U7065 ( .A(n5596), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5800) );
  INV_X1 U7066 ( .A(n5739), .ZN(n5700) );
  AOI211_X1 U7067 ( .C1(n5679), .C2(n5561), .A(n7293), .B(n5700), .ZN(n5583)
         );
  INV_X1 U7068 ( .A(n9159), .ZN(n9135) );
  NAND2_X1 U7069 ( .A1(n5727), .A2(n9133), .ZN(n9190) );
  NAND2_X1 U7070 ( .A1(n9216), .A2(n5723), .ZN(n9236) );
  NAND2_X1 U7071 ( .A1(n5720), .A2(n9127), .ZN(n9250) );
  NAND2_X1 U7072 ( .A1(n5641), .A2(n5585), .ZN(n9262) );
  NAND2_X1 U7073 ( .A1(n9125), .A2(n5584), .ZN(n9285) );
  NAND2_X1 U7074 ( .A1(n5562), .A2(n9124), .ZN(n9300) );
  INV_X1 U7075 ( .A(n9300), .ZN(n9293) );
  NAND2_X1 U7076 ( .A1(n9120), .A2(n9121), .ZN(n5633) );
  NAND2_X1 U7077 ( .A1(n5563), .A2(n9119), .ZN(n9355) );
  NAND2_X1 U7078 ( .A1(n9115), .A2(n5564), .ZN(n9380) );
  INV_X1 U7079 ( .A(n7168), .ZN(n5567) );
  NAND2_X1 U7080 ( .A1(n4531), .A2(n8987), .ZN(n5705) );
  AND2_X1 U7081 ( .A1(n6686), .A2(n5705), .ZN(n6652) );
  NAND2_X1 U7082 ( .A1(n5565), .A2(n5704), .ZN(n6682) );
  INV_X1 U7083 ( .A(n6682), .ZN(n5566) );
  NAND4_X1 U7084 ( .A1(n5567), .A2(n6652), .A3(n5566), .A4(n5708), .ZN(n5569)
         );
  NAND2_X1 U7085 ( .A1(n7395), .A2(n5711), .ZN(n7344) );
  OR4_X1 U7086 ( .A1(n5569), .A2(n5568), .A3(n7344), .A4(n7328), .ZN(n5570) );
  NAND2_X1 U7087 ( .A1(n7741), .A2(n5607), .ZN(n9549) );
  NAND2_X1 U7088 ( .A1(n9547), .A2(n7737), .ZN(n7607) );
  NAND2_X1 U7089 ( .A1(n7605), .A2(n7603), .ZN(n7397) );
  NOR4_X1 U7090 ( .A1(n5570), .A2(n9549), .A3(n7607), .A4(n7397), .ZN(n5573)
         );
  NAND2_X1 U7091 ( .A1(n5618), .A2(n9111), .ZN(n9495) );
  INV_X1 U7092 ( .A(n9495), .ZN(n5572) );
  XNOR2_X1 U7093 ( .A(n9074), .B(n9555), .ZN(n7742) );
  INV_X1 U7094 ( .A(n7742), .ZN(n5571) );
  NAND4_X1 U7095 ( .A1(n5573), .A2(n9399), .A3(n5572), .A4(n5571), .ZN(n5574)
         );
  NOR4_X1 U7096 ( .A1(n4616), .A2(n9355), .A3(n9380), .A4(n5574), .ZN(n5575)
         );
  NAND4_X1 U7097 ( .A1(n9293), .A2(n9313), .A3(n9339), .A4(n5575), .ZN(n5576)
         );
  NOR4_X1 U7098 ( .A1(n9250), .A2(n9262), .A3(n9285), .A4(n5576), .ZN(n5577)
         );
  NAND2_X1 U7099 ( .A1(n9225), .A2(n9239), .ZN(n9097) );
  INV_X1 U7100 ( .A(n9222), .ZN(n5662) );
  NAND4_X1 U7101 ( .A1(n9205), .A2(n9128), .A3(n5577), .A4(n5662), .ZN(n5578)
         );
  NOR4_X1 U7102 ( .A1(n9135), .A2(n9174), .A3(n9190), .A4(n5578), .ZN(n5580)
         );
  XNOR2_X1 U7103 ( .A(n9417), .B(n8974), .ZN(n9109) );
  NAND2_X1 U7104 ( .A1(n9412), .A2(n5579), .ZN(n5733) );
  NAND4_X1 U7105 ( .A1(n5739), .A2(n5580), .A3(n9109), .A4(n5733), .ZN(n5581)
         );
  OAI21_X1 U7106 ( .B1(n5581), .B2(n5738), .A(n7293), .ZN(n5696) );
  INV_X1 U7107 ( .A(n5696), .ZN(n5582) );
  NOR2_X1 U7108 ( .A1(n5583), .A2(n5582), .ZN(n5697) );
  NAND2_X1 U7109 ( .A1(n5584), .A2(n9124), .ZN(n5640) );
  INV_X1 U7110 ( .A(n7153), .ZN(n5587) );
  NAND2_X1 U7111 ( .A1(n5588), .A2(n5587), .ZN(n5589) );
  INV_X1 U7112 ( .A(n7524), .ZN(n5590) );
  NAND2_X1 U7113 ( .A1(n5590), .A2(n7265), .ZN(n7273) );
  INV_X1 U7114 ( .A(n7273), .ZN(n5592) );
  INV_X1 U7115 ( .A(n7395), .ZN(n5594) );
  INV_X1 U7116 ( .A(n5603), .ZN(n5593) );
  AOI211_X1 U7117 ( .C1(n5602), .C2(n5604), .A(n5594), .B(n5593), .ZN(n5601)
         );
  INV_X1 U7118 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7119 ( .A1(n5596), .A2(n5595), .ZN(n5597) );
  NAND4_X1 U7120 ( .A1(n7737), .A2(n7603), .A3(n5711), .A4(n5689), .ZN(n5599)
         );
  NOR3_X1 U7121 ( .A1(n5601), .A2(n5600), .A3(n5599), .ZN(n5617) );
  INV_X1 U7122 ( .A(n5602), .ZN(n7377) );
  INV_X1 U7123 ( .A(n5604), .ZN(n5605) );
  INV_X1 U7124 ( .A(n5689), .ZN(n5644) );
  NAND4_X1 U7125 ( .A1(n7605), .A2(n7395), .A3(n7739), .A4(n5644), .ZN(n5611)
         );
  MUX2_X1 U7126 ( .A(n7741), .B(n5607), .S(n5689), .Z(n5610) );
  NAND2_X1 U7127 ( .A1(n7605), .A2(n9547), .ZN(n5608) );
  NAND4_X1 U7128 ( .A1(n5608), .A2(n7741), .A3(n7737), .A4(n5689), .ZN(n5609)
         );
  OAI211_X1 U7129 ( .C1(n5612), .C2(n5611), .A(n5610), .B(n5609), .ZN(n5616)
         );
  INV_X1 U7130 ( .A(n7739), .ZN(n5614) );
  NOR3_X1 U7131 ( .A1(n5614), .A2(n5613), .A3(n5689), .ZN(n5615) );
  OAI211_X1 U7132 ( .C1(n5624), .C2(n5620), .A(n5619), .B(n5618), .ZN(n5622)
         );
  INV_X1 U7133 ( .A(n9115), .ZN(n5621) );
  AOI21_X1 U7134 ( .B1(n5624), .B2(n9111), .A(n5623), .ZN(n5627) );
  INV_X1 U7135 ( .A(n5625), .ZN(n5626) );
  INV_X1 U7136 ( .A(n5628), .ZN(n5630) );
  INV_X1 U7137 ( .A(n9118), .ZN(n5629) );
  MUX2_X1 U7138 ( .A(n5630), .B(n5629), .S(n5689), .Z(n5631) );
  INV_X1 U7139 ( .A(n9481), .ZN(n9354) );
  INV_X1 U7140 ( .A(n9363), .ZN(n9085) );
  MUX2_X1 U7141 ( .A(n9481), .B(n9085), .S(n5689), .Z(n5632) );
  AOI21_X1 U7142 ( .B1(n9354), .B2(n9363), .A(n5632), .ZN(n5634) );
  MUX2_X1 U7143 ( .A(n5636), .B(n5635), .S(n5689), .Z(n5637) );
  NOR2_X1 U7144 ( .A1(n5638), .A2(n5637), .ZN(n5647) );
  INV_X1 U7145 ( .A(n5641), .ZN(n9251) );
  INV_X1 U7146 ( .A(n5643), .ZN(n5645) );
  AND2_X1 U7147 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  AOI21_X1 U7148 ( .B1(n5654), .B2(n9127), .A(n5652), .ZN(n5656) );
  AOI21_X1 U7149 ( .B1(n5654), .B2(n5720), .A(n5653), .ZN(n5655) );
  MUX2_X1 U7150 ( .A(n5656), .B(n5655), .S(n5689), .Z(n5663) );
  OAI21_X1 U7151 ( .B1(n9222), .B2(n5723), .A(n5702), .ZN(n5660) );
  INV_X1 U7152 ( .A(n5657), .ZN(n5659) );
  INV_X1 U7153 ( .A(n9129), .ZN(n5658) );
  OAI211_X1 U7154 ( .C1(n5659), .C2(n9216), .A(n9131), .B(n5658), .ZN(n5725)
         );
  MUX2_X1 U7155 ( .A(n5660), .B(n5725), .S(n5689), .Z(n5661) );
  AOI21_X2 U7156 ( .B1(n5663), .B2(n5662), .A(n5661), .ZN(n5671) );
  MUX2_X1 U7157 ( .A(n9430), .B(n9103), .S(n5689), .Z(n5665) );
  INV_X1 U7158 ( .A(n5665), .ZN(n5670) );
  MUX2_X1 U7159 ( .A(n9131), .B(n9130), .S(n5689), .Z(n5664) );
  OAI21_X1 U7160 ( .B1(n9131), .B2(n9430), .A(n9175), .ZN(n5667) );
  OAI21_X1 U7161 ( .B1(n9134), .B2(n9130), .A(n9189), .ZN(n5666) );
  MUX2_X1 U7162 ( .A(n5667), .B(n5666), .S(n5689), .Z(n5668) );
  AOI22_X1 U7163 ( .A1(n5671), .A2(n5670), .B1(n5669), .B2(n5668), .ZN(n5675)
         );
  MUX2_X1 U7164 ( .A(n5673), .B(n5672), .S(n5689), .Z(n5674) );
  OAI211_X1 U7165 ( .C1(n5675), .C2(n9174), .A(n9159), .B(n5674), .ZN(n5678)
         );
  MUX2_X1 U7166 ( .A(n9136), .B(n5676), .S(n5689), .Z(n5677) );
  NAND2_X1 U7167 ( .A1(n5678), .A2(n5677), .ZN(n5687) );
  INV_X1 U7168 ( .A(n5679), .ZN(n5680) );
  AOI21_X1 U7169 ( .B1(n5684), .B2(n8974), .A(n5680), .ZN(n5686) );
  INV_X1 U7170 ( .A(n5681), .ZN(n5683) );
  AOI22_X1 U7171 ( .A1(n5684), .A2(n9417), .B1(n5683), .B2(n5682), .ZN(n5685)
         );
  NAND3_X1 U7172 ( .A1(n5687), .A2(n9144), .A3(n5690), .ZN(n5693) );
  INV_X1 U7173 ( .A(n5688), .ZN(n5692) );
  MUX2_X1 U7174 ( .A(n9144), .B(n5690), .S(n5689), .Z(n5691) );
  NAND3_X1 U7175 ( .A1(n5693), .A2(n5692), .A3(n5691), .ZN(n5694) );
  NAND2_X1 U7176 ( .A1(n6687), .A2(n5800), .ZN(n6125) );
  NOR3_X1 U7177 ( .A1(n5700), .A2(n6687), .A3(n7293), .ZN(n5701) );
  INV_X1 U7178 ( .A(n5702), .ZN(n5729) );
  NAND4_X1 U7179 ( .A1(n5705), .A2(n5704), .A3(n5703), .A4(n5800), .ZN(n5707)
         );
  NAND2_X1 U7180 ( .A1(n5707), .A2(n5706), .ZN(n5709) );
  OAI21_X1 U7181 ( .B1(n5588), .B2(n5709), .A(n5708), .ZN(n5710) );
  NAND3_X1 U7182 ( .A1(n5710), .A2(n7329), .A3(n7265), .ZN(n5713) );
  INV_X1 U7183 ( .A(n7328), .ZN(n5712) );
  NAND3_X1 U7184 ( .A1(n5713), .A2(n5712), .A3(n5711), .ZN(n5714) );
  NAND3_X1 U7185 ( .A1(n5715), .A2(n7395), .A3(n5714), .ZN(n5716) );
  AND2_X1 U7186 ( .A1(n5717), .A2(n5716), .ZN(n5721) );
  INV_X1 U7187 ( .A(n5718), .ZN(n5719) );
  OAI211_X1 U7188 ( .C1(n5722), .C2(n5721), .A(n5720), .B(n5719), .ZN(n5724)
         );
  NAND2_X1 U7189 ( .A1(n5724), .A2(n5723), .ZN(n5728) );
  NAND2_X1 U7190 ( .A1(n5725), .A2(n9130), .ZN(n5726) );
  OAI211_X1 U7191 ( .C1(n5729), .C2(n5728), .A(n5727), .B(n5726), .ZN(n5730)
         );
  OR3_X1 U7192 ( .A1(n5731), .A2(n9174), .A3(n5730), .ZN(n5732) );
  NAND2_X1 U7193 ( .A1(n5733), .A2(n5732), .ZN(n5736) );
  INV_X1 U7194 ( .A(n5734), .ZN(n5735) );
  NOR2_X1 U7195 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  OR2_X1 U7196 ( .A1(n5738), .A2(n5737), .ZN(n5740) );
  NAND2_X1 U7197 ( .A1(n5740), .A2(n5739), .ZN(n5751) );
  NAND2_X1 U7198 ( .A1(n7164), .A2(n9274), .ZN(n6058) );
  NAND2_X1 U7199 ( .A1(n7164), .A2(n9061), .ZN(n5793) );
  NAND2_X1 U7200 ( .A1(n5751), .A2(n7152), .ZN(n5750) );
  INV_X1 U7201 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5742) );
  INV_X1 U7202 ( .A(n5748), .ZN(n5745) );
  NAND2_X1 U7203 ( .A1(n5745), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5746) );
  MUX2_X1 U7204 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5746), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5749) );
  INV_X1 U7205 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U7206 ( .A1(n5748), .A2(n5747), .ZN(n5757) );
  NAND2_X1 U7207 ( .A1(n5749), .A2(n5757), .ZN(n6148) );
  NOR2_X1 U7208 ( .A1(n6148), .A2(P1_U3084), .ZN(n5752) );
  OAI211_X1 U7209 ( .C1(n5751), .C2(n6058), .A(n5750), .B(n5752), .ZN(n5767)
         );
  INV_X1 U7210 ( .A(n5752), .ZN(n7499) );
  INV_X1 U7211 ( .A(n6125), .ZN(n6048) );
  INV_X1 U7212 ( .A(n5754), .ZN(n6139) );
  NOR2_X1 U7213 ( .A1(n5757), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7214 ( .A1(n5757), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5758) );
  MUX2_X1 U7215 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5758), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5759) );
  NAND2_X1 U7216 ( .A1(n5760), .A2(n5759), .ZN(n5787) );
  NAND2_X1 U7217 ( .A1(n5755), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5762) );
  NOR2_X1 U7218 ( .A1(n5787), .A2(n7759), .ZN(n5763) );
  NAND2_X2 U7219 ( .A1(n5786), .A2(n5763), .ZN(n6150) );
  NAND2_X1 U7220 ( .A1(n6148), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6067) );
  INV_X1 U7221 ( .A(n6067), .ZN(n5764) );
  INV_X1 U7222 ( .A(n6058), .ZN(n5792) );
  INV_X1 U7223 ( .A(n7789), .ZN(n6350) );
  NAND4_X1 U7224 ( .A1(n9304), .A2(n7140), .A3(n5792), .A4(n6350), .ZN(n5765)
         );
  OAI211_X1 U7225 ( .C1(n6687), .C2(n7499), .A(n5765), .B(P1_B_REG_SCAN_IN), 
        .ZN(n5766) );
  OAI21_X1 U7226 ( .B1(n4353), .B2(n5767), .A(n5766), .ZN(P1_U3240) );
  NAND2_X1 U7227 ( .A1(n7530), .A2(n7535), .ZN(n7531) );
  NAND2_X1 U7228 ( .A1(n7400), .A2(n9703), .ZN(n7610) );
  INV_X1 U7229 ( .A(n9596), .ZN(n5768) );
  OR2_X2 U7230 ( .A1(n9348), .A2(n9476), .ZN(n9333) );
  OR2_X2 U7231 ( .A1(n9185), .A2(n9424), .ZN(n9167) );
  NOR2_X2 U7232 ( .A1(n9167), .A2(n9420), .ZN(n9154) );
  INV_X1 U7233 ( .A(n7164), .ZN(n6688) );
  AND2_X2 U7234 ( .A1(n6650), .A2(n6058), .ZN(n9712) );
  AND2_X1 U7235 ( .A1(n6350), .A2(P1_B_REG_SCAN_IN), .ZN(n5770) );
  NOR2_X1 U7236 ( .A1(n9556), .A2(n5770), .ZN(n9141) );
  INV_X1 U7237 ( .A(n5771), .ZN(n6548) );
  AND2_X1 U7238 ( .A1(n9141), .A2(n6548), .ZN(n9411) );
  NOR4_X1 U7239 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5779) );
  NOR4_X1 U7240 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5778) );
  NOR4_X1 U7241 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5777) );
  NOR4_X1 U7242 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5776) );
  NAND4_X1 U7243 ( .A1(n5779), .A2(n5778), .A3(n5777), .A4(n5776), .ZN(n5785)
         );
  NOR2_X1 U7244 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .ZN(
        n5783) );
  NOR4_X1 U7245 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5782) );
  NOR4_X1 U7246 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5781) );
  NOR4_X1 U7247 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5780) );
  NAND4_X1 U7248 ( .A1(n5783), .A2(n5782), .A3(n5781), .A4(n5780), .ZN(n5784)
         );
  NOR2_X1 U7249 ( .A1(n5785), .A2(n5784), .ZN(n6043) );
  NAND3_X1 U7250 ( .A1(n7725), .A2(P1_B_REG_SCAN_IN), .A3(n5787), .ZN(n5790)
         );
  INV_X1 U7251 ( .A(n5787), .ZN(n5788) );
  INV_X1 U7252 ( .A(P1_B_REG_SCAN_IN), .ZN(n10106) );
  AOI21_X1 U7253 ( .B1(n5788), .B2(n10106), .A(n7759), .ZN(n5789) );
  OAI21_X1 U7254 ( .B1(n6043), .B2(n6329), .A(n7140), .ZN(n5791) );
  INV_X1 U7255 ( .A(n5791), .ZN(n5796) );
  OR2_X1 U7256 ( .A1(n6654), .A2(n5793), .ZN(n5795) );
  NAND2_X1 U7257 ( .A1(n7725), .A2(n7759), .ZN(n6330) );
  OAI21_X1 U7258 ( .B1(n6329), .B2(P1_D_REG_1__SCAN_IN), .A(n6330), .ZN(n5794)
         );
  NAND4_X1 U7259 ( .A1(n5796), .A2(n7139), .A3(n5795), .A4(n5794), .ZN(n6696)
         );
  INV_X1 U7260 ( .A(n6329), .ZN(n5797) );
  INV_X1 U7261 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U7262 ( .A1(n5797), .A2(n10122), .ZN(n5798) );
  NAND2_X1 U7263 ( .A1(n5787), .A2(n7759), .ZN(n9534) );
  NAND2_X1 U7264 ( .A1(n5798), .A2(n9534), .ZN(n7138) );
  INV_X1 U7265 ( .A(n7138), .ZN(n6046) );
  INV_X1 U7266 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5799) );
  NAND2_X2 U7267 ( .A1(n5800), .A2(n7164), .ZN(n5805) );
  NAND2_X1 U7268 ( .A1(n9434), .A2(n8192), .ZN(n5803) );
  NAND2_X1 U7269 ( .A1(n8975), .A2(n4319), .ZN(n5802) );
  NAND2_X1 U7270 ( .A1(n5803), .A2(n5802), .ZN(n5807) );
  NAND2_X1 U7271 ( .A1(n5805), .A2(n9061), .ZN(n5806) );
  XNOR2_X1 U7272 ( .A(n5807), .B(n8195), .ZN(n6027) );
  OR2_X1 U7273 ( .A1(n5769), .A2(n6058), .ZN(n5809) );
  NOR2_X1 U7274 ( .A1(n9100), .A2(n8197), .ZN(n5810) );
  AOI21_X1 U7275 ( .B1(n9434), .B2(n8199), .A(n5810), .ZN(n6025) );
  INV_X1 U7276 ( .A(n6025), .ZN(n6026) );
  INV_X1 U7277 ( .A(n9541), .ZN(n5811) );
  NOR2_X1 U7278 ( .A1(n6150), .A2(n5811), .ZN(n5812) );
  AOI21_X1 U7279 ( .B1(n4319), .B2(n7144), .A(n5812), .ZN(n5813) );
  INV_X1 U7280 ( .A(n5813), .ZN(n5817) );
  INV_X1 U7281 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7282 ( .A1(n8987), .A2(n4319), .ZN(n5819) );
  NAND2_X1 U7283 ( .A1(n7144), .A2(n8192), .ZN(n5818) );
  OAI211_X1 U7284 ( .C1(n5820), .C2(n6150), .A(n5819), .B(n5818), .ZN(n6129)
         );
  NAND2_X1 U7285 ( .A1(n6130), .A2(n6129), .ZN(n6128) );
  INV_X1 U7286 ( .A(n6129), .ZN(n5821) );
  NAND2_X1 U7287 ( .A1(n5821), .A2(n8195), .ZN(n5822) );
  NAND2_X1 U7288 ( .A1(n5823), .A2(n4319), .ZN(n5825) );
  OR2_X1 U7289 ( .A1(n8236), .A2(n5808), .ZN(n5828) );
  NAND2_X1 U7290 ( .A1(n6037), .A2(n5823), .ZN(n5827) );
  NAND2_X1 U7291 ( .A1(n5828), .A2(n5827), .ZN(n5831) );
  NAND2_X1 U7292 ( .A1(n5830), .A2(n5831), .ZN(n5829) );
  NAND2_X1 U7293 ( .A1(n6676), .A2(n5829), .ZN(n5833) );
  INV_X1 U7294 ( .A(n5830), .ZN(n6674) );
  INV_X1 U7295 ( .A(n5831), .ZN(n6675) );
  NAND2_X1 U7296 ( .A1(n6674), .A2(n6675), .ZN(n5832) );
  NAND2_X1 U7297 ( .A1(n5833), .A2(n5832), .ZN(n6818) );
  NAND2_X1 U7298 ( .A1(n5838), .A2(n4319), .ZN(n5835) );
  OR2_X1 U7299 ( .A1(n9670), .A2(n5808), .ZN(n5840) );
  NAND2_X1 U7300 ( .A1(n6037), .A2(n5838), .ZN(n5839) );
  NAND2_X1 U7301 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  XNOR2_X1 U7302 ( .A(n5843), .B(n5841), .ZN(n6819) );
  NAND2_X1 U7303 ( .A1(n6818), .A2(n6819), .ZN(n5845) );
  INV_X1 U7304 ( .A(n5841), .ZN(n5842) );
  NAND2_X1 U7305 ( .A1(n5843), .A2(n5842), .ZN(n5844) );
  NAND2_X1 U7306 ( .A1(n5845), .A2(n5844), .ZN(n9624) );
  NAND2_X1 U7307 ( .A1(n8985), .A2(n4319), .ZN(n5846) );
  OAI21_X1 U7308 ( .B1(n5848), .B2(n6035), .A(n5846), .ZN(n5847) );
  XNOR2_X1 U7309 ( .A(n5847), .B(n6006), .ZN(n5853) );
  OR2_X1 U7310 ( .A1(n5848), .A2(n5808), .ZN(n5850) );
  NAND2_X1 U7311 ( .A1(n6037), .A2(n8985), .ZN(n5849) );
  NAND2_X1 U7312 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  XNOR2_X1 U7313 ( .A(n5853), .B(n5851), .ZN(n9625) );
  NAND2_X1 U7314 ( .A1(n9624), .A2(n9625), .ZN(n5855) );
  INV_X1 U7315 ( .A(n5851), .ZN(n5852) );
  NAND2_X1 U7316 ( .A1(n5853), .A2(n5852), .ZN(n5854) );
  NAND2_X1 U7317 ( .A1(n5855), .A2(n5854), .ZN(n6248) );
  INV_X1 U7318 ( .A(n6248), .ZN(n5861) );
  NAND2_X1 U7319 ( .A1(n8984), .A2(n8199), .ZN(n5856) );
  OAI21_X1 U7320 ( .B1(n7535), .B2(n6035), .A(n5856), .ZN(n5857) );
  XNOR2_X1 U7321 ( .A(n5857), .B(n8195), .ZN(n5863) );
  OR2_X1 U7322 ( .A1(n7535), .A2(n5808), .ZN(n5859) );
  NAND2_X1 U7323 ( .A1(n6037), .A2(n8984), .ZN(n5858) );
  NAND2_X1 U7324 ( .A1(n5859), .A2(n5858), .ZN(n5862) );
  XNOR2_X1 U7325 ( .A(n5863), .B(n5862), .ZN(n6249) );
  NAND2_X1 U7326 ( .A1(n5861), .A2(n5860), .ZN(n6246) );
  NAND2_X1 U7327 ( .A1(n5863), .A2(n5862), .ZN(n5864) );
  NAND2_X1 U7328 ( .A1(n6246), .A2(n5864), .ZN(n7318) );
  OR2_X1 U7329 ( .A1(n7494), .A2(n5808), .ZN(n5866) );
  NAND2_X1 U7330 ( .A1(n6037), .A2(n8983), .ZN(n5865) );
  AND2_X1 U7331 ( .A1(n5866), .A2(n5865), .ZN(n7321) );
  NAND2_X1 U7332 ( .A1(n8983), .A2(n4319), .ZN(n5867) );
  OAI21_X1 U7333 ( .B1(n7494), .B2(n6035), .A(n5867), .ZN(n5868) );
  NAND2_X1 U7334 ( .A1(n8982), .A2(n8199), .ZN(n5869) );
  OAI21_X1 U7335 ( .B1(n9641), .B2(n6035), .A(n5869), .ZN(n5870) );
  XNOR2_X1 U7336 ( .A(n5870), .B(n6006), .ZN(n9638) );
  OR2_X1 U7337 ( .A1(n9641), .A2(n5808), .ZN(n5872) );
  NAND2_X1 U7338 ( .A1(n6037), .A2(n8982), .ZN(n5871) );
  AND2_X1 U7339 ( .A1(n5872), .A2(n5871), .ZN(n5882) );
  AOI22_X1 U7340 ( .A1(n7321), .A2(n7319), .B1(n9638), .B2(n5882), .ZN(n5896)
         );
  NAND2_X1 U7341 ( .A1(n8981), .A2(n4319), .ZN(n5873) );
  OAI21_X1 U7342 ( .B1(n9697), .B2(n6035), .A(n5873), .ZN(n5874) );
  INV_X1 U7343 ( .A(n5879), .ZN(n5877) );
  OR2_X1 U7344 ( .A1(n9697), .A2(n5808), .ZN(n5876) );
  NAND2_X1 U7345 ( .A1(n6037), .A2(n8981), .ZN(n5875) );
  NAND2_X1 U7346 ( .A1(n5876), .A2(n5875), .ZN(n5878) );
  NAND2_X1 U7347 ( .A1(n5877), .A2(n5878), .ZN(n5887) );
  INV_X1 U7348 ( .A(n5887), .ZN(n5880) );
  XNOR2_X1 U7349 ( .A(n5879), .B(n5878), .ZN(n7297) );
  AND2_X1 U7350 ( .A1(n5896), .A2(n5899), .ZN(n5881) );
  NAND2_X1 U7351 ( .A1(n7318), .A2(n5881), .ZN(n5890) );
  INV_X1 U7352 ( .A(n5899), .ZN(n5888) );
  OAI21_X1 U7353 ( .B1(n7319), .B2(n7321), .A(n5882), .ZN(n5886) );
  INV_X1 U7354 ( .A(n9638), .ZN(n5885) );
  INV_X1 U7355 ( .A(n7319), .ZN(n9636) );
  INV_X1 U7356 ( .A(n7321), .ZN(n5883) );
  INV_X1 U7357 ( .A(n5882), .ZN(n9637) );
  AND2_X1 U7358 ( .A1(n5883), .A2(n9637), .ZN(n5884) );
  AOI22_X1 U7359 ( .A1(n5886), .A2(n5885), .B1(n9636), .B2(n5884), .ZN(n7294)
         );
  AND2_X1 U7360 ( .A1(n7294), .A2(n5887), .ZN(n5898) );
  NAND2_X1 U7361 ( .A1(n5890), .A2(n5889), .ZN(n5893) );
  OR2_X1 U7362 ( .A1(n9703), .A2(n5808), .ZN(n5892) );
  NAND2_X1 U7363 ( .A1(n6037), .A2(n8980), .ZN(n5891) );
  NAND2_X1 U7364 ( .A1(n5892), .A2(n5891), .ZN(n5900) );
  NAND2_X1 U7365 ( .A1(n5893), .A2(n5900), .ZN(n7306) );
  NAND2_X1 U7366 ( .A1(n8980), .A2(n4319), .ZN(n5894) );
  OAI21_X1 U7367 ( .B1(n9703), .B2(n6035), .A(n5894), .ZN(n5895) );
  XNOR2_X1 U7368 ( .A(n5895), .B(n6006), .ZN(n7308) );
  NAND2_X1 U7369 ( .A1(n7306), .A2(n7308), .ZN(n5902) );
  NAND2_X1 U7370 ( .A1(n7318), .A2(n5896), .ZN(n7295) );
  INV_X1 U7371 ( .A(n5900), .ZN(n5897) );
  AND2_X1 U7372 ( .A1(n5898), .A2(n5897), .ZN(n5901) );
  AOI21_X2 U7373 ( .B1(n7295), .B2(n5901), .A(n4361), .ZN(n7307) );
  NAND2_X1 U7374 ( .A1(n5902), .A2(n7307), .ZN(n6068) );
  NAND2_X1 U7375 ( .A1(n9711), .A2(n8192), .ZN(n5904) );
  NAND2_X1 U7376 ( .A1(n8979), .A2(n8199), .ZN(n5903) );
  NAND2_X1 U7377 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  XNOR2_X1 U7378 ( .A(n5905), .B(n6006), .ZN(n5908) );
  NAND2_X1 U7379 ( .A1(n6037), .A2(n8979), .ZN(n5907) );
  NAND2_X1 U7380 ( .A1(n9711), .A2(n8199), .ZN(n5906) );
  AND2_X1 U7381 ( .A1(n5907), .A2(n5906), .ZN(n5909) );
  NAND2_X1 U7382 ( .A1(n5908), .A2(n5909), .ZN(n5913) );
  INV_X1 U7383 ( .A(n5908), .ZN(n5911) );
  INV_X1 U7384 ( .A(n5909), .ZN(n5910) );
  NAND2_X1 U7385 ( .A1(n5911), .A2(n5910), .ZN(n5912) );
  AND2_X1 U7386 ( .A1(n5913), .A2(n5912), .ZN(n6070) );
  NAND2_X1 U7387 ( .A1(n9561), .A2(n8192), .ZN(n5915) );
  OR2_X1 U7388 ( .A1(n7746), .A2(n5808), .ZN(n5914) );
  NAND2_X1 U7389 ( .A1(n5915), .A2(n5914), .ZN(n5916) );
  XNOR2_X1 U7390 ( .A(n5916), .B(n8195), .ZN(n5919) );
  NAND2_X1 U7391 ( .A1(n9561), .A2(n4319), .ZN(n5918) );
  OR2_X1 U7392 ( .A1(n7746), .A2(n8197), .ZN(n5917) );
  NAND2_X1 U7393 ( .A1(n5918), .A2(n5917), .ZN(n5920) );
  NAND2_X1 U7394 ( .A1(n5919), .A2(n5920), .ZN(n6106) );
  INV_X1 U7395 ( .A(n5919), .ZN(n5922) );
  INV_X1 U7396 ( .A(n5920), .ZN(n5921) );
  NAND2_X1 U7397 ( .A1(n5922), .A2(n5921), .ZN(n6105) );
  INV_X1 U7398 ( .A(n6115), .ZN(n5929) );
  NAND2_X1 U7399 ( .A1(n9074), .A2(n8192), .ZN(n5925) );
  NAND2_X1 U7400 ( .A1(n9073), .A2(n4319), .ZN(n5924) );
  NAND2_X1 U7401 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  XNOR2_X1 U7402 ( .A(n5926), .B(n6006), .ZN(n5930) );
  AND2_X1 U7403 ( .A1(n6037), .A2(n9073), .ZN(n5927) );
  AOI21_X1 U7404 ( .B1(n9074), .B2(n8199), .A(n5927), .ZN(n5931) );
  XNOR2_X1 U7405 ( .A(n5930), .B(n5931), .ZN(n6118) );
  INV_X1 U7406 ( .A(n6118), .ZN(n5928) );
  INV_X1 U7407 ( .A(n5930), .ZN(n5933) );
  INV_X1 U7408 ( .A(n5931), .ZN(n5932) );
  NAND2_X1 U7409 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  NAND2_X1 U7410 ( .A1(n9596), .A2(n8192), .ZN(n5936) );
  OR2_X1 U7411 ( .A1(n8977), .A2(n5808), .ZN(n5935) );
  NAND2_X1 U7412 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  XNOR2_X1 U7413 ( .A(n5937), .B(n6006), .ZN(n7778) );
  NOR2_X1 U7414 ( .A1(n8977), .A2(n8197), .ZN(n5938) );
  AOI21_X1 U7415 ( .B1(n9596), .B2(n8199), .A(n5938), .ZN(n5940) );
  NAND2_X1 U7416 ( .A1(n7778), .A2(n5940), .ZN(n5939) );
  INV_X1 U7417 ( .A(n7778), .ZN(n5941) );
  INV_X1 U7418 ( .A(n5940), .ZN(n7777) );
  INV_X1 U7419 ( .A(n7709), .ZN(n5948) );
  NAND2_X1 U7420 ( .A1(n9612), .A2(n8192), .ZN(n5943) );
  NAND2_X1 U7421 ( .A1(n9078), .A2(n8199), .ZN(n5942) );
  NAND2_X1 U7422 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  XNOR2_X1 U7423 ( .A(n5944), .B(n8195), .ZN(n5949) );
  NAND2_X1 U7424 ( .A1(n9612), .A2(n8199), .ZN(n5946) );
  NAND2_X1 U7425 ( .A1(n6037), .A2(n9078), .ZN(n5945) );
  NAND2_X1 U7426 ( .A1(n5946), .A2(n5945), .ZN(n5950) );
  AND2_X1 U7427 ( .A1(n5949), .A2(n5950), .ZN(n7706) );
  INV_X1 U7428 ( .A(n7706), .ZN(n5947) );
  NAND2_X1 U7429 ( .A1(n5948), .A2(n5947), .ZN(n5953) );
  INV_X1 U7430 ( .A(n5949), .ZN(n5952) );
  INV_X1 U7431 ( .A(n5950), .ZN(n5951) );
  NAND2_X1 U7432 ( .A1(n5952), .A2(n5951), .ZN(n7705) );
  NAND2_X1 U7433 ( .A1(n9387), .A2(n8192), .ZN(n5955) );
  OR2_X1 U7434 ( .A1(n9364), .A2(n5808), .ZN(n5954) );
  NAND2_X1 U7435 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  XNOR2_X1 U7436 ( .A(n5956), .B(n6006), .ZN(n5960) );
  NAND2_X1 U7437 ( .A1(n5959), .A2(n5960), .ZN(n8836) );
  NAND2_X1 U7438 ( .A1(n9387), .A2(n8199), .ZN(n5958) );
  OR2_X1 U7439 ( .A1(n9364), .A2(n8197), .ZN(n5957) );
  NAND2_X1 U7440 ( .A1(n5958), .A2(n5957), .ZN(n8839) );
  NAND2_X1 U7441 ( .A1(n8836), .A2(n8839), .ZN(n5963) );
  NAND2_X1 U7442 ( .A1(n9488), .A2(n8192), .ZN(n5965) );
  NAND2_X1 U7443 ( .A1(n9083), .A2(n8199), .ZN(n5964) );
  NAND2_X1 U7444 ( .A1(n5965), .A2(n5964), .ZN(n5966) );
  XNOR2_X1 U7445 ( .A(n5966), .B(n8195), .ZN(n8960) );
  NAND2_X1 U7446 ( .A1(n9488), .A2(n8199), .ZN(n5968) );
  NAND2_X1 U7447 ( .A1(n6037), .A2(n9083), .ZN(n5967) );
  NAND2_X1 U7448 ( .A1(n5968), .A2(n5967), .ZN(n8961) );
  NAND2_X1 U7449 ( .A1(n9481), .A2(n8192), .ZN(n5970) );
  OR2_X1 U7450 ( .A1(n9363), .A2(n5808), .ZN(n5969) );
  NAND2_X1 U7451 ( .A1(n5970), .A2(n5969), .ZN(n5971) );
  XNOR2_X1 U7452 ( .A(n5971), .B(n8195), .ZN(n5974) );
  NAND2_X1 U7453 ( .A1(n9481), .A2(n8199), .ZN(n5973) );
  OR2_X1 U7454 ( .A1(n9363), .A2(n8197), .ZN(n5972) );
  NAND2_X1 U7455 ( .A1(n5973), .A2(n5972), .ZN(n5975) );
  AND2_X1 U7456 ( .A1(n5974), .A2(n5975), .ZN(n8889) );
  INV_X1 U7457 ( .A(n5974), .ZN(n5977) );
  INV_X1 U7458 ( .A(n5975), .ZN(n5976) );
  OAI22_X1 U7459 ( .A1(n9338), .A2(n6035), .B1(n9323), .B2(n5808), .ZN(n5978)
         );
  XNOR2_X1 U7460 ( .A(n5978), .B(n8195), .ZN(n5980) );
  OAI22_X1 U7461 ( .A1(n9338), .A2(n5808), .B1(n9323), .B2(n8197), .ZN(n5979)
         );
  NAND2_X1 U7462 ( .A1(n5980), .A2(n5979), .ZN(n8899) );
  OR2_X1 U7463 ( .A1(n5980), .A2(n5979), .ZN(n8900) );
  NOR2_X1 U7464 ( .A1(n8902), .A2(n8197), .ZN(n5982) );
  AOI21_X1 U7465 ( .B1(n9472), .B2(n8199), .A(n5982), .ZN(n8938) );
  NAND2_X1 U7466 ( .A1(n9472), .A2(n8192), .ZN(n5984) );
  OR2_X1 U7467 ( .A1(n8902), .A2(n5808), .ZN(n5983) );
  NAND2_X1 U7468 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  XNOR2_X1 U7469 ( .A(n5985), .B(n8195), .ZN(n8937) );
  NAND2_X1 U7470 ( .A1(n9467), .A2(n8192), .ZN(n5987) );
  NAND2_X1 U7471 ( .A1(n9090), .A2(n8199), .ZN(n5986) );
  NAND2_X1 U7472 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  XNOR2_X1 U7473 ( .A(n5988), .B(n6006), .ZN(n5990) );
  AND2_X1 U7474 ( .A1(n6037), .A2(n9090), .ZN(n5989) );
  AOI21_X1 U7475 ( .B1(n9467), .B2(n8199), .A(n5989), .ZN(n5991) );
  NAND2_X1 U7476 ( .A1(n5990), .A2(n5991), .ZN(n5995) );
  INV_X1 U7477 ( .A(n5990), .ZN(n5993) );
  INV_X1 U7478 ( .A(n5991), .ZN(n5992) );
  NAND2_X1 U7479 ( .A1(n5993), .A2(n5992), .ZN(n5994) );
  NAND2_X1 U7480 ( .A1(n8858), .A2(n5995), .ZN(n8916) );
  NAND2_X1 U7481 ( .A1(n9461), .A2(n8192), .ZN(n5997) );
  NAND2_X1 U7482 ( .A1(n9307), .A2(n8199), .ZN(n5996) );
  NAND2_X1 U7483 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  XNOR2_X1 U7484 ( .A(n5998), .B(n6006), .ZN(n6000) );
  AND2_X1 U7485 ( .A1(n6037), .A2(n9307), .ZN(n5999) );
  AOI21_X1 U7486 ( .B1(n9461), .B2(n8199), .A(n5999), .ZN(n6001) );
  INV_X1 U7487 ( .A(n6000), .ZN(n6003) );
  INV_X1 U7488 ( .A(n6001), .ZN(n6002) );
  NAND2_X1 U7489 ( .A1(n6003), .A2(n6002), .ZN(n8917) );
  NAND2_X1 U7490 ( .A1(n9458), .A2(n8192), .ZN(n6005) );
  NAND2_X1 U7491 ( .A1(n9255), .A2(n8199), .ZN(n6004) );
  NAND2_X1 U7492 ( .A1(n6005), .A2(n6004), .ZN(n6007) );
  XNOR2_X1 U7493 ( .A(n6007), .B(n6006), .ZN(n6012) );
  INV_X1 U7494 ( .A(n6012), .ZN(n6010) );
  NOR2_X1 U7495 ( .A1(n8920), .A2(n8197), .ZN(n6008) );
  AOI21_X1 U7496 ( .B1(n9458), .B2(n8199), .A(n6008), .ZN(n6011) );
  INV_X1 U7497 ( .A(n6011), .ZN(n6009) );
  NAND2_X1 U7498 ( .A1(n6010), .A2(n6009), .ZN(n8868) );
  OR2_X1 U7499 ( .A1(n9249), .A2(n5808), .ZN(n6014) );
  OR2_X1 U7500 ( .A1(n9273), .A2(n8197), .ZN(n6013) );
  OAI22_X1 U7501 ( .A1(n9249), .A2(n6035), .B1(n9273), .B2(n5808), .ZN(n6015)
         );
  XNOR2_X1 U7502 ( .A(n6015), .B(n8195), .ZN(n8927) );
  INV_X1 U7503 ( .A(n8927), .ZN(n6016) );
  AOI21_X1 U7504 ( .B1(n8926), .B2(n4340), .A(n6016), .ZN(n6017) );
  INV_X1 U7505 ( .A(n6017), .ZN(n6019) );
  OR2_X2 U7506 ( .A1(n8926), .A2(n4340), .ZN(n6018) );
  NAND2_X1 U7507 ( .A1(n6019), .A2(n6018), .ZN(n8850) );
  AOI22_X1 U7508 ( .A1(n9446), .A2(n8192), .B1(n8199), .B2(n9256), .ZN(n6020)
         );
  XOR2_X1 U7509 ( .A(n8195), .B(n6020), .Z(n8848) );
  AOI22_X1 U7510 ( .A1(n9446), .A2(n8199), .B1(n6037), .B2(n9256), .ZN(n8847)
         );
  AOI22_X1 U7511 ( .A1(n9225), .A2(n8192), .B1(n8199), .B2(n9239), .ZN(n6021)
         );
  XNOR2_X1 U7512 ( .A(n6021), .B(n8195), .ZN(n6023) );
  AOI22_X1 U7513 ( .A1(n9225), .A2(n4319), .B1(n6037), .B2(n9239), .ZN(n6022)
         );
  NAND2_X1 U7514 ( .A1(n6023), .A2(n6022), .ZN(n6024) );
  OAI21_X1 U7515 ( .B1(n6023), .B2(n6022), .A(n6024), .ZN(n8908) );
  INV_X1 U7516 ( .A(n6024), .ZN(n8877) );
  XNOR2_X1 U7517 ( .A(n6027), .B(n6025), .ZN(n8876) );
  OAI21_X1 U7518 ( .B1(n6027), .B2(n6026), .A(n8875), .ZN(n8948) );
  AND2_X1 U7519 ( .A1(n9103), .A2(n6037), .ZN(n6028) );
  AOI21_X1 U7520 ( .B1(n9430), .B2(n8199), .A(n6028), .ZN(n6032) );
  NAND2_X1 U7521 ( .A1(n9430), .A2(n8192), .ZN(n6030) );
  NAND2_X1 U7522 ( .A1(n9103), .A2(n8199), .ZN(n6029) );
  NAND2_X1 U7523 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  XNOR2_X1 U7524 ( .A(n6031), .B(n8195), .ZN(n6034) );
  XOR2_X1 U7525 ( .A(n6032), .B(n6034), .Z(n8947) );
  INV_X1 U7526 ( .A(n6032), .ZN(n6033) );
  INV_X1 U7527 ( .A(n9424), .ZN(n9171) );
  OAI22_X1 U7528 ( .A1(n9171), .A2(n6035), .B1(n8951), .B2(n5808), .ZN(n6036)
         );
  XOR2_X1 U7529 ( .A(n8195), .B(n6036), .Z(n6039) );
  INV_X1 U7530 ( .A(n8951), .ZN(n9106) );
  AOI22_X1 U7531 ( .A1(n9424), .A2(n4319), .B1(n6037), .B2(n9106), .ZN(n6038)
         );
  NAND2_X1 U7532 ( .A1(n6039), .A2(n6038), .ZN(n8209) );
  OAI21_X1 U7533 ( .B1(n6039), .B2(n6038), .A(n8209), .ZN(n6040) );
  NOR3_X2 U7534 ( .A1(n8946), .A2(n6041), .A3(n6040), .ZN(n8215) );
  INV_X1 U7535 ( .A(n6042), .ZN(n6049) );
  AND2_X1 U7536 ( .A1(n6043), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6044) );
  OR2_X1 U7537 ( .A1(n6329), .A2(n6044), .ZN(n6045) );
  NAND2_X1 U7538 ( .A1(n6046), .A2(n7141), .ZN(n6052) );
  INV_X1 U7539 ( .A(n6052), .ZN(n6047) );
  NAND2_X1 U7540 ( .A1(n6047), .A2(n7140), .ZN(n6057) );
  OAI21_X1 U7541 ( .B1(n8215), .B2(n6049), .A(n9643), .ZN(n6066) );
  NAND2_X1 U7542 ( .A1(n6057), .A2(n9559), .ZN(n9642) );
  NAND2_X1 U7543 ( .A1(n9702), .A2(n6052), .ZN(n6055) );
  OR2_X1 U7544 ( .A1(n6654), .A2(n7164), .ZN(n7142) );
  INV_X1 U7545 ( .A(n7142), .ZN(n6051) );
  NAND2_X1 U7546 ( .A1(n6052), .A2(n6051), .ZN(n6054) );
  AND3_X1 U7547 ( .A1(n7139), .A2(n6150), .A3(n6148), .ZN(n6053) );
  NAND3_X1 U7548 ( .A1(n6055), .A2(n6054), .A3(n6053), .ZN(n6056) );
  INV_X1 U7549 ( .A(n9648), .ZN(n8930) );
  INV_X1 U7550 ( .A(n6057), .ZN(n6059) );
  OR2_X1 U7551 ( .A1(n6125), .A2(n6058), .ZN(n7346) );
  INV_X1 U7552 ( .A(n7346), .ZN(n6651) );
  NAND2_X1 U7553 ( .A1(n9633), .A2(n6139), .ZN(n7301) );
  OAI22_X1 U7554 ( .A1(n9175), .A2(n7301), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6060), .ZN(n6062) );
  NAND2_X1 U7555 ( .A1(n9633), .A2(n5754), .ZN(n8964) );
  NOR2_X1 U7556 ( .A1(n9176), .A2(n8964), .ZN(n6061) );
  AOI211_X1 U7557 ( .C1(n8930), .C2(n9169), .A(n6062), .B(n6061), .ZN(n6063)
         );
  NAND2_X1 U7558 ( .A1(n6066), .A2(n6065), .ZN(P1_U3212) );
  NOR2_X2 U7559 ( .A1(n6150), .A2(n6067), .ZN(P1_U4006) );
  OAI21_X1 U7560 ( .B1(n6070), .B2(n6068), .A(n6069), .ZN(n6071) );
  AND2_X1 U7561 ( .A1(n6071), .A2(n9643), .ZN(n6077) );
  NOR2_X1 U7562 ( .A1(n8959), .A2(n7730), .ZN(n6076) );
  NOR2_X1 U7563 ( .A1(n9648), .A2(n7611), .ZN(n6075) );
  INV_X1 U7564 ( .A(n8980), .ZN(n7299) );
  OR2_X1 U7565 ( .A1(n7301), .A2(n7299), .ZN(n6073) );
  AND2_X1 U7566 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6641) );
  INV_X1 U7567 ( .A(n6641), .ZN(n6072) );
  OAI211_X1 U7568 ( .C1(n8964), .C2(n7746), .A(n6073), .B(n6072), .ZN(n6074)
         );
  OR4_X1 U7569 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(P1_U3229)
         );
  NOR2_X1 U7570 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6081) );
  NAND4_X1 U7571 ( .A1(n6081), .A2(n6080), .A3(n6312), .A4(n6079), .ZN(n6084)
         );
  INV_X2 U7572 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6333) );
  NAND4_X1 U7573 ( .A1(n6434), .A2(n6333), .A3(n6335), .A4(n6082), .ZN(n6083)
         );
  INV_X1 U7574 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7575 ( .A1(n6197), .A2(n6086), .ZN(n6087) );
  INV_X1 U7576 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7577 ( .A1(n6104), .A2(n6103), .ZN(n6088) );
  NAND2_X1 U7578 ( .A1(n6088), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6090) );
  INV_X1 U7579 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6089) );
  NOR2_X1 U7580 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6094) );
  NOR2_X1 U7581 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6093) );
  NOR2_X1 U7582 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n6092) );
  NOR2_X1 U7583 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n6091) );
  NAND2_X1 U7584 ( .A1(n6097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6096) );
  MUX2_X1 U7585 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6096), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6098) );
  NAND2_X1 U7586 ( .A1(n6098), .A2(n6167), .ZN(n7771) );
  INV_X1 U7587 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8826) );
  OR2_X1 U7588 ( .A1(n6099), .A2(n8826), .ZN(n6101) );
  MUX2_X1 U7589 ( .A(n6101), .B(P2_IR_REG_31__SCAN_IN), .S(n6100), .Z(n6102)
         );
  NAND2_X1 U7590 ( .A1(n6102), .A2(n6097), .ZN(n7728) );
  XNOR2_X1 U7591 ( .A(n6104), .B(n6103), .ZN(n6762) );
  NAND2_X1 U7592 ( .A1(n6762), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9873) );
  NOR2_X2 U7593 ( .A1(n6262), .A2(n9873), .ZN(P2_U3966) );
  NAND2_X1 U7594 ( .A1(n6106), .A2(n6105), .ZN(n6107) );
  XNOR2_X1 U7595 ( .A(n6108), .B(n6107), .ZN(n6109) );
  NOR2_X1 U7596 ( .A1(n6109), .A2(n8972), .ZN(n6114) );
  INV_X1 U7597 ( .A(n9561), .ZN(n9570) );
  NOR2_X1 U7598 ( .A1(n8959), .A2(n9570), .ZN(n6113) );
  NOR2_X1 U7599 ( .A1(n9648), .A2(n9558), .ZN(n6112) );
  OR2_X1 U7600 ( .A1(n7301), .A2(n9551), .ZN(n6110) );
  NAND2_X1 U7601 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10165) );
  OAI211_X1 U7602 ( .C1(n8964), .C2(n9555), .A(n6110), .B(n10165), .ZN(n6111)
         );
  OR4_X1 U7603 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .ZN(P1_U3215)
         );
  INV_X1 U7604 ( .A(n6116), .ZN(n6117) );
  AOI211_X1 U7605 ( .C1(n6118), .C2(n6115), .A(n8972), .B(n6117), .ZN(n6124)
         );
  NOR2_X1 U7606 ( .A1(n8959), .A2(n9507), .ZN(n6123) );
  NOR2_X1 U7607 ( .A1(n9648), .A2(n7752), .ZN(n6122) );
  OR2_X1 U7608 ( .A1(n7301), .A2(n7746), .ZN(n6120) );
  AND2_X1 U7609 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6578) );
  INV_X1 U7610 ( .A(n6578), .ZN(n6119) );
  OAI211_X1 U7611 ( .C1(n8964), .C2(n8977), .A(n6120), .B(n6119), .ZN(n6121)
         );
  OR4_X1 U7612 ( .A1(n6124), .A2(n6123), .A3(n6122), .A4(n6121), .ZN(P1_U3234)
         );
  NAND2_X1 U7613 ( .A1(n6125), .A2(n6150), .ZN(n6126) );
  NAND2_X1 U7614 ( .A1(n6126), .A2(n6148), .ZN(n6134) );
  NAND2_X1 U7615 ( .A1(n6134), .A2(n5356), .ZN(n6127) );
  NAND2_X1 U7616 ( .A1(n6127), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AOI21_X1 U7617 ( .B1(n6350), .B2(n5348), .A(n5754), .ZN(n6349) );
  AND2_X1 U7618 ( .A1(n9541), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9652) );
  OAI21_X1 U7619 ( .B1(n6130), .B2(n6129), .A(n6128), .ZN(n6699) );
  INV_X1 U7620 ( .A(n6699), .ZN(n6131) );
  MUX2_X1 U7621 ( .A(n9652), .B(n6131), .S(n7789), .Z(n6132) );
  NAND2_X1 U7622 ( .A1(n6132), .A2(n6139), .ZN(n6133) );
  CLKBUF_X1 U7623 ( .A(P1_U4006), .Z(n8986) );
  OAI211_X1 U7624 ( .C1(n9541), .C2(n6349), .A(n6133), .B(n8986), .ZN(n9016)
         );
  INV_X1 U7625 ( .A(n9016), .ZN(n6156) );
  NAND2_X1 U7626 ( .A1(n6134), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6141) );
  OR2_X1 U7627 ( .A1(n6141), .A2(n7789), .ZN(n9056) );
  XNOR2_X1 U7628 ( .A(n6527), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6137) );
  XNOR2_X1 U7629 ( .A(n9655), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U7630 ( .A1(n9653), .A2(n9652), .ZN(n9650) );
  INV_X1 U7631 ( .A(n9655), .ZN(n6143) );
  NAND2_X1 U7632 ( .A1(n6143), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7633 ( .A1(n9650), .A2(n6135), .ZN(n6136) );
  NAND2_X1 U7634 ( .A1(n6137), .A2(n6136), .ZN(n6525) );
  OAI21_X1 U7635 ( .B1(n6137), .B2(n6136), .A(n6525), .ZN(n6138) );
  NOR2_X1 U7636 ( .A1(n10154), .A2(n6138), .ZN(n6155) );
  OR2_X1 U7637 ( .A1(n6141), .A2(n6140), .ZN(n6348) );
  MUX2_X1 U7638 ( .A(n6142), .B(P1_REG1_REG_2__SCAN_IN), .S(n6527), .Z(n6146)
         );
  XNOR2_X1 U7639 ( .A(n9655), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9662) );
  AND2_X1 U7640 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(n9541), .ZN(n9661) );
  NAND2_X1 U7641 ( .A1(n9662), .A2(n9661), .ZN(n9659) );
  NAND2_X1 U7642 ( .A1(n6143), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7643 ( .A1(n9659), .A2(n6144), .ZN(n6145) );
  NAND2_X1 U7644 ( .A1(n6146), .A2(n6145), .ZN(n8989) );
  OAI21_X1 U7645 ( .B1(n6146), .B2(n6145), .A(n8989), .ZN(n6147) );
  OAI22_X1 U7646 ( .A1(n6527), .A2(n10163), .B1(n10162), .B2(n6147), .ZN(n6154) );
  INV_X1 U7647 ( .A(n6148), .ZN(n6149) );
  NOR2_X1 U7648 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  OAI22_X1 U7649 ( .A1(n10167), .A2(n7426), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6152), .ZN(n6153) );
  OR4_X1 U7650 ( .A1(n6156), .A2(n6155), .A3(n6154), .A4(n6153), .ZN(P1_U3243)
         );
  INV_X1 U7651 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6157) );
  INV_X1 U7652 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7653 ( .A1(n6171), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6160) );
  MUX2_X1 U7654 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6160), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6161) );
  AND2_X4 U7655 ( .A1(n8239), .A2(n8833), .ZN(n7958) );
  NAND2_X1 U7656 ( .A1(n7958), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7657 ( .A1(n4341), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7658 ( .A1(n6741), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6164) );
  AND2_X2 U7659 ( .A1(n8239), .A2(n6162), .ZN(n6738) );
  NAND2_X1 U7660 ( .A1(n6738), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7661 ( .A1(n6168), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6169) );
  NAND2_X4 U7662 ( .A1(n7955), .A2(n6205), .ZN(n7832) );
  NAND2_X1 U7663 ( .A1(n6839), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6176) );
  OR2_X1 U7664 ( .A1(n6174), .A2(n8826), .ZN(n6291) );
  XNOR2_X1 U7665 ( .A(n6291), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U7666 ( .A1(n7641), .A2(n6410), .ZN(n6175) );
  NAND2_X1 U7667 ( .A1(n9820), .A2(n6797), .ZN(n8000) );
  NAND2_X1 U7668 ( .A1(n6738), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7669 ( .A1(n4341), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7670 ( .A1(n7958), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7671 ( .A1(n6741), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6179) );
  NAND3_X2 U7672 ( .A1(n6181), .A2(n6180), .A3(n6179), .ZN(n6206) );
  NAND2_X1 U7673 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6182) );
  XNOR2_X1 U7674 ( .A(n6182), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U7675 ( .A1(n7641), .A2(n6459), .ZN(n6184) );
  NAND2_X1 U7676 ( .A1(n6738), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7677 ( .A1(n4341), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7678 ( .A1(n7958), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7679 ( .A1(n6741), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6187) );
  INV_X1 U7680 ( .A(SI_0_), .ZN(n6191) );
  INV_X1 U7681 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6190) );
  OAI21_X1 U7682 ( .B1(n6304), .B2(n6191), .A(n6190), .ZN(n6193) );
  AND2_X1 U7683 ( .A1(n6193), .A2(n6192), .ZN(n8835) );
  MUX2_X1 U7684 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8835), .S(n7832), .Z(n6990) );
  NAND2_X1 U7685 ( .A1(n6899), .A2(n6990), .ZN(n6982) );
  NAND2_X1 U7686 ( .A1(n8145), .A2(n8143), .ZN(n6195) );
  INV_X1 U7687 ( .A(n6195), .ZN(n6194) );
  NAND2_X1 U7688 ( .A1(n6195), .A2(n6238), .ZN(n6196) );
  NAND2_X1 U7689 ( .A1(n6805), .A2(n6196), .ZN(n6204) );
  NAND2_X1 U7690 ( .A1(n4365), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6198) );
  XNOR2_X1 U7691 ( .A(n6198), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U7692 ( .A1(n6234), .A2(n7985), .ZN(n8171) );
  INV_X1 U7693 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7694 ( .A1(n6200), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6201) );
  MUX2_X1 U7695 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6201), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6203) );
  NAND2_X1 U7696 ( .A1(n6203), .A2(n6202), .ZN(n7128) );
  OR2_X1 U7697 ( .A1(n7260), .A2(n7128), .ZN(n7983) );
  NAND2_X1 U7698 ( .A1(n8171), .A2(n7983), .ZN(n9816) );
  NAND2_X1 U7699 ( .A1(n6204), .A2(n9816), .ZN(n6212) );
  INV_X1 U7700 ( .A(n6205), .ZN(n6260) );
  NAND2_X1 U7701 ( .A1(n7958), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7702 ( .A1(n4341), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7703 ( .A1(n6741), .A2(n9833), .ZN(n6208) );
  NAND2_X1 U7704 ( .A1(n6738), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6207) );
  AOI22_X1 U7705 ( .A1(n9821), .A2(n6206), .B1(n6771), .B2(n9818), .ZN(n6211)
         );
  NAND2_X1 U7706 ( .A1(n6212), .A2(n6211), .ZN(n6542) );
  NOR4_X1 U7707 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6221) );
  INV_X1 U7708 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9991) );
  INV_X1 U7709 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9843) );
  INV_X1 U7710 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10089) );
  INV_X1 U7711 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10092) );
  NAND4_X1 U7712 ( .A1(n9991), .A2(n9843), .A3(n10089), .A4(n10092), .ZN(n6218) );
  NOR4_X1 U7713 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6216) );
  NOR4_X1 U7714 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6215) );
  NOR4_X1 U7715 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6214) );
  NOR4_X1 U7716 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6213) );
  NAND4_X1 U7717 ( .A1(n6216), .A2(n6215), .A3(n6214), .A4(n6213), .ZN(n6217)
         );
  NOR4_X1 U7718 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        n6218), .A4(n6217), .ZN(n6220) );
  NOR4_X1 U7719 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6219) );
  NAND3_X1 U7720 ( .A1(n6221), .A2(n6220), .A3(n6219), .ZN(n6226) );
  INV_X1 U7721 ( .A(n7771), .ZN(n6225) );
  INV_X1 U7722 ( .A(P2_B_REG_SCAN_IN), .ZN(n6222) );
  XOR2_X1 U7723 ( .A(n7622), .B(n6222), .Z(n6223) );
  NAND2_X1 U7724 ( .A1(n7728), .A2(n6223), .ZN(n6224) );
  INV_X1 U7725 ( .A(n6276), .ZN(n6758) );
  OR2_X1 U7726 ( .A1(n6758), .A2(n8178), .ZN(n6227) );
  NAND2_X1 U7727 ( .A1(n7622), .A2(n7771), .ZN(n9870) );
  INV_X1 U7728 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7729 ( .A1(n9841), .A2(n6228), .ZN(n6229) );
  NAND2_X1 U7730 ( .A1(n9870), .A2(n6229), .ZN(n6755) );
  NAND3_X1 U7731 ( .A1(n6763), .A2(n6597), .A3(n6755), .ZN(n6230) );
  INV_X1 U7732 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U7733 ( .A1(n9841), .A2(n6231), .ZN(n6232) );
  NAND2_X1 U7734 ( .A1(n7771), .A2(n7728), .ZN(n9872) );
  NAND2_X1 U7735 ( .A1(n6232), .A2(n9872), .ZN(n6754) );
  INV_X1 U7736 ( .A(n6754), .ZN(n6233) );
  NAND2_X1 U7737 ( .A1(n6546), .A2(n6233), .ZN(n6235) );
  NAND2_X1 U7738 ( .A1(n6262), .A2(n6597), .ZN(n9840) );
  INV_X1 U7739 ( .A(n6234), .ZN(n8189) );
  INV_X1 U7740 ( .A(n7128), .ZN(n8172) );
  MUX2_X1 U7741 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6542), .S(n9838), .Z(n6245)
         );
  OR2_X1 U7742 ( .A1(n6235), .A2(n7985), .ZN(n7045) );
  NOR2_X2 U7743 ( .A1(n7045), .A2(n9915), .ZN(n8716) );
  INV_X1 U7744 ( .A(n8716), .ZN(n7564) );
  OAI21_X1 U7745 ( .B1(n6989), .B2(n6797), .A(n9826), .ZN(n6541) );
  INV_X1 U7746 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6280) );
  OAI22_X1 U7747 ( .A1(n7564), .A2(n6541), .B1(n6280), .B2(n7366), .ZN(n6244)
         );
  NAND2_X1 U7748 ( .A1(n6236), .A2(n8143), .ZN(n6981) );
  INV_X1 U7749 ( .A(n6899), .ZN(n6986) );
  NAND2_X1 U7750 ( .A1(n6986), .A2(n6990), .ZN(n6997) );
  NAND2_X1 U7751 ( .A1(n6981), .A2(n6997), .ZN(n6996) );
  NAND2_X1 U7752 ( .A1(n6883), .A2(n9883), .ZN(n6237) );
  NAND2_X1 U7753 ( .A1(n6996), .A2(n6237), .ZN(n6239) );
  NAND2_X1 U7754 ( .A1(n6239), .A2(n6238), .ZN(n6800) );
  OAI21_X1 U7755 ( .B1(n6239), .B2(n6238), .A(n6800), .ZN(n6544) );
  INV_X1 U7756 ( .A(n6544), .ZN(n6242) );
  NAND2_X1 U7757 ( .A1(n8173), .A2(n7128), .ZN(n6720) );
  XNOR2_X1 U7758 ( .A(n6234), .B(n6720), .ZN(n6240) );
  NAND2_X1 U7759 ( .A1(n6240), .A2(n7982), .ZN(n8670) );
  OR2_X1 U7760 ( .A1(n6720), .A2(n7982), .ZN(n7197) );
  NAND2_X1 U7761 ( .A1(n8670), .A2(n7197), .ZN(n9824) );
  OR2_X1 U7762 ( .A1(n6722), .A2(n7128), .ZN(n6767) );
  INV_X1 U7763 ( .A(n6767), .ZN(n6241) );
  OAI22_X1 U7764 ( .A1(n6242), .A2(n8718), .B1(n8704), .B2(n6797), .ZN(n6243)
         );
  OR3_X1 U7765 ( .A1(n6245), .A2(n6244), .A3(n6243), .ZN(P2_U3294) );
  INV_X1 U7766 ( .A(n6246), .ZN(n6247) );
  AOI211_X1 U7767 ( .C1(n6249), .C2(n6248), .A(n8972), .B(n6247), .ZN(n6256)
         );
  NOR2_X1 U7768 ( .A1(n9648), .A2(n7534), .ZN(n6255) );
  INV_X1 U7769 ( .A(n8985), .ZN(n6251) );
  AND2_X1 U7770 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9013) );
  INV_X1 U7771 ( .A(n9013), .ZN(n6250) );
  OAI21_X1 U7772 ( .B1(n7301), .B2(n6251), .A(n6250), .ZN(n6254) );
  INV_X1 U7773 ( .A(n8983), .ZN(n6252) );
  OAI22_X1 U7774 ( .A1(n8964), .A2(n6252), .B1(n7535), .B2(n8959), .ZN(n6253)
         );
  OR4_X1 U7775 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(P1_U3228)
         );
  INV_X1 U7776 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6257) );
  MUX2_X1 U7777 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6257), .S(n6459), .Z(n6461)
         );
  AND2_X1 U7778 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6462) );
  NAND2_X1 U7779 ( .A1(n6461), .A2(n6462), .ZN(n6460) );
  NAND2_X1 U7780 ( .A1(n6459), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6258) );
  AND2_X1 U7781 ( .A1(n6460), .A2(n6258), .ZN(n6269) );
  INV_X1 U7782 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6259) );
  MUX2_X1 U7783 ( .A(n6259), .B(P2_REG2_REG_2__SCAN_IN), .S(n6410), .Z(n6268)
         );
  NOR2_X1 U7784 ( .A1(n6269), .A2(n6268), .ZN(n6409) );
  NAND2_X1 U7785 ( .A1(n6260), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7786) );
  OR2_X1 U7786 ( .A1(n6762), .A2(P2_U3152), .ZN(n8183) );
  OAI21_X1 U7787 ( .B1(n6262), .B2(n7786), .A(n8183), .ZN(n6263) );
  INV_X1 U7788 ( .A(n6263), .ZN(n6265) );
  OR2_X1 U7789 ( .A1(n9840), .A2(n6276), .ZN(n6264) );
  NAND2_X1 U7790 ( .A1(n6265), .A2(n6264), .ZN(n6272) );
  NAND2_X1 U7791 ( .A1(n6272), .A2(n7832), .ZN(n6266) );
  INV_X2 U7792 ( .A(P2_U3966), .ZN(n8448) );
  NAND2_X1 U7793 ( .A1(n6266), .A2(n8448), .ZN(n6275) );
  NOR2_X1 U7794 ( .A1(n6205), .A2(n7955), .ZN(n6267) );
  NAND2_X1 U7795 ( .A1(n6275), .A2(n6267), .ZN(n9736) );
  AOI211_X1 U7796 ( .C1(n6269), .C2(n6268), .A(n6409), .B(n9736), .ZN(n6285)
         );
  INV_X1 U7797 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9925) );
  XNOR2_X1 U7798 ( .A(n6459), .B(n9925), .ZN(n6455) );
  AND2_X1 U7799 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n6454) );
  NAND2_X1 U7800 ( .A1(n6455), .A2(n6454), .ZN(n6453) );
  NAND2_X1 U7801 ( .A1(n6459), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6270) );
  AND2_X1 U7802 ( .A1(n6453), .A2(n6270), .ZN(n6274) );
  INV_X1 U7803 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6602) );
  MUX2_X1 U7804 ( .A(n6602), .B(P2_REG1_REG_2__SCAN_IN), .S(n6410), .Z(n6273)
         );
  NOR2_X1 U7805 ( .A1(n6273), .A2(n6274), .ZN(n6388) );
  AND2_X1 U7806 ( .A1(n7832), .A2(n7955), .ZN(n6271) );
  AOI211_X1 U7807 ( .C1(n6274), .C2(n6273), .A(n6388), .B(n8475), .ZN(n6284)
         );
  NAND2_X1 U7808 ( .A1(n6275), .A2(n6205), .ZN(n9734) );
  INV_X1 U7809 ( .A(n6410), .ZN(n6288) );
  NOR2_X1 U7810 ( .A1(n9734), .A2(n6288), .ZN(n6283) );
  NOR2_X1 U7811 ( .A1(n6276), .A2(n7641), .ZN(n6277) );
  OR2_X1 U7812 ( .A1(n9840), .A2(n6277), .ZN(n6279) );
  OR2_X1 U7813 ( .A1(n8183), .A2(n7832), .ZN(n6278) );
  AND2_X1 U7814 ( .A1(n6279), .A2(n6278), .ZN(n8484) );
  INV_X1 U7815 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6281) );
  OAI22_X1 U7816 ( .A1(n8484), .A2(n6281), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6280), .ZN(n6282) );
  OR4_X1 U7817 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(P2_U3247)
         );
  AND2_X1 U7818 ( .A1(n6304), .A2(P2_U3152), .ZN(n8828) );
  AOI22_X1 U7819 ( .A1(n8828), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n6459), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6287) );
  OAI21_X1 U7820 ( .B1(n6314), .B2(n8830), .A(n6287), .ZN(P2_U3357) );
  INV_X1 U7821 ( .A(n8828), .ZN(n8831) );
  OAI222_X1 U7822 ( .A1(n8831), .A2(n6289), .B1(n8830), .B2(n6305), .C1(
        P2_U3152), .C2(n6288), .ZN(P2_U3356) );
  INV_X1 U7823 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7824 ( .A1(n6291), .A2(n6290), .ZN(n6292) );
  NAND2_X1 U7825 ( .A1(n6292), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6293) );
  XNOR2_X1 U7826 ( .A(n6293), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9742) );
  AOI22_X1 U7827 ( .A1(n9742), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n8828), .ZN(n6294) );
  OAI21_X1 U7828 ( .B1(n6736), .B2(n8830), .A(n6294), .ZN(P2_U3355) );
  NAND2_X1 U7829 ( .A1(n6295), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6296) );
  XNOR2_X1 U7830 ( .A(n6296), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9757) );
  INV_X1 U7831 ( .A(n9757), .ZN(n6412) );
  OAI222_X1 U7832 ( .A1(n8831), .A2(n6297), .B1(n8830), .B2(n6748), .C1(
        P2_U3152), .C2(n6412), .ZN(P2_U3354) );
  NAND2_X1 U7833 ( .A1(n6298), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6299) );
  MUX2_X1 U7834 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6299), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n6302) );
  INV_X1 U7835 ( .A(n6300), .ZN(n6301) );
  AND2_X1 U7836 ( .A1(n6302), .A2(n6301), .ZN(n6850) );
  AOI22_X1 U7837 ( .A1(n6850), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n8828), .ZN(n6303) );
  OAI21_X1 U7838 ( .B1(n6853), .B2(n8830), .A(n6303), .ZN(P2_U3353) );
  NOR2_X1 U7839 ( .A1(n6304), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9537) );
  INV_X2 U7840 ( .A(n9537), .ZN(n8242) );
  NAND2_X1 U7841 ( .A1(n6304), .A2(P1_U3084), .ZN(n9539) );
  OAI222_X1 U7842 ( .A1(n8242), .A2(n6306), .B1(n9539), .B2(n6305), .C1(n6527), 
        .C2(P1_U3084), .ZN(P1_U3351) );
  OAI222_X1 U7843 ( .A1(n8242), .A2(n6307), .B1(n9539), .B2(n6736), .C1(n6529), 
        .C2(P1_U3084), .ZN(P1_U3350) );
  OAI222_X1 U7844 ( .A1(n8242), .A2(n6308), .B1(n9539), .B2(n6748), .C1(
        P1_U3084), .C2(n9002), .ZN(P1_U3349) );
  OAI222_X1 U7845 ( .A1(n6512), .A2(P1_U3084), .B1(n9539), .B2(n6842), .C1(
        n6309), .C2(n8242), .ZN(P1_U3347) );
  OR2_X1 U7846 ( .A1(n6300), .A2(n8826), .ZN(n6310) );
  XNOR2_X1 U7847 ( .A(n6310), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9769) );
  INV_X1 U7848 ( .A(n9769), .ZN(n6311) );
  OAI222_X1 U7849 ( .A1(n8831), .A2(n10140), .B1(n8830), .B2(n6842), .C1(
        P2_U3152), .C2(n6311), .ZN(P2_U3352) );
  NAND2_X1 U7850 ( .A1(n6300), .A2(n6312), .ZN(n6318) );
  NAND2_X1 U7851 ( .A1(n6318), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6313) );
  XNOR2_X1 U7852 ( .A(n6313), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9782) );
  INV_X1 U7853 ( .A(n9782), .ZN(n6908) );
  OAI222_X1 U7854 ( .A1(n8831), .A2(n6909), .B1(n8830), .B2(n6906), .C1(
        P2_U3152), .C2(n6908), .ZN(P2_U3351) );
  INV_X1 U7855 ( .A(n9539), .ZN(n7498) );
  INV_X1 U7856 ( .A(n7498), .ZN(n8245) );
  OAI222_X1 U7857 ( .A1(n8242), .A2(n6315), .B1(n8245), .B2(n6314), .C1(n9655), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  OAI222_X1 U7858 ( .A1(n6558), .A2(P1_U3084), .B1(n8245), .B2(n6906), .C1(
        n6316), .C2(n8242), .ZN(P1_U3346) );
  OAI222_X1 U7859 ( .A1(n8242), .A2(n6317), .B1(n8245), .B2(n6853), .C1(n6595), 
        .C2(P1_U3084), .ZN(P1_U3348) );
  INV_X1 U7860 ( .A(n6334), .ZN(n6322) );
  NAND2_X1 U7861 ( .A1(n6319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6320) );
  MUX2_X1 U7862 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6320), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n6321) );
  INV_X1 U7863 ( .A(n6471), .ZN(n7010) );
  OAI222_X1 U7864 ( .A1(n8831), .A2(n7011), .B1(n8830), .B2(n7009), .C1(
        P2_U3152), .C2(n7010), .ZN(P2_U3350) );
  OAI222_X1 U7865 ( .A1(n6518), .A2(P1_U3084), .B1(n8245), .B2(n7009), .C1(
        n6323), .C2(n8242), .ZN(P1_U3345) );
  OR2_X1 U7866 ( .A1(n6334), .A2(n8826), .ZN(n6324) );
  XNOR2_X1 U7867 ( .A(n6324), .B(n6333), .ZN(n8454) );
  OAI222_X1 U7868 ( .A1(n8831), .A2(n7057), .B1(n8830), .B2(n7056), .C1(n8454), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U7869 ( .A1(P1_U3084), .A2(n6326), .B1(n9539), .B2(n7056), .C1(
        n6325), .C2(n8242), .ZN(P1_U3344) );
  INV_X1 U7870 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7871 ( .A1(n6986), .A2(P2_U3966), .ZN(n6327) );
  OAI21_X1 U7872 ( .B1(P2_U3966), .B2(n6328), .A(n6327), .ZN(P2_U3552) );
  INV_X1 U7873 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6332) );
  INV_X1 U7874 ( .A(n6330), .ZN(n6331) );
  AOI22_X1 U7875 ( .A1(n9666), .A2(n6332), .B1(n7140), .B2(n6331), .ZN(
        P1_U3441) );
  INV_X1 U7876 ( .A(n7076), .ZN(n6339) );
  NAND2_X1 U7877 ( .A1(n6334), .A2(n6333), .ZN(n6356) );
  NAND2_X1 U7878 ( .A1(n6356), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7879 ( .A1(n6336), .A2(n6335), .ZN(n6340) );
  OR2_X1 U7880 ( .A1(n6336), .A2(n6335), .ZN(n6337) );
  INV_X1 U7881 ( .A(n6488), .ZN(n7077) );
  OAI222_X1 U7882 ( .A1(n8831), .A2(n7078), .B1(n8830), .B2(n6339), .C1(n7077), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7883 ( .A(n6575), .ZN(n10164) );
  OAI222_X1 U7884 ( .A1(P1_U3084), .A2(n10164), .B1(n8245), .B2(n6339), .C1(
        n6338), .C2(n8242), .ZN(P1_U3343) );
  INV_X1 U7885 ( .A(n8484), .ZN(n9795) );
  NOR2_X1 U7886 ( .A1(n9795), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7887 ( .A(n7241), .ZN(n6343) );
  NAND2_X1 U7888 ( .A1(n6340), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6341) );
  XNOR2_X1 U7889 ( .A(n6341), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6450) );
  INV_X1 U7890 ( .A(n6450), .ZN(n7242) );
  OAI222_X1 U7891 ( .A1(n8831), .A2(n7243), .B1(n8830), .B2(n6343), .C1(n7242), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7892 ( .A(n6610), .ZN(n6604) );
  OAI222_X1 U7893 ( .A1(P1_U3084), .A2(n6604), .B1(n9539), .B2(n6343), .C1(
        n6342), .C2(n8242), .ZN(P1_U3342) );
  INV_X2 U7894 ( .A(n7875), .ZN(n7957) );
  NAND2_X1 U7895 ( .A1(n7957), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6346) );
  INV_X2 U7896 ( .A(n7912), .ZN(n7882) );
  NAND2_X1 U7897 ( .A1(n7882), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U7898 ( .A1(n7958), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6344) );
  AND3_X1 U7899 ( .A1(n6346), .A2(n6345), .A3(n6344), .ZN(n7978) );
  INV_X1 U7900 ( .A(n7978), .ZN(n8487) );
  NAND2_X1 U7901 ( .A1(n8487), .A2(P2_U3966), .ZN(n6347) );
  OAI21_X1 U7902 ( .B1(P2_U3966), .B2(n5068), .A(n6347), .ZN(P2_U3583) );
  INV_X1 U7903 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6355) );
  INV_X1 U7904 ( .A(n6348), .ZN(n6353) );
  OAI21_X1 U7905 ( .B1(n6350), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6349), .ZN(
        n6351) );
  XNOR2_X1 U7906 ( .A(n6351), .B(n9541), .ZN(n6352) );
  AOI22_X1 U7907 ( .A1(n6353), .A2(n6352), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3084), .ZN(n6354) );
  OAI21_X1 U7908 ( .B1(n10167), .B2(n6355), .A(n6354), .ZN(P1_U3241) );
  INV_X1 U7909 ( .A(n7454), .ZN(n6358) );
  NAND2_X1 U7910 ( .A1(n6380), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6357) );
  XNOR2_X1 U7911 ( .A(n6357), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6508) );
  INV_X1 U7912 ( .A(n6508), .ZN(n7455) );
  OAI222_X1 U7913 ( .A1(n8831), .A2(n10117), .B1(n8830), .B2(n6358), .C1(
        P2_U3152), .C2(n7455), .ZN(P2_U3346) );
  INV_X1 U7914 ( .A(n6709), .ZN(n6605) );
  OAI222_X1 U7915 ( .A1(n6605), .A2(P1_U3084), .B1(n8245), .B2(n6358), .C1(
        n10104), .C2(n8242), .ZN(P1_U3341) );
  NAND2_X1 U7916 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6773) );
  INV_X1 U7917 ( .A(n6773), .ZN(n6359) );
  NAND2_X1 U7918 ( .A1(n6359), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6833) );
  INV_X1 U7919 ( .A(n6833), .ZN(n6360) );
  NAND2_X1 U7920 ( .A1(n6360), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6864) );
  INV_X1 U7921 ( .A(n6864), .ZN(n6361) );
  NAND2_X1 U7922 ( .A1(n6361), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6915) );
  INV_X1 U7923 ( .A(n6915), .ZN(n6362) );
  NAND2_X1 U7924 ( .A1(n6362), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7017) );
  INV_X1 U7925 ( .A(n7017), .ZN(n6363) );
  NAND2_X1 U7926 ( .A1(n6363), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7083) );
  INV_X1 U7927 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7082) );
  INV_X1 U7928 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7247) );
  INV_X1 U7929 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7509) );
  INV_X1 U7930 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U7931 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n6368) );
  NAND2_X1 U7932 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n6370) );
  NAND2_X1 U7933 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n6372) );
  INV_X1 U7934 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9968) );
  INV_X1 U7935 ( .A(n7929), .ZN(n6374) );
  AND2_X1 U7936 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6373) );
  NAND2_X1 U7937 ( .A1(n6374), .A2(n6373), .ZN(n7931) );
  INV_X1 U7938 ( .A(n7931), .ZN(n7941) );
  INV_X1 U7939 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U7940 ( .A1(n7882), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U7941 ( .A1(n7957), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6375) );
  OAI211_X1 U7942 ( .C1(n7934), .C2(n6377), .A(n6376), .B(n6375), .ZN(n6378)
         );
  AOI21_X1 U7943 ( .B1(n7941), .B2(n7937), .A(n6378), .ZN(n8313) );
  NAND2_X1 U7944 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8448), .ZN(n6379) );
  OAI21_X1 U7945 ( .B1(n8313), .B2(n8448), .A(n6379), .ZN(P2_U3581) );
  INV_X1 U7946 ( .A(n7504), .ZN(n6382) );
  OAI21_X1 U7947 ( .B1(n6380), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6432) );
  XNOR2_X1 U7948 ( .A(n6432), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6663) );
  OAI222_X1 U7949 ( .A1(n8831), .A2(n9967), .B1(n8830), .B2(n6382), .C1(n7505), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7950 ( .A(n7120), .ZN(n7115) );
  OAI222_X1 U7951 ( .A1(P1_U3084), .A2(n7115), .B1(n9539), .B2(n6382), .C1(
        n6381), .C2(n8242), .ZN(P1_U3340) );
  INV_X1 U7952 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10119) );
  INV_X1 U7953 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9932) );
  MUX2_X1 U7954 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9932), .S(n6450), .Z(n6441)
         );
  INV_X1 U7955 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6383) );
  MUX2_X1 U7956 ( .A(n6383), .B(P2_REG1_REG_9__SCAN_IN), .S(n8454), .Z(n8458)
         );
  NAND2_X1 U7957 ( .A1(n6471), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6393) );
  INV_X1 U7958 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6384) );
  MUX2_X1 U7959 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6384), .S(n6471), .Z(n6466)
         );
  NAND2_X1 U7960 ( .A1(n9782), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6392) );
  INV_X1 U7961 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6385) );
  MUX2_X1 U7962 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6385), .S(n9782), .Z(n9787)
         );
  NAND2_X1 U7963 ( .A1(n9769), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6391) );
  INV_X1 U7964 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6386) );
  MUX2_X1 U7965 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6386), .S(n9769), .Z(n9771)
         );
  NAND2_X1 U7966 ( .A1(n6850), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6390) );
  INV_X1 U7967 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6387) );
  MUX2_X1 U7968 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6387), .S(n6850), .Z(n6478)
         );
  INV_X1 U7969 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6817) );
  MUX2_X1 U7970 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6817), .S(n9757), .Z(n9759)
         );
  NAND2_X1 U7971 ( .A1(n9742), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6389) );
  AOI21_X1 U7972 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n6410), .A(n6388), .ZN(
        n9748) );
  INV_X1 U7973 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9990) );
  MUX2_X1 U7974 ( .A(n9990), .B(P2_REG1_REG_3__SCAN_IN), .S(n9742), .Z(n9747)
         );
  OR2_X1 U7975 ( .A1(n9748), .A2(n9747), .ZN(n9750) );
  NAND2_X1 U7976 ( .A1(n6389), .A2(n9750), .ZN(n9760) );
  NAND2_X1 U7977 ( .A1(n9759), .A2(n9760), .ZN(n9758) );
  OAI21_X1 U7978 ( .B1(n6412), .B2(n6817), .A(n9758), .ZN(n6479) );
  NAND2_X1 U7979 ( .A1(n6478), .A2(n6479), .ZN(n6477) );
  NAND2_X1 U7980 ( .A1(n6390), .A2(n6477), .ZN(n9772) );
  NAND2_X1 U7981 ( .A1(n9771), .A2(n9772), .ZN(n9770) );
  NAND2_X1 U7982 ( .A1(n6391), .A2(n9770), .ZN(n9788) );
  NAND2_X1 U7983 ( .A1(n9787), .A2(n9788), .ZN(n9786) );
  NAND2_X1 U7984 ( .A1(n6392), .A2(n9786), .ZN(n6467) );
  NAND2_X1 U7985 ( .A1(n6466), .A2(n6467), .ZN(n6465) );
  NAND2_X1 U7986 ( .A1(n6393), .A2(n6465), .ZN(n8457) );
  NAND2_X1 U7987 ( .A1(n8458), .A2(n8457), .ZN(n8456) );
  OR2_X1 U7988 ( .A1(n8454), .A2(n6383), .ZN(n6489) );
  NAND2_X1 U7989 ( .A1(n8456), .A2(n6489), .ZN(n6396) );
  INV_X1 U7990 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6394) );
  MUX2_X1 U7991 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6394), .S(n6488), .Z(n6395)
         );
  NAND2_X1 U7992 ( .A1(n6396), .A2(n6395), .ZN(n6492) );
  NAND2_X1 U7993 ( .A1(n6488), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U7994 ( .A1(n6492), .A2(n6397), .ZN(n6442) );
  NAND2_X1 U7995 ( .A1(n6441), .A2(n6442), .ZN(n6440) );
  OAI21_X1 U7996 ( .B1(n9932), .B2(n7242), .A(n6440), .ZN(n6502) );
  AOI22_X1 U7997 ( .A1(n6508), .A2(n10119), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n7455), .ZN(n6501) );
  NOR2_X1 U7998 ( .A1(n6502), .A2(n6501), .ZN(n6500) );
  AOI21_X1 U7999 ( .B1(n7455), .B2(n10119), .A(n6500), .ZN(n6399) );
  INV_X1 U8000 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6659) );
  AOI22_X1 U8001 ( .A1(n6663), .A2(n6659), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7505), .ZN(n6398) );
  NOR2_X1 U8002 ( .A1(n6399), .A2(n6398), .ZN(n6658) );
  AOI21_X1 U8003 ( .B1(n6399), .B2(n6398), .A(n6658), .ZN(n6431) );
  NAND2_X1 U8004 ( .A1(n6508), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6421) );
  INV_X1 U8005 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6400) );
  MUX2_X1 U8006 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6400), .S(n6508), .Z(n6504)
         );
  NAND2_X1 U8007 ( .A1(n6488), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6418) );
  INV_X1 U8008 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6401) );
  MUX2_X1 U8009 ( .A(n6401), .B(P2_REG2_REG_10__SCAN_IN), .S(n6488), .Z(n6402)
         );
  INV_X1 U8010 ( .A(n6402), .ZN(n6496) );
  INV_X1 U8011 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8012 ( .A1(n6471), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6416) );
  INV_X1 U8013 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6403) );
  MUX2_X1 U8014 ( .A(n6403), .B(P2_REG2_REG_8__SCAN_IN), .S(n6471), .Z(n6404)
         );
  INV_X1 U8015 ( .A(n6404), .ZN(n6473) );
  NAND2_X1 U8016 ( .A1(n9782), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6415) );
  INV_X1 U8017 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6405) );
  MUX2_X1 U8018 ( .A(n6405), .B(P2_REG2_REG_7__SCAN_IN), .S(n9782), .Z(n6406)
         );
  INV_X1 U8019 ( .A(n6406), .ZN(n9784) );
  NAND2_X1 U8020 ( .A1(n9769), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6414) );
  INV_X1 U8021 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6407) );
  MUX2_X1 U8022 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6407), .S(n9769), .Z(n9774)
         );
  NAND2_X1 U8023 ( .A1(n6850), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6413) );
  INV_X1 U8024 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6408) );
  MUX2_X1 U8025 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6408), .S(n6850), .Z(n6484)
         );
  INV_X1 U8026 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7051) );
  MUX2_X1 U8027 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7051), .S(n9757), .Z(n9762)
         );
  NAND2_X1 U8028 ( .A1(n9742), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6411) );
  AOI21_X1 U8029 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n6410), .A(n6409), .ZN(
        n9744) );
  INV_X1 U8030 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9837) );
  MUX2_X1 U8031 ( .A(n9837), .B(P2_REG2_REG_3__SCAN_IN), .S(n9742), .Z(n9743)
         );
  OR2_X1 U8032 ( .A1(n9744), .A2(n9743), .ZN(n9746) );
  NAND2_X1 U8033 ( .A1(n6411), .A2(n9746), .ZN(n9763) );
  NAND2_X1 U8034 ( .A1(n9762), .A2(n9763), .ZN(n9761) );
  OAI21_X1 U8035 ( .B1(n6412), .B2(n7051), .A(n9761), .ZN(n6485) );
  NAND2_X1 U8036 ( .A1(n6484), .A2(n6485), .ZN(n6483) );
  NAND2_X1 U8037 ( .A1(n6413), .A2(n6483), .ZN(n9775) );
  NAND2_X1 U8038 ( .A1(n9774), .A2(n9775), .ZN(n9773) );
  NAND2_X1 U8039 ( .A1(n6414), .A2(n9773), .ZN(n9785) );
  NAND2_X1 U8040 ( .A1(n9784), .A2(n9785), .ZN(n9783) );
  NAND2_X1 U8041 ( .A1(n6415), .A2(n9783), .ZN(n6474) );
  NAND2_X1 U8042 ( .A1(n6473), .A2(n6474), .ZN(n6472) );
  NAND2_X1 U8043 ( .A1(n6416), .A2(n6472), .ZN(n8451) );
  MUX2_X1 U8044 ( .A(n6417), .B(P2_REG2_REG_9__SCAN_IN), .S(n8454), .Z(n8450)
         );
  NAND2_X1 U8045 ( .A1(n8451), .A2(n8450), .ZN(n8449) );
  OAI21_X1 U8046 ( .B1(n6417), .B2(n8454), .A(n8449), .ZN(n6497) );
  NAND2_X1 U8047 ( .A1(n6496), .A2(n6497), .ZN(n6495) );
  NAND2_X1 U8048 ( .A1(n6418), .A2(n6495), .ZN(n6446) );
  INV_X1 U8049 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6419) );
  AOI22_X1 U8050 ( .A1(n6450), .A2(n6419), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n7242), .ZN(n6445) );
  NOR2_X1 U8051 ( .A1(n6446), .A2(n6445), .ZN(n6444) );
  NOR2_X1 U8052 ( .A1(n6450), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6420) );
  NOR2_X1 U8053 ( .A1(n6444), .A2(n6420), .ZN(n6505) );
  NAND2_X1 U8054 ( .A1(n6504), .A2(n6505), .ZN(n6503) );
  NAND2_X1 U8055 ( .A1(n6421), .A2(n6503), .ZN(n6424) );
  INV_X1 U8056 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6422) );
  AOI22_X1 U8057 ( .A1(n6663), .A2(n6422), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7505), .ZN(n6423) );
  NOR2_X1 U8058 ( .A1(n6424), .A2(n6423), .ZN(n6664) );
  AOI21_X1 U8059 ( .B1(n6424), .B2(n6423), .A(n6664), .ZN(n6425) );
  NOR2_X1 U8060 ( .A1(n6425), .A2(n9736), .ZN(n6429) );
  INV_X1 U8061 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10135) );
  NOR2_X1 U8062 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10135), .ZN(n6426) );
  AOI21_X1 U8063 ( .B1(n9795), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n6426), .ZN(
        n6427) );
  OAI21_X1 U8064 ( .B1(n9734), .B2(n7505), .A(n6427), .ZN(n6428) );
  NOR2_X1 U8065 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  OAI21_X1 U8066 ( .B1(n6431), .B2(n8475), .A(n6430), .ZN(P2_U3258) );
  INV_X1 U8067 ( .A(n7625), .ZN(n6439) );
  INV_X1 U8068 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U8069 ( .A1(n6432), .A2(n10133), .ZN(n6433) );
  NAND2_X1 U8070 ( .A1(n6433), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U8071 ( .A1(n6435), .A2(n6434), .ZN(n6618) );
  OR2_X1 U8072 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  INV_X1 U8073 ( .A(n7626), .ZN(n6787) );
  OAI222_X1 U8074 ( .A1(n8831), .A2(n6437), .B1(n8830), .B2(n6439), .C1(n6787), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8075 ( .A(n7124), .ZN(n7415) );
  OAI222_X1 U8076 ( .A1(P1_U3084), .A2(n7415), .B1(n9539), .B2(n6439), .C1(
        n6438), .C2(n8242), .ZN(P1_U3339) );
  INV_X1 U8077 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10125) );
  OAI211_X1 U8078 ( .C1(n6442), .C2(n6441), .A(n9804), .B(n6440), .ZN(n6443)
         );
  NAND2_X1 U8079 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7254) );
  OAI211_X1 U8080 ( .C1(n8484), .C2(n10125), .A(n6443), .B(n7254), .ZN(n6449)
         );
  AOI21_X1 U8081 ( .B1(n6446), .B2(n6445), .A(n6444), .ZN(n6447) );
  NOR2_X1 U8082 ( .A1(n6447), .A2(n9736), .ZN(n6448) );
  AOI211_X1 U8083 ( .C1(n9802), .C2(n6450), .A(n6449), .B(n6448), .ZN(n6451)
         );
  INV_X1 U8084 ( .A(n6451), .ZN(P2_U3256) );
  INV_X1 U8085 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6452) );
  INV_X1 U8086 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6993) );
  OAI22_X1 U8087 ( .A1(n8484), .A2(n6452), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6993), .ZN(n6458) );
  OAI211_X1 U8088 ( .C1(n6455), .C2(n6454), .A(n9804), .B(n6453), .ZN(n6456)
         );
  INV_X1 U8089 ( .A(n6456), .ZN(n6457) );
  AOI211_X1 U8090 ( .C1(n9802), .C2(n6459), .A(n6458), .B(n6457), .ZN(n6464)
         );
  OAI211_X1 U8091 ( .C1(n6462), .C2(n6461), .A(n9797), .B(n6460), .ZN(n6463)
         );
  NAND2_X1 U8092 ( .A1(n6464), .A2(n6463), .ZN(P2_U3246) );
  INV_X1 U8093 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6469) );
  OAI211_X1 U8094 ( .C1(n6467), .C2(n6466), .A(n9804), .B(n6465), .ZN(n6468)
         );
  NAND2_X1 U8095 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7015) );
  OAI211_X1 U8096 ( .C1(n8484), .C2(n6469), .A(n6468), .B(n7015), .ZN(n6470)
         );
  AOI21_X1 U8097 ( .B1(n6471), .B2(n9802), .A(n6470), .ZN(n6476) );
  OAI211_X1 U8098 ( .C1(n6474), .C2(n6473), .A(n9797), .B(n6472), .ZN(n6475)
         );
  NAND2_X1 U8099 ( .A1(n6476), .A2(n6475), .ZN(P2_U3253) );
  INV_X1 U8100 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6481) );
  OAI211_X1 U8101 ( .C1(n6479), .C2(n6478), .A(n9804), .B(n6477), .ZN(n6480)
         );
  NAND2_X1 U8102 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n6888) );
  OAI211_X1 U8103 ( .C1(n8484), .C2(n6481), .A(n6480), .B(n6888), .ZN(n6482)
         );
  AOI21_X1 U8104 ( .B1(n6850), .B2(n9802), .A(n6482), .ZN(n6487) );
  OAI211_X1 U8105 ( .C1(n6485), .C2(n6484), .A(n9797), .B(n6483), .ZN(n6486)
         );
  NAND2_X1 U8106 ( .A1(n6487), .A2(n6486), .ZN(P2_U3250) );
  NAND2_X1 U8107 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7096) );
  INV_X1 U8108 ( .A(n7096), .ZN(n6494) );
  MUX2_X1 U8109 ( .A(n6394), .B(P2_REG1_REG_10__SCAN_IN), .S(n6488), .Z(n6490)
         );
  NAND3_X1 U8110 ( .A1(n6490), .A2(n8456), .A3(n6489), .ZN(n6491) );
  AND3_X1 U8111 ( .A1(n9804), .A2(n6492), .A3(n6491), .ZN(n6493) );
  AOI211_X1 U8112 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9795), .A(n6494), .B(
        n6493), .ZN(n6499) );
  OAI211_X1 U8113 ( .C1(n6497), .C2(n6496), .A(n9797), .B(n6495), .ZN(n6498)
         );
  OAI211_X1 U8114 ( .C1(n9734), .C2(n7077), .A(n6499), .B(n6498), .ZN(P2_U3255) );
  AOI21_X1 U8115 ( .B1(n6502), .B2(n6501), .A(n6500), .ZN(n6511) );
  OAI211_X1 U8116 ( .C1(n6505), .C2(n6504), .A(n9797), .B(n6503), .ZN(n6510)
         );
  INV_X1 U8117 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8118 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7482) );
  OAI21_X1 U8119 ( .B1(n8484), .B2(n6506), .A(n7482), .ZN(n6507) );
  AOI21_X1 U8120 ( .B1(n9802), .B2(n6508), .A(n6507), .ZN(n6509) );
  OAI211_X1 U8121 ( .C1(n6511), .C2(n8475), .A(n6510), .B(n6509), .ZN(P2_U3257) );
  NOR2_X1 U8122 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6533), .ZN(n6517) );
  NOR2_X1 U8123 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n6630), .ZN(n6515) );
  AOI22_X1 U8124 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n6512), .B1(n6630), .B2(
        n5391), .ZN(n6624) );
  INV_X1 U8125 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10108) );
  INV_X1 U8126 ( .A(n6529), .ZN(n8994) );
  INV_X1 U8127 ( .A(n6527), .ZN(n6513) );
  NAND2_X1 U8128 ( .A1(n6513), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8988) );
  MUX2_X1 U8129 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n5436), .S(n6529), .Z(n8990)
         );
  AOI21_X1 U8130 ( .B1(n8994), .B2(P1_REG1_REG_3__SCAN_IN), .A(n8992), .ZN(
        n9005) );
  MUX2_X1 U8131 ( .A(n10108), .B(P1_REG1_REG_4__SCAN_IN), .S(n9002), .Z(n9004)
         );
  NAND2_X1 U8132 ( .A1(n9005), .A2(n9004), .ZN(n9003) );
  MUX2_X1 U8133 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6589), .S(n6595), .Z(n6514)
         );
  OAI21_X1 U8134 ( .B1(n6589), .B2(n6595), .A(n6590), .ZN(n6625) );
  NOR2_X1 U8135 ( .A1(n6624), .A2(n6625), .ZN(n6623) );
  MUX2_X1 U8136 ( .A(n6516), .B(P1_REG1_REG_7__SCAN_IN), .S(n6533), .Z(n6555)
         );
  NOR2_X1 U8137 ( .A1(n6556), .A2(n6555), .ZN(n6554) );
  NOR2_X1 U8138 ( .A1(n6517), .A2(n6554), .ZN(n6520) );
  AOI22_X1 U8139 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6518), .B1(n6573), .B2(
        n5305), .ZN(n6519) );
  NOR2_X1 U8140 ( .A1(n6520), .A2(n6519), .ZN(n6563) );
  AOI21_X1 U8141 ( .B1(n6520), .B2(n6519), .A(n6563), .ZN(n6539) );
  INV_X1 U8142 ( .A(n10163), .ZN(n9036) );
  INV_X1 U8143 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U8144 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7314) );
  OAI21_X1 U8145 ( .B1(n10167), .B2(n6521), .A(n7314), .ZN(n6522) );
  AOI21_X1 U8146 ( .B1(n6573), .B2(n9036), .A(n6522), .ZN(n6538) );
  INV_X1 U8147 ( .A(n10154), .ZN(n9651) );
  NOR2_X1 U8148 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6573), .ZN(n6523) );
  AOI21_X1 U8149 ( .B1(n6573), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6523), .ZN(
        n6535) );
  NOR2_X1 U8150 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6533), .ZN(n6524) );
  AOI21_X1 U8151 ( .B1(n6533), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6524), .ZN(
        n6552) );
  OAI21_X1 U8152 ( .B1(n6527), .B2(n6526), .A(n6525), .ZN(n8997) );
  XNOR2_X1 U8153 ( .A(n6529), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U8154 ( .A1(n8997), .A2(n8998), .ZN(n8996) );
  OAI21_X1 U8155 ( .B1(n6529), .B2(n6528), .A(n8996), .ZN(n9009) );
  MUX2_X1 U8156 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7529), .S(n9002), .Z(n9010)
         );
  NOR2_X1 U8157 ( .A1(n9009), .A2(n9010), .ZN(n9008) );
  AOI21_X1 U8158 ( .B1(n9002), .B2(n7529), .A(n9008), .ZN(n6585) );
  XNOR2_X1 U8159 ( .A(n6595), .B(n6530), .ZN(n6584) );
  INV_X1 U8160 ( .A(n6595), .ZN(n6531) );
  OAI22_X1 U8161 ( .A1(n6585), .A2(n6584), .B1(n6531), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U8162 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n6630), .ZN(n6532) );
  OAI21_X1 U8163 ( .B1(n6630), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6532), .ZN(
        n6628) );
  NOR2_X1 U8164 ( .A1(n6627), .A2(n6628), .ZN(n6626) );
  AOI21_X1 U8165 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6630), .A(n6626), .ZN(
        n6553) );
  NAND2_X1 U8166 ( .A1(n6552), .A2(n6553), .ZN(n6551) );
  OAI21_X1 U8167 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6533), .A(n6551), .ZN(
        n6534) );
  NAND2_X1 U8168 ( .A1(n6535), .A2(n6534), .ZN(n6572) );
  OAI21_X1 U8169 ( .B1(n6535), .B2(n6534), .A(n6572), .ZN(n6536) );
  NAND2_X1 U8170 ( .A1(n9651), .A2(n6536), .ZN(n6537) );
  OAI211_X1 U8171 ( .C1(n6539), .C2(n10162), .A(n6538), .B(n6537), .ZN(
        P1_U3249) );
  NAND2_X1 U8172 ( .A1(n7128), .A2(n7985), .ZN(n6540) );
  OR2_X1 U8173 ( .A1(n6234), .A2(n6540), .ZN(n9905) );
  INV_X1 U8174 ( .A(n9877), .ZN(n9919) );
  OAI22_X1 U8175 ( .A1(n6541), .A2(n9915), .B1(n6797), .B2(n9914), .ZN(n6543)
         );
  AOI211_X1 U8176 ( .C1(n9919), .C2(n6544), .A(n6543), .B(n6542), .ZN(n6600)
         );
  NAND2_X1 U8177 ( .A1(n9921), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6547) );
  OAI21_X1 U8178 ( .B1(n6600), .B2(n9921), .A(n6547), .ZN(P2_U3457) );
  INV_X1 U8179 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U8180 ( .A1(n6548), .A2(n8986), .ZN(n6549) );
  OAI21_X1 U8181 ( .B1(n8986), .B2(n6550), .A(n6549), .ZN(P1_U3586) );
  OAI21_X1 U8182 ( .B1(n6553), .B2(n6552), .A(n6551), .ZN(n6561) );
  INV_X1 U8183 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U8184 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7300) );
  OAI21_X1 U8185 ( .B1(n10167), .B2(n10077), .A(n7300), .ZN(n6560) );
  AOI21_X1 U8186 ( .B1(n6556), .B2(n6555), .A(n6554), .ZN(n6557) );
  OAI22_X1 U8187 ( .A1(n6558), .A2(n10163), .B1(n10162), .B2(n6557), .ZN(n6559) );
  AOI211_X1 U8188 ( .C1(n9651), .C2(n6561), .A(n6560), .B(n6559), .ZN(n6562)
         );
  INV_X1 U8189 ( .A(n6562), .ZN(P1_U3248) );
  OR2_X1 U8190 ( .A1(n6642), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6567) );
  NOR2_X1 U8191 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6573), .ZN(n6564) );
  MUX2_X1 U8192 ( .A(n6565), .B(P1_REG1_REG_9__SCAN_IN), .S(n6642), .Z(n6635)
         );
  NOR2_X1 U8193 ( .A1(n6636), .A2(n6635), .ZN(n6634) );
  INV_X1 U8194 ( .A(n6634), .ZN(n6566) );
  MUX2_X1 U8195 ( .A(n6568), .B(P1_REG1_REG_10__SCAN_IN), .S(n6575), .Z(n10160) );
  NOR2_X1 U8196 ( .A1(n10159), .A2(n10160), .ZN(n10158) );
  AOI22_X1 U8197 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6604), .B1(n6610), .B2(
        n5257), .ZN(n6569) );
  NOR2_X1 U8198 ( .A1(n6570), .A2(n6569), .ZN(n6603) );
  AOI21_X1 U8199 ( .B1(n6570), .B2(n6569), .A(n6603), .ZN(n6583) );
  AOI22_X1 U8200 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6610), .B1(n6604), .B2(
        n5261), .ZN(n6577) );
  NAND2_X1 U8201 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6642), .ZN(n6571) );
  OAI21_X1 U8202 ( .B1(n6642), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6571), .ZN(
        n6638) );
  OAI21_X1 U8203 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6573), .A(n6572), .ZN(
        n6639) );
  NOR2_X1 U8204 ( .A1(n6638), .A2(n6639), .ZN(n6637) );
  AOI21_X1 U8205 ( .B1(n6642), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6637), .ZN(
        n10157) );
  NAND2_X1 U8206 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6575), .ZN(n6574) );
  OAI21_X1 U8207 ( .B1(n6575), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6574), .ZN(
        n10156) );
  NOR2_X1 U8208 ( .A1(n10157), .A2(n10156), .ZN(n10155) );
  AOI21_X1 U8209 ( .B1(n6575), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10155), .ZN(
        n6576) );
  NAND2_X1 U8210 ( .A1(n6577), .A2(n6576), .ZN(n6609) );
  OAI21_X1 U8211 ( .B1(n6577), .B2(n6576), .A(n6609), .ZN(n6581) );
  INV_X1 U8212 ( .A(n10167), .ZN(n9658) );
  AOI21_X1 U8213 ( .B1(n9658), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n6578), .ZN(
        n6579) );
  OAI21_X1 U8214 ( .B1(n6604), .B2(n10163), .A(n6579), .ZN(n6580) );
  AOI21_X1 U8215 ( .B1(n6581), .B2(n9651), .A(n6580), .ZN(n6582) );
  OAI21_X1 U8216 ( .B1(n6583), .B2(n10162), .A(n6582), .ZN(P1_U3252) );
  XNOR2_X1 U8217 ( .A(n6585), .B(n6584), .ZN(n6588) );
  NOR2_X1 U8218 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10094), .ZN(n7325) );
  INV_X1 U8219 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6586) );
  NOR2_X1 U8220 ( .A1(n10167), .A2(n6586), .ZN(n6587) );
  AOI211_X1 U8221 ( .C1(n9651), .C2(n6588), .A(n7325), .B(n6587), .ZN(n6594)
         );
  MUX2_X1 U8222 ( .A(n6589), .B(P1_REG1_REG_5__SCAN_IN), .S(n6595), .Z(n6591)
         );
  INV_X1 U8223 ( .A(n10162), .ZN(n9660) );
  OAI211_X1 U8224 ( .C1(n6592), .C2(n6591), .A(n9660), .B(n6590), .ZN(n6593)
         );
  OAI211_X1 U8225 ( .C1(n10163), .C2(n6595), .A(n6594), .B(n6593), .ZN(
        P1_U3246) );
  INV_X1 U8226 ( .A(n6755), .ZN(n6598) );
  NAND4_X1 U8227 ( .A1(n6598), .A2(n6597), .A3(n6763), .A4(n6596), .ZN(n6599)
         );
  OR2_X1 U8228 ( .A1(n6600), .A2(n9931), .ZN(n6601) );
  OAI21_X1 U8229 ( .B1(n9934), .B2(n6602), .A(n6601), .ZN(P2_U3522) );
  AOI21_X1 U8230 ( .B1(n5257), .B2(n6604), .A(n6603), .ZN(n6607) );
  AOI22_X1 U8231 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6605), .B1(n6709), .B2(
        n5243), .ZN(n6606) );
  NOR2_X1 U8232 ( .A1(n6607), .A2(n6606), .ZN(n6703) );
  AOI21_X1 U8233 ( .B1(n6607), .B2(n6606), .A(n6703), .ZN(n6617) );
  INV_X1 U8234 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U8235 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7774) );
  OAI21_X1 U8236 ( .B1(n10167), .B2(n6608), .A(n7774), .ZN(n6615) );
  OAI21_X1 U8237 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6610), .A(n6609), .ZN(
        n6613) );
  NAND2_X1 U8238 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6709), .ZN(n6611) );
  OAI21_X1 U8239 ( .B1(n6709), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6611), .ZN(
        n6612) );
  NOR2_X1 U8240 ( .A1(n6613), .A2(n6612), .ZN(n6708) );
  AOI211_X1 U8241 ( .C1(n6613), .C2(n6612), .A(n6708), .B(n10154), .ZN(n6614)
         );
  AOI211_X1 U8242 ( .C1(n9036), .C2(n6709), .A(n6615), .B(n6614), .ZN(n6616)
         );
  OAI21_X1 U8243 ( .B1(n6617), .B2(n10162), .A(n6616), .ZN(P1_U3253) );
  INV_X1 U8244 ( .A(n7640), .ZN(n6622) );
  NAND2_X1 U8245 ( .A1(n6618), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6619) );
  XNOR2_X1 U8246 ( .A(n6619), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7642) );
  INV_X1 U8247 ( .A(n7642), .ZN(n6791) );
  OAI222_X1 U8248 ( .A1(n8831), .A2(n6620), .B1(n8830), .B2(n6622), .C1(
        P2_U3152), .C2(n6791), .ZN(P2_U3343) );
  OAI222_X1 U8249 ( .A1(n7587), .A2(P1_U3084), .B1(n8245), .B2(n6622), .C1(
        n6621), .C2(n8242), .ZN(P1_U3338) );
  AOI21_X1 U8250 ( .B1(n6625), .B2(n6624), .A(n6623), .ZN(n6633) );
  AND2_X1 U8251 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9632) );
  AOI211_X1 U8252 ( .C1(n6628), .C2(n6627), .A(n6626), .B(n10154), .ZN(n6629)
         );
  AOI211_X1 U8253 ( .C1(n9658), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9632), .B(
        n6629), .ZN(n6632) );
  NAND2_X1 U8254 ( .A1(n9036), .A2(n6630), .ZN(n6631) );
  OAI211_X1 U8255 ( .C1(n6633), .C2(n10162), .A(n6632), .B(n6631), .ZN(
        P1_U3247) );
  AOI21_X1 U8256 ( .B1(n6636), .B2(n6635), .A(n6634), .ZN(n6645) );
  AOI211_X1 U8257 ( .C1(n6639), .C2(n6638), .A(n6637), .B(n10154), .ZN(n6640)
         );
  AOI211_X1 U8258 ( .C1(n9658), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n6641), .B(
        n6640), .ZN(n6644) );
  NAND2_X1 U8259 ( .A1(n9036), .A2(n6642), .ZN(n6643) );
  OAI211_X1 U8260 ( .C1(n6645), .C2(n10162), .A(n6644), .B(n6643), .ZN(
        P1_U3250) );
  INV_X1 U8261 ( .A(n7801), .ZN(n6648) );
  NAND2_X1 U8262 ( .A1(n6646), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6647) );
  XNOR2_X1 U8263 ( .A(n6647), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7543) );
  INV_X1 U8264 ( .A(n7543), .ZN(n7802) );
  OAI222_X1 U8265 ( .A1(n8831), .A2(n7803), .B1(n8830), .B2(n6648), .C1(n7802), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  OAI222_X1 U8266 ( .A1(n8242), .A2(n6649), .B1(n9539), .B2(n6648), .C1(
        P1_U3084), .C2(n9023), .ZN(P1_U3337) );
  INV_X1 U8267 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6656) );
  NOR3_X1 U8268 ( .A1(n6652), .A2(n6651), .A3(n6650), .ZN(n6653) );
  AOI21_X1 U8269 ( .B1(n9306), .B2(n5823), .A(n6653), .ZN(n7147) );
  OAI21_X1 U8270 ( .B1(n4531), .B2(n6654), .A(n7147), .ZN(n9513) );
  NAND2_X1 U8271 ( .A1(n9513), .A2(n9724), .ZN(n6655) );
  OAI21_X1 U8272 ( .B1(n9724), .B2(n6656), .A(n6655), .ZN(P1_U3454) );
  INV_X1 U8273 ( .A(n7808), .ZN(n6719) );
  AOI22_X1 U8274 ( .A1(n9031), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9537), .ZN(n6657) );
  OAI21_X1 U8275 ( .B1(n6719), .B2(n8245), .A(n6657), .ZN(P1_U3336) );
  AOI21_X1 U8276 ( .B1(n7505), .B2(n6659), .A(n6658), .ZN(n6661) );
  INV_X1 U8277 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10138) );
  AOI22_X1 U8278 ( .A1(n7626), .A2(n10138), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n6787), .ZN(n6660) );
  NOR2_X1 U8279 ( .A1(n6661), .A2(n6660), .ZN(n6786) );
  AOI21_X1 U8280 ( .B1(n6661), .B2(n6660), .A(n6786), .ZN(n6673) );
  INV_X1 U8281 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U8282 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7698) );
  OAI21_X1 U8283 ( .B1(n8484), .B2(n6662), .A(n7698), .ZN(n6671) );
  NOR2_X1 U8284 ( .A1(n6663), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6665) );
  NOR2_X1 U8285 ( .A1(n6665), .A2(n6664), .ZN(n6668) );
  INV_X1 U8286 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6666) );
  AOI22_X1 U8287 ( .A1(n7626), .A2(n6666), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n6787), .ZN(n6667) );
  NOR2_X1 U8288 ( .A1(n6668), .A2(n6667), .ZN(n6783) );
  AOI21_X1 U8289 ( .B1(n6668), .B2(n6667), .A(n6783), .ZN(n6669) );
  NOR2_X1 U8290 ( .A1(n6669), .A2(n9736), .ZN(n6670) );
  AOI211_X1 U8291 ( .C1(n9802), .C2(n7626), .A(n6671), .B(n6670), .ZN(n6672)
         );
  OAI21_X1 U8292 ( .B1(n6673), .B2(n8475), .A(n6672), .ZN(P2_U3259) );
  XNOR2_X1 U8293 ( .A(n6676), .B(n6675), .ZN(n6677) );
  XNOR2_X1 U8294 ( .A(n6674), .B(n6677), .ZN(n6681) );
  INV_X1 U8295 ( .A(n8964), .ZN(n6698) );
  NAND2_X1 U8296 ( .A1(n5357), .A2(n9712), .ZN(n6694) );
  INV_X1 U8297 ( .A(n6694), .ZN(n6678) );
  AOI22_X1 U8298 ( .A1(n6698), .A2(n5838), .B1(n6678), .B2(n9642), .ZN(n6680)
         );
  INV_X1 U8299 ( .A(n7301), .ZN(n8967) );
  NAND2_X1 U8300 ( .A1(n9642), .A2(n7139), .ZN(n6823) );
  AOI22_X1 U8301 ( .A1(n8967), .A2(n8987), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6823), .ZN(n6679) );
  OAI211_X1 U8302 ( .C1(n6681), .C2(n8972), .A(n6680), .B(n6679), .ZN(P1_U3220) );
  NAND2_X1 U8303 ( .A1(n6682), .A2(n6683), .ZN(n7149) );
  OAI21_X1 U8304 ( .B1(n6682), .B2(n6683), .A(n7149), .ZN(n8229) );
  AND2_X1 U8305 ( .A1(n6684), .A2(n9274), .ZN(n6685) );
  NAND2_X1 U8306 ( .A1(n7346), .A2(n6685), .ZN(n9497) );
  AOI22_X1 U8307 ( .A1(n9306), .A2(n5838), .B1(n9304), .B2(n8987), .ZN(n6693)
         );
  XNOR2_X1 U8308 ( .A(n6682), .B(n6686), .ZN(n6691) );
  NAND2_X1 U8309 ( .A1(n6687), .A2(n9061), .ZN(n6690) );
  NAND2_X1 U8310 ( .A1(n5800), .A2(n6688), .ZN(n6689) );
  NAND2_X1 U8311 ( .A1(n6691), .A2(n9501), .ZN(n6692) );
  OAI211_X1 U8312 ( .C1(n8229), .C2(n9497), .A(n6693), .B(n6692), .ZN(n8233)
         );
  NAND2_X1 U8313 ( .A1(n5804), .A2(n7152), .ZN(n9718) );
  OAI211_X1 U8314 ( .C1(n4531), .C2(n8236), .A(n9713), .B(n7172), .ZN(n8231)
         );
  OAI211_X1 U8315 ( .C1(n8229), .C2(n9718), .A(n6694), .B(n8231), .ZN(n6695)
         );
  NOR2_X1 U8316 ( .A1(n8233), .A2(n6695), .ZN(n9668) );
  NAND2_X1 U8317 ( .A1(n9731), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6697) );
  OAI21_X1 U8318 ( .B1(n9668), .B2(n9731), .A(n6697), .ZN(P1_U3524) );
  AOI22_X1 U8319 ( .A1(n6698), .A2(n5823), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6823), .ZN(n6701) );
  NAND2_X1 U8320 ( .A1(n6699), .A2(n9643), .ZN(n6700) );
  OAI211_X1 U8321 ( .C1(n8959), .C2(n4531), .A(n6701), .B(n6700), .ZN(P1_U3230) );
  NOR2_X1 U8322 ( .A1(n6709), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6702) );
  MUX2_X1 U8323 ( .A(n6704), .B(P1_REG1_REG_13__SCAN_IN), .S(n7120), .Z(n6705)
         );
  NOR2_X1 U8324 ( .A1(n6706), .A2(n6705), .ZN(n7114) );
  AOI21_X1 U8325 ( .B1(n6706), .B2(n6705), .A(n7114), .ZN(n6716) );
  AND2_X1 U8326 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6707) );
  AOI21_X1 U8327 ( .B1(n9658), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n6707), .ZN(
        n6715) );
  AOI21_X1 U8328 ( .B1(n6709), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6708), .ZN(
        n6712) );
  NAND2_X1 U8329 ( .A1(n7120), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6710) );
  OAI21_X1 U8330 ( .B1(n7120), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6710), .ZN(
        n6711) );
  NOR2_X1 U8331 ( .A1(n6712), .A2(n6711), .ZN(n7119) );
  AOI211_X1 U8332 ( .C1(n6712), .C2(n6711), .A(n7119), .B(n10154), .ZN(n6713)
         );
  AOI21_X1 U8333 ( .B1(n9036), .B2(n7120), .A(n6713), .ZN(n6714) );
  OAI211_X1 U8334 ( .C1(n6716), .C2(n10162), .A(n6715), .B(n6714), .ZN(
        P1_U3254) );
  NAND2_X1 U8335 ( .A1(n6095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6717) );
  MUX2_X1 U8336 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6717), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6718) );
  NAND2_X1 U8337 ( .A1(n6718), .A2(n6978), .ZN(n9800) );
  OAI222_X1 U8338 ( .A1(n8831), .A2(n7809), .B1(n8830), .B2(n6719), .C1(n9800), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND3_X1 U8339 ( .A1(n8171), .A2(n6722), .A3(n7260), .ZN(n6721) );
  XNOR2_X1 U8340 ( .A(n4321), .B(n6998), .ZN(n6725) );
  INV_X1 U8341 ( .A(n6722), .ZN(n6723) );
  AND2_X2 U8342 ( .A1(n6723), .A2(n8178), .ZN(n8306) );
  NAND2_X1 U8343 ( .A1(n6206), .A2(n8301), .ZN(n6724) );
  NAND2_X1 U8344 ( .A1(n6727), .A2(n6726), .ZN(n6897) );
  OAI22_X1 U8345 ( .A1(n6997), .A2(n8306), .B1(n6990), .B2(n4322), .ZN(n6896)
         );
  AND2_X1 U8346 ( .A1(n9820), .A2(n8301), .ZN(n6728) );
  XNOR2_X1 U8347 ( .A(n6876), .B(n4322), .ZN(n6729) );
  NAND2_X1 U8348 ( .A1(n6728), .A2(n6729), .ZN(n6732) );
  INV_X1 U8349 ( .A(n6728), .ZN(n6731) );
  INV_X1 U8350 ( .A(n6729), .ZN(n6730) );
  NAND2_X1 U8351 ( .A1(n6731), .A2(n6730), .ZN(n6733) );
  AND2_X1 U8352 ( .A1(n6732), .A2(n6733), .ZN(n6879) );
  NAND2_X1 U8353 ( .A1(n6771), .A2(n8301), .ZN(n6737) );
  NAND2_X1 U8354 ( .A1(n6839), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U8355 ( .A1(n7641), .A2(n9742), .ZN(n6734) );
  NAND2_X1 U8356 ( .A1(n6738), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6745) );
  NAND2_X1 U8357 ( .A1(n4341), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6744) );
  INV_X1 U8358 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6739) );
  NAND2_X1 U8359 ( .A1(n9833), .A2(n6739), .ZN(n6740) );
  AND2_X1 U8360 ( .A1(n6740), .A2(n6773), .ZN(n7046) );
  NAND2_X1 U8361 ( .A1(n6741), .A2(n7046), .ZN(n6743) );
  NAND2_X1 U8362 ( .A1(n7958), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6742) );
  NAND4_X1 U8363 ( .A1(n6745), .A2(n6744), .A3(n6743), .A4(n6742), .ZN(n9819)
         );
  NAND2_X1 U8364 ( .A1(n9819), .A2(n8301), .ZN(n6750) );
  NAND2_X1 U8365 ( .A1(n7970), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6747) );
  NAND2_X1 U8366 ( .A1(n7641), .A2(n9757), .ZN(n6746) );
  XNOR2_X1 U8367 ( .A(n7048), .B(n8300), .ZN(n6749) );
  NAND2_X1 U8368 ( .A1(n6750), .A2(n6749), .ZN(n6848) );
  OAI21_X1 U8369 ( .B1(n6750), .B2(n6749), .A(n6848), .ZN(n6753) );
  OR2_X1 U8370 ( .A1(n6751), .A2(n6753), .ZN(n6849) );
  INV_X1 U8371 ( .A(n6849), .ZN(n6752) );
  AOI21_X1 U8372 ( .B1(n6751), .B2(n6753), .A(n6752), .ZN(n6782) );
  OR2_X1 U8373 ( .A1(n6755), .A2(n6754), .ZN(n6756) );
  INV_X1 U8374 ( .A(n9840), .ZN(n8180) );
  NAND2_X1 U8375 ( .A1(n9914), .A2(n6758), .ZN(n6759) );
  INV_X1 U8376 ( .A(n6760), .ZN(n6761) );
  NAND2_X1 U8377 ( .A1(n6761), .A2(n8172), .ZN(n6765) );
  NAND2_X1 U8378 ( .A1(n6761), .A2(n9914), .ZN(n6764) );
  NAND4_X1 U8379 ( .A1(n6765), .A2(n6764), .A3(n6763), .A4(n6762), .ZN(n6766)
         );
  OR2_X1 U8380 ( .A1(n6768), .A2(n6767), .ZN(n6769) );
  INV_X1 U8381 ( .A(n8421), .ZN(n8436) );
  AND2_X1 U8382 ( .A1(n6770), .A2(n8178), .ZN(n8407) );
  INV_X1 U8383 ( .A(n6771), .ZN(n6796) );
  INV_X1 U8384 ( .A(n9821), .ZN(n8664) );
  NAND2_X1 U8385 ( .A1(n7882), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8386 ( .A1(n7958), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6777) );
  INV_X1 U8387 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U8388 ( .A1(n6773), .A2(n6772), .ZN(n6774) );
  AND2_X1 U8389 ( .A1(n6833), .A2(n6774), .ZN(n6887) );
  NAND2_X1 U8390 ( .A1(n7937), .A2(n6887), .ZN(n6776) );
  NAND2_X1 U8391 ( .A1(n7957), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6775) );
  NAND4_X1 U8392 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n8447)
         );
  INV_X1 U8393 ( .A(n8447), .ZN(n6936) );
  INV_X1 U8394 ( .A(n9818), .ZN(n8662) );
  OAI22_X1 U8395 ( .A1(n6796), .A2(n8664), .B1(n6936), .B2(n8662), .ZN(n6807)
         );
  NAND2_X1 U8396 ( .A1(n8407), .A2(n6807), .ZN(n6779) );
  NAND2_X1 U8397 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9755) );
  OAI211_X1 U8398 ( .C1(n8436), .C2(n6933), .A(n6779), .B(n9755), .ZN(n6780)
         );
  AOI21_X1 U8399 ( .B1(n7046), .B2(n8433), .A(n6780), .ZN(n6781) );
  OAI21_X1 U8400 ( .B1(n6782), .B2(n8423), .A(n6781), .ZN(P2_U3232) );
  NOR2_X1 U8401 ( .A1(n7626), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6784) );
  NOR2_X1 U8402 ( .A1(n6784), .A2(n6783), .ZN(n6968) );
  XNOR2_X1 U8403 ( .A(n7642), .B(n6968), .ZN(n6785) );
  NOR2_X1 U8404 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n6785), .ZN(n6969) );
  AOI21_X1 U8405 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n6785), .A(n6969), .ZN(
        n6795) );
  AOI21_X1 U8406 ( .B1(n6787), .B2(n10138), .A(n6786), .ZN(n6961) );
  XOR2_X1 U8407 ( .A(n7642), .B(n6961), .Z(n6788) );
  NAND2_X1 U8408 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n6788), .ZN(n6962) );
  OAI211_X1 U8409 ( .C1(n6788), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9804), .B(
        n6962), .ZN(n6794) );
  AND2_X1 U8410 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6789) );
  AOI21_X1 U8411 ( .B1(n9795), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n6789), .ZN(
        n6790) );
  OAI21_X1 U8412 ( .B1(n9734), .B2(n6791), .A(n6790), .ZN(n6792) );
  INV_X1 U8413 ( .A(n6792), .ZN(n6793) );
  OAI211_X1 U8414 ( .C1(n6795), .C2(n9736), .A(n6794), .B(n6793), .ZN(P2_U3260) );
  INV_X2 U8415 ( .A(n9921), .ZN(n9923) );
  INV_X1 U8416 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U8417 ( .A1(n6796), .A2(n9830), .ZN(n6798) );
  NAND2_X1 U8418 ( .A1(n6796), .A2(n9825), .ZN(n6940) );
  NAND2_X1 U8419 ( .A1(n6928), .A2(n6797), .ZN(n9811) );
  AND2_X1 U8420 ( .A1(n9811), .A2(n6798), .ZN(n6799) );
  NAND2_X1 U8421 ( .A1(n6800), .A2(n6799), .ZN(n6803) );
  AND2_X1 U8422 ( .A1(n6801), .A2(n6803), .ZN(n6804) );
  NAND2_X1 U8423 ( .A1(n7033), .A2(n7048), .ZN(n7988) );
  NAND2_X1 U8424 ( .A1(n9819), .A2(n6933), .ZN(n7029) );
  NAND2_X1 U8425 ( .A1(n7988), .A2(n7029), .ZN(n8146) );
  AND2_X1 U8426 ( .A1(n6801), .A2(n8146), .ZN(n6802) );
  NAND2_X1 U8427 ( .A1(n6803), .A2(n6802), .ZN(n6935) );
  OAI21_X1 U8428 ( .B1(n6804), .B2(n8146), .A(n6935), .ZN(n7053) );
  INV_X1 U8429 ( .A(n7053), .ZN(n6812) );
  NAND2_X1 U8430 ( .A1(n6805), .A2(n7999), .ZN(n9815) );
  NAND2_X1 U8431 ( .A1(n9814), .A2(n6940), .ZN(n6806) );
  XOR2_X1 U8432 ( .A(n8146), .B(n6806), .Z(n6808) );
  AOI21_X1 U8433 ( .B1(n6808), .B2(n9816), .A(n6807), .ZN(n7055) );
  NAND2_X1 U8434 ( .A1(n9831), .A2(n7048), .ZN(n6809) );
  NAND2_X1 U8435 ( .A1(n6809), .A2(n9827), .ZN(n6810) );
  NOR2_X1 U8436 ( .A1(n7037), .A2(n6810), .ZN(n7047) );
  AOI21_X1 U8437 ( .B1(n8804), .B2(n7048), .A(n7047), .ZN(n6811) );
  OAI211_X1 U8438 ( .C1(n9877), .C2(n6812), .A(n7055), .B(n6811), .ZN(n6815)
         );
  NAND2_X1 U8439 ( .A1(n6815), .A2(n9923), .ZN(n6813) );
  OAI21_X1 U8440 ( .B1(n9923), .B2(n6814), .A(n6813), .ZN(P2_U3463) );
  NAND2_X1 U8441 ( .A1(n6815), .A2(n9934), .ZN(n6816) );
  OAI21_X1 U8442 ( .B1(n9934), .B2(n6817), .A(n6816), .ZN(P2_U3524) );
  XNOR2_X1 U8443 ( .A(n6819), .B(n6818), .ZN(n6820) );
  NAND2_X1 U8444 ( .A1(n6820), .A2(n9643), .ZN(n6825) );
  NAND2_X1 U8445 ( .A1(n9306), .A2(n8985), .ZN(n6822) );
  NAND2_X1 U8446 ( .A1(n9304), .A2(n5823), .ZN(n6821) );
  NAND2_X1 U8447 ( .A1(n6822), .A2(n6821), .ZN(n7169) );
  AOI22_X1 U8448 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n6823), .B1(n9633), .B2(
        n7169), .ZN(n6824) );
  OAI211_X1 U8449 ( .C1(n9670), .C2(n8959), .A(n6825), .B(n6824), .ZN(P1_U3235) );
  NAND2_X1 U8450 ( .A1(n8416), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6902) );
  INV_X1 U8451 ( .A(n6902), .ZN(n6831) );
  INV_X1 U8452 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6830) );
  INV_X1 U8453 ( .A(n8415), .ZN(n8325) );
  INV_X1 U8454 ( .A(n6990), .ZN(n9876) );
  NAND2_X1 U8455 ( .A1(n6986), .A2(n9876), .ZN(n8142) );
  NOR3_X1 U8456 ( .A1(n8423), .A2(n8306), .A3(n8142), .ZN(n6828) );
  OAI21_X1 U8457 ( .B1(n8306), .B2(n6899), .A(n8425), .ZN(n6826) );
  AOI21_X1 U8458 ( .B1(n6826), .B2(n8436), .A(n9876), .ZN(n6827) );
  AOI211_X1 U8459 ( .C1(n8325), .C2(n6206), .A(n6828), .B(n6827), .ZN(n6829)
         );
  OAI21_X1 U8460 ( .B1(n6831), .B2(n6830), .A(n6829), .ZN(P2_U3234) );
  INV_X1 U8461 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U8462 ( .A1(n6833), .A2(n6832), .ZN(n6834) );
  AND2_X1 U8463 ( .A1(n6864), .A2(n6834), .ZN(n7129) );
  INV_X1 U8464 ( .A(n7129), .ZN(n6875) );
  NAND2_X1 U8465 ( .A1(n7882), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8466 ( .A1(n7958), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U8467 ( .A1(n7937), .A2(n7129), .ZN(n6836) );
  NAND2_X1 U8468 ( .A1(n7957), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6835) );
  NAND4_X1 U8469 ( .A1(n6838), .A2(n6837), .A3(n6836), .A4(n6835), .ZN(n8446)
         );
  AND2_X1 U8470 ( .A1(n8446), .A2(n8301), .ZN(n6843) );
  CLKBUF_X3 U8471 ( .A(n6839), .Z(n7970) );
  NAND2_X1 U8472 ( .A1(n7970), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U8473 ( .A1(n7641), .A2(n9769), .ZN(n6840) );
  OAI211_X1 U8474 ( .C1(n6842), .C2(n7977), .A(n6841), .B(n6840), .ZN(n7135)
         );
  XNOR2_X1 U8475 ( .A(n7135), .B(n4322), .ZN(n6844) );
  NAND2_X1 U8476 ( .A1(n6843), .A2(n6844), .ZN(n6847) );
  INV_X1 U8477 ( .A(n6843), .ZN(n6846) );
  INV_X1 U8478 ( .A(n6844), .ZN(n6845) );
  NAND2_X1 U8479 ( .A1(n6846), .A2(n6845), .ZN(n6904) );
  AND2_X1 U8480 ( .A1(n6847), .A2(n6904), .ZN(n6861) );
  AND2_X1 U8481 ( .A1(n8447), .A2(n8301), .ZN(n6854) );
  NAND2_X1 U8482 ( .A1(n7970), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U8483 ( .A1(n7641), .A2(n6850), .ZN(n6851) );
  OAI211_X1 U8484 ( .C1(n6853), .C2(n7977), .A(n6852), .B(n6851), .ZN(n7040)
         );
  XNOR2_X1 U8485 ( .A(n7040), .B(n4322), .ZN(n6855) );
  NAND2_X1 U8486 ( .A1(n6854), .A2(n6855), .ZN(n6858) );
  INV_X1 U8487 ( .A(n6854), .ZN(n6857) );
  INV_X1 U8488 ( .A(n6855), .ZN(n6856) );
  NAND2_X1 U8489 ( .A1(n6857), .A2(n6856), .ZN(n6859) );
  AND2_X1 U8490 ( .A1(n6858), .A2(n6859), .ZN(n6886) );
  OAI21_X1 U8491 ( .B1(n6861), .B2(n6860), .A(n6905), .ZN(n6862) );
  NAND2_X1 U8492 ( .A1(n6862), .A2(n8425), .ZN(n6874) );
  NAND2_X1 U8493 ( .A1(n7882), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6869) );
  NAND2_X1 U8494 ( .A1(n7958), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6868) );
  INV_X1 U8495 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6863) );
  NAND2_X1 U8496 ( .A1(n6864), .A2(n6863), .ZN(n6865) );
  AND2_X1 U8497 ( .A1(n6915), .A2(n6865), .ZN(n7212) );
  NAND2_X1 U8498 ( .A1(n7937), .A2(n7212), .ZN(n6867) );
  NAND2_X1 U8499 ( .A1(n7957), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6866) );
  NAND4_X1 U8500 ( .A1(n6869), .A2(n6868), .A3(n6867), .A4(n6866), .ZN(n8445)
         );
  NAND2_X1 U8501 ( .A1(n8445), .A2(n9818), .ZN(n6871) );
  NAND2_X1 U8502 ( .A1(n8447), .A2(n9821), .ZN(n6870) );
  NAND2_X1 U8503 ( .A1(n6871), .A2(n6870), .ZN(n6945) );
  AND2_X1 U8504 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9768) );
  INV_X1 U8505 ( .A(n7135), .ZN(n7181) );
  NOR2_X1 U8506 ( .A1(n8436), .A2(n7181), .ZN(n6872) );
  AOI211_X1 U8507 ( .C1(n8407), .C2(n6945), .A(n9768), .B(n6872), .ZN(n6873)
         );
  OAI211_X1 U8508 ( .C1(n8416), .C2(n6875), .A(n6874), .B(n6873), .ZN(P2_U3241) );
  NAND2_X1 U8509 ( .A1(n8407), .A2(n9821), .ZN(n8418) );
  AOI22_X1 U8510 ( .A1(n8325), .A2(n6771), .B1(n6876), .B2(n8421), .ZN(n6882)
         );
  OAI21_X1 U8511 ( .B1(n6879), .B2(n6878), .A(n6877), .ZN(n6880) );
  AOI22_X1 U8512 ( .A1(n6902), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8425), .B2(
        n6880), .ZN(n6881) );
  OAI211_X1 U8513 ( .C1(n6883), .C2(n8418), .A(n6882), .B(n6881), .ZN(P2_U3239) );
  OAI21_X1 U8514 ( .B1(n6886), .B2(n6885), .A(n6884), .ZN(n6892) );
  OAI22_X1 U8515 ( .A1(n7033), .A2(n8418), .B1(n8415), .B2(n7182), .ZN(n6891)
         );
  INV_X1 U8516 ( .A(n6887), .ZN(n7038) );
  NAND2_X1 U8517 ( .A1(n8421), .A2(n7040), .ZN(n6889) );
  OAI211_X1 U8518 ( .C1(n8416), .C2(n7038), .A(n6889), .B(n6888), .ZN(n6890)
         );
  AOI211_X1 U8519 ( .C1(n6892), .C2(n8425), .A(n6891), .B(n6890), .ZN(n6893)
         );
  INV_X1 U8520 ( .A(n6893), .ZN(P2_U3229) );
  INV_X1 U8521 ( .A(n6894), .ZN(n6895) );
  AOI21_X1 U8522 ( .B1(n6897), .B2(n6896), .A(n6895), .ZN(n6898) );
  OAI22_X1 U8523 ( .A1(n8436), .A2(n9883), .B1(n6898), .B2(n8423), .ZN(n6901)
         );
  OAI22_X1 U8524 ( .A1(n6899), .A2(n8418), .B1(n8415), .B2(n6928), .ZN(n6900)
         );
  AOI211_X1 U8525 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(n6902), .A(n6901), .B(
        n6900), .ZN(n6903) );
  INV_X1 U8526 ( .A(n6903), .ZN(P2_U3224) );
  OR2_X1 U8527 ( .A1(n7977), .A2(n6906), .ZN(n6912) );
  OAI22_X1 U8528 ( .A1(n6907), .A2(n6909), .B1(n7832), .B2(n6908), .ZN(n6910)
         );
  INV_X1 U8529 ( .A(n6910), .ZN(n6911) );
  XNOR2_X1 U8530 ( .A(n7199), .B(n8300), .ZN(n7006) );
  NAND2_X1 U8531 ( .A1(n8445), .A2(n8301), .ZN(n7005) );
  XNOR2_X1 U8532 ( .A(n7006), .B(n7005), .ZN(n7002) );
  XNOR2_X1 U8533 ( .A(n7001), .B(n7002), .ZN(n6924) );
  NAND2_X1 U8534 ( .A1(n8421), .A2(n7199), .ZN(n6913) );
  NAND2_X1 U8535 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9780) );
  NAND2_X1 U8536 ( .A1(n6913), .A2(n9780), .ZN(n6922) );
  NAND2_X1 U8537 ( .A1(n7882), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U8538 ( .A1(n7958), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6919) );
  INV_X1 U8539 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6914) );
  NAND2_X1 U8540 ( .A1(n6915), .A2(n6914), .ZN(n6916) );
  AND2_X1 U8541 ( .A1(n7017), .A2(n6916), .ZN(n7202) );
  NAND2_X1 U8542 ( .A1(n7937), .A2(n7202), .ZN(n6918) );
  NAND2_X1 U8543 ( .A1(n7957), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6917) );
  NAND4_X1 U8544 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(n8444)
         );
  INV_X1 U8545 ( .A(n8444), .ZN(n7186) );
  OAI22_X1 U8546 ( .A1(n7182), .A2(n8418), .B1(n8415), .B2(n7186), .ZN(n6921)
         );
  AOI211_X1 U8547 ( .C1(n7212), .C2(n8433), .A(n6922), .B(n6921), .ZN(n6923)
         );
  OAI21_X1 U8548 ( .B1(n6924), .B2(n8423), .A(n6923), .ZN(P2_U3215) );
  XNOR2_X1 U8549 ( .A(n6926), .B(n6925), .ZN(n6932) );
  INV_X1 U8550 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9833) );
  NAND2_X1 U8551 ( .A1(n8421), .A2(n9825), .ZN(n6927) );
  OAI21_X1 U8552 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n9833), .A(n6927), .ZN(n6930) );
  OAI22_X1 U8553 ( .A1(n6928), .A2(n8418), .B1(n8415), .B2(n7033), .ZN(n6929)
         );
  AOI211_X1 U8554 ( .C1(n8433), .C2(n9833), .A(n6930), .B(n6929), .ZN(n6931)
         );
  OAI21_X1 U8555 ( .B1(n6932), .B2(n8423), .A(n6931), .ZN(P2_U3220) );
  INV_X1 U8556 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U8557 ( .A1(n7033), .A2(n6933), .ZN(n6934) );
  NAND2_X1 U8558 ( .A1(n6935), .A2(n6934), .ZN(n7035) );
  NAND2_X1 U8559 ( .A1(n6936), .A2(n7040), .ZN(n7991) );
  NAND2_X1 U8560 ( .A1(n7991), .A2(n8006), .ZN(n8148) );
  NAND2_X1 U8561 ( .A1(n7035), .A2(n8148), .ZN(n7034) );
  NAND2_X1 U8562 ( .A1(n6936), .A2(n9894), .ZN(n6937) );
  NAND2_X1 U8563 ( .A1(n7034), .A2(n6937), .ZN(n6938) );
  NAND2_X1 U8564 ( .A1(n7182), .A2(n7135), .ZN(n8014) );
  NAND2_X1 U8565 ( .A1(n8446), .A2(n7181), .ZN(n8012) );
  NAND2_X1 U8566 ( .A1(n6938), .A2(n8149), .ZN(n7184) );
  OAI21_X1 U8567 ( .B1(n6938), .B2(n8149), .A(n7184), .ZN(n6939) );
  INV_X1 U8568 ( .A(n6939), .ZN(n7137) );
  AND2_X1 U8569 ( .A1(n6940), .A2(n7988), .ZN(n7992) );
  NAND2_X1 U8570 ( .A1(n9814), .A2(n7992), .ZN(n7030) );
  AND2_X1 U8571 ( .A1(n8006), .A2(n7029), .ZN(n8008) );
  NAND2_X1 U8572 ( .A1(n7030), .A2(n8008), .ZN(n6943) );
  NAND2_X1 U8573 ( .A1(n6943), .A2(n7991), .ZN(n6942) );
  INV_X1 U8574 ( .A(n8149), .ZN(n6941) );
  NAND3_X1 U8575 ( .A1(n6943), .A2(n8149), .A3(n7991), .ZN(n6944) );
  INV_X1 U8576 ( .A(n9816), .ZN(n8605) );
  AOI21_X1 U8577 ( .B1(n7190), .B2(n6944), .A(n8605), .ZN(n6946) );
  NOR2_X1 U8578 ( .A1(n6946), .A2(n6945), .ZN(n7132) );
  NAND2_X1 U8579 ( .A1(n7037), .A2(n9894), .ZN(n7036) );
  OR2_X1 U8580 ( .A1(n7036), .A2(n7135), .ZN(n7200) );
  INV_X1 U8581 ( .A(n7200), .ZN(n7211) );
  AOI211_X1 U8582 ( .C1(n7135), .C2(n7036), .A(n9915), .B(n7211), .ZN(n7130)
         );
  AOI21_X1 U8583 ( .B1(n8804), .B2(n7135), .A(n7130), .ZN(n6947) );
  OAI211_X1 U8584 ( .C1(n7137), .C2(n9877), .A(n7132), .B(n6947), .ZN(n6949)
         );
  NAND2_X1 U8585 ( .A1(n6949), .A2(n9923), .ZN(n6948) );
  OAI21_X1 U8586 ( .B1(n9923), .B2(n10091), .A(n6948), .ZN(P2_U3469) );
  NAND2_X1 U8587 ( .A1(n6949), .A2(n9934), .ZN(n6950) );
  OAI21_X1 U8588 ( .B1(n9934), .B2(n6386), .A(n6950), .ZN(P2_U3526) );
  NAND2_X1 U8589 ( .A1(n7564), .A2(n8704), .ZN(n9835) );
  NAND2_X1 U8590 ( .A1(n6982), .A2(n8142), .ZN(n6951) );
  INV_X1 U8591 ( .A(n6951), .ZN(n9878) );
  NAND2_X1 U8592 ( .A1(n6951), .A2(n9816), .ZN(n6953) );
  NAND2_X1 U8593 ( .A1(n6206), .A2(n9818), .ZN(n6952) );
  NAND2_X1 U8594 ( .A1(n6953), .A2(n6952), .ZN(n9879) );
  INV_X2 U8595 ( .A(n7366), .ZN(n9834) );
  AOI22_X1 U8596 ( .A1(n9838), .A2(n9879), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n9834), .ZN(n6956) );
  INV_X1 U8597 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6954) );
  OR2_X1 U8598 ( .A1(n9838), .A2(n6954), .ZN(n6955) );
  OAI211_X1 U8599 ( .C1(n8718), .C2(n9878), .A(n6956), .B(n6955), .ZN(n6957)
         );
  AOI21_X1 U8600 ( .B1(n9835), .B2(n6990), .A(n6957), .ZN(n6958) );
  INV_X1 U8601 ( .A(n6958), .ZN(P2_U3296) );
  INV_X1 U8602 ( .A(n7820), .ZN(n6980) );
  AOI22_X1 U8603 ( .A1(n9051), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9537), .ZN(n6959) );
  OAI21_X1 U8604 ( .B1(n6980), .B2(n8245), .A(n6959), .ZN(P1_U3335) );
  INV_X1 U8605 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6960) );
  AOI22_X1 U8606 ( .A1(n7543), .A2(n6960), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n7802), .ZN(n6965) );
  NAND2_X1 U8607 ( .A1(n7642), .A2(n6961), .ZN(n6963) );
  NAND2_X1 U8608 ( .A1(n6963), .A2(n6962), .ZN(n6964) );
  NOR2_X1 U8609 ( .A1(n6965), .A2(n6964), .ZN(n7545) );
  AOI21_X1 U8610 ( .B1(n6965), .B2(n6964), .A(n7545), .ZN(n6977) );
  INV_X1 U8611 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U8612 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8369) );
  OAI21_X1 U8613 ( .B1(n8484), .B2(n6966), .A(n8369), .ZN(n6967) );
  AOI21_X1 U8614 ( .B1(n9802), .B2(n7543), .A(n6967), .ZN(n6976) );
  NOR2_X1 U8615 ( .A1(n7642), .A2(n6968), .ZN(n6970) );
  NOR2_X1 U8616 ( .A1(n6970), .A2(n6969), .ZN(n6974) );
  INV_X1 U8617 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6972) );
  NAND2_X1 U8618 ( .A1(n7543), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7540) );
  INV_X1 U8619 ( .A(n7540), .ZN(n6971) );
  AOI21_X1 U8620 ( .B1(n6972), .B2(n7802), .A(n6971), .ZN(n6973) );
  NAND2_X1 U8621 ( .A1(n6973), .A2(n6974), .ZN(n7539) );
  OAI211_X1 U8622 ( .C1(n6974), .C2(n6973), .A(n9797), .B(n7539), .ZN(n6975)
         );
  OAI211_X1 U8623 ( .C1(n6977), .C2(n8475), .A(n6976), .B(n6975), .ZN(P2_U3261) );
  INV_X1 U8624 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U8625 ( .A1(n6978), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6979) );
  XNOR2_X1 U8626 ( .A(n6979), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8464) );
  INV_X1 U8627 ( .A(n8464), .ZN(n8470) );
  OAI222_X1 U8628 ( .A1(n8831), .A2(n7821), .B1(n8830), .B2(n6980), .C1(
        P2_U3152), .C2(n8470), .ZN(P2_U3340) );
  INV_X1 U8629 ( .A(n8143), .ZN(n6985) );
  INV_X1 U8630 ( .A(n6982), .ZN(n6983) );
  NAND2_X1 U8631 ( .A1(n6981), .A2(n6983), .ZN(n6984) );
  OAI211_X1 U8632 ( .C1(n8145), .C2(n6985), .A(n6984), .B(n9816), .ZN(n6988)
         );
  AOI22_X1 U8633 ( .A1(n9821), .A2(n6986), .B1(n9820), .B2(n9818), .ZN(n6987)
         );
  NAND2_X1 U8634 ( .A1(n6988), .A2(n6987), .ZN(n9884) );
  NOR2_X1 U8635 ( .A1(n9838), .A2(n6257), .ZN(n6995) );
  INV_X1 U8636 ( .A(n6989), .ZN(n6992) );
  AOI21_X1 U8637 ( .B1(n6998), .B2(n6990), .A(n9915), .ZN(n6991) );
  NAND2_X1 U8638 ( .A1(n6992), .A2(n6991), .ZN(n9882) );
  OAI22_X1 U8639 ( .A1(n7045), .A2(n9882), .B1(n6993), .B2(n7366), .ZN(n6994)
         );
  AOI211_X1 U8640 ( .C1(n9838), .C2(n9884), .A(n6995), .B(n6994), .ZN(n7000)
         );
  INV_X1 U8641 ( .A(n8718), .ZN(n8566) );
  OAI21_X1 U8642 ( .B1(n6981), .B2(n6997), .A(n6996), .ZN(n9886) );
  INV_X1 U8643 ( .A(n8704), .ZN(n7684) );
  AOI22_X1 U8644 ( .A1(n8566), .A2(n9886), .B1(n7684), .B2(n6998), .ZN(n6999)
         );
  NAND2_X1 U8645 ( .A1(n7000), .A2(n6999), .ZN(P2_U3295) );
  INV_X1 U8646 ( .A(n7005), .ZN(n7008) );
  INV_X1 U8647 ( .A(n7006), .ZN(n7007) );
  NAND2_X1 U8648 ( .A1(n7008), .A2(n7007), .ZN(n7070) );
  NAND2_X1 U8649 ( .A1(n7072), .A2(n7070), .ZN(n7102) );
  OR2_X1 U8650 ( .A1(n7009), .A2(n7977), .ZN(n7014) );
  OAI22_X1 U8651 ( .A1(n6907), .A2(n7011), .B1(n7832), .B2(n7010), .ZN(n7012)
         );
  INV_X1 U8652 ( .A(n7012), .ZN(n7013) );
  XNOR2_X1 U8653 ( .A(n7282), .B(n4322), .ZN(n7068) );
  NAND2_X1 U8654 ( .A1(n8444), .A2(n8301), .ZN(n7066) );
  XNOR2_X1 U8655 ( .A(n7068), .B(n7066), .ZN(n7101) );
  XNOR2_X1 U8656 ( .A(n7102), .B(n7101), .ZN(n7026) );
  INV_X1 U8657 ( .A(n7282), .ZN(n7205) );
  OAI21_X1 U8658 ( .B1(n8436), .B2(n7205), .A(n7015), .ZN(n7024) );
  INV_X1 U8659 ( .A(n8445), .ZN(n7194) );
  NAND2_X1 U8660 ( .A1(n7957), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U8661 ( .A1(n7882), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7021) );
  INV_X1 U8662 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7016) );
  NAND2_X1 U8663 ( .A1(n7017), .A2(n7016), .ZN(n7018) );
  AND2_X1 U8664 ( .A1(n7083), .A2(n7018), .ZN(n7232) );
  NAND2_X1 U8665 ( .A1(n7937), .A2(n7232), .ZN(n7020) );
  NAND2_X1 U8666 ( .A1(n7958), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7019) );
  NAND4_X1 U8667 ( .A1(n7022), .A2(n7021), .A3(n7020), .A4(n7019), .ZN(n8443)
         );
  OAI22_X1 U8668 ( .A1(n7194), .A2(n8418), .B1(n8415), .B2(n7356), .ZN(n7023)
         );
  AOI211_X1 U8669 ( .C1(n7202), .C2(n8433), .A(n7024), .B(n7023), .ZN(n7025)
         );
  OAI21_X1 U8670 ( .B1(n7026), .B2(n8423), .A(n7025), .ZN(P2_U3223) );
  INV_X1 U8671 ( .A(n7831), .ZN(n7028) );
  OAI222_X1 U8672 ( .A1(n8831), .A2(n7833), .B1(n8830), .B2(n7028), .C1(n7982), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8673 ( .A1(n9274), .A2(P1_U3084), .B1(n9539), .B2(n7028), .C1(
        n7027), .C2(n8242), .ZN(P1_U3334) );
  NAND2_X1 U8674 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  XOR2_X1 U8675 ( .A(n8148), .B(n7031), .Z(n7032) );
  OAI222_X1 U8676 ( .A1(n8662), .A2(n7182), .B1(n8664), .B2(n7033), .C1(n8605), 
        .C2(n7032), .ZN(n9895) );
  INV_X1 U8677 ( .A(n9895), .ZN(n7044) );
  INV_X2 U8678 ( .A(n9838), .ZN(n8713) );
  OAI21_X1 U8679 ( .B1(n7035), .B2(n8148), .A(n7034), .ZN(n9897) );
  OAI211_X1 U8680 ( .C1(n7037), .C2(n9894), .A(n7036), .B(n9827), .ZN(n9893)
         );
  OAI22_X1 U8681 ( .A1(n9838), .A2(n6408), .B1(n7038), .B2(n7366), .ZN(n7039)
         );
  AOI21_X1 U8682 ( .B1(n7684), .B2(n7040), .A(n7039), .ZN(n7041) );
  OAI21_X1 U8683 ( .B1(n7045), .B2(n9893), .A(n7041), .ZN(n7042) );
  AOI21_X1 U8684 ( .B1(n8566), .B2(n9897), .A(n7042), .ZN(n7043) );
  OAI21_X1 U8685 ( .B1(n7044), .B2(n8713), .A(n7043), .ZN(P2_U3291) );
  INV_X1 U8686 ( .A(n7045), .ZN(n8681) );
  AOI22_X1 U8687 ( .A1(n8681), .A2(n7047), .B1(n7046), .B2(n9834), .ZN(n7050)
         );
  NAND2_X1 U8688 ( .A1(n7684), .A2(n7048), .ZN(n7049) );
  OAI211_X1 U8689 ( .C1(n7051), .C2(n9838), .A(n7050), .B(n7049), .ZN(n7052)
         );
  AOI21_X1 U8690 ( .B1(n8566), .B2(n7053), .A(n7052), .ZN(n7054) );
  OAI21_X1 U8691 ( .B1(n7055), .B2(n8713), .A(n7054), .ZN(P2_U3292) );
  OR2_X1 U8692 ( .A1(n7056), .A2(n7977), .ZN(n7060) );
  OAI22_X1 U8693 ( .A1(n6907), .A2(n7057), .B1(n7832), .B2(n8454), .ZN(n7058)
         );
  INV_X1 U8694 ( .A(n7058), .ZN(n7059) );
  XNOR2_X1 U8695 ( .A(n7350), .B(n8300), .ZN(n7061) );
  NAND2_X1 U8696 ( .A1(n8443), .A2(n8301), .ZN(n7062) );
  NAND2_X1 U8697 ( .A1(n7061), .A2(n7062), .ZN(n7074) );
  INV_X1 U8698 ( .A(n7061), .ZN(n7064) );
  INV_X1 U8699 ( .A(n7062), .ZN(n7063) );
  NAND2_X1 U8700 ( .A1(n7064), .A2(n7063), .ZN(n7065) );
  NAND2_X1 U8701 ( .A1(n7074), .A2(n7065), .ZN(n7108) );
  INV_X1 U8702 ( .A(n7108), .ZN(n7069) );
  INV_X1 U8703 ( .A(n7066), .ZN(n7067) );
  NAND2_X1 U8704 ( .A1(n7068), .A2(n7067), .ZN(n7103) );
  AND2_X1 U8705 ( .A1(n7070), .A2(n7073), .ZN(n7071) );
  AND2_X1 U8706 ( .A1(n7074), .A2(n7105), .ZN(n7075) );
  NAND2_X1 U8707 ( .A1(n7076), .A2(n7969), .ZN(n7081) );
  OAI22_X1 U8708 ( .A1(n6907), .A2(n7078), .B1(n7832), .B2(n7077), .ZN(n7079)
         );
  INV_X1 U8709 ( .A(n7079), .ZN(n7080) );
  XNOR2_X1 U8710 ( .A(n7569), .B(n8300), .ZN(n7238) );
  NAND2_X1 U8711 ( .A1(n7882), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7088) );
  NAND2_X1 U8712 ( .A1(n7957), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7087) );
  NAND2_X1 U8713 ( .A1(n7083), .A2(n7082), .ZN(n7084) );
  AND2_X1 U8714 ( .A1(n7090), .A2(n7084), .ZN(n7365) );
  NAND2_X1 U8715 ( .A1(n7937), .A2(n7365), .ZN(n7086) );
  NAND2_X1 U8716 ( .A1(n7958), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7085) );
  NAND4_X1 U8717 ( .A1(n7088), .A2(n7087), .A3(n7086), .A4(n7085), .ZN(n8442)
         );
  NAND2_X1 U8718 ( .A1(n8442), .A2(n8301), .ZN(n7237) );
  XNOR2_X1 U8719 ( .A(n7238), .B(n7237), .ZN(n7239) );
  XNOR2_X1 U8720 ( .A(n7240), .B(n7239), .ZN(n7100) );
  NAND2_X1 U8721 ( .A1(n7882), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7095) );
  NAND2_X1 U8722 ( .A1(n7958), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7094) );
  INV_X1 U8723 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7089) );
  NAND2_X1 U8724 ( .A1(n7090), .A2(n7089), .ZN(n7091) );
  AND2_X1 U8725 ( .A1(n7248), .A2(n7091), .ZN(n7561) );
  NAND2_X1 U8726 ( .A1(n7937), .A2(n7561), .ZN(n7093) );
  NAND2_X1 U8727 ( .A1(n7957), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7092) );
  NAND4_X1 U8728 ( .A1(n7095), .A2(n7094), .A3(n7093), .A4(n7092), .ZN(n8441)
         );
  INV_X1 U8729 ( .A(n8418), .ZN(n8376) );
  AOI22_X1 U8730 ( .A1(n8376), .A2(n8443), .B1(n7365), .B2(n8433), .ZN(n7097)
         );
  OAI211_X1 U8731 ( .C1(n7555), .C2(n8415), .A(n7097), .B(n7096), .ZN(n7098)
         );
  AOI21_X1 U8732 ( .B1(n7569), .B2(n8421), .A(n7098), .ZN(n7099) );
  OAI21_X1 U8733 ( .B1(n7100), .B2(n8423), .A(n7099), .ZN(P2_U3219) );
  NAND2_X1 U8734 ( .A1(n7102), .A2(n7101), .ZN(n7104) );
  NAND2_X1 U8735 ( .A1(n7104), .A2(n7103), .ZN(n7109) );
  NAND2_X1 U8736 ( .A1(n7106), .A2(n7105), .ZN(n7107) );
  AOI21_X1 U8737 ( .B1(n7109), .B2(n7108), .A(n7107), .ZN(n7113) );
  AOI22_X1 U8738 ( .A1(n8376), .A2(n8444), .B1(n7232), .B2(n8433), .ZN(n7110)
         );
  NAND2_X1 U8739 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8452) );
  OAI211_X1 U8740 ( .C1(n7558), .C2(n8415), .A(n7110), .B(n8452), .ZN(n7111)
         );
  AOI21_X1 U8741 ( .B1(n7350), .B2(n8421), .A(n7111), .ZN(n7112) );
  OAI21_X1 U8742 ( .B1(n7113), .B2(n8423), .A(n7112), .ZN(P2_U3233) );
  AOI21_X1 U8743 ( .B1(n7115), .B2(n6704), .A(n7114), .ZN(n7117) );
  AOI22_X1 U8744 ( .A1(n7124), .A2(n5214), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n7415), .ZN(n7116) );
  NOR2_X1 U8745 ( .A1(n7117), .A2(n7116), .ZN(n7414) );
  AOI21_X1 U8746 ( .B1(n7117), .B2(n7116), .A(n7414), .ZN(n7126) );
  INV_X1 U8747 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7118) );
  NAND2_X1 U8748 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8842) );
  OAI21_X1 U8749 ( .B1(n10167), .B2(n7118), .A(n8842), .ZN(n7123) );
  AOI21_X1 U8750 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7120), .A(n7119), .ZN(
        n7408) );
  XNOR2_X1 U8751 ( .A(n7415), .B(n7408), .ZN(n7121) );
  NOR2_X1 U8752 ( .A1(n9385), .A2(n7121), .ZN(n7409) );
  AOI211_X1 U8753 ( .C1(n7121), .C2(n9385), .A(n7409), .B(n10154), .ZN(n7122)
         );
  AOI211_X1 U8754 ( .C1(n9036), .C2(n7124), .A(n7123), .B(n7122), .ZN(n7125)
         );
  OAI21_X1 U8755 ( .B1(n7126), .B2(n10162), .A(n7125), .ZN(P1_U3255) );
  INV_X1 U8756 ( .A(n7847), .ZN(n7163) );
  OAI222_X1 U8757 ( .A1(n8830), .A2(n7163), .B1(P2_U3152), .B2(n7128), .C1(
        n7127), .C2(n8831), .ZN(P2_U3338) );
  AOI22_X1 U8758 ( .A1(n7130), .A2(n8681), .B1(n7129), .B2(n9834), .ZN(n7131)
         );
  OAI21_X1 U8759 ( .B1(n6407), .B2(n9838), .A(n7131), .ZN(n7134) );
  NOR2_X1 U8760 ( .A1(n7132), .A2(n8713), .ZN(n7133) );
  AOI211_X1 U8761 ( .C1(n7684), .C2(n7135), .A(n7134), .B(n7133), .ZN(n7136)
         );
  OAI21_X1 U8762 ( .B1(n7137), .B2(n8718), .A(n7136), .ZN(P2_U3290) );
  NAND4_X1 U8763 ( .A1(n7141), .A2(n7140), .A3(n7139), .A4(n7138), .ZN(n7143)
         );
  AOI22_X1 U8764 ( .A1(n9377), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9594), .ZN(n7146) );
  NOR2_X2 U8765 ( .A1(n9377), .A2(n7142), .ZN(n9595) );
  NOR2_X1 U8766 ( .A1(n7143), .A2(n9061), .ZN(n9599) );
  NAND2_X1 U8767 ( .A1(n9599), .A2(n9713), .ZN(n9389) );
  OAI21_X1 U8768 ( .B1(n9595), .B2(n9566), .A(n7144), .ZN(n7145) );
  OAI211_X1 U8769 ( .C1(n7147), .C2(n9605), .A(n7146), .B(n7145), .ZN(P1_U3291) );
  NAND2_X1 U8770 ( .A1(n5823), .A2(n5357), .ZN(n7148) );
  NAND2_X1 U8771 ( .A1(n7166), .A2(n7168), .ZN(n7165) );
  OR2_X1 U8772 ( .A1(n5838), .A2(n7177), .ZN(n7150) );
  NAND2_X1 U8773 ( .A1(n7165), .A2(n7150), .ZN(n7151) );
  NAND2_X1 U8774 ( .A1(n7151), .A2(n7153), .ZN(n7264) );
  OAI21_X1 U8775 ( .B1(n7151), .B2(n7153), .A(n7264), .ZN(n9679) );
  INV_X1 U8776 ( .A(n9679), .ZN(n7161) );
  NAND3_X1 U8777 ( .A1(n9327), .A2(n7152), .A3(n5800), .ZN(n9373) );
  XNOR2_X1 U8778 ( .A(n7153), .B(n5588), .ZN(n7155) );
  INV_X1 U8779 ( .A(n9497), .ZN(n9721) );
  NAND2_X1 U8780 ( .A1(n9679), .A2(n9721), .ZN(n7154) );
  AOI22_X1 U8781 ( .A1(n9306), .A2(n8984), .B1(n9304), .B2(n5838), .ZN(n9622)
         );
  OAI211_X1 U8782 ( .C1(n9553), .C2(n7155), .A(n7154), .B(n9622), .ZN(n9677)
         );
  NAND2_X1 U8783 ( .A1(n9677), .A2(n9327), .ZN(n7160) );
  AND2_X1 U8784 ( .A1(n7173), .A2(n9626), .ZN(n7156) );
  OR2_X1 U8785 ( .A1(n7156), .A2(n7530), .ZN(n9676) );
  AOI22_X1 U8786 ( .A1(n9605), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9594), .B2(
        n5419), .ZN(n7157) );
  OAI21_X1 U8787 ( .B1(n9676), .B2(n9389), .A(n7157), .ZN(n7158) );
  AOI21_X1 U8788 ( .B1(n9595), .B2(n9626), .A(n7158), .ZN(n7159) );
  OAI211_X1 U8789 ( .C1(n7161), .C2(n9373), .A(n7160), .B(n7159), .ZN(P1_U3288) );
  OAI222_X1 U8790 ( .A1(P1_U3084), .A2(n7164), .B1(n8245), .B2(n7163), .C1(
        n7162), .C2(n8242), .ZN(P1_U3333) );
  OAI21_X1 U8791 ( .B1(n7166), .B2(n7168), .A(n7165), .ZN(n9673) );
  INV_X1 U8792 ( .A(n9673), .ZN(n7180) );
  XNOR2_X1 U8793 ( .A(n7167), .B(n7168), .ZN(n7171) );
  AOI21_X1 U8794 ( .B1(n9673), .B2(n9721), .A(n7169), .ZN(n7170) );
  OAI21_X1 U8795 ( .B1(n9553), .B2(n7171), .A(n7170), .ZN(n9671) );
  NAND2_X1 U8796 ( .A1(n9671), .A2(n9327), .ZN(n7179) );
  INV_X1 U8797 ( .A(n9599), .ZN(n7336) );
  NAND2_X1 U8798 ( .A1(n7177), .A2(n7172), .ZN(n7174) );
  NAND3_X1 U8799 ( .A1(n7174), .A2(n7173), .A3(n9713), .ZN(n9669) );
  INV_X2 U8800 ( .A(n9327), .ZN(n9605) );
  AOI22_X1 U8801 ( .A1(n9594), .A2(P1_REG3_REG_2__SCAN_IN), .B1(
        P1_REG2_REG_2__SCAN_IN), .B2(n9605), .ZN(n7175) );
  OAI21_X1 U8802 ( .B1(n7336), .B2(n9669), .A(n7175), .ZN(n7176) );
  AOI21_X1 U8803 ( .B1(n9595), .B2(n7177), .A(n7176), .ZN(n7178) );
  OAI211_X1 U8804 ( .C1(n7180), .C2(n9373), .A(n7179), .B(n7178), .ZN(P1_U3289) );
  NAND2_X1 U8805 ( .A1(n7182), .A2(n7181), .ZN(n7183) );
  NAND2_X1 U8806 ( .A1(n7184), .A2(n7183), .ZN(n7217) );
  NAND2_X1 U8807 ( .A1(n7194), .A2(n7199), .ZN(n8018) );
  INV_X1 U8808 ( .A(n7199), .ZN(n9901) );
  NAND2_X1 U8809 ( .A1(n8445), .A2(n9901), .ZN(n8019) );
  NAND2_X1 U8810 ( .A1(n8018), .A2(n8019), .ZN(n8150) );
  NAND2_X1 U8811 ( .A1(n7194), .A2(n9901), .ZN(n7185) );
  NAND2_X1 U8812 ( .A1(n7205), .A2(n8444), .ZN(n8021) );
  NAND2_X1 U8813 ( .A1(n7186), .A2(n7282), .ZN(n8022) );
  INV_X1 U8814 ( .A(n8152), .ZN(n7187) );
  NAND2_X1 U8815 ( .A1(n7188), .A2(n8152), .ZN(n7189) );
  AND2_X1 U8816 ( .A1(n7221), .A2(n7189), .ZN(n7281) );
  INV_X1 U8817 ( .A(n8670), .ZN(n7681) );
  INV_X1 U8818 ( .A(n8018), .ZN(n7191) );
  NAND2_X1 U8819 ( .A1(n7192), .A2(n7187), .ZN(n7193) );
  AOI21_X1 U8820 ( .B1(n7225), .B2(n7193), .A(n8605), .ZN(n7196) );
  OAI22_X1 U8821 ( .A1(n7194), .A2(n8664), .B1(n7356), .B2(n8662), .ZN(n7195)
         );
  AOI211_X1 U8822 ( .C1(n7281), .C2(n7681), .A(n7196), .B(n7195), .ZN(n7285)
         );
  INV_X1 U8823 ( .A(n7197), .ZN(n7198) );
  NAND2_X1 U8824 ( .A1(n9838), .A2(n7198), .ZN(n8678) );
  INV_X1 U8825 ( .A(n8678), .ZN(n7689) );
  NOR2_X1 U8826 ( .A1(n7200), .A2(n7199), .ZN(n7201) );
  INV_X1 U8827 ( .A(n7201), .ZN(n7210) );
  AND2_X2 U8828 ( .A1(n7201), .A2(n7205), .ZN(n7230) );
  AOI21_X1 U8829 ( .B1(n7282), .B2(n7210), .A(n7230), .ZN(n7283) );
  NAND2_X1 U8830 ( .A1(n7283), .A2(n8716), .ZN(n7204) );
  AOI22_X1 U8831 ( .A1(n8713), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7202), .B2(
        n9834), .ZN(n7203) );
  OAI211_X1 U8832 ( .C1(n7205), .C2(n8704), .A(n7204), .B(n7203), .ZN(n7206)
         );
  AOI21_X1 U8833 ( .B1(n7281), .B2(n7689), .A(n7206), .ZN(n7207) );
  OAI21_X1 U8834 ( .B1(n7285), .B2(n8713), .A(n7207), .ZN(P2_U3288) );
  XOR2_X1 U8835 ( .A(n8150), .B(n7208), .Z(n7209) );
  AOI222_X1 U8836 ( .A1(n9816), .A2(n7209), .B1(n8444), .B2(n9818), .C1(n8446), 
        .C2(n9821), .ZN(n9900) );
  OAI211_X1 U8837 ( .C1(n9901), .C2(n7211), .A(n7210), .B(n9827), .ZN(n9899)
         );
  INV_X1 U8838 ( .A(n9899), .ZN(n7215) );
  AOI22_X1 U8839 ( .A1(n8713), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7212), .B2(
        n9834), .ZN(n7213) );
  OAI21_X1 U8840 ( .B1(n9901), .B2(n8704), .A(n7213), .ZN(n7214) );
  AOI21_X1 U8841 ( .B1(n7215), .B2(n8681), .A(n7214), .ZN(n7219) );
  OAI21_X1 U8842 ( .B1(n7217), .B2(n8150), .A(n7216), .ZN(n9903) );
  NAND2_X1 U8843 ( .A1(n9903), .A2(n8566), .ZN(n7218) );
  OAI211_X1 U8844 ( .C1(n9900), .C2(n8713), .A(n7219), .B(n7218), .ZN(P2_U3289) );
  NAND2_X1 U8845 ( .A1(n7282), .A2(n8444), .ZN(n7220) );
  NAND2_X1 U8846 ( .A1(n7221), .A2(n7220), .ZN(n7223) );
  INV_X1 U8847 ( .A(n7223), .ZN(n7222) );
  NAND2_X1 U8848 ( .A1(n7350), .A2(n7356), .ZN(n8023) );
  NAND2_X1 U8849 ( .A1(n7223), .A2(n8153), .ZN(n7224) );
  NAND2_X1 U8850 ( .A1(n7352), .A2(n7224), .ZN(n9910) );
  INV_X1 U8851 ( .A(n8153), .ZN(n7226) );
  XNOR2_X1 U8852 ( .A(n7357), .B(n7226), .ZN(n7228) );
  AOI22_X1 U8853 ( .A1(n9821), .A2(n8444), .B1(n8442), .B2(n9818), .ZN(n7227)
         );
  OAI21_X1 U8854 ( .B1(n7228), .B2(n8605), .A(n7227), .ZN(n7229) );
  AOI21_X1 U8855 ( .B1(n9910), .B2(n7681), .A(n7229), .ZN(n9912) );
  INV_X1 U8856 ( .A(n7350), .ZN(n9906) );
  OR2_X1 U8857 ( .A1(n7230), .A2(n9906), .ZN(n7231) );
  NAND2_X1 U8858 ( .A1(n7363), .A2(n7231), .ZN(n9907) );
  AOI22_X1 U8859 ( .A1(n8713), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7232), .B2(
        n9834), .ZN(n7234) );
  NAND2_X1 U8860 ( .A1(n7684), .A2(n7350), .ZN(n7233) );
  OAI211_X1 U8861 ( .C1(n9907), .C2(n7564), .A(n7234), .B(n7233), .ZN(n7235)
         );
  AOI21_X1 U8862 ( .B1(n9910), .B2(n7689), .A(n7235), .ZN(n7236) );
  OAI21_X1 U8863 ( .B1(n9912), .B2(n8713), .A(n7236), .ZN(P2_U3287) );
  NAND2_X1 U8864 ( .A1(n7241), .A2(n7969), .ZN(n7246) );
  OAI22_X1 U8865 ( .A1(n6907), .A2(n7243), .B1(n7832), .B2(n7242), .ZN(n7244)
         );
  INV_X1 U8866 ( .A(n7244), .ZN(n7245) );
  XNOR2_X1 U8867 ( .A(n8041), .B(n4322), .ZN(n7468) );
  NAND2_X1 U8868 ( .A1(n8441), .A2(n8301), .ZN(n7466) );
  XNOR2_X1 U8869 ( .A(n7468), .B(n7466), .ZN(n7464) );
  XNOR2_X1 U8870 ( .A(n7465), .B(n7464), .ZN(n7258) );
  NAND2_X1 U8871 ( .A1(n7957), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7253) );
  NAND2_X1 U8872 ( .A1(n7882), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7252) );
  NAND2_X1 U8873 ( .A1(n7248), .A2(n7247), .ZN(n7249) );
  AND2_X1 U8874 ( .A1(n7476), .A2(n7249), .ZN(n7760) );
  NAND2_X1 U8875 ( .A1(n7937), .A2(n7760), .ZN(n7251) );
  NAND2_X1 U8876 ( .A1(n7958), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7250) );
  NAND4_X1 U8877 ( .A1(n7253), .A2(n7252), .A3(n7251), .A4(n7250), .ZN(n8440)
         );
  AOI22_X1 U8878 ( .A1(n8376), .A2(n8442), .B1(n7561), .B2(n8433), .ZN(n7255)
         );
  OAI211_X1 U8879 ( .C1(n7678), .C2(n8415), .A(n7255), .B(n7254), .ZN(n7256)
         );
  AOI21_X1 U8880 ( .B1(n8041), .B2(n8421), .A(n7256), .ZN(n7257) );
  OAI21_X1 U8881 ( .B1(n7258), .B2(n8423), .A(n7257), .ZN(P2_U3238) );
  INV_X1 U8882 ( .A(n7796), .ZN(n7292) );
  OAI222_X1 U8883 ( .A1(n8830), .A2(n7292), .B1(P2_U3152), .B2(n7260), .C1(
        n7259), .C2(n8831), .ZN(P2_U3337) );
  INV_X1 U8884 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7278) );
  OR2_X1 U8885 ( .A1(n8985), .A2(n9626), .ZN(n7263) );
  NAND2_X1 U8886 ( .A1(n7264), .A2(n7263), .ZN(n7522) );
  NAND2_X1 U8887 ( .A1(n7522), .A2(n7523), .ZN(n7521) );
  INV_X1 U8888 ( .A(n7535), .ZN(n9682) );
  OR2_X1 U8889 ( .A1(n8984), .A2(n9682), .ZN(n7266) );
  INV_X1 U8890 ( .A(n7341), .ZN(n7268) );
  AOI21_X1 U8891 ( .B1(n7274), .B2(n7269), .A(n7268), .ZN(n7489) );
  AOI21_X1 U8892 ( .B1(n7531), .B2(n7339), .A(n9704), .ZN(n7270) );
  NAND2_X1 U8893 ( .A1(n7270), .A2(n7379), .ZN(n7488) );
  OAI21_X1 U8894 ( .B1(n7494), .B2(n9702), .A(n7488), .ZN(n7271) );
  AOI21_X1 U8895 ( .B1(n7489), .B2(n9708), .A(n7271), .ZN(n7276) );
  NAND2_X1 U8896 ( .A1(n7273), .A2(n7272), .ZN(n7330) );
  XOR2_X1 U8897 ( .A(n7274), .B(n7330), .Z(n7275) );
  AOI222_X1 U8898 ( .A1(n9501), .A2(n7275), .B1(n8982), .B2(n9306), .C1(n8984), 
        .C2(n9304), .ZN(n7487) );
  NAND2_X1 U8899 ( .A1(n7276), .A2(n7487), .ZN(n7279) );
  NAND2_X1 U8900 ( .A1(n7279), .A2(n9724), .ZN(n7277) );
  OAI21_X1 U8901 ( .B1(n9724), .B2(n7278), .A(n7277), .ZN(P1_U3469) );
  NAND2_X1 U8902 ( .A1(n7279), .A2(n9733), .ZN(n7280) );
  OAI21_X1 U8903 ( .B1(n9733), .B2(n6589), .A(n7280), .ZN(P1_U3528) );
  INV_X1 U8904 ( .A(n7281), .ZN(n7286) );
  AOI22_X1 U8905 ( .A1(n7283), .A2(n9827), .B1(n8804), .B2(n7282), .ZN(n7284)
         );
  OAI211_X1 U8906 ( .C1(n9905), .C2(n7286), .A(n7285), .B(n7284), .ZN(n7288)
         );
  NAND2_X1 U8907 ( .A1(n7288), .A2(n9934), .ZN(n7287) );
  OAI21_X1 U8908 ( .B1(n9934), .B2(n6384), .A(n7287), .ZN(P2_U3528) );
  INV_X1 U8909 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7290) );
  NAND2_X1 U8910 ( .A1(n7288), .A2(n9923), .ZN(n7289) );
  OAI21_X1 U8911 ( .B1(n9923), .B2(n7290), .A(n7289), .ZN(P2_U3475) );
  OAI222_X1 U8912 ( .A1(n7293), .A2(P1_U3084), .B1(n9539), .B2(n7292), .C1(
        n7291), .C2(n8242), .ZN(P1_U3332) );
  NAND2_X1 U8913 ( .A1(n7295), .A2(n7294), .ZN(n7296) );
  XOR2_X1 U8914 ( .A(n7297), .B(n7296), .Z(n7298) );
  NAND2_X1 U8915 ( .A1(n7298), .A2(n9643), .ZN(n7305) );
  OAI22_X1 U8916 ( .A1(n8964), .A2(n7299), .B1(n9697), .B2(n8959), .ZN(n7303)
         );
  INV_X1 U8917 ( .A(n8982), .ZN(n7323) );
  OAI21_X1 U8918 ( .B1(n7301), .B2(n7323), .A(n7300), .ZN(n7302) );
  NOR2_X1 U8919 ( .A1(n7303), .A2(n7302), .ZN(n7304) );
  OAI211_X1 U8920 ( .C1(n9648), .C2(n7333), .A(n7305), .B(n7304), .ZN(P1_U3211) );
  NAND2_X1 U8921 ( .A1(n7307), .A2(n7306), .ZN(n7309) );
  XNOR2_X1 U8922 ( .A(n7309), .B(n7308), .ZN(n7317) );
  INV_X1 U8923 ( .A(n9703), .ZN(n7600) );
  INV_X1 U8924 ( .A(n9633), .ZN(n8884) );
  NAND2_X1 U8925 ( .A1(n9306), .A2(n8979), .ZN(n7311) );
  NAND2_X1 U8926 ( .A1(n9304), .A2(n8981), .ZN(n7310) );
  AND2_X1 U8927 ( .A1(n7311), .A2(n7310), .ZN(n7398) );
  INV_X1 U8928 ( .A(n7312), .ZN(n7401) );
  NAND2_X1 U8929 ( .A1(n8930), .A2(n7401), .ZN(n7313) );
  OAI211_X1 U8930 ( .C1(n8884), .C2(n7398), .A(n7314), .B(n7313), .ZN(n7315)
         );
  AOI21_X1 U8931 ( .B1(n8970), .B2(n7600), .A(n7315), .ZN(n7316) );
  OAI21_X1 U8932 ( .B1(n7317), .B2(n8972), .A(n7316), .ZN(P1_U3219) );
  XNOR2_X1 U8933 ( .A(n7318), .B(n7319), .ZN(n7320) );
  NAND2_X1 U8934 ( .A1(n7320), .A2(n7321), .ZN(n9635) );
  OAI21_X1 U8935 ( .B1(n7321), .B2(n7320), .A(n9635), .ZN(n7322) );
  NAND2_X1 U8936 ( .A1(n7322), .A2(n9643), .ZN(n7327) );
  OAI22_X1 U8937 ( .A1(n8964), .A2(n7323), .B1(n7494), .B2(n8959), .ZN(n7324)
         );
  AOI211_X1 U8938 ( .C1(n8967), .C2(n8984), .A(n7325), .B(n7324), .ZN(n7326)
         );
  OAI211_X1 U8939 ( .C1(n9648), .C2(n7490), .A(n7327), .B(n7326), .ZN(P1_U3225) );
  INV_X1 U8940 ( .A(n7344), .ZN(n7393) );
  XNOR2_X1 U8941 ( .A(n7394), .B(n7393), .ZN(n7331) );
  AOI222_X1 U8942 ( .A1(n9501), .A2(n7331), .B1(n8980), .B2(n9306), .C1(n8982), 
        .C2(n9304), .ZN(n9696) );
  NAND2_X1 U8943 ( .A1(n9377), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7332) );
  OAI21_X1 U8944 ( .B1(n9559), .B2(n7333), .A(n7332), .ZN(n7338) );
  INV_X1 U8945 ( .A(n7380), .ZN(n7335) );
  INV_X1 U8946 ( .A(n7400), .ZN(n7334) );
  OAI211_X1 U8947 ( .C1(n9697), .C2(n7335), .A(n7334), .B(n9713), .ZN(n9695)
         );
  NOR2_X1 U8948 ( .A1(n9695), .A2(n7336), .ZN(n7337) );
  AOI211_X1 U8949 ( .C1(n9595), .C2(n7389), .A(n7338), .B(n7337), .ZN(n7349)
         );
  NAND2_X1 U8950 ( .A1(n8983), .A2(n7339), .ZN(n7340) );
  OR2_X1 U8951 ( .A1(n8982), .A2(n7384), .ZN(n7343) );
  NAND2_X1 U8952 ( .A1(n7374), .A2(n7343), .ZN(n7345) );
  OAI21_X1 U8953 ( .B1(n7345), .B2(n7344), .A(n7391), .ZN(n9699) );
  NAND2_X1 U8954 ( .A1(n8195), .A2(n7346), .ZN(n7347) );
  INV_X1 U8955 ( .A(n9392), .ZN(n9224) );
  NAND2_X1 U8956 ( .A1(n9699), .A2(n9224), .ZN(n7348) );
  OAI211_X1 U8957 ( .C1(n9696), .C2(n9605), .A(n7349), .B(n7348), .ZN(P1_U3284) );
  OR2_X1 U8958 ( .A1(n7350), .A2(n8443), .ZN(n7351) );
  NAND2_X1 U8959 ( .A1(n7569), .A2(n7558), .ZN(n8031) );
  NAND2_X1 U8960 ( .A1(n7354), .A2(n8154), .ZN(n7355) );
  OAI22_X1 U8961 ( .A1(n7356), .A2(n8664), .B1(n7555), .B2(n8662), .ZN(n7362)
         );
  AND2_X1 U8962 ( .A1(n8031), .A2(n8023), .ZN(n8029) );
  INV_X1 U8963 ( .A(n7556), .ZN(n7360) );
  AOI21_X1 U8964 ( .B1(n7358), .B2(n8023), .A(n8154), .ZN(n7359) );
  AOI211_X1 U8965 ( .C1(n7360), .C2(n8032), .A(n8605), .B(n7359), .ZN(n7361)
         );
  AOI211_X1 U8966 ( .C1(n7568), .C2(n7681), .A(n7362), .B(n7361), .ZN(n7572)
         );
  NAND2_X1 U8967 ( .A1(n7363), .A2(n7569), .ZN(n7364) );
  AND2_X1 U8968 ( .A1(n7559), .A2(n7364), .ZN(n7570) );
  NAND2_X1 U8969 ( .A1(n7570), .A2(n8716), .ZN(n7370) );
  INV_X1 U8970 ( .A(n7365), .ZN(n7367) );
  OAI22_X1 U8971 ( .A1(n9838), .A2(n6401), .B1(n7367), .B2(n7366), .ZN(n7368)
         );
  AOI21_X1 U8972 ( .B1(n7684), .B2(n7569), .A(n7368), .ZN(n7369) );
  NAND2_X1 U8973 ( .A1(n7370), .A2(n7369), .ZN(n7371) );
  AOI21_X1 U8974 ( .B1(n7568), .B2(n7689), .A(n7371), .ZN(n7372) );
  OAI21_X1 U8975 ( .B1(n7572), .B2(n8713), .A(n7372), .ZN(P2_U3286) );
  INV_X1 U8976 ( .A(n7856), .ZN(n8190) );
  OAI222_X1 U8977 ( .A1(P1_U3084), .A2(n5804), .B1(n8245), .B2(n8190), .C1(
        n7373), .C2(n8242), .ZN(P1_U3331) );
  OAI21_X1 U8978 ( .B1(n9605), .B2(n9497), .A(n9373), .ZN(n9400) );
  INV_X1 U8979 ( .A(n9400), .ZN(n7618) );
  OAI21_X1 U8980 ( .B1(n7375), .B2(n7342), .A(n7374), .ZN(n9693) );
  INV_X1 U8981 ( .A(n9693), .ZN(n7388) );
  XNOR2_X1 U8982 ( .A(n7377), .B(n7376), .ZN(n7378) );
  AOI22_X1 U8983 ( .A1(n9306), .A2(n8981), .B1(n9304), .B2(n8983), .ZN(n9631)
         );
  OAI21_X1 U8984 ( .B1(n7378), .B2(n9553), .A(n9631), .ZN(n9691) );
  INV_X1 U8985 ( .A(n7379), .ZN(n7381) );
  OAI21_X1 U8986 ( .B1(n7381), .B2(n9641), .A(n7380), .ZN(n9690) );
  OAI22_X1 U8987 ( .A1(n9327), .A2(n7382), .B1(n9647), .B2(n9559), .ZN(n7383)
         );
  AOI21_X1 U8988 ( .B1(n9595), .B2(n7384), .A(n7383), .ZN(n7385) );
  OAI21_X1 U8989 ( .B1(n9690), .B2(n9389), .A(n7385), .ZN(n7386) );
  AOI21_X1 U8990 ( .B1(n9691), .B2(n9327), .A(n7386), .ZN(n7387) );
  OAI21_X1 U8991 ( .B1(n7618), .B2(n7388), .A(n7387), .ZN(P1_U3285) );
  OR2_X1 U8992 ( .A1(n8981), .A2(n7389), .ZN(n7390) );
  OAI21_X1 U8993 ( .B1(n7392), .B2(n7397), .A(n7601), .ZN(n9701) );
  NAND2_X1 U8994 ( .A1(n7394), .A2(n7393), .ZN(n7396) );
  NAND2_X1 U8995 ( .A1(n7396), .A2(n7395), .ZN(n7602) );
  XNOR2_X1 U8996 ( .A(n7602), .B(n7397), .ZN(n7399) );
  OAI21_X1 U8997 ( .B1(n7399), .B2(n9553), .A(n7398), .ZN(n9707) );
  OAI21_X1 U8998 ( .B1(n7400), .B2(n9703), .A(n7610), .ZN(n9705) );
  AOI22_X1 U8999 ( .A1(n9605), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7401), .B2(
        n9594), .ZN(n7403) );
  NAND2_X1 U9000 ( .A1(n9595), .A2(n7600), .ZN(n7402) );
  OAI211_X1 U9001 ( .C1(n9705), .C2(n9389), .A(n7403), .B(n7402), .ZN(n7404)
         );
  AOI21_X1 U9002 ( .B1(n9707), .B2(n9327), .A(n7404), .ZN(n7405) );
  OAI21_X1 U9003 ( .B1(n9701), .B2(n7618), .A(n7405), .ZN(P1_U3283) );
  INV_X1 U9004 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7407) );
  AND2_X1 U9005 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8966) );
  INV_X1 U9006 ( .A(n8966), .ZN(n7406) );
  OAI21_X1 U9007 ( .B1(n10167), .B2(n7407), .A(n7406), .ZN(n7413) );
  NOR2_X1 U9008 ( .A1(n7408), .A2(n7415), .ZN(n7410) );
  NOR2_X1 U9009 ( .A1(n7410), .A2(n7409), .ZN(n7588) );
  XNOR2_X1 U9010 ( .A(n7588), .B(n7587), .ZN(n7411) );
  NOR2_X1 U9011 ( .A1(n5202), .A2(n7411), .ZN(n7589) );
  AOI211_X1 U9012 ( .C1(n7411), .C2(n5202), .A(n7589), .B(n10154), .ZN(n7412)
         );
  AOI211_X1 U9013 ( .C1(n9036), .C2(n7579), .A(n7413), .B(n7412), .ZN(n7418)
         );
  XNOR2_X1 U9014 ( .A(n7578), .B(n7587), .ZN(n7416) );
  NAND2_X1 U9015 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7416), .ZN(n7580) );
  OAI211_X1 U9016 ( .C1(n7416), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9660), .B(
        n7580), .ZN(n7417) );
  NAND2_X1 U9017 ( .A1(n7418), .A2(n7417), .ZN(P1_U3256) );
  INV_X1 U9018 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10179) );
  NOR2_X1 U9019 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7419) );
  AOI21_X1 U9020 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7419), .ZN(n9941) );
  NOR2_X1 U9021 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7420) );
  AOI21_X1 U9022 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7420), .ZN(n9944) );
  NOR2_X1 U9023 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7421) );
  AOI21_X1 U9024 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7421), .ZN(n9947) );
  NOR2_X1 U9025 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7422) );
  AOI21_X1 U9026 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7422), .ZN(n9950) );
  NOR2_X1 U9027 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7423) );
  AOI21_X1 U9028 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7423), .ZN(n9953) );
  NOR2_X1 U9029 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7432) );
  INV_X1 U9030 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7424) );
  XOR2_X1 U9031 ( .A(n7424), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10192) );
  NAND2_X1 U9032 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7430) );
  INV_X1 U9033 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7425) );
  XNOR2_X1 U9034 ( .A(n7425), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U9035 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7428) );
  XNOR2_X1 U9036 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n7426), .ZN(n10188) );
  AOI21_X1 U9037 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9935) );
  NAND3_X1 U9038 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9937) );
  OAI21_X1 U9039 ( .B1(n9935), .B2(n6452), .A(n9937), .ZN(n10187) );
  NAND2_X1 U9040 ( .A1(n10188), .A2(n10187), .ZN(n7427) );
  NAND2_X1 U9041 ( .A1(n7428), .A2(n7427), .ZN(n10189) );
  NAND2_X1 U9042 ( .A1(n10190), .A2(n10189), .ZN(n7429) );
  NAND2_X1 U9043 ( .A1(n7430), .A2(n7429), .ZN(n10191) );
  NOR2_X1 U9044 ( .A1(n10192), .A2(n10191), .ZN(n7431) );
  NOR2_X1 U9045 ( .A1(n7432), .A2(n7431), .ZN(n7433) );
  NOR2_X1 U9046 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7433), .ZN(n10174) );
  AND2_X1 U9047 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7433), .ZN(n10175) );
  NOR2_X1 U9048 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10175), .ZN(n7434) );
  NOR2_X1 U9049 ( .A1(n10174), .A2(n7434), .ZN(n7435) );
  NAND2_X1 U9050 ( .A1(n7435), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7437) );
  XOR2_X1 U9051 ( .A(n7435), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10173) );
  NAND2_X1 U9052 ( .A1(n10173), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7436) );
  NAND2_X1 U9053 ( .A1(n7437), .A2(n7436), .ZN(n7438) );
  NAND2_X1 U9054 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7438), .ZN(n7440) );
  XNOR2_X1 U9055 ( .A(n10077), .B(n7438), .ZN(n10186) );
  NAND2_X1 U9056 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10186), .ZN(n7439) );
  NAND2_X1 U9057 ( .A1(n7440), .A2(n7439), .ZN(n7441) );
  NAND2_X1 U9058 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7441), .ZN(n7443) );
  XOR2_X1 U9059 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7441), .Z(n10185) );
  NAND2_X1 U9060 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10185), .ZN(n7442) );
  NAND2_X1 U9061 ( .A1(n7443), .A2(n7442), .ZN(n7444) );
  AND2_X1 U9062 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7444), .ZN(n7445) );
  INV_X1 U9063 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10184) );
  XNOR2_X1 U9064 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7444), .ZN(n10183) );
  NOR2_X1 U9065 ( .A1(n10184), .A2(n10183), .ZN(n10182) );
  NAND2_X1 U9066 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7446) );
  OAI21_X1 U9067 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n7446), .ZN(n9961) );
  AOI21_X1 U9068 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9960), .ZN(n9959) );
  NAND2_X1 U9069 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7447) );
  OAI21_X1 U9070 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7447), .ZN(n9958) );
  NOR2_X1 U9071 ( .A1(n9959), .A2(n9958), .ZN(n9957) );
  AOI21_X1 U9072 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9957), .ZN(n9956) );
  NOR2_X1 U9073 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7448) );
  AOI21_X1 U9074 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7448), .ZN(n9955) );
  NAND2_X1 U9075 ( .A1(n9956), .A2(n9955), .ZN(n9954) );
  OAI21_X1 U9076 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9954), .ZN(n9952) );
  NAND2_X1 U9077 ( .A1(n9953), .A2(n9952), .ZN(n9951) );
  OAI21_X1 U9078 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9951), .ZN(n9949) );
  NAND2_X1 U9079 ( .A1(n9950), .A2(n9949), .ZN(n9948) );
  OAI21_X1 U9080 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9948), .ZN(n9946) );
  NAND2_X1 U9081 ( .A1(n9947), .A2(n9946), .ZN(n9945) );
  OAI21_X1 U9082 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9945), .ZN(n9943) );
  NAND2_X1 U9083 ( .A1(n9944), .A2(n9943), .ZN(n9942) );
  OAI21_X1 U9084 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9942), .ZN(n9940) );
  NAND2_X1 U9085 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  OAI21_X1 U9086 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9939), .ZN(n10178) );
  NOR2_X1 U9087 ( .A1(n10179), .A2(n10178), .ZN(n7449) );
  NAND2_X1 U9088 ( .A1(n10179), .A2(n10178), .ZN(n10177) );
  OAI21_X1 U9089 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7449), .A(n10177), .ZN(
        n7451) );
  XNOR2_X1 U9090 ( .A(n4809), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7450) );
  XNOR2_X1 U9091 ( .A(n7451), .B(n7450), .ZN(ADD_1071_U4) );
  INV_X1 U9092 ( .A(n7867), .ZN(n7453) );
  NAND2_X1 U9093 ( .A1(n8828), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7452) );
  OAI211_X1 U9094 ( .C1(n7453), .C2(n8830), .A(n8183), .B(n7452), .ZN(P2_U3335) );
  NAND2_X1 U9095 ( .A1(n7454), .A2(n7969), .ZN(n7458) );
  OAI22_X1 U9096 ( .A1(n6907), .A2(n10117), .B1(n7832), .B2(n7455), .ZN(n7456)
         );
  INV_X1 U9097 ( .A(n7456), .ZN(n7457) );
  XNOR2_X1 U9098 ( .A(n7718), .B(n8300), .ZN(n7459) );
  NAND2_X1 U9099 ( .A1(n8440), .A2(n8301), .ZN(n7460) );
  NAND2_X1 U9100 ( .A1(n7459), .A2(n7460), .ZN(n7502) );
  INV_X1 U9101 ( .A(n7459), .ZN(n7462) );
  INV_X1 U9102 ( .A(n7460), .ZN(n7461) );
  NAND2_X1 U9103 ( .A1(n7462), .A2(n7461), .ZN(n7463) );
  NAND2_X1 U9104 ( .A1(n7502), .A2(n7463), .ZN(n7475) );
  INV_X1 U9105 ( .A(n7466), .ZN(n7467) );
  NAND2_X1 U9106 ( .A1(n7468), .A2(n7467), .ZN(n7469) );
  NAND2_X1 U9107 ( .A1(n7470), .A2(n7469), .ZN(n7471) );
  INV_X1 U9108 ( .A(n7471), .ZN(n7473) );
  INV_X1 U9109 ( .A(n7475), .ZN(n7472) );
  INV_X1 U9110 ( .A(n7503), .ZN(n7474) );
  AOI21_X1 U9111 ( .B1(n7475), .B2(n7471), .A(n7474), .ZN(n7486) );
  NAND2_X1 U9112 ( .A1(n7882), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7481) );
  NAND2_X1 U9113 ( .A1(n7957), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7480) );
  NAND2_X1 U9114 ( .A1(n7476), .A2(n10135), .ZN(n7477) );
  AND2_X1 U9115 ( .A1(n7510), .A2(n7477), .ZN(n7685) );
  NAND2_X1 U9116 ( .A1(n7937), .A2(n7685), .ZN(n7479) );
  NAND2_X1 U9117 ( .A1(n7958), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7478) );
  NAND4_X1 U9118 ( .A1(n7481), .A2(n7480), .A3(n7479), .A4(n7478), .ZN(n8711)
         );
  INV_X1 U9119 ( .A(n8711), .ZN(n7700) );
  AOI22_X1 U9120 ( .A1(n8376), .A2(n8441), .B1(n7760), .B2(n8433), .ZN(n7483)
         );
  OAI211_X1 U9121 ( .C1(n7700), .C2(n8415), .A(n7483), .B(n7482), .ZN(n7484)
         );
  AOI21_X1 U9122 ( .B1(n7718), .B2(n8421), .A(n7484), .ZN(n7485) );
  OAI21_X1 U9123 ( .B1(n7486), .B2(n8423), .A(n7485), .ZN(P2_U3226) );
  OAI21_X1 U9124 ( .B1(n9061), .B2(n7488), .A(n7487), .ZN(n7496) );
  NAND2_X1 U9125 ( .A1(n7489), .A2(n9224), .ZN(n7493) );
  INV_X1 U9126 ( .A(n7490), .ZN(n7491) );
  AOI22_X1 U9127 ( .A1(n9605), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7491), .B2(
        n9594), .ZN(n7492) );
  OAI211_X1 U9128 ( .C1(n7494), .C2(n9401), .A(n7493), .B(n7492), .ZN(n7495)
         );
  AOI21_X1 U9129 ( .B1(n7496), .B2(n9327), .A(n7495), .ZN(n7497) );
  INV_X1 U9130 ( .A(n7497), .ZN(P1_U3286) );
  NAND2_X1 U9131 ( .A1(n7867), .A2(n7498), .ZN(n7500) );
  OAI211_X1 U9132 ( .C1(n7501), .C2(n8242), .A(n7500), .B(n7499), .ZN(P1_U3330) );
  NAND2_X1 U9133 ( .A1(n7504), .A2(n7969), .ZN(n7508) );
  OAI22_X1 U9134 ( .A1(n6907), .A2(n9967), .B1(n7505), .B2(n7832), .ZN(n7506)
         );
  INV_X1 U9135 ( .A(n7506), .ZN(n7507) );
  XNOR2_X1 U9136 ( .A(n8803), .B(n8300), .ZN(n7634) );
  NAND2_X1 U9137 ( .A1(n8711), .A2(n8301), .ZN(n7635) );
  XNOR2_X1 U9138 ( .A(n7634), .B(n7635), .ZN(n7623) );
  XNOR2_X1 U9139 ( .A(n7624), .B(n7623), .ZN(n7520) );
  NAND2_X1 U9140 ( .A1(n7882), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7515) );
  NAND2_X1 U9141 ( .A1(n7957), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7514) );
  NAND2_X1 U9142 ( .A1(n7510), .A2(n7509), .ZN(n7511) );
  AND2_X1 U9143 ( .A1(n7645), .A2(n7511), .ZN(n8702) );
  NAND2_X1 U9144 ( .A1(n7937), .A2(n8702), .ZN(n7513) );
  NAND2_X1 U9145 ( .A1(n7958), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7512) );
  NAND4_X1 U9146 ( .A1(n7515), .A2(n7514), .A3(n7513), .A4(n7512), .ZN(n8692)
         );
  OAI22_X1 U9147 ( .A1(n8415), .A2(n7800), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10135), .ZN(n7518) );
  INV_X1 U9148 ( .A(n7685), .ZN(n7516) );
  OAI22_X1 U9149 ( .A1(n8418), .A2(n7678), .B1(n7516), .B2(n8416), .ZN(n7517)
         );
  AOI211_X1 U9150 ( .C1(n8803), .C2(n8421), .A(n7518), .B(n7517), .ZN(n7519)
         );
  OAI21_X1 U9151 ( .B1(n7520), .B2(n8423), .A(n7519), .ZN(P2_U3236) );
  OAI21_X1 U9152 ( .B1(n7522), .B2(n7523), .A(n7521), .ZN(n7528) );
  INV_X1 U9153 ( .A(n7528), .ZN(n9686) );
  XNOR2_X1 U9154 ( .A(n7524), .B(n7523), .ZN(n7526) );
  AOI22_X1 U9155 ( .A1(n9306), .A2(n8983), .B1(n9304), .B2(n8985), .ZN(n7525)
         );
  OAI21_X1 U9156 ( .B1(n7526), .B2(n9553), .A(n7525), .ZN(n7527) );
  AOI21_X1 U9157 ( .B1(n7528), .B2(n9721), .A(n7527), .ZN(n9685) );
  MUX2_X1 U9158 ( .A(n7529), .B(n9685), .S(n9327), .Z(n7538) );
  INV_X1 U9159 ( .A(n7530), .ZN(n7533) );
  INV_X1 U9160 ( .A(n7531), .ZN(n7532) );
  AOI21_X1 U9161 ( .B1(n9682), .B2(n7533), .A(n7532), .ZN(n9683) );
  OAI22_X1 U9162 ( .A1(n9401), .A2(n7535), .B1(n7534), .B2(n9559), .ZN(n7536)
         );
  AOI21_X1 U9163 ( .B1(n9566), .B2(n9683), .A(n7536), .ZN(n7537) );
  OAI211_X1 U9164 ( .C1(n9686), .C2(n9373), .A(n7538), .B(n7537), .ZN(P1_U3287) );
  INV_X1 U9165 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10141) );
  XNOR2_X1 U9166 ( .A(n9800), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U9167 ( .A1(n7540), .A2(n7539), .ZN(n9799) );
  NAND2_X1 U9168 ( .A1(n9798), .A2(n9799), .ZN(n9796) );
  OAI21_X1 U9169 ( .B1(n10141), .B2(n9800), .A(n9796), .ZN(n8463) );
  XOR2_X1 U9170 ( .A(n8463), .B(n8470), .Z(n7541) );
  NOR2_X1 U9171 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n7541), .ZN(n8466) );
  AOI21_X1 U9172 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n7541), .A(n8466), .ZN(
        n7553) );
  NAND2_X1 U9173 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3152), .ZN(n7542) );
  OAI21_X1 U9174 ( .B1(n8484), .B2(n10179), .A(n7542), .ZN(n7551) );
  INV_X1 U9175 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7546) );
  XNOR2_X1 U9176 ( .A(n9800), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9805) );
  NOR2_X1 U9177 ( .A1(n7543), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7544) );
  NOR2_X1 U9178 ( .A1(n7545), .A2(n7544), .ZN(n9806) );
  NAND2_X1 U9179 ( .A1(n9805), .A2(n9806), .ZN(n9803) );
  OAI21_X1 U9180 ( .B1(n7546), .B2(n9800), .A(n9803), .ZN(n7548) );
  INV_X1 U9181 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8469) );
  AOI22_X1 U9182 ( .A1(n8464), .A2(n8469), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8470), .ZN(n7547) );
  NOR2_X1 U9183 ( .A1(n7548), .A2(n7547), .ZN(n8468) );
  AOI21_X1 U9184 ( .B1(n7548), .B2(n7547), .A(n8468), .ZN(n7549) );
  NOR2_X1 U9185 ( .A1(n7549), .A2(n8475), .ZN(n7550) );
  AOI211_X1 U9186 ( .C1(n9802), .C2(n8464), .A(n7551), .B(n7550), .ZN(n7552)
         );
  OAI21_X1 U9187 ( .B1(n7553), .B2(n9736), .A(n7552), .ZN(P2_U3263) );
  NAND2_X1 U9188 ( .A1(n8041), .A2(n7555), .ZN(n8025) );
  NAND2_X1 U9189 ( .A1(n8033), .A2(n8025), .ZN(n8156) );
  XOR2_X1 U9190 ( .A(n7665), .B(n8156), .Z(n9920) );
  INV_X1 U9191 ( .A(n9920), .ZN(n7567) );
  XOR2_X1 U9192 ( .A(n8156), .B(n7672), .Z(n7557) );
  OAI222_X1 U9193 ( .A1(n8662), .A2(n7678), .B1(n8664), .B2(n7558), .C1(n8605), 
        .C2(n7557), .ZN(n9917) );
  INV_X1 U9194 ( .A(n7559), .ZN(n7560) );
  OAI21_X1 U9195 ( .B1(n4590), .B2(n7560), .A(n4395), .ZN(n9916) );
  AOI22_X1 U9196 ( .A1(n8713), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7561), .B2(
        n9834), .ZN(n7563) );
  NAND2_X1 U9197 ( .A1(n7684), .A2(n8041), .ZN(n7562) );
  OAI211_X1 U9198 ( .C1(n9916), .C2(n7564), .A(n7563), .B(n7562), .ZN(n7565)
         );
  AOI21_X1 U9199 ( .B1(n9917), .B2(n9838), .A(n7565), .ZN(n7566) );
  OAI21_X1 U9200 ( .B1(n7567), .B2(n8718), .A(n7566), .ZN(P2_U3285) );
  INV_X1 U9201 ( .A(n7568), .ZN(n7573) );
  AOI22_X1 U9202 ( .A1(n7570), .A2(n9827), .B1(n8804), .B2(n7569), .ZN(n7571)
         );
  OAI211_X1 U9203 ( .C1(n9905), .C2(n7573), .A(n7572), .B(n7571), .ZN(n7575)
         );
  NAND2_X1 U9204 ( .A1(n7575), .A2(n9934), .ZN(n7574) );
  OAI21_X1 U9205 ( .B1(n9934), .B2(n6394), .A(n7574), .ZN(P2_U3530) );
  INV_X1 U9206 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7577) );
  NAND2_X1 U9207 ( .A1(n7575), .A2(n9923), .ZN(n7576) );
  OAI21_X1 U9208 ( .B1(n9923), .B2(n7577), .A(n7576), .ZN(P2_U3481) );
  NAND2_X1 U9209 ( .A1(n7579), .A2(n7578), .ZN(n7581) );
  XNOR2_X1 U9210 ( .A(n7592), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9017) );
  INV_X1 U9211 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7583) );
  XNOR2_X1 U9212 ( .A(n9031), .B(n7583), .ZN(n9032) );
  XNOR2_X1 U9213 ( .A(n9033), .B(n9032), .ZN(n7599) );
  NOR2_X1 U9214 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5169), .ZN(n7586) );
  INV_X1 U9215 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7584) );
  NOR2_X1 U9216 ( .A1(n10167), .A2(n7584), .ZN(n7585) );
  AOI211_X1 U9217 ( .C1(n9036), .C2(n9031), .A(n7586), .B(n7585), .ZN(n7598)
         );
  NOR2_X1 U9218 ( .A1(n7588), .A2(n7587), .ZN(n7590) );
  NOR2_X1 U9219 ( .A1(n7590), .A2(n7589), .ZN(n9022) );
  MUX2_X1 U9220 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n7591), .S(n9023), .Z(n9021)
         );
  NAND2_X1 U9221 ( .A1(n7592), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9222 ( .A1(n9019), .A2(n7593), .ZN(n7596) );
  OR2_X1 U9223 ( .A1(n9031), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7594) );
  NAND2_X1 U9224 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9031), .ZN(n9041) );
  AND2_X1 U9225 ( .A1(n7594), .A2(n9041), .ZN(n7595) );
  NAND2_X1 U9226 ( .A1(n7596), .A2(n7595), .ZN(n9042) );
  OAI211_X1 U9227 ( .C1(n7596), .C2(n7595), .A(n9042), .B(n9651), .ZN(n7597)
         );
  OAI211_X1 U9228 ( .C1(n7599), .C2(n10162), .A(n7598), .B(n7597), .ZN(
        P1_U3258) );
  XNOR2_X1 U9229 ( .A(n7736), .B(n7607), .ZN(n9717) );
  INV_X1 U9230 ( .A(n7602), .ZN(n7606) );
  XOR2_X1 U9231 ( .A(n7738), .B(n7607), .Z(n7608) );
  INV_X1 U9232 ( .A(n7746), .ZN(n8978) );
  AOI222_X1 U9233 ( .A1(n9501), .A2(n7608), .B1(n8978), .B2(n9306), .C1(n8980), 
        .C2(n9304), .ZN(n9716) );
  INV_X1 U9234 ( .A(n9716), .ZN(n7616) );
  INV_X1 U9235 ( .A(n7609), .ZN(n9564) );
  AOI21_X1 U9236 ( .B1(n9711), .B2(n7610), .A(n9564), .ZN(n9714) );
  NAND2_X1 U9237 ( .A1(n9714), .A2(n9566), .ZN(n7614) );
  INV_X1 U9238 ( .A(n7611), .ZN(n7612) );
  AOI22_X1 U9239 ( .A1(n9605), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7612), .B2(
        n9594), .ZN(n7613) );
  OAI211_X1 U9240 ( .C1(n7730), .C2(n9401), .A(n7614), .B(n7613), .ZN(n7615)
         );
  AOI21_X1 U9241 ( .B1(n7616), .B2(n9327), .A(n7615), .ZN(n7617) );
  OAI21_X1 U9242 ( .B1(n7618), .B2(n9717), .A(n7617), .ZN(P1_U3282) );
  INV_X1 U9243 ( .A(n7879), .ZN(n7620) );
  OAI222_X1 U9244 ( .A1(n5787), .A2(P1_U3084), .B1(n9539), .B2(n7620), .C1(
        n7619), .C2(n8242), .ZN(P1_U3329) );
  OAI222_X1 U9245 ( .A1(P2_U3152), .A2(n7622), .B1(n8831), .B2(n7621), .C1(
        n8830), .C2(n7620), .ZN(P2_U3334) );
  NAND2_X1 U9246 ( .A1(n7625), .A2(n7969), .ZN(n7628) );
  AOI22_X1 U9247 ( .A1(n7970), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7641), .B2(
        n7626), .ZN(n7627) );
  XNOR2_X1 U9248 ( .A(n8797), .B(n8300), .ZN(n7629) );
  NAND2_X1 U9249 ( .A1(n8692), .A2(n8301), .ZN(n7630) );
  NAND2_X1 U9250 ( .A1(n7629), .A2(n7630), .ZN(n7639) );
  INV_X1 U9251 ( .A(n7629), .ZN(n7632) );
  INV_X1 U9252 ( .A(n7630), .ZN(n7631) );
  NAND2_X1 U9253 ( .A1(n7632), .A2(n7631), .ZN(n7633) );
  AND2_X1 U9254 ( .A1(n7639), .A2(n7633), .ZN(n7696) );
  INV_X1 U9255 ( .A(n7634), .ZN(n7637) );
  INV_X1 U9256 ( .A(n7635), .ZN(n7636) );
  NAND2_X1 U9257 ( .A1(n7637), .A2(n7636), .ZN(n7692) );
  AND2_X1 U9258 ( .A1(n7696), .A2(n7692), .ZN(n7638) );
  NAND2_X1 U9259 ( .A1(n7640), .A2(n7969), .ZN(n7644) );
  AOI22_X1 U9260 ( .A1(n7642), .A2(n7641), .B1(n7970), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n7643) );
  XNOR2_X1 U9261 ( .A(n8792), .B(n8300), .ZN(n8246) );
  INV_X1 U9262 ( .A(n8246), .ZN(n8249) );
  NAND2_X1 U9263 ( .A1(n7957), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7650) );
  NAND2_X1 U9264 ( .A1(n7882), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U9265 ( .A1(n7645), .A2(n7659), .ZN(n7646) );
  AND2_X1 U9266 ( .A1(n7653), .A2(n7646), .ZN(n8689) );
  NAND2_X1 U9267 ( .A1(n7937), .A2(n8689), .ZN(n7648) );
  NAND2_X1 U9268 ( .A1(n7958), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7647) );
  NAND4_X1 U9269 ( .A1(n7650), .A2(n7649), .A3(n7648), .A4(n7647), .ZN(n8710)
         );
  AND2_X1 U9270 ( .A1(n8710), .A2(n8301), .ZN(n8247) );
  XNOR2_X1 U9271 ( .A(n8249), .B(n8247), .ZN(n7651) );
  XNOR2_X1 U9272 ( .A(n8248), .B(n7651), .ZN(n7664) );
  NAND2_X1 U9273 ( .A1(n7882), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U9274 ( .A1(n7957), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7657) );
  INV_X1 U9275 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7652) );
  NAND2_X1 U9276 ( .A1(n7653), .A2(n7652), .ZN(n7654) );
  AND2_X1 U9277 ( .A1(n7814), .A2(n7654), .ZN(n8675) );
  NAND2_X1 U9278 ( .A1(n7937), .A2(n8675), .ZN(n7656) );
  NAND2_X1 U9279 ( .A1(n7958), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7655) );
  NAND4_X1 U9280 ( .A1(n7658), .A2(n7657), .A3(n7656), .A4(n7655), .ZN(n8693)
         );
  INV_X1 U9281 ( .A(n8693), .ZN(n8059) );
  OAI22_X1 U9282 ( .A1(n8415), .A2(n8059), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7659), .ZN(n7662) );
  INV_X1 U9283 ( .A(n8689), .ZN(n7660) );
  OAI22_X1 U9284 ( .A1(n8418), .A2(n7800), .B1(n8416), .B2(n7660), .ZN(n7661)
         );
  AOI211_X1 U9285 ( .C1(n8792), .C2(n8421), .A(n7662), .B(n7661), .ZN(n7663)
         );
  OAI21_X1 U9286 ( .B1(n7664), .B2(n8423), .A(n7663), .ZN(P2_U3243) );
  NAND2_X1 U9287 ( .A1(n8041), .A2(n8441), .ZN(n7666) );
  NAND2_X1 U9288 ( .A1(n7667), .A2(n7666), .ZN(n7714) );
  NAND2_X1 U9289 ( .A1(n7718), .A2(n7678), .ZN(n7987) );
  OR2_X1 U9290 ( .A1(n7718), .A2(n8440), .ZN(n7668) );
  OR2_X1 U9291 ( .A1(n8803), .A2(n7700), .ZN(n8048) );
  NAND2_X1 U9292 ( .A1(n8803), .A2(n7700), .ZN(n8706) );
  NAND2_X1 U9293 ( .A1(n7670), .A2(n8045), .ZN(n7671) );
  INV_X1 U9294 ( .A(n7676), .ZN(n7673) );
  INV_X1 U9295 ( .A(n8040), .ZN(n7674) );
  OAI21_X1 U9296 ( .B1(n7673), .B2(n7674), .A(n7669), .ZN(n7677) );
  NOR2_X1 U9297 ( .A1(n7669), .A2(n7674), .ZN(n7675) );
  AOI21_X1 U9298 ( .B1(n7677), .B2(n8707), .A(n8605), .ZN(n7680) );
  OAI22_X1 U9299 ( .A1(n7678), .A2(n8664), .B1(n7800), .B2(n8662), .ZN(n7679)
         );
  AOI211_X1 U9300 ( .C1(n8802), .C2(n7681), .A(n7680), .B(n7679), .ZN(n8807)
         );
  INV_X1 U9301 ( .A(n7718), .ZN(n7762) );
  INV_X1 U9302 ( .A(n8803), .ZN(n7682) );
  NAND2_X1 U9303 ( .A1(n7717), .A2(n7682), .ZN(n8701) );
  OR2_X1 U9304 ( .A1(n7717), .A2(n7682), .ZN(n7683) );
  AND2_X1 U9305 ( .A1(n8701), .A2(n7683), .ZN(n8805) );
  NAND2_X1 U9306 ( .A1(n8803), .A2(n7684), .ZN(n7687) );
  NAND2_X1 U9307 ( .A1(n9834), .A2(n7685), .ZN(n7686) );
  OAI211_X1 U9308 ( .C1(n9838), .C2(n6422), .A(n7687), .B(n7686), .ZN(n7688)
         );
  AOI21_X1 U9309 ( .B1(n8805), .B2(n8716), .A(n7688), .ZN(n7691) );
  NAND2_X1 U9310 ( .A1(n8802), .A2(n7689), .ZN(n7690) );
  OAI211_X1 U9311 ( .C1(n8807), .C2(n8713), .A(n7691), .B(n7690), .ZN(P2_U3283) );
  INV_X1 U9312 ( .A(n8797), .ZN(n8705) );
  AND2_X1 U9313 ( .A1(n7693), .A2(n7692), .ZN(n7695) );
  OAI21_X1 U9314 ( .B1(n7696), .B2(n7695), .A(n7694), .ZN(n7697) );
  NAND2_X1 U9315 ( .A1(n7697), .A2(n8425), .ZN(n7704) );
  INV_X1 U9316 ( .A(n7698), .ZN(n7702) );
  INV_X1 U9317 ( .A(n8702), .ZN(n7699) );
  OAI22_X1 U9318 ( .A1(n8418), .A2(n7700), .B1(n7699), .B2(n8416), .ZN(n7701)
         );
  AOI211_X1 U9319 ( .C1(n8325), .C2(n8710), .A(n7702), .B(n7701), .ZN(n7703)
         );
  OAI211_X1 U9320 ( .C1(n8705), .C2(n8436), .A(n7704), .B(n7703), .ZN(P2_U3217) );
  INV_X1 U9321 ( .A(n7705), .ZN(n7707) );
  NOR2_X1 U9322 ( .A1(n7707), .A2(n7706), .ZN(n7708) );
  XNOR2_X1 U9323 ( .A(n7709), .B(n7708), .ZN(n7713) );
  OAI22_X1 U9324 ( .A1(n9552), .A2(n8977), .B1(n9364), .B2(n9556), .ZN(n9396)
         );
  AOI22_X1 U9325 ( .A1(n9633), .A2(n9396), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3084), .ZN(n7710) );
  OAI21_X1 U9326 ( .B1(n9403), .B2(n9648), .A(n7710), .ZN(n7711) );
  AOI21_X1 U9327 ( .B1(n8970), .B2(n9612), .A(n7711), .ZN(n7712) );
  OAI21_X1 U9328 ( .B1(n7713), .B2(n8972), .A(n7712), .ZN(P1_U3232) );
  INV_X2 U9329 ( .A(n9931), .ZN(n9934) );
  INV_X1 U9330 ( .A(n8042), .ZN(n8157) );
  XNOR2_X1 U9331 ( .A(n7714), .B(n8157), .ZN(n7768) );
  XNOR2_X1 U9332 ( .A(n7715), .B(n8157), .ZN(n7716) );
  AOI222_X1 U9333 ( .A1(n9816), .A2(n7716), .B1(n8711), .B2(n9818), .C1(n8441), 
        .C2(n9821), .ZN(n7763) );
  AOI21_X1 U9334 ( .B1(n7718), .B2(n4395), .A(n7717), .ZN(n7766) );
  AOI22_X1 U9335 ( .A1(n7766), .A2(n9827), .B1(n8804), .B2(n7718), .ZN(n7719)
         );
  OAI211_X1 U9336 ( .C1(n7768), .C2(n9877), .A(n7763), .B(n7719), .ZN(n7721)
         );
  NAND2_X1 U9337 ( .A1(n7721), .A2(n9934), .ZN(n7720) );
  OAI21_X1 U9338 ( .B1(n9934), .B2(n10119), .A(n7720), .ZN(P2_U3532) );
  INV_X1 U9339 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U9340 ( .A1(n7721), .A2(n9923), .ZN(n7722) );
  OAI21_X1 U9341 ( .B1(n9923), .B2(n7723), .A(n7722), .ZN(P2_U3487) );
  INV_X1 U9342 ( .A(n7892), .ZN(n7727) );
  OAI222_X1 U9343 ( .A1(P1_U3084), .A2(n7725), .B1(n8245), .B2(n7727), .C1(
        n7724), .C2(n8242), .ZN(P1_U3328) );
  OAI222_X1 U9344 ( .A1(n7728), .A2(P2_U3152), .B1(n8830), .B2(n7727), .C1(
        n7726), .C2(n8831), .ZN(P2_U3333) );
  AND2_X1 U9345 ( .A1(n9711), .A2(n8979), .ZN(n9543) );
  INV_X1 U9346 ( .A(n7731), .ZN(n7729) );
  NOR2_X1 U9347 ( .A1(n7729), .A2(n9549), .ZN(n7733) );
  OR2_X1 U9348 ( .A1(n9543), .A2(n7733), .ZN(n7735) );
  NAND2_X1 U9349 ( .A1(n9551), .A2(n7730), .ZN(n9544) );
  AND2_X1 U9350 ( .A1(n9544), .A2(n7731), .ZN(n7732) );
  OR2_X1 U9351 ( .A1(n7733), .A2(n7732), .ZN(n7734) );
  OAI21_X1 U9352 ( .B1(n7736), .B2(n7735), .A(n7734), .ZN(n9076) );
  XNOR2_X1 U9353 ( .A(n9076), .B(n7742), .ZN(n9510) );
  INV_X1 U9354 ( .A(n9493), .ZN(n7745) );
  NAND3_X1 U9355 ( .A1(n7743), .A2(n7742), .A3(n7741), .ZN(n7744) );
  OAI211_X1 U9356 ( .C1(n9494), .C2(n7745), .A(n7744), .B(n9501), .ZN(n7749)
         );
  OAI22_X1 U9357 ( .A1(n9552), .A2(n7746), .B1(n8977), .B2(n9556), .ZN(n7747)
         );
  INV_X1 U9358 ( .A(n7747), .ZN(n7748) );
  NAND2_X1 U9359 ( .A1(n7749), .A2(n7748), .ZN(n7750) );
  AOI21_X1 U9360 ( .B1(n9510), .B2(n9721), .A(n7750), .ZN(n9512) );
  INV_X1 U9361 ( .A(n9373), .ZN(n9600) );
  NOR2_X1 U9362 ( .A1(n9562), .A2(n9507), .ZN(n7751) );
  OR2_X1 U9363 ( .A1(n9502), .A2(n7751), .ZN(n9508) );
  INV_X1 U9364 ( .A(n7752), .ZN(n7753) );
  AOI22_X1 U9365 ( .A1(n9605), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7753), .B2(
        n9594), .ZN(n7755) );
  NAND2_X1 U9366 ( .A1(n9595), .A2(n9074), .ZN(n7754) );
  OAI211_X1 U9367 ( .C1(n9508), .C2(n9389), .A(n7755), .B(n7754), .ZN(n7756)
         );
  AOI21_X1 U9368 ( .B1(n9510), .B2(n9600), .A(n7756), .ZN(n7757) );
  OAI21_X1 U9369 ( .B1(n9512), .B2(n9377), .A(n7757), .ZN(P1_U3280) );
  INV_X1 U9370 ( .A(n7904), .ZN(n7769) );
  OAI222_X1 U9371 ( .A1(n7759), .A2(P1_U3084), .B1(n8245), .B2(n7769), .C1(
        n7758), .C2(n8242), .ZN(P1_U3327) );
  AOI22_X1 U9372 ( .A1(n8713), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7760), .B2(
        n9834), .ZN(n7761) );
  OAI21_X1 U9373 ( .B1(n7762), .B2(n8704), .A(n7761), .ZN(n7765) );
  NOR2_X1 U9374 ( .A1(n7763), .A2(n8713), .ZN(n7764) );
  AOI211_X1 U9375 ( .C1(n7766), .C2(n8716), .A(n7765), .B(n7764), .ZN(n7767)
         );
  OAI21_X1 U9376 ( .B1(n8718), .B2(n7768), .A(n7767), .ZN(P2_U3284) );
  OAI222_X1 U9377 ( .A1(P2_U3152), .A2(n7771), .B1(n8831), .B2(n7770), .C1(
        n8830), .C2(n7769), .ZN(P2_U3332) );
  NAND2_X1 U9378 ( .A1(n9306), .A2(n9078), .ZN(n7773) );
  NAND2_X1 U9379 ( .A1(n9304), .A2(n9073), .ZN(n7772) );
  NAND2_X1 U9380 ( .A1(n7773), .A2(n7772), .ZN(n9499) );
  NAND2_X1 U9381 ( .A1(n9633), .A2(n9499), .ZN(n7775) );
  OAI211_X1 U9382 ( .C1(n9648), .C2(n9592), .A(n7775), .B(n7774), .ZN(n7782)
         );
  XNOR2_X1 U9383 ( .A(n7778), .B(n7777), .ZN(n7779) );
  XNOR2_X1 U9384 ( .A(n7776), .B(n7779), .ZN(n7780) );
  NOR2_X1 U9385 ( .A1(n7780), .A2(n8972), .ZN(n7781) );
  AOI211_X1 U9386 ( .C1(n8970), .C2(n9596), .A(n7782), .B(n7781), .ZN(n7783)
         );
  INV_X1 U9387 ( .A(n7783), .ZN(P1_U3222) );
  INV_X1 U9388 ( .A(n7916), .ZN(n7788) );
  OAI222_X1 U9389 ( .A1(n8830), .A2(n7788), .B1(P2_U3152), .B2(n7955), .C1(
        n7784), .C2(n8831), .ZN(P2_U3331) );
  INV_X1 U9390 ( .A(n7925), .ZN(n8237) );
  NAND2_X1 U9391 ( .A1(n8828), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7785) );
  OAI211_X1 U9392 ( .C1(n8237), .C2(n8830), .A(n7786), .B(n7785), .ZN(P2_U3330) );
  OAI222_X1 U9393 ( .A1(P1_U3084), .A2(n7789), .B1(n8245), .B2(n7788), .C1(
        n7787), .C2(n8242), .ZN(P1_U3326) );
  XNOR2_X1 U9394 ( .A(n7859), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U9395 ( .A1(n8591), .A2(n7937), .ZN(n7795) );
  INV_X1 U9396 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U9397 ( .A1(n7882), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U9398 ( .A1(n7957), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7790) );
  OAI211_X1 U9399 ( .C1(n7934), .C2(n7792), .A(n7791), .B(n7790), .ZN(n7793)
         );
  INV_X1 U9400 ( .A(n7793), .ZN(n7794) );
  NAND2_X1 U9401 ( .A1(n7795), .A2(n7794), .ZN(n8439) );
  NAND2_X1 U9402 ( .A1(n7796), .A2(n7969), .ZN(n7798) );
  NAND2_X1 U9403 ( .A1(n7970), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U9404 ( .A1(n8797), .A2(n7800), .ZN(n8052) );
  INV_X1 U9405 ( .A(n8710), .ZN(n8665) );
  OR2_X1 U9406 ( .A1(n8792), .A2(n8665), .ZN(n8055) );
  NAND2_X1 U9407 ( .A1(n8792), .A2(n8665), .ZN(n8054) );
  NAND2_X1 U9408 ( .A1(n8055), .A2(n8054), .ZN(n8684) );
  NAND2_X1 U9409 ( .A1(n7801), .A2(n7969), .ZN(n7806) );
  OAI22_X1 U9410 ( .A1(n6907), .A2(n7803), .B1(n7832), .B2(n7802), .ZN(n7804)
         );
  INV_X1 U9411 ( .A(n7804), .ZN(n7805) );
  XNOR2_X1 U9412 ( .A(n8788), .B(n8693), .ZN(n8666) );
  NAND2_X1 U9413 ( .A1(n7808), .A2(n7969), .ZN(n7812) );
  OAI22_X1 U9414 ( .A1(n6907), .A2(n7809), .B1(n7832), .B2(n9800), .ZN(n7810)
         );
  INV_X1 U9415 ( .A(n7810), .ZN(n7811) );
  NAND2_X1 U9416 ( .A1(n7882), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U9417 ( .A1(n7957), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7818) );
  INV_X1 U9418 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U9419 ( .A1(n7814), .A2(n7813), .ZN(n7815) );
  AND2_X1 U9420 ( .A1(n7838), .A2(n7815), .ZN(n8655) );
  NAND2_X1 U9421 ( .A1(n7937), .A2(n8655), .ZN(n7817) );
  NAND2_X1 U9422 ( .A1(n7958), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7816) );
  NAND4_X1 U9423 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), .ZN(n8637)
         );
  INV_X1 U9424 ( .A(n8637), .ZN(n8663) );
  NAND2_X1 U9425 ( .A1(n8784), .A2(n8663), .ZN(n8064) );
  NAND2_X1 U9426 ( .A1(n8063), .A2(n8064), .ZN(n8644) );
  NAND2_X1 U9427 ( .A1(n7820), .A2(n7969), .ZN(n7824) );
  OAI22_X1 U9428 ( .A1(n6907), .A2(n7821), .B1(n7832), .B2(n8470), .ZN(n7822)
         );
  INV_X1 U9429 ( .A(n7822), .ZN(n7823) );
  XNOR2_X1 U9430 ( .A(n7838), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U9431 ( .A1(n8633), .A2(n7937), .ZN(n7828) );
  NAND2_X1 U9432 ( .A1(n7882), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U9433 ( .A1(n7958), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7826) );
  NAND2_X1 U9434 ( .A1(n7957), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7825) );
  NAND4_X1 U9435 ( .A1(n7828), .A2(n7827), .A3(n7826), .A4(n7825), .ZN(n8649)
         );
  NAND2_X1 U9436 ( .A1(n8777), .A2(n8649), .ZN(n7830) );
  INV_X1 U9437 ( .A(n8649), .ZN(n8378) );
  INV_X1 U9438 ( .A(n8777), .ZN(n8635) );
  AOI21_X1 U9439 ( .B1(n8630), .B2(n7830), .A(n7829), .ZN(n8618) );
  NAND2_X1 U9440 ( .A1(n7831), .A2(n7969), .ZN(n7836) );
  OAI22_X1 U9441 ( .A1(n6907), .A2(n7833), .B1(n7982), .B2(n7832), .ZN(n7834)
         );
  INV_X1 U9442 ( .A(n7834), .ZN(n7835) );
  INV_X1 U9443 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n7844) );
  INV_X1 U9444 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8414) );
  INV_X1 U9445 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7837) );
  OAI21_X1 U9446 ( .B1(n7838), .B2(n8414), .A(n7837), .ZN(n7839) );
  AND2_X1 U9447 ( .A1(n7839), .A2(n7850), .ZN(n8620) );
  NAND2_X1 U9448 ( .A1(n8620), .A2(n7937), .ZN(n7843) );
  NAND2_X1 U9449 ( .A1(n7957), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U9450 ( .A1(n7882), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7840) );
  AND2_X1 U9451 ( .A1(n7841), .A2(n7840), .ZN(n7842) );
  OAI211_X1 U9452 ( .C1(n7934), .C2(n7844), .A(n7843), .B(n7842), .ZN(n8638)
         );
  INV_X1 U9453 ( .A(n8638), .ZN(n8607) );
  NAND2_X1 U9454 ( .A1(n7847), .A2(n7969), .ZN(n7849) );
  NAND2_X1 U9455 ( .A1(n7970), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7848) );
  INV_X1 U9456 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n7854) );
  INV_X1 U9457 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U9458 ( .A1(n7850), .A2(n10095), .ZN(n7851) );
  NAND2_X1 U9459 ( .A1(n7859), .A2(n7851), .ZN(n8611) );
  OR2_X1 U9460 ( .A1(n8611), .A2(n4666), .ZN(n7853) );
  AOI22_X1 U9461 ( .A1(n7958), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n7882), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n7852) );
  OAI211_X1 U9462 ( .C1(n7875), .C2(n7854), .A(n7853), .B(n7852), .ZN(n8625)
         );
  INV_X1 U9463 ( .A(n8625), .ZN(n8349) );
  NAND2_X1 U9464 ( .A1(n8769), .A2(n8349), .ZN(n8081) );
  NAND2_X1 U9465 ( .A1(n8079), .A2(n8081), .ZN(n8603) );
  INV_X1 U9466 ( .A(n8762), .ZN(n8593) );
  INV_X1 U9467 ( .A(n8439), .ZN(n8608) );
  NAND2_X1 U9468 ( .A1(n7856), .A2(n7969), .ZN(n7858) );
  NAND2_X1 U9469 ( .A1(n7970), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7857) );
  INV_X1 U9470 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8346) );
  INV_X1 U9471 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8408) );
  OAI21_X1 U9472 ( .B1(n7859), .B2(n8346), .A(n8408), .ZN(n7860) );
  AND2_X1 U9473 ( .A1(n7860), .A2(n7870), .ZN(n8582) );
  NAND2_X1 U9474 ( .A1(n8582), .A2(n7937), .ZN(n7866) );
  INV_X1 U9475 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U9476 ( .A1(n7957), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U9477 ( .A1(n7882), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7861) );
  OAI211_X1 U9478 ( .C1(n7863), .C2(n7934), .A(n7862), .B(n7861), .ZN(n7864)
         );
  INV_X1 U9479 ( .A(n7864), .ZN(n7865) );
  NAND2_X1 U9480 ( .A1(n7866), .A2(n7865), .ZN(n8596) );
  NAND2_X1 U9481 ( .A1(n8759), .A2(n8347), .ZN(n8097) );
  NAND2_X1 U9482 ( .A1(n8085), .A2(n8097), .ZN(n8162) );
  INV_X1 U9483 ( .A(n8759), .ZN(n8585) );
  NAND2_X1 U9484 ( .A1(n7867), .A2(n7969), .ZN(n7869) );
  NAND2_X1 U9485 ( .A1(n7970), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7868) );
  INV_X1 U9486 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U9487 ( .A1(n7870), .A2(n8331), .ZN(n7871) );
  NAND2_X1 U9488 ( .A1(n7896), .A2(n7871), .ZN(n8568) );
  OR2_X1 U9489 ( .A1(n8568), .A2(n4666), .ZN(n7878) );
  INV_X1 U9490 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U9491 ( .A1(n7882), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7873) );
  NAND2_X1 U9492 ( .A1(n7958), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7872) );
  OAI211_X1 U9493 ( .C1(n7875), .C2(n7874), .A(n7873), .B(n7872), .ZN(n7876)
         );
  INV_X1 U9494 ( .A(n7876), .ZN(n7877) );
  NAND2_X1 U9495 ( .A1(n7878), .A2(n7877), .ZN(n8549) );
  INV_X1 U9496 ( .A(n8549), .ZN(n8392) );
  OR2_X1 U9497 ( .A1(n8752), .A2(n8392), .ZN(n8099) );
  NAND2_X1 U9498 ( .A1(n8752), .A2(n8392), .ZN(n8089) );
  NAND2_X1 U9499 ( .A1(n8099), .A2(n8089), .ZN(n8564) );
  INV_X1 U9500 ( .A(n8752), .ZN(n8571) );
  NAND2_X1 U9501 ( .A1(n7879), .A2(n7969), .ZN(n7881) );
  NAND2_X1 U9502 ( .A1(n7970), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7880) );
  XNOR2_X1 U9503 ( .A(n7896), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U9504 ( .A1(n8553), .A2(n7937), .ZN(n7888) );
  INV_X1 U9505 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U9506 ( .A1(n7957), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U9507 ( .A1(n7882), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7883) );
  OAI211_X1 U9508 ( .C1(n7885), .C2(n7934), .A(n7884), .B(n7883), .ZN(n7886)
         );
  INV_X1 U9509 ( .A(n7886), .ZN(n7887) );
  NAND2_X1 U9510 ( .A1(n8745), .A2(n8562), .ZN(n7889) );
  NAND2_X1 U9511 ( .A1(n7890), .A2(n7889), .ZN(n8540) );
  INV_X1 U9512 ( .A(n7890), .ZN(n7891) );
  NAND2_X1 U9513 ( .A1(n7892), .A2(n7969), .ZN(n7894) );
  NAND2_X1 U9514 ( .A1(n7970), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7893) );
  INV_X1 U9515 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8389) );
  INV_X1 U9516 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7895) );
  OAI21_X1 U9517 ( .B1(n7896), .B2(n8389), .A(n7895), .ZN(n7897) );
  NAND2_X1 U9518 ( .A1(n7897), .A2(n7907), .ZN(n8525) );
  OR2_X1 U9519 ( .A1(n8525), .A2(n4666), .ZN(n7903) );
  INV_X1 U9520 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U9521 ( .A1(n7957), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n7899) );
  NAND2_X1 U9522 ( .A1(n7882), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7898) );
  OAI211_X1 U9523 ( .C1(n7900), .C2(n7934), .A(n7899), .B(n7898), .ZN(n7901)
         );
  INV_X1 U9524 ( .A(n7901), .ZN(n7902) );
  NAND2_X1 U9525 ( .A1(n7903), .A2(n7902), .ZN(n8550) );
  INV_X1 U9526 ( .A(n8550), .ZN(n8390) );
  NAND2_X1 U9527 ( .A1(n8741), .A2(n8390), .ZN(n8094) );
  NAND2_X1 U9528 ( .A1(n7904), .A2(n7969), .ZN(n7906) );
  NAND2_X1 U9529 ( .A1(n7970), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7905) );
  NAND2_X1 U9530 ( .A1(n7907), .A2(n9968), .ZN(n7908) );
  NAND2_X1 U9531 ( .A1(n7929), .A2(n7908), .ZN(n8429) );
  INV_X1 U9532 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U9533 ( .A1(n7957), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7910) );
  NAND2_X1 U9534 ( .A1(n7958), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7909) );
  OAI211_X1 U9535 ( .C1(n7912), .C2(n7911), .A(n7910), .B(n7909), .ZN(n7913)
         );
  INV_X1 U9536 ( .A(n7913), .ZN(n7914) );
  NAND2_X1 U9537 ( .A1(n8737), .A2(n8109), .ZN(n7915) );
  INV_X1 U9538 ( .A(n8737), .ZN(n8517) );
  NAND2_X1 U9539 ( .A1(n7970), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7917) );
  XNOR2_X1 U9540 ( .A(n7929), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8497) );
  NAND2_X1 U9541 ( .A1(n8497), .A2(n7937), .ZN(n7924) );
  INV_X1 U9542 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U9543 ( .A1(n7882), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U9544 ( .A1(n7957), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7919) );
  OAI211_X1 U9545 ( .C1(n7921), .C2(n7934), .A(n7920), .B(n7919), .ZN(n7922)
         );
  INV_X1 U9546 ( .A(n7922), .ZN(n7923) );
  NAND2_X1 U9547 ( .A1(n7925), .A2(n7969), .ZN(n7927) );
  NAND2_X1 U9548 ( .A1(n7970), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7926) );
  INV_X1 U9549 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7928) );
  INV_X1 U9550 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8312) );
  OAI21_X1 U9551 ( .B1(n7929), .B2(n7928), .A(n8312), .ZN(n7930) );
  INV_X1 U9552 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U9553 ( .A1(n7957), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7933) );
  NAND2_X1 U9554 ( .A1(n7882), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n7932) );
  OAI211_X1 U9555 ( .C1(n7935), .C2(n7934), .A(n7933), .B(n7932), .ZN(n7936)
         );
  AOI21_X1 U9556 ( .B1(n8314), .B2(n7937), .A(n7936), .ZN(n8324) );
  NAND2_X1 U9557 ( .A1(n8724), .A2(n8324), .ZN(n8122) );
  INV_X1 U9558 ( .A(n8724), .ZN(n8223) );
  NAND2_X1 U9559 ( .A1(n8241), .A2(n7969), .ZN(n7939) );
  NAND2_X1 U9560 ( .A1(n7970), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U9561 ( .A1(n8719), .A2(n8313), .ZN(n8128) );
  NAND2_X1 U9562 ( .A1(n8127), .A2(n8128), .ZN(n8120) );
  XNOR2_X1 U9563 ( .A(n7940), .B(n8120), .ZN(n8722) );
  INV_X1 U9564 ( .A(n8784), .ZN(n8658) );
  OR2_X2 U9565 ( .A1(n8652), .A2(n8777), .ZN(n8631) );
  INV_X1 U9566 ( .A(n8769), .ZN(n8615) );
  NOR2_X2 U9567 ( .A1(n8581), .A2(n8752), .ZN(n8567) );
  INV_X1 U9568 ( .A(n8745), .ZN(n8544) );
  AND2_X2 U9569 ( .A1(n8567), .A2(n8544), .ZN(n8541) );
  AOI21_X1 U9570 ( .B1(n8719), .B2(n8219), .A(n8490), .ZN(n8720) );
  INV_X1 U9571 ( .A(n8719), .ZN(n7943) );
  AOI22_X1 U9572 ( .A1(n8713), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n7941), .B2(
        n9834), .ZN(n7942) );
  OAI21_X1 U9573 ( .B1(n7943), .B2(n8704), .A(n7942), .ZN(n7966) );
  INV_X1 U9574 ( .A(n8708), .ZN(n8698) );
  INV_X1 U9575 ( .A(n8706), .ZN(n7944) );
  NOR2_X1 U9576 ( .A1(n8698), .A2(n7944), .ZN(n7946) );
  INV_X1 U9577 ( .A(n8051), .ZN(n7945) );
  OR2_X1 U9578 ( .A1(n8788), .A2(n8059), .ZN(n7947) );
  INV_X1 U9579 ( .A(n8644), .ZN(n8647) );
  OR2_X1 U9580 ( .A1(n8777), .A2(n8378), .ZN(n8076) );
  NAND2_X1 U9581 ( .A1(n8777), .A2(n8378), .ZN(n8070) );
  OR2_X1 U9582 ( .A1(n8773), .A2(n8607), .ZN(n8078) );
  NAND2_X1 U9583 ( .A1(n8773), .A2(n8607), .ZN(n8602) );
  NAND2_X1 U9584 ( .A1(n8623), .A2(n8624), .ZN(n8622) );
  INV_X1 U9585 ( .A(n8602), .ZN(n8075) );
  NOR2_X1 U9586 ( .A1(n8603), .A2(n8075), .ZN(n7949) );
  NAND2_X1 U9587 ( .A1(n8622), .A2(n7949), .ZN(n7950) );
  OR2_X1 U9588 ( .A1(n8762), .A2(n8608), .ZN(n8084) );
  NAND2_X1 U9589 ( .A1(n8762), .A2(n8608), .ZN(n8080) );
  NAND2_X1 U9590 ( .A1(n8084), .A2(n8080), .ZN(n8594) );
  INV_X1 U9591 ( .A(n8162), .ZN(n8578) );
  INV_X1 U9592 ( .A(n8085), .ZN(n8558) );
  NOR2_X1 U9593 ( .A1(n8564), .A2(n8558), .ZN(n8091) );
  NAND2_X1 U9594 ( .A1(n8576), .A2(n8091), .ZN(n8560) );
  NAND2_X1 U9595 ( .A1(n8560), .A2(n8089), .ZN(n8546) );
  INV_X1 U9596 ( .A(n8546), .ZN(n7951) );
  INV_X1 U9597 ( .A(n8540), .ZN(n8545) );
  OR2_X1 U9598 ( .A1(n8745), .A2(n8358), .ZN(n8528) );
  INV_X1 U9599 ( .A(n8107), .ZN(n7952) );
  INV_X1 U9600 ( .A(n8438), .ZN(n8316) );
  NOR2_X1 U9601 ( .A1(n8730), .A2(n8316), .ZN(n8113) );
  INV_X1 U9602 ( .A(n8121), .ZN(n7953) );
  NAND2_X1 U9603 ( .A1(n7954), .A2(n7968), .ZN(n7964) );
  INV_X1 U9604 ( .A(n7955), .ZN(n8179) );
  NAND2_X1 U9605 ( .A1(n8179), .A2(P2_B_REG_SCAN_IN), .ZN(n7956) );
  AND2_X1 U9606 ( .A1(n9818), .A2(n7956), .ZN(n8486) );
  NAND2_X1 U9607 ( .A1(n7957), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U9608 ( .A1(n7882), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7960) );
  NAND2_X1 U9609 ( .A1(n7958), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7959) );
  NAND3_X1 U9610 ( .A1(n7961), .A2(n7960), .A3(n7959), .ZN(n8437) );
  AOI21_X2 U9611 ( .B1(n7964), .B2(n9816), .A(n7963), .ZN(n8721) );
  NOR2_X1 U9612 ( .A1(n8721), .A2(n8713), .ZN(n7965) );
  AOI211_X1 U9613 ( .C1(n8720), .C2(n8716), .A(n7966), .B(n7965), .ZN(n7967)
         );
  OAI21_X1 U9614 ( .B1(n8722), .B2(n8718), .A(n7967), .ZN(P2_U3267) );
  NAND2_X1 U9615 ( .A1(n8216), .A2(n7969), .ZN(n7972) );
  NAND2_X1 U9616 ( .A1(n7970), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U9617 ( .A1(n7978), .A2(n8173), .ZN(n7973) );
  OAI21_X1 U9618 ( .B1(n9584), .B2(n7973), .A(n8128), .ZN(n7975) );
  INV_X1 U9619 ( .A(n7973), .ZN(n7974) );
  INV_X1 U9620 ( .A(n8437), .ZN(n7979) );
  OAI22_X1 U9621 ( .A1(n9540), .A2(n7977), .B1(n6907), .B2(n6550), .ZN(n7980)
         );
  NOR2_X1 U9622 ( .A1(n7980), .A2(n7978), .ZN(n8136) );
  NOR2_X1 U9623 ( .A1(n8136), .A2(n8125), .ZN(n8168) );
  INV_X1 U9624 ( .A(n7980), .ZN(n9579) );
  NOR2_X1 U9625 ( .A1(n9579), .A2(n8487), .ZN(n8135) );
  INV_X1 U9626 ( .A(n8131), .ZN(n7984) );
  NOR2_X1 U9627 ( .A1(n8135), .A2(n7984), .ZN(n8169) );
  NAND2_X1 U9628 ( .A1(n8173), .A2(n7985), .ZN(n7986) );
  MUX2_X1 U9629 ( .A(n8168), .B(n8169), .S(n8137), .Z(n8134) );
  NAND2_X1 U9630 ( .A1(n7991), .A2(n7988), .ZN(n7990) );
  INV_X1 U9631 ( .A(n8008), .ZN(n7989) );
  MUX2_X1 U9632 ( .A(n7990), .B(n7989), .S(n8137), .Z(n7994) );
  OAI211_X1 U9633 ( .C1(n7994), .C2(n7992), .A(n8014), .B(n7991), .ZN(n7993)
         );
  NAND2_X1 U9634 ( .A1(n7993), .A2(n8137), .ZN(n8005) );
  INV_X1 U9635 ( .A(n7994), .ZN(n8011) );
  AND2_X1 U9636 ( .A1(n8142), .A2(n8173), .ZN(n7995) );
  OAI211_X1 U9637 ( .C1(n8145), .C2(n7995), .A(n8000), .B(n8143), .ZN(n7996)
         );
  NAND3_X1 U9638 ( .A1(n7996), .A2(n7999), .A3(n8137), .ZN(n7997) );
  NAND3_X1 U9639 ( .A1(n8011), .A2(n4741), .A3(n7997), .ZN(n8004) );
  NAND2_X1 U9640 ( .A1(n8143), .A2(n8142), .ZN(n7998) );
  NAND3_X1 U9641 ( .A1(n7999), .A2(n6236), .A3(n7998), .ZN(n8001) );
  INV_X1 U9642 ( .A(n8137), .ZN(n8126) );
  NAND3_X1 U9643 ( .A1(n8001), .A2(n8126), .A3(n8000), .ZN(n8002) );
  NAND2_X1 U9644 ( .A1(n8002), .A2(n8012), .ZN(n8003) );
  AOI21_X1 U9645 ( .B1(n8005), .B2(n8004), .A(n8003), .ZN(n8017) );
  INV_X1 U9646 ( .A(n8006), .ZN(n8010) );
  NAND2_X1 U9647 ( .A1(n8008), .A2(n8007), .ZN(n8009) );
  OAI21_X1 U9648 ( .B1(n8011), .B2(n8010), .A(n8009), .ZN(n8013) );
  AOI21_X1 U9649 ( .B1(n8013), .B2(n8012), .A(n8137), .ZN(n8016) );
  NOR2_X1 U9650 ( .A1(n8014), .A2(n8137), .ZN(n8015) );
  MUX2_X1 U9651 ( .A(n8019), .B(n8018), .S(n8137), .Z(n8020) );
  MUX2_X1 U9652 ( .A(n8022), .B(n8021), .S(n8137), .Z(n8024) );
  NAND3_X1 U9653 ( .A1(n8030), .A2(n8032), .A3(n8027), .ZN(n8026) );
  NAND3_X1 U9654 ( .A1(n8026), .A2(n8025), .A3(n8031), .ZN(n8037) );
  INV_X1 U9655 ( .A(n8027), .ZN(n8028) );
  INV_X1 U9656 ( .A(n8031), .ZN(n8034) );
  OAI211_X1 U9657 ( .C1(n8035), .C2(n8034), .A(n8033), .B(n8032), .ZN(n8036)
         );
  MUX2_X1 U9658 ( .A(n8037), .B(n8036), .S(n8137), .Z(n8039) );
  NAND2_X1 U9659 ( .A1(n8039), .A2(n4590), .ZN(n8038) );
  INV_X1 U9660 ( .A(n8039), .ZN(n8047) );
  NAND2_X1 U9661 ( .A1(n8040), .A2(n8126), .ZN(n8044) );
  NAND2_X1 U9662 ( .A1(n8042), .A2(n8041), .ZN(n8043) );
  MUX2_X1 U9663 ( .A(n8044), .B(n8043), .S(n8441), .Z(n8046) );
  MUX2_X1 U9664 ( .A(n8048), .B(n8706), .S(n8137), .Z(n8049) );
  MUX2_X1 U9665 ( .A(n8052), .B(n8051), .S(n8137), .Z(n8053) );
  MUX2_X1 U9666 ( .A(n8055), .B(n8054), .S(n8137), .Z(n8056) );
  NAND2_X1 U9667 ( .A1(n8057), .A2(n8056), .ZN(n8058) );
  NAND2_X1 U9668 ( .A1(n8693), .A2(n8126), .ZN(n8061) );
  NAND2_X1 U9669 ( .A1(n8059), .A2(n8137), .ZN(n8060) );
  MUX2_X1 U9670 ( .A(n8061), .B(n8060), .S(n8788), .Z(n8062) );
  INV_X1 U9671 ( .A(n8063), .ZN(n8066) );
  NAND2_X1 U9672 ( .A1(n8070), .A2(n8064), .ZN(n8065) );
  MUX2_X1 U9673 ( .A(n8066), .B(n8065), .S(n8126), .Z(n8068) );
  INV_X1 U9674 ( .A(n8076), .ZN(n8067) );
  NOR2_X1 U9675 ( .A1(n8068), .A2(n8067), .ZN(n8069) );
  NAND2_X1 U9676 ( .A1(n8071), .A2(n8078), .ZN(n8072) );
  NAND3_X1 U9677 ( .A1(n8072), .A2(n8081), .A3(n8602), .ZN(n8073) );
  NAND3_X1 U9678 ( .A1(n8073), .A2(n8079), .A3(n8084), .ZN(n8074) );
  NAND3_X1 U9679 ( .A1(n8074), .A2(n8097), .A3(n8080), .ZN(n8088) );
  AOI21_X1 U9680 ( .B1(n8077), .B2(n8076), .A(n8075), .ZN(n8083) );
  NAND2_X1 U9681 ( .A1(n8079), .A2(n8078), .ZN(n8082) );
  OAI211_X1 U9682 ( .C1(n8083), .C2(n8082), .A(n8081), .B(n8080), .ZN(n8086)
         );
  NAND3_X1 U9683 ( .A1(n8086), .A2(n8085), .A3(n8084), .ZN(n8087) );
  INV_X1 U9684 ( .A(n8089), .ZN(n8090) );
  AOI21_X1 U9685 ( .B1(n8098), .B2(n8091), .A(n8090), .ZN(n8095) );
  NAND2_X1 U9686 ( .A1(n8745), .A2(n8358), .ZN(n8092) );
  MUX2_X1 U9687 ( .A(n8092), .B(n8528), .S(n8137), .Z(n8093) );
  NAND2_X1 U9688 ( .A1(n8530), .A2(n8093), .ZN(n8101) );
  INV_X1 U9689 ( .A(n8509), .ZN(n8507) );
  OAI211_X1 U9690 ( .C1(n8095), .C2(n8101), .A(n8507), .B(n8094), .ZN(n8096)
         );
  NAND2_X1 U9691 ( .A1(n8096), .A2(n8137), .ZN(n8106) );
  INV_X1 U9692 ( .A(n8564), .ZN(n8164) );
  NAND3_X1 U9693 ( .A1(n8098), .A2(n8164), .A3(n8097), .ZN(n8100) );
  AOI21_X1 U9694 ( .B1(n8100), .B2(n8099), .A(n8137), .ZN(n8103) );
  INV_X1 U9695 ( .A(n8101), .ZN(n8102) );
  OAI21_X1 U9696 ( .B1(n8103), .B2(n8545), .A(n8102), .ZN(n8105) );
  INV_X1 U9697 ( .A(n8108), .ZN(n8104) );
  AOI21_X1 U9698 ( .B1(n8106), .B2(n8105), .A(n8104), .ZN(n8112) );
  AOI21_X1 U9699 ( .B1(n8108), .B2(n8107), .A(n8137), .ZN(n8111) );
  NAND3_X1 U9700 ( .A1(n8737), .A2(n8109), .A3(n8126), .ZN(n8110) );
  OAI211_X1 U9701 ( .C1(n8112), .C2(n8111), .A(n8501), .B(n8110), .ZN(n8119)
         );
  INV_X1 U9702 ( .A(n8113), .ZN(n8114) );
  AND2_X1 U9703 ( .A1(n8114), .A2(n8121), .ZN(n8117) );
  AND2_X1 U9704 ( .A1(n8730), .A2(n8316), .ZN(n8115) );
  NOR2_X1 U9705 ( .A1(n8225), .A2(n8115), .ZN(n8116) );
  MUX2_X1 U9706 ( .A(n8117), .B(n8116), .S(n8137), .Z(n8118) );
  NAND2_X1 U9707 ( .A1(n8119), .A2(n8118), .ZN(n8124) );
  MUX2_X1 U9708 ( .A(n8122), .B(n8121), .S(n8137), .Z(n8123) );
  NAND3_X1 U9709 ( .A1(n8124), .A2(n4649), .A3(n8123), .ZN(n8132) );
  INV_X1 U9710 ( .A(n8125), .ZN(n8130) );
  MUX2_X1 U9711 ( .A(n8128), .B(n8127), .S(n8126), .Z(n8129) );
  NAND4_X1 U9712 ( .A1(n8132), .A2(n8131), .A3(n8130), .A4(n8129), .ZN(n8133)
         );
  NAND2_X1 U9713 ( .A1(n8134), .A2(n8133), .ZN(n8141) );
  INV_X1 U9714 ( .A(n8135), .ZN(n8139) );
  INV_X1 U9715 ( .A(n8136), .ZN(n8138) );
  MUX2_X1 U9716 ( .A(n8139), .B(n8138), .S(n8137), .Z(n8140) );
  INV_X1 U9717 ( .A(n8501), .ZN(n8166) );
  NAND4_X1 U9718 ( .A1(n8144), .A2(n8172), .A3(n8143), .A4(n8142), .ZN(n8147)
         );
  OR4_X1 U9719 ( .A1(n8147), .A2(n8146), .A3(n9813), .A4(n8145), .ZN(n8151) );
  NOR4_X1 U9720 ( .A1(n8151), .A2(n8150), .A3(n8149), .A4(n8148), .ZN(n8155)
         );
  NAND4_X1 U9721 ( .A1(n8155), .A2(n8154), .A3(n8153), .A4(n8152), .ZN(n8158)
         );
  OR4_X1 U9722 ( .A1(n7669), .A2(n8158), .A3(n8157), .A4(n8156), .ZN(n8159) );
  NOR4_X1 U9723 ( .A1(n8644), .A2(n8684), .A3(n8698), .A4(n8159), .ZN(n8160)
         );
  NAND4_X1 U9724 ( .A1(n8624), .A2(n4338), .A3(n8160), .A4(n8666), .ZN(n8161)
         );
  NOR4_X1 U9725 ( .A1(n8162), .A2(n8603), .A3(n8594), .A4(n8161), .ZN(n8163)
         );
  NAND4_X1 U9726 ( .A1(n8530), .A2(n8164), .A3(n8163), .A4(n8540), .ZN(n8165)
         );
  NOR4_X1 U9727 ( .A1(n8225), .A2(n8166), .A3(n8509), .A4(n8165), .ZN(n8167)
         );
  NAND4_X1 U9728 ( .A1(n8169), .A2(n8168), .A3(n4649), .A4(n8167), .ZN(n8170)
         );
  XNOR2_X1 U9729 ( .A(n8170), .B(n7982), .ZN(n8174) );
  OAI22_X1 U9730 ( .A1(n8174), .A2(n8173), .B1(n8172), .B2(n8171), .ZN(n8175)
         );
  NAND4_X1 U9731 ( .A1(n8180), .A2(n8179), .A3(n8178), .A4(n9821), .ZN(n8181)
         );
  OAI211_X1 U9732 ( .C1(n6234), .C2(n8183), .A(n8181), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8182) );
  NOR2_X1 U9733 ( .A1(n9327), .A2(n8184), .ZN(n8185) );
  NOR2_X1 U9734 ( .A1(n5772), .A2(n9605), .ZN(n9069) );
  AOI211_X1 U9735 ( .C1(n8186), .C2(n9595), .A(n8185), .B(n9069), .ZN(n8187)
         );
  OAI21_X1 U9736 ( .B1(n8188), .B2(n9389), .A(n8187), .ZN(P1_U3261) );
  OAI222_X1 U9737 ( .A1(n8831), .A2(n8191), .B1(n8830), .B2(n8190), .C1(n8189), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U9738 ( .A1(n9420), .A2(n8192), .ZN(n8194) );
  NAND2_X1 U9739 ( .A1(n9108), .A2(n8199), .ZN(n8193) );
  NAND2_X1 U9740 ( .A1(n8194), .A2(n8193), .ZN(n8196) );
  XNOR2_X1 U9741 ( .A(n8196), .B(n8195), .ZN(n8201) );
  NOR2_X1 U9742 ( .A1(n9176), .A2(n8197), .ZN(n8198) );
  AOI21_X1 U9743 ( .B1(n9420), .B2(n8199), .A(n8198), .ZN(n8200) );
  XNOR2_X1 U9744 ( .A(n8201), .B(n8200), .ZN(n8202) );
  INV_X1 U9745 ( .A(n8202), .ZN(n8208) );
  NAND3_X1 U9746 ( .A1(n8209), .A2(n9643), .A3(n8208), .ZN(n8214) );
  NAND3_X1 U9747 ( .A1(n8215), .A2(n9643), .A3(n8202), .ZN(n8213) );
  OR2_X1 U9748 ( .A1(n8951), .A2(n9552), .ZN(n8204) );
  NAND2_X1 U9749 ( .A1(n8974), .A2(n9306), .ZN(n8203) );
  NAND2_X1 U9750 ( .A1(n8204), .A2(n8203), .ZN(n9161) );
  INV_X1 U9751 ( .A(n9161), .ZN(n8207) );
  INV_X1 U9752 ( .A(n8205), .ZN(n9155) );
  AOI22_X1 U9753 ( .A1(n9155), .A2(n8930), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8206) );
  OAI21_X1 U9754 ( .B1(n8207), .B2(n8884), .A(n8206), .ZN(n8211) );
  NOR3_X1 U9755 ( .A1(n8209), .A2(n8208), .A3(n8972), .ZN(n8210) );
  AOI211_X1 U9756 ( .C1(n8970), .C2(n9420), .A(n8211), .B(n8210), .ZN(n8212)
         );
  OAI211_X1 U9757 ( .C1(n8215), .C2(n8214), .A(n8213), .B(n8212), .ZN(P1_U3218) );
  INV_X1 U9758 ( .A(n8216), .ZN(n8240) );
  OAI222_X1 U9759 ( .A1(n8242), .A2(n8217), .B1(n9539), .B2(n8240), .C1(
        P1_U3084), .C2(n5076), .ZN(P1_U3323) );
  XNOR2_X1 U9760 ( .A(n8218), .B(n4472), .ZN(n8723) );
  INV_X1 U9761 ( .A(n8219), .ZN(n8220) );
  AOI21_X1 U9762 ( .B1(n8724), .B2(n8221), .A(n8220), .ZN(n8725) );
  AOI22_X1 U9763 ( .A1(n8713), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8314), .B2(
        n9834), .ZN(n8222) );
  OAI21_X1 U9764 ( .B1(n8223), .B2(n8704), .A(n8222), .ZN(n8228) );
  AOI211_X1 U9765 ( .C1(n8226), .C2(n8225), .A(n8605), .B(n8224), .ZN(n8227)
         );
  INV_X1 U9766 ( .A(n8229), .ZN(n8230) );
  AOI22_X1 U9767 ( .A1(n9600), .A2(n8230), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9377), .ZN(n8235) );
  INV_X1 U9768 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9649) );
  OAI22_X1 U9769 ( .A1(n8231), .A2(n9061), .B1(n9559), .B2(n9649), .ZN(n8232)
         );
  OAI21_X1 U9770 ( .B1(n8233), .B2(n8232), .A(n9327), .ZN(n8234) );
  OAI211_X1 U9771 ( .C1(n8236), .C2(n9401), .A(n8235), .B(n8234), .ZN(P1_U3290) );
  OAI222_X1 U9772 ( .A1(n8242), .A2(n8238), .B1(P1_U3084), .B2(n5754), .C1(
        n8237), .C2(n8245), .ZN(P1_U3325) );
  OAI222_X1 U9773 ( .A1(n8831), .A2(n10137), .B1(n8830), .B2(n8240), .C1(n8239), .C2(P2_U3152), .ZN(P2_U3328) );
  INV_X1 U9774 ( .A(n8241), .ZN(n8834) );
  XNOR2_X1 U9775 ( .A(n8788), .B(n8300), .ZN(n8250) );
  NAND2_X1 U9776 ( .A1(n8693), .A2(n8301), .ZN(n8251) );
  NAND2_X1 U9777 ( .A1(n8250), .A2(n8251), .ZN(n8257) );
  INV_X1 U9778 ( .A(n8250), .ZN(n8253) );
  INV_X1 U9779 ( .A(n8251), .ZN(n8252) );
  NAND2_X1 U9780 ( .A1(n8253), .A2(n8252), .ZN(n8254) );
  NAND2_X1 U9781 ( .A1(n8257), .A2(n8254), .ZN(n8368) );
  INV_X1 U9782 ( .A(n8368), .ZN(n8255) );
  XNOR2_X1 U9783 ( .A(n8784), .B(n8300), .ZN(n8259) );
  NAND2_X1 U9784 ( .A1(n8637), .A2(n8301), .ZN(n8258) );
  XNOR2_X1 U9785 ( .A(n8259), .B(n8258), .ZN(n8374) );
  XNOR2_X1 U9786 ( .A(n8777), .B(n4322), .ZN(n8263) );
  NAND2_X1 U9787 ( .A1(n8649), .A2(n8301), .ZN(n8261) );
  XNOR2_X1 U9788 ( .A(n8263), .B(n8261), .ZN(n8412) );
  INV_X1 U9789 ( .A(n8261), .ZN(n8262) );
  INV_X1 U9790 ( .A(n8339), .ZN(n8270) );
  XNOR2_X1 U9791 ( .A(n8773), .B(n8300), .ZN(n8264) );
  NAND2_X1 U9792 ( .A1(n8638), .A2(n8301), .ZN(n8265) );
  NAND2_X1 U9793 ( .A1(n8264), .A2(n8265), .ZN(n8271) );
  INV_X1 U9794 ( .A(n8264), .ZN(n8267) );
  INV_X1 U9795 ( .A(n8265), .ZN(n8266) );
  NAND2_X1 U9796 ( .A1(n8267), .A2(n8266), .ZN(n8268) );
  NAND2_X1 U9797 ( .A1(n8271), .A2(n8268), .ZN(n8338) );
  XNOR2_X1 U9798 ( .A(n8769), .B(n8300), .ZN(n8273) );
  NAND2_X1 U9799 ( .A1(n8625), .A2(n8301), .ZN(n8272) );
  XNOR2_X1 U9800 ( .A(n8273), .B(n8272), .ZN(n8397) );
  XNOR2_X1 U9801 ( .A(n8762), .B(n4322), .ZN(n8277) );
  NAND2_X1 U9802 ( .A1(n8439), .A2(n8301), .ZN(n8275) );
  XNOR2_X1 U9803 ( .A(n8277), .B(n8275), .ZN(n8344) );
  INV_X1 U9804 ( .A(n8275), .ZN(n8276) );
  XNOR2_X1 U9805 ( .A(n8759), .B(n8300), .ZN(n8279) );
  XNOR2_X1 U9806 ( .A(n8278), .B(n8279), .ZN(n8405) );
  NAND2_X1 U9807 ( .A1(n8596), .A2(n8301), .ZN(n8404) );
  NAND2_X1 U9808 ( .A1(n8405), .A2(n8404), .ZN(n8403) );
  INV_X1 U9809 ( .A(n8279), .ZN(n8280) );
  INV_X1 U9810 ( .A(n8330), .ZN(n8286) );
  INV_X1 U9811 ( .A(n8386), .ZN(n8283) );
  NAND2_X1 U9812 ( .A1(n8549), .A2(n8301), .ZN(n8384) );
  INV_X1 U9813 ( .A(n8384), .ZN(n8282) );
  OAI21_X1 U9814 ( .B1(n8283), .B2(n8562), .A(n8282), .ZN(n8284) );
  INV_X1 U9815 ( .A(n8284), .ZN(n8285) );
  AND2_X1 U9816 ( .A1(n8562), .A2(n8301), .ZN(n8385) );
  INV_X1 U9817 ( .A(n8385), .ZN(n8288) );
  NAND2_X1 U9818 ( .A1(n8386), .A2(n8288), .ZN(n8290) );
  XNOR2_X1 U9819 ( .A(n8741), .B(n4322), .ZN(n8293) );
  INV_X1 U9820 ( .A(n8293), .ZN(n8355) );
  NAND2_X1 U9821 ( .A1(n8294), .A2(n8293), .ZN(n8295) );
  NAND2_X1 U9822 ( .A1(n8550), .A2(n8301), .ZN(n8354) );
  XNOR2_X1 U9823 ( .A(n8737), .B(n8300), .ZN(n8297) );
  NAND2_X1 U9824 ( .A1(n8502), .A2(n8301), .ZN(n8296) );
  NOR2_X1 U9825 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  AOI21_X1 U9826 ( .B1(n8297), .B2(n8296), .A(n8298), .ZN(n8427) );
  NAND2_X1 U9827 ( .A1(n8428), .A2(n8427), .ZN(n8426) );
  INV_X1 U9828 ( .A(n8298), .ZN(n8299) );
  NAND2_X1 U9829 ( .A1(n8426), .A2(n8299), .ZN(n8323) );
  XNOR2_X1 U9830 ( .A(n8730), .B(n8300), .ZN(n8303) );
  NAND2_X1 U9831 ( .A1(n8438), .A2(n8301), .ZN(n8302) );
  NOR2_X1 U9832 ( .A1(n8303), .A2(n8302), .ZN(n8304) );
  AOI21_X1 U9833 ( .B1(n8303), .B2(n8302), .A(n8304), .ZN(n8322) );
  NAND2_X1 U9834 ( .A1(n8323), .A2(n8322), .ZN(n8321) );
  INV_X1 U9835 ( .A(n8304), .ZN(n8305) );
  NAND2_X1 U9836 ( .A1(n8321), .A2(n8305), .ZN(n8311) );
  NOR2_X1 U9837 ( .A1(n8324), .A2(n8306), .ZN(n8307) );
  XOR2_X1 U9838 ( .A(n4322), .B(n8307), .Z(n8309) );
  XNOR2_X1 U9839 ( .A(n8724), .B(n8309), .ZN(n8310) );
  XNOR2_X1 U9840 ( .A(n8311), .B(n8310), .ZN(n8320) );
  OAI22_X1 U9841 ( .A1(n8415), .A2(n8313), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8312), .ZN(n8318) );
  INV_X1 U9842 ( .A(n8314), .ZN(n8315) );
  OAI22_X1 U9843 ( .A1(n8418), .A2(n8316), .B1(n8416), .B2(n8315), .ZN(n8317)
         );
  AOI211_X1 U9844 ( .C1(n8724), .C2(n8421), .A(n8318), .B(n8317), .ZN(n8319)
         );
  OAI21_X1 U9845 ( .B1(n8320), .B2(n8423), .A(n8319), .ZN(P2_U3222) );
  OAI211_X1 U9846 ( .C1(n8323), .C2(n8322), .A(n8321), .B(n8425), .ZN(n8329)
         );
  AOI22_X1 U9847 ( .A1(n4484), .A2(n8325), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8328) );
  AOI22_X1 U9848 ( .A1(n8376), .A2(n8502), .B1(n8497), .B2(n8433), .ZN(n8327)
         );
  NAND2_X1 U9849 ( .A1(n8730), .A2(n8421), .ZN(n8326) );
  NAND4_X1 U9850 ( .A1(n8329), .A2(n8328), .A3(n8327), .A4(n8326), .ZN(
        P2_U3216) );
  XNOR2_X1 U9851 ( .A(n8330), .B(n8384), .ZN(n8335) );
  OAI22_X1 U9852 ( .A1(n8415), .A2(n8358), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8331), .ZN(n8333) );
  OAI22_X1 U9853 ( .A1(n8418), .A2(n8347), .B1(n8416), .B2(n8568), .ZN(n8332)
         );
  AOI211_X1 U9854 ( .C1(n8752), .C2(n8421), .A(n8333), .B(n8332), .ZN(n8334)
         );
  OAI21_X1 U9855 ( .B1(n8335), .B2(n8423), .A(n8334), .ZN(P2_U3218) );
  INV_X1 U9856 ( .A(n8336), .ZN(n8337) );
  AOI21_X1 U9857 ( .B1(n8339), .B2(n8338), .A(n8337), .ZN(n8343) );
  AOI22_X1 U9858 ( .A1(n8376), .A2(n8649), .B1(n8620), .B2(n8433), .ZN(n8340)
         );
  NAND2_X1 U9859 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8481) );
  OAI211_X1 U9860 ( .C1(n8349), .C2(n8415), .A(n8340), .B(n8481), .ZN(n8341)
         );
  AOI21_X1 U9861 ( .B1(n8773), .B2(n8421), .A(n8341), .ZN(n8342) );
  OAI21_X1 U9862 ( .B1(n8343), .B2(n8423), .A(n8342), .ZN(P2_U3221) );
  XNOR2_X1 U9863 ( .A(n8345), .B(n8344), .ZN(n8353) );
  OAI22_X1 U9864 ( .A1(n8415), .A2(n8347), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8346), .ZN(n8351) );
  INV_X1 U9865 ( .A(n8591), .ZN(n8348) );
  OAI22_X1 U9866 ( .A1(n8418), .A2(n8349), .B1(n8348), .B2(n8416), .ZN(n8350)
         );
  AOI211_X1 U9867 ( .C1(n8762), .C2(n8421), .A(n8351), .B(n8350), .ZN(n8352)
         );
  OAI21_X1 U9868 ( .B1(n8353), .B2(n8423), .A(n8352), .ZN(P2_U3225) );
  XNOR2_X1 U9869 ( .A(n8355), .B(n8354), .ZN(n8356) );
  XNOR2_X1 U9870 ( .A(n8357), .B(n8356), .ZN(n8364) );
  NAND2_X1 U9871 ( .A1(n8502), .A2(n9818), .ZN(n8360) );
  OR2_X1 U9872 ( .A1(n8358), .A2(n8664), .ZN(n8359) );
  NAND2_X1 U9873 ( .A1(n8360), .A2(n8359), .ZN(n8533) );
  AOI22_X1 U9874 ( .A1(n8533), .A2(n8407), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8361) );
  OAI21_X1 U9875 ( .B1(n8525), .B2(n8416), .A(n8361), .ZN(n8362) );
  AOI21_X1 U9876 ( .B1(n8741), .B2(n8421), .A(n8362), .ZN(n8363) );
  OAI21_X1 U9877 ( .B1(n8364), .B2(n8423), .A(n8363), .ZN(P2_U3227) );
  INV_X1 U9878 ( .A(n4405), .ZN(n8367) );
  AOI21_X1 U9879 ( .B1(n8368), .B2(n8365), .A(n8367), .ZN(n8373) );
  AOI22_X1 U9880 ( .A1(n8376), .A2(n8710), .B1(n8675), .B2(n8433), .ZN(n8370)
         );
  OAI211_X1 U9881 ( .C1(n8663), .C2(n8415), .A(n8370), .B(n8369), .ZN(n8371)
         );
  AOI21_X1 U9882 ( .B1(n8788), .B2(n8421), .A(n8371), .ZN(n8372) );
  OAI21_X1 U9883 ( .B1(n8373), .B2(n8423), .A(n8372), .ZN(P2_U3228) );
  XNOR2_X1 U9884 ( .A(n8375), .B(n8374), .ZN(n8381) );
  AOI22_X1 U9885 ( .A1(n8376), .A2(n8693), .B1(n8655), .B2(n8433), .ZN(n8377)
         );
  NAND2_X1 U9886 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9793) );
  OAI211_X1 U9887 ( .C1(n8378), .C2(n8415), .A(n8377), .B(n9793), .ZN(n8379)
         );
  AOI21_X1 U9888 ( .B1(n8784), .B2(n8421), .A(n8379), .ZN(n8380) );
  OAI21_X1 U9889 ( .B1(n8381), .B2(n8423), .A(n8380), .ZN(P2_U3230) );
  INV_X1 U9890 ( .A(n8382), .ZN(n8383) );
  OAI21_X1 U9891 ( .B1(n8330), .B2(n8384), .A(n8383), .ZN(n8388) );
  XNOR2_X1 U9892 ( .A(n8386), .B(n8385), .ZN(n8387) );
  XNOR2_X1 U9893 ( .A(n8388), .B(n8387), .ZN(n8396) );
  OAI22_X1 U9894 ( .A1(n8415), .A2(n8390), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8389), .ZN(n8394) );
  INV_X1 U9895 ( .A(n8553), .ZN(n8391) );
  OAI22_X1 U9896 ( .A1(n8418), .A2(n8392), .B1(n8391), .B2(n8416), .ZN(n8393)
         );
  AOI211_X1 U9897 ( .C1(n8745), .C2(n8421), .A(n8394), .B(n8393), .ZN(n8395)
         );
  OAI21_X1 U9898 ( .B1(n8396), .B2(n8423), .A(n8395), .ZN(P2_U3231) );
  XNOR2_X1 U9899 ( .A(n8398), .B(n8397), .ZN(n8402) );
  OAI22_X1 U9900 ( .A1(n8415), .A2(n8608), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10095), .ZN(n8400) );
  OAI22_X1 U9901 ( .A1(n8418), .A2(n8607), .B1(n8611), .B2(n8416), .ZN(n8399)
         );
  AOI211_X1 U9902 ( .C1(n8769), .C2(n8421), .A(n8400), .B(n8399), .ZN(n8401)
         );
  OAI21_X1 U9903 ( .B1(n8402), .B2(n8423), .A(n8401), .ZN(P2_U3235) );
  OAI21_X1 U9904 ( .B1(n8405), .B2(n8404), .A(n8403), .ZN(n8406) );
  NAND2_X1 U9905 ( .A1(n8406), .A2(n8425), .ZN(n8411) );
  INV_X1 U9906 ( .A(n8407), .ZN(n8431) );
  AOI22_X1 U9907 ( .A1(n8549), .A2(n9818), .B1(n9821), .B2(n8439), .ZN(n8579)
         );
  OAI22_X1 U9908 ( .A1(n8431), .A2(n8579), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8408), .ZN(n8409) );
  AOI21_X1 U9909 ( .B1(n8582), .B2(n8433), .A(n8409), .ZN(n8410) );
  OAI211_X1 U9910 ( .C1(n8585), .C2(n8436), .A(n8411), .B(n8410), .ZN(P2_U3237) );
  XNOR2_X1 U9911 ( .A(n8413), .B(n8412), .ZN(n8424) );
  OAI22_X1 U9912 ( .A1(n8415), .A2(n8607), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8414), .ZN(n8420) );
  INV_X1 U9913 ( .A(n8633), .ZN(n8417) );
  OAI22_X1 U9914 ( .A1(n8418), .A2(n8663), .B1(n8417), .B2(n8416), .ZN(n8419)
         );
  AOI211_X1 U9915 ( .C1(n8777), .C2(n8421), .A(n8420), .B(n8419), .ZN(n8422)
         );
  OAI21_X1 U9916 ( .B1(n8424), .B2(n8423), .A(n8422), .ZN(P2_U3240) );
  OAI211_X1 U9917 ( .C1(n8428), .C2(n8427), .A(n8426), .B(n8425), .ZN(n8435)
         );
  INV_X1 U9918 ( .A(n8429), .ZN(n8514) );
  AND2_X1 U9919 ( .A1(n8550), .A2(n9821), .ZN(n8430) );
  AOI21_X1 U9920 ( .B1(n8438), .B2(n9818), .A(n8430), .ZN(n8511) );
  OAI22_X1 U9921 ( .A1(n8511), .A2(n8431), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9968), .ZN(n8432) );
  AOI21_X1 U9922 ( .B1(n8514), .B2(n8433), .A(n8432), .ZN(n8434) );
  OAI211_X1 U9923 ( .C1(n8517), .C2(n8436), .A(n8435), .B(n8434), .ZN(P2_U3242) );
  MUX2_X1 U9924 ( .A(n8437), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8448), .Z(
        P2_U3582) );
  MUX2_X1 U9925 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n4484), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9926 ( .A(n8438), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8448), .Z(
        P2_U3579) );
  MUX2_X1 U9927 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8502), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9928 ( .A(n8550), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8448), .Z(
        P2_U3577) );
  MUX2_X1 U9929 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8562), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9930 ( .A(n8549), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8448), .Z(
        P2_U3575) );
  MUX2_X1 U9931 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8596), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9932 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8439), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9933 ( .A(n8625), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8448), .Z(
        P2_U3572) );
  MUX2_X1 U9934 ( .A(n8638), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8448), .Z(
        P2_U3571) );
  MUX2_X1 U9935 ( .A(n8649), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8448), .Z(
        P2_U3570) );
  MUX2_X1 U9936 ( .A(n8637), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8448), .Z(
        P2_U3569) );
  MUX2_X1 U9937 ( .A(n8693), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8448), .Z(
        P2_U3568) );
  MUX2_X1 U9938 ( .A(n8710), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8448), .Z(
        P2_U3567) );
  MUX2_X1 U9939 ( .A(n8692), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8448), .Z(
        P2_U3566) );
  MUX2_X1 U9940 ( .A(n8711), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8448), .Z(
        P2_U3565) );
  MUX2_X1 U9941 ( .A(n8440), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8448), .Z(
        P2_U3564) );
  MUX2_X1 U9942 ( .A(n8441), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8448), .Z(
        P2_U3563) );
  MUX2_X1 U9943 ( .A(n8442), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8448), .Z(
        P2_U3562) );
  MUX2_X1 U9944 ( .A(n8443), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8448), .Z(
        P2_U3561) );
  MUX2_X1 U9945 ( .A(n8444), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8448), .Z(
        P2_U3560) );
  MUX2_X1 U9946 ( .A(n8445), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8448), .Z(
        P2_U3559) );
  MUX2_X1 U9947 ( .A(n8446), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8448), .Z(
        P2_U3558) );
  MUX2_X1 U9948 ( .A(n8447), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8448), .Z(
        P2_U3557) );
  MUX2_X1 U9949 ( .A(n9819), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8448), .Z(
        P2_U3556) );
  MUX2_X1 U9950 ( .A(n6771), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8448), .Z(
        P2_U3555) );
  MUX2_X1 U9951 ( .A(n9820), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8448), .Z(
        P2_U3554) );
  MUX2_X1 U9952 ( .A(n6206), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8448), .Z(
        P2_U3553) );
  OAI211_X1 U9953 ( .C1(n8451), .C2(n8450), .A(n9797), .B(n8449), .ZN(n8462)
         );
  INV_X1 U9954 ( .A(n8452), .ZN(n8453) );
  AOI21_X1 U9955 ( .B1(n9795), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8453), .ZN(
        n8461) );
  INV_X1 U9956 ( .A(n8454), .ZN(n8455) );
  NAND2_X1 U9957 ( .A1(n9802), .A2(n8455), .ZN(n8460) );
  OAI211_X1 U9958 ( .C1(n8458), .C2(n8457), .A(n9804), .B(n8456), .ZN(n8459)
         );
  NAND4_X1 U9959 ( .A1(n8462), .A2(n8461), .A3(n8460), .A4(n8459), .ZN(
        P2_U3254) );
  NOR2_X1 U9960 ( .A1(n8464), .A2(n8463), .ZN(n8465) );
  NOR2_X1 U9961 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  INV_X1 U9962 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9965) );
  XOR2_X1 U9963 ( .A(n8467), .B(n9965), .Z(n8477) );
  INV_X1 U9964 ( .A(n8477), .ZN(n8474) );
  INV_X1 U9965 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8472) );
  AOI21_X1 U9966 ( .B1(n8470), .B2(n8469), .A(n8468), .ZN(n8471) );
  XOR2_X1 U9967 ( .A(n8472), .B(n8471), .Z(n8476) );
  NAND2_X1 U9968 ( .A1(n8476), .A2(n9804), .ZN(n8473) );
  OAI211_X1 U9969 ( .C1(n8474), .C2(n9736), .A(n9734), .B(n8473), .ZN(n8479)
         );
  OAI22_X1 U9970 ( .A1(n8477), .A2(n9736), .B1(n8476), .B2(n8475), .ZN(n8478)
         );
  MUX2_X1 U9971 ( .A(n8479), .B(n8478), .S(n7982), .Z(n8480) );
  INV_X1 U9972 ( .A(n8480), .ZN(n8482) );
  OAI211_X1 U9973 ( .C1(n8484), .C2(n8483), .A(n8482), .B(n8481), .ZN(P2_U3264) );
  NAND2_X1 U9974 ( .A1(n9584), .A2(n8490), .ZN(n8485) );
  XNOR2_X1 U9975 ( .A(n9579), .B(n8485), .ZN(n9581) );
  NAND2_X1 U9976 ( .A1(n9581), .A2(n8716), .ZN(n8489) );
  NAND2_X1 U9977 ( .A1(n8487), .A2(n8486), .ZN(n9583) );
  NOR2_X1 U9978 ( .A1(n8713), .A2(n9583), .ZN(n8492) );
  AOI21_X1 U9979 ( .B1(n8713), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8492), .ZN(
        n8488) );
  OAI211_X1 U9980 ( .C1(n9579), .C2(n8704), .A(n8489), .B(n8488), .ZN(P2_U3265) );
  XNOR2_X1 U9981 ( .A(n8491), .B(n8490), .ZN(n9586) );
  NAND2_X1 U9982 ( .A1(n9586), .A2(n8716), .ZN(n8494) );
  AOI21_X1 U9983 ( .B1(n8713), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8492), .ZN(
        n8493) );
  OAI211_X1 U9984 ( .C1(n9584), .C2(n8704), .A(n8494), .B(n8493), .ZN(P2_U3266) );
  XOR2_X1 U9985 ( .A(n8501), .B(n8495), .Z(n8734) );
  AOI21_X1 U9986 ( .B1(n8730), .B2(n8513), .A(n8496), .ZN(n8731) );
  INV_X1 U9987 ( .A(n8730), .ZN(n8499) );
  AOI22_X1 U9988 ( .A1(n8713), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8497), .B2(
        n9834), .ZN(n8498) );
  OAI21_X1 U9989 ( .B1(n8499), .B2(n8704), .A(n8498), .ZN(n8505) );
  XOR2_X1 U9990 ( .A(n8501), .B(n8500), .Z(n8503) );
  AOI222_X1 U9991 ( .A1(n9816), .A2(n8503), .B1(n8502), .B2(n9821), .C1(n4484), 
        .C2(n9818), .ZN(n8733) );
  NOR2_X1 U9992 ( .A1(n8733), .A2(n8713), .ZN(n8504) );
  AOI211_X1 U9993 ( .C1(n8716), .C2(n8731), .A(n8505), .B(n8504), .ZN(n8506)
         );
  OAI21_X1 U9994 ( .B1(n8734), .B2(n8718), .A(n8506), .ZN(P2_U3269) );
  XNOR2_X1 U9995 ( .A(n8508), .B(n8507), .ZN(n8739) );
  XNOR2_X1 U9996 ( .A(n8510), .B(n8509), .ZN(n8512) );
  OAI21_X1 U9997 ( .B1(n8512), .B2(n8605), .A(n8511), .ZN(n8735) );
  AOI211_X1 U9998 ( .C1(n8737), .C2(n8522), .A(n9915), .B(n4577), .ZN(n8736)
         );
  NAND2_X1 U9999 ( .A1(n8736), .A2(n8681), .ZN(n8516) );
  AOI22_X1 U10000 ( .A1(n8713), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8514), .B2(
        n9834), .ZN(n8515) );
  OAI211_X1 U10001 ( .C1(n8517), .C2(n8704), .A(n8516), .B(n8515), .ZN(n8518)
         );
  AOI21_X1 U10002 ( .B1(n8735), .B2(n9838), .A(n8518), .ZN(n8519) );
  OAI21_X1 U10003 ( .B1(n8739), .B2(n8718), .A(n8519), .ZN(P2_U3270) );
  XNOR2_X1 U10004 ( .A(n8521), .B(n8520), .ZN(n8744) );
  INV_X1 U10005 ( .A(n8541), .ZN(n8524) );
  INV_X1 U10006 ( .A(n8522), .ZN(n8523) );
  AOI211_X1 U10007 ( .C1(n8741), .C2(n8524), .A(n9915), .B(n8523), .ZN(n8740)
         );
  INV_X1 U10008 ( .A(n8525), .ZN(n8526) );
  AOI22_X1 U10009 ( .A1(n8713), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8526), .B2(
        n9834), .ZN(n8527) );
  OAI21_X1 U10010 ( .B1(n4486), .B2(n8704), .A(n8527), .ZN(n8536) );
  INV_X1 U10011 ( .A(n8528), .ZN(n8529) );
  NOR2_X1 U10012 ( .A1(n8530), .A2(n8529), .ZN(n8532) );
  AOI211_X1 U10013 ( .C1(n8532), .C2(n8548), .A(n8605), .B(n8531), .ZN(n8534)
         );
  NOR2_X1 U10014 ( .A1(n8534), .A2(n8533), .ZN(n8743) );
  NOR2_X1 U10015 ( .A1(n8743), .A2(n8713), .ZN(n8535) );
  AOI211_X1 U10016 ( .C1(n8681), .C2(n8740), .A(n8536), .B(n8535), .ZN(n8537)
         );
  OAI21_X1 U10017 ( .B1(n8744), .B2(n8718), .A(n8537), .ZN(P2_U3271) );
  AOI21_X1 U10018 ( .B1(n8540), .B2(n8539), .A(n8538), .ZN(n8749) );
  INV_X1 U10019 ( .A(n8567), .ZN(n8542) );
  AOI21_X1 U10020 ( .B1(n8745), .B2(n8542), .A(n8541), .ZN(n8746) );
  INV_X1 U10021 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8543) );
  OAI22_X1 U10022 ( .A1(n8544), .A2(n8704), .B1(n8543), .B2(n9838), .ZN(n8556)
         );
  NAND2_X1 U10023 ( .A1(n8546), .A2(n8545), .ZN(n8547) );
  NAND3_X1 U10024 ( .A1(n8548), .A2(n9816), .A3(n8547), .ZN(n8552) );
  AOI22_X1 U10025 ( .A1(n8550), .A2(n9818), .B1(n9821), .B2(n8549), .ZN(n8551)
         );
  AND2_X1 U10026 ( .A1(n8552), .A2(n8551), .ZN(n8748) );
  NAND2_X1 U10027 ( .A1(n8553), .A2(n9834), .ZN(n8554) );
  AOI21_X1 U10028 ( .B1(n8748), .B2(n8554), .A(n8713), .ZN(n8555) );
  AOI211_X1 U10029 ( .C1(n8746), .C2(n8716), .A(n8556), .B(n8555), .ZN(n8557)
         );
  OAI21_X1 U10030 ( .B1(n8749), .B2(n8718), .A(n8557), .ZN(P2_U3272) );
  INV_X1 U10031 ( .A(n8576), .ZN(n8559) );
  OAI21_X1 U10032 ( .B1(n8559), .B2(n8558), .A(n8564), .ZN(n8561) );
  NAND2_X1 U10033 ( .A1(n8561), .A2(n8560), .ZN(n8563) );
  AOI222_X1 U10034 ( .A1(n9816), .A2(n8563), .B1(n8596), .B2(n9821), .C1(n8562), .C2(n9818), .ZN(n8755) );
  OR2_X1 U10035 ( .A1(n8565), .A2(n8564), .ZN(n8751) );
  NAND3_X1 U10036 ( .A1(n8751), .A2(n8750), .A3(n8566), .ZN(n8574) );
  AOI21_X1 U10037 ( .B1(n8752), .B2(n8581), .A(n8567), .ZN(n8753) );
  INV_X1 U10038 ( .A(n8568), .ZN(n8569) );
  AOI22_X1 U10039 ( .A1(n8713), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8569), .B2(
        n9834), .ZN(n8570) );
  OAI21_X1 U10040 ( .B1(n8571), .B2(n8704), .A(n8570), .ZN(n8572) );
  AOI21_X1 U10041 ( .B1(n8753), .B2(n8716), .A(n8572), .ZN(n8573) );
  OAI211_X1 U10042 ( .C1(n8713), .C2(n8755), .A(n8574), .B(n8573), .ZN(
        P2_U3273) );
  XNOR2_X1 U10043 ( .A(n8575), .B(n8578), .ZN(n8761) );
  OAI211_X1 U10044 ( .C1(n8578), .C2(n8577), .A(n8576), .B(n9816), .ZN(n8580)
         );
  NAND2_X1 U10045 ( .A1(n8580), .A2(n8579), .ZN(n8757) );
  AOI211_X1 U10046 ( .C1(n8759), .C2(n8589), .A(n9915), .B(n4592), .ZN(n8758)
         );
  NAND2_X1 U10047 ( .A1(n8758), .A2(n8681), .ZN(n8584) );
  AOI22_X1 U10048 ( .A1(n8713), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8582), .B2(
        n9834), .ZN(n8583) );
  OAI211_X1 U10049 ( .C1(n8585), .C2(n8704), .A(n8584), .B(n8583), .ZN(n8586)
         );
  AOI21_X1 U10050 ( .B1(n8757), .B2(n9838), .A(n8586), .ZN(n8587) );
  OAI21_X1 U10051 ( .B1(n8761), .B2(n8718), .A(n8587), .ZN(P2_U3274) );
  XOR2_X1 U10052 ( .A(n8588), .B(n8594), .Z(n8766) );
  INV_X1 U10053 ( .A(n8609), .ZN(n8590) );
  AOI21_X1 U10054 ( .B1(n8762), .B2(n8590), .A(n4593), .ZN(n8763) );
  AOI22_X1 U10055 ( .A1(n8713), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8591), .B2(
        n9834), .ZN(n8592) );
  OAI21_X1 U10056 ( .B1(n8593), .B2(n8704), .A(n8592), .ZN(n8599) );
  XNOR2_X1 U10057 ( .A(n8595), .B(n8594), .ZN(n8597) );
  AOI222_X1 U10058 ( .A1(n9816), .A2(n8597), .B1(n8596), .B2(n9818), .C1(n8625), .C2(n9821), .ZN(n8765) );
  NOR2_X1 U10059 ( .A1(n8765), .A2(n8713), .ZN(n8598) );
  AOI211_X1 U10060 ( .C1(n8763), .C2(n8716), .A(n8599), .B(n8598), .ZN(n8600)
         );
  OAI21_X1 U10061 ( .B1(n8766), .B2(n8718), .A(n8600), .ZN(P2_U3275) );
  XNOR2_X1 U10062 ( .A(n8601), .B(n8603), .ZN(n8771) );
  NAND2_X1 U10063 ( .A1(n8622), .A2(n8602), .ZN(n8604) );
  XNOR2_X1 U10064 ( .A(n8604), .B(n8603), .ZN(n8606) );
  OAI222_X1 U10065 ( .A1(n8662), .A2(n8608), .B1(n8664), .B2(n8607), .C1(n8606), .C2(n8605), .ZN(n8767) );
  INV_X1 U10066 ( .A(n8619), .ZN(n8610) );
  AOI211_X1 U10067 ( .C1(n8769), .C2(n8610), .A(n9915), .B(n8609), .ZN(n8768)
         );
  NAND2_X1 U10068 ( .A1(n8768), .A2(n8681), .ZN(n8614) );
  INV_X1 U10069 ( .A(n8611), .ZN(n8612) );
  AOI22_X1 U10070 ( .A1(n8713), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8612), .B2(
        n9834), .ZN(n8613) );
  OAI211_X1 U10071 ( .C1(n8615), .C2(n8704), .A(n8614), .B(n8613), .ZN(n8616)
         );
  AOI21_X1 U10072 ( .B1(n8767), .B2(n9838), .A(n8616), .ZN(n8617) );
  OAI21_X1 U10073 ( .B1(n8771), .B2(n8718), .A(n8617), .ZN(P2_U3276) );
  XOR2_X1 U10074 ( .A(n8618), .B(n8624), .Z(n8776) );
  AOI211_X1 U10075 ( .C1(n8773), .C2(n8631), .A(n9915), .B(n8619), .ZN(n8772)
         );
  AOI22_X1 U10076 ( .A1(n8713), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8620), .B2(
        n9834), .ZN(n8621) );
  OAI21_X1 U10077 ( .B1(n4597), .B2(n8704), .A(n8621), .ZN(n8628) );
  OAI21_X1 U10078 ( .B1(n8624), .B2(n8623), .A(n8622), .ZN(n8626) );
  AOI222_X1 U10079 ( .A1(n9816), .A2(n8626), .B1(n8625), .B2(n9818), .C1(n8649), .C2(n9821), .ZN(n8775) );
  NOR2_X1 U10080 ( .A1(n8775), .A2(n8713), .ZN(n8627) );
  AOI211_X1 U10081 ( .C1(n8772), .C2(n8681), .A(n8628), .B(n8627), .ZN(n8629)
         );
  OAI21_X1 U10082 ( .B1(n8776), .B2(n8718), .A(n8629), .ZN(P2_U3277) );
  XNOR2_X1 U10083 ( .A(n8630), .B(n4338), .ZN(n8781) );
  INV_X1 U10084 ( .A(n8631), .ZN(n8632) );
  AOI21_X1 U10085 ( .B1(n8777), .B2(n8652), .A(n8632), .ZN(n8778) );
  AOI22_X1 U10086 ( .A1(n8713), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8633), .B2(
        n9834), .ZN(n8634) );
  OAI21_X1 U10087 ( .B1(n8635), .B2(n8704), .A(n8634), .ZN(n8641) );
  OAI21_X1 U10088 ( .B1(n4390), .B2(n4338), .A(n8636), .ZN(n8639) );
  AOI222_X1 U10089 ( .A1(n9816), .A2(n8639), .B1(n8638), .B2(n9818), .C1(n8637), .C2(n9821), .ZN(n8780) );
  NOR2_X1 U10090 ( .A1(n8780), .A2(n8713), .ZN(n8640) );
  AOI211_X1 U10091 ( .C1(n8778), .C2(n8716), .A(n8641), .B(n8640), .ZN(n8642)
         );
  OAI21_X1 U10092 ( .B1(n8781), .B2(n8718), .A(n8642), .ZN(P2_U3278) );
  OAI21_X1 U10093 ( .B1(n4394), .B2(n8644), .A(n8643), .ZN(n8645) );
  INV_X1 U10094 ( .A(n8645), .ZN(n8786) );
  OAI211_X1 U10095 ( .C1(n8648), .C2(n8647), .A(n8646), .B(n9816), .ZN(n8651)
         );
  AOI22_X1 U10096 ( .A1(n8649), .A2(n9818), .B1(n8693), .B2(n9821), .ZN(n8650)
         );
  NAND2_X1 U10097 ( .A1(n8651), .A2(n8650), .ZN(n8782) );
  INV_X1 U10098 ( .A(n8674), .ZN(n8654) );
  INV_X1 U10099 ( .A(n8652), .ZN(n8653) );
  AOI211_X1 U10100 ( .C1(n8784), .C2(n8654), .A(n9915), .B(n8653), .ZN(n8783)
         );
  NAND2_X1 U10101 ( .A1(n8783), .A2(n8681), .ZN(n8657) );
  AOI22_X1 U10102 ( .A1(n8713), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8655), .B2(
        n9834), .ZN(n8656) );
  OAI211_X1 U10103 ( .C1(n8658), .C2(n8704), .A(n8657), .B(n8656), .ZN(n8659)
         );
  AOI21_X1 U10104 ( .B1(n8782), .B2(n9838), .A(n8659), .ZN(n8660) );
  OAI21_X1 U10105 ( .B1(n8786), .B2(n8718), .A(n8660), .ZN(P2_U3279) );
  XNOR2_X1 U10106 ( .A(n8661), .B(n8666), .ZN(n8673) );
  OAI22_X1 U10107 ( .A1(n8665), .A2(n8664), .B1(n8663), .B2(n8662), .ZN(n8672)
         );
  AND2_X1 U10108 ( .A1(n8667), .A2(n8666), .ZN(n8668) );
  NOR2_X1 U10109 ( .A1(n8791), .A2(n8670), .ZN(n8671) );
  AOI211_X1 U10110 ( .C1(n9816), .C2(n8673), .A(n8672), .B(n8671), .ZN(n8790)
         );
  AOI211_X1 U10111 ( .C1(n8788), .C2(n8687), .A(n9915), .B(n8674), .ZN(n8787)
         );
  INV_X1 U10112 ( .A(n8788), .ZN(n8677) );
  AOI22_X1 U10113 ( .A1(n8713), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8675), .B2(
        n9834), .ZN(n8676) );
  OAI21_X1 U10114 ( .B1(n8677), .B2(n8704), .A(n8676), .ZN(n8680) );
  NOR2_X1 U10115 ( .A1(n8791), .A2(n8678), .ZN(n8679) );
  AOI211_X1 U10116 ( .C1(n8787), .C2(n8681), .A(n8680), .B(n8679), .ZN(n8682)
         );
  OAI21_X1 U10117 ( .B1(n8790), .B2(n8713), .A(n8682), .ZN(P2_U3280) );
  OAI21_X1 U10118 ( .B1(n8685), .B2(n8684), .A(n8683), .ZN(n8686) );
  INV_X1 U10119 ( .A(n8686), .ZN(n8796) );
  INV_X1 U10120 ( .A(n8687), .ZN(n8688) );
  AOI21_X1 U10121 ( .B1(n8792), .B2(n8700), .A(n8688), .ZN(n8793) );
  AOI22_X1 U10122 ( .A1(n8713), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8689), .B2(
        n9834), .ZN(n8690) );
  OAI21_X1 U10123 ( .B1(n4581), .B2(n8704), .A(n8690), .ZN(n8696) );
  XNOR2_X1 U10124 ( .A(n8691), .B(n4462), .ZN(n8694) );
  AOI222_X1 U10125 ( .A1(n9816), .A2(n8694), .B1(n8693), .B2(n9818), .C1(n8692), .C2(n9821), .ZN(n8795) );
  NOR2_X1 U10126 ( .A1(n8795), .A2(n8713), .ZN(n8695) );
  AOI211_X1 U10127 ( .C1(n8793), .C2(n8716), .A(n8696), .B(n8695), .ZN(n8697)
         );
  OAI21_X1 U10128 ( .B1(n8796), .B2(n8718), .A(n8697), .ZN(P2_U3281) );
  XNOR2_X1 U10129 ( .A(n8699), .B(n8698), .ZN(n8801) );
  AOI21_X1 U10130 ( .B1(n8797), .B2(n8701), .A(n4582), .ZN(n8798) );
  AOI22_X1 U10131 ( .A1(n8713), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8702), .B2(
        n9834), .ZN(n8703) );
  OAI21_X1 U10132 ( .B1(n8705), .B2(n8704), .A(n8703), .ZN(n8715) );
  NAND2_X1 U10133 ( .A1(n8707), .A2(n8706), .ZN(n8709) );
  XNOR2_X1 U10134 ( .A(n8709), .B(n8708), .ZN(n8712) );
  AOI222_X1 U10135 ( .A1(n9816), .A2(n8712), .B1(n8711), .B2(n9821), .C1(n8710), .C2(n9818), .ZN(n8800) );
  NOR2_X1 U10136 ( .A1(n8800), .A2(n8713), .ZN(n8714) );
  AOI211_X1 U10137 ( .C1(n8798), .C2(n8716), .A(n8715), .B(n8714), .ZN(n8717)
         );
  OAI21_X1 U10138 ( .B1(n8718), .B2(n8801), .A(n8717), .ZN(P2_U3282) );
  AOI22_X1 U10139 ( .A1(n8725), .A2(n9827), .B1(n8804), .B2(n8724), .ZN(n8726)
         );
  NAND2_X1 U10140 ( .A1(n8729), .A2(n8728), .ZN(n8810) );
  MUX2_X1 U10141 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8810), .S(n9934), .Z(
        P2_U3548) );
  AOI22_X1 U10142 ( .A1(n8731), .A2(n9827), .B1(n8804), .B2(n8730), .ZN(n8732)
         );
  OAI211_X1 U10143 ( .C1(n8734), .C2(n9877), .A(n8733), .B(n8732), .ZN(n8811)
         );
  MUX2_X1 U10144 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8811), .S(n9934), .Z(
        P2_U3547) );
  AOI211_X1 U10145 ( .C1(n8804), .C2(n8737), .A(n8736), .B(n8735), .ZN(n8738)
         );
  OAI21_X1 U10146 ( .B1(n8739), .B2(n9877), .A(n8738), .ZN(n8812) );
  MUX2_X1 U10147 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8812), .S(n9934), .Z(
        P2_U3546) );
  AOI21_X1 U10148 ( .B1(n8804), .B2(n8741), .A(n8740), .ZN(n8742) );
  OAI211_X1 U10149 ( .C1(n8744), .C2(n9877), .A(n8743), .B(n8742), .ZN(n8813)
         );
  MUX2_X1 U10150 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8813), .S(n9934), .Z(
        P2_U3545) );
  AOI22_X1 U10151 ( .A1(n8746), .A2(n9827), .B1(n8804), .B2(n8745), .ZN(n8747)
         );
  OAI211_X1 U10152 ( .C1(n8749), .C2(n9877), .A(n8748), .B(n8747), .ZN(n8814)
         );
  MUX2_X1 U10153 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8814), .S(n9934), .Z(
        P2_U3544) );
  NAND3_X1 U10154 ( .A1(n8751), .A2(n8750), .A3(n9919), .ZN(n8756) );
  AOI22_X1 U10155 ( .A1(n8753), .A2(n9827), .B1(n8804), .B2(n8752), .ZN(n8754)
         );
  NAND3_X1 U10156 ( .A1(n8756), .A2(n8755), .A3(n8754), .ZN(n8815) );
  MUX2_X1 U10157 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8815), .S(n9934), .Z(
        P2_U3543) );
  AOI211_X1 U10158 ( .C1(n8804), .C2(n8759), .A(n8758), .B(n8757), .ZN(n8760)
         );
  OAI21_X1 U10159 ( .B1(n8761), .B2(n9877), .A(n8760), .ZN(n8816) );
  MUX2_X1 U10160 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8816), .S(n9934), .Z(
        P2_U3542) );
  AOI22_X1 U10161 ( .A1(n8763), .A2(n9827), .B1(n8804), .B2(n8762), .ZN(n8764)
         );
  OAI211_X1 U10162 ( .C1(n8766), .C2(n9877), .A(n8765), .B(n8764), .ZN(n8817)
         );
  MUX2_X1 U10163 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8817), .S(n9934), .Z(
        P2_U3541) );
  AOI211_X1 U10164 ( .C1(n8804), .C2(n8769), .A(n8768), .B(n8767), .ZN(n8770)
         );
  OAI21_X1 U10165 ( .B1(n8771), .B2(n9877), .A(n8770), .ZN(n8818) );
  MUX2_X1 U10166 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8818), .S(n9934), .Z(
        P2_U3540) );
  AOI21_X1 U10167 ( .B1(n8804), .B2(n8773), .A(n8772), .ZN(n8774) );
  OAI211_X1 U10168 ( .C1(n8776), .C2(n9877), .A(n8775), .B(n8774), .ZN(n8819)
         );
  MUX2_X1 U10169 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8819), .S(n9934), .Z(
        P2_U3539) );
  AOI22_X1 U10170 ( .A1(n8778), .A2(n9827), .B1(n8804), .B2(n8777), .ZN(n8779)
         );
  OAI211_X1 U10171 ( .C1(n8781), .C2(n9877), .A(n8780), .B(n8779), .ZN(n8820)
         );
  MUX2_X1 U10172 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8820), .S(n9934), .Z(
        P2_U3538) );
  AOI211_X1 U10173 ( .C1(n8804), .C2(n8784), .A(n8783), .B(n8782), .ZN(n8785)
         );
  OAI21_X1 U10174 ( .B1(n8786), .B2(n9877), .A(n8785), .ZN(n8821) );
  MUX2_X1 U10175 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8821), .S(n9934), .Z(
        P2_U3537) );
  AOI21_X1 U10176 ( .B1(n8804), .B2(n8788), .A(n8787), .ZN(n8789) );
  OAI211_X1 U10177 ( .C1(n9905), .C2(n8791), .A(n8790), .B(n8789), .ZN(n8822)
         );
  MUX2_X1 U10178 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8822), .S(n9934), .Z(
        P2_U3536) );
  AOI22_X1 U10179 ( .A1(n8793), .A2(n9827), .B1(n8804), .B2(n8792), .ZN(n8794)
         );
  OAI211_X1 U10180 ( .C1(n8796), .C2(n9877), .A(n8795), .B(n8794), .ZN(n8823)
         );
  MUX2_X1 U10181 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8823), .S(n9934), .Z(
        P2_U3535) );
  AOI22_X1 U10182 ( .A1(n8798), .A2(n9827), .B1(n8804), .B2(n8797), .ZN(n8799)
         );
  OAI211_X1 U10183 ( .C1(n8801), .C2(n9877), .A(n8800), .B(n8799), .ZN(n8824)
         );
  MUX2_X1 U10184 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8824), .S(n9934), .Z(
        P2_U3534) );
  INV_X1 U10185 ( .A(n8802), .ZN(n8808) );
  AOI22_X1 U10186 ( .A1(n8805), .A2(n9827), .B1(n8804), .B2(n8803), .ZN(n8806)
         );
  OAI211_X1 U10187 ( .C1(n9905), .C2(n8808), .A(n8807), .B(n8806), .ZN(n8825)
         );
  MUX2_X1 U10188 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8825), .S(n9934), .Z(
        P2_U3533) );
  MUX2_X1 U10189 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8810), .S(n9923), .Z(
        P2_U3516) );
  MUX2_X1 U10190 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8811), .S(n9923), .Z(
        P2_U3515) );
  MUX2_X1 U10191 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8812), .S(n9923), .Z(
        P2_U3514) );
  MUX2_X1 U10192 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8813), .S(n9923), .Z(
        P2_U3513) );
  MUX2_X1 U10193 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8814), .S(n9923), .Z(
        P2_U3512) );
  MUX2_X1 U10194 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8815), .S(n9923), .Z(
        P2_U3511) );
  MUX2_X1 U10195 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8816), .S(n9923), .Z(
        P2_U3510) );
  MUX2_X1 U10196 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8817), .S(n9923), .Z(
        P2_U3509) );
  MUX2_X1 U10197 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8818), .S(n9923), .Z(
        P2_U3508) );
  MUX2_X1 U10198 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8819), .S(n9923), .Z(
        P2_U3507) );
  MUX2_X1 U10199 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8820), .S(n9923), .Z(
        P2_U3505) );
  MUX2_X1 U10200 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8821), .S(n9923), .Z(
        P2_U3502) );
  MUX2_X1 U10201 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8822), .S(n9923), .Z(
        P2_U3499) );
  MUX2_X1 U10202 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8823), .S(n9923), .Z(
        P2_U3496) );
  MUX2_X1 U10203 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8824), .S(n9923), .Z(
        P2_U3493) );
  MUX2_X1 U10204 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8825), .S(n9923), .Z(
        P2_U3490) );
  NOR4_X1 U10205 ( .A1(n4323), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8826), .A4(
        P2_U3152), .ZN(n8827) );
  AOI21_X1 U10206 ( .B1(n8828), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8827), .ZN(
        n8829) );
  OAI21_X1 U10207 ( .B1(n9540), .B2(n8830), .A(n8829), .ZN(P2_U3327) );
  INV_X1 U10208 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8832) );
  OAI222_X1 U10209 ( .A1(n8830), .A2(n8834), .B1(P2_U3152), .B2(n8833), .C1(
        n8832), .C2(n8831), .ZN(P2_U3329) );
  MUX2_X1 U10210 ( .A(n8835), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10211 ( .A1(n8837), .A2(n8836), .ZN(n8838) );
  XOR2_X1 U10212 ( .A(n8839), .B(n8838), .Z(n8846) );
  NOR2_X1 U10213 ( .A1(n9648), .A2(n9384), .ZN(n8844) );
  NAND2_X1 U10214 ( .A1(n9306), .A2(n9083), .ZN(n8841) );
  NAND2_X1 U10215 ( .A1(n9304), .A2(n9078), .ZN(n8840) );
  AND2_X1 U10216 ( .A1(n8841), .A2(n8840), .ZN(n9382) );
  OAI21_X1 U10217 ( .B1(n8884), .B2(n9382), .A(n8842), .ZN(n8843) );
  AOI211_X1 U10218 ( .C1(n8970), .C2(n9387), .A(n8844), .B(n8843), .ZN(n8845)
         );
  OAI21_X1 U10219 ( .B1(n8846), .B2(n8972), .A(n8845), .ZN(P1_U3213) );
  XNOR2_X1 U10220 ( .A(n8848), .B(n8847), .ZN(n8849) );
  XNOR2_X1 U10221 ( .A(n8850), .B(n8849), .ZN(n8857) );
  INV_X1 U10222 ( .A(n9273), .ZN(n8976) );
  AOI22_X1 U10223 ( .A1(n8967), .A2(n8976), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8853) );
  INV_X1 U10224 ( .A(n8851), .ZN(n9231) );
  NAND2_X1 U10225 ( .A1(n8930), .A2(n9231), .ZN(n8852) );
  OAI211_X1 U10226 ( .C1(n8854), .C2(n8964), .A(n8853), .B(n8852), .ZN(n8855)
         );
  AOI21_X1 U10227 ( .B1(n9446), .B2(n8970), .A(n8855), .ZN(n8856) );
  OAI21_X1 U10228 ( .B1(n8857), .B2(n8972), .A(n8856), .ZN(P1_U3214) );
  INV_X1 U10229 ( .A(n9467), .ZN(n9298) );
  OAI21_X1 U10230 ( .B1(n8860), .B2(n8859), .A(n8858), .ZN(n8861) );
  NAND2_X1 U10231 ( .A1(n8861), .A2(n9643), .ZN(n8866) );
  INV_X1 U10232 ( .A(n8862), .ZN(n9296) );
  INV_X1 U10233 ( .A(n8902), .ZN(n9305) );
  NOR2_X1 U10234 ( .A1(n10120), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9064) );
  AOI21_X1 U10235 ( .B1(n8967), .B2(n9305), .A(n9064), .ZN(n8863) );
  OAI21_X1 U10236 ( .B1(n9092), .B2(n8964), .A(n8863), .ZN(n8864) );
  AOI21_X1 U10237 ( .B1(n9296), .B2(n8930), .A(n8864), .ZN(n8865) );
  OAI211_X1 U10238 ( .C1(n9298), .C2(n8959), .A(n8866), .B(n8865), .ZN(
        P1_U3217) );
  NAND2_X1 U10239 ( .A1(n4909), .A2(n8868), .ZN(n8869) );
  XNOR2_X1 U10240 ( .A(n8867), .B(n8869), .ZN(n8874) );
  NOR2_X1 U10241 ( .A1(n9648), .A2(n9264), .ZN(n8872) );
  AOI22_X1 U10242 ( .A1(n8967), .A2(n9307), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8870) );
  OAI21_X1 U10243 ( .B1(n9273), .B2(n8964), .A(n8870), .ZN(n8871) );
  AOI211_X1 U10244 ( .C1(n9458), .C2(n8970), .A(n8872), .B(n8871), .ZN(n8873)
         );
  OAI21_X1 U10245 ( .B1(n8874), .B2(n8972), .A(n8873), .ZN(P1_U3221) );
  INV_X1 U10246 ( .A(n8875), .ZN(n8879) );
  NOR3_X1 U10247 ( .A1(n4351), .A2(n8877), .A3(n8876), .ZN(n8878) );
  OAI21_X1 U10248 ( .B1(n8879), .B2(n8878), .A(n9643), .ZN(n8888) );
  INV_X1 U10249 ( .A(n8880), .ZN(n9201) );
  NAND2_X1 U10250 ( .A1(n9103), .A2(n9306), .ZN(n8882) );
  NAND2_X1 U10251 ( .A1(n9239), .A2(n9304), .ZN(n8881) );
  NAND2_X1 U10252 ( .A1(n8882), .A2(n8881), .ZN(n9206) );
  INV_X1 U10253 ( .A(n9206), .ZN(n8885) );
  OAI22_X1 U10254 ( .A1(n8885), .A2(n8884), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8883), .ZN(n8886) );
  AOI21_X1 U10255 ( .B1(n9201), .B2(n8930), .A(n8886), .ZN(n8887) );
  OAI211_X1 U10256 ( .C1(n9203), .C2(n8959), .A(n8888), .B(n8887), .ZN(
        P1_U3223) );
  NOR2_X1 U10257 ( .A1(n4398), .A2(n8889), .ZN(n8890) );
  XNOR2_X1 U10258 ( .A(n8891), .B(n8890), .ZN(n8897) );
  OR2_X1 U10259 ( .A1(n9323), .A2(n9556), .ZN(n8893) );
  NAND2_X1 U10260 ( .A1(n9304), .A2(n9083), .ZN(n8892) );
  NAND2_X1 U10261 ( .A1(n8893), .A2(n8892), .ZN(n9357) );
  AOI22_X1 U10262 ( .A1(n9633), .A2(n9357), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8894) );
  OAI21_X1 U10263 ( .B1(n9351), .B2(n9648), .A(n8894), .ZN(n8895) );
  AOI21_X1 U10264 ( .B1(n9481), .B2(n8970), .A(n8895), .ZN(n8896) );
  OAI21_X1 U10265 ( .B1(n8897), .B2(n8972), .A(n8896), .ZN(P1_U3224) );
  NAND2_X1 U10266 ( .A1(n8900), .A2(n8899), .ZN(n8901) );
  XNOR2_X1 U10267 ( .A(n8898), .B(n8901), .ZN(n8906) );
  OAI22_X1 U10268 ( .A1(n9552), .A2(n9363), .B1(n8902), .B2(n9556), .ZN(n9341)
         );
  AOI22_X1 U10269 ( .A1(n9633), .A2(n9341), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n8903) );
  OAI21_X1 U10270 ( .B1(n9335), .B2(n9648), .A(n8903), .ZN(n8904) );
  AOI21_X1 U10271 ( .B1(n9476), .B2(n8970), .A(n8904), .ZN(n8905) );
  OAI21_X1 U10272 ( .B1(n8906), .B2(n8972), .A(n8905), .ZN(P1_U3226) );
  AOI21_X1 U10273 ( .B1(n8908), .B2(n8907), .A(n4351), .ZN(n8915) );
  NAND2_X1 U10274 ( .A1(n9225), .A2(n9712), .ZN(n9439) );
  INV_X1 U10275 ( .A(n9439), .ZN(n8913) );
  AND2_X1 U10276 ( .A1(n9256), .A2(n9304), .ZN(n8909) );
  AOI21_X1 U10277 ( .B1(n8975), .B2(n9306), .A(n8909), .ZN(n9440) );
  INV_X1 U10278 ( .A(n9440), .ZN(n8910) );
  AOI22_X1 U10279 ( .A1(n8910), .A2(n9633), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8911) );
  OAI21_X1 U10280 ( .B1(n9214), .B2(n9648), .A(n8911), .ZN(n8912) );
  AOI21_X1 U10281 ( .B1(n8913), .B2(n9642), .A(n8912), .ZN(n8914) );
  OAI21_X1 U10282 ( .B1(n8915), .B2(n8972), .A(n8914), .ZN(P1_U3227) );
  NAND2_X1 U10283 ( .A1(n4910), .A2(n8917), .ZN(n8918) );
  XNOR2_X1 U10284 ( .A(n8916), .B(n8918), .ZN(n8925) );
  INV_X1 U10285 ( .A(n9282), .ZN(n8922) );
  NAND2_X1 U10286 ( .A1(n9304), .A2(n9090), .ZN(n8919) );
  OAI21_X1 U10287 ( .B1(n8920), .B2(n9556), .A(n8919), .ZN(n9287) );
  AOI22_X1 U10288 ( .A1(n9633), .A2(n9287), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8921) );
  OAI21_X1 U10289 ( .B1(n8922), .B2(n9648), .A(n8921), .ZN(n8923) );
  AOI21_X1 U10290 ( .B1(n9461), .B2(n8970), .A(n8923), .ZN(n8924) );
  OAI21_X1 U10291 ( .B1(n8925), .B2(n8972), .A(n8924), .ZN(P1_U3231) );
  INV_X1 U10292 ( .A(n8926), .ZN(n8929) );
  XNOR2_X1 U10293 ( .A(n8927), .B(n4340), .ZN(n8928) );
  XNOR2_X1 U10294 ( .A(n8929), .B(n8928), .ZN(n8936) );
  AOI22_X1 U10295 ( .A1(n8967), .A2(n9255), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8932) );
  NAND2_X1 U10296 ( .A1(n8930), .A2(n9247), .ZN(n8931) );
  OAI211_X1 U10297 ( .C1(n8933), .C2(n8964), .A(n8932), .B(n8931), .ZN(n8934)
         );
  AOI21_X1 U10298 ( .B1(n9452), .B2(n8970), .A(n8934), .ZN(n8935) );
  OAI21_X1 U10299 ( .B1(n8936), .B2(n8972), .A(n8935), .ZN(P1_U3233) );
  XOR2_X1 U10300 ( .A(n8938), .B(n8937), .Z(n8939) );
  XNOR2_X1 U10301 ( .A(n8940), .B(n8939), .ZN(n8945) );
  INV_X1 U10302 ( .A(n9323), .ZN(n9088) );
  NAND2_X1 U10303 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9037) );
  OAI21_X1 U10304 ( .B1(n8964), .B2(n9322), .A(n9037), .ZN(n8941) );
  AOI21_X1 U10305 ( .B1(n8967), .B2(n9088), .A(n8941), .ZN(n8942) );
  OAI21_X1 U10306 ( .B1(n9326), .B2(n9648), .A(n8942), .ZN(n8943) );
  AOI21_X1 U10307 ( .B1(n9472), .B2(n8970), .A(n8943), .ZN(n8944) );
  OAI21_X1 U10308 ( .B1(n8945), .B2(n8972), .A(n8944), .ZN(P1_U3236) );
  OR2_X1 U10309 ( .A1(n8951), .A2(n9556), .ZN(n8953) );
  NAND2_X1 U10310 ( .A1(n8975), .A2(n9304), .ZN(n8952) );
  NAND2_X1 U10311 ( .A1(n8953), .A2(n8952), .ZN(n9192) );
  INV_X1 U10312 ( .A(n9187), .ZN(n8955) );
  OAI22_X1 U10313 ( .A1(n8955), .A2(n9648), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8954), .ZN(n8956) );
  AOI21_X1 U10314 ( .B1(n9192), .B2(n9633), .A(n8956), .ZN(n8957) );
  OAI211_X1 U10315 ( .C1(n9189), .C2(n8959), .A(n8958), .B(n8957), .ZN(
        P1_U3238) );
  XOR2_X1 U10316 ( .A(n8961), .B(n8960), .Z(n8962) );
  XNOR2_X1 U10317 ( .A(n8963), .B(n8962), .ZN(n8973) );
  INV_X1 U10318 ( .A(n9364), .ZN(n9081) );
  NOR2_X1 U10319 ( .A1(n8964), .A2(n9363), .ZN(n8965) );
  AOI211_X1 U10320 ( .C1(n8967), .C2(n9081), .A(n8966), .B(n8965), .ZN(n8968)
         );
  OAI21_X1 U10321 ( .B1(n9369), .B2(n9648), .A(n8968), .ZN(n8969) );
  AOI21_X1 U10322 ( .B1(n8970), .B2(n9488), .A(n8969), .ZN(n8971) );
  OAI21_X1 U10323 ( .B1(n8973), .B2(n8972), .A(n8971), .ZN(P1_U3239) );
  MUX2_X1 U10324 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9140), .S(n8986), .Z(
        P1_U3585) );
  MUX2_X1 U10325 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8974), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10326 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9108), .S(n8986), .Z(
        P1_U3583) );
  MUX2_X1 U10327 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9106), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10328 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9103), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10329 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8975), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10330 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9239), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10331 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9256), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10332 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n8976), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10333 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9255), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10334 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9307), .S(n8986), .Z(
        P1_U3575) );
  MUX2_X1 U10335 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9090), .S(n8986), .Z(
        P1_U3574) );
  MUX2_X1 U10336 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9305), .S(n8986), .Z(
        P1_U3573) );
  MUX2_X1 U10337 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9088), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10338 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9085), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10339 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9083), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10340 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9081), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10341 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9078), .S(P1_U4006), .Z(
        P1_U3568) );
  INV_X1 U10342 ( .A(n8977), .ZN(n9077) );
  MUX2_X1 U10343 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9077), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10344 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9073), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10345 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8978), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10346 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8979), .S(n8986), .Z(
        P1_U3564) );
  MUX2_X1 U10347 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8980), .S(n8986), .Z(
        P1_U3563) );
  MUX2_X1 U10348 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8981), .S(n8986), .Z(
        P1_U3562) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8982), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10350 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8983), .S(n8986), .Z(
        P1_U3560) );
  MUX2_X1 U10351 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8984), .S(n8986), .Z(
        P1_U3559) );
  MUX2_X1 U10352 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8985), .S(n8986), .Z(
        P1_U3558) );
  MUX2_X1 U10353 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5838), .S(n8986), .Z(
        P1_U3557) );
  MUX2_X1 U10354 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5823), .S(n8986), .Z(
        P1_U3556) );
  MUX2_X1 U10355 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n8987), .S(n8986), .Z(
        P1_U3555) );
  AND3_X1 U10356 ( .A1(n8990), .A2(n8989), .A3(n8988), .ZN(n8991) );
  NOR3_X1 U10357 ( .A1(n10162), .A2(n8992), .A3(n8991), .ZN(n8993) );
  AOI21_X1 U10358 ( .B1(n9036), .B2(n8994), .A(n8993), .ZN(n9001) );
  NOR2_X1 U10359 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5419), .ZN(n8995) );
  AOI21_X1 U10360 ( .B1(n9658), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n8995), .ZN(
        n9000) );
  OAI211_X1 U10361 ( .C1(n8998), .C2(n8997), .A(n9651), .B(n8996), .ZN(n8999)
         );
  NAND3_X1 U10362 ( .A1(n9001), .A2(n9000), .A3(n8999), .ZN(P1_U3244) );
  INV_X1 U10363 ( .A(n9002), .ZN(n9007) );
  OAI21_X1 U10364 ( .B1(n9005), .B2(n9004), .A(n9003), .ZN(n9006) );
  AOI22_X1 U10365 ( .A1(n9036), .A2(n9007), .B1(n9660), .B2(n9006), .ZN(n9015)
         );
  AOI21_X1 U10366 ( .B1(n9010), .B2(n9009), .A(n9008), .ZN(n9011) );
  NOR2_X1 U10367 ( .A1(n10154), .A2(n9011), .ZN(n9012) );
  AOI211_X1 U10368 ( .C1(n9658), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9013), .B(
        n9012), .ZN(n9014) );
  NAND3_X1 U10369 ( .A1(n9016), .A2(n9015), .A3(n9014), .ZN(P1_U3245) );
  XNOR2_X1 U10370 ( .A(n9018), .B(n9017), .ZN(n9030) );
  INV_X1 U10371 ( .A(n9019), .ZN(n9020) );
  AOI211_X1 U10372 ( .C1(n9022), .C2(n9021), .A(n10154), .B(n9020), .ZN(n9028)
         );
  NOR2_X1 U10373 ( .A1(n10163), .A2(n9023), .ZN(n9027) );
  NOR2_X1 U10374 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9964), .ZN(n9026) );
  INV_X1 U10375 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9024) );
  NOR2_X1 U10376 ( .A1(n10167), .A2(n9024), .ZN(n9025) );
  NOR4_X1 U10377 ( .A1(n9028), .A2(n9027), .A3(n9026), .A4(n9025), .ZN(n9029)
         );
  OAI21_X1 U10378 ( .B1(n10162), .B2(n9030), .A(n9029), .ZN(P1_U3257) );
  AOI22_X1 U10379 ( .A1(n9033), .A2(n9032), .B1(P1_REG1_REG_17__SCAN_IN), .B2(
        n9031), .ZN(n9035) );
  NOR2_X1 U10380 ( .A1(n9051), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9047) );
  AOI21_X1 U10381 ( .B1(n9051), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9047), .ZN(
        n9034) );
  NAND2_X1 U10382 ( .A1(n9035), .A2(n9034), .ZN(n9049) );
  OAI21_X1 U10383 ( .B1(n9035), .B2(n9034), .A(n9049), .ZN(n9040) );
  INV_X1 U10384 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10180) );
  NAND2_X1 U10385 ( .A1(n9036), .A2(n9051), .ZN(n9038) );
  OAI211_X1 U10386 ( .C1(n10180), .C2(n10167), .A(n9038), .B(n9037), .ZN(n9039) );
  AOI21_X1 U10387 ( .B1(n9040), .B2(n9660), .A(n9039), .ZN(n9046) );
  NAND2_X1 U10388 ( .A1(n9042), .A2(n9041), .ZN(n9044) );
  MUX2_X1 U10389 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9316), .S(n9051), .Z(n9043) );
  NAND2_X1 U10390 ( .A1(n9044), .A2(n9043), .ZN(n9053) );
  OAI211_X1 U10391 ( .C1(n9044), .C2(n9043), .A(n9053), .B(n9651), .ZN(n9045)
         );
  NAND2_X1 U10392 ( .A1(n9046), .A2(n9045), .ZN(P1_U3259) );
  INV_X1 U10393 ( .A(n9047), .ZN(n9048) );
  NAND2_X1 U10394 ( .A1(n9049), .A2(n9048), .ZN(n9050) );
  XNOR2_X1 U10395 ( .A(n9050), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U10396 ( .A1(n9051), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U10397 ( .A1(n9053), .A2(n9052), .ZN(n9054) );
  XNOR2_X1 U10398 ( .A(n9054), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9059) );
  INV_X1 U10399 ( .A(n9059), .ZN(n9055) );
  AOI22_X1 U10400 ( .A1(n9057), .A2(n9660), .B1(n9055), .B2(n9651), .ZN(n9063)
         );
  INV_X1 U10401 ( .A(n9056), .ZN(n9060) );
  OAI21_X1 U10402 ( .B1(n9057), .B2(n10162), .A(n10163), .ZN(n9058) );
  AOI21_X1 U10403 ( .B1(n9060), .B2(n9059), .A(n9058), .ZN(n9062) );
  MUX2_X1 U10404 ( .A(n9063), .B(n9062), .S(n9061), .Z(n9066) );
  INV_X1 U10405 ( .A(n9064), .ZN(n9065) );
  OAI211_X1 U10406 ( .C1(n4809), .C2(n10167), .A(n9066), .B(n9065), .ZN(
        P1_U3260) );
  INV_X1 U10407 ( .A(n9412), .ZN(n9072) );
  INV_X1 U10408 ( .A(n9143), .ZN(n9067) );
  NOR2_X1 U10409 ( .A1(n9067), .A2(n9072), .ZN(n9410) );
  OR3_X1 U10410 ( .A1(n9410), .A2(n9409), .A3(n9389), .ZN(n9071) );
  AND2_X1 U10411 ( .A1(n9605), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9068) );
  NOR2_X1 U10412 ( .A1(n9069), .A2(n9068), .ZN(n9070) );
  OAI211_X1 U10413 ( .C1(n9072), .C2(n9401), .A(n9071), .B(n9070), .ZN(
        P1_U3262) );
  NOR2_X1 U10414 ( .A1(n9074), .A2(n9073), .ZN(n9075) );
  AND2_X1 U10415 ( .A1(n9612), .A2(n9078), .ZN(n9080) );
  OR2_X1 U10416 ( .A1(n9612), .A2(n9078), .ZN(n9079) );
  NOR2_X1 U10417 ( .A1(n9387), .A2(n9081), .ZN(n9082) );
  NOR2_X1 U10418 ( .A1(n9467), .A2(n9090), .ZN(n9091) );
  NAND2_X1 U10419 ( .A1(n9458), .A2(n9255), .ZN(n9093) );
  NAND2_X1 U10420 ( .A1(n9249), .A2(n9273), .ZN(n9095) );
  NOR2_X1 U10421 ( .A1(n9249), .A2(n9273), .ZN(n9094) );
  NAND2_X1 U10422 ( .A1(n9203), .A2(n9100), .ZN(n9183) );
  OR2_X1 U10423 ( .A1(n9430), .A2(n9103), .ZN(n9101) );
  AND2_X1 U10424 ( .A1(n9183), .A2(n9101), .ZN(n9102) );
  NAND2_X1 U10425 ( .A1(n9430), .A2(n9103), .ZN(n9104) );
  NAND2_X1 U10426 ( .A1(n9105), .A2(n9104), .ZN(n9166) );
  INV_X1 U10427 ( .A(n9420), .ZN(n9157) );
  INV_X1 U10428 ( .A(n9414), .ZN(n9150) );
  NAND2_X1 U10429 ( .A1(n9494), .A2(n9110), .ZN(n9112) );
  NAND2_X1 U10430 ( .A1(n9112), .A2(n9111), .ZN(n9395) );
  NAND2_X1 U10431 ( .A1(n9395), .A2(n9399), .ZN(n9394) );
  NOR2_X1 U10432 ( .A1(n9380), .A2(n9113), .ZN(n9114) );
  NAND2_X1 U10433 ( .A1(n9394), .A2(n9114), .ZN(n9116) );
  NAND2_X1 U10434 ( .A1(n9340), .A2(n9120), .ZN(n9122) );
  NAND2_X1 U10435 ( .A1(n9122), .A2(n9121), .ZN(n9320) );
  INV_X1 U10436 ( .A(n9313), .ZN(n9321) );
  NOR2_X1 U10437 ( .A1(n9300), .A2(n9301), .ZN(n9123) );
  NAND2_X1 U10438 ( .A1(n9288), .A2(n9125), .ZN(n9269) );
  INV_X1 U10439 ( .A(n9262), .ZN(n9270) );
  NOR2_X1 U10440 ( .A1(n9250), .A2(n9251), .ZN(n9126) );
  INV_X1 U10441 ( .A(n9130), .ZN(n9132) );
  NOR3_X1 U10442 ( .A1(n9172), .A2(n9158), .A3(n9135), .ZN(n9138) );
  INV_X1 U10443 ( .A(n9136), .ZN(n9137) );
  NOR2_X1 U10444 ( .A1(n9138), .A2(n9137), .ZN(n9139) );
  AOI22_X1 U10445 ( .A1(n9108), .A2(n9304), .B1(n9141), .B2(n9140), .ZN(n9142)
         );
  AOI22_X1 U10446 ( .A1(n9145), .A2(n9594), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9377), .ZN(n9147) );
  NAND2_X1 U10447 ( .A1(n9417), .A2(n9595), .ZN(n9146) );
  OAI211_X1 U10448 ( .C1(n9415), .C2(n9389), .A(n9147), .B(n9146), .ZN(n9148)
         );
  AOI21_X1 U10449 ( .B1(n9416), .B2(n9327), .A(n9148), .ZN(n9149) );
  OAI21_X1 U10450 ( .B1(n9150), .B2(n9392), .A(n9149), .ZN(P1_U3355) );
  NAND2_X1 U10451 ( .A1(n9152), .A2(n9159), .ZN(n9153) );
  AOI211_X1 U10452 ( .C1(n9420), .C2(n9167), .A(n9704), .B(n9154), .ZN(n9419)
         );
  AOI22_X1 U10453 ( .A1(n9155), .A2(n9594), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9377), .ZN(n9156) );
  OAI21_X1 U10454 ( .B1(n9157), .B2(n9401), .A(n9156), .ZN(n9164) );
  NOR2_X1 U10455 ( .A1(n9172), .A2(n9158), .ZN(n9160) );
  XNOR2_X1 U10456 ( .A(n9160), .B(n9159), .ZN(n9162) );
  AOI21_X2 U10457 ( .B1(n9162), .B2(n9501), .A(n9161), .ZN(n9422) );
  NOR2_X1 U10458 ( .A1(n9422), .A2(n9605), .ZN(n9163) );
  AOI211_X1 U10459 ( .C1(n9419), .C2(n9599), .A(n9164), .B(n9163), .ZN(n9165)
         );
  OAI21_X1 U10460 ( .B1(n9423), .B2(n9392), .A(n9165), .ZN(P1_U3263) );
  XNOR2_X1 U10461 ( .A(n9166), .B(n9174), .ZN(n9428) );
  INV_X1 U10462 ( .A(n9167), .ZN(n9168) );
  AOI21_X1 U10463 ( .B1(n9424), .B2(n9185), .A(n9168), .ZN(n9425) );
  AOI22_X1 U10464 ( .A1(n9169), .A2(n9594), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9377), .ZN(n9170) );
  OAI21_X1 U10465 ( .B1(n9171), .B2(n9401), .A(n9170), .ZN(n9180) );
  AOI211_X1 U10466 ( .C1(n9174), .C2(n9173), .A(n9553), .B(n9172), .ZN(n9178)
         );
  OAI22_X1 U10467 ( .A1(n9176), .A2(n9556), .B1(n9175), .B2(n9552), .ZN(n9177)
         );
  NOR2_X1 U10468 ( .A1(n9178), .A2(n9177), .ZN(n9427) );
  NOR2_X1 U10469 ( .A1(n9427), .A2(n9605), .ZN(n9179) );
  AOI211_X1 U10470 ( .C1(n9566), .C2(n9425), .A(n9180), .B(n9179), .ZN(n9181)
         );
  OAI21_X1 U10471 ( .B1(n9428), .B2(n9392), .A(n9181), .ZN(P1_U3264) );
  NAND2_X1 U10472 ( .A1(n9182), .A2(n9183), .ZN(n9184) );
  XOR2_X1 U10473 ( .A(n9190), .B(n9184), .Z(n9433) );
  INV_X1 U10474 ( .A(n9199), .ZN(n9186) );
  AOI211_X1 U10475 ( .C1(n9430), .C2(n9186), .A(n9704), .B(n4538), .ZN(n9429)
         );
  AOI22_X1 U10476 ( .A1(n9187), .A2(n9594), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9605), .ZN(n9188) );
  OAI21_X1 U10477 ( .B1(n9189), .B2(n9401), .A(n9188), .ZN(n9195) );
  XNOR2_X1 U10478 ( .A(n9191), .B(n9190), .ZN(n9193) );
  NOR2_X1 U10479 ( .A1(n9432), .A2(n9377), .ZN(n9194) );
  AOI211_X1 U10480 ( .C1(n9429), .C2(n9599), .A(n9195), .B(n9194), .ZN(n9196)
         );
  OAI21_X1 U10481 ( .B1(n9433), .B2(n9392), .A(n9196), .ZN(P1_U3265) );
  INV_X1 U10482 ( .A(n9182), .ZN(n9198) );
  AOI21_X1 U10483 ( .B1(n9205), .B2(n9197), .A(n9198), .ZN(n9438) );
  INV_X1 U10484 ( .A(n9212), .ZN(n9200) );
  AOI21_X1 U10485 ( .B1(n9434), .B2(n9200), .A(n9199), .ZN(n9435) );
  AOI22_X1 U10486 ( .A1(n9201), .A2(n9594), .B1(n9605), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n9202) );
  OAI21_X1 U10487 ( .B1(n9203), .B2(n9401), .A(n9202), .ZN(n9209) );
  XNOR2_X1 U10488 ( .A(n9204), .B(n9205), .ZN(n9207) );
  AOI21_X1 U10489 ( .B1(n9207), .B2(n9501), .A(n9206), .ZN(n9437) );
  NOR2_X1 U10490 ( .A1(n9437), .A2(n9605), .ZN(n9208) );
  AOI211_X1 U10491 ( .C1(n9435), .C2(n9566), .A(n9209), .B(n9208), .ZN(n9210)
         );
  OAI21_X1 U10492 ( .B1(n9438), .B2(n9392), .A(n9210), .ZN(P1_U3266) );
  NAND2_X1 U10493 ( .A1(n9230), .A2(n9225), .ZN(n9211) );
  NAND2_X1 U10494 ( .A1(n9211), .A2(n9713), .ZN(n9213) );
  OR2_X1 U10495 ( .A1(n9213), .A2(n9212), .ZN(n9441) );
  INV_X1 U10496 ( .A(n9441), .ZN(n9221) );
  OAI21_X1 U10497 ( .B1(n9214), .B2(n9559), .A(n9440), .ZN(n9220) );
  NAND3_X1 U10498 ( .A1(n9215), .A2(n9222), .A3(n9216), .ZN(n9217) );
  NAND2_X1 U10499 ( .A1(n9217), .A2(n9501), .ZN(n9218) );
  NOR2_X1 U10500 ( .A1(n9219), .A2(n9218), .ZN(n9443) );
  AOI211_X1 U10501 ( .C1(n9221), .C2(n9274), .A(n9220), .B(n9443), .ZN(n9228)
         );
  XOR2_X1 U10502 ( .A(n9223), .B(n9222), .Z(n9444) );
  NAND2_X1 U10503 ( .A1(n9444), .A2(n9224), .ZN(n9227) );
  AOI22_X1 U10504 ( .A1(n9225), .A2(n9595), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9377), .ZN(n9226) );
  OAI211_X1 U10505 ( .C1(n9605), .C2(n9228), .A(n9227), .B(n9226), .ZN(
        P1_U3267) );
  XNOR2_X1 U10506 ( .A(n9229), .B(n9128), .ZN(n9450) );
  AOI21_X1 U10507 ( .B1(n9446), .B2(n9244), .A(n4543), .ZN(n9447) );
  INV_X1 U10508 ( .A(n9446), .ZN(n9233) );
  AOI22_X1 U10509 ( .A1(n9377), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9231), .B2(
        n9594), .ZN(n9232) );
  OAI21_X1 U10510 ( .B1(n9233), .B2(n9401), .A(n9232), .ZN(n9241) );
  NOR2_X1 U10511 ( .A1(n9273), .A2(n9552), .ZN(n9238) );
  INV_X1 U10512 ( .A(n9215), .ZN(n9234) );
  AOI211_X1 U10513 ( .C1(n9236), .C2(n9235), .A(n9553), .B(n9234), .ZN(n9237)
         );
  AOI211_X1 U10514 ( .C1(n9306), .C2(n9239), .A(n9238), .B(n9237), .ZN(n9449)
         );
  NOR2_X1 U10515 ( .A1(n9449), .A2(n9605), .ZN(n9240) );
  AOI211_X1 U10516 ( .C1(n9447), .C2(n9566), .A(n9241), .B(n9240), .ZN(n9242)
         );
  OAI21_X1 U10517 ( .B1(n9450), .B2(n9392), .A(n9242), .ZN(P1_U3268) );
  XNOR2_X1 U10518 ( .A(n9243), .B(n9250), .ZN(n9455) );
  INV_X1 U10519 ( .A(n9266), .ZN(n9246) );
  INV_X1 U10520 ( .A(n9244), .ZN(n9245) );
  AOI211_X1 U10521 ( .C1(n9452), .C2(n9246), .A(n9704), .B(n9245), .ZN(n9451)
         );
  AOI22_X1 U10522 ( .A1(n9377), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9247), .B2(
        n9594), .ZN(n9248) );
  OAI21_X1 U10523 ( .B1(n9249), .B2(n9401), .A(n9248), .ZN(n9259) );
  INV_X1 U10524 ( .A(n9268), .ZN(n9252) );
  OAI21_X1 U10525 ( .B1(n9252), .B2(n9251), .A(n9250), .ZN(n9254) );
  NAND2_X1 U10526 ( .A1(n9254), .A2(n9253), .ZN(n9257) );
  AOI222_X1 U10527 ( .A1(n9501), .A2(n9257), .B1(n9256), .B2(n9306), .C1(n9255), .C2(n9304), .ZN(n9454) );
  NOR2_X1 U10528 ( .A1(n9454), .A2(n9605), .ZN(n9258) );
  AOI211_X1 U10529 ( .C1(n9451), .C2(n9599), .A(n9259), .B(n9258), .ZN(n9260)
         );
  OAI21_X1 U10530 ( .B1(n9455), .B2(n9392), .A(n9260), .ZN(P1_U3269) );
  OAI21_X1 U10531 ( .B1(n9263), .B2(n9262), .A(n9261), .ZN(n9460) );
  INV_X1 U10532 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9265) );
  OAI22_X1 U10533 ( .A1(n9327), .A2(n9265), .B1(n9264), .B2(n9559), .ZN(n9277)
         );
  INV_X1 U10534 ( .A(n9280), .ZN(n9267) );
  AOI211_X1 U10535 ( .C1(n9458), .C2(n9267), .A(n9704), .B(n9266), .ZN(n9457)
         );
  OAI211_X1 U10536 ( .C1(n9270), .C2(n9269), .A(n9268), .B(n9501), .ZN(n9272)
         );
  NAND2_X1 U10537 ( .A1(n9304), .A2(n9307), .ZN(n9271) );
  OAI211_X1 U10538 ( .C1(n9273), .C2(n9556), .A(n9272), .B(n9271), .ZN(n9456)
         );
  AOI21_X1 U10539 ( .B1(n9457), .B2(n9274), .A(n9456), .ZN(n9275) );
  NOR2_X1 U10540 ( .A1(n9275), .A2(n9377), .ZN(n9276) );
  AOI211_X1 U10541 ( .C1(n9595), .C2(n9458), .A(n9277), .B(n9276), .ZN(n9278)
         );
  OAI21_X1 U10542 ( .B1(n9460), .B2(n9392), .A(n9278), .ZN(P1_U3270) );
  XNOR2_X1 U10543 ( .A(n9279), .B(n9285), .ZN(n9465) );
  INV_X1 U10544 ( .A(n9295), .ZN(n9281) );
  AOI21_X1 U10545 ( .B1(n9461), .B2(n9281), .A(n9280), .ZN(n9462) );
  AOI22_X1 U10546 ( .A1(n9377), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9282), .B2(
        n9594), .ZN(n9283) );
  OAI21_X1 U10547 ( .B1(n9284), .B2(n9401), .A(n9283), .ZN(n9291) );
  AOI21_X1 U10548 ( .B1(n9286), .B2(n9285), .A(n9553), .ZN(n9289) );
  AOI21_X1 U10549 ( .B1(n9289), .B2(n9288), .A(n9287), .ZN(n9464) );
  NOR2_X1 U10550 ( .A1(n9464), .A2(n9377), .ZN(n9290) );
  AOI211_X1 U10551 ( .C1(n9462), .C2(n9566), .A(n9291), .B(n9290), .ZN(n9292)
         );
  OAI21_X1 U10552 ( .B1(n9465), .B2(n9392), .A(n9292), .ZN(P1_U3271) );
  XNOR2_X1 U10553 ( .A(n9294), .B(n9293), .ZN(n9470) );
  AOI211_X1 U10554 ( .C1(n9467), .C2(n9315), .A(n9704), .B(n9295), .ZN(n9466)
         );
  AOI22_X1 U10555 ( .A1(n9377), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9296), .B2(
        n9594), .ZN(n9297) );
  OAI21_X1 U10556 ( .B1(n9298), .B2(n9401), .A(n9297), .ZN(n9310) );
  INV_X1 U10557 ( .A(n9299), .ZN(n9319) );
  OAI21_X1 U10558 ( .B1(n9319), .B2(n9301), .A(n9300), .ZN(n9303) );
  NAND2_X1 U10559 ( .A1(n9303), .A2(n9302), .ZN(n9308) );
  AOI222_X1 U10560 ( .A1(n9501), .A2(n9308), .B1(n9307), .B2(n9306), .C1(n9305), .C2(n9304), .ZN(n9469) );
  NOR2_X1 U10561 ( .A1(n9469), .A2(n9605), .ZN(n9309) );
  AOI211_X1 U10562 ( .C1(n9466), .C2(n9599), .A(n9310), .B(n9309), .ZN(n9311)
         );
  OAI21_X1 U10563 ( .B1(n9470), .B2(n9392), .A(n9311), .ZN(P1_U3272) );
  AOI21_X1 U10564 ( .B1(n9313), .B2(n9312), .A(n4391), .ZN(n9314) );
  INV_X1 U10565 ( .A(n9314), .ZN(n9475) );
  AOI211_X1 U10566 ( .C1(n9472), .C2(n9333), .A(n9704), .B(n4537), .ZN(n9471)
         );
  INV_X1 U10567 ( .A(n9472), .ZN(n9317) );
  OAI22_X1 U10568 ( .A1(n9317), .A2(n9401), .B1(n9316), .B2(n9327), .ZN(n9318)
         );
  AOI21_X1 U10569 ( .B1(n9471), .B2(n9599), .A(n9318), .ZN(n9330) );
  AOI211_X1 U10570 ( .C1(n9321), .C2(n9320), .A(n9553), .B(n9319), .ZN(n9325)
         );
  OAI22_X1 U10571 ( .A1(n9552), .A2(n9323), .B1(n9322), .B2(n9556), .ZN(n9324)
         );
  NOR2_X1 U10572 ( .A1(n9325), .A2(n9324), .ZN(n9474) );
  OAI21_X1 U10573 ( .B1(n9326), .B2(n9559), .A(n9474), .ZN(n9328) );
  NAND2_X1 U10574 ( .A1(n9328), .A2(n9327), .ZN(n9329) );
  OAI211_X1 U10575 ( .C1(n9475), .C2(n9392), .A(n9330), .B(n9329), .ZN(
        P1_U3273) );
  XNOR2_X1 U10576 ( .A(n9332), .B(n9339), .ZN(n9480) );
  INV_X1 U10577 ( .A(n9333), .ZN(n9334) );
  AOI21_X1 U10578 ( .B1(n9476), .B2(n9348), .A(n9334), .ZN(n9477) );
  INV_X1 U10579 ( .A(n9335), .ZN(n9336) );
  AOI22_X1 U10580 ( .A1(n9377), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9336), .B2(
        n9594), .ZN(n9337) );
  OAI21_X1 U10581 ( .B1(n9338), .B2(n9401), .A(n9337), .ZN(n9344) );
  XNOR2_X1 U10582 ( .A(n9340), .B(n9339), .ZN(n9342) );
  AOI21_X1 U10583 ( .B1(n9342), .B2(n9501), .A(n9341), .ZN(n9479) );
  NOR2_X1 U10584 ( .A1(n9479), .A2(n9377), .ZN(n9343) );
  AOI211_X1 U10585 ( .C1(n9477), .C2(n9566), .A(n9344), .B(n9343), .ZN(n9345)
         );
  OAI21_X1 U10586 ( .B1(n9480), .B2(n9392), .A(n9345), .ZN(P1_U3274) );
  XNOR2_X1 U10587 ( .A(n9346), .B(n9355), .ZN(n9486) );
  INV_X1 U10588 ( .A(n9347), .ZN(n9350) );
  INV_X1 U10589 ( .A(n9348), .ZN(n9349) );
  AOI21_X1 U10590 ( .B1(n9481), .B2(n9350), .A(n9349), .ZN(n9482) );
  INV_X1 U10591 ( .A(n9351), .ZN(n9352) );
  AOI22_X1 U10592 ( .A1(n9377), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9352), .B2(
        n9594), .ZN(n9353) );
  OAI21_X1 U10593 ( .B1(n9354), .B2(n9401), .A(n9353), .ZN(n9360) );
  XNOR2_X1 U10594 ( .A(n9356), .B(n9355), .ZN(n9358) );
  AOI21_X1 U10595 ( .B1(n9358), .B2(n9501), .A(n9357), .ZN(n9484) );
  NOR2_X1 U10596 ( .A1(n9484), .A2(n9377), .ZN(n9359) );
  AOI211_X1 U10597 ( .C1(n9482), .C2(n9566), .A(n9360), .B(n9359), .ZN(n9361)
         );
  OAI21_X1 U10598 ( .B1(n9486), .B2(n9392), .A(n9361), .ZN(P1_U3275) );
  XNOR2_X1 U10599 ( .A(n9362), .B(n4616), .ZN(n9368) );
  OAI22_X1 U10600 ( .A1(n9552), .A2(n9364), .B1(n9363), .B2(n9556), .ZN(n9367)
         );
  XNOR2_X1 U10601 ( .A(n9365), .B(n4616), .ZN(n9491) );
  NOR2_X1 U10602 ( .A1(n9491), .A2(n9497), .ZN(n9366) );
  AOI211_X1 U10603 ( .C1(n9501), .C2(n9368), .A(n9367), .B(n9366), .ZN(n9490)
         );
  AOI211_X1 U10604 ( .C1(n9488), .C2(n4339), .A(n9704), .B(n9347), .ZN(n9487)
         );
  INV_X1 U10605 ( .A(n9369), .ZN(n9370) );
  AOI22_X1 U10606 ( .A1(n9377), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9370), .B2(
        n9594), .ZN(n9371) );
  OAI21_X1 U10607 ( .B1(n9372), .B2(n9401), .A(n9371), .ZN(n9375) );
  NOR2_X1 U10608 ( .A1(n9491), .A2(n9373), .ZN(n9374) );
  AOI211_X1 U10609 ( .C1(n9487), .C2(n9599), .A(n9375), .B(n9374), .ZN(n9376)
         );
  OAI21_X1 U10610 ( .B1(n9490), .B2(n9377), .A(n9376), .ZN(P1_U3276) );
  XNOR2_X1 U10611 ( .A(n9378), .B(n9380), .ZN(n9610) );
  INV_X1 U10612 ( .A(n9610), .ZN(n9393) );
  NAND2_X1 U10613 ( .A1(n9394), .A2(n9379), .ZN(n9381) );
  XNOR2_X1 U10614 ( .A(n9381), .B(n9380), .ZN(n9383) );
  OAI21_X1 U10615 ( .B1(n9383), .B2(n9553), .A(n9382), .ZN(n9609) );
  INV_X1 U10616 ( .A(n9387), .ZN(n9606) );
  OAI21_X1 U10617 ( .B1(n9606), .B2(n4384), .A(n4339), .ZN(n9607) );
  OAI22_X1 U10618 ( .A1(n9327), .A2(n9385), .B1(n9384), .B2(n9559), .ZN(n9386)
         );
  AOI21_X1 U10619 ( .B1(n9387), .B2(n9595), .A(n9386), .ZN(n9388) );
  OAI21_X1 U10620 ( .B1(n9607), .B2(n9389), .A(n9388), .ZN(n9390) );
  AOI21_X1 U10621 ( .B1(n9609), .B2(n9327), .A(n9390), .ZN(n9391) );
  OAI21_X1 U10622 ( .B1(n9393), .B2(n9392), .A(n9391), .ZN(P1_U3277) );
  OAI21_X1 U10623 ( .B1(n9399), .B2(n9395), .A(n9394), .ZN(n9397) );
  AOI21_X1 U10624 ( .B1(n9397), .B2(n9501), .A(n9396), .ZN(n9614) );
  XOR2_X1 U10625 ( .A(n9399), .B(n9398), .Z(n9615) );
  INV_X1 U10626 ( .A(n9615), .ZN(n9617) );
  NAND2_X1 U10627 ( .A1(n9617), .A2(n9400), .ZN(n9408) );
  AOI211_X1 U10628 ( .C1(n9612), .C2(n9503), .A(n9704), .B(n4384), .ZN(n9611)
         );
  INV_X1 U10629 ( .A(n9612), .ZN(n9402) );
  NOR2_X1 U10630 ( .A1(n9402), .A2(n9401), .ZN(n9406) );
  OAI22_X1 U10631 ( .A1(n9327), .A2(n9404), .B1(n9403), .B2(n9559), .ZN(n9405)
         );
  AOI211_X1 U10632 ( .C1(n9611), .C2(n9599), .A(n9406), .B(n9405), .ZN(n9407)
         );
  OAI211_X1 U10633 ( .C1(n9605), .C2(n9614), .A(n9408), .B(n9407), .ZN(
        P1_U3278) );
  MUX2_X1 U10634 ( .A(n5086), .B(n9514), .S(n9733), .Z(n9413) );
  INV_X1 U10635 ( .A(n9413), .ZN(P1_U3553) );
  NAND2_X1 U10636 ( .A1(n9414), .A2(n9708), .ZN(n9418) );
  MUX2_X1 U10637 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9517), .S(n9733), .Z(
        P1_U3552) );
  AOI21_X1 U10638 ( .B1(n9712), .B2(n9420), .A(n9419), .ZN(n9421) );
  OAI211_X1 U10639 ( .C1(n9423), .C2(n9485), .A(n9422), .B(n9421), .ZN(n9518)
         );
  MUX2_X1 U10640 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9518), .S(n9733), .Z(
        P1_U3551) );
  AOI22_X1 U10641 ( .A1(n9425), .A2(n9713), .B1(n9712), .B2(n9424), .ZN(n9426)
         );
  OAI211_X1 U10642 ( .C1(n9428), .C2(n9485), .A(n9427), .B(n9426), .ZN(n9519)
         );
  MUX2_X1 U10643 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9519), .S(n9733), .Z(
        P1_U3550) );
  AOI21_X1 U10644 ( .B1(n9712), .B2(n9430), .A(n9429), .ZN(n9431) );
  OAI211_X1 U10645 ( .C1(n9433), .C2(n9485), .A(n9432), .B(n9431), .ZN(n9520)
         );
  MUX2_X1 U10646 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9520), .S(n9733), .Z(
        P1_U3549) );
  AOI22_X1 U10647 ( .A1(n9435), .A2(n9713), .B1(n9712), .B2(n9434), .ZN(n9436)
         );
  OAI211_X1 U10648 ( .C1(n9438), .C2(n9485), .A(n9437), .B(n9436), .ZN(n9521)
         );
  MUX2_X1 U10649 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9521), .S(n9733), .Z(
        P1_U3548) );
  NAND3_X1 U10650 ( .A1(n9441), .A2(n9440), .A3(n9439), .ZN(n9442) );
  AOI211_X1 U10651 ( .C1(n9444), .C2(n9708), .A(n9443), .B(n9442), .ZN(n9445)
         );
  INV_X1 U10652 ( .A(n9445), .ZN(n9522) );
  MUX2_X1 U10653 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9522), .S(n9733), .Z(
        P1_U3547) );
  AOI22_X1 U10654 ( .A1(n9447), .A2(n9713), .B1(n9712), .B2(n9446), .ZN(n9448)
         );
  OAI211_X1 U10655 ( .C1(n9450), .C2(n9485), .A(n9449), .B(n9448), .ZN(n9523)
         );
  MUX2_X1 U10656 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9523), .S(n9733), .Z(
        P1_U3546) );
  AOI21_X1 U10657 ( .B1(n9712), .B2(n9452), .A(n9451), .ZN(n9453) );
  OAI211_X1 U10658 ( .C1(n9455), .C2(n9485), .A(n9454), .B(n9453), .ZN(n9524)
         );
  MUX2_X1 U10659 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9524), .S(n9733), .Z(
        P1_U3545) );
  AOI211_X1 U10660 ( .C1(n9712), .C2(n9458), .A(n9457), .B(n9456), .ZN(n9459)
         );
  OAI21_X1 U10661 ( .B1(n9460), .B2(n9485), .A(n9459), .ZN(n9525) );
  MUX2_X1 U10662 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9525), .S(n9733), .Z(
        P1_U3544) );
  AOI22_X1 U10663 ( .A1(n9462), .A2(n9713), .B1(n9712), .B2(n9461), .ZN(n9463)
         );
  OAI211_X1 U10664 ( .C1(n9465), .C2(n9485), .A(n9464), .B(n9463), .ZN(n9526)
         );
  MUX2_X1 U10665 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9526), .S(n9733), .Z(
        P1_U3543) );
  AOI21_X1 U10666 ( .B1(n9712), .B2(n9467), .A(n9466), .ZN(n9468) );
  OAI211_X1 U10667 ( .C1(n9470), .C2(n9485), .A(n9469), .B(n9468), .ZN(n9527)
         );
  MUX2_X1 U10668 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9527), .S(n9733), .Z(
        P1_U3542) );
  AOI21_X1 U10669 ( .B1(n9712), .B2(n9472), .A(n9471), .ZN(n9473) );
  OAI211_X1 U10670 ( .C1(n9475), .C2(n9485), .A(n9474), .B(n9473), .ZN(n9528)
         );
  MUX2_X1 U10671 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9528), .S(n9733), .Z(
        P1_U3541) );
  AOI22_X1 U10672 ( .A1(n9477), .A2(n9713), .B1(n9712), .B2(n9476), .ZN(n9478)
         );
  OAI211_X1 U10673 ( .C1(n9480), .C2(n9485), .A(n9479), .B(n9478), .ZN(n9529)
         );
  MUX2_X1 U10674 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9529), .S(n9733), .Z(
        P1_U3540) );
  AOI22_X1 U10675 ( .A1(n9482), .A2(n9713), .B1(n9712), .B2(n9481), .ZN(n9483)
         );
  OAI211_X1 U10676 ( .C1(n9486), .C2(n9485), .A(n9484), .B(n9483), .ZN(n9530)
         );
  MUX2_X1 U10677 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9530), .S(n9733), .Z(
        P1_U3539) );
  AOI21_X1 U10678 ( .B1(n9712), .B2(n9488), .A(n9487), .ZN(n9489) );
  OAI211_X1 U10679 ( .C1(n9491), .C2(n9718), .A(n9490), .B(n9489), .ZN(n9531)
         );
  MUX2_X1 U10680 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9531), .S(n9733), .Z(
        P1_U3538) );
  XNOR2_X1 U10681 ( .A(n9492), .B(n9495), .ZN(n9597) );
  NAND2_X1 U10682 ( .A1(n9494), .A2(n9493), .ZN(n9496) );
  XNOR2_X1 U10683 ( .A(n9496), .B(n9495), .ZN(n9500) );
  NOR2_X1 U10684 ( .A1(n9597), .A2(n9497), .ZN(n9498) );
  AOI211_X1 U10685 ( .C1(n9501), .C2(n9500), .A(n9499), .B(n9498), .ZN(n9604)
         );
  INV_X1 U10686 ( .A(n9502), .ZN(n9505) );
  INV_X1 U10687 ( .A(n9503), .ZN(n9504) );
  AOI211_X1 U10688 ( .C1(n9596), .C2(n9505), .A(n9704), .B(n9504), .ZN(n9598)
         );
  AOI21_X1 U10689 ( .B1(n9712), .B2(n9596), .A(n9598), .ZN(n9506) );
  OAI211_X1 U10690 ( .C1(n9718), .C2(n9597), .A(n9604), .B(n9506), .ZN(n9532)
         );
  MUX2_X1 U10691 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9532), .S(n9733), .Z(
        P1_U3535) );
  INV_X1 U10692 ( .A(n9718), .ZN(n9680) );
  OAI22_X1 U10693 ( .A1(n9508), .A2(n9704), .B1(n9507), .B2(n9702), .ZN(n9509)
         );
  AOI21_X1 U10694 ( .B1(n9510), .B2(n9680), .A(n9509), .ZN(n9511) );
  NAND2_X1 U10695 ( .A1(n9512), .A2(n9511), .ZN(n9533) );
  MUX2_X1 U10696 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9533), .S(n9733), .Z(
        P1_U3534) );
  MUX2_X1 U10697 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9513), .S(n9733), .Z(
        P1_U3523) );
  INV_X1 U10698 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9515) );
  MUX2_X1 U10699 ( .A(n9515), .B(n9514), .S(n9724), .Z(n9516) );
  INV_X1 U10700 ( .A(n9516), .ZN(P1_U3521) );
  MUX2_X1 U10701 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9517), .S(n9724), .Z(
        P1_U3520) );
  MUX2_X1 U10702 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9518), .S(n9724), .Z(
        P1_U3519) );
  MUX2_X1 U10703 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9519), .S(n9724), .Z(
        P1_U3518) );
  MUX2_X1 U10704 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9520), .S(n9724), .Z(
        P1_U3517) );
  MUX2_X1 U10705 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9521), .S(n9724), .Z(
        P1_U3516) );
  MUX2_X1 U10706 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9522), .S(n9724), .Z(
        P1_U3515) );
  MUX2_X1 U10707 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9523), .S(n9724), .Z(
        P1_U3514) );
  MUX2_X1 U10708 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9524), .S(n9724), .Z(
        P1_U3513) );
  MUX2_X1 U10709 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9525), .S(n9724), .Z(
        P1_U3512) );
  MUX2_X1 U10710 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9526), .S(n9724), .Z(
        P1_U3511) );
  MUX2_X1 U10711 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9527), .S(n9724), .Z(
        P1_U3510) );
  MUX2_X1 U10712 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9528), .S(n9724), .Z(
        P1_U3508) );
  MUX2_X1 U10713 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9529), .S(n9724), .Z(
        P1_U3505) );
  MUX2_X1 U10714 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9530), .S(n9724), .Z(
        P1_U3502) );
  MUX2_X1 U10715 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9531), .S(n9724), .Z(
        P1_U3499) );
  MUX2_X1 U10716 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9532), .S(n9724), .Z(
        P1_U3490) );
  MUX2_X1 U10717 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9533), .S(n9724), .Z(
        P1_U3487) );
  MUX2_X1 U10718 ( .A(n9534), .B(P1_D_REG_0__SCAN_IN), .S(n9666), .Z(P1_U3440)
         );
  NOR4_X1 U10719 ( .A1(n4628), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9535), .ZN(n9536) );
  AOI21_X1 U10720 ( .B1(n9537), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9536), .ZN(
        n9538) );
  OAI21_X1 U10721 ( .B1(n9540), .B2(n9539), .A(n9538), .ZN(P1_U3322) );
  MUX2_X1 U10722 ( .A(n9542), .B(n9541), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  OR2_X1 U10723 ( .A1(n7736), .A2(n9543), .ZN(n9545) );
  NAND2_X1 U10724 ( .A1(n9545), .A2(n9544), .ZN(n9546) );
  XNOR2_X1 U10725 ( .A(n9546), .B(n9549), .ZN(n9574) );
  NAND2_X1 U10726 ( .A1(n9548), .A2(n9547), .ZN(n9550) );
  XNOR2_X1 U10727 ( .A(n9550), .B(n9549), .ZN(n9554) );
  OAI222_X1 U10728 ( .A1(n9556), .A2(n9555), .B1(n9554), .B2(n9553), .C1(n9552), .C2(n9551), .ZN(n9572) );
  AOI21_X1 U10729 ( .B1(n9574), .B2(n9721), .A(n9572), .ZN(n9569) );
  NAND2_X1 U10730 ( .A1(n9605), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9557) );
  OAI21_X1 U10731 ( .B1(n9559), .B2(n9558), .A(n9557), .ZN(n9560) );
  AOI21_X1 U10732 ( .B1(n9595), .B2(n9561), .A(n9560), .ZN(n9568) );
  INV_X1 U10733 ( .A(n9562), .ZN(n9563) );
  OAI21_X1 U10734 ( .B1(n9570), .B2(n9564), .A(n9563), .ZN(n9571) );
  INV_X1 U10735 ( .A(n9571), .ZN(n9565) );
  AOI22_X1 U10736 ( .A1(n9574), .A2(n9600), .B1(n9566), .B2(n9565), .ZN(n9567)
         );
  OAI211_X1 U10737 ( .C1(n9605), .C2(n9569), .A(n9568), .B(n9567), .ZN(
        P1_U3281) );
  OAI22_X1 U10738 ( .A1(n9571), .A2(n9704), .B1(n9570), .B2(n9702), .ZN(n9573)
         );
  AOI211_X1 U10739 ( .C1(n9574), .C2(n9708), .A(n9573), .B(n9572), .ZN(n9576)
         );
  INV_X1 U10740 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9575) );
  AOI22_X1 U10741 ( .A1(n9724), .A2(n9576), .B1(n9575), .B2(n9722), .ZN(
        P1_U3484) );
  AOI22_X1 U10742 ( .A1(n9733), .A2(n9576), .B1(n6568), .B2(n9731), .ZN(
        P1_U3533) );
  AOI22_X1 U10743 ( .A1(n9733), .A2(n9578), .B1(n9577), .B2(n9731), .ZN(
        P1_U3554) );
  OAI21_X1 U10744 ( .B1(n9579), .B2(n9914), .A(n9583), .ZN(n9580) );
  AOI21_X1 U10745 ( .B1(n9581), .B2(n9827), .A(n9580), .ZN(n9589) );
  INV_X1 U10746 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9582) );
  AOI22_X1 U10747 ( .A1(n9934), .A2(n9589), .B1(n9582), .B2(n9931), .ZN(
        P2_U3551) );
  OAI21_X1 U10748 ( .B1(n9584), .B2(n9914), .A(n9583), .ZN(n9585) );
  AOI21_X1 U10749 ( .B1(n9586), .B2(n9827), .A(n9585), .ZN(n9591) );
  INV_X1 U10750 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9587) );
  AOI22_X1 U10751 ( .A1(n9934), .A2(n9591), .B1(n9587), .B2(n9931), .ZN(
        P2_U3550) );
  INV_X1 U10752 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9588) );
  AOI22_X1 U10753 ( .A1(n9923), .A2(n9589), .B1(n9588), .B2(n9921), .ZN(
        P2_U3519) );
  INV_X1 U10754 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9590) );
  AOI22_X1 U10755 ( .A1(n9923), .A2(n9591), .B1(n9590), .B2(n9921), .ZN(
        P2_U3518) );
  INV_X1 U10756 ( .A(n9592), .ZN(n9593) );
  AOI222_X1 U10757 ( .A1(n9596), .A2(n9595), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9605), .C1(n9594), .C2(n9593), .ZN(n9603) );
  INV_X1 U10758 ( .A(n9597), .ZN(n9601) );
  AOI22_X1 U10759 ( .A1(n9601), .A2(n9600), .B1(n9599), .B2(n9598), .ZN(n9602)
         );
  OAI211_X1 U10760 ( .C1(n9605), .C2(n9604), .A(n9603), .B(n9602), .ZN(
        P1_U3279) );
  OAI22_X1 U10761 ( .A1(n9607), .A2(n9704), .B1(n9606), .B2(n9702), .ZN(n9608)
         );
  AOI211_X1 U10762 ( .C1(n9610), .C2(n9708), .A(n9609), .B(n9608), .ZN(n9619)
         );
  AOI22_X1 U10763 ( .A1(n9733), .A2(n9619), .B1(n5214), .B2(n9731), .ZN(
        P1_U3537) );
  AOI21_X1 U10764 ( .B1(n9712), .B2(n9612), .A(n9611), .ZN(n9613) );
  OAI211_X1 U10765 ( .C1(n9615), .C2(n9718), .A(n9614), .B(n9613), .ZN(n9616)
         );
  AOI21_X1 U10766 ( .B1(n9721), .B2(n9617), .A(n9616), .ZN(n9621) );
  AOI22_X1 U10767 ( .A1(n9733), .A2(n9621), .B1(n6704), .B2(n9731), .ZN(
        P1_U3536) );
  INV_X1 U10768 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9618) );
  AOI22_X1 U10769 ( .A1(n9724), .A2(n9619), .B1(n9618), .B2(n9722), .ZN(
        P1_U3496) );
  INV_X1 U10770 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U10771 ( .A1(n9724), .A2(n9621), .B1(n9620), .B2(n9722), .ZN(
        P1_U3493) );
  XNOR2_X1 U10772 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10773 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10774 ( .A(n9622), .ZN(n9623) );
  AOI22_X1 U10775 ( .A1(n9623), .A2(n9633), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3084), .ZN(n9630) );
  XNOR2_X1 U10776 ( .A(n9625), .B(n9624), .ZN(n9628) );
  NAND2_X1 U10777 ( .A1(n9626), .A2(n9712), .ZN(n9675) );
  INV_X1 U10778 ( .A(n9675), .ZN(n9627) );
  AOI22_X1 U10779 ( .A1(n9628), .A2(n9643), .B1(n9627), .B2(n9642), .ZN(n9629)
         );
  OAI211_X1 U10780 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9648), .A(n9630), .B(
        n9629), .ZN(P1_U3216) );
  INV_X1 U10781 ( .A(n9631), .ZN(n9634) );
  AOI21_X1 U10782 ( .B1(n9634), .B2(n9633), .A(n9632), .ZN(n9646) );
  OAI21_X1 U10783 ( .B1(n9636), .B2(n7318), .A(n9635), .ZN(n9640) );
  XNOR2_X1 U10784 ( .A(n9638), .B(n9637), .ZN(n9639) );
  XNOR2_X1 U10785 ( .A(n9640), .B(n9639), .ZN(n9644) );
  NOR2_X1 U10786 ( .A1(n9702), .A2(n9641), .ZN(n9688) );
  AOI22_X1 U10787 ( .A1(n9644), .A2(n9643), .B1(n9688), .B2(n9642), .ZN(n9645)
         );
  OAI211_X1 U10788 ( .C1(n9648), .C2(n9647), .A(n9646), .B(n9645), .ZN(
        P1_U3237) );
  NOR2_X1 U10789 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9649), .ZN(n9657) );
  OAI211_X1 U10790 ( .C1(n9653), .C2(n9652), .A(n9651), .B(n9650), .ZN(n9654)
         );
  OAI21_X1 U10791 ( .B1(n10163), .B2(n9655), .A(n9654), .ZN(n9656) );
  AOI211_X1 U10792 ( .C1(n9658), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n9657), .B(
        n9656), .ZN(n9664) );
  OAI211_X1 U10793 ( .C1(n9662), .C2(n9661), .A(n9660), .B(n9659), .ZN(n9663)
         );
  NAND2_X1 U10794 ( .A1(n9664), .A2(n9663), .ZN(P1_U3242) );
  AND2_X1 U10795 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9666), .ZN(P1_U3292) );
  AND2_X1 U10796 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9666), .ZN(P1_U3293) );
  AND2_X1 U10797 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9666), .ZN(P1_U3294) );
  AND2_X1 U10798 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9666), .ZN(P1_U3295) );
  AND2_X1 U10799 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9666), .ZN(P1_U3296) );
  AND2_X1 U10800 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9666), .ZN(P1_U3297) );
  AND2_X1 U10801 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9666), .ZN(P1_U3298) );
  AND2_X1 U10802 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9666), .ZN(P1_U3299) );
  AND2_X1 U10803 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9666), .ZN(P1_U3300) );
  AND2_X1 U10804 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9666), .ZN(P1_U3301) );
  AND2_X1 U10805 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9666), .ZN(P1_U3302) );
  INV_X1 U10806 ( .A(n9666), .ZN(n9665) );
  INV_X1 U10807 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9975) );
  NOR2_X1 U10808 ( .A1(n9665), .A2(n9975), .ZN(P1_U3303) );
  AND2_X1 U10809 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9666), .ZN(P1_U3304) );
  AND2_X1 U10810 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9666), .ZN(P1_U3305) );
  AND2_X1 U10811 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9666), .ZN(P1_U3306) );
  AND2_X1 U10812 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9666), .ZN(P1_U3307) );
  AND2_X1 U10813 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9666), .ZN(P1_U3308) );
  INV_X1 U10814 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10132) );
  NOR2_X1 U10815 ( .A1(n9665), .A2(n10132), .ZN(P1_U3309) );
  AND2_X1 U10816 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9666), .ZN(P1_U3310) );
  INV_X1 U10817 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10001) );
  NOR2_X1 U10818 ( .A1(n9665), .A2(n10001), .ZN(P1_U3311) );
  AND2_X1 U10819 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9666), .ZN(P1_U3312) );
  AND2_X1 U10820 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9666), .ZN(P1_U3313) );
  AND2_X1 U10821 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9666), .ZN(P1_U3314) );
  AND2_X1 U10822 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9666), .ZN(P1_U3315) );
  AND2_X1 U10823 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9666), .ZN(P1_U3316) );
  INV_X1 U10824 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9974) );
  NOR2_X1 U10825 ( .A1(n9665), .A2(n9974), .ZN(P1_U3317) );
  AND2_X1 U10826 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9666), .ZN(P1_U3318) );
  AND2_X1 U10827 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9666), .ZN(P1_U3319) );
  AND2_X1 U10828 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9666), .ZN(P1_U3320) );
  AND2_X1 U10829 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9666), .ZN(P1_U3321) );
  INV_X1 U10830 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9667) );
  AOI22_X1 U10831 ( .A1(n9724), .A2(n9668), .B1(n9667), .B2(n9722), .ZN(
        P1_U3457) );
  OAI21_X1 U10832 ( .B1(n9670), .B2(n9702), .A(n9669), .ZN(n9672) );
  AOI211_X1 U10833 ( .C1(n9680), .C2(n9673), .A(n9672), .B(n9671), .ZN(n9725)
         );
  INV_X1 U10834 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9674) );
  AOI22_X1 U10835 ( .A1(n9724), .A2(n9725), .B1(n9674), .B2(n9722), .ZN(
        P1_U3460) );
  OAI21_X1 U10836 ( .B1(n9676), .B2(n9704), .A(n9675), .ZN(n9678) );
  AOI211_X1 U10837 ( .C1(n9680), .C2(n9679), .A(n9678), .B(n9677), .ZN(n9726)
         );
  INV_X1 U10838 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9681) );
  AOI22_X1 U10839 ( .A1(n9724), .A2(n9726), .B1(n9681), .B2(n9722), .ZN(
        P1_U3463) );
  AOI22_X1 U10840 ( .A1(n9683), .A2(n9713), .B1(n9712), .B2(n9682), .ZN(n9684)
         );
  OAI211_X1 U10841 ( .C1(n9686), .C2(n9718), .A(n9685), .B(n9684), .ZN(n9687)
         );
  INV_X1 U10842 ( .A(n9687), .ZN(n9727) );
  AOI22_X1 U10843 ( .A1(n9724), .A2(n9727), .B1(n5417), .B2(n9722), .ZN(
        P1_U3466) );
  INV_X1 U10844 ( .A(n9688), .ZN(n9689) );
  OAI21_X1 U10845 ( .B1(n9690), .B2(n9704), .A(n9689), .ZN(n9692) );
  AOI211_X1 U10846 ( .C1(n9708), .C2(n9693), .A(n9692), .B(n9691), .ZN(n9728)
         );
  INV_X1 U10847 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9694) );
  AOI22_X1 U10848 ( .A1(n9724), .A2(n9728), .B1(n9694), .B2(n9722), .ZN(
        P1_U3472) );
  OAI211_X1 U10849 ( .C1(n9697), .C2(n9702), .A(n9696), .B(n9695), .ZN(n9698)
         );
  AOI21_X1 U10850 ( .B1(n9708), .B2(n9699), .A(n9698), .ZN(n9729) );
  INV_X1 U10851 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9700) );
  AOI22_X1 U10852 ( .A1(n9724), .A2(n9729), .B1(n9700), .B2(n9722), .ZN(
        P1_U3475) );
  INV_X1 U10853 ( .A(n9701), .ZN(n9709) );
  OAI22_X1 U10854 ( .A1(n9705), .A2(n9704), .B1(n9703), .B2(n9702), .ZN(n9706)
         );
  AOI211_X1 U10855 ( .C1(n9709), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9730)
         );
  INV_X1 U10856 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9710) );
  AOI22_X1 U10857 ( .A1(n9724), .A2(n9730), .B1(n9710), .B2(n9722), .ZN(
        P1_U3478) );
  INV_X1 U10858 ( .A(n9717), .ZN(n9720) );
  AOI22_X1 U10859 ( .A1(n9714), .A2(n9713), .B1(n9712), .B2(n9711), .ZN(n9715)
         );
  OAI211_X1 U10860 ( .C1(n9718), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9719)
         );
  AOI21_X1 U10861 ( .B1(n9721), .B2(n9720), .A(n9719), .ZN(n9732) );
  INV_X1 U10862 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9723) );
  AOI22_X1 U10863 ( .A1(n9724), .A2(n9732), .B1(n9723), .B2(n9722), .ZN(
        P1_U3481) );
  AOI22_X1 U10864 ( .A1(n9733), .A2(n9725), .B1(n6142), .B2(n9731), .ZN(
        P1_U3525) );
  AOI22_X1 U10865 ( .A1(n9733), .A2(n9726), .B1(n5436), .B2(n9731), .ZN(
        P1_U3526) );
  AOI22_X1 U10866 ( .A1(n9733), .A2(n9727), .B1(n10108), .B2(n9731), .ZN(
        P1_U3527) );
  AOI22_X1 U10867 ( .A1(n9733), .A2(n9728), .B1(n5391), .B2(n9731), .ZN(
        P1_U3529) );
  AOI22_X1 U10868 ( .A1(n9733), .A2(n9729), .B1(n6516), .B2(n9731), .ZN(
        P1_U3530) );
  AOI22_X1 U10869 ( .A1(n9733), .A2(n9730), .B1(n5305), .B2(n9731), .ZN(
        P1_U3531) );
  AOI22_X1 U10870 ( .A1(n9733), .A2(n9732), .B1(n6565), .B2(n9731), .ZN(
        P1_U3532) );
  AOI22_X1 U10871 ( .A1(n9797), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9804), .ZN(n9741) );
  INV_X1 U10872 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9740) );
  INV_X1 U10873 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10103) );
  NAND2_X1 U10874 ( .A1(n9804), .A2(n10103), .ZN(n9735) );
  OAI211_X1 U10875 ( .C1(n9736), .C2(P2_REG2_REG_0__SCAN_IN), .A(n9735), .B(
        n9734), .ZN(n9737) );
  INV_X1 U10876 ( .A(n9737), .ZN(n9739) );
  AOI22_X1 U10877 ( .A1(n9795), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9738) );
  OAI221_X1 U10878 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9741), .C1(n9740), .C2(
        n9739), .A(n9738), .ZN(P2_U3245) );
  AOI22_X1 U10879 ( .A1(n9795), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n9754) );
  NAND2_X1 U10880 ( .A1(n9802), .A2(n9742), .ZN(n9753) );
  NAND2_X1 U10881 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  NAND3_X1 U10882 ( .A1(n9797), .A2(n9746), .A3(n9745), .ZN(n9752) );
  NAND2_X1 U10883 ( .A1(n9748), .A2(n9747), .ZN(n9749) );
  NAND3_X1 U10884 ( .A1(n9804), .A2(n9750), .A3(n9749), .ZN(n9751) );
  NAND4_X1 U10885 ( .A1(n9754), .A2(n9753), .A3(n9752), .A4(n9751), .ZN(
        P2_U3248) );
  INV_X1 U10886 ( .A(n9755), .ZN(n9756) );
  AOI21_X1 U10887 ( .B1(n9795), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n9756), .ZN(
        n9767) );
  NAND2_X1 U10888 ( .A1(n9802), .A2(n9757), .ZN(n9766) );
  OAI211_X1 U10889 ( .C1(n9760), .C2(n9759), .A(n9804), .B(n9758), .ZN(n9765)
         );
  OAI211_X1 U10890 ( .C1(n9763), .C2(n9762), .A(n9797), .B(n9761), .ZN(n9764)
         );
  NAND4_X1 U10891 ( .A1(n9767), .A2(n9766), .A3(n9765), .A4(n9764), .ZN(
        P2_U3249) );
  AOI21_X1 U10892 ( .B1(n9795), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9768), .ZN(
        n9779) );
  NAND2_X1 U10893 ( .A1(n9802), .A2(n9769), .ZN(n9778) );
  OAI211_X1 U10894 ( .C1(n9772), .C2(n9771), .A(n9804), .B(n9770), .ZN(n9777)
         );
  OAI211_X1 U10895 ( .C1(n9775), .C2(n9774), .A(n9797), .B(n9773), .ZN(n9776)
         );
  NAND4_X1 U10896 ( .A1(n9779), .A2(n9778), .A3(n9777), .A4(n9776), .ZN(
        P2_U3251) );
  INV_X1 U10897 ( .A(n9780), .ZN(n9781) );
  AOI21_X1 U10898 ( .B1(n9795), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n9781), .ZN(
        n9792) );
  NAND2_X1 U10899 ( .A1(n9802), .A2(n9782), .ZN(n9791) );
  OAI211_X1 U10900 ( .C1(n9785), .C2(n9784), .A(n9797), .B(n9783), .ZN(n9790)
         );
  OAI211_X1 U10901 ( .C1(n9788), .C2(n9787), .A(n9804), .B(n9786), .ZN(n9789)
         );
  NAND4_X1 U10902 ( .A1(n9792), .A2(n9791), .A3(n9790), .A4(n9789), .ZN(
        P2_U3252) );
  INV_X1 U10903 ( .A(n9793), .ZN(n9794) );
  AOI21_X1 U10904 ( .B1(n9795), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9794), .ZN(
        n9810) );
  OAI211_X1 U10905 ( .C1(n9799), .C2(n9798), .A(n9797), .B(n9796), .ZN(n9809)
         );
  INV_X1 U10906 ( .A(n9800), .ZN(n9801) );
  NAND2_X1 U10907 ( .A1(n9802), .A2(n9801), .ZN(n9808) );
  OAI211_X1 U10908 ( .C1(n9806), .C2(n9805), .A(n9804), .B(n9803), .ZN(n9807)
         );
  NAND4_X1 U10909 ( .A1(n9810), .A2(n9809), .A3(n9808), .A4(n9807), .ZN(
        P2_U3262) );
  NAND2_X1 U10910 ( .A1(n6800), .A2(n9811), .ZN(n9812) );
  XNOR2_X1 U10911 ( .A(n9813), .B(n9812), .ZN(n9888) );
  OAI21_X1 U10912 ( .B1(n4741), .B2(n9815), .A(n9814), .ZN(n9817) );
  NAND2_X1 U10913 ( .A1(n9817), .A2(n9816), .ZN(n9823) );
  AOI22_X1 U10914 ( .A1(n9821), .A2(n9820), .B1(n9819), .B2(n9818), .ZN(n9822)
         );
  NAND2_X1 U10915 ( .A1(n9823), .A2(n9822), .ZN(n9891) );
  AOI21_X1 U10916 ( .B1(n9824), .B2(n9888), .A(n9891), .ZN(n9839) );
  NAND2_X1 U10917 ( .A1(n9826), .A2(n9825), .ZN(n9828) );
  NAND2_X1 U10918 ( .A1(n9828), .A2(n9827), .ZN(n9829) );
  OAI21_X1 U10919 ( .B1(n9830), .B2(n9914), .A(n9829), .ZN(n9832) );
  AND2_X1 U10920 ( .A1(n9832), .A2(n9831), .ZN(n9889) );
  AOI22_X1 U10921 ( .A1(n9835), .A2(n9889), .B1(n9834), .B2(n9833), .ZN(n9836)
         );
  OAI221_X1 U10922 ( .B1(n8713), .B2(n9839), .C1(n9838), .C2(n9837), .A(n9836), 
        .ZN(P2_U3293) );
  INV_X1 U10923 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9842) );
  NOR2_X1 U10924 ( .A1(n9874), .A2(n9842), .ZN(P2_U3297) );
  NOR2_X1 U10925 ( .A1(n9874), .A2(n9843), .ZN(P2_U3298) );
  INV_X1 U10926 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9844) );
  NOR2_X1 U10927 ( .A1(n9874), .A2(n9844), .ZN(P2_U3299) );
  INV_X1 U10928 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9845) );
  NOR2_X1 U10929 ( .A1(n9874), .A2(n9845), .ZN(P2_U3300) );
  INV_X1 U10930 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9846) );
  NOR2_X1 U10931 ( .A1(n9854), .A2(n9846), .ZN(P2_U3301) );
  INV_X1 U10932 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9847) );
  NOR2_X1 U10933 ( .A1(n9854), .A2(n9847), .ZN(P2_U3302) );
  INV_X1 U10934 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9848) );
  NOR2_X1 U10935 ( .A1(n9854), .A2(n9848), .ZN(P2_U3303) );
  INV_X1 U10936 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9849) );
  NOR2_X1 U10937 ( .A1(n9854), .A2(n9849), .ZN(P2_U3304) );
  NOR2_X1 U10938 ( .A1(n9854), .A2(n10089), .ZN(P2_U3305) );
  INV_X1 U10939 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9850) );
  NOR2_X1 U10940 ( .A1(n9854), .A2(n9850), .ZN(P2_U3306) );
  INV_X1 U10941 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9851) );
  NOR2_X1 U10942 ( .A1(n9854), .A2(n9851), .ZN(P2_U3307) );
  INV_X1 U10943 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9852) );
  NOR2_X1 U10944 ( .A1(n9854), .A2(n9852), .ZN(P2_U3308) );
  NOR2_X1 U10945 ( .A1(n9854), .A2(n9991), .ZN(P2_U3309) );
  INV_X1 U10946 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9853) );
  NOR2_X1 U10947 ( .A1(n9854), .A2(n9853), .ZN(P2_U3310) );
  INV_X1 U10948 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9855) );
  NOR2_X1 U10949 ( .A1(n9874), .A2(n9855), .ZN(P2_U3311) );
  INV_X1 U10950 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9856) );
  NOR2_X1 U10951 ( .A1(n9874), .A2(n9856), .ZN(P2_U3312) );
  INV_X1 U10952 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9857) );
  NOR2_X1 U10953 ( .A1(n9874), .A2(n9857), .ZN(P2_U3313) );
  INV_X1 U10954 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9858) );
  NOR2_X1 U10955 ( .A1(n9874), .A2(n9858), .ZN(P2_U3314) );
  INV_X1 U10956 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9859) );
  NOR2_X1 U10957 ( .A1(n9874), .A2(n9859), .ZN(P2_U3315) );
  INV_X1 U10958 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U10959 ( .A1(n9874), .A2(n9860), .ZN(P2_U3316) );
  INV_X1 U10960 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9861) );
  NOR2_X1 U10961 ( .A1(n9874), .A2(n9861), .ZN(P2_U3317) );
  INV_X1 U10962 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9862) );
  NOR2_X1 U10963 ( .A1(n9874), .A2(n9862), .ZN(P2_U3318) );
  INV_X1 U10964 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9863) );
  NOR2_X1 U10965 ( .A1(n9874), .A2(n9863), .ZN(P2_U3319) );
  INV_X1 U10966 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9864) );
  NOR2_X1 U10967 ( .A1(n9874), .A2(n9864), .ZN(P2_U3320) );
  NOR2_X1 U10968 ( .A1(n9874), .A2(n10092), .ZN(P2_U3321) );
  INV_X1 U10969 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9865) );
  NOR2_X1 U10970 ( .A1(n9874), .A2(n9865), .ZN(P2_U3322) );
  INV_X1 U10971 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9866) );
  NOR2_X1 U10972 ( .A1(n9874), .A2(n9866), .ZN(P2_U3323) );
  INV_X1 U10973 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9867) );
  NOR2_X1 U10974 ( .A1(n9874), .A2(n9867), .ZN(P2_U3324) );
  INV_X1 U10975 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9868) );
  NOR2_X1 U10976 ( .A1(n9874), .A2(n9868), .ZN(P2_U3325) );
  INV_X1 U10977 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9869) );
  NOR2_X1 U10978 ( .A1(n9874), .A2(n9869), .ZN(P2_U3326) );
  OAI22_X1 U10979 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9874), .B1(n9873), .B2(
        n9870), .ZN(n9871) );
  INV_X1 U10980 ( .A(n9871), .ZN(P2_U3437) );
  OAI22_X1 U10981 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n9874), .B1(n9873), .B2(
        n9872), .ZN(n9875) );
  INV_X1 U10982 ( .A(n9875), .ZN(P2_U3438) );
  OAI22_X1 U10983 ( .A1(n9878), .A2(n9877), .B1(n6722), .B2(n9876), .ZN(n9880)
         );
  NOR2_X1 U10984 ( .A1(n9880), .A2(n9879), .ZN(n9924) );
  INV_X1 U10985 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9881) );
  AOI22_X1 U10986 ( .A1(n9923), .A2(n9924), .B1(n9881), .B2(n9921), .ZN(
        P2_U3451) );
  OAI21_X1 U10987 ( .B1(n9883), .B2(n9914), .A(n9882), .ZN(n9885) );
  AOI211_X1 U10988 ( .C1(n9919), .C2(n9886), .A(n9885), .B(n9884), .ZN(n9926)
         );
  INV_X1 U10989 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9887) );
  AOI22_X1 U10990 ( .A1(n9923), .A2(n9926), .B1(n9887), .B2(n9921), .ZN(
        P2_U3454) );
  AND2_X1 U10991 ( .A1(n9888), .A2(n9919), .ZN(n9890) );
  NOR3_X1 U10992 ( .A1(n9891), .A2(n9890), .A3(n9889), .ZN(n9927) );
  INV_X1 U10993 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9892) );
  AOI22_X1 U10994 ( .A1(n9923), .A2(n9927), .B1(n9892), .B2(n9921), .ZN(
        P2_U3460) );
  OAI21_X1 U10995 ( .B1(n9894), .B2(n9914), .A(n9893), .ZN(n9896) );
  AOI211_X1 U10996 ( .C1(n9919), .C2(n9897), .A(n9896), .B(n9895), .ZN(n9928)
         );
  INV_X1 U10997 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9898) );
  AOI22_X1 U10998 ( .A1(n9923), .A2(n9928), .B1(n9898), .B2(n9921), .ZN(
        P2_U3466) );
  OAI211_X1 U10999 ( .C1(n9901), .C2(n9914), .A(n9900), .B(n9899), .ZN(n9902)
         );
  AOI21_X1 U11000 ( .B1(n9919), .B2(n9903), .A(n9902), .ZN(n9929) );
  INV_X1 U11001 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9904) );
  AOI22_X1 U11002 ( .A1(n9923), .A2(n9929), .B1(n9904), .B2(n9921), .ZN(
        P2_U3472) );
  INV_X1 U11003 ( .A(n9905), .ZN(n9909) );
  OAI22_X1 U11004 ( .A1(n9907), .A2(n9915), .B1(n9906), .B2(n9914), .ZN(n9908)
         );
  AOI21_X1 U11005 ( .B1(n9910), .B2(n9909), .A(n9908), .ZN(n9911) );
  AND2_X1 U11006 ( .A1(n9912), .A2(n9911), .ZN(n9930) );
  INV_X1 U11007 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9913) );
  AOI22_X1 U11008 ( .A1(n9923), .A2(n9930), .B1(n9913), .B2(n9921), .ZN(
        P2_U3478) );
  OAI22_X1 U11009 ( .A1(n9916), .A2(n9915), .B1(n4590), .B2(n9914), .ZN(n9918)
         );
  AOI211_X1 U11010 ( .C1(n9920), .C2(n9919), .A(n9918), .B(n9917), .ZN(n9933)
         );
  INV_X1 U11011 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9922) );
  AOI22_X1 U11012 ( .A1(n9923), .A2(n9933), .B1(n9922), .B2(n9921), .ZN(
        P2_U3484) );
  AOI22_X1 U11013 ( .A1(n9934), .A2(n9924), .B1(n10103), .B2(n9931), .ZN(
        P2_U3520) );
  AOI22_X1 U11014 ( .A1(n9934), .A2(n9926), .B1(n9925), .B2(n9931), .ZN(
        P2_U3521) );
  AOI22_X1 U11015 ( .A1(n9934), .A2(n9927), .B1(n9990), .B2(n9931), .ZN(
        P2_U3523) );
  AOI22_X1 U11016 ( .A1(n9934), .A2(n9928), .B1(n6387), .B2(n9931), .ZN(
        P2_U3525) );
  AOI22_X1 U11017 ( .A1(n9934), .A2(n9929), .B1(n6385), .B2(n9931), .ZN(
        P2_U3527) );
  AOI22_X1 U11018 ( .A1(n9934), .A2(n9930), .B1(n6383), .B2(n9931), .ZN(
        P2_U3529) );
  AOI22_X1 U11019 ( .A1(n9934), .A2(n9933), .B1(n9932), .B2(n9931), .ZN(
        P2_U3531) );
  INV_X1 U11020 ( .A(n9935), .ZN(n9936) );
  NAND2_X1 U11021 ( .A1(n9937), .A2(n9936), .ZN(n9938) );
  XOR2_X1 U11022 ( .A(n6452), .B(n9938), .Z(ADD_1071_U5) );
  XOR2_X1 U11023 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11024 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(ADD_1071_U56) );
  OAI21_X1 U11025 ( .B1(n9944), .B2(n9943), .A(n9942), .ZN(ADD_1071_U57) );
  OAI21_X1 U11026 ( .B1(n9947), .B2(n9946), .A(n9945), .ZN(ADD_1071_U58) );
  OAI21_X1 U11027 ( .B1(n9950), .B2(n9949), .A(n9948), .ZN(ADD_1071_U59) );
  OAI21_X1 U11028 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(ADD_1071_U60) );
  OAI21_X1 U11029 ( .B1(n9956), .B2(n9955), .A(n9954), .ZN(ADD_1071_U61) );
  AOI21_X1 U11030 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(ADD_1071_U62) );
  AOI21_X1 U11031 ( .B1(n9962), .B2(n9961), .A(n9960), .ZN(ADD_1071_U63) );
  AOI22_X1 U11032 ( .A1(n9965), .A2(keyinput125), .B1(n9964), .B2(keyinput72), 
        .ZN(n9963) );
  OAI221_X1 U11033 ( .B1(n9965), .B2(keyinput125), .C1(n9964), .C2(keyinput72), 
        .A(n9963), .ZN(n9973) );
  AOI22_X1 U11034 ( .A1(n9968), .A2(keyinput97), .B1(n9967), .B2(keyinput115), 
        .ZN(n9966) );
  OAI221_X1 U11035 ( .B1(n9968), .B2(keyinput97), .C1(n9967), .C2(keyinput115), 
        .A(n9966), .ZN(n9972) );
  XOR2_X1 U11036 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput78), .Z(n9971) );
  XNOR2_X1 U11037 ( .A(n9969), .B(keyinput69), .ZN(n9970) );
  OR4_X1 U11038 ( .A1(n9973), .A2(n9972), .A3(n9971), .A4(n9970), .ZN(n9978)
         );
  XNOR2_X1 U11039 ( .A(n9974), .B(keyinput110), .ZN(n9977) );
  XNOR2_X1 U11040 ( .A(n9975), .B(keyinput100), .ZN(n9976) );
  NOR3_X1 U11041 ( .A1(n9978), .A2(n9977), .A3(n9976), .ZN(n10013) );
  INV_X1 U11042 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U11043 ( .A1(n10125), .A2(keyinput118), .B1(n10107), .B2(
        keyinput122), .ZN(n9979) );
  OAI221_X1 U11044 ( .B1(n10125), .B2(keyinput118), .C1(n10107), .C2(
        keyinput122), .A(n9979), .ZN(n9987) );
  AOI22_X1 U11045 ( .A1(n10135), .A2(keyinput93), .B1(n10122), .B2(keyinput94), 
        .ZN(n9980) );
  OAI221_X1 U11046 ( .B1(n10135), .B2(keyinput93), .C1(n10122), .C2(keyinput94), .A(n9980), .ZN(n9986) );
  XNOR2_X1 U11047 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput121), .ZN(n9984)
         );
  XNOR2_X1 U11048 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput103), .ZN(n9983)
         );
  XNOR2_X1 U11049 ( .A(P2_IR_REG_30__SCAN_IN), .B(keyinput106), .ZN(n9982) );
  XNOR2_X1 U11050 ( .A(P1_REG0_REG_28__SCAN_IN), .B(keyinput109), .ZN(n9981)
         );
  NAND4_X1 U11051 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), .ZN(n9985)
         );
  NOR3_X1 U11052 ( .A1(n9987), .A2(n9986), .A3(n9985), .ZN(n10012) );
  AOI22_X1 U11053 ( .A1(n10106), .A2(keyinput90), .B1(keyinput64), .B2(n5169), 
        .ZN(n9988) );
  OAI221_X1 U11054 ( .B1(n10106), .B2(keyinput90), .C1(n5169), .C2(keyinput64), 
        .A(n9988), .ZN(n9998) );
  AOI22_X1 U11055 ( .A1(n9991), .A2(keyinput107), .B1(keyinput91), .B2(n9990), 
        .ZN(n9989) );
  OAI221_X1 U11056 ( .B1(n9991), .B2(keyinput107), .C1(n9990), .C2(keyinput91), 
        .A(n9989), .ZN(n9997) );
  INV_X1 U11057 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U11058 ( .A1(n10094), .A2(keyinput67), .B1(keyinput68), .B2(n9993), 
        .ZN(n9992) );
  OAI221_X1 U11059 ( .B1(n10094), .B2(keyinput67), .C1(n9993), .C2(keyinput68), 
        .A(n9992), .ZN(n9996) );
  AOI22_X1 U11060 ( .A1(n10137), .A2(keyinput79), .B1(n10089), .B2(keyinput66), 
        .ZN(n9994) );
  OAI221_X1 U11061 ( .B1(n10137), .B2(keyinput79), .C1(n10089), .C2(keyinput66), .A(n9994), .ZN(n9995) );
  NOR4_X1 U11062 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n10011)
         );
  AOI22_X1 U11063 ( .A1(n10108), .A2(keyinput116), .B1(keyinput82), .B2(n7911), 
        .ZN(n9999) );
  OAI221_X1 U11064 ( .B1(n10108), .B2(keyinput116), .C1(n7911), .C2(keyinput82), .A(n9999), .ZN(n10009) );
  AOI22_X1 U11065 ( .A1(n10001), .A2(keyinput124), .B1(keyinput96), .B2(n6400), 
        .ZN(n10000) );
  OAI221_X1 U11066 ( .B1(n10001), .B2(keyinput124), .C1(n6400), .C2(keyinput96), .A(n10000), .ZN(n10008) );
  AOI22_X1 U11067 ( .A1(n10132), .A2(keyinput98), .B1(keyinput92), .B2(n10003), 
        .ZN(n10002) );
  OAI221_X1 U11068 ( .B1(n10132), .B2(keyinput98), .C1(n10003), .C2(keyinput92), .A(n10002), .ZN(n10007) );
  XNOR2_X1 U11069 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput85), .ZN(n10005)
         );
  XNOR2_X1 U11070 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput74), .ZN(n10004)
         );
  NAND2_X1 U11071 ( .A1(n10005), .A2(n10004), .ZN(n10006) );
  NOR4_X1 U11072 ( .A1(n10009), .A2(n10008), .A3(n10007), .A4(n10006), .ZN(
        n10010) );
  AND4_X1 U11073 ( .A1(n10013), .A2(n10012), .A3(n10011), .A4(n10010), .ZN(
        n10153) );
  OAI22_X1 U11074 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(keyinput123), .B1(
        keyinput114), .B2(P1_ADDR_REG_0__SCAN_IN), .ZN(n10014) );
  AOI221_X1 U11075 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(keyinput123), .C1(
        P1_ADDR_REG_0__SCAN_IN), .C2(keyinput114), .A(n10014), .ZN(n10021) );
  OAI22_X1 U11076 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput102), .B1(
        P2_REG2_REG_31__SCAN_IN), .B2(keyinput117), .ZN(n10015) );
  AOI221_X1 U11077 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput102), .C1(
        keyinput117), .C2(P2_REG2_REG_31__SCAN_IN), .A(n10015), .ZN(n10020) );
  OAI22_X1 U11078 ( .A1(P2_D_REG_30__SCAN_IN), .A2(keyinput70), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput126), .ZN(n10016) );
  AOI221_X1 U11079 ( .B1(P2_D_REG_30__SCAN_IN), .B2(keyinput70), .C1(
        keyinput126), .C2(P2_REG3_REG_20__SCAN_IN), .A(n10016), .ZN(n10019) );
  OAI22_X1 U11080 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(keyinput84), .B1(
        P2_REG0_REG_2__SCAN_IN), .B2(keyinput75), .ZN(n10017) );
  AOI221_X1 U11081 ( .B1(P1_REG3_REG_19__SCAN_IN), .B2(keyinput84), .C1(
        keyinput75), .C2(P2_REG0_REG_2__SCAN_IN), .A(n10017), .ZN(n10018) );
  NAND4_X1 U11082 ( .A1(n10021), .A2(n10020), .A3(n10019), .A4(n10018), .ZN(
        n10049) );
  OAI22_X1 U11083 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(keyinput86), .B1(
        keyinput65), .B2(P2_REG2_REG_15__SCAN_IN), .ZN(n10022) );
  AOI221_X1 U11084 ( .B1(P1_DATAO_REG_12__SCAN_IN), .B2(keyinput86), .C1(
        P2_REG2_REG_15__SCAN_IN), .C2(keyinput65), .A(n10022), .ZN(n10029) );
  OAI22_X1 U11085 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(keyinput81), .B1(
        keyinput112), .B2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10023) );
  AOI221_X1 U11086 ( .B1(P2_IR_REG_26__SCAN_IN), .B2(keyinput81), .C1(
        P1_ADDR_REG_7__SCAN_IN), .C2(keyinput112), .A(n10023), .ZN(n10028) );
  OAI22_X1 U11087 ( .A1(P2_D_REG_7__SCAN_IN), .A2(keyinput120), .B1(
        keyinput127), .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10024) );
  AOI221_X1 U11088 ( .B1(P2_D_REG_7__SCAN_IN), .B2(keyinput120), .C1(
        P2_REG1_REG_0__SCAN_IN), .C2(keyinput127), .A(n10024), .ZN(n10027) );
  OAI22_X1 U11089 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(keyinput76), .B1(
        keyinput113), .B2(P1_ADDR_REG_12__SCAN_IN), .ZN(n10025) );
  AOI221_X1 U11090 ( .B1(P1_REG3_REG_18__SCAN_IN), .B2(keyinput76), .C1(
        P1_ADDR_REG_12__SCAN_IN), .C2(keyinput113), .A(n10025), .ZN(n10026) );
  NAND4_X1 U11091 ( .A1(n10029), .A2(n10028), .A3(n10027), .A4(n10026), .ZN(
        n10048) );
  OAI22_X1 U11092 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(keyinput77), .B1(
        keyinput105), .B2(P2_REG1_REG_7__SCAN_IN), .ZN(n10030) );
  AOI221_X1 U11093 ( .B1(P2_IR_REG_9__SCAN_IN), .B2(keyinput77), .C1(
        P2_REG1_REG_7__SCAN_IN), .C2(keyinput105), .A(n10030), .ZN(n10037) );
  OAI22_X1 U11094 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(keyinput88), .B1(
        keyinput73), .B2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10031) );
  AOI221_X1 U11095 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(keyinput88), .C1(
        P1_ADDR_REG_2__SCAN_IN), .C2(keyinput73), .A(n10031), .ZN(n10036) );
  OAI22_X1 U11096 ( .A1(n5261), .A2(keyinput89), .B1(n10141), .B2(keyinput119), 
        .ZN(n10032) );
  AOI221_X1 U11097 ( .B1(n5261), .B2(keyinput89), .C1(keyinput119), .C2(n10141), .A(n10032), .ZN(n10035) );
  OAI22_X1 U11098 ( .A1(n10104), .A2(keyinput101), .B1(keyinput111), .B2(
        P1_DATAO_REG_22__SCAN_IN), .ZN(n10033) );
  AOI221_X1 U11099 ( .B1(n10104), .B2(keyinput101), .C1(
        P1_DATAO_REG_22__SCAN_IN), .C2(keyinput111), .A(n10033), .ZN(n10034)
         );
  NAND4_X1 U11100 ( .A1(n10037), .A2(n10036), .A3(n10035), .A4(n10034), .ZN(
        n10047) );
  OAI22_X1 U11101 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(keyinput95), .B1(
        P2_REG0_REG_6__SCAN_IN), .B2(keyinput80), .ZN(n10038) );
  AOI221_X1 U11102 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(keyinput95), .C1(
        keyinput80), .C2(P2_REG0_REG_6__SCAN_IN), .A(n10038), .ZN(n10045) );
  OAI22_X1 U11103 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(keyinput108), .B1(
        P2_REG2_REG_8__SCAN_IN), .B2(keyinput99), .ZN(n10039) );
  AOI221_X1 U11104 ( .B1(P1_REG0_REG_29__SCAN_IN), .B2(keyinput108), .C1(
        keyinput99), .C2(P2_REG2_REG_8__SCAN_IN), .A(n10039), .ZN(n10044) );
  OAI22_X1 U11105 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(keyinput87), .B1(
        keyinput83), .B2(P2_REG1_REG_23__SCAN_IN), .ZN(n10040) );
  AOI221_X1 U11106 ( .B1(P2_IR_REG_11__SCAN_IN), .B2(keyinput87), .C1(
        P2_REG1_REG_23__SCAN_IN), .C2(keyinput83), .A(n10040), .ZN(n10043) );
  OAI22_X1 U11107 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(keyinput104), .B1(
        keyinput71), .B2(P1_REG2_REG_31__SCAN_IN), .ZN(n10041) );
  AOI221_X1 U11108 ( .B1(P2_IR_REG_13__SCAN_IN), .B2(keyinput104), .C1(
        P1_REG2_REG_31__SCAN_IN), .C2(keyinput71), .A(n10041), .ZN(n10042) );
  NAND4_X1 U11109 ( .A1(n10045), .A2(n10044), .A3(n10043), .A4(n10042), .ZN(
        n10046) );
  NOR4_X1 U11110 ( .A1(n10049), .A2(n10048), .A3(n10047), .A4(n10046), .ZN(
        n10152) );
  AOI22_X1 U11111 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(keyinput50), .B1(
        P1_REG3_REG_16__SCAN_IN), .B2(keyinput8), .ZN(n10050) );
  OAI221_X1 U11112 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(keyinput50), .C1(
        P1_REG3_REG_16__SCAN_IN), .C2(keyinput8), .A(n10050), .ZN(n10057) );
  AOI22_X1 U11113 ( .A1(P1_REG2_REG_31__SCAN_IN), .A2(keyinput7), .B1(
        P1_REG3_REG_18__SCAN_IN), .B2(keyinput12), .ZN(n10051) );
  OAI221_X1 U11114 ( .B1(P1_REG2_REG_31__SCAN_IN), .B2(keyinput7), .C1(
        P1_REG3_REG_18__SCAN_IN), .C2(keyinput12), .A(n10051), .ZN(n10056) );
  AOI22_X1 U11115 ( .A1(P1_D_REG_12__SCAN_IN), .A2(keyinput60), .B1(
        P1_D_REG_6__SCAN_IN), .B2(keyinput46), .ZN(n10052) );
  OAI221_X1 U11116 ( .B1(P1_D_REG_12__SCAN_IN), .B2(keyinput60), .C1(
        P1_D_REG_6__SCAN_IN), .C2(keyinput46), .A(n10052), .ZN(n10055) );
  AOI22_X1 U11117 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(keyinput49), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput14), .ZN(n10053) );
  OAI221_X1 U11118 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(keyinput49), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput14), .A(n10053), .ZN(n10054) );
  NOR4_X1 U11119 ( .A1(n10057), .A2(n10056), .A3(n10055), .A4(n10054), .ZN(
        n10087) );
  AOI22_X1 U11120 ( .A1(P2_REG1_REG_23__SCAN_IN), .A2(keyinput19), .B1(
        P2_REG2_REG_12__SCAN_IN), .B2(keyinput32), .ZN(n10058) );
  OAI221_X1 U11121 ( .B1(P2_REG1_REG_23__SCAN_IN), .B2(keyinput19), .C1(
        P2_REG2_REG_12__SCAN_IN), .C2(keyinput32), .A(n10058), .ZN(n10065) );
  AOI22_X1 U11122 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput57), .B1(
        P2_D_REG_19__SCAN_IN), .B2(keyinput43), .ZN(n10059) );
  OAI221_X1 U11123 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput57), .C1(
        P2_D_REG_19__SCAN_IN), .C2(keyinput43), .A(n10059), .ZN(n10064) );
  AOI22_X1 U11124 ( .A1(P2_D_REG_30__SCAN_IN), .A2(keyinput6), .B1(
        P2_IR_REG_26__SCAN_IN), .B2(keyinput17), .ZN(n10060) );
  OAI221_X1 U11125 ( .B1(P2_D_REG_30__SCAN_IN), .B2(keyinput6), .C1(
        P2_IR_REG_26__SCAN_IN), .C2(keyinput17), .A(n10060), .ZN(n10063) );
  AOI22_X1 U11126 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(keyinput1), .B1(
        P2_REG1_REG_3__SCAN_IN), .B2(keyinput27), .ZN(n10061) );
  OAI221_X1 U11127 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(keyinput1), .C1(
        P2_REG1_REG_3__SCAN_IN), .C2(keyinput27), .A(n10061), .ZN(n10062) );
  NOR4_X1 U11128 ( .A1(n10065), .A2(n10064), .A3(n10063), .A4(n10062), .ZN(
        n10086) );
  AOI22_X1 U11129 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput38), .B1(SI_25_), 
        .B2(keyinput28), .ZN(n10066) );
  OAI221_X1 U11130 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput38), .C1(SI_25_), .C2(keyinput28), .A(n10066), .ZN(n10073) );
  AOI22_X1 U11131 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(keyinput61), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(keyinput47), .ZN(n10067) );
  OAI221_X1 U11132 ( .B1(P2_REG2_REG_19__SCAN_IN), .B2(keyinput61), .C1(
        P1_DATAO_REG_22__SCAN_IN), .C2(keyinput47), .A(n10067), .ZN(n10072) );
  AOI22_X1 U11133 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput33), .B1(
        P2_IR_REG_11__SCAN_IN), .B2(keyinput23), .ZN(n10068) );
  OAI221_X1 U11134 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput33), .C1(
        P2_IR_REG_11__SCAN_IN), .C2(keyinput23), .A(n10068), .ZN(n10071) );
  AOI22_X1 U11135 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(keyinput51), .B1(
        P1_IR_REG_28__SCAN_IN), .B2(keyinput5), .ZN(n10069) );
  OAI221_X1 U11136 ( .B1(P1_DATAO_REG_13__SCAN_IN), .B2(keyinput51), .C1(
        P1_IR_REG_28__SCAN_IN), .C2(keyinput5), .A(n10069), .ZN(n10070) );
  NOR4_X1 U11137 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10085) );
  AOI22_X1 U11138 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(keyinput9), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(keyinput42), .ZN(n10074) );
  OAI221_X1 U11139 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(keyinput9), .C1(
        P2_IR_REG_30__SCAN_IN), .C2(keyinput42), .A(n10074), .ZN(n10083) );
  AOI22_X1 U11140 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(keyinput35), .B1(
        P1_D_REG_20__SCAN_IN), .B2(keyinput36), .ZN(n10075) );
  OAI221_X1 U11141 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(keyinput35), .C1(
        P1_D_REG_20__SCAN_IN), .C2(keyinput36), .A(n10075), .ZN(n10082) );
  AOI22_X1 U11142 ( .A1(n5169), .A2(keyinput0), .B1(keyinput48), .B2(n10077), 
        .ZN(n10076) );
  OAI221_X1 U11143 ( .B1(n5169), .B2(keyinput0), .C1(n10077), .C2(keyinput48), 
        .A(n10076), .ZN(n10081) );
  INV_X1 U11144 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10079) );
  AOI22_X1 U11145 ( .A1(n10079), .A2(keyinput11), .B1(n5305), .B2(keyinput59), 
        .ZN(n10078) );
  OAI221_X1 U11146 ( .B1(n10079), .B2(keyinput11), .C1(n5305), .C2(keyinput59), 
        .A(n10078), .ZN(n10080) );
  NOR4_X1 U11147 ( .A1(n10083), .A2(n10082), .A3(n10081), .A4(n10080), .ZN(
        n10084) );
  NAND4_X1 U11148 ( .A1(n10087), .A2(n10086), .A3(n10085), .A4(n10084), .ZN(
        n10151) );
  AOI22_X1 U11149 ( .A1(n5261), .A2(keyinput25), .B1(keyinput2), .B2(n10089), 
        .ZN(n10088) );
  OAI221_X1 U11150 ( .B1(n5261), .B2(keyinput25), .C1(n10089), .C2(keyinput2), 
        .A(n10088), .ZN(n10101) );
  AOI22_X1 U11151 ( .A1(n10092), .A2(keyinput56), .B1(keyinput16), .B2(n10091), 
        .ZN(n10090) );
  OAI221_X1 U11152 ( .B1(n10092), .B2(keyinput56), .C1(n10091), .C2(keyinput16), .A(n10090), .ZN(n10100) );
  AOI22_X1 U11153 ( .A1(n10095), .A2(keyinput62), .B1(n10094), .B2(keyinput3), 
        .ZN(n10093) );
  OAI221_X1 U11154 ( .B1(n10095), .B2(keyinput62), .C1(n10094), .C2(keyinput3), 
        .A(n10093), .ZN(n10099) );
  XNOR2_X1 U11155 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput13), .ZN(n10097) );
  XNOR2_X1 U11156 ( .A(keyinput4), .B(P1_REG0_REG_11__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U11157 ( .A1(n10097), .A2(n10096), .ZN(n10098) );
  NOR4_X1 U11158 ( .A1(n10101), .A2(n10100), .A3(n10099), .A4(n10098), .ZN(
        n10149) );
  AOI22_X1 U11159 ( .A1(n10104), .A2(keyinput37), .B1(keyinput63), .B2(n10103), 
        .ZN(n10102) );
  OAI221_X1 U11160 ( .B1(n10104), .B2(keyinput37), .C1(n10103), .C2(keyinput63), .A(n10102), .ZN(n10115) );
  AOI22_X1 U11161 ( .A1(n10107), .A2(keyinput58), .B1(n10106), .B2(keyinput26), 
        .ZN(n10105) );
  OAI221_X1 U11162 ( .B1(n10107), .B2(keyinput58), .C1(n10106), .C2(keyinput26), .A(n10105), .ZN(n10114) );
  XOR2_X1 U11163 ( .A(n10108), .B(keyinput52), .Z(n10112) );
  XNOR2_X1 U11164 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput10), .ZN(n10111)
         );
  XNOR2_X1 U11165 ( .A(P1_REG0_REG_29__SCAN_IN), .B(keyinput44), .ZN(n10110)
         );
  XNOR2_X1 U11166 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput39), .ZN(n10109)
         );
  NAND4_X1 U11167 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .ZN(
        n10113) );
  NOR3_X1 U11168 ( .A1(n10115), .A2(n10114), .A3(n10113), .ZN(n10148) );
  AOI22_X1 U11169 ( .A1(n7911), .A2(keyinput18), .B1(n10117), .B2(keyinput22), 
        .ZN(n10116) );
  OAI221_X1 U11170 ( .B1(n7911), .B2(keyinput18), .C1(n10117), .C2(keyinput22), 
        .A(n10116), .ZN(n10130) );
  AOI22_X1 U11171 ( .A1(n10120), .A2(keyinput20), .B1(keyinput24), .B2(n10119), 
        .ZN(n10118) );
  OAI221_X1 U11172 ( .B1(n10120), .B2(keyinput20), .C1(n10119), .C2(keyinput24), .A(n10118), .ZN(n10129) );
  INV_X1 U11173 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n10123) );
  AOI22_X1 U11174 ( .A1(n10123), .A2(keyinput53), .B1(n10122), .B2(keyinput30), 
        .ZN(n10121) );
  OAI221_X1 U11175 ( .B1(n10123), .B2(keyinput53), .C1(n10122), .C2(keyinput30), .A(n10121), .ZN(n10128) );
  AOI22_X1 U11176 ( .A1(n10126), .A2(keyinput45), .B1(keyinput54), .B2(n10125), 
        .ZN(n10124) );
  OAI221_X1 U11177 ( .B1(n10126), .B2(keyinput45), .C1(n10125), .C2(keyinput54), .A(n10124), .ZN(n10127) );
  NOR4_X1 U11178 ( .A1(n10130), .A2(n10129), .A3(n10128), .A4(n10127), .ZN(
        n10147) );
  AOI22_X1 U11179 ( .A1(n10133), .A2(keyinput40), .B1(n10132), .B2(keyinput34), 
        .ZN(n10131) );
  OAI221_X1 U11180 ( .B1(n10133), .B2(keyinput40), .C1(n10132), .C2(keyinput34), .A(n10131), .ZN(n10145) );
  AOI22_X1 U11181 ( .A1(n10135), .A2(keyinput29), .B1(keyinput41), .B2(n6385), 
        .ZN(n10134) );
  OAI221_X1 U11182 ( .B1(n10135), .B2(keyinput29), .C1(n6385), .C2(keyinput41), 
        .A(n10134), .ZN(n10144) );
  AOI22_X1 U11183 ( .A1(n10138), .A2(keyinput31), .B1(keyinput15), .B2(n10137), 
        .ZN(n10136) );
  OAI221_X1 U11184 ( .B1(n10138), .B2(keyinput31), .C1(n10137), .C2(keyinput15), .A(n10136), .ZN(n10143) );
  AOI22_X1 U11185 ( .A1(n10141), .A2(keyinput55), .B1(n10140), .B2(keyinput21), 
        .ZN(n10139) );
  OAI221_X1 U11186 ( .B1(n10141), .B2(keyinput55), .C1(n10140), .C2(keyinput21), .A(n10139), .ZN(n10142) );
  NOR4_X1 U11187 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        n10146) );
  NAND4_X1 U11188 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10150) );
  AOI211_X1 U11189 ( .C1(n10153), .C2(n10152), .A(n10151), .B(n10150), .ZN(
        n10172) );
  AOI211_X1 U11190 ( .C1(n10157), .C2(n10156), .A(n10155), .B(n10154), .ZN(
        n10170) );
  AOI21_X1 U11191 ( .B1(n10160), .B2(n10159), .A(n10158), .ZN(n10161) );
  OAI22_X1 U11192 ( .A1(n10164), .A2(n10163), .B1(n10162), .B2(n10161), .ZN(
        n10169) );
  INV_X1 U11193 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10166) );
  OAI21_X1 U11194 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(n10168) );
  OR3_X1 U11195 ( .A1(n10170), .A2(n10169), .A3(n10168), .ZN(n10171) );
  XOR2_X1 U11196 ( .A(n10172), .B(n10171), .Z(P1_U3251) );
  XOR2_X1 U11197 ( .A(n10173), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11198 ( .A1(n10175), .A2(n10174), .ZN(n10176) );
  XOR2_X1 U11199 ( .A(n10176), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  OAI21_X1 U11200 ( .B1(n10179), .B2(n10178), .A(n10177), .ZN(n10181) );
  XOR2_X1 U11201 ( .A(n10181), .B(n10180), .Z(ADD_1071_U55) );
  AOI21_X1 U11202 ( .B1(n10184), .B2(n10183), .A(n10182), .ZN(ADD_1071_U47) );
  XOR2_X1 U11203 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10185), .Z(ADD_1071_U48) );
  XOR2_X1 U11204 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10186), .Z(ADD_1071_U49) );
  XOR2_X1 U11205 ( .A(n10188), .B(n10187), .Z(ADD_1071_U54) );
  XOR2_X1 U11206 ( .A(n10190), .B(n10189), .Z(ADD_1071_U53) );
  XNOR2_X1 U11207 ( .A(n10192), .B(n10191), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4844 ( .A(n5366), .Z(n5548) );
endmodule

