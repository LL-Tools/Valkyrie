

module b14_C_AntiSAT_k_128_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2053, n2054, n2055, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726;

  INV_X1 U2296 ( .A(n3394), .ZN(n3407) );
  CLKBUF_X3 U2298 ( .A(n2067), .Z(n2452) );
  AND2_X1 U2299 ( .A1(n3857), .A2(n3856), .ZN(n3859) );
  CLKBUF_X3 U2300 ( .A(n3591), .Z(n2053) );
  BUF_X1 U2301 ( .A(n2818), .Z(n2916) );
  XNOR2_X1 U2302 ( .A(n3859), .B(n3858), .ZN(n4171) );
  AND4_X1 U2303 ( .A1(n2303), .A2(n2302), .A3(n2301), .A4(n2300), .ZN(n2939)
         );
  NAND2_X1 U2304 ( .A1(n3476), .A2(n2216), .ZN(n2215) );
  INV_X1 U2305 ( .A(n3065), .ZN(n3754) );
  XNOR2_X1 U2306 ( .A(n2278), .B(IR_REG_30__SCAN_IN), .ZN(n4350) );
  BUF_X1 U2308 ( .A(n2410), .Z(n3591) );
  NOR2_X2 U2309 ( .A1(n4121), .A2(n4235), .ZN(n4090) );
  OAI21_X2 U2310 ( .B1(n3170), .B2(n3169), .A(n3168), .ZN(n3221) );
  NOR2_X1 U2312 ( .A1(n4350), .A2(n2282), .ZN(n2307) );
  NAND2_X1 U2313 ( .A1(n2177), .A2(n2182), .ZN(n3894) );
  NAND2_X1 U2314 ( .A1(n4530), .A2(n4021), .ZN(n4348) );
  INV_X2 U2315 ( .A(n2057), .ZN(n2932) );
  AND4_X2 U2317 ( .A1(n2287), .A2(n2286), .A3(n2285), .A4(n2284), .ZN(n2298)
         );
  AND2_X1 U2318 ( .A1(n4350), .A2(n2282), .ZN(n2306) );
  XNOR2_X1 U2319 ( .A(n2206), .B(n2205), .ZN(n4361) );
  OAI21_X1 U2320 ( .B1(n2687), .B2(n2135), .A(n2133), .ZN(n2691) );
  NOR2_X1 U2321 ( .A1(n2069), .A2(n2686), .ZN(n2137) );
  NAND2_X1 U2322 ( .A1(n2223), .A2(n2227), .ZN(n3441) );
  AND2_X1 U2323 ( .A1(n4045), .A2(n4053), .ZN(n4047) );
  NOR2_X1 U2324 ( .A1(n3884), .A2(n3383), .ZN(n3868) );
  AOI21_X1 U2325 ( .B1(n2227), .B2(n2226), .A(n2225), .ZN(n2224) );
  AOI21_X1 U2326 ( .B1(n3004), .B2(n3692), .A(n3003), .ZN(n3050) );
  NAND2_X2 U2327 ( .A1(n4536), .A2(n4021), .ZN(n4272) );
  OR2_X1 U2328 ( .A1(n3640), .A2(n3664), .ZN(n2697) );
  AND2_X1 U2329 ( .A1(n2153), .A2(n2152), .ZN(n2807) );
  AND2_X1 U2330 ( .A1(n3674), .A2(n3678), .ZN(n3651) );
  NAND2_X1 U2331 ( .A1(n2107), .A2(n2106), .ZN(n3549) );
  AND4_X1 U2332 ( .A1(n2333), .A2(n2332), .A3(n2331), .A4(n2330), .ZN(n3093)
         );
  AND4_X1 U2333 ( .A1(n2322), .A2(n2321), .A3(n2320), .A4(n2319), .ZN(n3065)
         );
  INV_X1 U2334 ( .A(n2939), .ZN(n3036) );
  NAND3_X1 U2335 ( .A1(n2297), .A2(n2296), .A3(n2295), .ZN(n3756) );
  BUF_X2 U2336 ( .A(n2307), .Z(n2534) );
  NAND2_X2 U2337 ( .A1(n2847), .A2(n2846), .ZN(n3394) );
  NAND2_X1 U2338 ( .A1(n4354), .A2(n3731), .ZN(n2846) );
  INV_X1 U2339 ( .A(n2641), .ZN(n4351) );
  XNOR2_X1 U2340 ( .A(n2638), .B(IR_REG_26__SCAN_IN), .ZN(n2642) );
  XNOR2_X1 U2341 ( .A(n2635), .B(n2634), .ZN(n2641) );
  NAND2_X1 U2342 ( .A1(n2629), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  XNOR2_X1 U2343 ( .A(n2579), .B(n2578), .ZN(n3731) );
  AND2_X4 U2344 ( .A1(n4350), .A2(n2283), .ZN(n2308) );
  NAND2_X1 U2345 ( .A1(n2577), .A2(IR_REG_31__SCAN_IN), .ZN(n2579) );
  INV_X1 U2346 ( .A(n2645), .ZN(n4354) );
  AND2_X1 U2347 ( .A1(n2160), .A2(n2085), .ZN(n2105) );
  OR2_X1 U2348 ( .A1(n2281), .A2(n2242), .ZN(n2160) );
  OR2_X1 U2349 ( .A1(n2279), .A2(n2725), .ZN(n2278) );
  AND2_X1 U2350 ( .A1(n2184), .A2(n2077), .ZN(n2279) );
  NOR2_X1 U2351 ( .A1(n2188), .A2(n2185), .ZN(n2184) );
  NAND2_X1 U2352 ( .A1(n2277), .A2(n2189), .ZN(n2188) );
  AND2_X1 U2353 ( .A1(n2272), .A2(n2245), .ZN(n2244) );
  AND2_X1 U2354 ( .A1(n2122), .A2(n2274), .ZN(n2121) );
  AND4_X1 U2355 ( .A1(n2384), .A2(n2271), .A3(n2270), .A4(n2269), .ZN(n2272)
         );
  AND2_X1 U2356 ( .A1(n2273), .A2(n2247), .ZN(n2245) );
  NOR2_X1 U2357 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2632)
         );
  NOR2_X1 U2358 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2262)
         );
  NOR3_X1 U2359 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .A3(
        IR_REG_15__SCAN_IN), .ZN(n2273) );
  BUF_X4 U2361 ( .A(n3369), .Z(n2057) );
  NAND2_X2 U2362 ( .A1(n2818), .A2(n2846), .ZN(n3369) );
  OAI21_X2 U2363 ( .B1(n3115), .B2(n3114), .A(n3113), .ZN(n3116) );
  OR2_X2 U2364 ( .A1(n3944), .A2(n3943), .ZN(n3942) );
  OAI21_X2 U2365 ( .B1(n3284), .B2(n2254), .A(n2251), .ZN(n3523) );
  AOI21_X2 U2366 ( .B1(n3968), .B2(n3634), .A(n3635), .ZN(n3950) );
  XNOR2_X2 U2367 ( .A(n2631), .B(n2630), .ZN(n2640) );
  NAND2_X4 U2368 ( .A1(n2818), .A2(n2817), .ZN(n2931) );
  INV_X2 U2369 ( .A(n2306), .ZN(n2059) );
  NOR2_X1 U2370 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2275)
         );
  NOR2_X1 U2371 ( .A1(n2068), .A2(n2182), .ZN(n2179) );
  INV_X1 U2372 ( .A(n2173), .ZN(n2169) );
  INV_X1 U2373 ( .A(n3201), .ZN(n3205) );
  OR2_X1 U2374 ( .A1(n3877), .A2(n2621), .ZN(n3861) );
  INV_X1 U2375 ( .A(IR_REG_23__SCAN_IN), .ZN(n2644) );
  INV_X1 U2376 ( .A(n2312), .ZN(n2268) );
  INV_X1 U2377 ( .A(n3525), .ZN(n3296) );
  OAI22_X1 U2378 ( .A1(n2298), .A2(n2931), .B1(n2058), .B2(n2904), .ZN(n2848)
         );
  NAND2_X1 U2379 ( .A1(n2158), .A2(n2157), .ZN(n2156) );
  INV_X1 U2380 ( .A(n2796), .ZN(n2157) );
  OR2_X1 U2381 ( .A1(n2788), .A2(n3106), .ZN(n2153) );
  NAND2_X1 U2382 ( .A1(n4372), .A2(n4371), .ZN(n4370) );
  NAND2_X1 U2383 ( .A1(n2093), .A2(n2092), .ZN(n2091) );
  INV_X1 U2384 ( .A(n4433), .ZN(n2092) );
  XNOR2_X1 U2385 ( .A(n3782), .B(n4502), .ZN(n4445) );
  NAND2_X1 U2386 ( .A1(n4454), .A2(n2203), .ZN(n2202) );
  NAND2_X1 U2387 ( .A1(n4501), .A2(n2204), .ZN(n2203) );
  INV_X1 U2388 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2204) );
  INV_X1 U2389 ( .A(n3629), .ZN(n3839) );
  NAND2_X1 U2390 ( .A1(n2624), .A2(n2132), .ZN(n3842) );
  OR2_X1 U2391 ( .A1(n4216), .A2(n4014), .ZN(n2488) );
  AOI21_X1 U2392 ( .B1(n2264), .B2(n2064), .A(n2082), .ZN(n2167) );
  NAND2_X1 U2393 ( .A1(n4047), .A2(n2064), .ZN(n2166) );
  NOR2_X1 U2394 ( .A1(n3839), .A2(n3614), .ZN(n2132) );
  NAND2_X1 U2395 ( .A1(n2687), .A2(n4145), .ZN(n2138) );
  NAND2_X1 U2396 ( .A1(n2497), .A2(IR_REG_31__SCAN_IN), .ZN(n2576) );
  NOR2_X1 U2397 ( .A1(n2202), .A2(n4465), .ZN(n4464) );
  NOR2_X1 U2398 ( .A1(n4460), .A2(n3813), .ZN(n4470) );
  NAND2_X1 U2399 ( .A1(n4470), .A2(n4471), .ZN(n4468) );
  INV_X1 U2400 ( .A(n3558), .ZN(n2240) );
  INV_X1 U2401 ( .A(n3559), .ZN(n2239) );
  INV_X1 U2402 ( .A(n2125), .ZN(n2124) );
  NOR2_X1 U2403 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2190)
         );
  INV_X1 U2404 ( .A(IR_REG_18__SCAN_IN), .ZN(n2122) );
  NAND2_X1 U2405 ( .A1(n2240), .A2(n2239), .ZN(n2238) );
  NOR2_X1 U2406 ( .A1(n3331), .A2(n2232), .ZN(n2231) );
  INV_X1 U2407 ( .A(n2238), .ZN(n2232) );
  AOI21_X1 U2408 ( .B1(n2258), .B2(n2257), .A(n2256), .ZN(n2255) );
  INV_X1 U2409 ( .A(n3464), .ZN(n2256) );
  INV_X1 U2410 ( .A(n2257), .ZN(n2253) );
  OR2_X1 U2411 ( .A1(n2837), .A2(n4356), .ZN(n2847) );
  AND3_X1 U2412 ( .A1(n2191), .A2(n2086), .A3(n2193), .ZN(n3771) );
  OAI21_X1 U2413 ( .B1(n4413), .B2(n4409), .A(n2197), .ZN(n3779) );
  OR2_X1 U2414 ( .A1(n3788), .A2(REG2_REG_13__SCAN_IN), .ZN(n2197) );
  NOR2_X1 U2415 ( .A1(n2068), .A2(n2181), .ZN(n2180) );
  INV_X1 U2416 ( .A(n2183), .ZN(n2181) );
  AND2_X1 U2417 ( .A1(n2063), .A2(n2520), .ZN(n2183) );
  NAND2_X1 U2418 ( .A1(n2063), .A2(n2080), .ZN(n2182) );
  INV_X1 U2419 ( .A(n3701), .ZN(n2115) );
  INV_X1 U2420 ( .A(n2117), .ZN(n2116) );
  OAI21_X1 U2421 ( .B1(n3684), .B2(n2118), .A(n3699), .ZN(n2117) );
  INV_X1 U2422 ( .A(n3700), .ZN(n2118) );
  OR2_X1 U2423 ( .A1(n3183), .A2(n3690), .ZN(n2597) );
  INV_X1 U2424 ( .A(n3045), .ZN(n2936) );
  NOR2_X1 U2425 ( .A1(n3126), .A2(n3205), .ZN(n2142) );
  OR2_X1 U2426 ( .A1(n2829), .A2(n2646), .ZN(n2704) );
  INV_X1 U2427 ( .A(n2121), .ZN(n2120) );
  INV_X1 U2428 ( .A(n2275), .ZN(n2185) );
  NAND2_X1 U2429 ( .A1(n2496), .A2(n2184), .ZN(n2289) );
  AND2_X1 U2430 ( .A1(n2569), .A2(n2571), .ZN(n2633) );
  INV_X1 U2431 ( .A(IR_REG_19__SCAN_IN), .ZN(n2575) );
  INV_X1 U2432 ( .A(IR_REG_15__SCAN_IN), .ZN(n2459) );
  INV_X1 U2433 ( .A(IR_REG_1__SCAN_IN), .ZN(n2139) );
  AND2_X1 U2434 ( .A1(n3282), .A2(n3283), .ZN(n2258) );
  OR2_X1 U2435 ( .A1(n3282), .A2(n3283), .ZN(n2257) );
  NAND2_X1 U2436 ( .A1(n3482), .A2(n3310), .ZN(n2250) );
  NAND2_X1 U2437 ( .A1(n3441), .A2(n3368), .ZN(n3503) );
  AND2_X1 U2438 ( .A1(n3371), .A2(n3372), .ZN(n3368) );
  INV_X1 U2439 ( .A(n3549), .ZN(n2974) );
  AOI21_X1 U2440 ( .B1(n2836), .B2(n2822), .A(n2819), .ZN(n2820) );
  NOR2_X1 U2441 ( .A1(n2916), .A2(n2140), .ZN(n2819) );
  NAND2_X1 U2442 ( .A1(n2825), .A2(n2824), .ZN(n2851) );
  OAI22_X1 U2443 ( .A1(n4253), .A2(n3358), .B1(n2931), .B2(n3267), .ZN(n3283)
         );
  INV_X1 U2444 ( .A(n2922), .ZN(n2220) );
  OR2_X1 U2445 ( .A1(n2441), .A2(n2440), .ZN(n2450) );
  NAND2_X1 U2446 ( .A1(n2310), .A2(n2111), .ZN(n2110) );
  NAND2_X1 U2447 ( .A1(n2534), .A2(REG0_REG_3__SCAN_IN), .ZN(n2111) );
  NOR2_X1 U2448 ( .A1(n2802), .A2(n3012), .ZN(n2103) );
  NAND2_X1 U2449 ( .A1(n4359), .A2(REG1_REG_5__SCAN_IN), .ZN(n2155) );
  NAND2_X1 U2450 ( .A1(n2783), .A2(n2194), .ZN(n2191) );
  NOR2_X1 U2451 ( .A1(n2811), .A2(n2195), .ZN(n2194) );
  INV_X1 U2452 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2195) );
  OR2_X1 U2453 ( .A1(n2196), .A2(n2811), .ZN(n2193) );
  OAI22_X1 U2454 ( .A1(n2807), .A2(n2753), .B1(n4534), .B2(n2809), .ZN(n3792)
         );
  NAND2_X1 U2455 ( .A1(n4370), .A2(n3773), .ZN(n3774) );
  NAND2_X1 U2456 ( .A1(n4380), .A2(REG2_REG_10__SCAN_IN), .ZN(n4379) );
  NAND2_X1 U2457 ( .A1(n4391), .A2(n3776), .ZN(n3777) );
  NAND2_X1 U2458 ( .A1(n4401), .A2(REG2_REG_12__SCAN_IN), .ZN(n4400) );
  XNOR2_X1 U2459 ( .A(n3779), .B(n4507), .ZN(n4424) );
  NAND2_X1 U2460 ( .A1(n4437), .A2(n3808), .ZN(n3809) );
  AND2_X1 U2461 ( .A1(n2091), .A2(n2088), .ZN(n3782) );
  NAND2_X1 U2462 ( .A1(n4445), .A2(n4443), .ZN(n4444) );
  OR2_X1 U2463 ( .A1(n2554), .A2(n2553), .ZN(n3856) );
  OR2_X1 U2464 ( .A1(n2527), .A2(n4551), .ZN(n2542) );
  NAND2_X1 U2465 ( .A1(n4196), .A2(n2519), .ZN(n2520) );
  AND2_X1 U2466 ( .A1(n3916), .A2(n2615), .ZN(n3943) );
  INV_X1 U2467 ( .A(n4356), .ZN(n3818) );
  INV_X1 U2468 ( .A(n4012), .ZN(n2487) );
  AND2_X1 U2469 ( .A1(n3992), .A2(n3993), .ZN(n4012) );
  NOR2_X1 U2470 ( .A1(n2174), .A2(n2389), .ZN(n2173) );
  INV_X1 U2471 ( .A(n3750), .ZN(n3246) );
  AND2_X1 U2472 ( .A1(n2837), .A2(n2645), .ZN(n2889) );
  AND2_X1 U2473 ( .A1(n3850), .A2(n3419), .ZN(n2690) );
  NAND2_X1 U2474 ( .A1(n2690), .A2(n2689), .ZN(n4154) );
  NAND2_X1 U2475 ( .A1(n3842), .A2(n2625), .ZN(n2678) );
  INV_X1 U2476 ( .A(n4160), .ZN(n3848) );
  AND2_X1 U2477 ( .A1(n3868), .A2(n3848), .ZN(n3850) );
  NAND2_X1 U2478 ( .A1(n3937), .A2(n2066), .ZN(n3884) );
  AND2_X1 U2479 ( .A1(n3252), .A2(n3251), .ZN(n3268) );
  NAND2_X1 U2480 ( .A1(n2843), .A2(n2738), .ZN(n4163) );
  AND2_X1 U2481 ( .A1(n2889), .A2(n3731), .ZN(n4021) );
  AND2_X1 U2482 ( .A1(n2639), .A2(n2642), .ZN(n2729) );
  OR2_X1 U2483 ( .A1(n2436), .A2(IR_REG_10__SCAN_IN), .ZN(n2406) );
  INV_X1 U2484 ( .A(IR_REG_7__SCAN_IN), .ZN(n2360) );
  INV_X1 U2485 ( .A(IR_REG_3__SCAN_IN), .ZN(n2313) );
  NOR2_X1 U2486 ( .A1(n2065), .A2(n2211), .ZN(n2208) );
  INV_X1 U2487 ( .A(n3402), .ZN(n2219) );
  NOR2_X1 U2488 ( .A1(n2218), .A2(n2217), .ZN(n2216) );
  INV_X1 U2489 ( .A(n2081), .ZN(n2218) );
  INV_X1 U2490 ( .A(n2221), .ZN(n2923) );
  OR2_X1 U2491 ( .A1(n2059), .A2(n2990), .ZN(n2319) );
  OAI21_X2 U2492 ( .B1(n2919), .B2(U3149), .A(n2918), .ZN(n3574) );
  INV_X1 U2493 ( .A(n4219), .ZN(n4228) );
  XNOR2_X1 U2494 ( .A(n2102), .B(n2101), .ZN(n2783) );
  INV_X1 U2495 ( .A(n4358), .ZN(n2101) );
  NAND2_X1 U2496 ( .A1(n4392), .A2(n4393), .ZN(n4391) );
  XNOR2_X1 U2497 ( .A(n3809), .B(n4502), .ZN(n4448) );
  NOR2_X1 U2498 ( .A1(n4448), .A2(REG1_REG_16__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U2499 ( .A1(n2201), .A2(n4411), .ZN(n2200) );
  NAND2_X1 U2500 ( .A1(n2202), .A2(n4465), .ZN(n2201) );
  AOI21_X1 U2501 ( .B1(n4467), .B2(ADDR_REG_18__SCAN_IN), .A(n4466), .ZN(n2199) );
  XNOR2_X1 U2502 ( .A(n2147), .B(n3815), .ZN(n3820) );
  NAND2_X1 U2503 ( .A1(n4468), .A2(n2090), .ZN(n2147) );
  AND2_X1 U2504 ( .A1(n2768), .A2(n2860), .ZN(n4469) );
  OR2_X1 U2505 ( .A1(n4464), .A2(n2089), .ZN(n2104) );
  AOI21_X1 U2506 ( .B1(n2624), .B2(n2131), .A(n2128), .ZN(n2679) );
  NAND2_X1 U2507 ( .A1(n2130), .A2(n2129), .ZN(n2128) );
  AND2_X1 U2508 ( .A1(n2132), .A2(n3612), .ZN(n2131) );
  NOR2_X1 U2509 ( .A1(n4533), .A2(n4145), .ZN(n2134) );
  NAND2_X1 U2510 ( .A1(n2137), .A2(n4536), .ZN(n2135) );
  OR2_X1 U2511 ( .A1(n3273), .A2(n4272), .ZN(n2670) );
  OAI21_X1 U2512 ( .B1(n2690), .B2(n2689), .A(n4154), .ZN(n3830) );
  XNOR2_X1 U2513 ( .A(n2576), .B(IR_REG_19__SCAN_IN), .ZN(n4356) );
  AND2_X1 U2514 ( .A1(n3442), .A2(n3443), .ZN(n3363) );
  NAND2_X1 U2515 ( .A1(n3356), .A2(n3451), .ZN(n2229) );
  INV_X1 U2516 ( .A(n3356), .ZN(n2226) );
  INV_X1 U2517 ( .A(n3371), .ZN(n2225) );
  OR2_X1 U2518 ( .A1(n3457), .A2(n2228), .ZN(n2222) );
  INV_X1 U2519 ( .A(n3358), .ZN(n3404) );
  NAND2_X1 U2520 ( .A1(n2055), .A2(REG2_REG_2__SCAN_IN), .ZN(n2096) );
  INV_X1 U2521 ( .A(n3905), .ZN(n2661) );
  OAI211_X1 U2522 ( .C1(n4054), .C2(n2124), .A(n3599), .B(n2123), .ZN(n2617)
         );
  NAND2_X1 U2523 ( .A1(n2125), .A2(n4053), .ZN(n2123) );
  NOR2_X1 U2524 ( .A1(n3712), .A2(n2126), .ZN(n2125) );
  NAND2_X1 U2525 ( .A1(n4054), .A2(n3655), .ZN(n2127) );
  OR2_X1 U2526 ( .A1(n2108), .A2(n2110), .ZN(n3673) );
  INV_X1 U2527 ( .A(n3870), .ZN(n3383) );
  NOR2_X1 U2528 ( .A1(n2661), .A2(n2618), .ZN(n2141) );
  NOR2_X1 U2529 ( .A1(n4215), .A2(n4056), .ZN(n2145) );
  NOR2_X1 U2530 ( .A1(n4119), .A2(n2438), .ZN(n2439) );
  NOR2_X1 U2531 ( .A1(n2188), .A2(n2187), .ZN(n2186) );
  NAND2_X1 U2532 ( .A1(n2190), .A2(n2275), .ZN(n2187) );
  INV_X1 U2533 ( .A(IR_REG_5__SCAN_IN), .ZN(n2247) );
  INV_X1 U2534 ( .A(IR_REG_11__SCAN_IN), .ZN(n2434) );
  NOR2_X1 U2535 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2384)
         );
  INV_X1 U2536 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2391) );
  NAND2_X1 U2537 ( .A1(n3557), .A2(n2238), .ZN(n2237) );
  NAND2_X1 U2538 ( .A1(n2081), .A2(n2213), .ZN(n2212) );
  NAND2_X1 U2539 ( .A1(n3566), .A2(n2214), .ZN(n2213) );
  INV_X1 U2540 ( .A(n3474), .ZN(n2214) );
  NOR2_X1 U2541 ( .A1(n2500), .A2(n3517), .ZN(n2506) );
  AND2_X1 U2542 ( .A1(n2506), .A2(REG3_REG_21__SCAN_IN), .ZN(n2513) );
  INV_X1 U2543 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2414) );
  NAND2_X1 U2544 ( .A1(n3290), .A2(n3291), .ZN(n3464) );
  AOI21_X1 U2545 ( .B1(n2236), .B2(n3329), .A(n2234), .ZN(n2233) );
  INV_X1 U2546 ( .A(n3338), .ZN(n2234) );
  INV_X1 U2547 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3517) );
  AOI21_X1 U2548 ( .B1(n2255), .B2(n2253), .A(n2252), .ZN(n2251) );
  INV_X1 U2549 ( .A(n2255), .ZN(n2254) );
  INV_X1 U2550 ( .A(n3463), .ZN(n2252) );
  OR2_X1 U2551 ( .A1(n3457), .A2(n3451), .ZN(n3534) );
  INV_X1 U2552 ( .A(n3433), .ZN(n2249) );
  OR3_X1 U2553 ( .A1(n2931), .A2(n4496), .A3(n2847), .ZN(n2841) );
  AND4_X1 U2554 ( .A1(n2405), .A2(n2404), .A3(n2403), .A4(n2402), .ZN(n4253)
         );
  AND2_X1 U2555 ( .A1(n2097), .A2(n2095), .ZN(n2869) );
  NAND2_X1 U2556 ( .A1(n2871), .A2(n3758), .ZN(n2097) );
  INV_X1 U2557 ( .A(n2870), .ZN(n2095) );
  OAI21_X1 U2558 ( .B1(n2055), .B2(REG2_REG_2__SCAN_IN), .A(n2096), .ZN(n2870)
         );
  NOR2_X1 U2559 ( .A1(n2869), .A2(n2094), .ZN(n2756) );
  INV_X1 U2560 ( .A(n2096), .ZN(n2094) );
  NAND2_X1 U2561 ( .A1(n2880), .A2(n2159), .ZN(n2158) );
  XNOR2_X1 U2562 ( .A(n3771), .B(n3793), .ZN(n3772) );
  OAI21_X1 U2563 ( .B1(n3772), .B2(n4478), .A(n2099), .ZN(n4372) );
  NAND2_X1 U2564 ( .A1(n2100), .A2(n2151), .ZN(n2099) );
  INV_X1 U2565 ( .A(n3771), .ZN(n2100) );
  OR2_X1 U2566 ( .A1(n4423), .A2(n3780), .ZN(n2093) );
  AND2_X1 U2567 ( .A1(n3591), .A2(n2739), .ZN(n2746) );
  AND2_X1 U2568 ( .A1(n2746), .A2(n2745), .ZN(n2768) );
  OR2_X1 U2569 ( .A1(n2178), .A2(n3943), .ZN(n2176) );
  OR2_X1 U2570 ( .A1(n2178), .A2(n2180), .ZN(n2175) );
  OR2_X1 U2571 ( .A1(n2261), .A2(n2179), .ZN(n2178) );
  INV_X1 U2572 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U2573 ( .A1(n3942), .A2(n2183), .ZN(n2177) );
  INV_X1 U2574 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3444) );
  AND2_X1 U2575 ( .A1(n3656), .A2(n3915), .ZN(n3949) );
  NAND2_X1 U2576 ( .A1(n2127), .A2(n2125), .ZN(n3953) );
  INV_X1 U2577 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2489) );
  OR2_X1 U2578 ( .A1(n2490), .A2(n2489), .ZN(n2500) );
  INV_X1 U2579 ( .A(n4014), .ZN(n4023) );
  AND2_X1 U2580 ( .A1(n2471), .A2(n2470), .ZN(n2479) );
  NAND2_X1 U2581 ( .A1(n2127), .A2(n3595), .ZN(n4030) );
  NOR2_X1 U2582 ( .A1(n2450), .A2(n2449), .ZN(n2471) );
  NAND2_X1 U2583 ( .A1(n2604), .A2(n3704), .ZN(n4082) );
  AOI21_X1 U2584 ( .B1(n2116), .B2(n2118), .A(n2115), .ZN(n2114) );
  NOR2_X1 U2585 ( .A1(n2415), .A2(n2414), .ZN(n2426) );
  OAI21_X1 U2586 ( .B1(n2377), .B2(n2171), .A(n2168), .ZN(n3259) );
  AOI21_X1 U2587 ( .B1(n2170), .B2(n2169), .A(n2076), .ZN(n2168) );
  OR2_X1 U2588 ( .A1(n2392), .A2(n2391), .ZN(n2400) );
  INV_X1 U2589 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2399) );
  AND2_X1 U2590 ( .A1(n4104), .A2(n4107), .ZN(n3650) );
  OAI21_X1 U2591 ( .B1(n2597), .B2(n2118), .A(n2116), .ZN(n4106) );
  NAND2_X1 U2592 ( .A1(n2597), .A2(n3684), .ZN(n3243) );
  AOI21_X1 U2593 ( .B1(n2165), .B2(n2060), .A(n2072), .ZN(n2164) );
  NAND2_X1 U2594 ( .A1(n2979), .A2(n2161), .ZN(n2163) );
  NOR2_X1 U2595 ( .A1(n2162), .A2(n2352), .ZN(n2161) );
  INV_X1 U2596 ( .A(n2341), .ZN(n2162) );
  AND2_X1 U2597 ( .A1(n2593), .A2(n3683), .ZN(n3680) );
  AND2_X1 U2598 ( .A1(n3673), .A2(n3670), .ZN(n3649) );
  NAND2_X1 U2599 ( .A1(n2292), .A2(n2855), .ZN(n2299) );
  NAND2_X1 U2600 ( .A1(n2697), .A2(n2589), .ZN(n2949) );
  NAND2_X1 U2601 ( .A1(n2306), .A2(REG3_REG_2__SCAN_IN), .ZN(n2300) );
  NAND2_X1 U2602 ( .A1(n2580), .A2(n3818), .ZN(n4088) );
  NAND2_X1 U2603 ( .A1(n2916), .A2(n2732), .ZN(n2839) );
  INV_X1 U2604 ( .A(n3609), .ZN(n2129) );
  NAND2_X1 U2605 ( .A1(n3608), .A2(n3612), .ZN(n2130) );
  NAND2_X1 U2606 ( .A1(n2626), .A2(n3735), .ZN(n4145) );
  NOR2_X1 U2607 ( .A1(n4154), .A2(n4157), .ZN(n4153) );
  AND2_X1 U2608 ( .A1(n2053), .A2(DATAI_30_), .ZN(n4157) );
  NAND2_X1 U2609 ( .A1(n2053), .A2(DATAI_28_), .ZN(n3419) );
  NAND2_X1 U2610 ( .A1(n3937), .A2(n2141), .ZN(n3904) );
  NAND2_X1 U2611 ( .A1(n2053), .A2(DATAI_24_), .ZN(n3905) );
  NAND2_X1 U2612 ( .A1(n3937), .A2(n3923), .ZN(n3922) );
  AND2_X1 U2613 ( .A1(n3956), .A2(n3939), .ZN(n3937) );
  NOR2_X1 U2614 ( .A1(n3985), .A2(n4195), .ZN(n3956) );
  INV_X1 U2615 ( .A(n3958), .ZN(n4195) );
  AND2_X1 U2616 ( .A1(n2053), .A2(DATAI_20_), .ZN(n3983) );
  OR2_X1 U2617 ( .A1(n4001), .A2(n3983), .ZN(n3985) );
  NOR2_X1 U2618 ( .A1(n4070), .A2(n2144), .ZN(n4020) );
  NAND2_X1 U2619 ( .A1(n4023), .A2(n2145), .ZN(n2144) );
  NAND2_X1 U2620 ( .A1(n4020), .A2(n4002), .ZN(n4001) );
  NOR2_X1 U2621 ( .A1(n4070), .A2(n2143), .ZN(n4034) );
  INV_X1 U2622 ( .A(n2145), .ZN(n2143) );
  INV_X1 U2623 ( .A(n4227), .ZN(n4071) );
  NAND2_X1 U2624 ( .A1(n4090), .A2(n4071), .ZN(n4070) );
  OR2_X1 U2625 ( .A1(n4132), .A2(n3530), .ZN(n4121) );
  OR2_X1 U2626 ( .A1(n4130), .A2(n4248), .ZN(n4132) );
  INV_X1 U2627 ( .A(n3244), .ZN(n3251) );
  AND2_X1 U2628 ( .A1(n3073), .A2(n2061), .ZN(n3252) );
  NAND2_X1 U2629 ( .A1(n3073), .A2(n2142), .ZN(n3200) );
  NAND2_X1 U2630 ( .A1(n3073), .A2(n3120), .ZN(n3199) );
  AND2_X1 U2631 ( .A1(n3052), .A2(n3100), .ZN(n3073) );
  OR2_X1 U2632 ( .A1(n2988), .A2(n2983), .ZN(n3010) );
  NOR2_X1 U2633 ( .A1(n3010), .A2(n3062), .ZN(n3052) );
  NOR2_X1 U2634 ( .A1(n2955), .A2(n3551), .ZN(n3042) );
  AND2_X1 U2635 ( .A1(n2889), .A2(n4355), .ZN(n4249) );
  INV_X1 U2636 ( .A(n4261), .ZN(n4161) );
  INV_X1 U2637 ( .A(n2705), .ZN(n2828) );
  NOR2_X1 U2638 ( .A1(n2120), .A2(n2241), .ZN(n2119) );
  NOR2_X1 U2639 ( .A1(n2289), .A2(IR_REG_27__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U2640 ( .A1(n2289), .A2(IR_REG_31__SCAN_IN), .ZN(n2683) );
  INV_X1 U2641 ( .A(IR_REG_25__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U2642 ( .A1(n2637), .A2(IR_REG_31__SCAN_IN), .ZN(n2635) );
  XNOR2_X1 U2643 ( .A(n2643), .B(n2644), .ZN(n2915) );
  XNOR2_X1 U2644 ( .A(n2572), .B(n2571), .ZN(n2837) );
  XNOR2_X1 U2645 ( .A(n2574), .B(n2189), .ZN(n2645) );
  INV_X1 U2646 ( .A(IR_REG_20__SCAN_IN), .ZN(n2578) );
  INV_X1 U2647 ( .A(IR_REG_17__SCAN_IN), .ZN(n2274) );
  INV_X1 U2648 ( .A(n2335), .ZN(n2246) );
  AND2_X1 U2649 ( .A1(n2468), .A2(n2461), .ZN(n3786) );
  OR2_X1 U2650 ( .A1(n2387), .A2(IR_REG_9__SCAN_IN), .ZN(n2436) );
  INV_X1 U2651 ( .A(IR_REG_8__SCAN_IN), .ZN(n4688) );
  NAND2_X1 U2652 ( .A1(n2150), .A2(n2148), .ZN(n2755) );
  NOR2_X1 U2653 ( .A1(n2288), .A2(n2149), .ZN(n2148) );
  NAND2_X1 U2654 ( .A1(n2075), .A2(IR_REG_1__SCAN_IN), .ZN(n2150) );
  NOR2_X1 U2655 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2149)
         );
  INV_X1 U2656 ( .A(n4235), .ZN(n4092) );
  NAND2_X1 U2657 ( .A1(n3534), .A2(n3356), .ZN(n3535) );
  NAND2_X1 U2658 ( .A1(n3545), .A2(n2930), .ZN(n2964) );
  XNOR2_X1 U2659 ( .A(n2966), .B(n2937), .ZN(n2963) );
  AND2_X1 U2660 ( .A1(n3829), .A2(n2562), .ZN(n3426) );
  NAND2_X1 U2661 ( .A1(n2852), .A2(n2851), .ZN(n2853) );
  INV_X1 U2662 ( .A(n3753), .ZN(n3123) );
  NAND2_X1 U2663 ( .A1(n3022), .A2(n3021), .ZN(n3026) );
  AND4_X1 U2664 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .ZN(n3498)
         );
  AND4_X1 U2665 ( .A1(n2371), .A2(n2370), .A3(n2369), .A4(n2368), .ZN(n3194)
         );
  INV_X1 U2666 ( .A(n2822), .ZN(n2891) );
  AND4_X1 U2667 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(n3899)
         );
  AND4_X1 U2668 ( .A1(n2511), .A2(n2510), .A3(n2509), .A4(n2508), .ZN(n3936)
         );
  INV_X1 U2669 ( .A(n3584), .ZN(n3550) );
  NOR2_X1 U2670 ( .A1(n2923), .A2(n2922), .ZN(n3546) );
  INV_X1 U2671 ( .A(n3585), .ZN(n3553) );
  AND4_X1 U2672 ( .A1(n2357), .A2(n2356), .A3(n2355), .A4(n2354), .ZN(n3121)
         );
  NAND2_X1 U2673 ( .A1(n2053), .A2(DATAI_26_), .ZN(n3870) );
  AND4_X1 U2674 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n4231)
         );
  AND4_X1 U2675 ( .A1(n2467), .A2(n2466), .A3(n2465), .A4(n2464), .ZN(n4219)
         );
  NAND2_X1 U2676 ( .A1(n2856), .A2(n2861), .ZN(n3585) );
  NAND2_X1 U2677 ( .A1(n2856), .A2(n2843), .ZN(n3584) );
  INV_X1 U2678 ( .A(n3570), .ZN(n3587) );
  INV_X1 U2679 ( .A(n3574), .ZN(n3590) );
  OAI211_X1 U2680 ( .C1(n3397), .C2(n2059), .A(n2549), .B(n2548), .ZN(n3745)
         );
  NAND2_X1 U2681 ( .A1(n2539), .A2(n2538), .ZN(n3901) );
  AND3_X1 U2682 ( .A1(n2537), .A2(n2536), .A3(n2535), .ZN(n2539) );
  OR2_X1 U2683 ( .A1(n2533), .A2(n2532), .ZN(n3746) );
  INV_X1 U2684 ( .A(n3936), .ZN(n3976) );
  INV_X1 U2685 ( .A(n3498), .ZN(n4216) );
  INV_X1 U2686 ( .A(n4253), .ZN(n4137) );
  INV_X1 U2687 ( .A(n3194), .ZN(n3751) );
  INV_X1 U2688 ( .A(n3121), .ZN(n3752) );
  NOR2_X1 U2689 ( .A1(n2109), .A2(n2112), .ZN(n2106) );
  INV_X1 U2690 ( .A(n2110), .ZN(n2107) );
  OR2_X1 U2691 ( .A1(n2916), .A2(n4496), .ZN(n3755) );
  OAI21_X1 U2692 ( .B1(n2755), .B2(REG2_REG_1__SCAN_IN), .A(n2098), .ZN(n3759)
         );
  NAND2_X1 U2693 ( .A1(n2755), .A2(REG2_REG_1__SCAN_IN), .ZN(n2098) );
  NAND2_X1 U2694 ( .A1(n3759), .A2(n3760), .ZN(n3758) );
  XNOR2_X1 U2695 ( .A(n2755), .B(REG1_REG_1__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U2696 ( .A1(n3763), .A2(n3762), .ZN(n3761) );
  NOR2_X1 U2697 ( .A1(n2800), .A2(n2799), .ZN(n2798) );
  INV_X1 U2698 ( .A(n2153), .ZN(n2787) );
  NAND2_X1 U2699 ( .A1(n2154), .A2(n4358), .ZN(n2152) );
  AND2_X1 U2700 ( .A1(n2192), .A2(n2196), .ZN(n2812) );
  NAND2_X1 U2701 ( .A1(n2191), .A2(n2193), .ZN(n2810) );
  NAND2_X1 U2702 ( .A1(n2783), .A2(REG2_REG_6__SCAN_IN), .ZN(n2192) );
  XNOR2_X1 U2703 ( .A(n3792), .B(n2151), .ZN(n3795) );
  NAND2_X1 U2704 ( .A1(n4379), .A2(n3775), .ZN(n4392) );
  NAND2_X1 U2705 ( .A1(n4400), .A2(n3778), .ZN(n4413) );
  INV_X1 U2706 ( .A(n2091), .ZN(n4432) );
  INV_X1 U2707 ( .A(n2093), .ZN(n4434) );
  NOR2_X1 U2708 ( .A1(n4449), .A2(n3810), .ZN(n4459) );
  NAND2_X1 U2709 ( .A1(n4444), .A2(n3783), .ZN(n4453) );
  OR2_X1 U2710 ( .A1(n2561), .A2(n2560), .ZN(n3829) );
  INV_X1 U2711 ( .A(n2686), .ZN(n2136) );
  NAND2_X1 U2712 ( .A1(n2624), .A2(n2623), .ZN(n3840) );
  NAND2_X1 U2713 ( .A1(n3942), .A2(n2520), .ZN(n3913) );
  NAND2_X1 U2714 ( .A1(n2166), .A2(n2167), .ZN(n4011) );
  NOR2_X1 U2715 ( .A1(n4047), .A2(n2264), .ZN(n4033) );
  NAND2_X1 U2716 ( .A1(n2172), .A2(n2390), .ZN(n3242) );
  NAND2_X1 U2717 ( .A1(n2377), .A2(n2173), .ZN(n2172) );
  AOI21_X1 U2718 ( .B1(n2979), .B2(n2341), .A(n2060), .ZN(n3049) );
  INV_X1 U2719 ( .A(n4476), .ZN(n4486) );
  INV_X1 U2720 ( .A(n4142), .ZN(n4488) );
  INV_X1 U2721 ( .A(n2855), .ZN(n2904) );
  OR2_X1 U2722 ( .A1(n2839), .A2(n2707), .ZN(n4476) );
  NOR2_X1 U2723 ( .A1(n4494), .A2(n3008), .ZN(n4489) );
  OR2_X1 U2724 ( .A1(n3273), .A2(n4348), .ZN(n2664) );
  OR2_X1 U2725 ( .A1(n3850), .A2(n3849), .ZN(n4283) );
  INV_X1 U2726 ( .A(n4496), .ZN(n2732) );
  INV_X1 U2727 ( .A(n2843), .ZN(n2861) );
  NAND2_X1 U2728 ( .A1(n2915), .A2(STATE_REG_SCAN_IN), .ZN(n4496) );
  AND2_X1 U2729 ( .A1(n2409), .A2(n2421), .ZN(n4511) );
  AND2_X1 U2730 ( .A1(n2372), .A2(n2362), .ZN(n4357) );
  AND2_X1 U2731 ( .A1(n2323), .A2(n2315), .ZN(n4360) );
  OAI211_X1 U2732 ( .C1(n2215), .C2(n2209), .A(n2207), .B(n3401), .ZN(U3211)
         );
  NAND2_X1 U2733 ( .A1(n2210), .A2(n2219), .ZN(n2209) );
  INV_X1 U2734 ( .A(n2198), .ZN(n4473) );
  OAI21_X1 U2735 ( .B1(n4464), .B2(n2200), .A(n2199), .ZN(n2198) );
  XNOR2_X1 U2736 ( .A(n2104), .B(n3784), .ZN(n3822) );
  AOI21_X1 U2737 ( .B1(n2137), .B2(n2134), .A(n2087), .ZN(n2133) );
  AND2_X1 U2738 ( .A1(n2670), .A2(n2669), .ZN(n2671) );
  AND2_X1 U2739 ( .A1(n3093), .A2(n3023), .ZN(n2060) );
  NAND2_X1 U2740 ( .A1(n2237), .A2(n2235), .ZN(n3330) );
  AND2_X1 U2741 ( .A1(n2142), .A2(n3151), .ZN(n2061) );
  AND2_X1 U2742 ( .A1(n2972), .A2(n2967), .ZN(n2062) );
  OR2_X1 U2743 ( .A1(n3899), .A2(n3923), .ZN(n2063) );
  OR2_X1 U2744 ( .A1(n4057), .A2(n4215), .ZN(n2064) );
  AND2_X1 U2745 ( .A1(n2219), .A2(n2212), .ZN(n2065) );
  OR2_X1 U2746 ( .A1(n2667), .A2(n2705), .ZN(n4533) );
  OR2_X1 U2747 ( .A1(n2842), .A2(n2832), .ZN(n3576) );
  INV_X1 U2748 ( .A(n3576), .ZN(n3582) );
  AND2_X1 U2749 ( .A1(n2141), .A2(n3885), .ZN(n2066) );
  NOR2_X1 U2750 ( .A1(n2335), .A2(IR_REG_5__SCAN_IN), .ZN(n2334) );
  NOR2_X1 U2751 ( .A1(n2573), .A2(IR_REG_21__SCAN_IN), .ZN(n2569) );
  NOR2_X1 U2752 ( .A1(n2283), .A2(n4350), .ZN(n2067) );
  NAND2_X1 U2753 ( .A1(n3835), .A2(n2550), .ZN(n2068) );
  NAND2_X1 U2754 ( .A1(n2156), .A2(n2155), .ZN(n2154) );
  NAND2_X1 U2755 ( .A1(n3322), .A2(n3493), .ZN(n3557) );
  AND2_X1 U2756 ( .A1(n3828), .A2(n4523), .ZN(n2069) );
  OR2_X1 U2757 ( .A1(n3749), .A2(n3244), .ZN(n2070) );
  INV_X1 U2758 ( .A(n3126), .ZN(n3120) );
  NAND2_X1 U2759 ( .A1(n2496), .A2(n2275), .ZN(n2573) );
  NAND2_X1 U2760 ( .A1(n2105), .A2(n2726), .ZN(n2283) );
  INV_X1 U2761 ( .A(n2283), .ZN(n2282) );
  NOR2_X1 U2762 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2288)
         );
  NAND2_X1 U2763 ( .A1(n2138), .A2(n2136), .ZN(n2071) );
  NOR2_X1 U2764 ( .A1(n3753), .A2(n3096), .ZN(n2072) );
  AND2_X1 U2765 ( .A1(n3330), .A2(n3329), .ZN(n2073) );
  INV_X1 U2766 ( .A(n2309), .ZN(n2112) );
  OR2_X1 U2767 ( .A1(n2798), .A2(n2103), .ZN(n2102) );
  AND2_X1 U2768 ( .A1(n2363), .A2(n2164), .ZN(n2074) );
  INV_X1 U2769 ( .A(n2171), .ZN(n2170) );
  NAND2_X1 U2770 ( .A1(n2390), .A2(n2070), .ZN(n2171) );
  AND2_X1 U2771 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2075)
         );
  NOR2_X1 U2772 ( .A1(n4262), .A2(n3251), .ZN(n2076) );
  NAND2_X1 U2773 ( .A1(n2230), .A2(n2233), .ZN(n3453) );
  AND3_X1 U2774 ( .A1(n2244), .A2(n2246), .A3(n2119), .ZN(n2077) );
  AND2_X1 U2775 ( .A1(n2246), .A2(n2121), .ZN(n2078) );
  INV_X1 U2776 ( .A(n2311), .ZN(n2109) );
  INV_X1 U2777 ( .A(IR_REG_2__SCAN_IN), .ZN(n2205) );
  INV_X1 U2778 ( .A(IR_REG_31__SCAN_IN), .ZN(n2725) );
  INV_X1 U2779 ( .A(IR_REG_0__SCAN_IN), .ZN(n2140) );
  INV_X1 U2780 ( .A(n3793), .ZN(n2151) );
  OR2_X1 U2781 ( .A1(n2633), .A2(n2725), .ZN(n2643) );
  AND3_X1 U2782 ( .A1(n2246), .A2(n2272), .A3(n2247), .ZN(n2079) );
  INV_X1 U2783 ( .A(IR_REG_21__SCAN_IN), .ZN(n2189) );
  INV_X1 U2784 ( .A(n3473), .ZN(n2217) );
  AND2_X1 U2785 ( .A1(n3899), .A2(n3923), .ZN(n2080) );
  INV_X1 U2786 ( .A(n3331), .ZN(n3329) );
  NAND2_X1 U2787 ( .A1(n3391), .A2(n3390), .ZN(n2081) );
  NOR2_X1 U2788 ( .A1(n4017), .A2(n4036), .ZN(n2082) );
  INV_X1 U2789 ( .A(n2211), .ZN(n2210) );
  OAI21_X1 U2790 ( .B1(n2212), .B2(n2219), .A(n3582), .ZN(n2211) );
  INV_X1 U2791 ( .A(IR_REG_27__SCAN_IN), .ZN(n2243) );
  INV_X1 U2792 ( .A(n2236), .ZN(n2235) );
  NOR2_X1 U2793 ( .A1(n2240), .A2(n2239), .ZN(n2236) );
  AND2_X1 U2794 ( .A1(n2167), .A2(n2487), .ZN(n2083) );
  NAND2_X1 U2795 ( .A1(n3301), .A2(n3300), .ZN(n3431) );
  NOR2_X1 U2796 ( .A1(n3433), .A2(n3307), .ZN(n2084) );
  INV_X1 U2797 ( .A(n2228), .ZN(n2227) );
  NAND2_X1 U2798 ( .A1(n2229), .A2(n3363), .ZN(n2228) );
  INV_X1 U2799 ( .A(IR_REG_22__SCAN_IN), .ZN(n2571) );
  OR2_X1 U2800 ( .A1(IR_REG_29__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2085)
         );
  INV_X1 U2801 ( .A(IR_REG_29__SCAN_IN), .ZN(n2242) );
  NAND2_X1 U2802 ( .A1(n4357), .A2(REG2_REG_7__SCAN_IN), .ZN(n2086) );
  INV_X1 U2803 ( .A(n3595), .ZN(n2126) );
  NAND2_X1 U2804 ( .A1(n2074), .A2(n2163), .ZN(n3078) );
  INV_X2 U2805 ( .A(n4528), .ZN(n4530) );
  INV_X1 U2806 ( .A(n4411), .ZN(n4463) );
  NAND2_X1 U2807 ( .A1(n2968), .A2(n2967), .ZN(n2970) );
  NAND2_X1 U2808 ( .A1(n2246), .A2(n2244), .ZN(n2477) );
  NAND2_X1 U2809 ( .A1(n2163), .A2(n2164), .ZN(n3079) );
  INV_X1 U2810 ( .A(n2146), .ZN(n4049) );
  NOR2_X1 U2811 ( .A1(n4070), .A2(n4056), .ZN(n2146) );
  INV_X1 U2812 ( .A(n2618), .ZN(n3923) );
  AND2_X1 U2813 ( .A1(n2053), .A2(DATAI_23_), .ZN(n2618) );
  AND2_X1 U2814 ( .A1(n4533), .A2(n2688), .ZN(n2087) );
  NAND2_X1 U2815 ( .A1(n2053), .A2(DATAI_25_), .ZN(n3885) );
  NAND2_X1 U2816 ( .A1(n3786), .A2(REG2_REG_15__SCAN_IN), .ZN(n2088) );
  AND2_X1 U2817 ( .A1(n4498), .A2(REG2_REG_18__SCAN_IN), .ZN(n2089) );
  OR2_X1 U2818 ( .A1(n4474), .A2(n4647), .ZN(n2090) );
  AND2_X1 U2819 ( .A1(n4006), .A2(n3009), .ZN(n4149) );
  NAND3_X1 U2820 ( .A1(n2311), .A2(n3045), .A3(n2309), .ZN(n2108) );
  NAND2_X1 U2821 ( .A1(n2597), .A2(n2116), .ZN(n2113) );
  NAND2_X1 U2822 ( .A1(n2113), .A2(n2114), .ZN(n2604) );
  AND2_X2 U2823 ( .A1(n2078), .A2(n2244), .ZN(n2496) );
  NAND3_X1 U2824 ( .A1(n2244), .A2(n2246), .A3(n2274), .ZN(n2485) );
  NAND2_X1 U2825 ( .A1(n2138), .A2(n2137), .ZN(n2692) );
  NAND3_X1 U2826 ( .A1(n2139), .A2(n2140), .A3(n2205), .ZN(n2312) );
  INV_X1 U2827 ( .A(n2158), .ZN(n2797) );
  INV_X1 U2828 ( .A(n2156), .ZN(n2795) );
  INV_X1 U2829 ( .A(n2154), .ZN(n2752) );
  NAND2_X1 U2830 ( .A1(n2751), .A2(n2760), .ZN(n2159) );
  INV_X1 U2831 ( .A(n2352), .ZN(n2165) );
  NAND2_X1 U2832 ( .A1(n2166), .A2(n2083), .ZN(n4009) );
  NAND2_X1 U2833 ( .A1(n2377), .A2(n2376), .ZN(n3176) );
  INV_X1 U2834 ( .A(n2376), .ZN(n2174) );
  OAI21_X1 U2835 ( .B1(n3944), .B2(n2176), .A(n2175), .ZN(n2674) );
  NAND2_X1 U2836 ( .A1(n2496), .A2(n2186), .ZN(n2280) );
  NAND2_X1 U2837 ( .A1(n2102), .A2(n4358), .ZN(n2196) );
  NOR2_X1 U2838 ( .A1(n2288), .A2(n2725), .ZN(n2206) );
  NAND2_X1 U2839 ( .A1(n2215), .A2(n2208), .ZN(n2207) );
  NAND2_X1 U2840 ( .A1(n2215), .A2(n2212), .ZN(n3403) );
  AOI21_X1 U2841 ( .B1(n3476), .B2(n3473), .A(n3474), .ZN(n3565) );
  NAND2_X1 U2842 ( .A1(n2854), .A2(n2853), .ZN(n2221) );
  NAND3_X1 U2843 ( .A1(n2221), .A2(n3547), .A3(n2220), .ZN(n3545) );
  NAND2_X1 U2844 ( .A1(n3457), .A2(n3356), .ZN(n2223) );
  NAND2_X1 U2845 ( .A1(n2222), .A2(n2224), .ZN(n3374) );
  NAND2_X1 U2846 ( .A1(n3557), .A2(n2231), .ZN(n2230) );
  NAND2_X1 U2847 ( .A1(n2968), .A2(n2062), .ZN(n3022) );
  NAND3_X1 U2848 ( .A1(n2582), .A2(n2243), .A3(n2242), .ZN(n2241) );
  NAND3_X1 U2849 ( .A1(n3301), .A2(n3300), .A3(n2249), .ZN(n2248) );
  NAND2_X1 U2850 ( .A1(n2248), .A2(n3306), .ZN(n3579) );
  NAND3_X1 U2851 ( .A1(n3301), .A2(n3300), .A3(n2084), .ZN(n3482) );
  NAND3_X1 U2852 ( .A1(n2250), .A2(n3579), .A3(n3486), .ZN(n3316) );
  OAI21_X1 U2853 ( .B1(n3284), .B2(n2258), .A(n2257), .ZN(n3466) );
  XNOR2_X1 U2854 ( .A(n2674), .B(n2673), .ZN(n3281) );
  AND2_X1 U2855 ( .A1(n2921), .A2(n2920), .ZN(n2922) );
  NAND2_X1 U2856 ( .A1(n3299), .A2(n3298), .ZN(n3300) );
  NAND2_X1 U2857 ( .A1(n3297), .A2(n3296), .ZN(n3301) );
  INV_X1 U2858 ( .A(n3523), .ZN(n3299) );
  NAND2_X1 U2859 ( .A1(n3523), .A2(n3524), .ZN(n3297) );
  AND2_X2 U2860 ( .A1(n2708), .A2(n4476), .ZN(n4494) );
  INV_X1 U2861 ( .A(n4196), .ZN(n3458) );
  OR2_X1 U2862 ( .A1(n3978), .A2(n4002), .ZN(n2259) );
  AND2_X1 U2863 ( .A1(n2313), .A2(n2267), .ZN(n2260) );
  NOR2_X1 U2864 ( .A1(n2559), .A2(n2558), .ZN(n2261) );
  INV_X1 U2865 ( .A(n3650), .ZN(n2411) );
  AND2_X1 U2866 ( .A1(n4251), .A2(n3530), .ZN(n2263) );
  NAND2_X1 U2867 ( .A1(n2053), .A2(DATAI_22_), .ZN(n3939) );
  INV_X1 U2868 ( .A(n3939), .ZN(n2519) );
  NAND2_X1 U2869 ( .A1(n2298), .A2(n2855), .ZN(n2589) );
  AND2_X1 U2870 ( .A1(n4228), .A2(n4056), .ZN(n2264) );
  OR2_X1 U2871 ( .A1(n3830), .A2(n4348), .ZN(n2265) );
  OR2_X1 U2872 ( .A1(n3830), .A2(n4272), .ZN(n2266) );
  INV_X1 U2873 ( .A(IR_REG_4__SCAN_IN), .ZN(n2267) );
  INV_X1 U2874 ( .A(n3680), .ZN(n2363) );
  AND2_X1 U2875 ( .A1(n2276), .A2(n2262), .ZN(n2277) );
  INV_X1 U2876 ( .A(n3524), .ZN(n3298) );
  AND2_X1 U2877 ( .A1(n3615), .A2(n3613), .ZN(n3630) );
  NAND2_X1 U2878 ( .A1(n3978), .A2(n4002), .ZN(n2498) );
  NAND2_X1 U2879 ( .A1(n3671), .A2(n3668), .ZN(n3642) );
  INV_X1 U2880 ( .A(n2965), .ZN(n2937) );
  OAI22_X1 U2881 ( .A1(n2298), .A2(n3358), .B1(n2931), .B2(n2904), .ZN(n2920)
         );
  INV_X1 U2882 ( .A(n2971), .ZN(n2972) );
  INV_X1 U2883 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2365) );
  INV_X1 U2884 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2440) );
  NAND2_X1 U2885 ( .A1(n2067), .A2(REG1_REG_1__SCAN_IN), .ZN(n2285) );
  OR2_X1 U2886 ( .A1(n2521), .A2(n3444), .ZN(n2527) );
  INV_X1 U2887 ( .A(n3651), .ZN(n2325) );
  AND2_X1 U2888 ( .A1(n2053), .A2(DATAI_27_), .ZN(n4160) );
  INV_X1 U2889 ( .A(n3096), .ZN(n3100) );
  INV_X1 U2890 ( .A(n4163), .ZN(n4250) );
  INV_X1 U2891 ( .A(n2829), .ZN(n2738) );
  INV_X1 U2892 ( .A(n2569), .ZN(n2570) );
  NAND2_X1 U2893 ( .A1(n2850), .A2(n3407), .ZN(n2852) );
  AND3_X1 U2894 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2342) );
  AND2_X1 U2895 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2470) );
  AOI22_X1 U2896 ( .A1(n3756), .A2(n3294), .B1(n2932), .B2(n2822), .ZN(n2850)
         );
  INV_X1 U2897 ( .A(n3749), .ZN(n4262) );
  INV_X1 U2898 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2449) );
  NOR2_X1 U2899 ( .A1(n2542), .A2(n2541), .ZN(n2546) );
  INV_X1 U2900 ( .A(IR_REG_28__SCAN_IN), .ZN(n2582) );
  INV_X1 U2901 ( .A(n2766), .ZN(n2860) );
  INV_X1 U2902 ( .A(n3746), .ZN(n4178) );
  AOI21_X1 U2903 ( .B1(n4069), .B2(n2463), .A(n2462), .ZN(n4045) );
  INV_X1 U2904 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2688) );
  INV_X1 U2905 ( .A(n4249), .ZN(n4113) );
  INV_X1 U2906 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2693) );
  INV_X1 U2907 ( .A(n3885), .ZN(n4174) );
  INV_X1 U2908 ( .A(DATAI_19_), .ZN(n4691) );
  INV_X1 U2909 ( .A(n4145), .ZN(n4117) );
  NAND2_X1 U2910 ( .A1(n2861), .A2(n2738), .ZN(n4261) );
  INV_X1 U2911 ( .A(IR_REG_24__SCAN_IN), .ZN(n2630) );
  AND2_X1 U2912 ( .A1(n2342), .A2(REG3_REG_6__SCAN_IN), .ZN(n2353) );
  INV_X1 U2913 ( .A(n3330), .ZN(n3332) );
  INV_X1 U2914 ( .A(n3023), .ZN(n3062) );
  OAI21_X1 U2915 ( .B1(n2821), .B2(n3358), .A(n2820), .ZN(n2825) );
  OR2_X1 U2916 ( .A1(n2400), .A2(n2399), .ZN(n2415) );
  AND3_X1 U2917 ( .A1(n2565), .A2(n2564), .A3(n2563), .ZN(n2566) );
  AND4_X1 U2918 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n3978)
         );
  INV_X1 U2919 ( .A(n3093), .ZN(n3103) );
  AND2_X1 U2920 ( .A1(n2294), .A2(n2293), .ZN(n2297) );
  XNOR2_X1 U2921 ( .A(n2583), .B(n2582), .ZN(n2843) );
  AND2_X1 U2922 ( .A1(n2768), .A2(n3739), .ZN(n4411) );
  OR2_X1 U2923 ( .A1(n3609), .A2(n2568), .ZN(n2673) );
  NAND2_X1 U2926 ( .A1(n4533), .A2(REG1_REG_28__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U2927 ( .A1(n2660), .A2(n2731), .ZN(n2705) );
  NAND2_X1 U2928 ( .A1(n3591), .A2(DATAI_21_), .ZN(n3958) );
  INV_X1 U2929 ( .A(n3262), .ZN(n3267) );
  NAND2_X1 U2930 ( .A1(n4088), .A2(n4263), .ZN(n4523) );
  AND2_X1 U2931 ( .A1(n2979), .A2(n2981), .ZN(n4521) );
  AND2_X1 U2932 ( .A1(n2894), .A2(n2837), .ZN(n4520) );
  INV_X1 U2933 ( .A(n2839), .ZN(n2838) );
  AND2_X1 U2934 ( .A1(n2740), .A2(n2745), .ZN(n4467) );
  NAND2_X1 U2935 ( .A1(n2567), .A2(n2566), .ZN(n3843) );
  INV_X1 U2936 ( .A(n3978), .ZN(n4015) );
  NAND2_X1 U2937 ( .A1(n2768), .A2(n2843), .ZN(n4475) );
  OR2_X1 U2938 ( .A1(n4024), .A2(n2711), .ZN(n4142) );
  INV_X1 U2939 ( .A(n4149), .ZN(n4063) );
  INV_X2 U2940 ( .A(n4533), .ZN(n4536) );
  AND2_X1 U2941 ( .A1(n2664), .A2(n2663), .ZN(n2665) );
  OR2_X1 U2942 ( .A1(n2667), .A2(n2828), .ZN(n4528) );
  INV_X1 U2943 ( .A(n4537), .ZN(n4495) );
  INV_X1 U2944 ( .A(D_REG_1__SCAN_IN), .ZN(n2737) );
  NAND2_X1 U2945 ( .A1(n2730), .A2(n2838), .ZN(n4537) );
  INV_X1 U2946 ( .A(n2837), .ZN(n4353) );
  AND2_X1 U2947 ( .A1(n2388), .A2(n2436), .ZN(n4366) );
  INV_X2 U2948 ( .A(n3755), .ZN(U4043) );
  OR4_X1 U2949 ( .A1(n2716), .A2(n2715), .A3(n2714), .A4(n2713), .ZN(U3289) );
  NAND2_X1 U2950 ( .A1(n2666), .A2(n2665), .ZN(U3514) );
  NAND2_X1 U2951 ( .A1(n2268), .A2(n2260), .ZN(n2335) );
  NOR2_X1 U2952 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2271)
         );
  NOR2_X1 U2953 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2270)
         );
  NOR2_X1 U2954 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2269)
         );
  AND2_X1 U2955 ( .A1(n2632), .A2(n2571), .ZN(n2276) );
  INV_X1 U2956 ( .A(n2279), .ZN(n2726) );
  NAND2_X1 U2957 ( .A1(n2280), .A2(IR_REG_31__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2958 ( .A1(n2307), .A2(REG0_REG_1__SCAN_IN), .ZN(n2287) );
  NAND2_X1 U2959 ( .A1(n2306), .A2(REG3_REG_1__SCAN_IN), .ZN(n2286) );
  NAND2_X1 U2960 ( .A1(n2308), .A2(REG2_REG_1__SCAN_IN), .ZN(n2284) );
  INV_X1 U2961 ( .A(n2298), .ZN(n2292) );
  INV_X1 U2962 ( .A(n2755), .ZN(n4362) );
  NAND2_X1 U2963 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2291) );
  NAND2_X1 U2964 ( .A1(n2243), .A2(n2582), .ZN(n2290) );
  MUX2_X1 U2965 ( .A(n2291), .B(n2290), .S(n2683), .Z(n2410) );
  MUX2_X1 U2966 ( .A(n4362), .B(DATAI_1_), .S(n2410), .Z(n2855) );
  NAND2_X1 U2967 ( .A1(n2292), .A2(n2904), .ZN(n3665) );
  NAND2_X1 U2968 ( .A1(n3665), .A2(n2589), .ZN(n2588) );
  NAND2_X1 U2969 ( .A1(n2308), .A2(REG2_REG_0__SCAN_IN), .ZN(n2294) );
  NAND2_X1 U2970 ( .A1(n2307), .A2(REG0_REG_0__SCAN_IN), .ZN(n2293) );
  NAND2_X1 U2971 ( .A1(n2067), .A2(REG1_REG_0__SCAN_IN), .ZN(n2296) );
  NAND2_X1 U2972 ( .A1(n2306), .A2(REG3_REG_0__SCAN_IN), .ZN(n2295) );
  MUX2_X1 U2973 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2410), .Z(n2822) );
  AND2_X1 U2974 ( .A1(n3756), .A2(n2822), .ZN(n2700) );
  NAND2_X1 U2975 ( .A1(n2588), .A2(n2700), .ZN(n2699) );
  NAND2_X1 U2976 ( .A1(n2699), .A2(n2299), .ZN(n2945) );
  INV_X1 U2977 ( .A(n2945), .ZN(n2304) );
  NAND2_X1 U2978 ( .A1(n2054), .A2(REG0_REG_2__SCAN_IN), .ZN(n2303) );
  NAND2_X1 U2979 ( .A1(n2067), .A2(REG1_REG_2__SCAN_IN), .ZN(n2302) );
  NAND2_X1 U2980 ( .A1(n2308), .A2(REG2_REG_2__SCAN_IN), .ZN(n2301) );
  MUX2_X1 U2981 ( .A(n2055), .B(DATAI_2_), .S(n2410), .Z(n3551) );
  INV_X1 U2982 ( .A(n3551), .ZN(n2924) );
  NAND2_X1 U2983 ( .A1(n3036), .A2(n2924), .ZN(n3671) );
  NAND2_X1 U2984 ( .A1(n2939), .A2(n3551), .ZN(n3668) );
  NAND2_X1 U2985 ( .A1(n2304), .A2(n3642), .ZN(n2944) );
  NAND2_X1 U2986 ( .A1(n2939), .A2(n2924), .ZN(n2305) );
  NAND2_X1 U2987 ( .A1(n2944), .A2(n2305), .ZN(n3032) );
  OR2_X1 U2988 ( .A1(n2059), .A2(REG3_REG_3__SCAN_IN), .ZN(n2311) );
  NAND2_X1 U2989 ( .A1(n2452), .A2(REG1_REG_3__SCAN_IN), .ZN(n2310) );
  NAND2_X1 U2990 ( .A1(n2308), .A2(REG2_REG_3__SCAN_IN), .ZN(n2309) );
  NAND2_X1 U2991 ( .A1(n2312), .A2(IR_REG_31__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U2992 ( .A1(n2314), .A2(n2313), .ZN(n2323) );
  OR2_X1 U2993 ( .A1(n2314), .A2(n2313), .ZN(n2315) );
  MUX2_X1 U2994 ( .A(n4360), .B(DATAI_3_), .S(n3591), .Z(n3045) );
  NAND2_X1 U2995 ( .A1(n3549), .A2(n3045), .ZN(n2316) );
  NAND2_X1 U2996 ( .A1(n3032), .A2(n2316), .ZN(n2318) );
  NAND2_X1 U2997 ( .A1(n2974), .A2(n2936), .ZN(n2317) );
  NAND2_X1 U2998 ( .A1(n2318), .A2(n2317), .ZN(n2980) );
  INV_X1 U2999 ( .A(n2980), .ZN(n2326) );
  NAND2_X1 U3000 ( .A1(n2308), .A2(REG2_REG_4__SCAN_IN), .ZN(n2322) );
  NAND2_X1 U3001 ( .A1(n2534), .A2(REG0_REG_4__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U3002 ( .A1(n2452), .A2(REG1_REG_4__SCAN_IN), .ZN(n2320) );
  XNOR2_X1 U3003 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n2990) );
  NAND2_X1 U3004 ( .A1(n2323), .A2(IR_REG_31__SCAN_IN), .ZN(n2324) );
  XNOR2_X1 U3005 ( .A(n2324), .B(IR_REG_4__SCAN_IN), .ZN(n2760) );
  MUX2_X1 U3006 ( .A(n2760), .B(DATAI_4_), .S(n2053), .Z(n2983) );
  NAND2_X1 U3007 ( .A1(n3065), .A2(n2983), .ZN(n3674) );
  INV_X1 U3008 ( .A(n2983), .ZN(n2989) );
  NAND2_X1 U3009 ( .A1(n3754), .A2(n2989), .ZN(n3678) );
  NAND2_X1 U3010 ( .A1(n2326), .A2(n2325), .ZN(n2979) );
  NAND2_X1 U3011 ( .A1(n3754), .A2(n2983), .ZN(n3006) );
  NAND2_X1 U3012 ( .A1(n2534), .A2(REG0_REG_5__SCAN_IN), .ZN(n2333) );
  NAND2_X1 U3013 ( .A1(n2452), .A2(REG1_REG_5__SCAN_IN), .ZN(n2332) );
  NAND2_X1 U3014 ( .A1(n2308), .A2(REG2_REG_5__SCAN_IN), .ZN(n2331) );
  INV_X1 U3015 ( .A(n2342), .ZN(n2344) );
  INV_X1 U3016 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2328) );
  NAND2_X1 U3017 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2327) );
  NAND2_X1 U3018 ( .A1(n2328), .A2(n2327), .ZN(n2329) );
  NAND2_X1 U3019 ( .A1(n2344), .A2(n2329), .ZN(n3031) );
  OR2_X1 U3020 ( .A1(n2059), .A2(n3031), .ZN(n2330) );
  INV_X1 U3021 ( .A(n2334), .ZN(n2338) );
  NAND2_X1 U3022 ( .A1(n2335), .A2(IR_REG_31__SCAN_IN), .ZN(n2336) );
  MUX2_X1 U3023 ( .A(IR_REG_31__SCAN_IN), .B(n2336), .S(IR_REG_5__SCAN_IN), 
        .Z(n2337) );
  NAND2_X1 U3024 ( .A1(n2338), .A2(n2337), .ZN(n2802) );
  INV_X1 U3025 ( .A(DATAI_5_), .ZN(n2339) );
  MUX2_X1 U3026 ( .A(n2802), .B(n2339), .S(n2053), .Z(n3023) );
  NAND2_X1 U3027 ( .A1(n3103), .A2(n3062), .ZN(n2340) );
  AND2_X1 U3028 ( .A1(n3006), .A2(n2340), .ZN(n2341) );
  INV_X1 U3029 ( .A(n2353), .ZN(n2346) );
  INV_X1 U3030 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2343) );
  NAND2_X1 U3031 ( .A1(n2344), .A2(n2343), .ZN(n2345) );
  NAND2_X1 U3032 ( .A1(n2346), .A2(n2345), .ZN(n3099) );
  OR2_X1 U3033 ( .A1(n2059), .A2(n3099), .ZN(n2350) );
  NAND2_X1 U3034 ( .A1(n2308), .A2(REG2_REG_6__SCAN_IN), .ZN(n2349) );
  NAND2_X1 U3035 ( .A1(n2534), .A2(REG0_REG_6__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U3036 ( .A1(n2452), .A2(REG1_REG_6__SCAN_IN), .ZN(n2347) );
  NAND4_X1 U3037 ( .A1(n2350), .A2(n2349), .A3(n2348), .A4(n2347), .ZN(n3753)
         );
  OR2_X1 U3038 ( .A1(n2334), .A2(n2725), .ZN(n2351) );
  XNOR2_X1 U3039 ( .A(n2351), .B(IR_REG_6__SCAN_IN), .ZN(n4358) );
  MUX2_X1 U3040 ( .A(n4358), .B(DATAI_6_), .S(n2053), .Z(n3096) );
  AND2_X1 U3041 ( .A1(n3753), .A2(n3096), .ZN(n2352) );
  NAND2_X1 U3042 ( .A1(n2308), .A2(REG2_REG_7__SCAN_IN), .ZN(n2357) );
  NAND2_X1 U3043 ( .A1(n2534), .A2(REG0_REG_7__SCAN_IN), .ZN(n2356) );
  NAND2_X1 U3044 ( .A1(n2452), .A2(REG1_REG_7__SCAN_IN), .ZN(n2355) );
  NAND2_X1 U3045 ( .A1(n2353), .A2(REG3_REG_7__SCAN_IN), .ZN(n2366) );
  OAI21_X1 U3046 ( .B1(n2353), .B2(REG3_REG_7__SCAN_IN), .A(n2366), .ZN(n3129)
         );
  OR2_X1 U3047 ( .A1(n2059), .A2(n3129), .ZN(n2354) );
  INV_X1 U3048 ( .A(IR_REG_6__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U3049 ( .A1(n2334), .A2(n2358), .ZN(n2359) );
  NAND2_X1 U3050 ( .A1(n2359), .A2(IR_REG_31__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U3051 ( .A1(n2361), .A2(n2360), .ZN(n2372) );
  OR2_X1 U3052 ( .A1(n2361), .A2(n2360), .ZN(n2362) );
  MUX2_X1 U3053 ( .A(n4357), .B(DATAI_7_), .S(n2053), .Z(n3126) );
  NAND2_X1 U3054 ( .A1(n3121), .A2(n3126), .ZN(n2593) );
  NAND2_X1 U3055 ( .A1(n3752), .A2(n3120), .ZN(n3683) );
  NAND2_X1 U3056 ( .A1(n3752), .A2(n3126), .ZN(n2364) );
  NAND2_X1 U3057 ( .A1(n3078), .A2(n2364), .ZN(n3203) );
  NAND2_X1 U3058 ( .A1(n2534), .A2(REG0_REG_8__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3059 ( .A1(n2452), .A2(REG1_REG_8__SCAN_IN), .ZN(n2370) );
  NAND2_X1 U3060 ( .A1(n2308), .A2(REG2_REG_8__SCAN_IN), .ZN(n2369) );
  AND2_X1 U3061 ( .A1(n2366), .A2(n2365), .ZN(n2367) );
  NOR2_X1 U3062 ( .A1(n2366), .A2(n2365), .ZN(n2378) );
  OR2_X1 U3063 ( .A1(n2367), .A2(n2378), .ZN(n4477) );
  OR2_X1 U3064 ( .A1(n2059), .A2(n4477), .ZN(n2368) );
  NAND2_X1 U3065 ( .A1(n2372), .A2(IR_REG_31__SCAN_IN), .ZN(n2373) );
  XNOR2_X1 U3066 ( .A(n2373), .B(n4688), .ZN(n3793) );
  INV_X1 U3067 ( .A(DATAI_8_), .ZN(n2374) );
  MUX2_X1 U3068 ( .A(n3793), .B(n2374), .S(n2053), .Z(n3201) );
  NAND2_X1 U3069 ( .A1(n3194), .A2(n3201), .ZN(n2375) );
  NAND2_X1 U3070 ( .A1(n3203), .A2(n2375), .ZN(n2377) );
  NAND2_X1 U3071 ( .A1(n3751), .A2(n3205), .ZN(n2376) );
  NAND2_X1 U3072 ( .A1(n2378), .A2(REG3_REG_9__SCAN_IN), .ZN(n2392) );
  OR2_X1 U3073 ( .A1(n2378), .A2(REG3_REG_9__SCAN_IN), .ZN(n2379) );
  NAND2_X1 U3074 ( .A1(n2392), .A2(n2379), .ZN(n3198) );
  OR2_X1 U3075 ( .A1(n2059), .A2(n3198), .ZN(n2383) );
  NAND2_X1 U3076 ( .A1(n2534), .A2(REG0_REG_9__SCAN_IN), .ZN(n2382) );
  NAND2_X1 U3077 ( .A1(n2452), .A2(REG1_REG_9__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3078 ( .A1(n2308), .A2(REG2_REG_9__SCAN_IN), .ZN(n2380) );
  NAND4_X1 U3079 ( .A1(n2383), .A2(n2382), .A3(n2381), .A4(n2380), .ZN(n3750)
         );
  AND2_X1 U3080 ( .A1(n2384), .A2(n4688), .ZN(n2385) );
  NAND2_X1 U3081 ( .A1(n2334), .A2(n2385), .ZN(n2387) );
  NAND2_X1 U3082 ( .A1(n2387), .A2(IR_REG_31__SCAN_IN), .ZN(n2386) );
  MUX2_X1 U3083 ( .A(IR_REG_31__SCAN_IN), .B(n2386), .S(IR_REG_9__SCAN_IN), 
        .Z(n2388) );
  MUX2_X1 U3084 ( .A(n4366), .B(DATAI_9_), .S(n2053), .Z(n3229) );
  AND2_X1 U3085 ( .A1(n3750), .A2(n3229), .ZN(n2389) );
  INV_X1 U3086 ( .A(n3229), .ZN(n3151) );
  NAND2_X1 U3087 ( .A1(n3246), .A2(n3151), .ZN(n2390) );
  NAND2_X1 U3088 ( .A1(n2392), .A2(n2391), .ZN(n2393) );
  NAND2_X1 U3089 ( .A1(n2400), .A2(n2393), .ZN(n3253) );
  OR2_X1 U3090 ( .A1(n2059), .A2(n3253), .ZN(n2397) );
  NAND2_X1 U3091 ( .A1(n2534), .A2(REG0_REG_10__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U3092 ( .A1(n2452), .A2(REG1_REG_10__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3093 ( .A1(n2308), .A2(REG2_REG_10__SCAN_IN), .ZN(n2394) );
  NAND4_X1 U3094 ( .A1(n2397), .A2(n2396), .A3(n2395), .A4(n2394), .ZN(n3749)
         );
  NAND2_X1 U3095 ( .A1(n2436), .A2(IR_REG_31__SCAN_IN), .ZN(n2398) );
  XNOR2_X1 U3096 ( .A(n2398), .B(IR_REG_10__SCAN_IN), .ZN(n3797) );
  MUX2_X1 U3097 ( .A(n3797), .B(DATAI_10_), .S(n2053), .Z(n3244) );
  INV_X1 U3098 ( .A(n3259), .ZN(n2412) );
  NAND2_X1 U3099 ( .A1(n2534), .A2(REG0_REG_11__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3100 ( .A1(n2452), .A2(REG1_REG_11__SCAN_IN), .ZN(n2404) );
  NAND2_X1 U3101 ( .A1(n2308), .A2(REG2_REG_11__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U3102 ( .A1(n2400), .A2(n2399), .ZN(n2401) );
  NAND2_X1 U3103 ( .A1(n2415), .A2(n2401), .ZN(n3266) );
  OR2_X1 U3104 ( .A1(n2059), .A2(n3266), .ZN(n2402) );
  NAND2_X1 U3105 ( .A1(n2406), .A2(IR_REG_31__SCAN_IN), .ZN(n2408) );
  INV_X1 U3106 ( .A(n2408), .ZN(n2407) );
  NAND2_X1 U3107 ( .A1(n2407), .A2(IR_REG_11__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U3108 ( .A1(n2408), .A2(n2434), .ZN(n2421) );
  MUX2_X1 U3109 ( .A(n4511), .B(DATAI_11_), .S(n2053), .Z(n3262) );
  NAND2_X1 U3110 ( .A1(n4253), .A2(n3262), .ZN(n4104) );
  NAND2_X1 U3111 ( .A1(n4137), .A2(n3267), .ZN(n4107) );
  NAND2_X1 U3112 ( .A1(n2412), .A2(n2411), .ZN(n3260) );
  NAND2_X1 U3113 ( .A1(n4253), .A2(n3267), .ZN(n2413) );
  NAND2_X1 U3114 ( .A1(n3260), .A2(n2413), .ZN(n4129) );
  AND2_X1 U3115 ( .A1(n2415), .A2(n2414), .ZN(n2416) );
  OR2_X1 U3116 ( .A1(n2416), .A2(n2426), .ZN(n4133) );
  OR2_X1 U3117 ( .A1(n2059), .A2(n4133), .ZN(n2420) );
  NAND2_X1 U3118 ( .A1(n2308), .A2(REG2_REG_12__SCAN_IN), .ZN(n2419) );
  NAND2_X1 U3119 ( .A1(n2534), .A2(REG0_REG_12__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U3120 ( .A1(n2452), .A2(REG1_REG_12__SCAN_IN), .ZN(n2417) );
  NAND4_X1 U3121 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .ZN(n4115)
         );
  NAND2_X1 U3122 ( .A1(n2421), .A2(IR_REG_31__SCAN_IN), .ZN(n2422) );
  XNOR2_X1 U3123 ( .A(n2422), .B(IR_REG_12__SCAN_IN), .ZN(n3801) );
  MUX2_X1 U3124 ( .A(n3801), .B(DATAI_12_), .S(n2053), .Z(n4248) );
  NAND2_X1 U3125 ( .A1(n4115), .A2(n4248), .ZN(n2423) );
  NAND2_X1 U3126 ( .A1(n4129), .A2(n2423), .ZN(n2425) );
  INV_X1 U3127 ( .A(n4115), .ZN(n3528) );
  INV_X1 U3128 ( .A(n4248), .ZN(n3468) );
  NAND2_X1 U3129 ( .A1(n3528), .A2(n3468), .ZN(n2424) );
  NAND2_X1 U3130 ( .A1(n2425), .A2(n2424), .ZN(n4119) );
  NAND2_X1 U3131 ( .A1(n2426), .A2(REG3_REG_13__SCAN_IN), .ZN(n2441) );
  OR2_X1 U3132 ( .A1(n2426), .A2(REG3_REG_13__SCAN_IN), .ZN(n2427) );
  NAND2_X1 U3133 ( .A1(n2441), .A2(n2427), .ZN(n4124) );
  OR2_X1 U3134 ( .A1(n2059), .A2(n4124), .ZN(n2431) );
  NAND2_X1 U3135 ( .A1(n2308), .A2(REG2_REG_13__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U3136 ( .A1(n2534), .A2(REG0_REG_13__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U3137 ( .A1(n2452), .A2(REG1_REG_13__SCAN_IN), .ZN(n2428) );
  NAND4_X1 U3138 ( .A1(n2431), .A2(n2430), .A3(n2429), .A4(n2428), .ZN(n4251)
         );
  INV_X1 U3139 ( .A(IR_REG_10__SCAN_IN), .ZN(n2433) );
  INV_X1 U3140 ( .A(IR_REG_12__SCAN_IN), .ZN(n2432) );
  NAND3_X1 U3141 ( .A1(n2434), .A2(n2433), .A3(n2432), .ZN(n2435) );
  OAI21_X1 U3142 ( .B1(n2436), .B2(n2435), .A(IR_REG_31__SCAN_IN), .ZN(n2437)
         );
  XNOR2_X1 U3143 ( .A(n2437), .B(IR_REG_13__SCAN_IN), .ZN(n3788) );
  MUX2_X1 U3144 ( .A(n3788), .B(DATAI_13_), .S(n2053), .Z(n3530) );
  NOR2_X1 U3145 ( .A1(n4251), .A2(n3530), .ZN(n2438) );
  NOR2_X1 U3146 ( .A1(n2439), .A2(n2263), .ZN(n4081) );
  NAND2_X1 U3147 ( .A1(n2534), .A2(REG0_REG_14__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U31480 ( .A1(n2452), .A2(REG1_REG_14__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U31490 ( .A1(n2308), .A2(REG2_REG_14__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3150 ( .A1(n2441), .A2(n2440), .ZN(n2442) );
  NAND2_X1 U3151 ( .A1(n2450), .A2(n2442), .ZN(n3436) );
  OR2_X1 U3152 ( .A1(n2059), .A2(n3436), .ZN(n2443) );
  OR2_X1 U3153 ( .A1(n2079), .A2(n2725), .ZN(n2447) );
  XNOR2_X1 U3154 ( .A(n2447), .B(IR_REG_14__SCAN_IN), .ZN(n3805) );
  MUX2_X1 U3155 ( .A(n3805), .B(DATAI_14_), .S(n2053), .Z(n4235) );
  NAND2_X1 U3156 ( .A1(n4231), .A2(n4235), .ZN(n4064) );
  INV_X1 U3157 ( .A(n4231), .ZN(n3748) );
  NAND2_X1 U3158 ( .A1(n3748), .A2(n4092), .ZN(n3592) );
  NAND2_X1 U3159 ( .A1(n4064), .A2(n3592), .ZN(n4085) );
  NAND2_X1 U3160 ( .A1(n4081), .A2(n4085), .ZN(n4080) );
  NAND2_X1 U3161 ( .A1(n4231), .A2(n4092), .ZN(n2448) );
  NAND2_X1 U3162 ( .A1(n4080), .A2(n2448), .ZN(n4069) );
  AND2_X1 U3163 ( .A1(n2450), .A2(n2449), .ZN(n2451) );
  OR2_X1 U3164 ( .A1(n2451), .A2(n2471), .ZN(n4072) );
  OR2_X1 U3165 ( .A1(n2059), .A2(n4072), .ZN(n2456) );
  NAND2_X1 U3166 ( .A1(n2308), .A2(REG2_REG_15__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U3167 ( .A1(n2534), .A2(REG0_REG_15__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U3168 ( .A1(n2452), .A2(REG1_REG_15__SCAN_IN), .ZN(n2453) );
  NAND4_X1 U3169 ( .A1(n2456), .A2(n2455), .A3(n2454), .A4(n2453), .ZN(n4236)
         );
  INV_X1 U3170 ( .A(IR_REG_14__SCAN_IN), .ZN(n2457) );
  NAND2_X1 U3171 ( .A1(n2079), .A2(n2457), .ZN(n2458) );
  NAND2_X1 U3172 ( .A1(n2458), .A2(IR_REG_31__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3173 ( .A1(n2460), .A2(n2459), .ZN(n2468) );
  OR2_X1 U3174 ( .A1(n2460), .A2(n2459), .ZN(n2461) );
  MUX2_X1 U3175 ( .A(n3786), .B(DATAI_15_), .S(n2053), .Z(n4227) );
  NAND2_X1 U3176 ( .A1(n4236), .A2(n4227), .ZN(n2463) );
  NOR2_X1 U3177 ( .A1(n4236), .A2(n4227), .ZN(n2462) );
  NAND2_X1 U3178 ( .A1(n2308), .A2(REG2_REG_16__SCAN_IN), .ZN(n2467) );
  NAND2_X1 U3179 ( .A1(n2534), .A2(REG0_REG_16__SCAN_IN), .ZN(n2466) );
  NAND2_X1 U3180 ( .A1(n2452), .A2(REG1_REG_16__SCAN_IN), .ZN(n2465) );
  XNOR2_X1 U3181 ( .A(n2471), .B(REG3_REG_16__SCAN_IN), .ZN(n4050) );
  OR2_X1 U3182 ( .A1(n2059), .A2(n4050), .ZN(n2464) );
  NAND2_X1 U3183 ( .A1(n2468), .A2(IR_REG_31__SCAN_IN), .ZN(n2469) );
  XNOR2_X1 U3184 ( .A(n2469), .B(IR_REG_16__SCAN_IN), .ZN(n4502) );
  MUX2_X1 U3185 ( .A(n4502), .B(DATAI_16_), .S(n2053), .Z(n4056) );
  NAND2_X1 U3186 ( .A1(n4219), .A2(n4056), .ZN(n3710) );
  INV_X1 U3187 ( .A(n4056), .ZN(n3488) );
  NAND2_X1 U3188 ( .A1(n4228), .A2(n3488), .ZN(n3595) );
  NAND2_X1 U3189 ( .A1(n3710), .A2(n3595), .ZN(n4053) );
  AOI21_X1 U3190 ( .B1(n2471), .B2(REG3_REG_16__SCAN_IN), .A(
        REG3_REG_17__SCAN_IN), .ZN(n2472) );
  OR2_X1 U3191 ( .A1(n2479), .A2(n2472), .ZN(n4037) );
  OR2_X1 U3192 ( .A1(n2059), .A2(n4037), .ZN(n2476) );
  NAND2_X1 U3193 ( .A1(n2534), .A2(REG0_REG_17__SCAN_IN), .ZN(n2475) );
  NAND2_X1 U3194 ( .A1(n2452), .A2(REG1_REG_17__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3195 ( .A1(n2308), .A2(REG2_REG_17__SCAN_IN), .ZN(n2473) );
  NAND4_X1 U3196 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(n2473), .ZN(n4057)
         );
  NAND2_X1 U3197 ( .A1(n2477), .A2(IR_REG_31__SCAN_IN), .ZN(n2478) );
  XNOR2_X1 U3198 ( .A(n2478), .B(IR_REG_17__SCAN_IN), .ZN(n3812) );
  MUX2_X1 U3199 ( .A(n3812), .B(DATAI_17_), .S(n2053), .Z(n4215) );
  INV_X1 U3200 ( .A(n4057), .ZN(n4017) );
  INV_X1 U3201 ( .A(n4215), .ZN(n4036) );
  NAND2_X1 U3202 ( .A1(n2534), .A2(REG0_REG_18__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3203 ( .A1(n2452), .A2(REG1_REG_18__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U3204 ( .A1(n2308), .A2(REG2_REG_18__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U3205 ( .A1(n2479), .A2(REG3_REG_18__SCAN_IN), .ZN(n2490) );
  OR2_X1 U3206 ( .A1(n2479), .A2(REG3_REG_18__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3207 ( .A1(n2490), .A2(n2480), .ZN(n4025) );
  OR2_X1 U3208 ( .A1(n2059), .A2(n4025), .ZN(n2481) );
  NAND2_X1 U3209 ( .A1(n2485), .A2(IR_REG_31__SCAN_IN), .ZN(n2486) );
  XNOR2_X1 U32100 ( .A(n2486), .B(IR_REG_18__SCAN_IN), .ZN(n4498) );
  MUX2_X1 U32110 ( .A(n4498), .B(DATAI_18_), .S(n2053), .Z(n4014) );
  NAND2_X1 U32120 ( .A1(n3498), .A2(n4014), .ZN(n3992) );
  NAND2_X1 U32130 ( .A1(n4216), .A2(n4023), .ZN(n3993) );
  NAND2_X1 U32140 ( .A1(n4009), .A2(n2488), .ZN(n3991) );
  NAND2_X1 U32150 ( .A1(n2308), .A2(REG2_REG_19__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U32160 ( .A1(n2534), .A2(REG0_REG_19__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U32170 ( .A1(n2452), .A2(REG1_REG_19__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U32180 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  NAND2_X1 U32190 ( .A1(n2500), .A2(n2491), .ZN(n4003) );
  OR2_X1 U32200 ( .A1(n2059), .A2(n4003), .ZN(n2492) );
  INV_X1 U32210 ( .A(n2496), .ZN(n2497) );
  MUX2_X1 U32220 ( .A(n3818), .B(n4691), .S(n2053), .Z(n4002) );
  NAND2_X1 U32230 ( .A1(n3991), .A2(n2259), .ZN(n2499) );
  INV_X1 U32240 ( .A(n4002), .ZN(n3647) );
  NAND2_X1 U32250 ( .A1(n2499), .A2(n2498), .ZN(n3968) );
  AND2_X1 U32260 ( .A1(n2500), .A2(n3517), .ZN(n2501) );
  OR2_X1 U32270 ( .A1(n2501), .A2(n2506), .ZN(n3516) );
  OR2_X1 U32280 ( .A1(n2059), .A2(n3516), .ZN(n2505) );
  NAND2_X1 U32290 ( .A1(n2308), .A2(REG2_REG_20__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U32300 ( .A1(n2534), .A2(REG0_REG_20__SCAN_IN), .ZN(n2503) );
  NAND2_X1 U32310 ( .A1(n2452), .A2(REG1_REG_20__SCAN_IN), .ZN(n2502) );
  NAND4_X1 U32320 ( .A1(n2505), .A2(n2504), .A3(n2503), .A4(n2502), .ZN(n3747)
         );
  NAND2_X1 U32330 ( .A1(n3747), .A2(n3983), .ZN(n3634) );
  NOR2_X1 U32340 ( .A1(n3747), .A2(n3983), .ZN(n3635) );
  NAND2_X1 U32350 ( .A1(n2308), .A2(REG2_REG_21__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U32360 ( .A1(n2534), .A2(REG0_REG_21__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U32370 ( .A1(n2452), .A2(REG1_REG_21__SCAN_IN), .ZN(n2509) );
  NOR2_X1 U32380 ( .A1(n2506), .A2(REG3_REG_21__SCAN_IN), .ZN(n2507) );
  OR2_X1 U32390 ( .A1(n2513), .A2(n2507), .ZN(n3960) );
  OR2_X1 U32400 ( .A1(n2059), .A2(n3960), .ZN(n2508) );
  NOR2_X1 U32410 ( .A1(n3936), .A2(n3958), .ZN(n2512) );
  OAI22_X1 U32420 ( .A1(n3950), .A2(n2512), .B1(n4195), .B2(n3976), .ZN(n3944)
         );
  NAND2_X1 U32430 ( .A1(n2513), .A2(REG3_REG_22__SCAN_IN), .ZN(n2521) );
  OR2_X1 U32440 ( .A1(n2513), .A2(REG3_REG_22__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U32450 ( .A1(n2521), .A2(n2514), .ZN(n3539) );
  OR2_X1 U32460 ( .A1(n2059), .A2(n3539), .ZN(n2518) );
  NAND2_X1 U32470 ( .A1(n2054), .A2(REG0_REG_22__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32480 ( .A1(n2452), .A2(REG1_REG_22__SCAN_IN), .ZN(n2516) );
  NAND2_X1 U32490 ( .A1(n2308), .A2(REG2_REG_22__SCAN_IN), .ZN(n2515) );
  NAND4_X1 U32500 ( .A1(n2518), .A2(n2517), .A3(n2516), .A4(n2515), .ZN(n4196)
         );
  NAND2_X1 U32510 ( .A1(n3458), .A2(n2519), .ZN(n3916) );
  NAND2_X1 U32520 ( .A1(n4196), .A2(n3939), .ZN(n2615) );
  NAND2_X1 U32530 ( .A1(n2308), .A2(REG2_REG_23__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U32540 ( .A1(n2054), .A2(REG0_REG_23__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U32550 ( .A1(n2452), .A2(REG1_REG_23__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U32560 ( .A1(n2521), .A2(n3444), .ZN(n2522) );
  NAND2_X1 U32570 ( .A1(n2527), .A2(n2522), .ZN(n3924) );
  OR2_X1 U32580 ( .A1(n2059), .A2(n3924), .ZN(n2523) );
  NAND2_X1 U32590 ( .A1(n2527), .A2(n4551), .ZN(n2528) );
  NAND2_X1 U32600 ( .A1(n2542), .A2(n2528), .ZN(n3907) );
  NAND2_X1 U32610 ( .A1(n2452), .A2(REG1_REG_24__SCAN_IN), .ZN(n2529) );
  OAI21_X1 U32620 ( .B1(n3907), .B2(n2059), .A(n2529), .ZN(n2533) );
  NAND2_X1 U32630 ( .A1(n2308), .A2(REG2_REG_24__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32640 ( .A1(n2534), .A2(REG0_REG_24__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U32650 ( .A1(n2531), .A2(n2530), .ZN(n2532) );
  NAND2_X1 U32660 ( .A1(n3746), .A2(n2661), .ZN(n3879) );
  NAND2_X1 U32670 ( .A1(n2452), .A2(REG1_REG_25__SCAN_IN), .ZN(n2537) );
  NAND2_X1 U32680 ( .A1(n2308), .A2(REG2_REG_25__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U32690 ( .A1(n2534), .A2(REG0_REG_25__SCAN_IN), .ZN(n2535) );
  XNOR2_X1 U32700 ( .A(n2542), .B(REG3_REG_25__SCAN_IN), .ZN(n3887) );
  NAND2_X1 U32710 ( .A1(n3887), .A2(n2306), .ZN(n2538) );
  NAND2_X1 U32720 ( .A1(n3901), .A2(n4174), .ZN(n2551) );
  AND2_X1 U32730 ( .A1(n3879), .A2(n2551), .ZN(n3855) );
  INV_X1 U32740 ( .A(n2542), .ZN(n2540) );
  AOI21_X1 U32750 ( .B1(n2540), .B2(REG3_REG_25__SCAN_IN), .A(
        REG3_REG_26__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U32760 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2541) );
  OR2_X1 U32770 ( .A1(n2543), .A2(n2546), .ZN(n3568) );
  AOI22_X1 U32780 ( .A1(n2308), .A2(REG2_REG_26__SCAN_IN), .B1(n2534), .B2(
        REG0_REG_26__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U32790 ( .A1(n2452), .A2(REG1_REG_26__SCAN_IN), .ZN(n2544) );
  OAI211_X2 U32800 ( .C1(n3568), .C2(n2059), .A(n2545), .B(n2544), .ZN(n4175)
         );
  INV_X1 U32810 ( .A(n4175), .ZN(n3847) );
  NOR2_X1 U32820 ( .A1(n3847), .A2(n3870), .ZN(n2555) );
  INV_X1 U32830 ( .A(n2555), .ZN(n3624) );
  AND2_X1 U32840 ( .A1(n3855), .A2(n3624), .ZN(n3835) );
  NAND2_X1 U32850 ( .A1(n2546), .A2(REG3_REG_27__SCAN_IN), .ZN(n2561) );
  OR2_X1 U32860 ( .A1(n2546), .A2(REG3_REG_27__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U32870 ( .A1(n2561), .A2(n2547), .ZN(n3397) );
  AOI22_X1 U32880 ( .A1(n2308), .A2(REG2_REG_27__SCAN_IN), .B1(n2054), .B2(
        REG0_REG_27__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U32890 ( .A1(n2452), .A2(REG1_REG_27__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32900 ( .A1(n3745), .A2(n4160), .ZN(n2550) );
  INV_X1 U32910 ( .A(n2550), .ZN(n2559) );
  OR2_X1 U32920 ( .A1(n3745), .A2(n4160), .ZN(n2557) );
  INV_X1 U32930 ( .A(n2551), .ZN(n2554) );
  NAND2_X1 U32940 ( .A1(n4178), .A2(n3905), .ZN(n3880) );
  OR2_X1 U32950 ( .A1(n3901), .A2(n4174), .ZN(n2552) );
  AND2_X1 U32960 ( .A1(n3880), .A2(n2552), .ZN(n2553) );
  OR2_X1 U32970 ( .A1(n2555), .A2(n3856), .ZN(n2556) );
  OR2_X1 U32980 ( .A1(n4175), .A2(n3383), .ZN(n3623) );
  AND2_X1 U32990 ( .A1(n2556), .A2(n3623), .ZN(n3836) );
  AND2_X1 U33000 ( .A1(n2557), .A2(n3836), .ZN(n2558) );
  INV_X1 U33010 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U33020 ( .A1(n2561), .A2(n2560), .ZN(n2562) );
  NAND2_X1 U33030 ( .A1(n3426), .A2(n2306), .ZN(n2567) );
  NAND2_X1 U33040 ( .A1(n2452), .A2(REG1_REG_28__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U33050 ( .A1(n2308), .A2(REG2_REG_28__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U33060 ( .A1(n2054), .A2(REG0_REG_28__SCAN_IN), .ZN(n2563) );
  NOR2_X1 U33070 ( .A1(n3843), .A2(n3419), .ZN(n3609) );
  NAND2_X1 U33080 ( .A1(n3843), .A2(n3419), .ZN(n3612) );
  INV_X1 U33090 ( .A(n3612), .ZN(n2568) );
  NAND2_X1 U33100 ( .A1(n2570), .A2(IR_REG_31__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U33110 ( .A1(n2573), .A2(IR_REG_31__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U33120 ( .A1(n2576), .A2(n2575), .ZN(n2577) );
  XNOR2_X1 U33130 ( .A(n4353), .B(n2846), .ZN(n2580) );
  AND2_X1 U33140 ( .A1(n3731), .A2(n4356), .ZN(n2894) );
  INV_X1 U33150 ( .A(n4520), .ZN(n4263) );
  INV_X1 U33160 ( .A(n4523), .ZN(n4213) );
  OR2_X1 U33170 ( .A1(n2581), .A2(n2725), .ZN(n2583) );
  NAND2_X1 U33180 ( .A1(n4353), .A2(n4354), .ZN(n2829) );
  AOI22_X1 U33190 ( .A1(n2308), .A2(REG2_REG_29__SCAN_IN), .B1(n2054), .B2(
        REG0_REG_29__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U33200 ( .A1(n2452), .A2(REG1_REG_29__SCAN_IN), .ZN(n2584) );
  OAI211_X1 U33210 ( .C1(n3829), .C2(n2059), .A(n2585), .B(n2584), .ZN(n3416)
         );
  INV_X1 U33220 ( .A(n3416), .ZN(n2586) );
  INV_X1 U33230 ( .A(n3731), .ZN(n4355) );
  OAI22_X1 U33240 ( .A1(n2586), .A2(n4163), .B1(n4113), .B2(n3419), .ZN(n2587)
         );
  AOI21_X1 U33250 ( .B1(n4161), .B2(n3745), .A(n2587), .ZN(n2628) );
  CLKBUF_X1 U33260 ( .A(n2588), .Z(n3640) );
  INV_X1 U33270 ( .A(n3756), .ZN(n2821) );
  NAND2_X1 U33280 ( .A1(n2821), .A2(n2822), .ZN(n3664) );
  INV_X1 U33290 ( .A(n3642), .ZN(n2950) );
  NAND2_X1 U33300 ( .A1(n2949), .A2(n2950), .ZN(n2948) );
  NAND2_X1 U33310 ( .A1(n2948), .A2(n3668), .ZN(n3034) );
  NAND2_X1 U33320 ( .A1(n3549), .A2(n2936), .ZN(n3670) );
  NAND2_X1 U33330 ( .A1(n3034), .A2(n3649), .ZN(n3033) );
  NAND2_X1 U33340 ( .A1(n3033), .A2(n3673), .ZN(n2982) );
  INV_X1 U33350 ( .A(n3674), .ZN(n2590) );
  OR2_X1 U33360 ( .A1(n2982), .A2(n2590), .ZN(n2591) );
  NAND2_X1 U33370 ( .A1(n2591), .A2(n3678), .ZN(n3004) );
  NAND2_X1 U33380 ( .A1(n3093), .A2(n3062), .ZN(n3692) );
  AND2_X1 U33390 ( .A1(n3103), .A2(n3023), .ZN(n3003) );
  NAND2_X1 U33400 ( .A1(n3753), .A2(n3100), .ZN(n3693) );
  NAND2_X1 U33410 ( .A1(n3050), .A2(n3693), .ZN(n2592) );
  NAND2_X1 U33420 ( .A1(n3123), .A2(n3096), .ZN(n3679) );
  NAND2_X1 U33430 ( .A1(n2592), .A2(n3679), .ZN(n3069) );
  INV_X1 U33440 ( .A(n2593), .ZN(n2594) );
  OR2_X1 U33450 ( .A1(n3069), .A2(n2594), .ZN(n2595) );
  NAND2_X1 U33460 ( .A1(n2595), .A2(n3683), .ZN(n3204) );
  NAND2_X1 U33470 ( .A1(n3194), .A2(n3205), .ZN(n3685) );
  NAND2_X1 U33480 ( .A1(n3204), .A2(n3685), .ZN(n2596) );
  NAND2_X1 U33490 ( .A1(n3751), .A2(n3201), .ZN(n3682) );
  NAND2_X1 U33500 ( .A1(n2596), .A2(n3682), .ZN(n3183) );
  AND2_X1 U33510 ( .A1(n3750), .A2(n3151), .ZN(n3690) );
  NAND2_X1 U33520 ( .A1(n3246), .A2(n3229), .ZN(n3684) );
  NAND2_X1 U3353 ( .A1(n3749), .A2(n3251), .ZN(n3700) );
  NAND2_X1 U33540 ( .A1(n4262), .A2(n3244), .ZN(n3699) );
  NAND2_X1 U3355 ( .A1(n4115), .A2(n3468), .ZN(n4109) );
  INV_X1 U3356 ( .A(n3530), .ZN(n4122) );
  NAND2_X1 U3357 ( .A1(n4251), .A2(n4122), .ZN(n2598) );
  NAND2_X1 U3358 ( .A1(n4109), .A2(n2598), .ZN(n2600) );
  INV_X1 U3359 ( .A(n4107), .ZN(n2599) );
  NOR2_X1 U3360 ( .A1(n2600), .A2(n2599), .ZN(n3701) );
  NAND2_X1 U3361 ( .A1(n3528), .A2(n4248), .ZN(n4111) );
  NAND2_X1 U3362 ( .A1(n4104), .A2(n4111), .ZN(n2603) );
  INV_X1 U3363 ( .A(n2600), .ZN(n2602) );
  NOR2_X1 U3364 ( .A1(n4251), .A2(n4122), .ZN(n2601) );
  AOI21_X1 U3365 ( .B1(n2603), .B2(n2602), .A(n2601), .ZN(n3704) );
  INV_X1 U3366 ( .A(n4085), .ZN(n2605) );
  NAND2_X1 U3367 ( .A1(n4082), .A2(n2605), .ZN(n4083) );
  INV_X1 U3368 ( .A(n4236), .ZN(n4060) );
  NAND2_X1 U3369 ( .A1(n4060), .A2(n4227), .ZN(n3594) );
  NAND2_X1 U3370 ( .A1(n4236), .A2(n4071), .ZN(n3593) );
  NAND2_X1 U3371 ( .A1(n3594), .A2(n3593), .ZN(n4068) );
  INV_X1 U3372 ( .A(n4064), .ZN(n2606) );
  NOR2_X1 U3373 ( .A1(n4068), .A2(n2606), .ZN(n2607) );
  NAND2_X1 U3374 ( .A1(n4083), .A2(n2607), .ZN(n2608) );
  NAND2_X1 U3375 ( .A1(n2608), .A2(n3593), .ZN(n4054) );
  INV_X1 U3376 ( .A(n4053), .ZN(n3655) );
  NAND2_X1 U3377 ( .A1(n4015), .A2(n4002), .ZN(n2609) );
  AND2_X1 U3378 ( .A1(n3993), .A2(n2609), .ZN(n3973) );
  NAND2_X1 U3379 ( .A1(n4057), .A2(n4036), .ZN(n3969) );
  INV_X1 U3380 ( .A(n3983), .ZN(n3518) );
  NAND2_X1 U3381 ( .A1(n3747), .A2(n3518), .ZN(n2613) );
  AND2_X1 U3382 ( .A1(n3969), .A2(n2613), .ZN(n2610) );
  NAND2_X1 U3383 ( .A1(n3973), .A2(n2610), .ZN(n3712) );
  INV_X1 U3384 ( .A(n3973), .ZN(n2611) );
  OAI22_X1 U3385 ( .A1(n2611), .A2(n3992), .B1(n4002), .B2(n4015), .ZN(n3972)
         );
  NAND2_X1 U3386 ( .A1(n4017), .A2(n4215), .ZN(n3970) );
  OAI22_X1 U3387 ( .A1(n2611), .A2(n3970), .B1(n3747), .B2(n3518), .ZN(n2612)
         );
  OR2_X1 U3388 ( .A1(n3972), .A2(n2612), .ZN(n2614) );
  NAND2_X1 U3389 ( .A1(n2614), .A2(n2613), .ZN(n3952) );
  NAND2_X1 U3390 ( .A1(n3936), .A2(n4195), .ZN(n3915) );
  AND2_X1 U3391 ( .A1(n3916), .A2(n3915), .ZN(n3716) );
  AND2_X1 U3392 ( .A1(n3952), .A2(n3716), .ZN(n3599) );
  AND2_X1 U3393 ( .A1(n3976), .A2(n3958), .ZN(n3717) );
  AND2_X1 U3394 ( .A1(n3916), .A2(n3717), .ZN(n3598) );
  OR2_X1 U3395 ( .A1(n3899), .A2(n2618), .ZN(n3637) );
  NAND2_X1 U3396 ( .A1(n3637), .A2(n2615), .ZN(n3601) );
  NOR2_X1 U3397 ( .A1(n3598), .A2(n3601), .ZN(n2616) );
  NAND2_X1 U3398 ( .A1(n2617), .A2(n2616), .ZN(n3896) );
  NAND2_X1 U3399 ( .A1(n4178), .A2(n2661), .ZN(n3632) );
  NAND2_X1 U3400 ( .A1(n3899), .A2(n2618), .ZN(n3895) );
  NAND2_X1 U3401 ( .A1(n3632), .A2(n3895), .ZN(n3721) );
  INV_X1 U3402 ( .A(n3721), .ZN(n2619) );
  NAND2_X1 U3403 ( .A1(n3896), .A2(n2619), .ZN(n2620) );
  NAND2_X1 U3404 ( .A1(n3746), .A2(n3905), .ZN(n3631) );
  NAND2_X1 U3405 ( .A1(n2620), .A2(n3631), .ZN(n3877) );
  NAND2_X1 U3406 ( .A1(n3901), .A2(n3885), .ZN(n3657) );
  INV_X1 U3407 ( .A(n3657), .ZN(n2621) );
  OR2_X1 U3408 ( .A1(n4175), .A2(n3870), .ZN(n2622) );
  OR2_X1 U3409 ( .A1(n3901), .A2(n3885), .ZN(n3860) );
  AND2_X1 U3410 ( .A1(n2622), .A2(n3860), .ZN(n3726) );
  NAND2_X1 U3411 ( .A1(n3861), .A2(n3726), .ZN(n2624) );
  AND2_X1 U3412 ( .A1(n4175), .A2(n3870), .ZN(n3614) );
  INV_X1 U3413 ( .A(n3614), .ZN(n2623) );
  XNOR2_X1 U3414 ( .A(n3745), .B(n4160), .ZN(n3629) );
  NOR2_X1 U3415 ( .A1(n3745), .A2(n3848), .ZN(n3608) );
  INV_X1 U3416 ( .A(n3608), .ZN(n2625) );
  INV_X1 U3417 ( .A(n2673), .ZN(n3645) );
  XNOR2_X1 U3418 ( .A(n2678), .B(n3645), .ZN(n2627) );
  NAND2_X1 U3419 ( .A1(n4353), .A2(n4356), .ZN(n2626) );
  NAND2_X1 U3420 ( .A1(n4354), .A2(n4355), .ZN(n3735) );
  NAND2_X1 U3421 ( .A1(n2627), .A2(n4145), .ZN(n3276) );
  OAI211_X1 U3422 ( .C1(n3281), .C2(n4213), .A(n2628), .B(n3276), .ZN(n2668)
         );
  NAND2_X1 U3423 ( .A1(n2643), .A2(n2644), .ZN(n2629) );
  NAND2_X1 U3424 ( .A1(n2633), .A2(n2632), .ZN(n2637) );
  NAND2_X1 U3425 ( .A1(n2640), .A2(n2641), .ZN(n2636) );
  MUX2_X1 U3426 ( .A(n2640), .B(n2636), .S(B_REG_SCAN_IN), .Z(n2639) );
  OAI21_X2 U3427 ( .B1(n2637), .B2(IR_REG_25__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2638) );
  NAND2_X1 U3428 ( .A1(n2729), .A2(n2737), .ZN(n2826) );
  INV_X1 U3429 ( .A(n2642), .ZN(n2735) );
  NAND2_X1 U3430 ( .A1(n2735), .A2(n2641), .ZN(n2702) );
  NAND2_X1 U3431 ( .A1(n2826), .A2(n2702), .ZN(n2659) );
  INV_X1 U3432 ( .A(n2640), .ZN(n4352) );
  NAND3_X2 U3433 ( .A1(n4352), .A2(n4351), .A3(n2642), .ZN(n2818) );
  NAND2_X1 U3434 ( .A1(n4520), .A2(n2645), .ZN(n2707) );
  AND2_X1 U3435 ( .A1(n3731), .A2(n3818), .ZN(n2646) );
  NAND2_X1 U3436 ( .A1(n2707), .A2(n2704), .ZN(n2647) );
  NOR2_X1 U3437 ( .A1(n2839), .A2(n2647), .ZN(n2658) );
  NOR4_X1 U3438 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2651) );
  NOR4_X1 U3439 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2650) );
  NOR4_X1 U3440 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2649) );
  NOR4_X1 U3441 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2648) );
  NAND4_X1 U3442 ( .A1(n2651), .A2(n2650), .A3(n2649), .A4(n2648), .ZN(n2657)
         );
  NOR2_X1 U3443 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_22__SCAN_IN), .ZN(n2655)
         );
  NOR4_X1 U3444 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2654) );
  NOR4_X1 U3445 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2653) );
  NOR4_X1 U3446 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2652) );
  NAND4_X1 U3447 ( .A1(n2655), .A2(n2654), .A3(n2653), .A4(n2652), .ZN(n2656)
         );
  OAI21_X1 U3448 ( .B1(n2657), .B2(n2656), .A(n2729), .ZN(n2703) );
  NAND3_X1 U3449 ( .A1(n2659), .A2(n2658), .A3(n2703), .ZN(n2667) );
  INV_X1 U3450 ( .A(D_REG_0__SCAN_IN), .ZN(n2734) );
  NAND2_X1 U3451 ( .A1(n2729), .A2(n2734), .ZN(n2660) );
  NAND2_X1 U3452 ( .A1(n2735), .A2(n2640), .ZN(n2731) );
  NAND2_X1 U3453 ( .A1(n2668), .A2(n4530), .ZN(n2666) );
  NAND2_X1 U3454 ( .A1(n2904), .A2(n2891), .ZN(n2955) );
  NAND2_X1 U3455 ( .A1(n3042), .A2(n2936), .ZN(n2988) );
  NAND2_X1 U3456 ( .A1(n3268), .A2(n3267), .ZN(n4130) );
  INV_X1 U3457 ( .A(n2690), .ZN(n2662) );
  OAI21_X1 U34580 ( .B1(n3850), .B2(n3419), .A(n2662), .ZN(n3273) );
  NAND2_X1 U34590 ( .A1(n4528), .A2(REG0_REG_28__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3460 ( .A1(n2668), .A2(n4536), .ZN(n2672) );
  NAND2_X1 U3461 ( .A1(n2672), .A2(n2671), .ZN(U3546) );
  NAND2_X1 U3462 ( .A1(n2674), .A2(n2673), .ZN(n2676) );
  INV_X1 U3463 ( .A(n3419), .ZN(n3409) );
  NAND2_X1 U3464 ( .A1(n3843), .A2(n3409), .ZN(n2675) );
  NAND2_X1 U3465 ( .A1(n2676), .A2(n2675), .ZN(n2677) );
  NAND2_X1 U3466 ( .A1(n3591), .A2(DATAI_29_), .ZN(n2689) );
  OR2_X1 U34670 ( .A1(n3416), .A2(n2689), .ZN(n3615) );
  NAND2_X1 U3468 ( .A1(n3416), .A2(n2689), .ZN(n3613) );
  XNOR2_X1 U34690 ( .A(n2677), .B(n3630), .ZN(n3828) );
  XOR2_X1 U3470 ( .A(n3630), .B(n2679), .Z(n2687) );
  INV_X1 U34710 ( .A(n3843), .ZN(n4164) );
  NAND2_X1 U3472 ( .A1(n2452), .A2(REG1_REG_30__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U34730 ( .A1(n2308), .A2(REG2_REG_30__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3474 ( .A1(n2054), .A2(REG0_REG_30__SCAN_IN), .ZN(n2680) );
  NAND3_X1 U34750 ( .A1(n2682), .A2(n2681), .A3(n2680), .ZN(n3744) );
  XNOR2_X1 U3476 ( .A(n2683), .B(IR_REG_27__SCAN_IN), .ZN(n2766) );
  AOI21_X1 U34770 ( .B1(n2766), .B2(B_REG_SCAN_IN), .A(n4163), .ZN(n3823) );
  INV_X1 U3478 ( .A(n2689), .ZN(n2684) );
  AOI22_X1 U34790 ( .A1(n3744), .A2(n3823), .B1(n4249), .B2(n2684), .ZN(n2685)
         );
  OAI21_X1 U3480 ( .B1(n4164), .B2(n4261), .A(n2685), .ZN(n2686) );
  NAND2_X1 U34810 ( .A1(n2691), .A2(n2266), .ZN(U3547) );
  OR2_X1 U3482 ( .A1(n2692), .A2(n4528), .ZN(n2695) );
  NAND2_X1 U34830 ( .A1(n4528), .A2(n2693), .ZN(n2694) );
  NAND2_X1 U3484 ( .A1(n2695), .A2(n2694), .ZN(n2696) );
  NAND2_X1 U34850 ( .A1(n2696), .A2(n2265), .ZN(U3515) );
  INV_X1 U3486 ( .A(n2697), .ZN(n2698) );
  AOI21_X1 U34870 ( .B1(n3640), .B2(n3664), .A(n2698), .ZN(n2701) );
  OAI21_X1 U3488 ( .B1(n3640), .B2(n2700), .A(n2699), .ZN(n2908) );
  OAI22_X1 U34890 ( .A1(n2701), .A2(n4117), .B1(n4088), .B2(n2908), .ZN(n2903)
         );
  AND2_X1 U3490 ( .A1(n2703), .A2(n2702), .ZN(n2827) );
  INV_X1 U34910 ( .A(n2704), .ZN(n2834) );
  NOR2_X1 U3492 ( .A1(n2839), .A2(n2834), .ZN(n2706) );
  NAND4_X1 U34930 ( .A1(n2827), .A2(n2706), .A3(n2705), .A4(n2826), .ZN(n2708)
         );
  MUX2_X1 U3494 ( .A(REG2_REG_1__SCAN_IN), .B(n2903), .S(n4006), .Z(n2716) );
  NAND2_X1 U34950 ( .A1(n4006), .A2(n4161), .ZN(n4097) );
  INV_X1 U3496 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2709) );
  OAI22_X1 U34970 ( .A1(n2821), .A2(n4097), .B1(n2709), .B2(n4476), .ZN(n2715)
         );
  AND2_X1 U3498 ( .A1(n4006), .A2(n4250), .ZN(n4138) );
  INV_X1 U34990 ( .A(n4138), .ZN(n3057) );
  AND2_X1 U3500 ( .A1(n4006), .A2(n4249), .ZN(n4139) );
  INV_X1 U35010 ( .A(n4139), .ZN(n2710) );
  OAI22_X1 U3502 ( .A1(n2939), .A2(n3057), .B1(n2710), .B2(n2904), .ZN(n2714)
         );
  OR2_X1 U35030 ( .A1(n2846), .A2(n3818), .ZN(n3008) );
  INV_X1 U3504 ( .A(n4489), .ZN(n4102) );
  NAND2_X1 U35050 ( .A1(n4006), .A2(n3818), .ZN(n4024) );
  INV_X1 U35060 ( .A(n4021), .ZN(n2711) );
  NAND2_X1 U35070 ( .A1(n2855), .A2(n2822), .ZN(n2712) );
  NAND2_X1 U35080 ( .A1(n2955), .A2(n2712), .ZN(n2911) );
  OAI22_X1 U35090 ( .A1(n2908), .A2(n4102), .B1(n4142), .B2(n2911), .ZN(n2713)
         );
  INV_X2 U35100 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U35110 ( .A(DATAI_4_), .ZN(n2717) );
  INV_X1 U35120 ( .A(n2760), .ZN(n2884) );
  MUX2_X1 U35130 ( .A(n2717), .B(n2884), .S(STATE_REG_SCAN_IN), .Z(n2718) );
  INV_X1 U35140 ( .A(n2718), .ZN(U3348) );
  MUX2_X1 U35150 ( .A(n2374), .B(n3793), .S(STATE_REG_SCAN_IN), .Z(n2719) );
  INV_X1 U35160 ( .A(n2719), .ZN(U3344) );
  INV_X1 U35170 ( .A(DATAI_27_), .ZN(n2721) );
  NAND2_X1 U35180 ( .A1(n2766), .A2(STATE_REG_SCAN_IN), .ZN(n2720) );
  OAI21_X1 U35190 ( .B1(STATE_REG_SCAN_IN), .B2(n2721), .A(n2720), .ZN(U3325)
         );
  INV_X1 U35200 ( .A(DATAI_29_), .ZN(n2723) );
  NAND2_X1 U35210 ( .A1(n2282), .A2(STATE_REG_SCAN_IN), .ZN(n2722) );
  OAI21_X1 U35220 ( .B1(STATE_REG_SCAN_IN), .B2(n2723), .A(n2722), .ZN(U3323)
         );
  INV_X1 U35230 ( .A(DATAI_28_), .ZN(n4692) );
  NAND2_X1 U35240 ( .A1(n2861), .A2(STATE_REG_SCAN_IN), .ZN(n2724) );
  OAI21_X1 U35250 ( .B1(STATE_REG_SCAN_IN), .B2(n4692), .A(n2724), .ZN(U3324)
         );
  INV_X1 U35260 ( .A(DATAI_31_), .ZN(n2728) );
  OR4_X1 U35270 ( .A1(n2726), .A2(IR_REG_30__SCAN_IN), .A3(U3149), .A4(n2725), 
        .ZN(n2727) );
  OAI21_X1 U35280 ( .B1(STATE_REG_SCAN_IN), .B2(n2728), .A(n2727), .ZN(U3321)
         );
  INV_X1 U35290 ( .A(n2729), .ZN(n2730) );
  INV_X1 U35300 ( .A(n2731), .ZN(n2733) );
  AOI22_X1 U35310 ( .A1(n4537), .A2(n2734), .B1(n2733), .B2(n2732), .ZN(U3458)
         );
  NOR2_X1 U35320 ( .A1(n4351), .A2(n4496), .ZN(n2736) );
  AOI22_X1 U35330 ( .A1(n4537), .A2(n2737), .B1(n2736), .B2(n2735), .ZN(U3459)
         );
  NAND2_X1 U35340 ( .A1(n2915), .A2(n2738), .ZN(n2739) );
  INV_X1 U35350 ( .A(n2746), .ZN(n2740) );
  OR2_X1 U35360 ( .A1(n2915), .A2(U3149), .ZN(n3742) );
  NAND2_X1 U35370 ( .A1(n2839), .A2(n3742), .ZN(n2745) );
  NOR2_X1 U35380 ( .A1(n4467), .A2(U4043), .ZN(U3148) );
  INV_X1 U35390 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U35400 ( .A1(n3549), .A2(U4043), .ZN(n2741) );
  OAI21_X1 U35410 ( .B1(U4043), .B2(n4710), .A(n2741), .ZN(U3553) );
  INV_X1 U35420 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4562) );
  NAND2_X1 U35430 ( .A1(n4057), .A2(U4043), .ZN(n2742) );
  OAI21_X1 U35440 ( .B1(U4043), .B2(n4562), .A(n2742), .ZN(U3567) );
  INV_X1 U35450 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4706) );
  NAND2_X1 U35460 ( .A1(n3103), .A2(U4043), .ZN(n2743) );
  OAI21_X1 U35470 ( .B1(U4043), .B2(n4706), .A(n2743), .ZN(U3555) );
  INV_X1 U35480 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4707) );
  NAND2_X1 U35490 ( .A1(n3036), .A2(U4043), .ZN(n2744) );
  OAI21_X1 U35500 ( .B1(U4043), .B2(n4707), .A(n2744), .ZN(U3552) );
  INV_X1 U35510 ( .A(n2802), .ZN(n4359) );
  AND2_X1 U35520 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3762) );
  NAND2_X1 U35530 ( .A1(n4362), .A2(REG1_REG_1__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U35540 ( .A1(n3761), .A2(n2747), .ZN(n2867) );
  INV_X1 U35550 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2956) );
  XNOR2_X1 U35560 ( .A(n2055), .B(n2956), .ZN(n2868) );
  NAND2_X1 U35570 ( .A1(n2867), .A2(n2868), .ZN(n2866) );
  NAND2_X1 U35580 ( .A1(n2055), .A2(REG1_REG_2__SCAN_IN), .ZN(n2748) );
  NAND2_X1 U35590 ( .A1(n2866), .A2(n2748), .ZN(n2749) );
  INV_X1 U35600 ( .A(n4360), .ZN(n2776) );
  XNOR2_X1 U35610 ( .A(n2749), .B(n2776), .ZN(n2779) );
  NAND2_X1 U35620 ( .A1(n2779), .A2(REG1_REG_3__SCAN_IN), .ZN(n2778) );
  NAND2_X1 U35630 ( .A1(n2749), .A2(n4360), .ZN(n2750) );
  NAND2_X1 U35640 ( .A1(n2778), .A2(n2750), .ZN(n2751) );
  XNOR2_X1 U35650 ( .A(n2751), .B(n2884), .ZN(n2881) );
  NAND2_X1 U35660 ( .A1(n2881), .A2(REG1_REG_4__SCAN_IN), .ZN(n2880) );
  XOR2_X1 U35670 ( .A(REG1_REG_5__SCAN_IN), .B(n2802), .Z(n2796) );
  XOR2_X1 U35680 ( .A(n4358), .B(n2752), .Z(n2788) );
  INV_X1 U35690 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3106) );
  NOR2_X1 U35700 ( .A1(n4357), .A2(REG1_REG_7__SCAN_IN), .ZN(n2753) );
  INV_X1 U35710 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4534) );
  INV_X1 U35720 ( .A(n4357), .ZN(n2809) );
  XNOR2_X1 U35730 ( .A(n3795), .B(REG1_REG_8__SCAN_IN), .ZN(n2754) );
  NAND2_X1 U35740 ( .A1(n2754), .A2(n4469), .ZN(n2765) );
  NOR2_X1 U35750 ( .A1(n2843), .A2(n2860), .ZN(n3739) );
  NAND2_X1 U35760 ( .A1(n4362), .A2(REG2_REG_1__SCAN_IN), .ZN(n2871) );
  XNOR2_X1 U35770 ( .A(n2756), .B(n4360), .ZN(n2775) );
  INV_X1 U35780 ( .A(n2756), .ZN(n2757) );
  AOI22_X1 U35790 ( .A1(n2775), .A2(REG2_REG_3__SCAN_IN), .B1(n4360), .B2(
        n2757), .ZN(n2758) );
  XNOR2_X1 U35800 ( .A(n2758), .B(n2760), .ZN(n2879) );
  INV_X1 U35810 ( .A(n2758), .ZN(n2759) );
  AOI22_X1 U3582 ( .A1(n2879), .A2(REG2_REG_4__SCAN_IN), .B1(n2760), .B2(n2759), .ZN(n2800) );
  INV_X1 U3583 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3012) );
  MUX2_X1 U3584 ( .A(REG2_REG_5__SCAN_IN), .B(n3012), .S(n2802), .Z(n2799) );
  INV_X1 U3585 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3074) );
  MUX2_X1 U3586 ( .A(n3074), .B(REG2_REG_7__SCAN_IN), .S(n4357), .Z(n2811) );
  XNOR2_X1 U3587 ( .A(REG2_REG_8__SCAN_IN), .B(n3772), .ZN(n2761) );
  NAND2_X1 U3588 ( .A1(n4411), .A2(n2761), .ZN(n2762) );
  NAND2_X1 U3589 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3142) );
  NAND2_X1 U3590 ( .A1(n2762), .A2(n3142), .ZN(n2763) );
  AOI21_X1 U3591 ( .B1(n4467), .B2(ADDR_REG_8__SCAN_IN), .A(n2763), .ZN(n2764)
         );
  OAI211_X1 U3592 ( .C1(n4475), .C2(n3793), .A(n2765), .B(n2764), .ZN(U3248)
         );
  INV_X1 U3593 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2898) );
  INV_X1 U3594 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2899) );
  NAND2_X1 U3595 ( .A1(n2766), .A2(n2899), .ZN(n2767) );
  NAND2_X1 U3596 ( .A1(n2861), .A2(n2767), .ZN(n2770) );
  INV_X1 U3597 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2823) );
  AOI21_X1 U3598 ( .B1(n2860), .B2(n2823), .A(IR_REG_0__SCAN_IN), .ZN(n2769)
         );
  NAND2_X1 U3599 ( .A1(n2770), .A2(n2140), .ZN(n2863) );
  OAI211_X1 U3600 ( .C1(n2770), .C2(n2769), .A(n2863), .B(n2768), .ZN(n2771)
         );
  OAI21_X1 U3601 ( .B1(STATE_REG_SCAN_IN), .B2(n2898), .A(n2771), .ZN(n2773)
         );
  INV_X1 U3602 ( .A(n4469), .ZN(n2794) );
  NOR3_X1 U3603 ( .A1(n2794), .A2(REG1_REG_0__SCAN_IN), .A3(n2140), .ZN(n2772)
         );
  AOI211_X1 U3604 ( .C1(n4467), .C2(ADDR_REG_0__SCAN_IN), .A(n2773), .B(n2772), 
        .ZN(n2774) );
  INV_X1 U3605 ( .A(n2774), .ZN(U3240) );
  XNOR2_X1 U3606 ( .A(n2775), .B(REG2_REG_3__SCAN_IN), .ZN(n2782) );
  INV_X1 U3607 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U3608 ( .A1(STATE_REG_SCAN_IN), .A2(n4689), .ZN(n2941) );
  NOR2_X1 U3609 ( .A1(n4475), .A2(n2776), .ZN(n2777) );
  AOI211_X1 U3610 ( .C1(n4467), .C2(ADDR_REG_3__SCAN_IN), .A(n2941), .B(n2777), 
        .ZN(n2781) );
  OAI211_X1 U3611 ( .C1(REG1_REG_3__SCAN_IN), .C2(n2779), .A(n4469), .B(n2778), 
        .ZN(n2780) );
  OAI211_X1 U3612 ( .C1(n2782), .C2(n4463), .A(n2781), .B(n2780), .ZN(U3243)
         );
  XNOR2_X1 U3613 ( .A(n2783), .B(REG2_REG_6__SCAN_IN), .ZN(n2792) );
  INV_X1 U3614 ( .A(n4475), .ZN(n3757) );
  INV_X1 U3615 ( .A(n4467), .ZN(n2786) );
  INV_X1 U3616 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n2785) );
  AND2_X1 U3617 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3095) );
  INV_X1 U3618 ( .A(n3095), .ZN(n2784) );
  OAI21_X1 U3619 ( .B1(n2786), .B2(n2785), .A(n2784), .ZN(n2790) );
  AOI211_X1 U3620 ( .C1(n3106), .C2(n2788), .A(n2794), .B(n2787), .ZN(n2789)
         );
  AOI211_X1 U3621 ( .C1(n3757), .C2(n4358), .A(n2790), .B(n2789), .ZN(n2791)
         );
  OAI21_X1 U3622 ( .B1(n2792), .B2(n4463), .A(n2791), .ZN(U3246) );
  INV_X1 U3623 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U3624 ( .A1(n3416), .A2(U4043), .ZN(n2793) );
  OAI21_X1 U3625 ( .B1(U4043), .B2(n4704), .A(n2793), .ZN(U3579) );
  AOI211_X1 U3626 ( .C1(n2797), .C2(n2796), .A(n2795), .B(n2794), .ZN(n2805)
         );
  AOI211_X1 U3627 ( .C1(n2800), .C2(n2799), .A(n2798), .B(n4463), .ZN(n2804)
         );
  AND2_X1 U3628 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3028) );
  AOI21_X1 U3629 ( .B1(n4467), .B2(ADDR_REG_5__SCAN_IN), .A(n3028), .ZN(n2801)
         );
  OAI21_X1 U3630 ( .B1(n2802), .B2(n4475), .A(n2801), .ZN(n2803) );
  OR3_X1 U3631 ( .A1(n2805), .A2(n2804), .A3(n2803), .ZN(U3245) );
  MUX2_X1 U3632 ( .A(REG1_REG_7__SCAN_IN), .B(n4534), .S(n4357), .Z(n2806) );
  XNOR2_X1 U3633 ( .A(n2807), .B(n2806), .ZN(n2815) );
  AND2_X1 U3634 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3125) );
  AOI21_X1 U3635 ( .B1(n4467), .B2(ADDR_REG_7__SCAN_IN), .A(n3125), .ZN(n2808)
         );
  OAI21_X1 U3636 ( .B1(n2809), .B2(n4475), .A(n2808), .ZN(n2814) );
  AOI211_X1 U3637 ( .C1(n2812), .C2(n2811), .A(n4463), .B(n2810), .ZN(n2813)
         );
  AOI211_X1 U3638 ( .C1(n4469), .C2(n2815), .A(n2814), .B(n2813), .ZN(n2816)
         );
  INV_X1 U3639 ( .A(n2816), .ZN(U3247) );
  INV_X1 U3641 ( .A(n2846), .ZN(n2817) );
  INV_X1 U3642 ( .A(n2931), .ZN(n2836) );
  INV_X1 U3643 ( .A(n2931), .ZN(n3294) );
  OAI21_X1 U3644 ( .B1(n2916), .B2(n2823), .A(n2850), .ZN(n2824) );
  OAI21_X1 U3645 ( .B1(n2825), .B2(n2824), .A(n2851), .ZN(n2862) );
  NAND3_X1 U3646 ( .A1(n2828), .A2(n2827), .A3(n2826), .ZN(n2842) );
  NAND2_X1 U3647 ( .A1(n2889), .A2(n4356), .ZN(n2830) );
  NAND2_X1 U3648 ( .A1(n2830), .A2(n2829), .ZN(n2831) );
  OR2_X1 U3649 ( .A1(n4249), .A2(n2831), .ZN(n2833) );
  OR2_X1 U3650 ( .A1(n2839), .A2(n2833), .ZN(n2832) );
  NAND2_X1 U3651 ( .A1(n2833), .A2(n4113), .ZN(n2835) );
  AOI21_X1 U3652 ( .B1(n2842), .B2(n2835), .A(n2834), .ZN(n2917) );
  INV_X1 U3653 ( .A(n2841), .ZN(n3738) );
  NAND2_X1 U3654 ( .A1(n2842), .A2(n3738), .ZN(n2918) );
  NAND3_X1 U3655 ( .A1(n2917), .A2(n2838), .A3(n2918), .ZN(n3552) );
  NOR3_X1 U3656 ( .A1(n2842), .A2(n4113), .A3(n2839), .ZN(n2840) );
  NOR2_X2 U3657 ( .A1(n2840), .A2(n4486), .ZN(n3570) );
  NOR2_X1 U3658 ( .A1(n2842), .A2(n2841), .ZN(n2856) );
  OAI22_X1 U3659 ( .A1(n3570), .A2(n2891), .B1(n2298), .B2(n3584), .ZN(n2844)
         );
  AOI21_X1 U3660 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3552), .A(n2844), .ZN(n2845)
         );
  OAI21_X1 U3661 ( .B1(n2862), .B2(n3576), .A(n2845), .ZN(U3229) );
  XNOR2_X1 U3662 ( .A(n2848), .B(n3394), .ZN(n2921) );
  INV_X1 U3663 ( .A(n2920), .ZN(n2849) );
  XNOR2_X1 U3664 ( .A(n2921), .B(n2849), .ZN(n2854) );
  OAI21_X1 U3665 ( .B1(n2854), .B2(n2853), .A(n3582), .ZN(n2859) );
  AOI22_X1 U3666 ( .A1(n3587), .A2(n2855), .B1(n3550), .B2(n3036), .ZN(n2858)
         );
  AOI22_X1 U3667 ( .A1(n3553), .A2(n3756), .B1(n3552), .B2(REG3_REG_1__SCAN_IN), .ZN(n2857) );
  OAI211_X1 U3668 ( .C1(n2859), .C2(n2923), .A(n2858), .B(n2857), .ZN(U3219)
         );
  NAND3_X1 U3669 ( .A1(n2862), .A2(n2861), .A3(n2860), .ZN(n2865) );
  AND2_X1 U3670 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3760)
         );
  AOI21_X1 U3671 ( .B1(n3739), .B2(n3760), .A(n3755), .ZN(n2864) );
  NAND3_X1 U3672 ( .A1(n2865), .A2(n2864), .A3(n2863), .ZN(n2888) );
  NAND2_X1 U3673 ( .A1(n3757), .A2(n2055), .ZN(n2877) );
  AOI22_X1 U3674 ( .A1(n4467), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2876) );
  OAI211_X1 U3675 ( .C1(n2868), .C2(n2867), .A(n4469), .B(n2866), .ZN(n2875)
         );
  INV_X1 U3676 ( .A(n2869), .ZN(n2873) );
  NAND3_X1 U3677 ( .A1(n3758), .A2(n2871), .A3(n2870), .ZN(n2872) );
  NAND3_X1 U3678 ( .A1(n4411), .A2(n2873), .A3(n2872), .ZN(n2874) );
  AND4_X1 U3679 ( .A1(n2877), .A2(n2876), .A3(n2875), .A4(n2874), .ZN(n2878)
         );
  NAND2_X1 U3680 ( .A1(n2888), .A2(n2878), .ZN(U3242) );
  XOR2_X1 U3681 ( .A(REG2_REG_4__SCAN_IN), .B(n2879), .Z(n2886) );
  OAI211_X1 U3682 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2881), .A(n4469), .B(n2880), 
        .ZN(n2883) );
  AND2_X1 U3683 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n2976) );
  AOI21_X1 U3684 ( .B1(n4467), .B2(ADDR_REG_4__SCAN_IN), .A(n2976), .ZN(n2882)
         );
  OAI211_X1 U3685 ( .C1(n4475), .C2(n2884), .A(n2883), .B(n2882), .ZN(n2885)
         );
  AOI21_X1 U3686 ( .B1(n4411), .B2(n2886), .A(n2885), .ZN(n2887) );
  NAND2_X1 U3687 ( .A1(n2888), .A2(n2887), .ZN(U3244) );
  NAND2_X1 U3688 ( .A1(n3756), .A2(n2891), .ZN(n3666) );
  NAND2_X1 U3689 ( .A1(n3664), .A2(n3666), .ZN(n3658) );
  INV_X1 U3690 ( .A(n2889), .ZN(n2890) );
  NOR2_X1 U3691 ( .A1(n2891), .A2(n2890), .ZN(n2897) );
  INV_X1 U3692 ( .A(n4088), .ZN(n3040) );
  OAI21_X1 U3693 ( .B1(n3040), .B2(n4145), .A(n3658), .ZN(n2892) );
  OAI21_X1 U3694 ( .B1(n2298), .B2(n4163), .A(n2892), .ZN(n2895) );
  AOI211_X1 U3695 ( .C1(n4520), .C2(n3658), .A(n2897), .B(n2895), .ZN(n4516)
         );
  NAND2_X1 U3696 ( .A1(n4533), .A2(REG1_REG_0__SCAN_IN), .ZN(n2893) );
  OAI21_X1 U3697 ( .B1(n4516), .B2(n4533), .A(n2893), .ZN(U3518) );
  INV_X1 U3698 ( .A(n2894), .ZN(n2896) );
  AOI21_X1 U3699 ( .B1(n2897), .B2(n2896), .A(n2895), .ZN(n2902) );
  OAI22_X1 U3700 ( .A1(n4006), .A2(n2899), .B1(n2898), .B2(n4476), .ZN(n2900)
         );
  AOI21_X1 U3701 ( .B1(n3658), .B2(n4489), .A(n2900), .ZN(n2901) );
  OAI21_X1 U3702 ( .B1(n2902), .B2(n4494), .A(n2901), .ZN(U3290) );
  INV_X1 U3703 ( .A(n2903), .ZN(n2907) );
  OAI22_X1 U3704 ( .A1(n2939), .A2(n4163), .B1(n4113), .B2(n2904), .ZN(n2905)
         );
  AOI21_X1 U3705 ( .B1(n4161), .B2(n3756), .A(n2905), .ZN(n2906) );
  OAI211_X1 U3706 ( .C1(n4263), .C2(n2908), .A(n2907), .B(n2906), .ZN(n2913)
         );
  NAND2_X1 U3707 ( .A1(n2913), .A2(n4536), .ZN(n2910) );
  NAND2_X1 U3708 ( .A1(n4533), .A2(REG1_REG_1__SCAN_IN), .ZN(n2909) );
  OAI211_X1 U3709 ( .C1(n2911), .C2(n4272), .A(n2910), .B(n2909), .ZN(U3519)
         );
  INV_X1 U3710 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4664) );
  OAI22_X1 U3711 ( .A1(n4348), .A2(n2911), .B1(n4530), .B2(n4664), .ZN(n2912)
         );
  AOI21_X1 U3712 ( .B1(n2913), .B2(n4530), .A(n2912), .ZN(n2914) );
  INV_X1 U3713 ( .A(n2914), .ZN(U3469) );
  AND3_X1 U3714 ( .A1(n2917), .A2(n2916), .A3(n2915), .ZN(n2919) );
  OAI22_X1 U3715 ( .A1(n2939), .A2(n3358), .B1(n2931), .B2(n2924), .ZN(n2927)
         );
  OAI22_X1 U3716 ( .A1(n2939), .A2(n2931), .B1(n2057), .B2(n2924), .ZN(n2925)
         );
  XNOR2_X1 U3717 ( .A(n2925), .B(n3394), .ZN(n2926) );
  XOR2_X1 U3718 ( .A(n2927), .B(n2926), .Z(n3547) );
  INV_X1 U3719 ( .A(n2926), .ZN(n2929) );
  INV_X1 U3720 ( .A(n2927), .ZN(n2928) );
  NAND2_X1 U3721 ( .A1(n2929), .A2(n2928), .ZN(n2930) );
  NAND2_X1 U3722 ( .A1(n3549), .A2(n2836), .ZN(n2934) );
  NAND2_X1 U3723 ( .A1(n3045), .A2(n2932), .ZN(n2933) );
  NAND2_X1 U3724 ( .A1(n2934), .A2(n2933), .ZN(n2935) );
  XNOR2_X1 U3725 ( .A(n2935), .B(n3394), .ZN(n2966) );
  OAI22_X1 U3726 ( .A1(n2974), .A2(n3358), .B1(n2931), .B2(n2936), .ZN(n2965)
         );
  XNOR2_X1 U3727 ( .A(n2964), .B(n2963), .ZN(n2938) );
  NAND2_X1 U3728 ( .A1(n2938), .A2(n3582), .ZN(n2943) );
  OAI22_X1 U3729 ( .A1(n2939), .A2(n3585), .B1(n3584), .B2(n3065), .ZN(n2940)
         );
  AOI211_X1 U3730 ( .C1(n3045), .C2(n3587), .A(n2941), .B(n2940), .ZN(n2942)
         );
  OAI211_X1 U3731 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3590), .A(n2943), .B(n2942), 
        .ZN(U3215) );
  NAND2_X1 U3732 ( .A1(n2945), .A2(n2950), .ZN(n2946) );
  NAND2_X1 U3733 ( .A1(n2944), .A2(n2946), .ZN(n3001) );
  AOI22_X1 U3734 ( .A1(n3549), .A2(n4250), .B1(n4249), .B2(n3551), .ZN(n2947)
         );
  OAI21_X1 U3735 ( .B1(n2298), .B2(n4261), .A(n2947), .ZN(n2954) );
  OAI21_X1 U3736 ( .B1(n2950), .B2(n2949), .A(n2948), .ZN(n2951) );
  NAND2_X1 U3737 ( .A1(n2951), .A2(n4145), .ZN(n2953) );
  NAND2_X1 U3738 ( .A1(n3001), .A2(n3040), .ZN(n2952) );
  NAND2_X1 U3739 ( .A1(n2953), .A2(n2952), .ZN(n2998) );
  AOI211_X1 U3740 ( .C1(n4520), .C2(n3001), .A(n2954), .B(n2998), .ZN(n2962)
         );
  XNOR2_X1 U3741 ( .A(n2955), .B(n3551), .ZN(n2997) );
  OAI22_X1 U3742 ( .A1(n4272), .A2(n2997), .B1(n4536), .B2(n2956), .ZN(n2957)
         );
  INV_X1 U3743 ( .A(n2957), .ZN(n2958) );
  OAI21_X1 U3744 ( .B1(n2962), .B2(n4533), .A(n2958), .ZN(U3520) );
  NAND2_X1 U3745 ( .A1(n4528), .A2(REG0_REG_2__SCAN_IN), .ZN(n2961) );
  INV_X1 U3746 ( .A(n4348), .ZN(n3235) );
  INV_X1 U3747 ( .A(n2997), .ZN(n2959) );
  NAND2_X1 U3748 ( .A1(n3235), .A2(n2959), .ZN(n2960) );
  OAI211_X1 U3749 ( .C1(n2962), .C2(n4528), .A(n2961), .B(n2960), .ZN(U3471)
         );
  NAND2_X1 U3750 ( .A1(n2964), .A2(n2963), .ZN(n2968) );
  OR2_X1 U3751 ( .A1(n2966), .A2(n2965), .ZN(n2967) );
  OAI22_X1 U3752 ( .A1(n3065), .A2(n2931), .B1(n2057), .B2(n2989), .ZN(n2969)
         );
  XNOR2_X1 U3753 ( .A(n2969), .B(n3394), .ZN(n3020) );
  OAI22_X1 U3754 ( .A1(n3065), .A2(n3358), .B1(n2931), .B2(n2989), .ZN(n3019)
         );
  XNOR2_X1 U3755 ( .A(n3020), .B(n3019), .ZN(n2971) );
  AOI21_X1 U3756 ( .B1(n2970), .B2(n2971), .A(n3576), .ZN(n2973) );
  NAND2_X1 U3757 ( .A1(n2973), .A2(n3022), .ZN(n2978) );
  OAI22_X1 U3758 ( .A1(n3093), .A2(n3584), .B1(n3585), .B2(n2974), .ZN(n2975)
         );
  AOI211_X1 U3759 ( .C1(n2983), .C2(n3587), .A(n2976), .B(n2975), .ZN(n2977)
         );
  OAI211_X1 U3760 ( .C1(n3590), .C2(n2990), .A(n2978), .B(n2977), .ZN(U3227)
         );
  NAND2_X1 U3761 ( .A1(n2980), .A2(n3651), .ZN(n2981) );
  INV_X1 U3762 ( .A(n4521), .ZN(n2994) );
  XOR2_X1 U3763 ( .A(n3651), .B(n2982), .Z(n2987) );
  AOI22_X1 U3764 ( .A1(n3549), .A2(n4161), .B1(n4249), .B2(n2983), .ZN(n2984)
         );
  OAI21_X1 U3765 ( .B1(n3093), .B2(n4163), .A(n2984), .ZN(n2985) );
  AOI21_X1 U3766 ( .B1(n4521), .B2(n3040), .A(n2985), .ZN(n2986) );
  OAI21_X1 U3767 ( .B1(n2987), .B2(n4117), .A(n2986), .ZN(n4518) );
  INV_X1 U3768 ( .A(n2988), .ZN(n3043) );
  OAI211_X1 U3769 ( .C1(n3043), .C2(n2989), .A(n4021), .B(n3010), .ZN(n4517)
         );
  OAI22_X1 U3770 ( .A1(n4517), .A2(n4356), .B1(n4476), .B2(n2990), .ZN(n2991)
         );
  OAI21_X1 U3771 ( .B1(n4518), .B2(n2991), .A(n4006), .ZN(n2993) );
  NAND2_X1 U3772 ( .A1(n4494), .A2(REG2_REG_4__SCAN_IN), .ZN(n2992) );
  OAI211_X1 U3773 ( .C1(n2994), .C2(n4102), .A(n2993), .B(n2992), .ZN(U3286)
         );
  INV_X1 U3774 ( .A(n4097), .ZN(n4136) );
  AOI22_X1 U3775 ( .A1(n2292), .A2(n4136), .B1(REG3_REG_2__SCAN_IN), .B2(n4486), .ZN(n2996) );
  AOI22_X1 U3776 ( .A1(n3551), .A2(n4139), .B1(n4138), .B2(n3549), .ZN(n2995)
         );
  OAI211_X1 U3777 ( .C1(n2997), .C2(n4142), .A(n2996), .B(n2995), .ZN(n3000)
         );
  MUX2_X1 U3778 ( .A(n2998), .B(REG2_REG_2__SCAN_IN), .S(n4494), .Z(n2999) );
  AOI211_X1 U3779 ( .C1(n4489), .C2(n3001), .A(n3000), .B(n2999), .ZN(n3002)
         );
  INV_X1 U3780 ( .A(n3002), .ZN(U3288) );
  INV_X1 U3781 ( .A(n3003), .ZN(n3676) );
  NAND2_X1 U3782 ( .A1(n3676), .A2(n3692), .ZN(n3641) );
  XNOR2_X1 U3783 ( .A(n3004), .B(n3641), .ZN(n3005) );
  NAND2_X1 U3784 ( .A1(n3005), .A2(n4145), .ZN(n3064) );
  NAND2_X1 U3785 ( .A1(n2979), .A2(n3006), .ZN(n3007) );
  XOR2_X1 U3786 ( .A(n3641), .B(n3007), .Z(n3067) );
  NAND2_X1 U3787 ( .A1(n4088), .A2(n3008), .ZN(n3009) );
  AND2_X1 U3788 ( .A1(n3010), .A2(n3062), .ZN(n3011) );
  NOR2_X1 U3789 ( .A1(n3052), .A2(n3011), .ZN(n3082) );
  INV_X1 U3790 ( .A(n3082), .ZN(n3016) );
  OAI22_X1 U3791 ( .A1(n4006), .A2(n3012), .B1(n3031), .B2(n4476), .ZN(n3013)
         );
  AOI21_X1 U3792 ( .B1(n3754), .B2(n4136), .A(n3013), .ZN(n3015) );
  AOI22_X1 U3793 ( .A1(n4139), .A2(n3062), .B1(n4138), .B2(n3753), .ZN(n3014)
         );
  OAI211_X1 U3794 ( .C1(n3016), .C2(n4142), .A(n3015), .B(n3014), .ZN(n3017)
         );
  AOI21_X1 U3795 ( .B1(n3067), .B2(n4149), .A(n3017), .ZN(n3018) );
  OAI21_X1 U3796 ( .B1(n4494), .B2(n3064), .A(n3018), .ZN(U3285) );
  NAND2_X1 U3797 ( .A1(n3020), .A2(n3019), .ZN(n3021) );
  OAI22_X1 U3798 ( .A1(n3093), .A2(n3358), .B1(n2931), .B2(n3023), .ZN(n3086)
         );
  OAI22_X1 U3799 ( .A1(n3093), .A2(n2931), .B1(n2058), .B2(n3023), .ZN(n3024)
         );
  XNOR2_X1 U3800 ( .A(n3024), .B(n3394), .ZN(n3087) );
  XOR2_X1 U3801 ( .A(n3086), .B(n3087), .Z(n3025) );
  OAI211_X1 U3803 ( .C1(n3026), .C2(n3025), .A(n3089), .B(n3582), .ZN(n3030)
         );
  OAI22_X1 U3804 ( .A1(n3065), .A2(n3585), .B1(n3584), .B2(n3123), .ZN(n3027)
         );
  AOI211_X1 U3805 ( .C1(n3062), .C2(n3587), .A(n3028), .B(n3027), .ZN(n3029)
         );
  OAI211_X1 U3806 ( .C1(n3590), .C2(n3031), .A(n3030), .B(n3029), .ZN(U3224)
         );
  XOR2_X1 U3807 ( .A(n3032), .B(n3649), .Z(n4490) );
  OAI21_X1 U3808 ( .B1(n3649), .B2(n3034), .A(n3033), .ZN(n3035) );
  NAND2_X1 U3809 ( .A1(n3035), .A2(n4145), .ZN(n3038) );
  AOI22_X1 U3810 ( .A1(n3036), .A2(n4161), .B1(n4249), .B2(n3045), .ZN(n3037)
         );
  OAI211_X1 U3811 ( .C1(n3065), .C2(n4163), .A(n3038), .B(n3037), .ZN(n3039)
         );
  AOI21_X1 U3812 ( .B1(n4490), .B2(n3040), .A(n3039), .ZN(n4493) );
  INV_X1 U3813 ( .A(n4493), .ZN(n3041) );
  AOI21_X1 U3814 ( .B1(n4520), .B2(n4490), .A(n3041), .ZN(n3048) );
  INV_X1 U3815 ( .A(n3042), .ZN(n3044) );
  AOI21_X1 U3816 ( .B1(n3045), .B2(n3044), .A(n3043), .ZN(n4487) );
  AOI22_X1 U3817 ( .A1(n4487), .A2(n3235), .B1(REG0_REG_3__SCAN_IN), .B2(n4528), .ZN(n3046) );
  OAI21_X1 U3818 ( .B1(n3048), .B2(n4528), .A(n3046), .ZN(U3473) );
  INV_X1 U3819 ( .A(n4272), .ZN(n3240) );
  AOI22_X1 U3820 ( .A1(n4487), .A2(n3240), .B1(REG1_REG_3__SCAN_IN), .B2(n4533), .ZN(n3047) );
  OAI21_X1 U3821 ( .B1(n3048), .B2(n4533), .A(n3047), .ZN(U3521) );
  NAND2_X1 U3822 ( .A1(n3679), .A2(n3693), .ZN(n3653) );
  XNOR2_X1 U3823 ( .A(n3049), .B(n3653), .ZN(n3105) );
  XNOR2_X1 U3824 ( .A(n3050), .B(n3653), .ZN(n3051) );
  NOR2_X1 U3825 ( .A1(n3051), .A2(n4117), .ZN(n3101) );
  NAND2_X1 U3826 ( .A1(n3101), .A2(n4006), .ZN(n3061) );
  NOR2_X1 U3827 ( .A1(n3052), .A2(n3100), .ZN(n3053) );
  OR2_X1 U3828 ( .A1(n3073), .A2(n3053), .ZN(n3109) );
  INV_X1 U3829 ( .A(n3109), .ZN(n3059) );
  AOI22_X1 U3830 ( .A1(n3103), .A2(n4136), .B1(n3096), .B2(n4139), .ZN(n3056)
         );
  INV_X1 U3831 ( .A(n3099), .ZN(n3054) );
  AOI22_X1 U3832 ( .A1(n4494), .A2(REG2_REG_6__SCAN_IN), .B1(n3054), .B2(n4486), .ZN(n3055) );
  OAI211_X1 U3833 ( .C1(n3121), .C2(n3057), .A(n3056), .B(n3055), .ZN(n3058)
         );
  AOI21_X1 U3834 ( .B1(n3059), .B2(n4488), .A(n3058), .ZN(n3060) );
  OAI211_X1 U3835 ( .C1(n4063), .C2(n3105), .A(n3061), .B(n3060), .ZN(U3284)
         );
  AOI22_X1 U3836 ( .A1(n3753), .A2(n4250), .B1(n4249), .B2(n3062), .ZN(n3063)
         );
  OAI211_X1 U3837 ( .C1(n3065), .C2(n4261), .A(n3064), .B(n3063), .ZN(n3066)
         );
  AOI21_X1 U3838 ( .B1(n3067), .B2(n4523), .A(n3066), .ZN(n3085) );
  AOI22_X1 U3839 ( .A1(n3082), .A2(n3235), .B1(REG0_REG_5__SCAN_IN), .B2(n4528), .ZN(n3068) );
  OAI21_X1 U3840 ( .B1(n3085), .B2(n4528), .A(n3068), .ZN(U3477) );
  XNOR2_X1 U3841 ( .A(n3069), .B(n3680), .ZN(n3072) );
  AOI22_X1 U3842 ( .A1(n3751), .A2(n4250), .B1(n4249), .B2(n3126), .ZN(n3070)
         );
  OAI21_X1 U3843 ( .B1(n3123), .B2(n4261), .A(n3070), .ZN(n3071) );
  AOI21_X1 U3844 ( .B1(n3072), .B2(n4145), .A(n3071), .ZN(n4527) );
  OAI211_X1 U3845 ( .C1(n3073), .C2(n3120), .A(n4021), .B(n3199), .ZN(n4526)
         );
  INV_X1 U3846 ( .A(n4526), .ZN(n3077) );
  INV_X1 U3847 ( .A(n4024), .ZN(n3076) );
  OAI22_X1 U3848 ( .A1(n4006), .A2(n3074), .B1(n3129), .B2(n4476), .ZN(n3075)
         );
  AOI21_X1 U3849 ( .B1(n3077), .B2(n3076), .A(n3075), .ZN(n3081) );
  NAND2_X1 U3850 ( .A1(n3079), .A2(n3680), .ZN(n4524) );
  NAND3_X1 U3851 ( .A1(n3078), .A2(n4524), .A3(n4149), .ZN(n3080) );
  OAI211_X1 U3852 ( .C1(n4527), .C2(n4494), .A(n3081), .B(n3080), .ZN(U3283)
         );
  NAND2_X1 U3853 ( .A1(n4533), .A2(REG1_REG_5__SCAN_IN), .ZN(n3084) );
  NAND2_X1 U3854 ( .A1(n3082), .A2(n3240), .ZN(n3083) );
  OAI211_X1 U3855 ( .C1(n3085), .C2(n4533), .A(n3084), .B(n3083), .ZN(U3523)
         );
  NAND2_X1 U3856 ( .A1(n3087), .A2(n3086), .ZN(n3088) );
  OAI22_X1 U3858 ( .A1(n3123), .A2(n2931), .B1(n2057), .B2(n3100), .ZN(n3090)
         );
  XNOR2_X1 U3859 ( .A(n3090), .B(n3394), .ZN(n3113) );
  OAI22_X1 U3860 ( .A1(n3123), .A2(n3358), .B1(n2931), .B2(n3100), .ZN(n3114)
         );
  XNOR2_X1 U3861 ( .A(n3113), .B(n3114), .ZN(n3091) );
  XNOR2_X1 U3862 ( .A(n3115), .B(n3091), .ZN(n3092) );
  NAND2_X1 U3863 ( .A1(n3092), .A2(n3582), .ZN(n3098) );
  OAI22_X1 U3864 ( .A1(n3121), .A2(n3584), .B1(n3585), .B2(n3093), .ZN(n3094)
         );
  AOI211_X1 U3865 ( .C1(n3096), .C2(n3587), .A(n3095), .B(n3094), .ZN(n3097)
         );
  OAI211_X1 U3866 ( .C1(n3590), .C2(n3099), .A(n3098), .B(n3097), .ZN(U3236)
         );
  OAI22_X1 U3867 ( .A1(n3121), .A2(n4163), .B1(n4113), .B2(n3100), .ZN(n3102)
         );
  AOI211_X1 U3868 ( .C1(n4161), .C2(n3103), .A(n3102), .B(n3101), .ZN(n3104)
         );
  OAI21_X1 U3869 ( .B1(n4213), .B2(n3105), .A(n3104), .ZN(n3111) );
  OAI22_X1 U3870 ( .A1(n3109), .A2(n4272), .B1(n4536), .B2(n3106), .ZN(n3107)
         );
  AOI21_X1 U3871 ( .B1(n3111), .B2(n4536), .A(n3107), .ZN(n3108) );
  INV_X1 U3872 ( .A(n3108), .ZN(U3524) );
  INV_X1 U3873 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4658) );
  OAI22_X1 U3874 ( .A1(n3109), .A2(n4348), .B1(n4530), .B2(n4658), .ZN(n3110)
         );
  AOI21_X1 U3875 ( .B1(n3111), .B2(n4530), .A(n3110), .ZN(n3112) );
  INV_X1 U3876 ( .A(n3112), .ZN(U3479) );
  INV_X1 U3877 ( .A(n3115), .ZN(n3118) );
  INV_X1 U3878 ( .A(n3114), .ZN(n3117) );
  OAI21_X1 U3879 ( .B1(n3118), .B2(n3117), .A(n3116), .ZN(n3131) );
  OAI22_X1 U3880 ( .A1(n3121), .A2(n2931), .B1(n2058), .B2(n3120), .ZN(n3119)
         );
  XNOR2_X1 U3881 ( .A(n3119), .B(n3407), .ZN(n3132) );
  OAI22_X1 U3882 ( .A1(n3121), .A2(n3358), .B1(n2931), .B2(n3120), .ZN(n3133)
         );
  XNOR2_X1 U3883 ( .A(n3132), .B(n3133), .ZN(n3130) );
  XOR2_X1 U3884 ( .A(n3131), .B(n3130), .Z(n3122) );
  NAND2_X1 U3885 ( .A1(n3122), .A2(n3582), .ZN(n3128) );
  OAI22_X1 U3886 ( .A1(n3123), .A2(n3585), .B1(n3584), .B2(n3194), .ZN(n3124)
         );
  AOI211_X1 U3887 ( .C1(n3126), .C2(n3587), .A(n3125), .B(n3124), .ZN(n3127)
         );
  OAI211_X1 U3888 ( .C1(n3590), .C2(n3129), .A(n3128), .B(n3127), .ZN(U3210)
         );
  NAND2_X1 U3889 ( .A1(n3131), .A2(n3130), .ZN(n3136) );
  INV_X1 U3890 ( .A(n3132), .ZN(n3134) );
  NAND2_X1 U3891 ( .A1(n3134), .A2(n3133), .ZN(n3135) );
  NAND2_X1 U3892 ( .A1(n3136), .A2(n3135), .ZN(n3170) );
  OAI22_X1 U3893 ( .A1(n3194), .A2(n2931), .B1(n2057), .B2(n3201), .ZN(n3137)
         );
  XNOR2_X1 U3894 ( .A(n3137), .B(n3394), .ZN(n3139) );
  OAI22_X1 U3895 ( .A1(n3194), .A2(n3358), .B1(n2931), .B2(n3201), .ZN(n3138)
         );
  OR2_X1 U3896 ( .A1(n3139), .A2(n3138), .ZN(n3189) );
  INV_X1 U3897 ( .A(n3189), .ZN(n3140) );
  AND2_X1 U3898 ( .A1(n3139), .A2(n3138), .ZN(n3188) );
  NOR2_X1 U3899 ( .A1(n3140), .A2(n3188), .ZN(n3141) );
  XNOR2_X1 U3900 ( .A(n3170), .B(n3141), .ZN(n3147) );
  INV_X1 U3901 ( .A(n4477), .ZN(n3145) );
  AOI22_X1 U3902 ( .A1(n3550), .A2(n3750), .B1(n3553), .B2(n3752), .ZN(n3143)
         );
  OAI211_X1 U3903 ( .C1(n3570), .C2(n3201), .A(n3143), .B(n3142), .ZN(n3144)
         );
  AOI21_X1 U3904 ( .B1(n3145), .B2(n3574), .A(n3144), .ZN(n3146) );
  OAI21_X1 U3905 ( .B1(n3147), .B2(n3576), .A(n3146), .ZN(U3218) );
  NAND2_X1 U3906 ( .A1(n3750), .A2(n2836), .ZN(n3149) );
  NAND2_X1 U3907 ( .A1(n3229), .A2(n2932), .ZN(n3148) );
  NAND2_X1 U3908 ( .A1(n3149), .A2(n3148), .ZN(n3150) );
  XNOR2_X1 U3909 ( .A(n3150), .B(n3394), .ZN(n3152) );
  OAI22_X1 U3910 ( .A1(n3246), .A2(n3358), .B1(n2931), .B2(n3151), .ZN(n3153)
         );
  XOR2_X1 U3911 ( .A(n3152), .B(n3153), .Z(n3191) );
  INV_X1 U3912 ( .A(n3191), .ZN(n3156) );
  OR2_X1 U3913 ( .A1(n3188), .A2(n3156), .ZN(n3169) );
  OR2_X1 U3914 ( .A1(n3170), .A2(n3169), .ZN(n3159) );
  INV_X1 U3915 ( .A(n3152), .ZN(n3155) );
  INV_X1 U3916 ( .A(n3153), .ZN(n3154) );
  NAND2_X1 U3917 ( .A1(n3155), .A2(n3154), .ZN(n3158) );
  OR2_X1 U3918 ( .A1(n3156), .A2(n3189), .ZN(n3157) );
  AND2_X1 U3919 ( .A1(n3158), .A2(n3157), .ZN(n3166) );
  NAND2_X1 U3920 ( .A1(n3159), .A2(n3166), .ZN(n3164) );
  NAND2_X1 U3921 ( .A1(n3749), .A2(n2836), .ZN(n3162) );
  NAND2_X1 U3922 ( .A1(n3244), .A2(n2932), .ZN(n3161) );
  NAND2_X1 U3923 ( .A1(n3162), .A2(n3161), .ZN(n3163) );
  XNOR2_X1 U3924 ( .A(n3163), .B(n3394), .ZN(n3217) );
  AOI22_X1 U3925 ( .A1(n3749), .A2(n3404), .B1(n2836), .B2(n3244), .ZN(n3218)
         );
  XOR2_X1 U3926 ( .A(n3217), .B(n3218), .Z(n3165) );
  AOI21_X1 U3927 ( .B1(n3164), .B2(n3165), .A(n3576), .ZN(n3171) );
  INV_X1 U3928 ( .A(n3165), .ZN(n3167) );
  AND2_X1 U3929 ( .A1(n3167), .A2(n3166), .ZN(n3168) );
  NAND2_X1 U3930 ( .A1(n3171), .A2(n3221), .ZN(n3175) );
  NAND2_X1 U3931 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4381) );
  INV_X1 U3932 ( .A(n4381), .ZN(n3173) );
  OAI22_X1 U3933 ( .A1(n3246), .A2(n3585), .B1(n3584), .B2(n4253), .ZN(n3172)
         );
  AOI211_X1 U3934 ( .C1(n3244), .C2(n3587), .A(n3173), .B(n3172), .ZN(n3174)
         );
  OAI211_X1 U3935 ( .C1(n3590), .C2(n3253), .A(n3175), .B(n3174), .ZN(U3214)
         );
  INV_X1 U3936 ( .A(n3690), .ZN(n3694) );
  NAND2_X1 U3937 ( .A1(n3694), .A2(n3684), .ZN(n3654) );
  INV_X1 U3938 ( .A(n3654), .ZN(n3177) );
  XNOR2_X1 U3939 ( .A(n3176), .B(n3177), .ZN(n3228) );
  AND2_X1 U3940 ( .A1(n3200), .A2(n3229), .ZN(n3178) );
  NOR2_X1 U3941 ( .A1(n3252), .A2(n3178), .ZN(n3239) );
  NAND2_X1 U3942 ( .A1(n3239), .A2(n4488), .ZN(n3182) );
  OAI22_X1 U3943 ( .A1(n3198), .A2(n4476), .B1(n3770), .B2(n4006), .ZN(n3179)
         );
  AOI21_X1 U3944 ( .B1(n3751), .B2(n4136), .A(n3179), .ZN(n3181) );
  AOI22_X1 U3945 ( .A1(n4139), .A2(n3229), .B1(n4138), .B2(n3749), .ZN(n3180)
         );
  NAND3_X1 U3946 ( .A1(n3182), .A2(n3181), .A3(n3180), .ZN(n3186) );
  XNOR2_X1 U3947 ( .A(n3183), .B(n3654), .ZN(n3184) );
  NAND2_X1 U3948 ( .A1(n3184), .A2(n4145), .ZN(n3231) );
  NOR2_X1 U3949 ( .A1(n3231), .A2(n4494), .ZN(n3185) );
  AOI211_X1 U3950 ( .C1(n3228), .C2(n4149), .A(n3186), .B(n3185), .ZN(n3187)
         );
  INV_X1 U3951 ( .A(n3187), .ZN(U3281) );
  OR2_X1 U3952 ( .A1(n3170), .A2(n3188), .ZN(n3190) );
  NAND2_X1 U3953 ( .A1(n3190), .A2(n3189), .ZN(n3192) );
  XNOR2_X1 U3954 ( .A(n3192), .B(n3191), .ZN(n3193) );
  NAND2_X1 U3955 ( .A1(n3193), .A2(n3582), .ZN(n3197) );
  AND2_X1 U3956 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4377) );
  OAI22_X1 U3957 ( .A1(n3194), .A2(n3585), .B1(n3584), .B2(n4262), .ZN(n3195)
         );
  AOI211_X1 U3958 ( .C1(n3229), .C2(n3587), .A(n4377), .B(n3195), .ZN(n3196)
         );
  OAI211_X1 U3959 ( .C1(n3590), .C2(n3198), .A(n3197), .B(n3196), .ZN(U3228)
         );
  INV_X1 U3960 ( .A(n3199), .ZN(n3202) );
  OAI21_X1 U3961 ( .B1(n3202), .B2(n3201), .A(n3200), .ZN(n4480) );
  INV_X1 U3962 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U3963 ( .A1(n3685), .A2(n3682), .ZN(n3652) );
  XNOR2_X1 U3964 ( .A(n3203), .B(n3652), .ZN(n3207) );
  INV_X1 U3965 ( .A(n3207), .ZN(n4482) );
  XNOR2_X1 U3966 ( .A(n3204), .B(n3652), .ZN(n3210) );
  AOI22_X1 U3967 ( .A1(n3752), .A2(n4161), .B1(n4249), .B2(n3205), .ZN(n3206)
         );
  OAI21_X1 U3968 ( .B1(n3246), .B2(n4163), .A(n3206), .ZN(n3209) );
  NOR2_X1 U3969 ( .A1(n3207), .A2(n4088), .ZN(n3208) );
  AOI211_X1 U3970 ( .C1(n4145), .C2(n3210), .A(n3209), .B(n3208), .ZN(n4485)
         );
  INV_X1 U3971 ( .A(n4485), .ZN(n3211) );
  AOI21_X1 U3972 ( .B1(n4520), .B2(n4482), .A(n3211), .ZN(n3214) );
  MUX2_X1 U3973 ( .A(n3212), .B(n3214), .S(n4536), .Z(n3213) );
  OAI21_X1 U3974 ( .B1(n4480), .B2(n4272), .A(n3213), .ZN(U3526) );
  INV_X1 U3975 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3215) );
  MUX2_X1 U3976 ( .A(n3215), .B(n3214), .S(n4530), .Z(n3216) );
  OAI21_X1 U3977 ( .B1(n4480), .B2(n4348), .A(n3216), .ZN(U3483) );
  INV_X1 U3978 ( .A(n3217), .ZN(n3219) );
  OR2_X1 U3979 ( .A1(n3219), .A2(n3218), .ZN(n3220) );
  NAND2_X1 U3980 ( .A1(n3221), .A2(n3220), .ZN(n3284) );
  OAI22_X1 U3981 ( .A1(n4253), .A2(n2931), .B1(n2058), .B2(n3267), .ZN(n3222)
         );
  XNOR2_X1 U3982 ( .A(n3222), .B(n3394), .ZN(n3282) );
  XNOR2_X1 U3983 ( .A(n3282), .B(n3283), .ZN(n3223) );
  XNOR2_X1 U3984 ( .A(n3284), .B(n3223), .ZN(n3224) );
  NAND2_X1 U3985 ( .A1(n3224), .A2(n3582), .ZN(n3227) );
  AND2_X1 U3986 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4398) );
  OAI22_X1 U3987 ( .A1(n4262), .A2(n3585), .B1(n3584), .B2(n3528), .ZN(n3225)
         );
  AOI211_X1 U3988 ( .C1(n3262), .C2(n3587), .A(n4398), .B(n3225), .ZN(n3226)
         );
  OAI211_X1 U3989 ( .C1(n3590), .C2(n3266), .A(n3227), .B(n3226), .ZN(U3233)
         );
  NAND2_X1 U3990 ( .A1(n3228), .A2(n4523), .ZN(n3233) );
  AOI22_X1 U3991 ( .A1(n3749), .A2(n4250), .B1(n4249), .B2(n3229), .ZN(n3232)
         );
  NAND2_X1 U3992 ( .A1(n3751), .A2(n4161), .ZN(n3230) );
  NAND4_X1 U3993 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n3237)
         );
  MUX2_X1 U3994 ( .A(REG0_REG_9__SCAN_IN), .B(n3237), .S(n4530), .Z(n3234) );
  AOI21_X1 U3995 ( .B1(n3239), .B2(n3235), .A(n3234), .ZN(n3236) );
  INV_X1 U3996 ( .A(n3236), .ZN(U3485) );
  MUX2_X1 U3997 ( .A(REG1_REG_9__SCAN_IN), .B(n3237), .S(n4536), .Z(n3238) );
  AOI21_X1 U3998 ( .B1(n3240), .B2(n3239), .A(n3238), .ZN(n3241) );
  INV_X1 U3999 ( .A(n3241), .ZN(U3527) );
  NAND2_X1 U4000 ( .A1(n3699), .A2(n3700), .ZN(n3639) );
  XOR2_X1 U4001 ( .A(n3639), .B(n3242), .Z(n4268) );
  XOR2_X1 U4002 ( .A(n3243), .B(n3639), .Z(n3248) );
  AOI22_X1 U4003 ( .A1(n4137), .A2(n4250), .B1(n4249), .B2(n3244), .ZN(n3245)
         );
  OAI21_X1 U4004 ( .B1(n3246), .B2(n4261), .A(n3245), .ZN(n3247) );
  AOI21_X1 U4005 ( .B1(n3248), .B2(n4145), .A(n3247), .ZN(n3249) );
  OAI21_X1 U4006 ( .B1(n4268), .B2(n4088), .A(n3249), .ZN(n4269) );
  NAND2_X1 U4007 ( .A1(n4269), .A2(n4006), .ZN(n3258) );
  INV_X1 U4008 ( .A(n3268), .ZN(n3250) );
  OAI21_X1 U4009 ( .B1(n3252), .B2(n3251), .A(n3250), .ZN(n4349) );
  INV_X1 U4010 ( .A(n4349), .ZN(n3256) );
  INV_X1 U4011 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3254) );
  OAI22_X1 U4012 ( .A1(n4006), .A2(n3254), .B1(n3253), .B2(n4476), .ZN(n3255)
         );
  AOI21_X1 U4013 ( .B1(n3256), .B2(n4488), .A(n3255), .ZN(n3257) );
  OAI211_X1 U4014 ( .C1(n4268), .C2(n4102), .A(n3258), .B(n3257), .ZN(U3280)
         );
  INV_X1 U4015 ( .A(n3260), .ZN(n3261) );
  AOI21_X1 U4016 ( .B1(n3650), .B2(n3259), .A(n3261), .ZN(n4264) );
  AOI22_X1 U4017 ( .A1(n4115), .A2(n4250), .B1(n4249), .B2(n3262), .ZN(n3265)
         );
  XNOR2_X1 U4018 ( .A(n4106), .B(n3650), .ZN(n3263) );
  NAND2_X1 U4019 ( .A1(n3263), .A2(n4145), .ZN(n3264) );
  OAI211_X1 U4020 ( .C1(n4264), .C2(n4088), .A(n3265), .B(n3264), .ZN(n4266)
         );
  NAND2_X1 U4021 ( .A1(n4266), .A2(n4006), .ZN(n3272) );
  OAI22_X1 U4022 ( .A1(n4006), .A2(n3769), .B1(n3266), .B2(n4476), .ZN(n3270)
         );
  OAI21_X1 U4023 ( .B1(n3268), .B2(n3267), .A(n4130), .ZN(n4344) );
  NOR2_X1 U4024 ( .A1(n4344), .A2(n4142), .ZN(n3269) );
  AOI211_X1 U4025 ( .C1(n4136), .C2(n3749), .A(n3270), .B(n3269), .ZN(n3271)
         );
  OAI211_X1 U4026 ( .C1(n4264), .C2(n4102), .A(n3272), .B(n3271), .ZN(U3279)
         );
  INV_X1 U4027 ( .A(n3273), .ZN(n3279) );
  INV_X1 U4028 ( .A(n3745), .ZN(n3864) );
  AOI22_X1 U4029 ( .A1(n3416), .A2(n4138), .B1(n4139), .B2(n3409), .ZN(n3275)
         );
  AOI22_X1 U4030 ( .A1(n3426), .A2(n4486), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4494), .ZN(n3274) );
  OAI211_X1 U4031 ( .C1(n3864), .C2(n4097), .A(n3275), .B(n3274), .ZN(n3278)
         );
  NOR2_X1 U4032 ( .A1(n3276), .A2(n4494), .ZN(n3277) );
  AOI211_X1 U4033 ( .C1(n4488), .C2(n3279), .A(n3278), .B(n3277), .ZN(n3280)
         );
  OAI21_X1 U4034 ( .B1(n3281), .B2(n4063), .A(n3280), .ZN(U3262) );
  NAND2_X1 U4035 ( .A1(n4115), .A2(n2836), .ZN(n3286) );
  NAND2_X1 U4036 ( .A1(n4248), .A2(n2932), .ZN(n3285) );
  NAND2_X1 U4037 ( .A1(n3286), .A2(n3285), .ZN(n3287) );
  XNOR2_X1 U4038 ( .A(n3287), .B(n3394), .ZN(n3290) );
  NAND2_X1 U4039 ( .A1(n4115), .A2(n3404), .ZN(n3289) );
  NAND2_X1 U4040 ( .A1(n4248), .A2(n3160), .ZN(n3288) );
  NAND2_X1 U4041 ( .A1(n3289), .A2(n3288), .ZN(n3291) );
  INV_X1 U4042 ( .A(n3290), .ZN(n3293) );
  INV_X1 U40430 ( .A(n3291), .ZN(n3292) );
  NAND2_X1 U4044 ( .A1(n3293), .A2(n3292), .ZN(n3463) );
  AOI22_X1 U4045 ( .A1(n4251), .A2(n3160), .B1(n2932), .B2(n3530), .ZN(n3295)
         );
  XNOR2_X1 U4046 ( .A(n3295), .B(n3394), .ZN(n3524) );
  AOI22_X1 U4047 ( .A1(n4251), .A2(n3404), .B1(n3160), .B2(n3530), .ZN(n3525)
         );
  OAI22_X1 U4048 ( .A1(n4231), .A2(n2931), .B1(n2057), .B2(n4092), .ZN(n3302)
         );
  XNOR2_X1 U4049 ( .A(n3302), .B(n3394), .ZN(n3304) );
  OAI22_X1 U4050 ( .A1(n4231), .A2(n3358), .B1(n2931), .B2(n4092), .ZN(n3303)
         );
  AND2_X1 U4051 ( .A1(n3304), .A2(n3303), .ZN(n3433) );
  OR2_X1 U4052 ( .A1(n3304), .A2(n3303), .ZN(n3432) );
  OAI22_X1 U4053 ( .A1(n4060), .A2(n2931), .B1(n2057), .B2(n4071), .ZN(n3305)
         );
  XNOR2_X1 U4054 ( .A(n3394), .B(n3305), .ZN(n3307) );
  AND2_X1 U4055 ( .A1(n3432), .A2(n3307), .ZN(n3306) );
  OR2_X1 U4056 ( .A1(n3307), .A2(n3432), .ZN(n3483) );
  NAND2_X1 U4057 ( .A1(n4236), .A2(n3404), .ZN(n3309) );
  NAND2_X1 U4058 ( .A1(n4227), .A2(n3160), .ZN(n3308) );
  NAND2_X1 U4059 ( .A1(n3309), .A2(n3308), .ZN(n3580) );
  AND2_X1 U4060 ( .A1(n3483), .A2(n3580), .ZN(n3310) );
  OAI22_X1 U4061 ( .A1(n4219), .A2(n2931), .B1(n2058), .B2(n3488), .ZN(n3311)
         );
  XNOR2_X1 U4062 ( .A(n3311), .B(n3394), .ZN(n3313) );
  OAI22_X1 U4063 ( .A1(n4219), .A2(n3358), .B1(n2931), .B2(n3488), .ZN(n3312)
         );
  NOR2_X1 U4064 ( .A1(n3313), .A2(n3312), .ZN(n3314) );
  AOI21_X1 U4065 ( .B1(n3313), .B2(n3312), .A(n3314), .ZN(n3486) );
  INV_X1 U4066 ( .A(n3314), .ZN(n3315) );
  NAND2_X1 U4067 ( .A1(n3316), .A2(n3315), .ZN(n3495) );
  NAND2_X1 U4068 ( .A1(n4057), .A2(n3160), .ZN(n3318) );
  NAND2_X1 U4069 ( .A1(n4215), .A2(n2932), .ZN(n3317) );
  NAND2_X1 U4070 ( .A1(n3318), .A2(n3317), .ZN(n3319) );
  XNOR2_X1 U4071 ( .A(n3319), .B(n3407), .ZN(n3321) );
  AOI22_X1 U4072 ( .A1(n4057), .A2(n3404), .B1(n3160), .B2(n4215), .ZN(n3320)
         );
  OR2_X1 U4073 ( .A1(n3321), .A2(n3320), .ZN(n3494) );
  NAND2_X1 U4074 ( .A1(n3495), .A2(n3494), .ZN(n3322) );
  NAND2_X1 U4075 ( .A1(n3321), .A2(n3320), .ZN(n3493) );
  AOI22_X1 U4076 ( .A1(n4216), .A2(n3404), .B1(n3160), .B2(n4014), .ZN(n3559)
         );
  OAI22_X1 U4077 ( .A1(n3498), .A2(n2931), .B1(n2057), .B2(n4023), .ZN(n3323)
         );
  XOR2_X1 U4078 ( .A(n3394), .B(n3323), .Z(n3558) );
  OAI22_X1 U4079 ( .A1(n3978), .A2(n2931), .B1(n2058), .B2(n4002), .ZN(n3324)
         );
  XNOR2_X1 U4080 ( .A(n3324), .B(n3394), .ZN(n3326) );
  INV_X1 U4081 ( .A(n3326), .ZN(n3328) );
  OAI22_X1 U4082 ( .A1(n3978), .A2(n3358), .B1(n2931), .B2(n4002), .ZN(n3325)
         );
  INV_X1 U4083 ( .A(n3325), .ZN(n3327) );
  OR2_X1 U4084 ( .A1(n3326), .A2(n3325), .ZN(n3338) );
  OAI21_X1 U4085 ( .B1(n3328), .B2(n3327), .A(n3338), .ZN(n3331) );
  AOI21_X1 U4086 ( .B1(n3332), .B2(n3331), .A(n2073), .ZN(n3337) );
  INV_X1 U4087 ( .A(n4003), .ZN(n3335) );
  AOI22_X1 U4088 ( .A1(n3553), .A2(n4216), .B1(n3550), .B2(n3747), .ZN(n3333)
         );
  NAND2_X1 U4089 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3817) );
  OAI211_X1 U4090 ( .C1(n3570), .C2(n4002), .A(n3333), .B(n3817), .ZN(n3334)
         );
  AOI21_X1 U4091 ( .B1(n3335), .B2(n3574), .A(n3334), .ZN(n3336) );
  OAI21_X1 U4092 ( .B1(n3337), .B2(n3576), .A(n3336), .ZN(U3216) );
  NAND2_X1 U4093 ( .A1(n3747), .A2(n3160), .ZN(n3340) );
  NAND2_X1 U4094 ( .A1(n3983), .A2(n2932), .ZN(n3339) );
  NAND2_X1 U4095 ( .A1(n3340), .A2(n3339), .ZN(n3341) );
  XNOR2_X1 U4096 ( .A(n3341), .B(n3394), .ZN(n3344) );
  NAND2_X1 U4097 ( .A1(n3747), .A2(n3404), .ZN(n3343) );
  NAND2_X1 U4098 ( .A1(n3983), .A2(n3160), .ZN(n3342) );
  NAND2_X1 U4099 ( .A1(n3343), .A2(n3342), .ZN(n3345) );
  NAND2_X1 U4100 ( .A1(n3344), .A2(n3345), .ZN(n3512) );
  NAND2_X1 U4101 ( .A1(n3453), .A2(n3512), .ZN(n3511) );
  INV_X1 U4102 ( .A(n3344), .ZN(n3347) );
  INV_X1 U4103 ( .A(n3345), .ZN(n3346) );
  NAND2_X1 U4104 ( .A1(n3347), .A2(n3346), .ZN(n3514) );
  NAND2_X2 U4105 ( .A1(n3511), .A2(n3514), .ZN(n3457) );
  OAI22_X1 U4106 ( .A1(n3936), .A2(n2931), .B1(n2057), .B2(n3958), .ZN(n3348)
         );
  XNOR2_X1 U4107 ( .A(n3348), .B(n3407), .ZN(n3351) );
  NOR2_X1 U4108 ( .A1(n3958), .A2(n2931), .ZN(n3349) );
  AOI21_X1 U4109 ( .B1(n3976), .B2(n3404), .A(n3349), .ZN(n3352) );
  AND2_X1 U4110 ( .A1(n3351), .A2(n3352), .ZN(n3451) );
  OAI22_X1 U4111 ( .A1(n3458), .A2(n2931), .B1(n2058), .B2(n3939), .ZN(n3350)
         );
  XNOR2_X1 U4112 ( .A(n3350), .B(n3394), .ZN(n3359) );
  OAI22_X1 U4113 ( .A1(n3458), .A2(n3358), .B1(n2931), .B2(n3939), .ZN(n3360)
         );
  XNOR2_X1 U4114 ( .A(n3359), .B(n3360), .ZN(n3538) );
  INV_X1 U4115 ( .A(n3538), .ZN(n3355) );
  INV_X1 U4116 ( .A(n3351), .ZN(n3354) );
  INV_X1 U4117 ( .A(n3352), .ZN(n3353) );
  NAND2_X1 U4118 ( .A1(n3354), .A2(n3353), .ZN(n3533) );
  AND2_X1 U4119 ( .A1(n3355), .A2(n3533), .ZN(n3356) );
  OAI22_X1 U4120 ( .A1(n3899), .A2(n2931), .B1(n2058), .B2(n3923), .ZN(n3357)
         );
  XNOR2_X1 U4121 ( .A(n3357), .B(n3407), .ZN(n3364) );
  OAI22_X1 U4122 ( .A1(n3899), .A2(n3358), .B1(n2931), .B2(n3923), .ZN(n3365)
         );
  XNOR2_X1 U4123 ( .A(n3364), .B(n3365), .ZN(n3442) );
  INV_X1 U4124 ( .A(n3359), .ZN(n3362) );
  INV_X1 U4125 ( .A(n3360), .ZN(n3361) );
  NAND2_X1 U4126 ( .A1(n3362), .A2(n3361), .ZN(n3443) );
  INV_X1 U4127 ( .A(n3364), .ZN(n3366) );
  NAND2_X1 U4128 ( .A1(n3366), .A2(n3365), .ZN(n3371) );
  NOR2_X1 U4129 ( .A1(n3905), .A2(n2931), .ZN(n3367) );
  AOI21_X1 U4130 ( .B1(n3746), .B2(n3404), .A(n3367), .ZN(n3372) );
  OAI22_X1 U4131 ( .A1(n4178), .A2(n2931), .B1(n2057), .B2(n3905), .ZN(n3370)
         );
  XNOR2_X1 U4132 ( .A(n3370), .B(n3394), .ZN(n3505) );
  NAND2_X1 U4133 ( .A1(n3503), .A2(n3505), .ZN(n3375) );
  INV_X1 U4134 ( .A(n3372), .ZN(n3373) );
  NAND2_X1 U4135 ( .A1(n3374), .A2(n3373), .ZN(n3502) );
  NAND2_X1 U4136 ( .A1(n3375), .A2(n3502), .ZN(n3476) );
  NAND2_X1 U4137 ( .A1(n3901), .A2(n3160), .ZN(n3377) );
  NAND2_X1 U4138 ( .A1(n4174), .A2(n2932), .ZN(n3376) );
  NAND2_X1 U4139 ( .A1(n3377), .A2(n3376), .ZN(n3378) );
  XNOR2_X1 U4140 ( .A(n3378), .B(n3407), .ZN(n3382) );
  NOR2_X1 U4141 ( .A1(n3885), .A2(n2931), .ZN(n3380) );
  AOI21_X1 U4142 ( .B1(n3901), .B2(n3404), .A(n3380), .ZN(n3381) );
  NAND2_X1 U4143 ( .A1(n3382), .A2(n3381), .ZN(n3473) );
  NOR2_X1 U4144 ( .A1(n3382), .A2(n3381), .ZN(n3474) );
  NAND2_X1 U4145 ( .A1(n4175), .A2(n3160), .ZN(n3385) );
  NAND2_X1 U4146 ( .A1(n3383), .A2(n2932), .ZN(n3384) );
  NAND2_X1 U4147 ( .A1(n3385), .A2(n3384), .ZN(n3386) );
  XNOR2_X1 U4148 ( .A(n3386), .B(n3407), .ZN(n3391) );
  INV_X1 U4149 ( .A(n3391), .ZN(n3389) );
  NOR2_X1 U4150 ( .A1(n3870), .A2(n2931), .ZN(n3387) );
  AOI21_X1 U4151 ( .B1(n4175), .B2(n3404), .A(n3387), .ZN(n3390) );
  INV_X1 U4152 ( .A(n3390), .ZN(n3388) );
  NAND2_X1 U4153 ( .A1(n3389), .A2(n3388), .ZN(n3566) );
  NAND2_X1 U4154 ( .A1(n3745), .A2(n3160), .ZN(n3393) );
  NAND2_X1 U4155 ( .A1(n4160), .A2(n2932), .ZN(n3392) );
  NAND2_X1 U4156 ( .A1(n3393), .A2(n3392), .ZN(n3395) );
  XNOR2_X1 U4157 ( .A(n3395), .B(n3394), .ZN(n3412) );
  AND2_X1 U4158 ( .A1(n4160), .A2(n3160), .ZN(n3396) );
  AOI21_X1 U4159 ( .B1(n3745), .B2(n3404), .A(n3396), .ZN(n3413) );
  XNOR2_X1 U4160 ( .A(n3412), .B(n3413), .ZN(n3402) );
  INV_X1 U4161 ( .A(n3397), .ZN(n3844) );
  INV_X1 U4162 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3398) );
  OAI22_X1 U4163 ( .A1(n3570), .A2(n3848), .B1(STATE_REG_SCAN_IN), .B2(n3398), 
        .ZN(n3400) );
  OAI22_X1 U4164 ( .A1(n4164), .A2(n3584), .B1(n3847), .B2(n3585), .ZN(n3399)
         );
  AOI211_X1 U4165 ( .C1(n3844), .C2(n3574), .A(n3400), .B(n3399), .ZN(n3401)
         );
  NAND2_X1 U4166 ( .A1(n3403), .A2(n3402), .ZN(n3430) );
  NAND2_X1 U4167 ( .A1(n3843), .A2(n3404), .ZN(n3406) );
  NAND2_X1 U4168 ( .A1(n3409), .A2(n3160), .ZN(n3405) );
  NAND2_X1 U4169 ( .A1(n3406), .A2(n3405), .ZN(n3408) );
  XNOR2_X1 U4170 ( .A(n3408), .B(n3407), .ZN(n3411) );
  AOI22_X1 U4171 ( .A1(n3843), .A2(n3160), .B1(n2932), .B2(n3409), .ZN(n3410)
         );
  XNOR2_X1 U4172 ( .A(n3411), .B(n3410), .ZN(n3420) );
  NAND2_X1 U4173 ( .A1(n3420), .A2(n3582), .ZN(n3429) );
  INV_X1 U4174 ( .A(n3412), .ZN(n3414) );
  NOR2_X1 U4175 ( .A1(n3414), .A2(n3413), .ZN(n3421) );
  NOR3_X1 U4176 ( .A1(n3421), .A2(n3420), .A3(n3576), .ZN(n3415) );
  NAND2_X1 U4177 ( .A1(n3430), .A2(n3415), .ZN(n3428) );
  AOI22_X1 U4178 ( .A1(n3550), .A2(n3416), .B1(n3745), .B2(n3553), .ZN(n3418)
         );
  NAND2_X1 U4179 ( .A1(U3149), .A2(REG3_REG_28__SCAN_IN), .ZN(n3417) );
  OAI211_X1 U4180 ( .C1(n3570), .C2(n3419), .A(n3418), .B(n3417), .ZN(n3425)
         );
  INV_X1 U4181 ( .A(n3420), .ZN(n3423) );
  INV_X1 U4182 ( .A(n3421), .ZN(n3422) );
  NOR3_X1 U4183 ( .A1(n3423), .A2(n3576), .A3(n3422), .ZN(n3424) );
  AOI211_X1 U4184 ( .C1(n3426), .C2(n3574), .A(n3425), .B(n3424), .ZN(n3427)
         );
  OAI211_X1 U4185 ( .C1(n3430), .C2(n3429), .A(n3428), .B(n3427), .ZN(U3217)
         );
  INV_X1 U4186 ( .A(n3432), .ZN(n3434) );
  NOR2_X1 U4187 ( .A1(n3434), .A2(n3433), .ZN(n3435) );
  XNOR2_X1 U4188 ( .A(n3431), .B(n3435), .ZN(n3440) );
  INV_X1 U4189 ( .A(n3436), .ZN(n4094) );
  AOI22_X1 U4190 ( .A1(n3553), .A2(n4251), .B1(n3550), .B2(n4236), .ZN(n3437)
         );
  NAND2_X1 U4191 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4422) );
  OAI211_X1 U4192 ( .C1(n3570), .C2(n4092), .A(n3437), .B(n4422), .ZN(n3438)
         );
  AOI21_X1 U4193 ( .B1(n4094), .B2(n3574), .A(n3438), .ZN(n3439) );
  OAI21_X1 U4194 ( .B1(n3440), .B2(n3576), .A(n3439), .ZN(U3212) );
  NAND2_X1 U4195 ( .A1(n3441), .A2(n3582), .ZN(n3450) );
  AOI21_X1 U4196 ( .B1(n3535), .B2(n3443), .A(n3442), .ZN(n3449) );
  INV_X1 U4197 ( .A(n3924), .ZN(n3447) );
  OAI22_X1 U4198 ( .A1(n4178), .A2(n3584), .B1(n3585), .B2(n3458), .ZN(n3446)
         );
  OAI22_X1 U4199 ( .A1(n3570), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n3444), 
        .ZN(n3445) );
  AOI211_X1 U4200 ( .C1(n3447), .C2(n3574), .A(n3446), .B(n3445), .ZN(n3448)
         );
  OAI21_X1 U4201 ( .B1(n3450), .B2(n3449), .A(n3448), .ZN(U3213) );
  INV_X1 U4202 ( .A(n3451), .ZN(n3452) );
  NAND2_X1 U4203 ( .A1(n3452), .A2(n3533), .ZN(n3456) );
  INV_X1 U4204 ( .A(n3514), .ZN(n3454) );
  OAI211_X1 U4205 ( .C1(n3453), .C2(n3454), .A(n3512), .B(n3456), .ZN(n3455)
         );
  OAI211_X1 U4206 ( .C1(n3457), .C2(n3456), .A(n3582), .B(n3455), .ZN(n3462)
         );
  INV_X1 U4207 ( .A(n3747), .ZN(n4198) );
  OAI22_X1 U4208 ( .A1(n4198), .A2(n3585), .B1(n3584), .B2(n3458), .ZN(n3460)
         );
  NOR2_X1 U4209 ( .A1(n3570), .A2(n3958), .ZN(n3459) );
  AOI211_X1 U4210 ( .C1(REG3_REG_21__SCAN_IN), .C2(U3149), .A(n3460), .B(n3459), .ZN(n3461) );
  OAI211_X1 U4211 ( .C1(n3590), .C2(n3960), .A(n3462), .B(n3461), .ZN(U3220)
         );
  NAND2_X1 U4212 ( .A1(n3464), .A2(n3463), .ZN(n3465) );
  XNOR2_X1 U4213 ( .A(n3466), .B(n3465), .ZN(n3472) );
  INV_X1 U4214 ( .A(n4133), .ZN(n3470) );
  AOI22_X1 U4215 ( .A1(n3553), .A2(n4137), .B1(n3550), .B2(n4251), .ZN(n3467)
         );
  NAND2_X1 U4216 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4402) );
  OAI211_X1 U4217 ( .C1(n3570), .C2(n3468), .A(n3467), .B(n4402), .ZN(n3469)
         );
  AOI21_X1 U4218 ( .B1(n3470), .B2(n3574), .A(n3469), .ZN(n3471) );
  OAI21_X1 U4219 ( .B1(n3472), .B2(n3576), .A(n3471), .ZN(U3221) );
  NOR2_X1 U4220 ( .A1(n3474), .A2(n2217), .ZN(n3475) );
  XNOR2_X1 U4221 ( .A(n3476), .B(n3475), .ZN(n3481) );
  INV_X1 U4222 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3477) );
  OAI22_X1 U4223 ( .A1(n3570), .A2(n3885), .B1(STATE_REG_SCAN_IN), .B2(n3477), 
        .ZN(n3479) );
  OAI22_X1 U4224 ( .A1(n3847), .A2(n3584), .B1(n4178), .B2(n3585), .ZN(n3478)
         );
  AOI211_X1 U4225 ( .C1(n3887), .C2(n3574), .A(n3479), .B(n3478), .ZN(n3480)
         );
  OAI21_X1 U4226 ( .B1(n3481), .B2(n3576), .A(n3480), .ZN(U3222) );
  INV_X1 U4227 ( .A(n3579), .ZN(n3484) );
  AND2_X1 U4228 ( .A1(n3482), .A2(n3483), .ZN(n3578) );
  OAI21_X1 U4229 ( .B1(n3484), .B2(n3580), .A(n3578), .ZN(n3485) );
  XOR2_X1 U4230 ( .A(n3486), .B(n3485), .Z(n3492) );
  INV_X1 U4231 ( .A(n4050), .ZN(n3490) );
  AOI22_X1 U4232 ( .A1(n3553), .A2(n4236), .B1(n3550), .B2(n4057), .ZN(n3487)
         );
  NAND2_X1 U4233 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4442) );
  OAI211_X1 U4234 ( .C1(n3570), .C2(n3488), .A(n3487), .B(n4442), .ZN(n3489)
         );
  AOI21_X1 U4235 ( .B1(n3490), .B2(n3574), .A(n3489), .ZN(n3491) );
  OAI21_X1 U4236 ( .B1(n3492), .B2(n3576), .A(n3491), .ZN(U3223) );
  NAND2_X1 U4237 ( .A1(n3494), .A2(n3493), .ZN(n3496) );
  XOR2_X1 U4238 ( .A(n3496), .B(n3495), .Z(n3497) );
  NAND2_X1 U4239 ( .A1(n3497), .A2(n3582), .ZN(n3501) );
  AND2_X1 U4240 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4457) );
  OAI22_X1 U4241 ( .A1(n3498), .A2(n3584), .B1(n3585), .B2(n4219), .ZN(n3499)
         );
  AOI211_X1 U4242 ( .C1(n4215), .C2(n3587), .A(n4457), .B(n3499), .ZN(n3500)
         );
  OAI211_X1 U4243 ( .C1(n3590), .C2(n4037), .A(n3501), .B(n3500), .ZN(U3225)
         );
  NAND2_X1 U4244 ( .A1(n3502), .A2(n3503), .ZN(n3504) );
  XOR2_X1 U4245 ( .A(n3505), .B(n3504), .Z(n3510) );
  INV_X1 U4246 ( .A(n3907), .ZN(n3508) );
  INV_X1 U4247 ( .A(n3901), .ZN(n3571) );
  OAI22_X1 U4248 ( .A1(n3571), .A2(n3584), .B1(n3585), .B2(n3899), .ZN(n3507)
         );
  OAI22_X1 U4249 ( .A1(n3570), .A2(n3905), .B1(STATE_REG_SCAN_IN), .B2(n4551), 
        .ZN(n3506) );
  AOI211_X1 U4250 ( .C1(n3508), .C2(n3574), .A(n3507), .B(n3506), .ZN(n3509)
         );
  OAI21_X1 U4251 ( .B1(n3510), .B2(n3576), .A(n3509), .ZN(U3226) );
  INV_X1 U4252 ( .A(n3511), .ZN(n3515) );
  AOI21_X1 U4253 ( .B1(n3512), .B2(n3514), .A(n3453), .ZN(n3513) );
  AOI21_X1 U4254 ( .B1(n3515), .B2(n3514), .A(n3513), .ZN(n3522) );
  INV_X1 U4255 ( .A(n3516), .ZN(n3986) );
  OAI22_X1 U4256 ( .A1(n3978), .A2(n3585), .B1(n3584), .B2(n3936), .ZN(n3520)
         );
  OAI22_X1 U4257 ( .A1(n3570), .A2(n3518), .B1(STATE_REG_SCAN_IN), .B2(n3517), 
        .ZN(n3519) );
  AOI211_X1 U4258 ( .C1(n3986), .C2(n3574), .A(n3520), .B(n3519), .ZN(n3521)
         );
  OAI21_X1 U4259 ( .B1(n3522), .B2(n3576), .A(n3521), .ZN(U3230) );
  XOR2_X1 U4260 ( .A(n3525), .B(n3524), .Z(n3526) );
  XNOR2_X1 U4261 ( .A(n3523), .B(n3526), .ZN(n3527) );
  NAND2_X1 U4262 ( .A1(n3527), .A2(n3582), .ZN(n3532) );
  INV_X1 U4263 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4679) );
  NOR2_X1 U4264 ( .A1(STATE_REG_SCAN_IN), .A2(n4679), .ZN(n4415) );
  OAI22_X1 U4265 ( .A1(n3528), .A2(n3585), .B1(n3584), .B2(n4231), .ZN(n3529)
         );
  AOI211_X1 U4266 ( .C1(n3530), .C2(n3587), .A(n4415), .B(n3529), .ZN(n3531)
         );
  OAI211_X1 U4267 ( .C1(n3590), .C2(n4124), .A(n3532), .B(n3531), .ZN(U3231)
         );
  NAND2_X1 U4268 ( .A1(n3534), .A2(n3533), .ZN(n3537) );
  INV_X1 U4269 ( .A(n3535), .ZN(n3536) );
  AOI21_X1 U4270 ( .B1(n3538), .B2(n3537), .A(n3536), .ZN(n3544) );
  INV_X1 U4271 ( .A(n3539), .ZN(n3940) );
  OAI22_X1 U4272 ( .A1(n3899), .A2(n3584), .B1(n3585), .B2(n3936), .ZN(n3542)
         );
  INV_X1 U4273 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3540) );
  OAI22_X1 U4274 ( .A1(n3570), .A2(n3939), .B1(STATE_REG_SCAN_IN), .B2(n3540), 
        .ZN(n3541) );
  AOI211_X1 U4275 ( .C1(n3940), .C2(n3574), .A(n3542), .B(n3541), .ZN(n3543)
         );
  OAI21_X1 U4276 ( .B1(n3544), .B2(n3576), .A(n3543), .ZN(U3232) );
  OAI21_X1 U4277 ( .B1(n3547), .B2(n3546), .A(n3545), .ZN(n3548) );
  NAND2_X1 U4278 ( .A1(n3548), .A2(n3582), .ZN(n3556) );
  AOI22_X1 U4279 ( .A1(n3587), .A2(n3551), .B1(n3550), .B2(n3549), .ZN(n3555)
         );
  AOI22_X1 U4280 ( .A1(n3553), .A2(n2292), .B1(n3552), .B2(REG3_REG_2__SCAN_IN), .ZN(n3554) );
  NAND3_X1 U4281 ( .A1(n3556), .A2(n3555), .A3(n3554), .ZN(U3234) );
  XOR2_X1 U4282 ( .A(n3559), .B(n3558), .Z(n3560) );
  XNOR2_X1 U4283 ( .A(n3557), .B(n3560), .ZN(n3561) );
  NAND2_X1 U4284 ( .A1(n3561), .A2(n3582), .ZN(n3564) );
  AND2_X1 U4285 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4466) );
  OAI22_X1 U4286 ( .A1(n4017), .A2(n3585), .B1(n3584), .B2(n3978), .ZN(n3562)
         );
  AOI211_X1 U4287 ( .C1(n4014), .C2(n3587), .A(n4466), .B(n3562), .ZN(n3563)
         );
  OAI211_X1 U4288 ( .C1(n3590), .C2(n4025), .A(n3564), .B(n3563), .ZN(U3235)
         );
  NAND2_X1 U4289 ( .A1(n2081), .A2(n3566), .ZN(n3567) );
  XNOR2_X1 U4290 ( .A(n3565), .B(n3567), .ZN(n3577) );
  INV_X1 U4291 ( .A(n3568), .ZN(n3872) );
  INV_X1 U4292 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3569) );
  OAI22_X1 U4293 ( .A1(n3570), .A2(n3870), .B1(STATE_REG_SCAN_IN), .B2(n3569), 
        .ZN(n3573) );
  OAI22_X1 U4294 ( .A1(n3864), .A2(n3584), .B1(n3571), .B2(n3585), .ZN(n3572)
         );
  AOI211_X1 U4295 ( .C1(n3872), .C2(n3574), .A(n3573), .B(n3572), .ZN(n3575)
         );
  OAI21_X1 U4296 ( .B1(n3577), .B2(n3576), .A(n3575), .ZN(U3237) );
  NAND2_X1 U4297 ( .A1(n3579), .A2(n3578), .ZN(n3581) );
  XNOR2_X1 U4298 ( .A(n3581), .B(n3580), .ZN(n3583) );
  NAND2_X1 U4299 ( .A1(n3583), .A2(n3582), .ZN(n3589) );
  AND2_X1 U4300 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4436) );
  OAI22_X1 U4301 ( .A1(n4231), .A2(n3585), .B1(n3584), .B2(n4219), .ZN(n3586)
         );
  AOI211_X1 U4302 ( .C1(n4227), .C2(n3587), .A(n4436), .B(n3586), .ZN(n3588)
         );
  OAI211_X1 U4303 ( .C1(n3590), .C2(n4072), .A(n3589), .B(n3588), .ZN(U3238)
         );
  NAND2_X1 U4304 ( .A1(n3591), .A2(DATAI_31_), .ZN(n3825) );
  NAND2_X1 U4305 ( .A1(n4064), .A2(n3594), .ZN(n3706) );
  NAND2_X1 U4306 ( .A1(n3593), .A2(n3592), .ZN(n3689) );
  NAND2_X1 U4307 ( .A1(n3689), .A2(n3594), .ZN(n3705) );
  OAI21_X1 U4308 ( .B1(n4082), .B2(n3706), .A(n3705), .ZN(n3596) );
  AOI211_X1 U4309 ( .C1(n3596), .C2(n3710), .A(n2126), .B(n3712), .ZN(n3597)
         );
  INV_X1 U4310 ( .A(n3597), .ZN(n3600) );
  AOI21_X1 U4311 ( .B1(n3600), .B2(n3599), .A(n3598), .ZN(n3604) );
  INV_X1 U4312 ( .A(n3601), .ZN(n3602) );
  OAI211_X1 U4313 ( .C1(n3602), .C2(n3721), .A(n3657), .B(n3631), .ZN(n3603)
         );
  INV_X1 U4314 ( .A(n3603), .ZN(n3719) );
  OAI21_X1 U4315 ( .B1(n3604), .B2(n3721), .A(n3719), .ZN(n3621) );
  INV_X1 U4316 ( .A(n3744), .ZN(n3610) );
  NAND2_X1 U4317 ( .A1(n2452), .A2(REG1_REG_31__SCAN_IN), .ZN(n3607) );
  NAND2_X1 U4318 ( .A1(n2308), .A2(REG2_REG_31__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4319 ( .A1(n2054), .A2(REG0_REG_31__SCAN_IN), .ZN(n3605) );
  NAND3_X1 U4320 ( .A1(n3607), .A2(n3606), .A3(n3605), .ZN(n3824) );
  AND2_X1 U4321 ( .A1(n3824), .A2(n3825), .ZN(n3728) );
  AOI21_X1 U4322 ( .B1(n3610), .B2(n4157), .A(n3728), .ZN(n3628) );
  NOR2_X1 U4323 ( .A1(n3609), .A2(n3608), .ZN(n3617) );
  AND4_X1 U4324 ( .A1(n3726), .A2(n3628), .A3(n3617), .A4(n3615), .ZN(n3620)
         );
  NOR2_X1 U4325 ( .A1(n3610), .A2(n4157), .ZN(n3625) );
  INV_X1 U4326 ( .A(n3625), .ZN(n3611) );
  AOI21_X1 U4327 ( .B1(n3611), .B2(n3824), .A(n3825), .ZN(n3619) );
  NAND2_X1 U4328 ( .A1(n3613), .A2(n3612), .ZN(n3616) );
  NOR2_X1 U4329 ( .A1(n3614), .A2(n3616), .ZN(n3722) );
  OAI211_X1 U4330 ( .C1(n3617), .C2(n3616), .A(n3628), .B(n3615), .ZN(n3729)
         );
  AOI21_X1 U4331 ( .B1(n3629), .B2(n3722), .A(n3729), .ZN(n3618) );
  AOI211_X1 U4332 ( .C1(n3621), .C2(n3620), .A(n3619), .B(n3618), .ZN(n3622)
         );
  AOI21_X1 U4333 ( .B1(n4157), .B2(n3825), .A(n3622), .ZN(n3736) );
  NAND2_X1 U4334 ( .A1(n3624), .A2(n3623), .ZN(n3858) );
  INV_X1 U4335 ( .A(n3858), .ZN(n3862) );
  INV_X1 U4336 ( .A(n3825), .ZN(n3627) );
  INV_X1 U4337 ( .A(n3824), .ZN(n3626) );
  AOI21_X1 U4338 ( .B1(n3627), .B2(n3626), .A(n3625), .ZN(n3727) );
  NAND4_X1 U4339 ( .A1(n3630), .A2(n3629), .A3(n3727), .A4(n3628), .ZN(n3633)
         );
  NAND2_X1 U4340 ( .A1(n3632), .A2(n3631), .ZN(n3897) );
  NOR4_X1 U4341 ( .A1(n3862), .A2(n4354), .A3(n3633), .A4(n3897), .ZN(n3646)
         );
  INV_X1 U4342 ( .A(n3634), .ZN(n3636) );
  OR2_X1 U4343 ( .A1(n3636), .A2(n3635), .ZN(n3975) );
  INV_X1 U4344 ( .A(n3975), .ZN(n3638) );
  NAND2_X1 U4345 ( .A1(n3637), .A2(n3895), .ZN(n3917) );
  NAND2_X1 U4346 ( .A1(n3970), .A2(n3969), .ZN(n4032) );
  NAND2_X1 U4347 ( .A1(n4111), .A2(n4109), .ZN(n4143) );
  NOR4_X1 U4348 ( .A1(n3638), .A2(n3917), .A3(n4032), .A4(n4143), .ZN(n3644)
         );
  NOR4_X1 U4349 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n3643)
         );
  NAND4_X1 U4350 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .ZN(n3648)
         );
  XNOR2_X1 U4351 ( .A(n3978), .B(n3647), .ZN(n3995) );
  XNOR2_X1 U4352 ( .A(n4251), .B(n4122), .ZN(n4120) );
  NOR3_X1 U4353 ( .A1(n3648), .A2(n3995), .A3(n4120), .ZN(n3663) );
  AND4_X1 U4354 ( .A1(n3651), .A2(n3650), .A3(n4012), .A4(n3649), .ZN(n3662)
         );
  NOR4_X1 U4355 ( .A1(n4085), .A2(n3654), .A3(n3653), .A4(n3652), .ZN(n3661)
         );
  INV_X1 U4356 ( .A(n4068), .ZN(n4065) );
  NAND4_X1 U4357 ( .A1(n3655), .A2(n4065), .A3(n3943), .A4(n3680), .ZN(n3659)
         );
  INV_X1 U4358 ( .A(n3717), .ZN(n3656) );
  INV_X1 U4359 ( .A(n3949), .ZN(n3951) );
  NAND2_X1 U4360 ( .A1(n3860), .A2(n3657), .ZN(n3882) );
  NOR4_X1 U4361 ( .A1(n3659), .A2(n3951), .A3(n3882), .A4(n3658), .ZN(n3660)
         );
  NAND4_X1 U4362 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3733)
         );
  INV_X1 U4363 ( .A(n3664), .ZN(n3667) );
  OAI211_X1 U4364 ( .C1(n3667), .C2(n4354), .A(n3666), .B(n3665), .ZN(n3669)
         );
  NAND3_X1 U4365 ( .A1(n3669), .A2(n3668), .A3(n2589), .ZN(n3672) );
  NAND3_X1 U4366 ( .A1(n3672), .A2(n3671), .A3(n3670), .ZN(n3675) );
  NAND3_X1 U4367 ( .A1(n3675), .A2(n3674), .A3(n3673), .ZN(n3677) );
  NAND4_X1 U4368 ( .A1(n3678), .A2(n3677), .A3(n3693), .A4(n3676), .ZN(n3681)
         );
  NAND3_X1 U4369 ( .A1(n3681), .A2(n3680), .A3(n3679), .ZN(n3688) );
  AND2_X1 U4370 ( .A1(n3683), .A2(n3682), .ZN(n3695) );
  INV_X1 U4371 ( .A(n3684), .ZN(n3687) );
  INV_X1 U4372 ( .A(n3685), .ZN(n3686) );
  AOI211_X1 U4373 ( .C1(n3688), .C2(n3695), .A(n3687), .B(n3686), .ZN(n3691)
         );
  NOR3_X1 U4374 ( .A1(n3691), .A2(n3690), .A3(n3689), .ZN(n3703) );
  INV_X1 U4375 ( .A(n3692), .ZN(n3696) );
  NAND4_X1 U4376 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(n3698)
         );
  INV_X1 U4377 ( .A(n3705), .ZN(n3697) );
  AOI21_X1 U4378 ( .B1(n3699), .B2(n3698), .A(n3697), .ZN(n3702) );
  OAI211_X1 U4379 ( .C1(n3703), .C2(n3702), .A(n3701), .B(n3700), .ZN(n3709)
         );
  INV_X1 U4380 ( .A(n3704), .ZN(n3707) );
  OAI21_X1 U4381 ( .B1(n3707), .B2(n3706), .A(n3705), .ZN(n3708) );
  AND2_X1 U4382 ( .A1(n3709), .A2(n3708), .ZN(n3711) );
  OAI21_X1 U4383 ( .B1(n3711), .B2(n2126), .A(n3710), .ZN(n3715) );
  INV_X1 U4384 ( .A(n3712), .ZN(n3714) );
  INV_X1 U4385 ( .A(n3952), .ZN(n3713) );
  AOI21_X1 U4386 ( .B1(n3715), .B2(n3714), .A(n3713), .ZN(n3718) );
  OAI21_X1 U4387 ( .B1(n3718), .B2(n3717), .A(n3716), .ZN(n3720) );
  OAI21_X1 U4388 ( .B1(n3721), .B2(n3720), .A(n3719), .ZN(n3725) );
  NOR2_X1 U4389 ( .A1(n3864), .A2(n4160), .ZN(n3724) );
  INV_X1 U4390 ( .A(n3722), .ZN(n3723) );
  AOI211_X1 U4391 ( .C1(n3726), .C2(n3725), .A(n3724), .B(n3723), .ZN(n3730)
         );
  OAI22_X1 U4392 ( .A1(n3730), .A2(n3729), .B1(n3728), .B2(n3727), .ZN(n3732)
         );
  MUX2_X1 U4393 ( .A(n3733), .B(n3732), .S(n3731), .Z(n3734) );
  OAI21_X1 U4394 ( .B1(n3736), .B2(n3735), .A(n3734), .ZN(n3737) );
  XNOR2_X1 U4395 ( .A(n3737), .B(n4356), .ZN(n3743) );
  NAND2_X1 U4396 ( .A1(n3739), .A2(n3738), .ZN(n3740) );
  OAI211_X1 U4397 ( .C1(n4353), .C2(n3742), .A(n3740), .B(B_REG_SCAN_IN), .ZN(
        n3741) );
  OAI21_X1 U4398 ( .B1(n3743), .B2(n3742), .A(n3741), .ZN(U3239) );
  MUX2_X1 U4399 ( .A(DATAO_REG_31__SCAN_IN), .B(n3824), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4400 ( .A(DATAO_REG_30__SCAN_IN), .B(n3744), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4401 ( .A(n3843), .B(DATAO_REG_28__SCAN_IN), .S(n3755), .Z(U3578)
         );
  MUX2_X1 U4402 ( .A(DATAO_REG_27__SCAN_IN), .B(n3745), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4403 ( .A(n4175), .B(DATAO_REG_26__SCAN_IN), .S(n3755), .Z(U3576)
         );
  MUX2_X1 U4404 ( .A(DATAO_REG_25__SCAN_IN), .B(n3901), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4405 ( .A(n3746), .B(DATAO_REG_24__SCAN_IN), .S(n3755), .Z(U3574)
         );
  INV_X1 U4406 ( .A(n3899), .ZN(n3933) );
  MUX2_X1 U4407 ( .A(DATAO_REG_23__SCAN_IN), .B(n3933), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4408 ( .A(n4196), .B(DATAO_REG_22__SCAN_IN), .S(n3755), .Z(U3572)
         );
  MUX2_X1 U4409 ( .A(DATAO_REG_21__SCAN_IN), .B(n3976), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4410 ( .A(n3747), .B(DATAO_REG_20__SCAN_IN), .S(n3755), .Z(U3570)
         );
  MUX2_X1 U4411 ( .A(DATAO_REG_19__SCAN_IN), .B(n4015), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4412 ( .A(DATAO_REG_18__SCAN_IN), .B(n4216), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4413 ( .A(DATAO_REG_16__SCAN_IN), .B(n4228), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4414 ( .A(n4236), .B(DATAO_REG_15__SCAN_IN), .S(n3755), .Z(U3565)
         );
  MUX2_X1 U4415 ( .A(DATAO_REG_14__SCAN_IN), .B(n3748), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4416 ( .A(n4251), .B(DATAO_REG_13__SCAN_IN), .S(n3755), .Z(U3563)
         );
  MUX2_X1 U4417 ( .A(n4115), .B(DATAO_REG_12__SCAN_IN), .S(n3755), .Z(U3562)
         );
  MUX2_X1 U4418 ( .A(DATAO_REG_11__SCAN_IN), .B(n4137), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4419 ( .A(n3749), .B(DATAO_REG_10__SCAN_IN), .S(n3755), .Z(U3560)
         );
  MUX2_X1 U4420 ( .A(n3750), .B(DATAO_REG_9__SCAN_IN), .S(n3755), .Z(U3559) );
  MUX2_X1 U4421 ( .A(DATAO_REG_8__SCAN_IN), .B(n3751), .S(U4043), .Z(U3558) );
  MUX2_X1 U4422 ( .A(DATAO_REG_7__SCAN_IN), .B(n3752), .S(U4043), .Z(U3557) );
  MUX2_X1 U4423 ( .A(n3753), .B(DATAO_REG_6__SCAN_IN), .S(n3755), .Z(U3556) );
  MUX2_X1 U4424 ( .A(DATAO_REG_4__SCAN_IN), .B(n3754), .S(U4043), .Z(U3554) );
  MUX2_X1 U4425 ( .A(DATAO_REG_1__SCAN_IN), .B(n2292), .S(U4043), .Z(U3551) );
  MUX2_X1 U4426 ( .A(n3756), .B(DATAO_REG_0__SCAN_IN), .S(n3755), .Z(U3550) );
  NAND2_X1 U4427 ( .A1(n3757), .A2(n4362), .ZN(n3767) );
  OAI211_X1 U4428 ( .C1(n3760), .C2(n3759), .A(n4411), .B(n3758), .ZN(n3766)
         );
  OAI211_X1 U4429 ( .C1(n3763), .C2(n3762), .A(n4469), .B(n3761), .ZN(n3765)
         );
  AOI22_X1 U4430 ( .A1(n4467), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3764) );
  NAND4_X1 U4431 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(U3241)
         );
  INV_X1 U4432 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4675) );
  MUX2_X1 U4433 ( .A(REG2_REG_19__SCAN_IN), .B(n4675), .S(n4356), .Z(n3784) );
  INV_X1 U4434 ( .A(n4498), .ZN(n4474) );
  INV_X1 U4435 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U4436 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4474), .B1(n4498), .B2(
        n4676), .ZN(n4465) );
  NOR2_X1 U4437 ( .A1(n3812), .A2(REG2_REG_17__SCAN_IN), .ZN(n3768) );
  AOI21_X1 U4438 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3812), .A(n3768), .ZN(n4455) );
  INV_X1 U4439 ( .A(n3805), .ZN(n4507) );
  INV_X1 U4440 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4410) );
  INV_X1 U4441 ( .A(n3788), .ZN(n4509) );
  NOR2_X1 U4442 ( .A1(n4410), .A2(n4509), .ZN(n4409) );
  NAND2_X1 U4443 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4511), .ZN(n3776) );
  INV_X1 U4444 ( .A(n4511), .ZN(n4396) );
  INV_X1 U4445 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4446 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4511), .B1(n4396), .B2(
        n3769), .ZN(n4393) );
  NAND2_X1 U4447 ( .A1(n4366), .A2(REG2_REG_9__SCAN_IN), .ZN(n3773) );
  INV_X1 U4448 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3770) );
  MUX2_X1 U4449 ( .A(REG2_REG_9__SCAN_IN), .B(n3770), .S(n4366), .Z(n4371) );
  INV_X1 U4450 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4478) );
  NAND2_X1 U4451 ( .A1(n3797), .A2(n3774), .ZN(n3775) );
  INV_X1 U4452 ( .A(n3797), .ZN(n4513) );
  XNOR2_X1 U4453 ( .A(n3774), .B(n4513), .ZN(n4380) );
  NAND2_X1 U4454 ( .A1(n3801), .A2(n3777), .ZN(n3778) );
  INV_X1 U4455 ( .A(n3801), .ZN(n4510) );
  XNOR2_X1 U4456 ( .A(n3777), .B(n4510), .ZN(n4401) );
  NOR2_X1 U4457 ( .A1(n4507), .A2(n3779), .ZN(n3780) );
  INV_X1 U4458 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4425) );
  NOR2_X1 U4459 ( .A1(n4425), .A2(n4424), .ZN(n4423) );
  NAND2_X1 U4460 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3786), .ZN(n3781) );
  OAI21_X1 U4461 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3786), .A(n3781), .ZN(n4433) );
  INV_X1 U4462 ( .A(n4502), .ZN(n4452) );
  NAND2_X1 U4463 ( .A1(n3782), .A2(n4452), .ZN(n3783) );
  INV_X1 U4464 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4443) );
  NAND2_X1 U4465 ( .A1(n4455), .A2(n4453), .ZN(n4454) );
  INV_X1 U4466 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4647) );
  AOI22_X1 U4467 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4498), .B1(n4474), .B2(
        n4647), .ZN(n4471) );
  NOR2_X1 U4468 ( .A1(n3812), .A2(REG1_REG_17__SCAN_IN), .ZN(n3813) );
  NAND2_X1 U4469 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3786), .ZN(n3808) );
  INV_X1 U4470 ( .A(n3786), .ZN(n4505) );
  INV_X1 U4471 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4472 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3786), .B1(n4505), .B2(
        n3785), .ZN(n4439) );
  NAND2_X1 U4473 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3788), .ZN(n3804) );
  INV_X1 U4474 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4475 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3788), .B1(n4509), .B2(
        n3787), .ZN(n4419) );
  NAND2_X1 U4476 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4511), .ZN(n3800) );
  INV_X1 U4477 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4478 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4511), .B1(n4396), .B2(
        n3789), .ZN(n4390) );
  NAND2_X1 U4479 ( .A1(n4366), .A2(REG1_REG_9__SCAN_IN), .ZN(n3796) );
  INV_X1 U4480 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3790) );
  MUX2_X1 U4481 ( .A(n3790), .B(REG1_REG_9__SCAN_IN), .S(n4366), .Z(n3791) );
  INV_X1 U4482 ( .A(n3791), .ZN(n4368) );
  INV_X1 U4483 ( .A(n3792), .ZN(n3794) );
  OAI22_X1 U4484 ( .A1(n3795), .A2(n3212), .B1(n3794), .B2(n3793), .ZN(n4369)
         );
  NAND2_X1 U4485 ( .A1(n4368), .A2(n4369), .ZN(n4367) );
  NAND2_X1 U4486 ( .A1(n3796), .A2(n4367), .ZN(n3798) );
  NAND2_X1 U4487 ( .A1(n3797), .A2(n3798), .ZN(n3799) );
  XNOR2_X1 U4488 ( .A(n3798), .B(n4513), .ZN(n4385) );
  NAND2_X1 U4489 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4385), .ZN(n4384) );
  NAND2_X1 U4490 ( .A1(n3799), .A2(n4384), .ZN(n4389) );
  NAND2_X1 U4491 ( .A1(n4390), .A2(n4389), .ZN(n4388) );
  NAND2_X1 U4492 ( .A1(n3800), .A2(n4388), .ZN(n3802) );
  NAND2_X1 U4493 ( .A1(n3801), .A2(n3802), .ZN(n3803) );
  XNOR2_X1 U4494 ( .A(n3802), .B(n4510), .ZN(n4406) );
  NAND2_X1 U4495 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4406), .ZN(n4405) );
  NAND2_X1 U4496 ( .A1(n3803), .A2(n4405), .ZN(n4418) );
  NAND2_X1 U4497 ( .A1(n4419), .A2(n4418), .ZN(n4417) );
  NAND2_X1 U4498 ( .A1(n3804), .A2(n4417), .ZN(n3806) );
  NAND2_X1 U4499 ( .A1(n3805), .A2(n3806), .ZN(n3807) );
  XNOR2_X1 U4500 ( .A(n3806), .B(n4507), .ZN(n4429) );
  NAND2_X1 U4501 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4429), .ZN(n4428) );
  NAND2_X1 U4502 ( .A1(n3807), .A2(n4428), .ZN(n4438) );
  NAND2_X1 U4503 ( .A1(n4439), .A2(n4438), .ZN(n4437) );
  NOR2_X1 U4504 ( .A1(n4502), .A2(n3809), .ZN(n3810) );
  INV_X1 U4505 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3811) );
  INV_X1 U4506 ( .A(n3812), .ZN(n4501) );
  AOI22_X1 U4507 ( .A1(n3812), .A2(n3811), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4501), .ZN(n4458) );
  NOR2_X1 U4508 ( .A1(n4459), .A2(n4458), .ZN(n4460) );
  INV_X1 U4509 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3814) );
  MUX2_X1 U4510 ( .A(n3814), .B(REG1_REG_19__SCAN_IN), .S(n4356), .Z(n3815) );
  NAND2_X1 U4511 ( .A1(n4467), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3816) );
  OAI211_X1 U4512 ( .C1(n4475), .C2(n3818), .A(n3817), .B(n3816), .ZN(n3819)
         );
  AOI21_X1 U4513 ( .B1(n3820), .B2(n4469), .A(n3819), .ZN(n3821) );
  OAI21_X1 U4514 ( .B1(n3822), .B2(n4463), .A(n3821), .ZN(U3259) );
  XNOR2_X1 U4515 ( .A(n4153), .B(n3825), .ZN(n4276) );
  NAND2_X1 U4516 ( .A1(n3824), .A2(n3823), .ZN(n4155) );
  OAI21_X1 U4517 ( .B1(n3825), .B2(n4113), .A(n4155), .ZN(n4273) );
  NAND2_X1 U4518 ( .A1(n4273), .A2(n4006), .ZN(n3827) );
  NAND2_X1 U4519 ( .A1(n4494), .A2(REG2_REG_31__SCAN_IN), .ZN(n3826) );
  OAI211_X1 U4520 ( .C1(n4276), .C2(n4142), .A(n3827), .B(n3826), .ZN(U3260)
         );
  INV_X1 U4521 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U4522 ( .A1(n3828), .A2(n4149), .ZN(n3833) );
  OAI22_X1 U4523 ( .A1(n3830), .A2(n4142), .B1(n4476), .B2(n3829), .ZN(n3831)
         );
  OAI21_X1 U4524 ( .B1(n2071), .B2(n3831), .A(n4006), .ZN(n3832) );
  OAI211_X1 U4525 ( .C1(n4006), .C2(n3834), .A(n3833), .B(n3832), .ZN(U3354)
         );
  NAND2_X1 U4526 ( .A1(n3894), .A2(n3835), .ZN(n3837) );
  NAND2_X1 U4527 ( .A1(n3837), .A2(n3836), .ZN(n3838) );
  XNOR2_X1 U4528 ( .A(n3838), .B(n3839), .ZN(n4167) );
  INV_X1 U4529 ( .A(n4167), .ZN(n3854) );
  NAND2_X1 U4530 ( .A1(n3840), .A2(n3839), .ZN(n3841) );
  AOI21_X1 U4531 ( .B1(n3842), .B2(n3841), .A(n4117), .ZN(n4166) );
  AOI22_X1 U4532 ( .A1(n3843), .A2(n4138), .B1(n4160), .B2(n4139), .ZN(n3846)
         );
  AOI22_X1 U4533 ( .A1(n3844), .A2(n4486), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4494), .ZN(n3845) );
  OAI211_X1 U4534 ( .C1(n3847), .C2(n4097), .A(n3846), .B(n3845), .ZN(n3852)
         );
  NOR2_X1 U4535 ( .A1(n3868), .A2(n3848), .ZN(n3849) );
  NOR2_X1 U4536 ( .A1(n4283), .A2(n4142), .ZN(n3851) );
  AOI211_X1 U4537 ( .C1(n4166), .C2(n4006), .A(n3852), .B(n3851), .ZN(n3853)
         );
  OAI21_X1 U4538 ( .B1(n3854), .B2(n4063), .A(n3853), .ZN(U3263) );
  NAND2_X1 U4539 ( .A1(n3894), .A2(n3855), .ZN(n3857) );
  INV_X1 U4540 ( .A(n4171), .ZN(n3876) );
  NAND2_X1 U4541 ( .A1(n3861), .A2(n3860), .ZN(n3863) );
  XNOR2_X1 U4542 ( .A(n3863), .B(n3862), .ZN(n3867) );
  OAI22_X1 U4543 ( .A1(n3864), .A2(n4163), .B1(n4113), .B2(n3870), .ZN(n3865)
         );
  AOI21_X1 U4544 ( .B1(n4161), .B2(n3901), .A(n3865), .ZN(n3866) );
  OAI21_X1 U4545 ( .B1(n3867), .B2(n4117), .A(n3866), .ZN(n4170) );
  INV_X1 U4546 ( .A(n3884), .ZN(n3871) );
  INV_X1 U4547 ( .A(n3868), .ZN(n3869) );
  OAI21_X1 U4548 ( .B1(n3871), .B2(n3870), .A(n3869), .ZN(n4287) );
  AOI22_X1 U4549 ( .A1(n3872), .A2(n4486), .B1(n4494), .B2(
        REG2_REG_26__SCAN_IN), .ZN(n3873) );
  OAI21_X1 U4550 ( .B1(n4287), .B2(n4142), .A(n3873), .ZN(n3874) );
  AOI21_X1 U4551 ( .B1(n4170), .B2(n4006), .A(n3874), .ZN(n3875) );
  OAI21_X1 U4552 ( .B1(n3876), .B2(n4063), .A(n3875), .ZN(U3264) );
  XNOR2_X1 U4553 ( .A(n3877), .B(n3882), .ZN(n3878) );
  NAND2_X1 U4554 ( .A1(n3878), .A2(n4145), .ZN(n4177) );
  NAND2_X1 U4555 ( .A1(n3894), .A2(n3879), .ZN(n3881) );
  NAND2_X1 U4556 ( .A1(n3881), .A2(n3880), .ZN(n3883) );
  XNOR2_X1 U4557 ( .A(n3883), .B(n3882), .ZN(n4180) );
  NAND2_X1 U4558 ( .A1(n4180), .A2(n4149), .ZN(n3893) );
  INV_X1 U4559 ( .A(n3904), .ZN(n3886) );
  OAI21_X1 U4560 ( .B1(n3886), .B2(n3885), .A(n3884), .ZN(n4291) );
  INV_X1 U4561 ( .A(n4291), .ZN(n3891) );
  AOI22_X1 U4562 ( .A1(n4175), .A2(n4138), .B1(n4139), .B2(n4174), .ZN(n3889)
         );
  AOI22_X1 U4563 ( .A1(n4494), .A2(REG2_REG_25__SCAN_IN), .B1(n3887), .B2(
        n4486), .ZN(n3888) );
  OAI211_X1 U4564 ( .C1(n4178), .C2(n4097), .A(n3889), .B(n3888), .ZN(n3890)
         );
  AOI21_X1 U4565 ( .B1(n3891), .B2(n4488), .A(n3890), .ZN(n3892) );
  OAI211_X1 U4566 ( .C1(n4494), .C2(n4177), .A(n3893), .B(n3892), .ZN(U3265)
         );
  XNOR2_X1 U4567 ( .A(n3894), .B(n3897), .ZN(n4184) );
  INV_X1 U4568 ( .A(n4184), .ZN(n3912) );
  NAND2_X1 U4569 ( .A1(n3896), .A2(n3895), .ZN(n3898) );
  XNOR2_X1 U4570 ( .A(n3898), .B(n3897), .ZN(n3903) );
  OAI22_X1 U4571 ( .A1(n3899), .A2(n4261), .B1(n4113), .B2(n3905), .ZN(n3900)
         );
  AOI21_X1 U4572 ( .B1(n4250), .B2(n3901), .A(n3900), .ZN(n3902) );
  OAI21_X1 U4573 ( .B1(n3903), .B2(n4117), .A(n3902), .ZN(n4183) );
  INV_X1 U4574 ( .A(n3922), .ZN(n3906) );
  OAI21_X1 U4575 ( .B1(n3906), .B2(n3905), .A(n3904), .ZN(n4295) );
  NOR2_X1 U4576 ( .A1(n4295), .A2(n4142), .ZN(n3910) );
  INV_X1 U4577 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3908) );
  OAI22_X1 U4578 ( .A1(n4006), .A2(n3908), .B1(n3907), .B2(n4476), .ZN(n3909)
         );
  AOI211_X1 U4579 ( .C1(n4183), .C2(n4006), .A(n3910), .B(n3909), .ZN(n3911)
         );
  OAI21_X1 U4580 ( .B1(n3912), .B2(n4063), .A(n3911), .ZN(U3266) );
  XOR2_X1 U4581 ( .A(n3917), .B(n3913), .Z(n4188) );
  INV_X1 U4582 ( .A(n4188), .ZN(n3929) );
  NAND2_X1 U4583 ( .A1(n3953), .A2(n3952), .ZN(n3914) );
  NAND2_X1 U4584 ( .A1(n3914), .A2(n3949), .ZN(n3955) );
  NAND2_X1 U4585 ( .A1(n3955), .A2(n3915), .ZN(n3931) );
  NAND2_X1 U4586 ( .A1(n3931), .A2(n3943), .ZN(n3930) );
  NAND2_X1 U4587 ( .A1(n3930), .A2(n3916), .ZN(n3918) );
  XNOR2_X1 U4588 ( .A(n3918), .B(n3917), .ZN(n3921) );
  OAI22_X1 U4589 ( .A1(n4178), .A2(n4163), .B1(n4113), .B2(n3923), .ZN(n3919)
         );
  AOI21_X1 U4590 ( .B1(n4161), .B2(n4196), .A(n3919), .ZN(n3920) );
  OAI21_X1 U4591 ( .B1(n3921), .B2(n4117), .A(n3920), .ZN(n4187) );
  OAI21_X1 U4592 ( .B1(n3937), .B2(n3923), .A(n3922), .ZN(n4299) );
  NOR2_X1 U4593 ( .A1(n4299), .A2(n4142), .ZN(n3927) );
  INV_X1 U4594 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3925) );
  OAI22_X1 U4595 ( .A1(n4006), .A2(n3925), .B1(n3924), .B2(n4476), .ZN(n3926)
         );
  AOI211_X1 U4596 ( .C1(n4187), .C2(n4006), .A(n3927), .B(n3926), .ZN(n3928)
         );
  OAI21_X1 U4597 ( .B1(n3929), .B2(n4063), .A(n3928), .ZN(U3267) );
  OAI21_X1 U4598 ( .B1(n3943), .B2(n3931), .A(n3930), .ZN(n3932) );
  NAND2_X1 U4599 ( .A1(n3932), .A2(n4145), .ZN(n3935) );
  AOI22_X1 U4600 ( .A1(n3933), .A2(n4250), .B1(n4249), .B2(n2519), .ZN(n3934)
         );
  OAI211_X1 U4601 ( .C1(n3936), .C2(n4261), .A(n3935), .B(n3934), .ZN(n4192)
         );
  INV_X1 U4602 ( .A(n3937), .ZN(n3938) );
  OAI21_X1 U4603 ( .B1(n3956), .B2(n3939), .A(n3938), .ZN(n4303) );
  AOI22_X1 U4604 ( .A1(n4494), .A2(REG2_REG_22__SCAN_IN), .B1(n3940), .B2(
        n4486), .ZN(n3941) );
  OAI21_X1 U4605 ( .B1(n4303), .B2(n4142), .A(n3941), .ZN(n3947) );
  INV_X1 U4606 ( .A(n3942), .ZN(n3945) );
  AND2_X1 U4607 ( .A1(n3944), .A2(n3943), .ZN(n4191) );
  NOR3_X1 U4608 ( .A1(n3945), .A2(n4191), .A3(n4063), .ZN(n3946) );
  AOI211_X1 U4609 ( .C1(n4006), .C2(n4192), .A(n3947), .B(n3946), .ZN(n3948)
         );
  INV_X1 U4610 ( .A(n3948), .ZN(U3268) );
  XNOR2_X1 U4611 ( .A(n3950), .B(n3949), .ZN(n4201) );
  INV_X1 U4612 ( .A(n4201), .ZN(n3967) );
  NAND3_X1 U4613 ( .A1(n3953), .A2(n3952), .A3(n3951), .ZN(n3954) );
  AOI21_X1 U4614 ( .B1(n3955), .B2(n3954), .A(n4117), .ZN(n4200) );
  INV_X1 U4615 ( .A(n3985), .ZN(n3959) );
  INV_X1 U4616 ( .A(n3956), .ZN(n3957) );
  OAI21_X1 U4617 ( .B1(n3959), .B2(n3958), .A(n3957), .ZN(n4307) );
  NOR2_X1 U4618 ( .A1(n4307), .A2(n4142), .ZN(n3965) );
  AOI22_X1 U4619 ( .A1(n4139), .A2(n4195), .B1(n4138), .B2(n4196), .ZN(n3963)
         );
  INV_X1 U4620 ( .A(n3960), .ZN(n3961) );
  AOI22_X1 U4621 ( .A1(n4494), .A2(REG2_REG_21__SCAN_IN), .B1(n3961), .B2(
        n4486), .ZN(n3962) );
  OAI211_X1 U4622 ( .C1(n4198), .C2(n4097), .A(n3963), .B(n3962), .ZN(n3964)
         );
  AOI211_X1 U4623 ( .C1(n4200), .C2(n4006), .A(n3965), .B(n3964), .ZN(n3966)
         );
  OAI21_X1 U4624 ( .B1(n3967), .B2(n4063), .A(n3966), .ZN(U3269) );
  XNOR2_X1 U4625 ( .A(n3968), .B(n3975), .ZN(n3982) );
  INV_X1 U4626 ( .A(n3969), .ZN(n3971) );
  OAI21_X1 U4627 ( .B1(n4030), .B2(n3971), .A(n3970), .ZN(n4013) );
  AOI21_X1 U4628 ( .B1(n4013), .B2(n3973), .A(n3972), .ZN(n3974) );
  XOR2_X1 U4629 ( .A(n3975), .B(n3974), .Z(n3980) );
  AOI22_X1 U4630 ( .A1(n3976), .A2(n4250), .B1(n4249), .B2(n3983), .ZN(n3977)
         );
  OAI21_X1 U4631 ( .B1(n3978), .B2(n4261), .A(n3977), .ZN(n3979) );
  AOI21_X1 U4632 ( .B1(n3980), .B2(n4145), .A(n3979), .ZN(n3981) );
  OAI21_X1 U4633 ( .B1(n3982), .B2(n4088), .A(n3981), .ZN(n4204) );
  INV_X1 U4634 ( .A(n4204), .ZN(n3990) );
  INV_X1 U4635 ( .A(n3982), .ZN(n4205) );
  NAND2_X1 U4636 ( .A1(n4001), .A2(n3983), .ZN(n3984) );
  NAND2_X1 U4637 ( .A1(n3985), .A2(n3984), .ZN(n4311) );
  AOI22_X1 U4638 ( .A1(n4494), .A2(REG2_REG_20__SCAN_IN), .B1(n3986), .B2(
        n4486), .ZN(n3987) );
  OAI21_X1 U4639 ( .B1(n4311), .B2(n4142), .A(n3987), .ZN(n3988) );
  AOI21_X1 U4640 ( .B1(n4205), .B2(n4489), .A(n3988), .ZN(n3989) );
  OAI21_X1 U4641 ( .B1(n3990), .B2(n4494), .A(n3989), .ZN(U3270) );
  XNOR2_X1 U4642 ( .A(n3991), .B(n3995), .ZN(n4209) );
  INV_X1 U4643 ( .A(n4209), .ZN(n4008) );
  INV_X1 U4644 ( .A(n3992), .ZN(n3994) );
  OAI21_X1 U4645 ( .B1(n4013), .B2(n3994), .A(n3993), .ZN(n3997) );
  INV_X1 U4646 ( .A(n3995), .ZN(n3996) );
  XNOR2_X1 U4647 ( .A(n3997), .B(n3996), .ZN(n4000) );
  OAI22_X1 U4648 ( .A1(n4198), .A2(n4163), .B1(n4113), .B2(n4002), .ZN(n3998)
         );
  AOI21_X1 U4649 ( .B1(n4161), .B2(n4216), .A(n3998), .ZN(n3999) );
  OAI21_X1 U4650 ( .B1(n4000), .B2(n4117), .A(n3999), .ZN(n4208) );
  OAI21_X1 U4651 ( .B1(n4020), .B2(n4002), .A(n4001), .ZN(n4315) );
  NOR2_X1 U4652 ( .A1(n4315), .A2(n4142), .ZN(n4005) );
  OAI22_X1 U4653 ( .A1(n4006), .A2(n4675), .B1(n4003), .B2(n4476), .ZN(n4004)
         );
  AOI211_X1 U4654 ( .C1(n4208), .C2(n4006), .A(n4005), .B(n4004), .ZN(n4007)
         );
  OAI21_X1 U4655 ( .B1(n4008), .B2(n4063), .A(n4007), .ZN(U3271) );
  INV_X1 U4656 ( .A(n4009), .ZN(n4010) );
  AOI21_X1 U4657 ( .B1(n4012), .B2(n4011), .A(n4010), .ZN(n4214) );
  XNOR2_X1 U4658 ( .A(n4013), .B(n4012), .ZN(n4019) );
  AOI22_X1 U4659 ( .A1(n4015), .A2(n4250), .B1(n4249), .B2(n4014), .ZN(n4016)
         );
  OAI21_X1 U4660 ( .B1(n4017), .B2(n4261), .A(n4016), .ZN(n4018) );
  AOI21_X1 U4661 ( .B1(n4019), .B2(n4145), .A(n4018), .ZN(n4212) );
  INV_X1 U4662 ( .A(n4212), .ZN(n4028) );
  INV_X1 U4663 ( .A(n4020), .ZN(n4022) );
  OAI211_X1 U4664 ( .C1(n4034), .C2(n4023), .A(n4022), .B(n4021), .ZN(n4211)
         );
  NOR2_X1 U4665 ( .A1(n4211), .A2(n4024), .ZN(n4027) );
  OAI22_X1 U4666 ( .A1(n4006), .A2(n4676), .B1(n4025), .B2(n4476), .ZN(n4026)
         );
  AOI211_X1 U4667 ( .C1(n4028), .C2(n4006), .A(n4027), .B(n4026), .ZN(n4029)
         );
  OAI21_X1 U4668 ( .B1(n4214), .B2(n4063), .A(n4029), .ZN(U3272) );
  XNOR2_X1 U4669 ( .A(n4030), .B(n4032), .ZN(n4031) );
  NAND2_X1 U4670 ( .A1(n4031), .A2(n4145), .ZN(n4218) );
  XNOR2_X1 U4671 ( .A(n4033), .B(n4032), .ZN(n4221) );
  NAND2_X1 U4672 ( .A1(n4221), .A2(n4149), .ZN(n4044) );
  INV_X1 U4673 ( .A(n4034), .ZN(n4035) );
  OAI21_X1 U4674 ( .B1(n2146), .B2(n4036), .A(n4035), .ZN(n4320) );
  INV_X1 U4675 ( .A(n4320), .ZN(n4042) );
  AOI22_X1 U4676 ( .A1(n4216), .A2(n4138), .B1(n4215), .B2(n4139), .ZN(n4040)
         );
  INV_X1 U4677 ( .A(n4037), .ZN(n4038) );
  AOI22_X1 U4678 ( .A1(n4494), .A2(REG2_REG_17__SCAN_IN), .B1(n4038), .B2(
        n4486), .ZN(n4039) );
  OAI211_X1 U4679 ( .C1(n4219), .C2(n4097), .A(n4040), .B(n4039), .ZN(n4041)
         );
  AOI21_X1 U4680 ( .B1(n4042), .B2(n4488), .A(n4041), .ZN(n4043) );
  OAI211_X1 U4681 ( .C1(n4494), .C2(n4218), .A(n4044), .B(n4043), .ZN(U3273)
         );
  NOR2_X1 U4682 ( .A1(n4045), .A2(n4053), .ZN(n4046) );
  OR2_X1 U4683 ( .A1(n4047), .A2(n4046), .ZN(n4223) );
  NAND2_X1 U4684 ( .A1(n4070), .A2(n4056), .ZN(n4048) );
  NAND2_X1 U4685 ( .A1(n4049), .A2(n4048), .ZN(n4324) );
  INV_X1 U4686 ( .A(n4324), .ZN(n4052) );
  OAI22_X1 U4687 ( .A1(n4006), .A2(n4443), .B1(n4050), .B2(n4476), .ZN(n4051)
         );
  AOI21_X1 U4688 ( .B1(n4052), .B2(n4488), .A(n4051), .ZN(n4062) );
  XNOR2_X1 U4689 ( .A(n4054), .B(n4053), .ZN(n4055) );
  NAND2_X1 U4690 ( .A1(n4055), .A2(n4145), .ZN(n4059) );
  AOI22_X1 U4691 ( .A1(n4057), .A2(n4250), .B1(n4249), .B2(n4056), .ZN(n4058)
         );
  OAI211_X1 U4692 ( .C1(n4060), .C2(n4261), .A(n4059), .B(n4058), .ZN(n4224)
         );
  NAND2_X1 U4693 ( .A1(n4224), .A2(n4006), .ZN(n4061) );
  OAI211_X1 U4694 ( .C1(n4223), .C2(n4063), .A(n4062), .B(n4061), .ZN(U3274)
         );
  NAND2_X1 U4695 ( .A1(n4083), .A2(n4064), .ZN(n4066) );
  XNOR2_X1 U4696 ( .A(n4066), .B(n4065), .ZN(n4067) );
  NAND2_X1 U4697 ( .A1(n4067), .A2(n4145), .ZN(n4230) );
  XNOR2_X1 U4698 ( .A(n4069), .B(n4068), .ZN(n4233) );
  NAND2_X1 U4699 ( .A1(n4233), .A2(n4149), .ZN(n4079) );
  OAI21_X1 U4700 ( .B1(n4090), .B2(n4071), .A(n4070), .ZN(n4328) );
  INV_X1 U4701 ( .A(n4328), .ZN(n4077) );
  AOI22_X1 U4702 ( .A1(n4228), .A2(n4138), .B1(n4139), .B2(n4227), .ZN(n4075)
         );
  INV_X1 U4703 ( .A(n4072), .ZN(n4073) );
  AOI22_X1 U4704 ( .A1(n4494), .A2(REG2_REG_15__SCAN_IN), .B1(n4073), .B2(
        n4486), .ZN(n4074) );
  OAI211_X1 U4705 ( .C1(n4231), .C2(n4097), .A(n4075), .B(n4074), .ZN(n4076)
         );
  AOI21_X1 U4706 ( .B1(n4077), .B2(n4488), .A(n4076), .ZN(n4078) );
  OAI211_X1 U4707 ( .C1(n4494), .C2(n4230), .A(n4079), .B(n4078), .ZN(U3275)
         );
  OAI21_X1 U4708 ( .B1(n4081), .B2(n4085), .A(n4080), .ZN(n4241) );
  INV_X1 U4709 ( .A(n4241), .ZN(n4103) );
  INV_X1 U4710 ( .A(n4082), .ZN(n4086) );
  INV_X1 U4711 ( .A(n4083), .ZN(n4084) );
  AOI21_X1 U4712 ( .B1(n4086), .B2(n4085), .A(n4084), .ZN(n4087) );
  OAI22_X1 U4713 ( .A1(n4103), .A2(n4088), .B1(n4117), .B2(n4087), .ZN(n4239)
         );
  NAND2_X1 U4714 ( .A1(n4239), .A2(n4006), .ZN(n4101) );
  INV_X1 U4715 ( .A(n4121), .ZN(n4093) );
  INV_X1 U4716 ( .A(n4090), .ZN(n4091) );
  OAI21_X1 U4717 ( .B1(n4093), .B2(n4092), .A(n4091), .ZN(n4332) );
  INV_X1 U4718 ( .A(n4332), .ZN(n4099) );
  INV_X1 U4719 ( .A(n4251), .ZN(n4238) );
  AOI22_X1 U4720 ( .A1(n4139), .A2(n4235), .B1(n4138), .B2(n4236), .ZN(n4096)
         );
  AOI22_X1 U4721 ( .A1(n4494), .A2(REG2_REG_14__SCAN_IN), .B1(n4094), .B2(
        n4486), .ZN(n4095) );
  OAI211_X1 U4722 ( .C1(n4238), .C2(n4097), .A(n4096), .B(n4095), .ZN(n4098)
         );
  AOI21_X1 U4723 ( .B1(n4099), .B2(n4488), .A(n4098), .ZN(n4100) );
  OAI211_X1 U4724 ( .C1(n4103), .C2(n4102), .A(n4101), .B(n4100), .ZN(U3276)
         );
  INV_X1 U4725 ( .A(n4104), .ZN(n4105) );
  OR2_X1 U4726 ( .A1(n4106), .A2(n4105), .ZN(n4108) );
  NAND2_X1 U4727 ( .A1(n4108), .A2(n4107), .ZN(n4144) );
  INV_X1 U4728 ( .A(n4109), .ZN(n4110) );
  AOI21_X1 U4729 ( .B1(n4144), .B2(n4111), .A(n4110), .ZN(n4112) );
  XNOR2_X1 U4730 ( .A(n4112), .B(n4120), .ZN(n4118) );
  OAI22_X1 U4731 ( .A1(n4231), .A2(n4163), .B1(n4113), .B2(n4122), .ZN(n4114)
         );
  AOI21_X1 U4732 ( .B1(n4161), .B2(n4115), .A(n4114), .ZN(n4116) );
  OAI21_X1 U4733 ( .B1(n4118), .B2(n4117), .A(n4116), .ZN(n4244) );
  INV_X1 U4734 ( .A(n4244), .ZN(n4128) );
  XNOR2_X1 U4735 ( .A(n4119), .B(n4120), .ZN(n4245) );
  INV_X1 U4736 ( .A(n4132), .ZN(n4123) );
  OAI21_X1 U4737 ( .B1(n4123), .B2(n4122), .A(n4121), .ZN(n4336) );
  NOR2_X1 U4738 ( .A1(n4336), .A2(n4142), .ZN(n4126) );
  OAI22_X1 U4739 ( .A1(n4006), .A2(n4410), .B1(n4124), .B2(n4476), .ZN(n4125)
         );
  AOI211_X1 U4740 ( .C1(n4245), .C2(n4149), .A(n4126), .B(n4125), .ZN(n4127)
         );
  OAI21_X1 U4741 ( .B1(n4128), .B2(n4494), .A(n4127), .ZN(U3277) );
  XNOR2_X1 U4742 ( .A(n4129), .B(n4143), .ZN(n4247) );
  NAND2_X1 U4743 ( .A1(n4130), .A2(n4248), .ZN(n4131) );
  NAND2_X1 U4744 ( .A1(n4132), .A2(n4131), .ZN(n4340) );
  INV_X1 U4745 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4134) );
  OAI22_X1 U4746 ( .A1(n4006), .A2(n4134), .B1(n4133), .B2(n4476), .ZN(n4135)
         );
  AOI21_X1 U4747 ( .B1(n4137), .B2(n4136), .A(n4135), .ZN(n4141) );
  AOI22_X1 U4748 ( .A1(n4139), .A2(n4248), .B1(n4138), .B2(n4251), .ZN(n4140)
         );
  OAI211_X1 U4749 ( .C1(n4340), .C2(n4142), .A(n4141), .B(n4140), .ZN(n4148)
         );
  XNOR2_X1 U4750 ( .A(n4144), .B(n4143), .ZN(n4146) );
  NAND2_X1 U4751 ( .A1(n4146), .A2(n4145), .ZN(n4256) );
  NOR2_X1 U4752 ( .A1(n4256), .A2(n4494), .ZN(n4147) );
  AOI211_X1 U4753 ( .C1(n4149), .C2(n4247), .A(n4148), .B(n4147), .ZN(n4150)
         );
  INV_X1 U4754 ( .A(n4150), .ZN(U3278) );
  NAND2_X1 U4755 ( .A1(n4273), .A2(n4536), .ZN(n4152) );
  NAND2_X1 U4756 ( .A1(n4533), .A2(REG1_REG_31__SCAN_IN), .ZN(n4151) );
  OAI211_X1 U4757 ( .C1(n4276), .C2(n4272), .A(n4152), .B(n4151), .ZN(U3549)
         );
  AOI21_X1 U4758 ( .B1(n4157), .B2(n4154), .A(n4153), .ZN(n4363) );
  INV_X1 U4759 ( .A(n4363), .ZN(n4279) );
  INV_X1 U4760 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4158) );
  INV_X1 U4761 ( .A(n4155), .ZN(n4156) );
  AOI21_X1 U4762 ( .B1(n4157), .B2(n4249), .A(n4156), .ZN(n4365) );
  MUX2_X1 U4763 ( .A(n4158), .B(n4365), .S(n4536), .Z(n4159) );
  OAI21_X1 U4764 ( .B1(n4279), .B2(n4272), .A(n4159), .ZN(U3548) );
  INV_X1 U4765 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U4766 ( .A1(n4175), .A2(n4161), .B1(n4249), .B2(n4160), .ZN(n4162)
         );
  OAI21_X1 U4767 ( .B1(n4164), .B2(n4163), .A(n4162), .ZN(n4165) );
  AOI211_X1 U4768 ( .C1(n4167), .C2(n4523), .A(n4166), .B(n4165), .ZN(n4280)
         );
  MUX2_X1 U4769 ( .A(n4168), .B(n4280), .S(n4536), .Z(n4169) );
  OAI21_X1 U4770 ( .B1(n4272), .B2(n4283), .A(n4169), .ZN(U3545) );
  INV_X1 U4771 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4172) );
  AOI21_X1 U4772 ( .B1(n4171), .B2(n4523), .A(n4170), .ZN(n4284) );
  MUX2_X1 U4773 ( .A(n4172), .B(n4284), .S(n4536), .Z(n4173) );
  OAI21_X1 U4774 ( .B1(n4272), .B2(n4287), .A(n4173), .ZN(U3544) );
  INV_X1 U4775 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U4776 ( .A1(n4175), .A2(n4250), .B1(n4249), .B2(n4174), .ZN(n4176)
         );
  OAI211_X1 U4777 ( .C1(n4178), .C2(n4261), .A(n4177), .B(n4176), .ZN(n4179)
         );
  AOI21_X1 U4778 ( .B1(n4180), .B2(n4523), .A(n4179), .ZN(n4288) );
  MUX2_X1 U4779 ( .A(n4181), .B(n4288), .S(n4536), .Z(n4182) );
  OAI21_X1 U4780 ( .B1(n4272), .B2(n4291), .A(n4182), .ZN(U3543) );
  INV_X1 U4781 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4185) );
  AOI21_X1 U4782 ( .B1(n4184), .B2(n4523), .A(n4183), .ZN(n4292) );
  MUX2_X1 U4783 ( .A(n4185), .B(n4292), .S(n4536), .Z(n4186) );
  OAI21_X1 U4784 ( .B1(n4272), .B2(n4295), .A(n4186), .ZN(U3542) );
  INV_X1 U4785 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4189) );
  AOI21_X1 U4786 ( .B1(n4188), .B2(n4523), .A(n4187), .ZN(n4296) );
  MUX2_X1 U4787 ( .A(n4189), .B(n4296), .S(n4536), .Z(n4190) );
  OAI21_X1 U4788 ( .B1(n4272), .B2(n4299), .A(n4190), .ZN(U3541) );
  INV_X1 U4789 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4695) );
  NOR2_X1 U4790 ( .A1(n4191), .A2(n4213), .ZN(n4193) );
  AOI21_X1 U4791 ( .B1(n4193), .B2(n3942), .A(n4192), .ZN(n4300) );
  MUX2_X1 U4792 ( .A(n4695), .B(n4300), .S(n4536), .Z(n4194) );
  OAI21_X1 U4793 ( .B1(n4272), .B2(n4303), .A(n4194), .ZN(U3540) );
  INV_X1 U4794 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U4795 ( .A1(n4196), .A2(n4250), .B1(n4249), .B2(n4195), .ZN(n4197)
         );
  OAI21_X1 U4796 ( .B1(n4198), .B2(n4261), .A(n4197), .ZN(n4199) );
  AOI211_X1 U4797 ( .C1(n4201), .C2(n4523), .A(n4200), .B(n4199), .ZN(n4304)
         );
  MUX2_X1 U4798 ( .A(n4202), .B(n4304), .S(n4536), .Z(n4203) );
  OAI21_X1 U4799 ( .B1(n4272), .B2(n4307), .A(n4203), .ZN(U3539) );
  INV_X1 U4800 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4206) );
  AOI21_X1 U4801 ( .B1(n4520), .B2(n4205), .A(n4204), .ZN(n4308) );
  MUX2_X1 U4802 ( .A(n4206), .B(n4308), .S(n4536), .Z(n4207) );
  OAI21_X1 U4803 ( .B1(n4272), .B2(n4311), .A(n4207), .ZN(U3538) );
  AOI21_X1 U4804 ( .B1(n4209), .B2(n4523), .A(n4208), .ZN(n4312) );
  MUX2_X1 U4805 ( .A(n3814), .B(n4312), .S(n4536), .Z(n4210) );
  OAI21_X1 U4806 ( .B1(n4272), .B2(n4315), .A(n4210), .ZN(U3537) );
  OAI211_X1 U4807 ( .C1(n4214), .C2(n4213), .A(n4212), .B(n4211), .ZN(n4316)
         );
  MUX2_X1 U4808 ( .A(REG1_REG_18__SCAN_IN), .B(n4316), .S(n4536), .Z(U3536) );
  AOI22_X1 U4809 ( .A1(n4216), .A2(n4250), .B1(n4249), .B2(n4215), .ZN(n4217)
         );
  OAI211_X1 U4810 ( .C1(n4219), .C2(n4261), .A(n4218), .B(n4217), .ZN(n4220)
         );
  AOI21_X1 U4811 ( .B1(n4221), .B2(n4523), .A(n4220), .ZN(n4317) );
  MUX2_X1 U4812 ( .A(n3811), .B(n4317), .S(n4536), .Z(n4222) );
  OAI21_X1 U4813 ( .B1(n4272), .B2(n4320), .A(n4222), .ZN(U3535) );
  INV_X1 U4814 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4661) );
  INV_X1 U4815 ( .A(n4223), .ZN(n4225) );
  AOI21_X1 U4816 ( .B1(n4225), .B2(n4523), .A(n4224), .ZN(n4321) );
  MUX2_X1 U4817 ( .A(n4661), .B(n4321), .S(n4536), .Z(n4226) );
  OAI21_X1 U4818 ( .B1(n4272), .B2(n4324), .A(n4226), .ZN(U3534) );
  AOI22_X1 U4819 ( .A1(n4228), .A2(n4250), .B1(n4249), .B2(n4227), .ZN(n4229)
         );
  OAI211_X1 U4820 ( .C1(n4231), .C2(n4261), .A(n4230), .B(n4229), .ZN(n4232)
         );
  AOI21_X1 U4821 ( .B1(n4233), .B2(n4523), .A(n4232), .ZN(n4326) );
  MUX2_X1 U4822 ( .A(n4326), .B(n3785), .S(n4533), .Z(n4234) );
  OAI21_X1 U4823 ( .B1(n4272), .B2(n4328), .A(n4234), .ZN(U3533) );
  INV_X1 U4824 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U4825 ( .A1(n4236), .A2(n4250), .B1(n4249), .B2(n4235), .ZN(n4237)
         );
  OAI21_X1 U4826 ( .B1(n4238), .B2(n4261), .A(n4237), .ZN(n4240) );
  AOI211_X1 U4827 ( .C1(n4520), .C2(n4241), .A(n4240), .B(n4239), .ZN(n4329)
         );
  MUX2_X1 U4828 ( .A(n4242), .B(n4329), .S(n4536), .Z(n4243) );
  OAI21_X1 U4829 ( .B1(n4272), .B2(n4332), .A(n4243), .ZN(U3532) );
  AOI21_X1 U4830 ( .B1(n4523), .B2(n4245), .A(n4244), .ZN(n4333) );
  MUX2_X1 U4831 ( .A(n3787), .B(n4333), .S(n4536), .Z(n4246) );
  OAI21_X1 U4832 ( .B1(n4272), .B2(n4336), .A(n4246), .ZN(U3531) );
  NAND2_X1 U4833 ( .A1(n4247), .A2(n4523), .ZN(n4258) );
  AOI22_X1 U4834 ( .A1(n4251), .A2(n4250), .B1(n4249), .B2(n4248), .ZN(n4252)
         );
  OAI21_X1 U4835 ( .B1(n4253), .B2(n4261), .A(n4252), .ZN(n4254) );
  INV_X1 U4836 ( .A(n4254), .ZN(n4255) );
  AND2_X1 U4837 ( .A1(n4256), .A2(n4255), .ZN(n4257) );
  NAND2_X1 U4838 ( .A1(n4258), .A2(n4257), .ZN(n4337) );
  MUX2_X1 U4839 ( .A(REG1_REG_12__SCAN_IN), .B(n4337), .S(n4536), .Z(n4259) );
  INV_X1 U4840 ( .A(n4259), .ZN(n4260) );
  OAI21_X1 U4841 ( .B1(n4272), .B2(n4340), .A(n4260), .ZN(U3530) );
  OAI22_X1 U4842 ( .A1(n4264), .A2(n4263), .B1(n4262), .B2(n4261), .ZN(n4265)
         );
  NOR2_X1 U4843 ( .A1(n4266), .A2(n4265), .ZN(n4341) );
  MUX2_X1 U4844 ( .A(n3789), .B(n4341), .S(n4536), .Z(n4267) );
  OAI21_X1 U4845 ( .B1(n4272), .B2(n4344), .A(n4267), .ZN(U3529) );
  INV_X1 U4846 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4568) );
  INV_X1 U4847 ( .A(n4268), .ZN(n4270) );
  AOI21_X1 U4848 ( .B1(n4520), .B2(n4270), .A(n4269), .ZN(n4345) );
  MUX2_X1 U4849 ( .A(n4568), .B(n4345), .S(n4536), .Z(n4271) );
  OAI21_X1 U4850 ( .B1(n4349), .B2(n4272), .A(n4271), .ZN(U3528) );
  NAND2_X1 U4851 ( .A1(n4273), .A2(n4530), .ZN(n4275) );
  NAND2_X1 U4852 ( .A1(n4528), .A2(REG0_REG_31__SCAN_IN), .ZN(n4274) );
  OAI211_X1 U4853 ( .C1(n4276), .C2(n4348), .A(n4275), .B(n4274), .ZN(U3517)
         );
  INV_X1 U4854 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4277) );
  MUX2_X1 U4855 ( .A(n4277), .B(n4365), .S(n4530), .Z(n4278) );
  OAI21_X1 U4856 ( .B1(n4279), .B2(n4348), .A(n4278), .ZN(U3516) );
  INV_X1 U4857 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4281) );
  MUX2_X1 U4858 ( .A(n4281), .B(n4280), .S(n4530), .Z(n4282) );
  OAI21_X1 U4859 ( .B1(n4283), .B2(n4348), .A(n4282), .ZN(U3513) );
  INV_X1 U4860 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4285) );
  MUX2_X1 U4861 ( .A(n4285), .B(n4284), .S(n4530), .Z(n4286) );
  OAI21_X1 U4862 ( .B1(n4287), .B2(n4348), .A(n4286), .ZN(U3512) );
  INV_X1 U4863 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4289) );
  MUX2_X1 U4864 ( .A(n4289), .B(n4288), .S(n4530), .Z(n4290) );
  OAI21_X1 U4865 ( .B1(n4291), .B2(n4348), .A(n4290), .ZN(U3511) );
  INV_X1 U4866 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4293) );
  MUX2_X1 U4867 ( .A(n4293), .B(n4292), .S(n4530), .Z(n4294) );
  OAI21_X1 U4868 ( .B1(n4295), .B2(n4348), .A(n4294), .ZN(U3510) );
  INV_X1 U4869 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4297) );
  MUX2_X1 U4870 ( .A(n4297), .B(n4296), .S(n4530), .Z(n4298) );
  OAI21_X1 U4871 ( .B1(n4299), .B2(n4348), .A(n4298), .ZN(U3509) );
  INV_X1 U4872 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4301) );
  MUX2_X1 U4873 ( .A(n4301), .B(n4300), .S(n4530), .Z(n4302) );
  OAI21_X1 U4874 ( .B1(n4303), .B2(n4348), .A(n4302), .ZN(U3508) );
  INV_X1 U4875 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4305) );
  MUX2_X1 U4876 ( .A(n4305), .B(n4304), .S(n4530), .Z(n4306) );
  OAI21_X1 U4877 ( .B1(n4307), .B2(n4348), .A(n4306), .ZN(U3507) );
  INV_X1 U4878 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4309) );
  MUX2_X1 U4879 ( .A(n4309), .B(n4308), .S(n4530), .Z(n4310) );
  OAI21_X1 U4880 ( .B1(n4311), .B2(n4348), .A(n4310), .ZN(U3506) );
  INV_X1 U4881 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4313) );
  MUX2_X1 U4882 ( .A(n4313), .B(n4312), .S(n4530), .Z(n4314) );
  OAI21_X1 U4883 ( .B1(n4315), .B2(n4348), .A(n4314), .ZN(U3505) );
  MUX2_X1 U4884 ( .A(REG0_REG_18__SCAN_IN), .B(n4316), .S(n4530), .Z(U3503) );
  INV_X1 U4885 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4318) );
  MUX2_X1 U4886 ( .A(n4318), .B(n4317), .S(n4530), .Z(n4319) );
  OAI21_X1 U4887 ( .B1(n4320), .B2(n4348), .A(n4319), .ZN(U3501) );
  INV_X1 U4888 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4322) );
  MUX2_X1 U4889 ( .A(n4322), .B(n4321), .S(n4530), .Z(n4323) );
  OAI21_X1 U4890 ( .B1(n4324), .B2(n4348), .A(n4323), .ZN(U3499) );
  INV_X1 U4891 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4325) );
  MUX2_X1 U4892 ( .A(n4326), .B(n4325), .S(n4528), .Z(n4327) );
  OAI21_X1 U4893 ( .B1(n4328), .B2(n4348), .A(n4327), .ZN(U3497) );
  INV_X1 U4894 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4330) );
  MUX2_X1 U4895 ( .A(n4330), .B(n4329), .S(n4530), .Z(n4331) );
  OAI21_X1 U4896 ( .B1(n4332), .B2(n4348), .A(n4331), .ZN(U3495) );
  INV_X1 U4897 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4334) );
  MUX2_X1 U4898 ( .A(n4334), .B(n4333), .S(n4530), .Z(n4335) );
  OAI21_X1 U4899 ( .B1(n4336), .B2(n4348), .A(n4335), .ZN(U3493) );
  MUX2_X1 U4900 ( .A(REG0_REG_12__SCAN_IN), .B(n4337), .S(n4530), .Z(n4338) );
  INV_X1 U4901 ( .A(n4338), .ZN(n4339) );
  OAI21_X1 U4902 ( .B1(n4340), .B2(n4348), .A(n4339), .ZN(U3491) );
  INV_X1 U4903 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4342) );
  MUX2_X1 U4904 ( .A(n4342), .B(n4341), .S(n4530), .Z(n4343) );
  OAI21_X1 U4905 ( .B1(n4344), .B2(n4348), .A(n4343), .ZN(U3489) );
  INV_X1 U4906 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4346) );
  MUX2_X1 U4907 ( .A(n4346), .B(n4345), .S(n4530), .Z(n4347) );
  OAI21_X1 U4908 ( .B1(n4349), .B2(n4348), .A(n4347), .ZN(U3487) );
  MUX2_X1 U4909 ( .A(n4350), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4910 ( .A(DATAI_26_), .B(n2642), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  MUX2_X1 U4911 ( .A(DATAI_25_), .B(n4351), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4912 ( .A(DATAI_24_), .B(n4352), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4913 ( .A(n4353), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4914 ( .A(DATAI_21_), .B(n4354), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U4915 ( .A(DATAI_20_), .B(n4355), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4916 ( .A(n4356), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4917 ( .A(n4366), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U4918 ( .A(n4357), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4919 ( .A(n4358), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4920 ( .A(n4359), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4921 ( .A(n4360), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4922 ( .A(n2055), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4923 ( .A(n4362), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4924 ( .A1(n4363), .A2(n4488), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4494), .ZN(n4364) );
  OAI21_X1 U4925 ( .B1(n4494), .B2(n4365), .A(n4364), .ZN(U3261) );
  INV_X1 U4926 ( .A(n4366), .ZN(n4375) );
  OAI211_X1 U4927 ( .C1(n4369), .C2(n4368), .A(n4469), .B(n4367), .ZN(n4374)
         );
  OAI211_X1 U4928 ( .C1(n4372), .C2(n4371), .A(n4411), .B(n4370), .ZN(n4373)
         );
  OAI211_X1 U4929 ( .C1(n4475), .C2(n4375), .A(n4374), .B(n4373), .ZN(n4376)
         );
  AOI211_X1 U4930 ( .C1(n4467), .C2(ADDR_REG_9__SCAN_IN), .A(n4377), .B(n4376), 
        .ZN(n4378) );
  INV_X1 U4931 ( .A(n4378), .ZN(U3249) );
  OAI211_X1 U4932 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4380), .A(n4411), .B(n4379), .ZN(n4382) );
  NAND2_X1 U4933 ( .A1(n4382), .A2(n4381), .ZN(n4383) );
  AOI21_X1 U4934 ( .B1(n4467), .B2(ADDR_REG_10__SCAN_IN), .A(n4383), .ZN(n4387) );
  OAI211_X1 U4935 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4385), .A(n4469), .B(n4384), .ZN(n4386) );
  OAI211_X1 U4936 ( .C1(n4475), .C2(n4513), .A(n4387), .B(n4386), .ZN(U3250)
         );
  OAI211_X1 U4937 ( .C1(n4390), .C2(n4389), .A(n4469), .B(n4388), .ZN(n4395)
         );
  OAI211_X1 U4938 ( .C1(n4393), .C2(n4392), .A(n4411), .B(n4391), .ZN(n4394)
         );
  OAI211_X1 U4939 ( .C1(n4475), .C2(n4396), .A(n4395), .B(n4394), .ZN(n4397)
         );
  AOI211_X1 U4940 ( .C1(n4467), .C2(ADDR_REG_11__SCAN_IN), .A(n4398), .B(n4397), .ZN(n4399) );
  INV_X1 U4941 ( .A(n4399), .ZN(U3251) );
  OAI211_X1 U4942 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4401), .A(n4411), .B(n4400), .ZN(n4403) );
  NAND2_X1 U4943 ( .A1(n4403), .A2(n4402), .ZN(n4404) );
  AOI21_X1 U4944 ( .B1(n4467), .B2(ADDR_REG_12__SCAN_IN), .A(n4404), .ZN(n4408) );
  OAI211_X1 U4945 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4406), .A(n4469), .B(n4405), .ZN(n4407) );
  OAI211_X1 U4946 ( .C1(n4475), .C2(n4510), .A(n4408), .B(n4407), .ZN(U3252)
         );
  AOI21_X1 U4947 ( .B1(n4410), .B2(n4509), .A(n4409), .ZN(n4414) );
  OAI21_X1 U4948 ( .B1(n4414), .B2(n4413), .A(n4411), .ZN(n4412) );
  AOI21_X1 U4949 ( .B1(n4414), .B2(n4413), .A(n4412), .ZN(n4416) );
  AOI211_X1 U4950 ( .C1(n4467), .C2(ADDR_REG_13__SCAN_IN), .A(n4416), .B(n4415), .ZN(n4421) );
  OAI211_X1 U4951 ( .C1(n4419), .C2(n4418), .A(n4469), .B(n4417), .ZN(n4420)
         );
  OAI211_X1 U4952 ( .C1(n4475), .C2(n4509), .A(n4421), .B(n4420), .ZN(U3253)
         );
  INV_X1 U4953 ( .A(n4422), .ZN(n4427) );
  AOI211_X1 U4954 ( .C1(n4425), .C2(n4424), .A(n4423), .B(n4463), .ZN(n4426)
         );
  AOI211_X1 U4955 ( .C1(n4467), .C2(ADDR_REG_14__SCAN_IN), .A(n4427), .B(n4426), .ZN(n4431) );
  OAI211_X1 U4956 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4429), .A(n4469), .B(n4428), .ZN(n4430) );
  OAI211_X1 U4957 ( .C1(n4475), .C2(n4507), .A(n4431), .B(n4430), .ZN(U3254)
         );
  AOI211_X1 U4958 ( .C1(n4434), .C2(n4433), .A(n4432), .B(n4463), .ZN(n4435)
         );
  AOI211_X1 U4959 ( .C1(n4467), .C2(ADDR_REG_15__SCAN_IN), .A(n4436), .B(n4435), .ZN(n4441) );
  OAI211_X1 U4960 ( .C1(n4439), .C2(n4438), .A(n4469), .B(n4437), .ZN(n4440)
         );
  OAI211_X1 U4961 ( .C1(n4475), .C2(n4505), .A(n4441), .B(n4440), .ZN(U3255)
         );
  INV_X1 U4962 ( .A(n4442), .ZN(n4447) );
  AOI221_X1 U4963 ( .B1(n4445), .B2(n4444), .C1(n4443), .C2(n4444), .A(n4463), 
        .ZN(n4446) );
  AOI211_X1 U4964 ( .C1(n4467), .C2(ADDR_REG_16__SCAN_IN), .A(n4447), .B(n4446), .ZN(n4451) );
  OAI221_X1 U4965 ( .B1(n4449), .B2(REG1_REG_16__SCAN_IN), .C1(n4449), .C2(
        n4448), .A(n4469), .ZN(n4450) );
  OAI211_X1 U4966 ( .C1(n4475), .C2(n4452), .A(n4451), .B(n4450), .ZN(U3256)
         );
  AOI221_X1 U4967 ( .B1(n4455), .B2(n4454), .C1(n4453), .C2(n4454), .A(n4463), 
        .ZN(n4456) );
  AOI211_X1 U4968 ( .C1(n4467), .C2(ADDR_REG_17__SCAN_IN), .A(n4457), .B(n4456), .ZN(n4462) );
  OAI221_X1 U4969 ( .B1(n4460), .B2(n4459), .C1(n4460), .C2(n4458), .A(n4469), 
        .ZN(n4461) );
  OAI211_X1 U4970 ( .C1(n4475), .C2(n4501), .A(n4462), .B(n4461), .ZN(U3257)
         );
  OAI211_X1 U4971 ( .C1(n4471), .C2(n4470), .A(n4469), .B(n4468), .ZN(n4472)
         );
  OAI211_X1 U4972 ( .C1(n4475), .C2(n4474), .A(n4473), .B(n4472), .ZN(U3258)
         );
  OAI22_X1 U4973 ( .A1(n4006), .A2(n4478), .B1(n4477), .B2(n4476), .ZN(n4479)
         );
  INV_X1 U4974 ( .A(n4479), .ZN(n4484) );
  INV_X1 U4975 ( .A(n4480), .ZN(n4481) );
  AOI22_X1 U4976 ( .A1(n4482), .A2(n4489), .B1(n4488), .B2(n4481), .ZN(n4483)
         );
  OAI211_X1 U4977 ( .C1(n4494), .C2(n4485), .A(n4484), .B(n4483), .ZN(U3282)
         );
  AOI22_X1 U4978 ( .A1(n4494), .A2(REG2_REG_3__SCAN_IN), .B1(n4486), .B2(n4689), .ZN(n4492) );
  AOI22_X1 U4979 ( .A1(n4490), .A2(n4489), .B1(n4488), .B2(n4487), .ZN(n4491)
         );
  OAI211_X1 U4980 ( .C1(n4494), .C2(n4493), .A(n4492), .B(n4491), .ZN(U3287)
         );
  AND2_X1 U4981 ( .A1(D_REG_31__SCAN_IN), .A2(n4537), .ZN(U3291) );
  AND2_X1 U4982 ( .A1(D_REG_30__SCAN_IN), .A2(n4537), .ZN(U3292) );
  AND2_X1 U4983 ( .A1(D_REG_29__SCAN_IN), .A2(n4537), .ZN(U3293) );
  AND2_X1 U4984 ( .A1(D_REG_28__SCAN_IN), .A2(n4537), .ZN(U3294) );
  AND2_X1 U4985 ( .A1(D_REG_27__SCAN_IN), .A2(n4537), .ZN(U3295) );
  AND2_X1 U4986 ( .A1(D_REG_26__SCAN_IN), .A2(n4537), .ZN(U3296) );
  AND2_X1 U4987 ( .A1(D_REG_25__SCAN_IN), .A2(n4537), .ZN(U3297) );
  AND2_X1 U4988 ( .A1(D_REG_24__SCAN_IN), .A2(n4537), .ZN(U3298) );
  AND2_X1 U4989 ( .A1(D_REG_23__SCAN_IN), .A2(n4537), .ZN(U3299) );
  INV_X1 U4990 ( .A(D_REG_22__SCAN_IN), .ZN(n4663) );
  NOR2_X1 U4991 ( .A1(n4495), .A2(n4663), .ZN(U3300) );
  AND2_X1 U4992 ( .A1(D_REG_21__SCAN_IN), .A2(n4537), .ZN(U3301) );
  AND2_X1 U4993 ( .A1(D_REG_20__SCAN_IN), .A2(n4537), .ZN(U3302) );
  INV_X1 U4994 ( .A(D_REG_19__SCAN_IN), .ZN(n4558) );
  NOR2_X1 U4995 ( .A1(n4495), .A2(n4558), .ZN(U3303) );
  AND2_X1 U4996 ( .A1(D_REG_18__SCAN_IN), .A2(n4537), .ZN(U3304) );
  AND2_X1 U4997 ( .A1(D_REG_17__SCAN_IN), .A2(n4537), .ZN(U3305) );
  INV_X1 U4998 ( .A(D_REG_16__SCAN_IN), .ZN(n4662) );
  NOR2_X1 U4999 ( .A1(n4495), .A2(n4662), .ZN(U3306) );
  AND2_X1 U5000 ( .A1(D_REG_15__SCAN_IN), .A2(n4537), .ZN(U3307) );
  AND2_X1 U5001 ( .A1(D_REG_14__SCAN_IN), .A2(n4537), .ZN(U3308) );
  AND2_X1 U5002 ( .A1(D_REG_13__SCAN_IN), .A2(n4537), .ZN(U3309) );
  INV_X1 U5003 ( .A(D_REG_12__SCAN_IN), .ZN(n4698) );
  NOR2_X1 U5004 ( .A1(n4495), .A2(n4698), .ZN(U3310) );
  AND2_X1 U5005 ( .A1(D_REG_10__SCAN_IN), .A2(n4537), .ZN(U3312) );
  AND2_X1 U5006 ( .A1(D_REG_9__SCAN_IN), .A2(n4537), .ZN(U3313) );
  AND2_X1 U5007 ( .A1(D_REG_8__SCAN_IN), .A2(n4537), .ZN(U3314) );
  AND2_X1 U5008 ( .A1(D_REG_7__SCAN_IN), .A2(n4537), .ZN(U3315) );
  AND2_X1 U5009 ( .A1(D_REG_6__SCAN_IN), .A2(n4537), .ZN(U3316) );
  AND2_X1 U5010 ( .A1(D_REG_5__SCAN_IN), .A2(n4537), .ZN(U3317) );
  AND2_X1 U5011 ( .A1(D_REG_4__SCAN_IN), .A2(n4537), .ZN(U3318) );
  AND2_X1 U5012 ( .A1(D_REG_3__SCAN_IN), .A2(n4537), .ZN(U3319) );
  AND2_X1 U5013 ( .A1(D_REG_2__SCAN_IN), .A2(n4537), .ZN(U3320) );
  OAI21_X1 U5014 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4496), .ZN(
        n4497) );
  INV_X1 U5015 ( .A(n4497), .ZN(U3329) );
  OAI22_X1 U5016 ( .A1(U3149), .A2(n4498), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4499) );
  INV_X1 U5017 ( .A(n4499), .ZN(U3334) );
  INV_X1 U5018 ( .A(DATAI_17_), .ZN(n4500) );
  AOI22_X1 U5019 ( .A1(STATE_REG_SCAN_IN), .A2(n4501), .B1(n4500), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U5020 ( .A1(U3149), .A2(n4502), .B1(DATAI_16_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4503) );
  INV_X1 U5021 ( .A(n4503), .ZN(U3336) );
  INV_X1 U5022 ( .A(DATAI_15_), .ZN(n4504) );
  AOI22_X1 U5023 ( .A1(STATE_REG_SCAN_IN), .A2(n4505), .B1(n4504), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5024 ( .A(DATAI_14_), .ZN(n4506) );
  AOI22_X1 U5025 ( .A1(STATE_REG_SCAN_IN), .A2(n4507), .B1(n4506), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5026 ( .A(DATAI_13_), .ZN(n4508) );
  AOI22_X1 U5027 ( .A1(STATE_REG_SCAN_IN), .A2(n4509), .B1(n4508), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5028 ( .A(DATAI_12_), .ZN(n4570) );
  AOI22_X1 U5029 ( .A1(STATE_REG_SCAN_IN), .A2(n4510), .B1(n4570), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5030 ( .A1(U3149), .A2(n4511), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4512) );
  INV_X1 U5031 ( .A(n4512), .ZN(U3341) );
  INV_X1 U5032 ( .A(DATAI_10_), .ZN(n4659) );
  AOI22_X1 U5033 ( .A1(STATE_REG_SCAN_IN), .A2(n4513), .B1(n4659), .B2(U3149), 
        .ZN(U3342) );
  OAI22_X1 U5034 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4514) );
  INV_X1 U5035 ( .A(n4514), .ZN(U3352) );
  INV_X1 U5036 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4515) );
  AOI22_X1 U5037 ( .A1(n4530), .A2(n4516), .B1(n4515), .B2(n4528), .ZN(U3467)
         );
  INV_X1 U5038 ( .A(n4517), .ZN(n4519) );
  AOI211_X1 U5039 ( .C1(n4521), .C2(n4520), .A(n4519), .B(n4518), .ZN(n4532)
         );
  INV_X1 U5040 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U5041 ( .A1(n4530), .A2(n4532), .B1(n4522), .B2(n4528), .ZN(U3475)
         );
  NAND3_X1 U5042 ( .A1(n3078), .A2(n4524), .A3(n4523), .ZN(n4525) );
  AND3_X1 U5043 ( .A1(n4527), .A2(n4526), .A3(n4525), .ZN(n4535) );
  INV_X1 U5044 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4529) );
  AOI22_X1 U5045 ( .A1(n4530), .A2(n4535), .B1(n4529), .B2(n4528), .ZN(U3481)
         );
  INV_X1 U5046 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4531) );
  AOI22_X1 U5047 ( .A1(n4536), .A2(n4532), .B1(n4531), .B2(n4533), .ZN(U3522)
         );
  AOI22_X1 U5048 ( .A1(n4536), .A2(n4535), .B1(n4534), .B2(n4533), .ZN(U3525)
         );
  NAND2_X1 U5049 ( .A1(n4537), .A2(D_REG_11__SCAN_IN), .ZN(n4726) );
  INV_X1 U5050 ( .A(DATAI_21_), .ZN(n4539) );
  AOI22_X1 U5051 ( .A1(n4539), .A2(keyinput117), .B1(keyinput93), .B2(n4691), 
        .ZN(n4538) );
  OAI221_X1 U5052 ( .B1(n4539), .B2(keyinput117), .C1(n4691), .C2(keyinput93), 
        .A(n4538), .ZN(n4547) );
  INV_X1 U5053 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4541) );
  AOI22_X1 U5054 ( .A1(n4541), .A2(keyinput105), .B1(n4692), .B2(keyinput97), 
        .ZN(n4540) );
  OAI221_X1 U5055 ( .B1(n4541), .B2(keyinput105), .C1(n4692), .C2(keyinput97), 
        .A(n4540), .ZN(n4546) );
  INV_X1 U5056 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4681) );
  AOI22_X1 U5057 ( .A1(n4681), .A2(keyinput75), .B1(n4679), .B2(keyinput119), 
        .ZN(n4542) );
  OAI221_X1 U5058 ( .B1(n4681), .B2(keyinput75), .C1(n4679), .C2(keyinput119), 
        .A(n4542), .ZN(n4545) );
  AOI22_X1 U5059 ( .A1(n2140), .A2(keyinput66), .B1(keyinput107), .B2(n2785), 
        .ZN(n4543) );
  OAI221_X1 U5060 ( .B1(n2140), .B2(keyinput66), .C1(n2785), .C2(keyinput107), 
        .A(n4543), .ZN(n4544) );
  NOR4_X1 U5061 ( .A1(n4547), .A2(n4546), .A3(n4545), .A4(n4544), .ZN(n4582)
         );
  AOI22_X1 U5062 ( .A1(ADDR_REG_14__SCAN_IN), .A2(keyinput65), .B1(
        IR_REG_29__SCAN_IN), .B2(keyinput95), .ZN(n4548) );
  OAI221_X1 U5063 ( .B1(ADDR_REG_14__SCAN_IN), .B2(keyinput65), .C1(
        IR_REG_29__SCAN_IN), .C2(keyinput95), .A(n4548), .ZN(n4556) );
  AOI22_X1 U5064 ( .A1(REG0_REG_20__SCAN_IN), .A2(keyinput72), .B1(
        REG3_REG_8__SCAN_IN), .B2(keyinput83), .ZN(n4549) );
  OAI221_X1 U5065 ( .B1(REG0_REG_20__SCAN_IN), .B2(keyinput72), .C1(
        REG3_REG_8__SCAN_IN), .C2(keyinput83), .A(n4549), .ZN(n4555) );
  AOI22_X1 U5066 ( .A1(DATAO_REG_29__SCAN_IN), .A2(keyinput96), .B1(n4551), 
        .B2(keyinput84), .ZN(n4550) );
  OAI221_X1 U5067 ( .B1(DATAO_REG_29__SCAN_IN), .B2(keyinput96), .C1(n4551), 
        .C2(keyinput84), .A(n4550), .ZN(n4554) );
  AOI22_X1 U5068 ( .A1(DATAO_REG_2__SCAN_IN), .A2(keyinput70), .B1(
        DATAO_REG_3__SCAN_IN), .B2(keyinput90), .ZN(n4552) );
  OAI221_X1 U5069 ( .B1(DATAO_REG_2__SCAN_IN), .B2(keyinput70), .C1(
        DATAO_REG_3__SCAN_IN), .C2(keyinput90), .A(n4552), .ZN(n4553) );
  NOR4_X1 U5070 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), .ZN(n4581)
         );
  AOI22_X1 U5071 ( .A1(n4662), .A2(keyinput92), .B1(n4558), .B2(keyinput89), 
        .ZN(n4557) );
  OAI221_X1 U5072 ( .B1(n4662), .B2(keyinput92), .C1(n4558), .C2(keyinput89), 
        .A(n4557), .ZN(n4566) );
  AOI22_X1 U5073 ( .A1(n4664), .A2(keyinput78), .B1(n4688), .B2(keyinput81), 
        .ZN(n4559) );
  OAI221_X1 U5074 ( .B1(n4664), .B2(keyinput78), .C1(n4688), .C2(keyinput81), 
        .A(n4559), .ZN(n4565) );
  INV_X1 U5075 ( .A(DATAI_9_), .ZN(n4709) );
  AOI22_X1 U5076 ( .A1(n4709), .A2(keyinput94), .B1(keyinput82), .B2(n4706), 
        .ZN(n4560) );
  OAI221_X1 U5077 ( .B1(n4709), .B2(keyinput94), .C1(n4706), .C2(keyinput82), 
        .A(n4560), .ZN(n4564) );
  AOI22_X1 U5078 ( .A1(n4695), .A2(keyinput68), .B1(keyinput67), .B2(n4562), 
        .ZN(n4561) );
  OAI221_X1 U5079 ( .B1(n4695), .B2(keyinput68), .C1(n4562), .C2(keyinput67), 
        .A(n4561), .ZN(n4563) );
  NOR4_X1 U5080 ( .A1(n4566), .A2(n4565), .A3(n4564), .A4(n4563), .ZN(n4580)
         );
  AOI22_X1 U5081 ( .A1(n4568), .A2(keyinput106), .B1(keyinput80), .B2(n4659), 
        .ZN(n4567) );
  OAI221_X1 U5082 ( .B1(n4568), .B2(keyinput106), .C1(n4659), .C2(keyinput80), 
        .A(n4567), .ZN(n4578) );
  INV_X1 U5083 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5084 ( .A1(n4570), .A2(keyinput102), .B1(keyinput87), .B2(n4678), 
        .ZN(n4569) );
  OAI221_X1 U5085 ( .B1(n4570), .B2(keyinput102), .C1(n4678), .C2(keyinput87), 
        .A(n4569), .ZN(n4577) );
  XOR2_X1 U5086 ( .A(n4325), .B(keyinput121), .Z(n4573) );
  XNOR2_X1 U5087 ( .A(REG1_REG_1__SCAN_IN), .B(keyinput116), .ZN(n4572) );
  XNOR2_X1 U5088 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput86), .ZN(n4571) );
  NAND3_X1 U5089 ( .A1(n4573), .A2(n4572), .A3(n4571), .ZN(n4576) );
  INV_X1 U5090 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4574) );
  XNOR2_X1 U5091 ( .A(n4574), .B(keyinput115), .ZN(n4575) );
  NOR4_X1 U5092 ( .A1(n4578), .A2(n4577), .A3(n4576), .A4(n4575), .ZN(n4579)
         );
  AND4_X1 U5093 ( .A1(n4582), .A2(n4581), .A3(n4580), .A4(n4579), .ZN(n4724)
         );
  OAI22_X1 U5094 ( .A1(REG0_REG_29__SCAN_IN), .A2(keyinput77), .B1(keyinput85), 
        .B2(REG2_REG_29__SCAN_IN), .ZN(n4583) );
  AOI221_X1 U5095 ( .B1(REG0_REG_29__SCAN_IN), .B2(keyinput77), .C1(
        REG2_REG_29__SCAN_IN), .C2(keyinput85), .A(n4583), .ZN(n4590) );
  OAI22_X1 U5096 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput79), .B1(
        DATAO_REG_9__SCAN_IN), .B2(keyinput109), .ZN(n4584) );
  AOI221_X1 U5097 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput79), .C1(keyinput109), .C2(DATAO_REG_9__SCAN_IN), .A(n4584), .ZN(n4589) );
  OAI22_X1 U5098 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput110), .B1(keyinput120), .B2(ADDR_REG_1__SCAN_IN), .ZN(n4585) );
  AOI221_X1 U5099 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput110), .C1(
        ADDR_REG_1__SCAN_IN), .C2(keyinput120), .A(n4585), .ZN(n4588) );
  OAI22_X1 U5100 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput101), .B1(
        REG3_REG_1__SCAN_IN), .B2(keyinput114), .ZN(n4586) );
  AOI221_X1 U5101 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput101), .C1(
        keyinput114), .C2(REG3_REG_1__SCAN_IN), .A(n4586), .ZN(n4587) );
  NAND4_X1 U5102 ( .A1(n4590), .A2(n4589), .A3(n4588), .A4(n4587), .ZN(n4618)
         );
  OAI22_X1 U5103 ( .A1(REG1_REG_18__SCAN_IN), .A2(keyinput71), .B1(
        REG2_REG_18__SCAN_IN), .B2(keyinput76), .ZN(n4591) );
  AOI221_X1 U5104 ( .B1(REG1_REG_18__SCAN_IN), .B2(keyinput71), .C1(keyinput76), .C2(REG2_REG_18__SCAN_IN), .A(n4591), .ZN(n4598) );
  OAI22_X1 U5105 ( .A1(REG2_REG_27__SCAN_IN), .A2(keyinput64), .B1(
        REG2_REG_17__SCAN_IN), .B2(keyinput98), .ZN(n4592) );
  AOI221_X1 U5106 ( .B1(REG2_REG_27__SCAN_IN), .B2(keyinput64), .C1(keyinput98), .C2(REG2_REG_17__SCAN_IN), .A(n4592), .ZN(n4597) );
  OAI22_X1 U5107 ( .A1(DATAI_29_), .A2(keyinput108), .B1(ADDR_REG_3__SCAN_IN), 
        .B2(keyinput122), .ZN(n4593) );
  AOI221_X1 U5108 ( .B1(DATAI_29_), .B2(keyinput108), .C1(keyinput122), .C2(
        ADDR_REG_3__SCAN_IN), .A(n4593), .ZN(n4596) );
  OAI22_X1 U5109 ( .A1(REG2_REG_19__SCAN_IN), .A2(keyinput74), .B1(DATAI_3_), 
        .B2(keyinput111), .ZN(n4594) );
  AOI221_X1 U5110 ( .B1(REG2_REG_19__SCAN_IN), .B2(keyinput74), .C1(
        keyinput111), .C2(DATAI_3_), .A(n4594), .ZN(n4595) );
  NAND4_X1 U5111 ( .A1(n4598), .A2(n4597), .A3(n4596), .A4(n4595), .ZN(n4617)
         );
  OAI22_X1 U5112 ( .A1(IR_REG_20__SCAN_IN), .A2(keyinput100), .B1(keyinput112), 
        .B2(D_REG_1__SCAN_IN), .ZN(n4599) );
  AOI221_X1 U5113 ( .B1(IR_REG_20__SCAN_IN), .B2(keyinput100), .C1(
        D_REG_1__SCAN_IN), .C2(keyinput112), .A(n4599), .ZN(n4606) );
  OAI22_X1 U5114 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput126), .B1(
        IR_REG_27__SCAN_IN), .B2(keyinput99), .ZN(n4600) );
  AOI221_X1 U5115 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput126), .C1(keyinput99), 
        .C2(IR_REG_27__SCAN_IN), .A(n4600), .ZN(n4605) );
  OAI22_X1 U5116 ( .A1(D_REG_22__SCAN_IN), .A2(keyinput124), .B1(
        REG1_REG_16__SCAN_IN), .B2(keyinput103), .ZN(n4601) );
  AOI221_X1 U5117 ( .B1(D_REG_22__SCAN_IN), .B2(keyinput124), .C1(keyinput103), 
        .C2(REG1_REG_16__SCAN_IN), .A(n4601), .ZN(n4604) );
  OAI22_X1 U5118 ( .A1(D_REG_12__SCAN_IN), .A2(keyinput125), .B1(
        D_REG_11__SCAN_IN), .B2(keyinput113), .ZN(n4602) );
  AOI221_X1 U5119 ( .B1(D_REG_12__SCAN_IN), .B2(keyinput125), .C1(keyinput113), 
        .C2(D_REG_11__SCAN_IN), .A(n4602), .ZN(n4603) );
  NAND4_X1 U5120 ( .A1(n4606), .A2(n4605), .A3(n4604), .A4(n4603), .ZN(n4616)
         );
  OAI22_X1 U5121 ( .A1(DATAI_13_), .A2(keyinput127), .B1(keyinput88), .B2(
        REG2_REG_5__SCAN_IN), .ZN(n4607) );
  AOI221_X1 U5122 ( .B1(DATAI_13_), .B2(keyinput127), .C1(REG2_REG_5__SCAN_IN), 
        .C2(keyinput88), .A(n4607), .ZN(n4614) );
  OAI22_X1 U5123 ( .A1(ADDR_REG_11__SCAN_IN), .A2(keyinput104), .B1(keyinput91), .B2(ADDR_REG_9__SCAN_IN), .ZN(n4608) );
  AOI221_X1 U5124 ( .B1(ADDR_REG_11__SCAN_IN), .B2(keyinput104), .C1(
        ADDR_REG_9__SCAN_IN), .C2(keyinput91), .A(n4608), .ZN(n4613) );
  OAI22_X1 U5125 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput69), .B1(keyinput123), 
        .B2(REG0_REG_6__SCAN_IN), .ZN(n4609) );
  AOI221_X1 U5126 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput69), .C1(
        REG0_REG_6__SCAN_IN), .C2(keyinput123), .A(n4609), .ZN(n4612) );
  OAI22_X1 U5127 ( .A1(REG1_REG_14__SCAN_IN), .A2(keyinput73), .B1(keyinput118), .B2(DATAI_7_), .ZN(n4610) );
  AOI221_X1 U5128 ( .B1(REG1_REG_14__SCAN_IN), .B2(keyinput73), .C1(DATAI_7_), 
        .C2(keyinput118), .A(n4610), .ZN(n4611) );
  NAND4_X1 U5129 ( .A1(n4614), .A2(n4613), .A3(n4612), .A4(n4611), .ZN(n4615)
         );
  NOR4_X1 U5130 ( .A1(n4618), .A2(n4617), .A3(n4616), .A4(n4615), .ZN(n4723)
         );
  AOI22_X1 U5131 ( .A1(REG1_REG_0__SCAN_IN), .A2(keyinput22), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput2), .ZN(n4619) );
  OAI221_X1 U5132 ( .B1(REG1_REG_0__SCAN_IN), .B2(keyinput22), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput2), .A(n4619), .ZN(n4626) );
  AOI22_X1 U5133 ( .A1(REG2_REG_17__SCAN_IN), .A2(keyinput34), .B1(
        REG3_REG_4__SCAN_IN), .B2(keyinput46), .ZN(n4620) );
  OAI221_X1 U5134 ( .B1(REG2_REG_17__SCAN_IN), .B2(keyinput34), .C1(
        REG3_REG_4__SCAN_IN), .C2(keyinput46), .A(n4620), .ZN(n4625) );
  AOI22_X1 U5135 ( .A1(DATAI_7_), .A2(keyinput54), .B1(DATAI_12_), .B2(
        keyinput38), .ZN(n4621) );
  OAI221_X1 U5136 ( .B1(DATAI_7_), .B2(keyinput54), .C1(DATAI_12_), .C2(
        keyinput38), .A(n4621), .ZN(n4624) );
  AOI22_X1 U5137 ( .A1(DATAI_3_), .A2(keyinput47), .B1(REG1_REG_10__SCAN_IN), 
        .B2(keyinput42), .ZN(n4622) );
  OAI221_X1 U5138 ( .B1(DATAI_3_), .B2(keyinput47), .C1(REG1_REG_10__SCAN_IN), 
        .C2(keyinput42), .A(n4622), .ZN(n4623) );
  NOR4_X1 U5139 ( .A1(n4626), .A2(n4625), .A3(n4624), .A4(n4623), .ZN(n4656)
         );
  AOI22_X1 U5140 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput15), .B1(DATAI_29_), 
        .B2(keyinput44), .ZN(n4627) );
  OAI221_X1 U5141 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput15), .C1(DATAI_29_), 
        .C2(keyinput44), .A(n4627), .ZN(n4634) );
  AOI22_X1 U5142 ( .A1(DATAO_REG_9__SCAN_IN), .A2(keyinput45), .B1(
        REG0_REG_29__SCAN_IN), .B2(keyinput13), .ZN(n4628) );
  OAI221_X1 U5143 ( .B1(DATAO_REG_9__SCAN_IN), .B2(keyinput45), .C1(
        REG0_REG_29__SCAN_IN), .C2(keyinput13), .A(n4628), .ZN(n4633) );
  AOI22_X1 U5144 ( .A1(REG2_REG_22__SCAN_IN), .A2(keyinput41), .B1(
        REG3_REG_24__SCAN_IN), .B2(keyinput20), .ZN(n4629) );
  OAI221_X1 U5145 ( .B1(REG2_REG_22__SCAN_IN), .B2(keyinput41), .C1(
        REG3_REG_24__SCAN_IN), .C2(keyinput20), .A(n4629), .ZN(n4632) );
  AOI22_X1 U5146 ( .A1(ADDR_REG_1__SCAN_IN), .A2(keyinput56), .B1(DATAI_21_), 
        .B2(keyinput53), .ZN(n4630) );
  OAI221_X1 U5147 ( .B1(ADDR_REG_1__SCAN_IN), .B2(keyinput56), .C1(DATAI_21_), 
        .C2(keyinput53), .A(n4630), .ZN(n4631) );
  NOR4_X1 U5148 ( .A1(n4634), .A2(n4633), .A3(n4632), .A4(n4631), .ZN(n4655)
         );
  AOI22_X1 U5149 ( .A1(ADDR_REG_6__SCAN_IN), .A2(keyinput43), .B1(
        ADDR_REG_9__SCAN_IN), .B2(keyinput27), .ZN(n4635) );
  OAI221_X1 U5150 ( .B1(ADDR_REG_6__SCAN_IN), .B2(keyinput43), .C1(
        ADDR_REG_9__SCAN_IN), .C2(keyinput27), .A(n4635), .ZN(n4642) );
  AOI22_X1 U5151 ( .A1(ADDR_REG_17__SCAN_IN), .A2(keyinput51), .B1(
        REG1_REG_1__SCAN_IN), .B2(keyinput52), .ZN(n4636) );
  OAI221_X1 U5152 ( .B1(ADDR_REG_17__SCAN_IN), .B2(keyinput51), .C1(
        REG1_REG_1__SCAN_IN), .C2(keyinput52), .A(n4636), .ZN(n4641) );
  AOI22_X1 U5153 ( .A1(REG2_REG_5__SCAN_IN), .A2(keyinput24), .B1(DATAI_13_), 
        .B2(keyinput63), .ZN(n4637) );
  OAI221_X1 U5154 ( .B1(REG2_REG_5__SCAN_IN), .B2(keyinput24), .C1(DATAI_13_), 
        .C2(keyinput63), .A(n4637), .ZN(n4640) );
  AOI22_X1 U5155 ( .A1(REG1_REG_14__SCAN_IN), .A2(keyinput9), .B1(
        REG0_REG_15__SCAN_IN), .B2(keyinput57), .ZN(n4638) );
  OAI221_X1 U5156 ( .B1(REG1_REG_14__SCAN_IN), .B2(keyinput9), .C1(
        REG0_REG_15__SCAN_IN), .C2(keyinput57), .A(n4638), .ZN(n4639) );
  NOR4_X1 U5157 ( .A1(n4642), .A2(n4641), .A3(n4640), .A4(n4639), .ZN(n4654)
         );
  AOI22_X1 U5158 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput48), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput5), .ZN(n4643) );
  OAI221_X1 U5159 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput48), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput5), .A(n4643), .ZN(n4652) );
  AOI22_X1 U5160 ( .A1(D_REG_19__SCAN_IN), .A2(keyinput25), .B1(
        IR_REG_20__SCAN_IN), .B2(keyinput36), .ZN(n4644) );
  OAI221_X1 U5161 ( .B1(D_REG_19__SCAN_IN), .B2(keyinput25), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput36), .A(n4644), .ZN(n4651) );
  AOI22_X1 U5162 ( .A1(DATAO_REG_17__SCAN_IN), .A2(keyinput3), .B1(
        REG3_REG_8__SCAN_IN), .B2(keyinput19), .ZN(n4645) );
  OAI221_X1 U5163 ( .B1(DATAO_REG_17__SCAN_IN), .B2(keyinput3), .C1(
        REG3_REG_8__SCAN_IN), .C2(keyinput19), .A(n4645), .ZN(n4650) );
  INV_X1 U5164 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4648) );
  AOI22_X1 U5165 ( .A1(n4648), .A2(keyinput0), .B1(keyinput7), .B2(n4647), 
        .ZN(n4646) );
  OAI221_X1 U5166 ( .B1(n4648), .B2(keyinput0), .C1(n4647), .C2(keyinput7), 
        .A(n4646), .ZN(n4649) );
  NOR4_X1 U5167 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(n4653)
         );
  NAND4_X1 U5168 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), .ZN(n4722)
         );
  AOI22_X1 U5169 ( .A1(n4659), .A2(keyinput16), .B1(keyinput59), .B2(n4658), 
        .ZN(n4657) );
  OAI221_X1 U5170 ( .B1(n4659), .B2(keyinput16), .C1(n4658), .C2(keyinput59), 
        .A(n4657), .ZN(n4671) );
  AOI22_X1 U5171 ( .A1(n4662), .A2(keyinput28), .B1(keyinput39), .B2(n4661), 
        .ZN(n4660) );
  OAI221_X1 U5172 ( .B1(n4662), .B2(keyinput28), .C1(n4661), .C2(keyinput39), 
        .A(n4660), .ZN(n4670) );
  XNOR2_X1 U5173 ( .A(n4663), .B(keyinput60), .ZN(n4669) );
  XOR2_X1 U5174 ( .A(n4664), .B(keyinput14), .Z(n4667) );
  XNOR2_X1 U5175 ( .A(IR_REG_9__SCAN_IN), .B(keyinput62), .ZN(n4666) );
  XNOR2_X1 U5176 ( .A(IR_REG_27__SCAN_IN), .B(keyinput35), .ZN(n4665) );
  NAND3_X1 U5177 ( .A1(n4667), .A2(n4666), .A3(n4665), .ZN(n4668) );
  NOR4_X1 U5178 ( .A1(n4671), .A2(n4670), .A3(n4669), .A4(n4668), .ZN(n4720)
         );
  INV_X1 U5179 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5180 ( .A1(n4673), .A2(keyinput58), .B1(n2709), .B2(keyinput50), 
        .ZN(n4672) );
  OAI221_X1 U5181 ( .B1(n4673), .B2(keyinput58), .C1(n2709), .C2(keyinput50), 
        .A(n4672), .ZN(n4686) );
  AOI22_X1 U5182 ( .A1(n4676), .A2(keyinput12), .B1(n4675), .B2(keyinput10), 
        .ZN(n4674) );
  OAI221_X1 U5183 ( .B1(n4676), .B2(keyinput12), .C1(n4675), .C2(keyinput10), 
        .A(n4674), .ZN(n4685) );
  AOI22_X1 U5184 ( .A1(n4679), .A2(keyinput55), .B1(keyinput23), .B2(n4678), 
        .ZN(n4677) );
  OAI221_X1 U5185 ( .B1(n4679), .B2(keyinput55), .C1(n4678), .C2(keyinput23), 
        .A(n4677), .ZN(n4684) );
  INV_X1 U5186 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n4682) );
  AOI22_X1 U5187 ( .A1(n4682), .A2(keyinput40), .B1(n4681), .B2(keyinput11), 
        .ZN(n4680) );
  OAI221_X1 U5188 ( .B1(n4682), .B2(keyinput40), .C1(n4681), .C2(keyinput11), 
        .A(n4680), .ZN(n4683) );
  NOR4_X1 U5189 ( .A1(n4686), .A2(n4685), .A3(n4684), .A4(n4683), .ZN(n4719)
         );
  AOI22_X1 U5190 ( .A1(n4689), .A2(keyinput37), .B1(n4688), .B2(keyinput17), 
        .ZN(n4687) );
  OAI221_X1 U5191 ( .B1(n4689), .B2(keyinput37), .C1(n4688), .C2(keyinput17), 
        .A(n4687), .ZN(n4702) );
  AOI22_X1 U5192 ( .A1(n4692), .A2(keyinput33), .B1(keyinput29), .B2(n4691), 
        .ZN(n4690) );
  OAI221_X1 U5193 ( .B1(n4692), .B2(keyinput33), .C1(n4691), .C2(keyinput29), 
        .A(n4690), .ZN(n4701) );
  INV_X1 U5194 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4694) );
  AOI22_X1 U5195 ( .A1(n4695), .A2(keyinput4), .B1(keyinput1), .B2(n4694), 
        .ZN(n4693) );
  OAI221_X1 U5196 ( .B1(n4695), .B2(keyinput4), .C1(n4694), .C2(keyinput1), 
        .A(n4693), .ZN(n4700) );
  INV_X1 U5197 ( .A(D_REG_11__SCAN_IN), .ZN(n4697) );
  AOI22_X1 U5198 ( .A1(n4698), .A2(keyinput61), .B1(keyinput49), .B2(n4697), 
        .ZN(n4696) );
  OAI221_X1 U5199 ( .B1(n4698), .B2(keyinput61), .C1(n4697), .C2(keyinput49), 
        .A(n4696), .ZN(n4699) );
  NOR4_X1 U5200 ( .A1(n4702), .A2(n4701), .A3(n4700), .A4(n4699), .ZN(n4718)
         );
  AOI22_X1 U5201 ( .A1(n4704), .A2(keyinput32), .B1(n3834), .B2(keyinput21), 
        .ZN(n4703) );
  OAI221_X1 U5202 ( .B1(n4704), .B2(keyinput32), .C1(n3834), .C2(keyinput21), 
        .A(n4703), .ZN(n4716) );
  AOI22_X1 U5203 ( .A1(n4707), .A2(keyinput6), .B1(n4706), .B2(keyinput18), 
        .ZN(n4705) );
  OAI221_X1 U5204 ( .B1(n4707), .B2(keyinput6), .C1(n4706), .C2(keyinput18), 
        .A(n4705), .ZN(n4715) );
  AOI22_X1 U5205 ( .A1(n4710), .A2(keyinput26), .B1(n4709), .B2(keyinput30), 
        .ZN(n4708) );
  OAI221_X1 U5206 ( .B1(n4710), .B2(keyinput26), .C1(n4709), .C2(keyinput30), 
        .A(n4708), .ZN(n4714) );
  XNOR2_X1 U5207 ( .A(REG0_REG_20__SCAN_IN), .B(keyinput8), .ZN(n4712) );
  XNOR2_X1 U5208 ( .A(IR_REG_29__SCAN_IN), .B(keyinput31), .ZN(n4711) );
  NAND2_X1 U5209 ( .A1(n4712), .A2(n4711), .ZN(n4713) );
  NOR4_X1 U5210 ( .A1(n4716), .A2(n4715), .A3(n4714), .A4(n4713), .ZN(n4717)
         );
  NAND4_X1 U5211 ( .A1(n4720), .A2(n4719), .A3(n4718), .A4(n4717), .ZN(n4721)
         );
  AOI211_X1 U5212 ( .C1(n4724), .C2(n4723), .A(n4722), .B(n4721), .ZN(n4725)
         );
  XNOR2_X1 U5213 ( .A(n4726), .B(n4725), .ZN(U3311) );
  NAND2_X1 U3857 ( .A1(n3089), .A2(n3088), .ZN(n3115) );
  NAND2_X1 U3802 ( .A1(n3026), .A2(n3025), .ZN(n3089) );
  CLKBUF_X1 U2295 ( .A(n3369), .Z(n2058) );
  OR2_X2 U2297 ( .A1(n3369), .A2(n4021), .ZN(n3358) );
  CLKBUF_X2 U2307 ( .A(n2307), .Z(n2054) );
  CLKBUF_X1 U2311 ( .A(n4361), .Z(n2055) );
  INV_X1 U2316 ( .A(n2931), .ZN(n3160) );
  INV_X2 U2360 ( .A(n4494), .ZN(n4006) );
endmodule

