

module b15_C_AntiSAT_k_256_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
         keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
         keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
         keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
         keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
         keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
         keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
         keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
         keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
         keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
         keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
         keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
         keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
         keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
         keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
         keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
         keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
         keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
         keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
         keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
         keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
         keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
         keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
         keyinput239, keyinput240, keyinput241, keyinput242, keyinput243,
         keyinput244, keyinput245, keyinput246, keyinput247, keyinput248,
         keyinput249, keyinput250, keyinput251, keyinput252, keyinput253,
         keyinput254, keyinput255;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168;

  OR2_X1 U3627 ( .A1(n3740), .A2(n3275), .ZN(n6099) );
  OR2_X1 U3628 ( .A1(n3201), .A2(n4988), .ZN(n5119) );
  AND2_X2 U3629 ( .A1(n3721), .A2(n3720), .ZN(n6131) );
  CLKBUF_X2 U3630 ( .A(n3506), .Z(n5476) );
  CLKBUF_X1 U3631 ( .A(n3435), .Z(n4294) );
  AND2_X1 U3632 ( .A1(n4032), .A2(n4172), .ZN(n3511) );
  AND2_X1 U3633 ( .A1(n4033), .A2(n4172), .ZN(n3526) );
  AND2_X2 U3634 ( .A1(n3311), .A2(n4033), .ZN(n3400) );
  AND2_X2 U3635 ( .A1(n3311), .A2(n3317), .ZN(n5398) );
  AND2_X1 U3636 ( .A1(n4174), .A2(n4032), .ZN(n3494) );
  AND2_X1 U3638 ( .A1(n3449), .A2(n3940), .ZN(n3464) );
  XNOR2_X1 U3639 ( .A(n3721), .B(n3710), .ZN(n4413) );
  AND4_X1 U3640 ( .A1(n3464), .A2(n3463), .A3(n3462), .A4(n3461), .ZN(n3470)
         );
  XNOR2_X1 U3641 ( .A(n3662), .B(n3663), .ZN(n4215) );
  AOI21_X1 U3642 ( .B1(n4060), .B2(n7028), .A(n3574), .ZN(n3600) );
  INV_X1 U3643 ( .A(n4097), .ZN(n3473) );
  AND2_X1 U3644 ( .A1(n4097), .A2(n3447), .ZN(n4144) );
  NOR2_X1 U3645 ( .A1(n3447), .A2(n4097), .ZN(n3826) );
  INV_X1 U3646 ( .A(n4144), .ZN(n5526) );
  INV_X1 U3647 ( .A(n6515), .ZN(n6503) );
  AND2_X1 U3648 ( .A1(n5179), .A2(n3210), .ZN(n5290) );
  INV_X1 U3649 ( .A(n6518), .ZN(n6541) );
  AND2_X1 U3650 ( .A1(n3284), .A2(n3206), .ZN(n3179) );
  AND2_X1 U3651 ( .A1(n6263), .A2(n5256), .ZN(n5095) );
  NAND3_X4 U3652 ( .A1(n3292), .A2(n3294), .A3(n3363), .ZN(n3444) );
  NAND2_X2 U3655 ( .A1(n3599), .A2(n3598), .ZN(n3639) );
  NAND2_X2 U3656 ( .A1(n3969), .A2(n3355), .ZN(n3452) );
  INV_X2 U3657 ( .A(n3446), .ZN(n3355) );
  NOR2_X2 U3658 ( .A1(n3740), .A2(n3186), .ZN(n5531) );
  NOR2_X2 U3659 ( .A1(n4986), .A2(n4985), .ZN(n5140) );
  OR2_X1 U3660 ( .A1(n5550), .A2(n5549), .ZN(n6139) );
  AND2_X1 U3661 ( .A1(n3215), .A2(n3193), .ZN(n3183) );
  AND3_X1 U3662 ( .A1(n4329), .A2(n4328), .A3(n4327), .ZN(n4503) );
  NAND2_X1 U3663 ( .A1(n6689), .A2(n3640), .ZN(n4255) );
  CLKBUF_X2 U3664 ( .A(n6648), .Z(n6658) );
  CLKBUF_X2 U3665 ( .A(n4263), .Z(n3196) );
  INV_X2 U3666 ( .A(n3913), .ZN(n5537) );
  BUF_X2 U3667 ( .A(n3387), .Z(n5478) );
  CLKBUF_X2 U3668 ( .A(n3365), .Z(n5307) );
  CLKBUF_X2 U3669 ( .A(n3489), .Z(n5480) );
  CLKBUF_X2 U3670 ( .A(n3488), .Z(n5332) );
  BUF_X2 U3671 ( .A(n5398), .Z(n5486) );
  BUF_X2 U3672 ( .A(n3526), .Z(n5487) );
  CLKBUF_X2 U3673 ( .A(n3494), .Z(n5477) );
  OR2_X1 U3674 ( .A1(n5558), .A2(n3228), .ZN(n3227) );
  NOR3_X1 U3675 ( .A1(n5551), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n6216), 
        .ZN(n5552) );
  NAND2_X1 U3676 ( .A1(n6139), .A2(n3198), .ZN(n5551) );
  OR2_X1 U3677 ( .A1(n5557), .A2(n6681), .ZN(n3228) );
  AOI21_X1 U3678 ( .B1(n6031), .B2(n6030), .A(n6029), .ZN(n6331) );
  NAND2_X1 U3679 ( .A1(n6030), .A2(n5933), .ZN(n6085) );
  NAND2_X1 U3680 ( .A1(n4743), .A2(n3183), .ZN(n3180) );
  NAND2_X1 U3681 ( .A1(n4583), .A2(n3727), .ZN(n4745) );
  AOI21_X1 U3682 ( .B1(n3234), .B2(n3232), .A(n3204), .ZN(n3231) );
  NOR2_X1 U3683 ( .A1(n5095), .A2(n3219), .ZN(n3218) );
  NOR2_X1 U3684 ( .A1(n3733), .A2(n3235), .ZN(n3234) );
  OR3_X1 U3685 ( .A1(n5300), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3185) );
  NAND2_X1 U3686 ( .A1(n6678), .A2(n6677), .ZN(n6676) );
  NAND2_X1 U3687 ( .A1(n4255), .A2(n4254), .ZN(n4253) );
  XNOR2_X1 U3688 ( .A(n3681), .B(n6751), .ZN(n6677) );
  NAND2_X1 U3689 ( .A1(n4243), .A2(n4242), .ZN(n4328) );
  NAND2_X1 U3690 ( .A1(n3593), .A2(n3592), .ZN(n4376) );
  OAI21_X1 U3691 ( .B1(n6817), .B2(n3762), .A(n3628), .ZN(n4076) );
  OR2_X1 U3692 ( .A1(n4895), .A2(n4894), .ZN(n4956) );
  AND2_X1 U3694 ( .A1(n4509), .A2(n4508), .ZN(n4589) );
  CLKBUF_X1 U3695 ( .A(n3971), .Z(n6995) );
  NAND2_X1 U3696 ( .A1(n3257), .A2(n3256), .ZN(n4447) );
  NAND2_X1 U3697 ( .A1(n3470), .A2(n3938), .ZN(n3503) );
  NAND2_X1 U3698 ( .A1(n4155), .A2(n3838), .ZN(n4249) );
  AND2_X1 U3699 ( .A1(n3469), .A2(n3468), .ZN(n3938) );
  NAND2_X1 U3700 ( .A1(n3438), .A2(n3437), .ZN(n3442) );
  OR2_X1 U3701 ( .A1(n3816), .A2(n3790), .ZN(n3290) );
  NAND2_X1 U3702 ( .A1(n3477), .A2(n3295), .ZN(n3926) );
  NAND2_X1 U3703 ( .A1(n3768), .A2(n4294), .ZN(n3790) );
  NOR2_X2 U3704 ( .A1(n3184), .A2(n6930), .ZN(n3972) );
  NAND3_X1 U3705 ( .A1(n3324), .A2(n3323), .A3(n3322), .ZN(n3435) );
  NAND2_X1 U3706 ( .A1(n3809), .A2(n4289), .ZN(n3932) );
  CLKBUF_X1 U3707 ( .A(n3446), .Z(n3430) );
  INV_X1 U3708 ( .A(n3446), .ZN(n4279) );
  AND2_X1 U3709 ( .A1(n4097), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3768) );
  OR2_X1 U3710 ( .A1(n3517), .A2(n3516), .ZN(n3723) );
  AND3_X1 U3711 ( .A1(n3310), .A2(n3309), .A3(n3308), .ZN(n3324) );
  OR2_X1 U3712 ( .A1(n3532), .A2(n3531), .ZN(n3626) );
  NAND2_X1 U3713 ( .A1(n3334), .A2(n3333), .ZN(n3434) );
  AND4_X1 U3714 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3334)
         );
  AND4_X1 U3715 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3333)
         );
  AND4_X1 U3716 ( .A1(n3369), .A2(n3368), .A3(n3367), .A4(n3366), .ZN(n3375)
         );
  AND4_X1 U3717 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n3354)
         );
  AND4_X1 U3718 ( .A1(n3342), .A2(n3341), .A3(n3340), .A4(n3339), .ZN(n3353)
         );
  AND4_X1 U3719 ( .A1(n3346), .A2(n3345), .A3(n3344), .A4(n3343), .ZN(n3352)
         );
  AND4_X1 U3720 ( .A1(n3350), .A2(n3349), .A3(n3348), .A4(n3347), .ZN(n3351)
         );
  AND4_X1 U3721 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3408)
         );
  AND4_X1 U3722 ( .A1(n3404), .A2(n3403), .A3(n3402), .A4(n3401), .ZN(n3405)
         );
  AND4_X1 U3723 ( .A1(n3425), .A2(n3424), .A3(n3423), .A4(n3422), .ZN(n3426)
         );
  AND4_X1 U3724 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(n3429)
         );
  AND4_X1 U3725 ( .A1(n3420), .A2(n3419), .A3(n3418), .A4(n3417), .ZN(n3427)
         );
  AND4_X1 U3726 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3428)
         );
  AND4_X1 U3727 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3323)
         );
  AND4_X1 U3728 ( .A1(n3321), .A2(n3320), .A3(n3319), .A4(n3318), .ZN(n3322)
         );
  AND4_X1 U3729 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3292)
         );
  BUF_X2 U3730 ( .A(n3519), .Z(n5485) );
  BUF_X2 U3731 ( .A(n3524), .Z(n3525) );
  BUF_X2 U3732 ( .A(n3370), .Z(n5475) );
  AND2_X2 U3733 ( .A1(n3317), .A2(n3312), .ZN(n3365) );
  AND2_X2 U3734 ( .A1(n3743), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4039)
         );
  INV_X1 U3735 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3298) );
  AOI21_X1 U3736 ( .B1(n3215), .B2(n3217), .A(n3203), .ZN(n3213) );
  NAND2_X2 U3737 ( .A1(n3180), .A2(n3181), .ZN(n5250) );
  INV_X1 U3739 ( .A(n3193), .ZN(n3182) );
  INV_X2 U3740 ( .A(n3969), .ZN(n3184) );
  NOR2_X1 U3741 ( .A1(n6114), .A2(n3185), .ZN(n5301) );
  NAND2_X1 U3742 ( .A1(n6090), .A2(n6115), .ZN(n6114) );
  OR2_X1 U3743 ( .A1(n3275), .A2(n3964), .ZN(n3186) );
  INV_X1 U3744 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3187) );
  AND2_X1 U3745 ( .A1(n3815), .A2(n3433), .ZN(n3450) );
  BUF_X8 U3746 ( .A(n3643), .Z(n5333) );
  XNOR2_X1 U3747 ( .A(n3660), .B(n6784), .ZN(n4254) );
  NAND3_X1 U3748 ( .A1(n3486), .A2(n3485), .A3(n3484), .ZN(n3551) );
  NAND2_X1 U3749 ( .A1(n6676), .A2(n3682), .ZN(n3188) );
  INV_X1 U3750 ( .A(n5250), .ZN(n3189) );
  INV_X1 U3751 ( .A(n3189), .ZN(n3190) );
  BUF_X1 U3752 ( .A(n3825), .Z(n3191) );
  NAND2_X1 U3753 ( .A1(n3813), .A2(n3479), .ZN(n3825) );
  NAND2_X1 U3754 ( .A1(n4253), .A2(n3661), .ZN(n3192) );
  OR2_X1 U3755 ( .A1(n3194), .A2(n3206), .ZN(n3193) );
  INV_X1 U3756 ( .A(n3731), .ZN(n3194) );
  AND2_X1 U3757 ( .A1(n3213), .A2(n3731), .ZN(n3195) );
  NAND2_X1 U3758 ( .A1(n3641), .A2(n3602), .ZN(n6284) );
  AND2_X4 U3759 ( .A1(n3479), .A2(n4097), .ZN(n3596) );
  INV_X2 U3760 ( .A(n3434), .ZN(n3969) );
  NAND2_X2 U3761 ( .A1(n4745), .A2(n4744), .ZN(n4743) );
  AND2_X1 U3762 ( .A1(n3740), .A2(n3277), .ZN(n5532) );
  NAND2_X2 U3763 ( .A1(n6114), .A2(n3739), .ZN(n3740) );
  NAND2_X2 U3764 ( .A1(n3736), .A2(n6147), .ZN(n6146) );
  NAND2_X1 U3765 ( .A1(n3618), .A2(n3617), .ZN(n4154) );
  AOI21_X2 U3766 ( .B1(n5531), .B2(n5518), .A(n5301), .ZN(n5302) );
  NOR2_X4 U3767 ( .A1(n3478), .A2(n3296), .ZN(n3813) );
  NAND3_X2 U3768 ( .A1(n3442), .A2(n3441), .A3(n3440), .ZN(n3478) );
  OAI21_X4 U3769 ( .B1(n5250), .B2(n3233), .A(n3231), .ZN(n6264) );
  AND2_X4 U3770 ( .A1(n3311), .A2(n4039), .ZN(n3488) );
  XNOR2_X1 U3771 ( .A(n3608), .B(n3612), .ZN(n4263) );
  XNOR2_X2 U3772 ( .A(n3641), .B(n4376), .ZN(n4208) );
  NAND2_X2 U3773 ( .A1(n3238), .A2(n3237), .ZN(n3641) );
  OAI211_X1 U3774 ( .C1(n4016), .C2(n3475), .A(n3926), .B(n3825), .ZN(n3480)
         );
  NAND2_X1 U3775 ( .A1(n3457), .A2(n3456), .ZN(n3505) );
  NAND2_X1 U3776 ( .A1(n3554), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3457) );
  AND2_X1 U3777 ( .A1(n6165), .A2(n3951), .ZN(n3735) );
  INV_X1 U3778 ( .A(n5019), .ZN(n3219) );
  AND2_X2 U3779 ( .A1(n3505), .A2(n3503), .ZN(n3553) );
  OR2_X1 U3780 ( .A1(n4040), .A2(n7033), .ZN(n4336) );
  NOR2_X1 U3781 ( .A1(n3444), .A2(n6930), .ZN(n5510) );
  INV_X1 U3782 ( .A(n4336), .ZN(n4340) );
  NAND2_X1 U3783 ( .A1(n3264), .A2(n3262), .ZN(n3261) );
  INV_X1 U3784 ( .A(n5538), .ZN(n3264) );
  NAND2_X1 U3785 ( .A1(n4173), .A2(n7028), .ZN(n3593) );
  NOR2_X1 U3786 ( .A1(n6227), .A2(n3957), .ZN(n6214) );
  OAI21_X1 U3787 ( .B1(n3458), .B2(n3460), .A(n3447), .ZN(n3461) );
  NAND2_X1 U3788 ( .A1(n3642), .A2(n4376), .ZN(n3662) );
  CLKBUF_X1 U3789 ( .A(n3421), .Z(n5338) );
  NOR2_X1 U3790 ( .A1(n3458), .A2(n3932), .ZN(n3815) );
  OR2_X1 U3791 ( .A1(n4294), .A2(n7028), .ZN(n3562) );
  OR2_X1 U3792 ( .A1(n4097), .A2(n7028), .ZN(n3561) );
  NOR2_X1 U3793 ( .A1(n5988), .A2(n3250), .ZN(n3249) );
  INV_X1 U3794 ( .A(n6002), .ZN(n3250) );
  NOR2_X1 U3795 ( .A1(n5202), .A2(n3244), .ZN(n3243) );
  INV_X1 U3796 ( .A(n5178), .ZN(n3244) );
  INV_X1 U3797 ( .A(n5369), .ZN(n5501) );
  NAND2_X1 U3798 ( .A1(n4504), .A2(n3255), .ZN(n3254) );
  INV_X1 U3799 ( .A(n4577), .ZN(n3255) );
  INV_X1 U3800 ( .A(n4507), .ZN(n4504) );
  NOR2_X1 U3801 ( .A1(n5945), .A2(n5524), .ZN(n5535) );
  NAND2_X1 U3802 ( .A1(n3708), .A2(n3707), .ZN(n3721) );
  AND2_X1 U3803 ( .A1(n6263), .A2(n3732), .ZN(n3733) );
  INV_X1 U3804 ( .A(n5247), .ZN(n3235) );
  INV_X1 U3805 ( .A(n5248), .ZN(n3232) );
  NAND2_X1 U3806 ( .A1(n4968), .A2(n3269), .ZN(n3268) );
  INV_X1 U3807 ( .A(n4957), .ZN(n3269) );
  NAND2_X1 U3808 ( .A1(n3830), .A2(n4097), .ZN(n3917) );
  OR2_X1 U3809 ( .A1(n3500), .A2(n3499), .ZN(n3613) );
  NAND2_X1 U3810 ( .A1(n3562), .A2(n3561), .ZN(n3781) );
  INV_X1 U3811 ( .A(n3576), .ZN(n3281) );
  OR2_X1 U3812 ( .A1(n3756), .A2(n3755), .ZN(n3758) );
  NOR2_X1 U3813 ( .A1(n3790), .A2(n3762), .ZN(n3791) );
  INV_X1 U3814 ( .A(n3596), .ZN(n7162) );
  NAND2_X1 U3815 ( .A1(n7157), .A2(n3980), .ZN(n6504) );
  AND2_X1 U3816 ( .A1(n6930), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5509) );
  AND2_X1 U3817 ( .A1(n3246), .A2(n3247), .ZN(n3245) );
  INV_X1 U3818 ( .A(n5964), .ZN(n3246) );
  NAND2_X1 U3819 ( .A1(n5318), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5364)
         );
  NOR2_X1 U3820 ( .A1(n5136), .A2(n5134), .ZN(n5175) );
  NAND2_X1 U3821 ( .A1(n5175), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5198)
         );
  NAND2_X1 U3822 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n4414), .ZN(n4486)
         );
  OR2_X1 U3823 ( .A1(n5535), .A2(n5537), .ZN(n3263) );
  AND2_X1 U3824 ( .A1(n6120), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5554)
         );
  INV_X1 U3825 ( .A(n5551), .ZN(n6121) );
  OR2_X1 U3826 ( .A1(n6263), .A2(n6388), .ZN(n5248) );
  OR2_X1 U3827 ( .A1(n6263), .A2(n5841), .ZN(n3729) );
  NAND2_X1 U3828 ( .A1(n3214), .A2(n3213), .ZN(n3284) );
  OAI21_X2 U3829 ( .B1(n3553), .B2(n3552), .A(n3551), .ZN(n3575) );
  AOI22_X1 U3830 ( .A1(n3365), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3363) );
  AND2_X1 U3831 ( .A1(n4096), .A2(n4095), .ZN(n6590) );
  OAI21_X1 U3832 ( .B1(n3261), .B2(n6775), .A(n3199), .ZN(n3260) );
  XNOR2_X1 U3833 ( .A(n3273), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6082)
         );
  NAND2_X1 U3834 ( .A1(n3276), .A2(n3274), .ZN(n3273) );
  NAND2_X1 U3835 ( .A1(n5532), .A2(n5539), .ZN(n3276) );
  NAND2_X1 U3836 ( .A1(n5531), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3274) );
  OR2_X1 U3837 ( .A1(n6369), .A2(n3955), .ZN(n6227) );
  OR2_X1 U3838 ( .A1(n6743), .A2(n6746), .ZN(n6750) );
  INV_X1 U3839 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7000) );
  NAND2_X1 U3840 ( .A1(n3534), .A2(n3622), .ZN(n3623) );
  NAND2_X1 U3841 ( .A1(n3620), .A2(n3621), .ZN(n3624) );
  INV_X1 U3842 ( .A(n3738), .ZN(n3287) );
  OR2_X1 U3843 ( .A1(n3695), .A2(n3694), .ZN(n3712) );
  NAND2_X1 U3844 ( .A1(n3445), .A2(n3444), .ZN(n3471) );
  NAND2_X1 U3845 ( .A1(n3816), .A2(n3596), .ZN(n3818) );
  AND2_X1 U3846 ( .A1(n4142), .A2(n3444), .ZN(n3364) );
  INV_X1 U3847 ( .A(n3452), .ZN(n3816) );
  NAND2_X1 U3848 ( .A1(n5398), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3307)
         );
  NAND2_X1 U3849 ( .A1(n5438), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U3850 ( .A1(n3370), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3313) );
  NOR2_X1 U3851 ( .A1(n5559), .A2(n3248), .ZN(n3247) );
  INV_X1 U3852 ( .A(n3249), .ZN(n3248) );
  NAND2_X1 U3853 ( .A1(n3680), .A2(n3679), .ZN(n3681) );
  XNOR2_X1 U3854 ( .A(n3683), .B(n3684), .ZN(n4236) );
  NAND2_X1 U3855 ( .A1(n3212), .A2(n3287), .ZN(n3286) );
  NAND2_X1 U3856 ( .A1(n4289), .A2(n3447), .ZN(n3877) );
  OR2_X1 U3857 ( .A1(n3591), .A2(n3590), .ZN(n3655) );
  XNOR2_X1 U3858 ( .A(n3505), .B(n3504), .ZN(n3971) );
  INV_X1 U3859 ( .A(n3503), .ZN(n3504) );
  AOI21_X1 U3860 ( .B1(n3452), .B2(n4289), .A(n4149), .ZN(n3440) );
  NAND2_X1 U3861 ( .A1(n3365), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U3862 ( .A1(n3488), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3387), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3369) );
  AOI21_X1 U3863 ( .B1(n3387), .B2(INSTQUEUE_REG_14__3__SCAN_IN), .A(n3376), 
        .ZN(n3379) );
  AND2_X1 U3864 ( .A1(n3519), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U3865 ( .A1(n5438), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3524), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U3866 ( .A1(n3519), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3332) );
  INV_X1 U3867 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7005) );
  INV_X1 U3868 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7010) );
  NAND2_X1 U3869 ( .A1(n3998), .A2(n3988), .ZN(n6507) );
  AND2_X1 U3870 ( .A1(n6504), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3998) );
  NAND2_X1 U3871 ( .A1(n5029), .A2(n4144), .ZN(n4155) );
  NAND2_X1 U3872 ( .A1(n5951), .A2(n5940), .ZN(n5939) );
  AND2_X1 U3873 ( .A1(n5428), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5449)
         );
  NAND2_X1 U3874 ( .A1(n5449), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5472)
         );
  AND2_X1 U3875 ( .A1(n5409), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5428)
         );
  OR3_X1 U3876 ( .A1(n5364), .A2(n5977), .A3(n6124), .ZN(n5388) );
  NAND2_X1 U3877 ( .A1(n6003), .A2(n3247), .ZN(n5963) );
  NAND2_X1 U3878 ( .A1(n6003), .A2(n3249), .ZN(n5986) );
  AND2_X1 U3879 ( .A1(n5321), .A2(n5320), .ZN(n6002) );
  NAND2_X1 U3880 ( .A1(n6003), .A2(n6002), .ZN(n6005) );
  INV_X1 U3881 ( .A(n5239), .ZN(n3242) );
  NAND2_X1 U3882 ( .A1(n5179), .A2(n3243), .ZN(n5240) );
  AND2_X1 U3883 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  NAND2_X1 U3884 ( .A1(n5179), .A2(n5178), .ZN(n5203) );
  NAND2_X1 U3885 ( .A1(n4981), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5136)
         );
  NAND2_X1 U3886 ( .A1(n4642), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4717)
         );
  NOR2_X1 U3887 ( .A1(n4717), .A2(n5820), .ZN(n4981) );
  AND2_X1 U3888 ( .A1(n4736), .A2(n3253), .ZN(n3252) );
  INV_X1 U3889 ( .A(n3254), .ZN(n3253) );
  AND2_X1 U3890 ( .A1(n4737), .A2(n4735), .ZN(n4736) );
  AND2_X1 U3891 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n4656), .ZN(n4642)
         );
  AND2_X1 U3892 ( .A1(n4900), .A2(n4899), .ZN(n5046) );
  AND2_X1 U3893 ( .A1(n4687), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4671)
         );
  AND2_X1 U3894 ( .A1(n4702), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4687)
         );
  AND3_X1 U3895 ( .A1(n4575), .A2(n4574), .A3(n4573), .ZN(n4577) );
  NOR2_X1 U3896 ( .A1(n4506), .A2(n3254), .ZN(n4898) );
  NAND2_X1 U3897 ( .A1(n3251), .A2(n4504), .ZN(n4576) );
  NAND2_X1 U3898 ( .A1(n4419), .A2(n4418), .ZN(n4502) );
  NOR2_X1 U3899 ( .A1(n4320), .A2(n4319), .ZN(n4414) );
  NAND2_X1 U3900 ( .A1(n4237), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4320)
         );
  NOR2_X1 U3901 ( .A1(n4219), .A2(n5013), .ZN(n4237) );
  INV_X1 U3902 ( .A(n4125), .ZN(n4209) );
  NAND2_X1 U3903 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4125) );
  AOI21_X1 U3904 ( .B1(n4154), .B2(n4153), .A(n3633), .ZN(n6697) );
  INV_X1 U3905 ( .A(n5300), .ZN(n3277) );
  NAND2_X1 U3906 ( .A1(n6262), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3275) );
  OR3_X1 U3907 ( .A1(n5294), .A2(n3200), .A3(n5999), .ZN(n3258) );
  NOR3_X1 U3908 ( .A1(n5242), .A2(n5294), .A3(n3200), .ZN(n6010) );
  NAND2_X1 U3909 ( .A1(n6139), .A2(n6138), .ZN(n6130) );
  NOR3_X1 U3910 ( .A1(n5242), .A2(n5294), .A3(n3894), .ZN(n6008) );
  INV_X1 U3911 ( .A(n3234), .ZN(n3233) );
  NAND2_X1 U3912 ( .A1(n3873), .A2(n3270), .ZN(n3267) );
  INV_X1 U3913 ( .A(n4740), .ZN(n3270) );
  NOR3_X1 U3914 ( .A1(n4956), .A2(n3271), .A3(n4957), .ZN(n5055) );
  NOR2_X1 U3915 ( .A1(n5023), .A2(n3947), .ZN(n5262) );
  INV_X1 U3916 ( .A(n3728), .ZN(n3216) );
  INV_X1 U3917 ( .A(n3218), .ZN(n3217) );
  NOR2_X1 U3918 ( .A1(n4956), .A2(n4957), .ZN(n5053) );
  NAND2_X1 U3919 ( .A1(n4589), .A2(n4588), .ZN(n4895) );
  NAND2_X1 U3920 ( .A1(n4743), .A2(n3728), .ZN(n5018) );
  NAND2_X1 U3921 ( .A1(n5018), .A2(n5019), .ZN(n5094) );
  INV_X1 U3922 ( .A(n4315), .ZN(n3256) );
  INV_X1 U3923 ( .A(n4316), .ZN(n3257) );
  NOR2_X1 U3924 ( .A1(n4250), .A2(n4206), .ZN(n4234) );
  NAND2_X1 U3925 ( .A1(n3266), .A2(n3265), .ZN(n4250) );
  NOR2_X1 U3926 ( .A1(n4247), .A2(n4248), .ZN(n3265) );
  INV_X1 U3927 ( .A(n4249), .ZN(n3266) );
  OR2_X1 U3928 ( .A1(n3945), .A2(n4061), .ZN(n6795) );
  INV_X1 U3929 ( .A(n3939), .ZN(n3477) );
  AND3_X1 U3930 ( .A1(n3544), .A2(n3543), .A3(n3542), .ZN(n3609) );
  INV_X1 U3931 ( .A(n3600), .ZN(n3237) );
  AND2_X1 U3933 ( .A1(n4265), .A2(n6923), .ZN(n6811) );
  AND2_X1 U3934 ( .A1(n4208), .A2(n6284), .ZN(n4838) );
  AND2_X1 U3935 ( .A1(n6281), .A2(n4060), .ZN(n4842) );
  INV_X1 U3936 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6930) );
  INV_X1 U3937 ( .A(n6817), .ZN(n4836) );
  NAND2_X1 U3938 ( .A1(n3281), .A2(n4841), .ZN(n3280) );
  NAND2_X1 U3939 ( .A1(n3283), .A2(n3576), .ZN(n3282) );
  AND2_X1 U3940 ( .A1(n4269), .A2(n4268), .ZN(n4295) );
  AND2_X1 U3941 ( .A1(n3807), .A2(n3806), .ZN(n4040) );
  OAI21_X1 U3942 ( .B1(n3805), .B2(n3804), .A(n3803), .ZN(n3806) );
  AND2_X1 U3943 ( .A1(n3983), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3822) );
  AND2_X1 U3944 ( .A1(n6504), .A2(n3999), .ZN(n6518) );
  INV_X1 U3945 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U3946 ( .A1(n3550), .A2(n3551), .ZN(n3487) );
  INV_X1 U3947 ( .A(n6543), .ZN(n6522) );
  INV_X1 U3948 ( .A(n6539), .ZN(n6527) );
  INV_X1 U3949 ( .A(n3261), .ZN(n6304) );
  OR2_X1 U3950 ( .A1(n4141), .A2(n7033), .ZN(n4148) );
  AND2_X1 U3951 ( .A1(n6064), .A2(n4344), .ZN(n6562) );
  AND2_X1 U3952 ( .A1(n6064), .A2(n4343), .ZN(n6559) );
  INV_X1 U3953 ( .A(n6064), .ZN(n6561) );
  OR2_X1 U3954 ( .A1(n6558), .A2(n6562), .ZN(n5004) );
  INV_X1 U3955 ( .A(n5004), .ZN(n5048) );
  INV_X1 U3956 ( .A(n6559), .ZN(n6345) );
  CLKBUF_X1 U3957 ( .A(n6578), .Z(n7160) );
  NAND2_X1 U3958 ( .A1(n4340), .A2(n4093), .ZN(n6660) );
  NOR2_X1 U3959 ( .A1(n3197), .A2(n5909), .ZN(n3223) );
  AND2_X1 U3960 ( .A1(n3197), .A2(n5909), .ZN(n3224) );
  INV_X1 U3961 ( .A(n6155), .ZN(n6350) );
  NAND2_X1 U3962 ( .A1(n6681), .A2(n4081), .ZN(n6162) );
  INV_X1 U3963 ( .A(n6704), .ZN(n6663) );
  INV_X1 U3964 ( .A(n6162), .ZN(n6694) );
  INV_X1 U3965 ( .A(n3263), .ZN(n5533) );
  INV_X1 U3966 ( .A(n3740), .ZN(n6089) );
  AND2_X1 U3967 ( .A1(n6197), .A2(n6199), .ZN(n6188) );
  NAND2_X1 U3968 ( .A1(n3230), .A2(n5247), .ZN(n6172) );
  NAND2_X1 U3969 ( .A1(n3190), .A2(n5248), .ZN(n3230) );
  NOR2_X1 U3970 ( .A1(n3945), .A2(n4182), .ZN(n5258) );
  INV_X1 U3971 ( .A(n6773), .ZN(n6801) );
  INV_X1 U3972 ( .A(n7026), .ZN(n6297) );
  CLKBUF_X1 U3973 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n6301) );
  NAND2_X1 U3974 ( .A1(n3278), .A2(n3576), .ZN(n4195) );
  INV_X1 U3975 ( .A(n3575), .ZN(n3278) );
  OR3_X1 U3976 ( .A1(n6863), .A2(n6862), .A3(n6861), .ZN(n6890) );
  INV_X1 U3977 ( .A(n6856), .ZN(n6888) );
  INV_X1 U3978 ( .A(n4802), .ZN(n6939) );
  INV_X1 U3979 ( .A(n4816), .ZN(n6945) );
  INV_X1 U3980 ( .A(n4828), .ZN(n6951) );
  INV_X1 U3981 ( .A(n4832), .ZN(n6957) );
  INV_X1 U3982 ( .A(n4905), .ZN(n6970) );
  AND2_X1 U3983 ( .A1(n4425), .A2(n6817), .ZN(n4885) );
  INV_X1 U3984 ( .A(n4824), .ZN(n6979) );
  INV_X1 U3985 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7028) );
  NOR2_X1 U3986 ( .A1(n3454), .A2(n4040), .ZN(n7026) );
  OAI21_X1 U3987 ( .B1(n6088), .B2(n6681), .A(n3239), .ZN(U2957) );
  INV_X1 U3988 ( .A(n3240), .ZN(n3239) );
  OAI21_X1 U3989 ( .B1(n6085), .B2(n6679), .A(n3241), .ZN(n3240) );
  AOI21_X1 U3990 ( .B1(n6663), .B2(n6087), .A(n6086), .ZN(n3241) );
  INV_X1 U3991 ( .A(n3260), .ZN(n5545) );
  INV_X2 U3992 ( .A(n6131), .ZN(n6262) );
  NAND2_X2 U3993 ( .A1(n3917), .A2(n3913), .ZN(n3852) );
  AND2_X2 U3994 ( .A1(n3317), .A2(n4172), .ZN(n3387) );
  NAND2_X1 U3995 ( .A1(n3518), .A2(n4279), .ZN(n3766) );
  NOR2_X1 U3996 ( .A1(n5563), .A2(n5562), .ZN(n3197) );
  AND2_X1 U3997 ( .A1(n6138), .A2(n3207), .ZN(n3198) );
  AND2_X2 U3998 ( .A1(n4039), .A2(n4172), .ZN(n3524) );
  NOR2_X1 U3999 ( .A1(n5541), .A2(n6079), .ZN(n3199) );
  OR2_X1 U4000 ( .A1(n3894), .A2(n3259), .ZN(n3200) );
  OR3_X1 U4001 ( .A1(n4956), .A2(n3268), .A3(n3267), .ZN(n3201) );
  OAI21_X1 U4002 ( .B1(n4294), .B2(n3452), .A(n3364), .ZN(n3458) );
  CLKBUF_X3 U4003 ( .A(n3877), .Z(n3913) );
  NAND2_X1 U4004 ( .A1(n3453), .A2(n3290), .ZN(n3554) );
  XOR2_X1 U4005 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .B(n5302), .Z(n3202) );
  INV_X1 U4006 ( .A(n3435), .ZN(n3518) );
  NOR2_X1 U4007 ( .A1(n4289), .A2(n3439), .ZN(n3476) );
  NOR2_X1 U4008 ( .A1(n3447), .A2(n3741), .ZN(n3475) );
  AND2_X1 U4009 ( .A1(n6263), .A2(n5841), .ZN(n3203) );
  NOR2_X1 U4010 ( .A1(n6263), .A2(n3732), .ZN(n3204) );
  NAND2_X1 U4011 ( .A1(n5093), .A2(n5096), .ZN(n3205) );
  AND2_X1 U4012 ( .A1(n3730), .A2(n3729), .ZN(n3206) );
  INV_X1 U4013 ( .A(n6775), .ZN(n6799) );
  NAND2_X1 U4014 ( .A1(n3284), .A2(n3729), .ZN(n5215) );
  NOR2_X1 U4015 ( .A1(n6262), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3207)
         );
  AND2_X1 U4016 ( .A1(n6131), .A2(n3286), .ZN(n3208) );
  NAND2_X1 U4017 ( .A1(n4503), .A2(n4502), .ZN(n4506) );
  NAND2_X1 U4018 ( .A1(n4279), .A2(n3447), .ZN(n3762) );
  INV_X1 U4019 ( .A(n3762), .ZN(n3794) );
  OR2_X1 U4020 ( .A1(n5242), .A2(n3894), .ZN(n3209) );
  AND2_X1 U4021 ( .A1(n3242), .A2(n3243), .ZN(n3210) );
  INV_X1 U4022 ( .A(n4841), .ZN(n3283) );
  INV_X1 U4023 ( .A(n3439), .ZN(n3809) );
  OR3_X1 U4024 ( .A1(n4956), .A2(n3268), .A3(n3271), .ZN(n3211) );
  NAND2_X1 U4025 ( .A1(n3446), .A2(n3434), .ZN(n4142) );
  AND3_X1 U4026 ( .A1(n6232), .A2(n6122), .A3(n6216), .ZN(n3212) );
  INV_X1 U4027 ( .A(n5909), .ZN(n3229) );
  AND2_X1 U4028 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4172) );
  NOR2_X2 U4029 ( .A1(n6679), .A2(n5896), .ZN(n6968) );
  OR2_X1 U4030 ( .A1(n7044), .A2(n6927), .ZN(n6679) );
  OAI21_X1 U4031 ( .B1(n4743), .B2(n3217), .A(n3215), .ZN(n5105) );
  NAND2_X1 U4032 ( .A1(n4743), .A2(n3215), .ZN(n3214) );
  AOI21_X2 U4033 ( .B1(n3218), .B2(n3216), .A(n3205), .ZN(n3215) );
  OR2_X1 U4034 ( .A1(n5558), .A2(n5557), .ZN(n3220) );
  NOR2_X1 U4035 ( .A1(n3220), .A2(n5552), .ZN(n6221) );
  OAI211_X1 U4036 ( .C1(n3225), .C2(n3227), .A(n3222), .B(n3221), .ZN(U2962)
         );
  NAND2_X1 U4037 ( .A1(n3227), .A2(n3224), .ZN(n3221) );
  AOI21_X1 U4038 ( .B1(n5552), .B2(n3224), .A(n3223), .ZN(n3222) );
  NAND2_X1 U4039 ( .A1(n3226), .A2(n3229), .ZN(n3225) );
  INV_X1 U4040 ( .A(n5552), .ZN(n3226) );
  NAND2_X1 U4041 ( .A1(n3236), .A2(n3607), .ZN(n6695) );
  NAND3_X1 U4042 ( .A1(n3641), .A2(n3794), .A3(n3602), .ZN(n3236) );
  INV_X1 U4043 ( .A(n3601), .ZN(n3238) );
  AND2_X2 U4044 ( .A1(n6003), .A2(n3245), .ZN(n6044) );
  INV_X1 U4045 ( .A(n4506), .ZN(n3251) );
  NAND2_X1 U4046 ( .A1(n3251), .A2(n3252), .ZN(n4986) );
  NAND4_X1 U4047 ( .A1(n6308), .A2(n6307), .A3(n6309), .A4(n6310), .ZN(U2797)
         );
  NOR2_X2 U4048 ( .A1(n4447), .A2(n4446), .ZN(n4509) );
  OR2_X2 U4049 ( .A1(n5242), .A2(n3258), .ZN(n5996) );
  INV_X1 U4050 ( .A(n6007), .ZN(n3259) );
  OAI211_X1 U4051 ( .C1(n5535), .C2(n5945), .A(n5536), .B(n3263), .ZN(n3262)
         );
  INV_X1 U4052 ( .A(n3873), .ZN(n3271) );
  INV_X1 U4053 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3272) );
  AND2_X2 U4054 ( .A1(n4174), .A2(n3317), .ZN(n3489) );
  AND2_X2 U4055 ( .A1(n3272), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3317)
         );
  NOR2_X4 U4056 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4174) );
  NAND2_X1 U4057 ( .A1(n3575), .A2(n4841), .ZN(n3279) );
  OAI211_X2 U4058 ( .C1(n3575), .C2(n3282), .A(n3280), .B(n3279), .ZN(n4173)
         );
  OR2_X1 U4059 ( .A1(n6264), .A2(n3285), .ZN(n3734) );
  NAND3_X1 U4060 ( .A1(n6381), .A2(n6391), .A3(n6374), .ZN(n3285) );
  NOR2_X1 U4061 ( .A1(n6146), .A2(n3738), .ZN(n5550) );
  OAI22_X2 U4062 ( .A1(n6146), .A2(n3208), .B1(n6131), .B2(n3737), .ZN(n6090)
         );
  XNOR2_X1 U4063 ( .A(n3289), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6088)
         );
  AOI21_X1 U4064 ( .B1(n6121), .B2(n6122), .A(n5555), .ZN(n5558) );
  INV_X1 U4065 ( .A(n3641), .ZN(n3642) );
  XNOR2_X1 U4066 ( .A(n3611), .B(n3610), .ZN(n3612) );
  NAND2_X1 U4067 ( .A1(n6668), .A2(n6670), .ZN(n6669) );
  CLKBUF_X1 U4068 ( .A(n6090), .Z(n6116) );
  AOI22_X1 U4069 ( .A1(n3365), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3380) );
  NAND2_X1 U4070 ( .A1(n7028), .A2(n4268), .ZN(n4600) );
  AND2_X1 U4071 ( .A1(n3968), .A2(n3967), .ZN(n3288) );
  OR2_X1 U4072 ( .A1(n5531), .A2(n5532), .ZN(n3289) );
  OR2_X1 U4073 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5499) );
  AND4_X1 U4074 ( .A1(n3374), .A2(n3373), .A3(n3372), .A4(n3371), .ZN(n3291)
         );
  INV_X1 U4075 ( .A(n3534), .ZN(n3621) );
  NOR2_X1 U4076 ( .A1(n4060), .A2(n4027), .ZN(n3293) );
  AND3_X1 U4077 ( .A1(n3362), .A2(n3361), .A3(n3360), .ZN(n3294) );
  INV_X1 U4078 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4319) );
  INV_X1 U4079 ( .A(n3444), .ZN(n4149) );
  AND2_X1 U4080 ( .A1(n4148), .A2(n4147), .ZN(n6055) );
  AND2_X1 U4081 ( .A1(n3184), .A2(n3444), .ZN(n3295) );
  OR2_X1 U4082 ( .A1(n3766), .A2(n4097), .ZN(n3296) );
  AND2_X1 U4083 ( .A1(n6504), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6525) );
  AND2_X1 U4084 ( .A1(n3465), .A2(n3432), .ZN(n3433) );
  AND2_X1 U4085 ( .A1(n3771), .A2(n3770), .ZN(n3775) );
  INV_X1 U4086 ( .A(n3766), .ZN(n3466) );
  INV_X1 U4087 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3743) );
  OR2_X1 U4088 ( .A1(n3674), .A2(n3673), .ZN(n3697) );
  AND3_X1 U4089 ( .A1(n3307), .A2(n3306), .A3(n3305), .ZN(n3308) );
  AOI22_X1 U4090 ( .A1(n3421), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3526), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3330) );
  INV_X1 U4091 ( .A(n3767), .ZN(n3744) );
  OR2_X1 U4092 ( .A1(n3653), .A2(n3652), .ZN(n3698) );
  INV_X1 U4093 ( .A(n5467), .ZN(n5503) );
  INV_X1 U4094 ( .A(n5510), .ZN(n5369) );
  XNOR2_X1 U4095 ( .A(n3706), .B(n3707), .ZN(n4318) );
  OR2_X1 U4096 ( .A1(n5554), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5555)
         );
  INV_X1 U4097 ( .A(n3781), .ZN(n3804) );
  NAND2_X1 U4098 ( .A1(n3447), .A2(n3473), .ZN(n3465) );
  NAND2_X1 U4099 ( .A1(n3560), .A2(n3559), .ZN(n3576) );
  AND2_X1 U4100 ( .A1(n3862), .A2(n3861), .ZN(n4588) );
  NOR2_X1 U4101 ( .A1(n4970), .A2(n7028), .ZN(n5467) );
  NOR2_X1 U4102 ( .A1(n5285), .A2(n6140), .ZN(n5318) );
  AND2_X1 U4103 ( .A1(n4671), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4656)
         );
  INV_X1 U4104 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4487) );
  OR4_X1 U4105 ( .A1(n6262), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A4(INSTADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n5300) );
  AND2_X1 U4106 ( .A1(n6120), .A2(n5556), .ZN(n5557) );
  INV_X1 U4107 ( .A(n5216), .ZN(n3730) );
  AND2_X1 U4108 ( .A1(n4917), .A2(n6923), .ZN(n4919) );
  OAI21_X1 U4109 ( .B1(n7163), .B2(n4171), .A(n6297), .ZN(n4268) );
  INV_X1 U4110 ( .A(n5198), .ZN(n3981) );
  NOR2_X1 U4111 ( .A1(n4486), .A2(n4487), .ZN(n4562) );
  INV_X1 U4112 ( .A(n6507), .ZN(n6532) );
  AND2_X1 U4113 ( .A1(n4716), .A2(n4897), .ZN(n4735) );
  OR2_X1 U4114 ( .A1(n5472), .A2(n6084), .ZN(n5505) );
  NOR2_X1 U4115 ( .A1(n5388), .A2(n6111), .ZN(n5409) );
  AND2_X1 U4116 ( .A1(n4562), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4702)
         );
  OR2_X1 U4117 ( .A1(n7147), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4080) );
  OR2_X1 U4118 ( .A1(n3945), .A2(n3929), .ZN(n6775) );
  NAND2_X1 U4119 ( .A1(n3580), .A2(n3579), .ZN(n4841) );
  INV_X1 U4120 ( .A(n3196), .ZN(n4751) );
  NOR2_X1 U4121 ( .A1(n6284), .A2(n4377), .ZN(n4804) );
  INV_X1 U4122 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7016) );
  NAND2_X1 U4123 ( .A1(n5236), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5285)
         );
  AND2_X1 U4124 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n3981), .ZN(n5236)
         );
  AND2_X1 U4125 ( .A1(n3995), .A2(n3993), .ZN(n6539) );
  INV_X1 U4126 ( .A(n6511), .ZN(n6524) );
  AND2_X1 U4127 ( .A1(n3998), .A2(n3997), .ZN(n6543) );
  INV_X1 U4128 ( .A(n6660), .ZN(n6653) );
  NAND2_X1 U4129 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n4209), .ZN(n4219)
         );
  INV_X1 U4130 ( .A(n6681), .ZN(n6700) );
  OR2_X1 U4131 ( .A1(n5258), .A2(n5263), .ZN(n6743) );
  INV_X1 U4132 ( .A(n6774), .ZN(n6803) );
  NAND2_X1 U4133 ( .A1(n3823), .A2(n7036), .ZN(n3945) );
  INV_X1 U4134 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n3983) );
  AND2_X1 U4135 ( .A1(n4528), .A2(n6294), .ZN(n5085) );
  INV_X1 U4136 ( .A(n4554), .ZN(n4298) );
  INV_X1 U4137 ( .A(n6822), .ZN(n6846) );
  INV_X1 U4138 ( .A(n6923), .ZN(n6927) );
  OR2_X1 U4139 ( .A1(n4605), .A2(n4604), .ZN(n4629) );
  AND2_X1 U4140 ( .A1(n4838), .A2(n4751), .ZN(n4351) );
  INV_X1 U4141 ( .A(n4450), .ZN(n4482) );
  AND2_X1 U4142 ( .A1(n3196), .A2(n6817), .ZN(n4527) );
  INV_X1 U4143 ( .A(n6974), .ZN(n6976) );
  INV_X1 U4144 ( .A(n4812), .ZN(n6920) );
  INV_X1 U4145 ( .A(n4820), .ZN(n6963) );
  AND2_X1 U4146 ( .A1(n4804), .A2(n4751), .ZN(n4425) );
  AND2_X1 U4147 ( .A1(n4804), .A2(n4527), .ZN(n4909) );
  NAND2_X1 U4148 ( .A1(n4340), .A2(n4009), .ZN(n6598) );
  AND2_X1 U4149 ( .A1(n6598), .A2(n4006), .ZN(n7157) );
  NAND2_X1 U4150 ( .A1(n6504), .A2(n3984), .ZN(n6515) );
  OR2_X1 U4151 ( .A1(n5047), .A2(n5046), .ZN(n6458) );
  NAND3_X1 U4152 ( .A1(n4342), .A2(n4341), .A3(n6656), .ZN(n6064) );
  INV_X1 U4153 ( .A(n6590), .ZN(n6596) );
  NAND2_X1 U4154 ( .A1(n4340), .A2(n4077), .ZN(n6681) );
  NAND2_X1 U4155 ( .A1(n6162), .A2(n4228), .ZN(n6704) );
  INV_X1 U4156 ( .A(n6785), .ZN(n6774) );
  OR2_X1 U4157 ( .A1(n3945), .A2(n3829), .ZN(n6773) );
  AND2_X1 U4158 ( .A1(n4759), .A2(n4758), .ZN(n4795) );
  NAND2_X1 U4159 ( .A1(n4753), .A2(n6817), .ZN(n4944) );
  INV_X1 U4160 ( .A(n5061), .ZN(n5092) );
  NAND2_X1 U4161 ( .A1(n6291), .A2(n4527), .ZN(n6917) );
  NAND2_X1 U4162 ( .A1(n4351), .A2(n6817), .ZN(n4632) );
  NAND2_X1 U4163 ( .A1(n4838), .A2(n4527), .ZN(n6985) );
  NOR2_X1 U4164 ( .A1(n4846), .A2(n4845), .ZN(n4893) );
  NAND2_X1 U4165 ( .A1(n4425), .A2(n4836), .ZN(n4445) );
  AND2_X1 U4166 ( .A1(n7025), .A2(n7024), .ZN(n7042) );
  OAI21_X1 U4167 ( .B1(n6088), .B2(n6773), .A(n3288), .ZN(U2989) );
  INV_X1 U4168 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3297) );
  AND2_X2 U4169 ( .A1(n3297), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3311)
         );
  NAND2_X1 U4170 ( .A1(n3488), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3300) );
  AND2_X2 U4171 ( .A1(n3298), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3312)
         );
  AND2_X2 U4172 ( .A1(n4039), .A2(n3312), .ZN(n3519) );
  NAND2_X1 U4173 ( .A1(n3519), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3299) );
  NAND2_X1 U4174 ( .A1(n3300), .A2(n3299), .ZN(n3304) );
  AND2_X4 U4175 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4032) );
  NAND2_X1 U4176 ( .A1(n3494), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3302) );
  NAND2_X1 U4177 ( .A1(n3387), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3301)
         );
  NAND2_X1 U4178 ( .A1(n3302), .A2(n3301), .ZN(n3303) );
  NOR2_X1 U4179 ( .A1(n3304), .A2(n3303), .ZN(n3310) );
  NOR2_X4 U4180 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4033) );
  AND2_X2 U4181 ( .A1(n4033), .A2(n4174), .ZN(n3421) );
  NAND2_X1 U4182 ( .A1(n3421), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3309) );
  NAND2_X1 U4183 ( .A1(n3526), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3306)
         );
  NAND2_X1 U4184 ( .A1(n3400), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3305) );
  AND2_X4 U4185 ( .A1(n3311), .A2(n4032), .ZN(n3643) );
  NAND2_X1 U4186 ( .A1(n3643), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3316)
         );
  AND2_X2 U4187 ( .A1(n3312), .A2(n4033), .ZN(n3506) );
  NAND2_X1 U4188 ( .A1(n3506), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U4189 ( .A1(n3365), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3314) );
  AND2_X2 U4190 ( .A1(n3312), .A2(n4032), .ZN(n3370) );
  AND2_X4 U4191 ( .A1(n4174), .A2(n4039), .ZN(n5438) );
  NAND2_X1 U4192 ( .A1(n3524), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3320)
         );
  NAND2_X1 U4193 ( .A1(n3489), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4194 ( .A1(n3511), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3318)
         );
  AOI22_X1 U4195 ( .A1(n3489), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3511), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4196 ( .A1(n3365), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4197 ( .A1(n3488), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3387), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4198 ( .A1(n5398), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4199 ( .A1(n3643), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3329) );
  NAND2_X1 U4200 ( .A1(n5438), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U4201 ( .A1(n3524), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3337)
         );
  NAND2_X1 U4202 ( .A1(n3489), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3336) );
  NAND2_X1 U4203 ( .A1(n3511), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3335)
         );
  NAND2_X1 U4204 ( .A1(n3643), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3342)
         );
  NAND2_X1 U4205 ( .A1(n3506), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3341) );
  NAND2_X1 U4206 ( .A1(n3365), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U4207 ( .A1(n3370), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4208 ( .A1(n3488), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3346) );
  NAND2_X1 U4209 ( .A1(n3519), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3345) );
  NAND2_X1 U4210 ( .A1(n3387), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3344)
         );
  NAND2_X1 U4211 ( .A1(n3494), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4212 ( .A1(n5398), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3350)
         );
  NAND2_X1 U4213 ( .A1(n3400), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3349) );
  NAND2_X1 U4214 ( .A1(n3421), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3348) );
  NAND2_X1 U4215 ( .A1(n3526), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3347)
         );
  AND4_X2 U4216 ( .A1(n3354), .A2(n3353), .A3(n3352), .A4(n3351), .ZN(n3446)
         );
  AOI22_X1 U4217 ( .A1(n3524), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4218 ( .A1(n5398), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4219 ( .A1(n5438), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3511), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4220 ( .A1(n3421), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3526), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4221 ( .A1(n3643), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4222 ( .A1(n3488), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4223 ( .A1(n3519), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3387), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4224 ( .A1(n3365), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4225 ( .A1(n3400), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3511), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4226 ( .A1(n3421), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3526), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4227 ( .A1(n3506), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4228 ( .A1(n5438), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4229 ( .A1(n5398), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3524), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4230 ( .A1(n3519), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3371) );
  NAND2_X1 U4231 ( .A1(n3375), .A2(n3291), .ZN(n3439) );
  AOI22_X1 U4232 ( .A1(n3488), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4233 ( .A1(n5333), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3377) );
  NAND4_X1 U4234 ( .A1(n3380), .A2(n3379), .A3(n3378), .A4(n3377), .ZN(n3386)
         );
  AOI22_X1 U4235 ( .A1(n5438), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3511), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4236 ( .A1(n5398), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4237 ( .A1(n3524), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4238 ( .A1(n3421), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3526), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3381) );
  NAND4_X1 U4239 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3385)
         );
  OR2_X2 U4240 ( .A1(n3386), .A2(n3385), .ZN(n4289) );
  NAND2_X1 U4241 ( .A1(n3488), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4242 ( .A1(n3519), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4243 ( .A1(n3387), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3389)
         );
  NAND2_X1 U4244 ( .A1(n3494), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3388) );
  NAND2_X1 U4245 ( .A1(n5333), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3395)
         );
  NAND2_X1 U4246 ( .A1(n3506), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U4247 ( .A1(n3365), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U4248 ( .A1(n3370), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3392) );
  AND4_X2 U4249 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3407)
         );
  NAND2_X1 U4250 ( .A1(n5438), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3398) );
  NAND2_X1 U4251 ( .A1(n3511), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3397)
         );
  NAND2_X1 U4252 ( .A1(n3524), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3396)
         );
  NAND3_X1 U4253 ( .A1(n3398), .A2(n3397), .A3(n3396), .ZN(n3399) );
  AOI21_X2 U4254 ( .B1(n3489), .B2(INSTQUEUE_REG_2__1__SCAN_IN), .A(n3399), 
        .ZN(n3406) );
  NAND2_X1 U4255 ( .A1(n5398), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3404)
         );
  NAND2_X1 U4256 ( .A1(n3400), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3403) );
  NAND2_X1 U4257 ( .A1(n3421), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3402) );
  NAND2_X1 U4258 ( .A1(n3526), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3401)
         );
  NAND4_X4 U4259 ( .A1(n3408), .A2(n3407), .A3(n3406), .A4(n3405), .ZN(n3447)
         );
  NAND2_X1 U4260 ( .A1(n3519), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3412) );
  NAND2_X1 U4261 ( .A1(n3488), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3411) );
  NAND2_X1 U4262 ( .A1(n3643), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3410)
         );
  NAND2_X1 U4263 ( .A1(n3506), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3409) );
  NAND2_X1 U4264 ( .A1(n3387), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3416)
         );
  NAND2_X1 U4265 ( .A1(n5438), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3415) );
  NAND2_X1 U4266 ( .A1(n3370), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3414) );
  NAND2_X1 U4267 ( .A1(n3494), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3413) );
  NAND2_X1 U4268 ( .A1(n3489), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3420) );
  NAND2_X1 U4269 ( .A1(n5398), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3419)
         );
  NAND2_X1 U4270 ( .A1(n3400), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U4271 ( .A1(n3511), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3417)
         );
  NAND2_X1 U4272 ( .A1(n3526), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3424)
         );
  NAND2_X1 U4273 ( .A1(n3421), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3423) );
  NAND2_X1 U4274 ( .A1(n3524), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3422)
         );
  NAND4_X4 U4275 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n4097)
         );
  INV_X1 U4276 ( .A(STATE_REG_1__SCAN_IN), .ZN(n7055) );
  XNOR2_X1 U4277 ( .A(n7055), .B(STATE_REG_2__SCAN_IN), .ZN(n3741) );
  INV_X1 U4278 ( .A(n3475), .ZN(n3431) );
  NAND2_X1 U4279 ( .A1(n3431), .A2(n3430), .ZN(n3432) );
  NAND2_X1 U4280 ( .A1(n3969), .A2(n3443), .ZN(n3438) );
  NAND2_X1 U4281 ( .A1(n4142), .A2(n3809), .ZN(n3436) );
  NAND2_X1 U4282 ( .A1(n3436), .A2(n3184), .ZN(n3437) );
  NAND2_X1 U4283 ( .A1(n3443), .A2(n3439), .ZN(n3441) );
  NAND2_X1 U4284 ( .A1(n3478), .A2(n3826), .ZN(n3468) );
  INV_X1 U4285 ( .A(n3443), .ZN(n3445) );
  INV_X2 U4286 ( .A(n3447), .ZN(n3479) );
  NAND2_X1 U4287 ( .A1(n3471), .A2(n3596), .ZN(n3449) );
  INV_X1 U4288 ( .A(n3877), .ZN(n3448) );
  NAND2_X1 U4289 ( .A1(n3466), .A2(n3448), .ZN(n3940) );
  NAND3_X1 U4290 ( .A1(n3450), .A2(n3468), .A3(n3464), .ZN(n3451) );
  NAND2_X1 U4291 ( .A1(n3451), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3453) );
  INV_X1 U4292 ( .A(n3822), .ZN(n4143) );
  INV_X1 U4293 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n3454) );
  NAND2_X1 U4294 ( .A1(n3454), .A2(n3983), .ZN(n7147) );
  INV_X1 U4295 ( .A(n4080), .ZN(n3558) );
  MUX2_X1 U4296 ( .A(n4143), .B(n3558), .S(n7000), .Z(n3455) );
  INV_X1 U4297 ( .A(n3455), .ZN(n3456) );
  OR2_X1 U4298 ( .A1(n7147), .A2(n7028), .ZN(n7035) );
  AOI21_X1 U4299 ( .B1(n3932), .B2(n4097), .A(n7035), .ZN(n3463) );
  NAND2_X1 U4300 ( .A1(n3476), .A2(n3969), .ZN(n3462) );
  NAND2_X1 U4301 ( .A1(n3452), .A2(n4294), .ZN(n3459) );
  NAND2_X1 U4302 ( .A1(n3459), .A2(n4289), .ZN(n3460) );
  OAI21_X1 U4303 ( .B1(n3466), .B2(n3465), .A(n3818), .ZN(n3467) );
  INV_X1 U4304 ( .A(n3467), .ZN(n3469) );
  INV_X1 U4305 ( .A(n3471), .ZN(n3817) );
  NOR2_X1 U4306 ( .A1(n3932), .A2(n4279), .ZN(n3472) );
  NAND2_X1 U4307 ( .A1(n3817), .A2(n3472), .ZN(n3761) );
  INV_X1 U4308 ( .A(n3761), .ZN(n3474) );
  NAND2_X1 U4309 ( .A1(n3474), .A2(n4097), .ZN(n4016) );
  NAND3_X1 U4310 ( .A1(n3826), .A2(n3476), .A3(n3430), .ZN(n3939) );
  NAND2_X1 U4311 ( .A1(n3480), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3486) );
  INV_X1 U4312 ( .A(n3486), .ZN(n3482) );
  NAND2_X1 U4313 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3556) );
  OAI21_X1 U4314 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n3556), .ZN(n4595) );
  OAI22_X1 U4315 ( .A1(n4080), .A2(n4595), .B1(n3822), .B2(n7005), .ZN(n3483)
         );
  OR2_X1 U4316 ( .A1(n3483), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3481)
         );
  NAND2_X1 U4317 ( .A1(n3482), .A2(n3481), .ZN(n3550) );
  INV_X1 U4318 ( .A(n3483), .ZN(n3485) );
  NAND2_X1 U4319 ( .A1(n3554), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3484) );
  XNOR2_X2 U4320 ( .A(n3553), .B(n3487), .ZN(n4027) );
  NAND2_X1 U4321 ( .A1(n4027), .A2(n7028), .ZN(n3502) );
  INV_X1 U4322 ( .A(n3562), .ZN(n4333) );
  AOI22_X1 U4323 ( .A1(n5332), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4324 ( .A1(n5333), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4325 ( .A1(n3365), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4326 ( .A1(n5460), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3490) );
  NAND4_X1 U4327 ( .A1(n3493), .A2(n3492), .A3(n3491), .A4(n3490), .ZN(n3500)
         );
  AOI22_X1 U4328 ( .A1(n5486), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4329 ( .A1(n5478), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3497) );
  INV_X1 U4330 ( .A(n3511), .ZN(n3581) );
  AOI22_X1 U4331 ( .A1(n5487), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4332 ( .A1(n5475), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3495) );
  NAND4_X1 U4333 ( .A1(n3498), .A2(n3497), .A3(n3496), .A4(n3495), .ZN(n3499)
         );
  NAND2_X1 U4334 ( .A1(n4333), .A2(n3613), .ZN(n3501) );
  NAND2_X2 U4335 ( .A1(n3502), .A2(n3501), .ZN(n3611) );
  NAND2_X1 U4336 ( .A1(n3971), .A2(n7028), .ZN(n3619) );
  INV_X1 U4337 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5818) );
  AOI22_X1 U4338 ( .A1(n5485), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4339 ( .A1(n5333), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4340 ( .A1(n3365), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4341 ( .A1(n5332), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3507) );
  NAND4_X1 U4342 ( .A1(n3510), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(n3517)
         );
  AOI22_X1 U4343 ( .A1(n3525), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4344 ( .A1(n5486), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4345 ( .A1(n5460), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4346 ( .A1(n3421), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3512) );
  NAND4_X1 U4347 ( .A1(n3515), .A2(n3514), .A3(n3513), .A4(n3512), .ZN(n3516)
         );
  NOR2_X1 U4348 ( .A1(n3562), .A2(n3723), .ZN(n3540) );
  NAND2_X1 U4349 ( .A1(n3518), .A2(n3723), .ZN(n3535) );
  NOR2_X1 U4350 ( .A1(n3535), .A2(n7028), .ZN(n3538) );
  AOI22_X1 U4351 ( .A1(n5478), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4352 ( .A1(n5307), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5333), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3522) );
  BUF_X1 U4353 ( .A(n5438), .Z(n5460) );
  AOI22_X1 U4354 ( .A1(n5486), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5460), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4355 ( .A1(n3519), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3520) );
  NAND4_X1 U4356 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3532)
         );
  AOI22_X1 U4357 ( .A1(n5332), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4358 ( .A1(n3525), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4359 ( .A1(n3489), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4360 ( .A1(n3421), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3527) );
  NAND4_X1 U4361 ( .A1(n3530), .A2(n3529), .A3(n3528), .A4(n3527), .ZN(n3531)
         );
  INV_X1 U4362 ( .A(n3626), .ZN(n3533) );
  MUX2_X1 U4363 ( .A(n3540), .B(n3538), .S(n3533), .Z(n3534) );
  NAND2_X1 U4364 ( .A1(n3619), .A2(n3621), .ZN(n3537) );
  INV_X1 U4365 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4784) );
  AOI21_X1 U4366 ( .B1(n3473), .B2(n3626), .A(n7028), .ZN(n3536) );
  OAI211_X1 U4367 ( .C1(n3790), .C2(n4784), .A(n3536), .B(n3535), .ZN(n3622)
         );
  NAND2_X1 U4368 ( .A1(n3537), .A2(n3622), .ZN(n3539) );
  INV_X1 U4369 ( .A(n3538), .ZN(n3719) );
  NAND2_X1 U4370 ( .A1(n3539), .A2(n3719), .ZN(n3608) );
  NAND2_X1 U4371 ( .A1(n3611), .A2(n3608), .ZN(n3545) );
  INV_X1 U4372 ( .A(n3790), .ZN(n3800) );
  NAND2_X1 U4373 ( .A1(n3800), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3544) );
  INV_X1 U4374 ( .A(n3540), .ZN(n3543) );
  INV_X1 U4375 ( .A(n3561), .ZN(n3541) );
  NAND2_X1 U4376 ( .A1(n3541), .A2(n3613), .ZN(n3542) );
  NAND2_X1 U4377 ( .A1(n3545), .A2(n3609), .ZN(n3549) );
  INV_X1 U4378 ( .A(n3611), .ZN(n3547) );
  INV_X1 U4379 ( .A(n3608), .ZN(n3546) );
  NAND2_X1 U4380 ( .A1(n3547), .A2(n3546), .ZN(n3548) );
  NAND2_X1 U4381 ( .A1(n3549), .A2(n3548), .ZN(n3601) );
  INV_X1 U4382 ( .A(n3550), .ZN(n3552) );
  NAND2_X1 U4383 ( .A1(n3554), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3560) );
  INV_X1 U4384 ( .A(n3556), .ZN(n3555) );
  NAND2_X1 U4385 ( .A1(n3555), .A2(n7010), .ZN(n6918) );
  NAND2_X1 U4386 ( .A1(n3556), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3557) );
  NAND2_X1 U4387 ( .A1(n6918), .A2(n3557), .ZN(n4262) );
  AOI22_X1 U4388 ( .A1(n3558), .A2(n4262), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n4143), .ZN(n3559) );
  XNOR2_X2 U4389 ( .A(n3575), .B(n3576), .ZN(n4060) );
  INV_X1 U4390 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4780) );
  AOI22_X1 U4391 ( .A1(n5485), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4392 ( .A1(n5333), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4393 ( .A1(n5307), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4394 ( .A1(n5332), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4395 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3572)
         );
  AOI22_X1 U4396 ( .A1(n3525), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4397 ( .A1(n5486), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4398 ( .A1(n5460), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4399 ( .A1(n5338), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4400 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3571)
         );
  OR2_X1 U4401 ( .A1(n3572), .A2(n3571), .ZN(n3594) );
  NAND2_X1 U4402 ( .A1(n3781), .A2(n3594), .ZN(n3573) );
  OAI21_X1 U4403 ( .B1(n3790), .B2(n4780), .A(n3573), .ZN(n3574) );
  NAND2_X1 U4404 ( .A1(n3554), .A2(n6301), .ZN(n3580) );
  NOR3_X1 U4405 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n7010), .A3(n7005), 
        .ZN(n6855) );
  NAND2_X1 U4406 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6855), .ZN(n4309) );
  NAND2_X1 U4407 ( .A1(n7016), .A2(n4309), .ZN(n3577) );
  NOR3_X1 U4408 ( .A1(n7016), .A2(n7010), .A3(n7005), .ZN(n4809) );
  NAND2_X1 U4409 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4809), .ZN(n4906) );
  NAND2_X1 U4410 ( .A1(n3577), .A2(n4906), .ZN(n4261) );
  OAI22_X1 U4411 ( .A1(n4080), .A2(n4261), .B1(n3822), .B2(n7016), .ZN(n3578)
         );
  INV_X1 U4412 ( .A(n3578), .ZN(n3579) );
  AOI22_X1 U4413 ( .A1(n5332), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4414 ( .A1(n5476), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4415 ( .A1(n5486), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3583) );
  INV_X2 U4416 ( .A(n3581), .ZN(n5479) );
  AOI22_X1 U4417 ( .A1(n5460), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3582) );
  NAND4_X1 U4418 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3591)
         );
  AOI22_X1 U4419 ( .A1(n5307), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4420 ( .A1(n3525), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4421 ( .A1(n5478), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4422 ( .A1(n5338), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3586) );
  NAND4_X1 U4423 ( .A1(n3589), .A2(n3588), .A3(n3587), .A4(n3586), .ZN(n3590)
         );
  AOI22_X1 U4424 ( .A1(n3800), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3781), 
        .B2(n3655), .ZN(n3592) );
  NAND2_X1 U4425 ( .A1(n4208), .A2(n3794), .ZN(n3599) );
  NAND2_X1 U4426 ( .A1(n3626), .A2(n3613), .ZN(n3604) );
  INV_X1 U4427 ( .A(n3594), .ZN(n3603) );
  NAND2_X1 U4428 ( .A1(n3604), .A2(n3603), .ZN(n3656) );
  INV_X1 U4429 ( .A(n3655), .ZN(n3595) );
  XNOR2_X1 U4430 ( .A(n3656), .B(n3595), .ZN(n3597) );
  NAND2_X1 U4431 ( .A1(n3597), .A2(n3596), .ZN(n3598) );
  INV_X1 U4432 ( .A(n6686), .ZN(n3638) );
  NAND2_X1 U4433 ( .A1(n3601), .A2(n3600), .ZN(n3602) );
  XNOR2_X1 U4434 ( .A(n3604), .B(n3603), .ZN(n3606) );
  NAND2_X1 U4435 ( .A1(n3473), .A2(n4289), .ZN(n3625) );
  INV_X1 U4436 ( .A(n3625), .ZN(n3605) );
  AOI21_X1 U4437 ( .B1(n3606), .B2(n3596), .A(n3605), .ZN(n3607) );
  NAND2_X1 U4438 ( .A1(n6695), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3634)
         );
  INV_X1 U4439 ( .A(n3609), .ZN(n3610) );
  NAND2_X1 U4440 ( .A1(n4263), .A2(n3794), .ZN(n3618) );
  XNOR2_X1 U4441 ( .A(n3626), .B(n3613), .ZN(n3615) );
  INV_X1 U4442 ( .A(n3932), .ZN(n3614) );
  OAI211_X1 U4443 ( .C1(n3615), .C2(n7162), .A(n3614), .B(n4279), .ZN(n3616)
         );
  INV_X1 U4444 ( .A(n3616), .ZN(n3617) );
  NAND2_X1 U4445 ( .A1(n3619), .A2(n3622), .ZN(n3620) );
  OAI21_X1 U4446 ( .B1(n7162), .B2(n3626), .A(n3625), .ZN(n3627) );
  INV_X1 U4447 ( .A(n3627), .ZN(n3628) );
  NAND2_X1 U4448 ( .A1(n4076), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3629)
         );
  INV_X1 U4449 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U4450 ( .A1(n3629), .A2(n6805), .ZN(n3631) );
  AND2_X1 U4451 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3630) );
  NAND2_X1 U4452 ( .A1(n4076), .A2(n3630), .ZN(n3632) );
  AND2_X1 U4453 ( .A1(n3631), .A2(n3632), .ZN(n4153) );
  INV_X1 U4454 ( .A(n3632), .ZN(n3633) );
  NAND2_X1 U4455 ( .A1(n3634), .A2(n6697), .ZN(n3636) );
  OR2_X1 U4456 ( .A1(n6695), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3635)
         );
  NAND2_X1 U4457 ( .A1(n3636), .A2(n3635), .ZN(n6687) );
  INV_X1 U4458 ( .A(n6687), .ZN(n3637) );
  NAND2_X1 U4459 ( .A1(n3638), .A2(n3637), .ZN(n6689) );
  NAND2_X1 U4460 ( .A1(n3639), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3640)
         );
  INV_X1 U4461 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5893) );
  AOI22_X1 U4462 ( .A1(n5485), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4463 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5476), .B1(n3643), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4464 ( .A1(n5307), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4465 ( .A1(n5332), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3644) );
  NAND4_X1 U4466 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3653)
         );
  AOI22_X1 U4467 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5480), .B1(n3525), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4468 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5486), .B1(n5221), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4469 ( .A1(n5460), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4470 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5338), .B1(n5487), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3648) );
  NAND4_X1 U4471 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3652)
         );
  NAND2_X1 U4472 ( .A1(n3781), .A2(n3698), .ZN(n3654) );
  OAI21_X1 U4473 ( .B1(n3790), .B2(n5893), .A(n3654), .ZN(n3663) );
  NAND2_X1 U4474 ( .A1(n4215), .A2(n3794), .ZN(n3659) );
  NAND2_X1 U4475 ( .A1(n3656), .A2(n3655), .ZN(n3700) );
  XNOR2_X1 U4476 ( .A(n3700), .B(n3698), .ZN(n3657) );
  NAND2_X1 U4477 ( .A1(n3657), .A2(n3596), .ZN(n3658) );
  NAND2_X1 U4478 ( .A1(n3659), .A2(n3658), .ZN(n3660) );
  INV_X1 U4479 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6784) );
  NAND2_X1 U4480 ( .A1(n3660), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3661)
         );
  NAND2_X1 U4481 ( .A1(n4253), .A2(n3661), .ZN(n6678) );
  INV_X1 U4482 ( .A(n3662), .ZN(n3664) );
  NAND2_X1 U4483 ( .A1(n3664), .A2(n3663), .ZN(n3683) );
  INV_X1 U4484 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4788) );
  AOI22_X1 U4485 ( .A1(n5478), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4486 ( .A1(n5333), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4487 ( .A1(n5460), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4488 ( .A1(n5485), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3665) );
  NAND4_X1 U4489 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(n3674)
         );
  AOI22_X1 U4490 ( .A1(n5332), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5307), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4491 ( .A1(n5486), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4492 ( .A1(n3525), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4493 ( .A1(n5338), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4494 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3673)
         );
  NAND2_X1 U4495 ( .A1(n3781), .A2(n3697), .ZN(n3675) );
  OAI21_X1 U4496 ( .B1(n3790), .B2(n4788), .A(n3675), .ZN(n3684) );
  NAND2_X1 U4497 ( .A1(n4236), .A2(n3794), .ZN(n3680) );
  INV_X1 U4498 ( .A(n3698), .ZN(n3676) );
  OR2_X1 U4499 ( .A1(n3700), .A2(n3676), .ZN(n3677) );
  XNOR2_X1 U4500 ( .A(n3677), .B(n3697), .ZN(n3678) );
  NAND2_X1 U4501 ( .A1(n3678), .A2(n3596), .ZN(n3679) );
  INV_X1 U4502 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6751) );
  NAND2_X1 U4503 ( .A1(n3681), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3682)
         );
  NAND2_X1 U4504 ( .A1(n6676), .A2(n3682), .ZN(n4513) );
  INV_X1 U4505 ( .A(n3683), .ZN(n3685) );
  NAND2_X1 U4506 ( .A1(n3685), .A2(n3684), .ZN(n3706) );
  INV_X1 U4507 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4794) );
  AOI22_X1 U4508 ( .A1(n5485), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4509 ( .A1(n5333), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4510 ( .A1(n5307), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4511 ( .A1(n5332), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3686) );
  NAND4_X1 U4512 ( .A1(n3689), .A2(n3688), .A3(n3687), .A4(n3686), .ZN(n3695)
         );
  INV_X1 U4513 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5853) );
  AOI22_X1 U4514 ( .A1(n3525), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4515 ( .A1(n5486), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4516 ( .A1(n5460), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4517 ( .A1(n5338), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3690) );
  NAND4_X1 U4518 ( .A1(n3693), .A2(n3692), .A3(n3691), .A4(n3690), .ZN(n3694)
         );
  NAND2_X1 U4519 ( .A1(n3781), .A2(n3712), .ZN(n3696) );
  OAI21_X1 U4520 ( .B1(n3790), .B2(n4794), .A(n3696), .ZN(n3707) );
  NAND2_X1 U4521 ( .A1(n4318), .A2(n3794), .ZN(n3703) );
  NAND2_X1 U4522 ( .A1(n3698), .A2(n3697), .ZN(n3699) );
  OR2_X1 U4523 ( .A1(n3700), .A2(n3699), .ZN(n3711) );
  XNOR2_X1 U4524 ( .A(n3711), .B(n3712), .ZN(n3701) );
  NAND2_X1 U4525 ( .A1(n3701), .A2(n3596), .ZN(n3702) );
  NAND2_X1 U4526 ( .A1(n3703), .A2(n3702), .ZN(n3704) );
  INV_X1 U4527 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6761) );
  XNOR2_X1 U4528 ( .A(n3704), .B(n6761), .ZN(n4515) );
  NAND2_X1 U4529 ( .A1(n4513), .A2(n4515), .ZN(n4514) );
  NAND2_X1 U4530 ( .A1(n3704), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3705)
         );
  NAND2_X1 U4531 ( .A1(n4514), .A2(n3705), .ZN(n6668) );
  INV_X1 U4532 ( .A(n3706), .ZN(n3708) );
  INV_X1 U4533 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4769) );
  NAND2_X1 U4534 ( .A1(n3781), .A2(n3723), .ZN(n3709) );
  OAI21_X1 U4535 ( .B1(n3790), .B2(n4769), .A(n3709), .ZN(n3710) );
  NAND2_X1 U4536 ( .A1(n4413), .A2(n3794), .ZN(n3716) );
  INV_X1 U4537 ( .A(n3711), .ZN(n3713) );
  NAND2_X1 U4538 ( .A1(n3713), .A2(n3712), .ZN(n3722) );
  XNOR2_X1 U4539 ( .A(n3722), .B(n3723), .ZN(n3714) );
  NAND2_X1 U4540 ( .A1(n3714), .A2(n3596), .ZN(n3715) );
  NAND2_X1 U4541 ( .A1(n3716), .A2(n3715), .ZN(n3717) );
  INV_X1 U4542 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6741) );
  XNOR2_X1 U4543 ( .A(n3717), .B(n6741), .ZN(n6670) );
  NAND2_X1 U4544 ( .A1(n3717), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3718)
         );
  NAND2_X1 U4545 ( .A1(n6669), .A2(n3718), .ZN(n4581) );
  NOR2_X1 U4546 ( .A1(n3719), .A2(n3762), .ZN(n3720) );
  INV_X4 U4547 ( .A(n6131), .ZN(n6263) );
  INV_X1 U4548 ( .A(n3722), .ZN(n3724) );
  NAND3_X1 U4549 ( .A1(n3724), .A2(n3596), .A3(n3723), .ZN(n3725) );
  NAND2_X1 U4550 ( .A1(n6263), .A2(n3725), .ZN(n3726) );
  INV_X1 U4551 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6734) );
  XNOR2_X1 U4552 ( .A(n3726), .B(n6734), .ZN(n4580) );
  NAND2_X1 U4553 ( .A1(n4581), .A2(n4580), .ZN(n4583) );
  NAND2_X1 U4554 ( .A1(n3726), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3727)
         );
  XNOR2_X1 U4555 ( .A(n6262), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4744)
         );
  INV_X1 U4556 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6724) );
  OR2_X1 U4557 ( .A1(n6263), .A2(n6724), .ZN(n3728) );
  INV_X1 U4558 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U4559 ( .A1(n6263), .A2(n5891), .ZN(n5019) );
  INV_X1 U4560 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5256) );
  OR2_X2 U4561 ( .A1(n6263), .A2(n5891), .ZN(n5093) );
  OR2_X1 U4562 ( .A1(n6263), .A2(n5256), .ZN(n5096) );
  INV_X1 U4563 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5841) );
  INV_X1 U4564 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5257) );
  XNOR2_X1 U4565 ( .A(n6262), .B(n5257), .ZN(n5216) );
  NAND2_X1 U4566 ( .A1(n6263), .A2(n5257), .ZN(n3731) );
  INV_X1 U4567 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U4568 ( .A1(n6263), .A2(n6388), .ZN(n5247) );
  INV_X1 U4569 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3732) );
  NAND2_X1 U4570 ( .A1(n3734), .A2(n6131), .ZN(n3736) );
  INV_X1 U4571 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U4572 ( .A1(n6263), .A2(n6391), .ZN(n6165) );
  AND2_X1 U4573 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3951) );
  NAND2_X1 U4574 ( .A1(n6264), .A2(n3735), .ZN(n6147) );
  AND2_X1 U4575 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6231) );
  AND2_X1 U4576 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3950) );
  NAND2_X1 U4577 ( .A1(n6231), .A2(n3950), .ZN(n5553) );
  NAND2_X1 U4578 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3956) );
  NOR2_X1 U4579 ( .A1(n5553), .A2(n3956), .ZN(n3737) );
  OR2_X1 U4580 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3738) );
  NOR2_X1 U4581 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6232) );
  INV_X1 U4582 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6122) );
  INV_X1 U4583 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6216) );
  XNOR2_X1 U4584 ( .A(n6262), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6115)
         );
  INV_X1 U4585 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U4586 ( .A1(n6263), .A2(n6212), .ZN(n3739) );
  INV_X1 U4587 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U4588 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3964) );
  INV_X1 U4589 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7063) );
  NAND2_X1 U4590 ( .A1(n3741), .A2(n7063), .ZN(n7060) );
  NAND2_X1 U4591 ( .A1(n3447), .A2(n7060), .ZN(n3760) );
  XNOR2_X1 U4592 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4593 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n7005), .B1(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3743), .ZN(n3745) );
  NAND2_X1 U4594 ( .A1(n7000), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3767) );
  NAND2_X1 U4595 ( .A1(n3745), .A2(n3744), .ZN(n3742) );
  OAI21_X1 U4596 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3743), .A(n3742), 
        .ZN(n3747) );
  XOR2_X1 U4597 ( .A(n3746), .B(n3747), .Z(n3784) );
  XOR2_X1 U4598 ( .A(n3745), .B(n3744), .Z(n3774) );
  NAND2_X1 U4599 ( .A1(n3747), .A2(n3746), .ZN(n3749) );
  NAND2_X1 U4600 ( .A1(n7010), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3748) );
  NAND2_X1 U4601 ( .A1(n3749), .A2(n3748), .ZN(n3752) );
  XNOR2_X1 U4602 ( .A(n6301), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3751)
         );
  INV_X1 U4603 ( .A(n3751), .ZN(n3750) );
  XNOR2_X1 U4604 ( .A(n3752), .B(n3750), .ZN(n3798) );
  NAND2_X1 U4605 ( .A1(n3752), .A2(n3751), .ZN(n3754) );
  NAND2_X1 U4606 ( .A1(n7016), .A2(n6301), .ZN(n3753) );
  NAND2_X1 U4607 ( .A1(n3754), .A2(n3753), .ZN(n3756) );
  INV_X1 U4608 ( .A(n3756), .ZN(n3793) );
  INV_X1 U4609 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7014) );
  NOR2_X1 U4610 ( .A1(n7014), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3792)
         );
  NAND2_X1 U4611 ( .A1(n3793), .A2(n3792), .ZN(n3799) );
  NAND4_X1 U4612 ( .A1(n3784), .A2(n3774), .A3(n3798), .A4(n3799), .ZN(n3759)
         );
  AND2_X1 U4613 ( .A1(n7014), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3755)
         );
  INV_X1 U4614 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U4615 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6407), .ZN(n3757) );
  NAND2_X1 U4616 ( .A1(n3758), .A2(n3757), .ZN(n3805) );
  NAND2_X1 U4617 ( .A1(n3759), .A2(n3805), .ZN(n4011) );
  NOR2_X1 U4618 ( .A1(READY_N), .A2(n4011), .ZN(n4048) );
  NAND2_X1 U4619 ( .A1(n3760), .A2(n4048), .ZN(n3811) );
  OR2_X1 U4620 ( .A1(n3761), .A2(READY_N), .ZN(n4338) );
  AND2_X1 U4621 ( .A1(n3596), .A2(n7060), .ZN(n3987) );
  AOI21_X1 U4622 ( .B1(n4338), .B2(n4097), .A(n3987), .ZN(n3808) );
  INV_X1 U4623 ( .A(n3805), .ZN(n3763) );
  NAND2_X1 U4624 ( .A1(n3763), .A2(n3791), .ZN(n3807) );
  INV_X1 U4625 ( .A(n3798), .ZN(n3789) );
  NAND2_X1 U4626 ( .A1(n3430), .A2(n4097), .ZN(n3764) );
  NAND2_X1 U4627 ( .A1(n3764), .A2(n3479), .ZN(n3783) );
  INV_X1 U4628 ( .A(n3783), .ZN(n3765) );
  NAND3_X1 U4629 ( .A1(n3765), .A2(n3781), .A3(n3784), .ZN(n3788) );
  NAND2_X1 U4630 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3774), .ZN(n3780) );
  AOI21_X1 U4631 ( .B1(n3781), .B2(n3447), .A(n3430), .ZN(n3779) );
  NAND2_X1 U4632 ( .A1(n3779), .A2(n3780), .ZN(n3771) );
  OAI21_X1 U4633 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7000), .A(n3767), 
        .ZN(n3772) );
  OAI21_X1 U4634 ( .B1(n3466), .B2(n3772), .A(n3768), .ZN(n3769) );
  NAND2_X1 U4635 ( .A1(n3769), .A2(n3783), .ZN(n3770) );
  NOR2_X1 U4636 ( .A1(n3804), .A2(n3772), .ZN(n3773) );
  NAND2_X1 U4637 ( .A1(n3775), .A2(n3773), .ZN(n3778) );
  INV_X1 U4638 ( .A(n3774), .ZN(n3776) );
  OAI21_X1 U4639 ( .B1(n3776), .B2(n3775), .A(n3791), .ZN(n3777) );
  OAI211_X1 U4640 ( .C1(n3780), .C2(n3779), .A(n3778), .B(n3777), .ZN(n3786)
         );
  NAND2_X1 U4641 ( .A1(n3781), .A2(n3784), .ZN(n3782) );
  OAI211_X1 U4642 ( .C1(n3784), .C2(n3790), .A(n3783), .B(n3782), .ZN(n3785)
         );
  NAND2_X1 U4643 ( .A1(n3786), .A2(n3785), .ZN(n3787) );
  AOI22_X1 U4644 ( .A1(n3790), .A2(n3789), .B1(n3788), .B2(n3787), .ZN(n3802)
         );
  INV_X1 U4645 ( .A(n3791), .ZN(n3797) );
  NAND2_X1 U4646 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n7028), .ZN(n3796) );
  NAND3_X1 U4647 ( .A1(n3794), .A2(n3793), .A3(n3792), .ZN(n3795) );
  OAI211_X1 U4648 ( .C1(n3798), .C2(n3797), .A(n3796), .B(n3795), .ZN(n3801)
         );
  OAI22_X1 U4649 ( .A1(n3802), .A2(n3801), .B1(n3800), .B2(n3799), .ZN(n3803)
         );
  INV_X1 U4650 ( .A(n4040), .ZN(n4046) );
  OAI21_X1 U4651 ( .B1(n3808), .B2(n3295), .A(n4046), .ZN(n3810) );
  MUX2_X1 U4652 ( .A(n3811), .B(n3810), .S(n3809), .Z(n3821) );
  NAND2_X1 U4653 ( .A1(n3444), .A2(n4294), .ZN(n3812) );
  OR2_X1 U4654 ( .A1(n3452), .A2(n3812), .ZN(n4970) );
  NOR2_X1 U4655 ( .A1(n4970), .A2(n3479), .ZN(n3944) );
  NAND2_X1 U4656 ( .A1(n4040), .A2(n3944), .ZN(n4052) );
  INV_X1 U4657 ( .A(n3813), .ZN(n3820) );
  NAND2_X1 U4658 ( .A1(n4970), .A2(n3473), .ZN(n3814) );
  AND2_X1 U4659 ( .A1(n3815), .A2(n3814), .ZN(n3827) );
  OR3_X1 U4660 ( .A1(n3817), .A2(n3473), .A3(n3816), .ZN(n3936) );
  NAND3_X1 U4661 ( .A1(n3827), .A2(n3818), .A3(n3936), .ZN(n3819) );
  NAND2_X1 U4662 ( .A1(n3820), .A2(n3819), .ZN(n4050) );
  NAND3_X1 U4663 ( .A1(n3821), .A2(n4052), .A3(n4050), .ZN(n3823) );
  AND2_X1 U4664 ( .A1(n3822), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7036) );
  AND2_X1 U4665 ( .A1(n3466), .A2(n3827), .ZN(n4077) );
  INV_X1 U4666 ( .A(n4077), .ZN(n6989) );
  OAI22_X1 U4667 ( .A1(n3761), .A2(n5526), .B1(n3518), .B2(n3926), .ZN(n3824)
         );
  INV_X1 U4668 ( .A(n3824), .ZN(n3828) );
  NAND2_X1 U4669 ( .A1(n3827), .A2(n3826), .ZN(n4335) );
  AND4_X1 U4670 ( .A1(n6989), .A2(n3828), .A3(n3191), .A4(n4335), .ZN(n3829)
         );
  INV_X1 U4671 ( .A(n4289), .ZN(n3830) );
  NAND2_X1 U4672 ( .A1(n3917), .A2(n6805), .ZN(n3832) );
  INV_X1 U4673 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4167) );
  NAND2_X1 U4674 ( .A1(n4144), .A2(n4167), .ZN(n3831) );
  NAND3_X1 U4675 ( .A1(n3832), .A2(n3913), .A3(n3831), .ZN(n3834) );
  NAND2_X1 U4676 ( .A1(n5537), .A2(n4167), .ZN(n3833) );
  NAND2_X1 U4677 ( .A1(n3834), .A2(n3833), .ZN(n3838) );
  NAND2_X1 U4678 ( .A1(n3917), .A2(EBX_REG_0__SCAN_IN), .ZN(n3837) );
  INV_X1 U4679 ( .A(EBX_REG_0__SCAN_IN), .ZN(n3835) );
  NAND2_X1 U4680 ( .A1(n3913), .A2(n3835), .ZN(n3836) );
  NAND2_X1 U4681 ( .A1(n3837), .A2(n3836), .ZN(n3989) );
  XNOR2_X1 U4682 ( .A(n3838), .B(n3989), .ZN(n5029) );
  NAND2_X1 U4683 ( .A1(n4144), .A2(n3913), .ZN(n3906) );
  MUX2_X1 U4684 ( .A(n3906), .B(n3913), .S(EBX_REG_3__SCAN_IN), .Z(n3840) );
  OR2_X1 U4685 ( .A1(n3852), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3839)
         );
  NAND2_X1 U4686 ( .A1(n3840), .A2(n3839), .ZN(n4247) );
  NAND2_X1 U4687 ( .A1(n3852), .A2(EBX_REG_2__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U4688 ( .A1(n5526), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3841)
         );
  NAND2_X1 U4689 ( .A1(n3842), .A2(n3841), .ZN(n3843) );
  XNOR2_X1 U4690 ( .A(n3843), .B(n5537), .ZN(n4248) );
  NAND2_X1 U4691 ( .A1(n3913), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3844)
         );
  AND2_X1 U4692 ( .A1(n3917), .A2(n3844), .ZN(n3846) );
  NOR2_X1 U4693 ( .A1(n5526), .A2(EBX_REG_4__SCAN_IN), .ZN(n3845) );
  MUX2_X1 U4694 ( .A(n3846), .B(n3913), .S(n3845), .Z(n4206) );
  MUX2_X1 U4695 ( .A(n3906), .B(n3913), .S(EBX_REG_5__SCAN_IN), .Z(n3848) );
  OR2_X1 U4696 ( .A1(n3852), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3847)
         );
  AND2_X1 U4697 ( .A1(n3848), .A2(n3847), .ZN(n4233) );
  NAND2_X1 U4698 ( .A1(n4234), .A2(n4233), .ZN(n4316) );
  NAND2_X1 U4699 ( .A1(n3913), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3849)
         );
  AND2_X1 U4700 ( .A1(n3917), .A2(n3849), .ZN(n3851) );
  NOR2_X1 U4701 ( .A1(n5526), .A2(EBX_REG_6__SCAN_IN), .ZN(n3850) );
  MUX2_X1 U4702 ( .A(n3851), .B(n3913), .S(n3850), .Z(n4315) );
  NAND2_X1 U4703 ( .A1(n3852), .A2(EBX_REG_7__SCAN_IN), .ZN(n3854) );
  NAND2_X1 U4704 ( .A1(n5526), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3853)
         );
  NAND2_X1 U4705 ( .A1(n3854), .A2(n3853), .ZN(n3855) );
  XNOR2_X1 U4706 ( .A(n3855), .B(n5537), .ZN(n4446) );
  NAND2_X1 U4707 ( .A1(n3917), .A2(n6734), .ZN(n3857) );
  INV_X1 U4708 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U4709 ( .A1(n4144), .A2(n5146), .ZN(n3856) );
  NAND3_X1 U4710 ( .A1(n3857), .A2(n3913), .A3(n3856), .ZN(n3859) );
  NAND2_X1 U4711 ( .A1(n5537), .A2(n5146), .ZN(n3858) );
  NAND2_X1 U4712 ( .A1(n3859), .A2(n3858), .ZN(n4508) );
  INV_X1 U4713 ( .A(n3906), .ZN(n3912) );
  INV_X1 U4714 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U4715 ( .A1(n3912), .A2(n6494), .ZN(n3862) );
  NAND2_X1 U4716 ( .A1(n3913), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3860)
         );
  OAI211_X1 U4717 ( .C1(n5526), .C2(EBX_REG_9__SCAN_IN), .A(n3917), .B(n3860), 
        .ZN(n3861) );
  NAND2_X1 U4718 ( .A1(n3852), .A2(EBX_REG_10__SCAN_IN), .ZN(n3864) );
  NAND2_X1 U4719 ( .A1(n5526), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3863) );
  NAND2_X1 U4720 ( .A1(n3864), .A2(n3863), .ZN(n3865) );
  XNOR2_X1 U4721 ( .A(n3865), .B(n5537), .ZN(n4894) );
  MUX2_X1 U4722 ( .A(n3906), .B(n3913), .S(EBX_REG_11__SCAN_IN), .Z(n3866) );
  OAI21_X1 U4723 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n3852), .A(n3866), 
        .ZN(n4957) );
  MUX2_X1 U4724 ( .A(n3906), .B(n3913), .S(EBX_REG_13__SCAN_IN), .Z(n3868) );
  OR2_X1 U4725 ( .A1(n3852), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3867)
         );
  NAND2_X1 U4726 ( .A1(n3868), .A2(n3867), .ZN(n5050) );
  NAND2_X1 U4727 ( .A1(n3917), .A2(n5841), .ZN(n3870) );
  INV_X1 U4728 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U4729 ( .A1(n4144), .A2(n6464), .ZN(n3869) );
  NAND3_X1 U4730 ( .A1(n3870), .A2(n3913), .A3(n3869), .ZN(n3872) );
  NAND2_X1 U4731 ( .A1(n5537), .A2(n6464), .ZN(n3871) );
  AND2_X1 U4732 ( .A1(n3872), .A2(n3871), .ZN(n5049) );
  NOR2_X1 U4733 ( .A1(n5050), .A2(n5049), .ZN(n3873) );
  NAND2_X1 U4734 ( .A1(n3852), .A2(EBX_REG_14__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U4735 ( .A1(n5526), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3874) );
  NAND2_X1 U4736 ( .A1(n3875), .A2(n3874), .ZN(n3876) );
  XNOR2_X1 U4737 ( .A(n3876), .B(n3913), .ZN(n4968) );
  MUX2_X1 U4738 ( .A(n3906), .B(n3877), .S(EBX_REG_15__SCAN_IN), .Z(n3878) );
  OAI21_X1 U4739 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n3852), .A(n3878), 
        .ZN(n4740) );
  NAND2_X1 U4740 ( .A1(n3913), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3879) );
  AND2_X1 U4741 ( .A1(n3917), .A2(n3879), .ZN(n3881) );
  NOR2_X1 U4742 ( .A1(n5526), .A2(EBX_REG_16__SCAN_IN), .ZN(n3880) );
  MUX2_X1 U4743 ( .A(n3881), .B(n3913), .S(n3880), .Z(n4988) );
  MUX2_X1 U4744 ( .A(n3906), .B(n3913), .S(EBX_REG_17__SCAN_IN), .Z(n3882) );
  OAI21_X1 U4745 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n3852), .A(n3882), 
        .ZN(n5118) );
  NOR2_X2 U4746 ( .A1(n5119), .A2(n5118), .ZN(n5159) );
  INV_X1 U4747 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U4748 ( .A1(n3917), .A2(n6246), .ZN(n3884) );
  INV_X1 U4749 ( .A(EBX_REG_19__SCAN_IN), .ZN(n3885) );
  NAND2_X1 U4750 ( .A1(n4144), .A2(n3885), .ZN(n3883) );
  NAND3_X1 U4751 ( .A1(n3884), .A2(n3913), .A3(n3883), .ZN(n3887) );
  NAND2_X1 U4752 ( .A1(n5537), .A2(n3885), .ZN(n3886) );
  NAND2_X1 U4753 ( .A1(n3887), .A2(n3886), .ZN(n5204) );
  NAND2_X1 U4754 ( .A1(n5159), .A2(n5204), .ZN(n5242) );
  OR2_X1 U4755 ( .A1(n3852), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3889)
         );
  INV_X1 U4756 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U4757 ( .A1(n4144), .A2(n5246), .ZN(n3888) );
  NAND2_X1 U4758 ( .A1(n3889), .A2(n3888), .ZN(n5244) );
  OR2_X1 U4759 ( .A1(n3852), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3890)
         );
  INV_X1 U4760 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U4761 ( .A1(n4144), .A2(n5182), .ZN(n5156) );
  NAND2_X1 U4762 ( .A1(n3890), .A2(n5156), .ZN(n5243) );
  MUX2_X1 U4763 ( .A(n5244), .B(n3913), .S(n5243), .Z(n3891) );
  INV_X1 U4764 ( .A(n3891), .ZN(n3893) );
  NAND2_X1 U4765 ( .A1(n5537), .A2(EBX_REG_20__SCAN_IN), .ZN(n3892) );
  NAND2_X1 U4766 ( .A1(n3893), .A2(n3892), .ZN(n3894) );
  NAND2_X1 U4767 ( .A1(n3852), .A2(EBX_REG_21__SCAN_IN), .ZN(n3896) );
  NAND2_X1 U4768 ( .A1(n5526), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3895) );
  NAND2_X1 U4769 ( .A1(n3896), .A2(n3895), .ZN(n3897) );
  XNOR2_X1 U4770 ( .A(n3897), .B(n5537), .ZN(n5294) );
  NAND2_X1 U4771 ( .A1(n3913), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3898) );
  NAND2_X1 U4772 ( .A1(n3917), .A2(n3898), .ZN(n3900) );
  INV_X1 U4773 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U4774 ( .A1(n4144), .A2(n6059), .ZN(n3899) );
  MUX2_X1 U4775 ( .A(n5537), .B(n3900), .S(n3899), .Z(n6007) );
  MUX2_X1 U4776 ( .A(n3906), .B(n3913), .S(EBX_REG_23__SCAN_IN), .Z(n3902) );
  OR2_X1 U4777 ( .A1(n3852), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3901)
         );
  NAND2_X1 U4778 ( .A1(n3902), .A2(n3901), .ZN(n5999) );
  NAND2_X1 U4779 ( .A1(n3852), .A2(EBX_REG_24__SCAN_IN), .ZN(n3904) );
  NAND2_X1 U4780 ( .A1(n5526), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3903) );
  NAND2_X1 U4781 ( .A1(n3904), .A2(n3903), .ZN(n3905) );
  XNOR2_X1 U4782 ( .A(n3905), .B(n5537), .ZN(n5975) );
  MUX2_X1 U4783 ( .A(n3906), .B(n3913), .S(EBX_REG_25__SCAN_IN), .Z(n3907) );
  OAI21_X1 U4784 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n3852), .A(n3907), 
        .ZN(n5966) );
  OR3_X2 U4785 ( .A1(n5996), .A2(n5975), .A3(n5966), .ZN(n6047) );
  NAND2_X1 U4786 ( .A1(n3917), .A2(n6204), .ZN(n3909) );
  INV_X1 U4787 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U4788 ( .A1(n4144), .A2(n6320), .ZN(n3908) );
  NAND3_X1 U4789 ( .A1(n3909), .A2(n3913), .A3(n3908), .ZN(n3911) );
  NAND2_X1 U4790 ( .A1(n5537), .A2(n6320), .ZN(n3910) );
  AND2_X1 U4791 ( .A1(n3911), .A2(n3910), .ZN(n6046) );
  NOR2_X2 U4792 ( .A1(n6047), .A2(n6046), .ZN(n6049) );
  INV_X1 U4793 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U4794 ( .A1(n3912), .A2(n6040), .ZN(n3916) );
  NAND2_X1 U4795 ( .A1(n3913), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3914) );
  OAI211_X1 U4796 ( .C1(n5526), .C2(EBX_REG_27__SCAN_IN), .A(n3917), .B(n3914), 
        .ZN(n3915) );
  AND2_X1 U4797 ( .A1(n3916), .A2(n3915), .ZN(n5954) );
  NAND2_X1 U4798 ( .A1(n6049), .A2(n5954), .ZN(n5956) );
  INV_X1 U4799 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U4800 ( .A1(n3917), .A2(n6179), .ZN(n3919) );
  INV_X1 U4801 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U4802 ( .A1(n4144), .A2(n6037), .ZN(n3918) );
  NAND3_X1 U4803 ( .A1(n3919), .A2(n3913), .A3(n3918), .ZN(n3921) );
  NAND2_X1 U4804 ( .A1(n5537), .A2(n6037), .ZN(n3920) );
  AND2_X1 U4805 ( .A1(n3921), .A2(n3920), .ZN(n5943) );
  OR2_X2 U4806 ( .A1(n5956), .A2(n5943), .ZN(n5945) );
  OR2_X1 U4807 ( .A1(n3852), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3923)
         );
  INV_X1 U4808 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U4809 ( .A1(n4144), .A2(n6035), .ZN(n3922) );
  NAND2_X1 U4810 ( .A1(n3923), .A2(n3922), .ZN(n5524) );
  MUX2_X1 U4811 ( .A(n5524), .B(EBX_REG_29__SCAN_IN), .S(n5537), .Z(n3924) );
  NOR2_X1 U4812 ( .A1(n5945), .A2(n3924), .ZN(n5525) );
  AND2_X1 U4813 ( .A1(n5945), .A2(n3924), .ZN(n3925) );
  NOR2_X1 U4814 ( .A1(n5525), .A2(n3925), .ZN(n6034) );
  OR2_X1 U4815 ( .A1(n3761), .A2(n7162), .ZN(n7023) );
  INV_X1 U4816 ( .A(n3926), .ZN(n3927) );
  NAND2_X1 U4817 ( .A1(n3927), .A2(n3518), .ZN(n3928) );
  AND2_X1 U4818 ( .A1(n7023), .A2(n3928), .ZN(n3929) );
  NOR2_X1 U4819 ( .A1(n4080), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U4820 ( .A1(n6803), .A2(REIP_REG_29__SCAN_IN), .ZN(n6083) );
  INV_X1 U4821 ( .A(n6083), .ZN(n3930) );
  AOI21_X1 U4822 ( .B1(n6034), .B2(n6799), .A(n3930), .ZN(n3968) );
  AOI21_X1 U4823 ( .B1(n3295), .B2(n3473), .A(n3809), .ZN(n3931) );
  AOI21_X1 U4824 ( .B1(n3458), .B2(n5537), .A(n3931), .ZN(n3935) );
  NOR2_X1 U4825 ( .A1(n3479), .A2(n3439), .ZN(n3933) );
  OAI21_X1 U4826 ( .B1(n3852), .B2(n3933), .A(n3932), .ZN(n3934) );
  AND3_X1 U4827 ( .A1(n3936), .A2(n3935), .A3(n3934), .ZN(n3937) );
  NAND2_X1 U4828 ( .A1(n3938), .A2(n3937), .ZN(n4029) );
  INV_X1 U4829 ( .A(n4970), .ZN(n6996) );
  NAND2_X1 U4830 ( .A1(n6996), .A2(n3476), .ZN(n4180) );
  INV_X1 U4831 ( .A(n3940), .ZN(n3941) );
  NAND2_X1 U4832 ( .A1(n3941), .A2(n3473), .ZN(n3942) );
  OAI211_X1 U4833 ( .C1(n3939), .C2(n3184), .A(n4180), .B(n3942), .ZN(n3943)
         );
  NOR2_X1 U4834 ( .A1(n4029), .A2(n3943), .ZN(n4054) );
  NAND2_X1 U4835 ( .A1(n4054), .A2(n3944), .ZN(n4061) );
  INV_X1 U4836 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6791) );
  NOR2_X1 U4837 ( .A1(n6791), .A2(n6784), .ZN(n6764) );
  INV_X1 U4838 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U4839 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6794) );
  NAND2_X1 U4840 ( .A1(n6793), .A2(n6794), .ZN(n6778) );
  NAND2_X1 U4841 ( .A1(n6764), .A2(n6778), .ZN(n6749) );
  NOR2_X1 U4842 ( .A1(n6795), .A2(n6749), .ZN(n6762) );
  NAND3_X1 U4843 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6762), .ZN(n5023) );
  NOR2_X1 U4844 ( .A1(n6741), .A2(n6734), .ZN(n6727) );
  NAND3_X1 U4845 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6727), .ZN(n3947) );
  NAND3_X1 U4846 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n6389) );
  NOR2_X1 U4847 ( .A1(n6388), .A2(n6389), .ZN(n6384) );
  NAND3_X1 U4848 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6384), .ZN(n3948) );
  INV_X1 U4849 ( .A(n3948), .ZN(n3962) );
  NAND2_X1 U4850 ( .A1(n5262), .A2(n3962), .ZN(n6242) );
  INV_X1 U4851 ( .A(n6795), .ZN(n6746) );
  NOR2_X1 U4852 ( .A1(n3945), .A2(n4054), .ZN(n5263) );
  NOR2_X1 U4853 ( .A1(n6746), .A2(n5263), .ZN(n5261) );
  NOR2_X1 U4854 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5261), .ZN(n4089)
         );
  AND2_X1 U4855 ( .A1(n3945), .A2(n6774), .ZN(n4086) );
  NOR2_X1 U4856 ( .A1(n4089), .A2(n4086), .ZN(n6745) );
  NAND2_X1 U4857 ( .A1(n6795), .A2(n6745), .ZN(n6241) );
  NAND2_X1 U4858 ( .A1(n6242), .A2(n6241), .ZN(n3954) );
  NAND2_X1 U4859 ( .A1(n3813), .A2(n3447), .ZN(n4182) );
  INV_X1 U4860 ( .A(n6764), .ZN(n6781) );
  NAND2_X1 U4861 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3946) );
  NAND2_X1 U4862 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6744) );
  OR3_X1 U4863 ( .A1(n6781), .A2(n3946), .A3(n6744), .ZN(n5022) );
  OR2_X1 U4864 ( .A1(n3947), .A2(n5022), .ZN(n3961) );
  NAND2_X1 U4865 ( .A1(n6743), .A2(n3961), .ZN(n5107) );
  NAND2_X1 U4866 ( .A1(n6743), .A2(n3948), .ZN(n3949) );
  AND2_X1 U4867 ( .A1(n5107), .A2(n3949), .ZN(n6244) );
  NAND2_X1 U4868 ( .A1(n3951), .A2(n3950), .ZN(n5546) );
  OAI21_X1 U4869 ( .B1(n6743), .B2(n6241), .A(n5546), .ZN(n3952) );
  AND2_X1 U4870 ( .A1(n6244), .A2(n3952), .ZN(n3953) );
  NAND2_X1 U4871 ( .A1(n3954), .A2(n3953), .ZN(n6369) );
  INV_X1 U4872 ( .A(n6231), .ZN(n6223) );
  AND2_X1 U4873 ( .A1(n6750), .A2(n6223), .ZN(n3955) );
  OR2_X1 U4874 ( .A1(n5258), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4160)
         );
  NAND2_X1 U4875 ( .A1(n6743), .A2(n4160), .ZN(n6804) );
  INV_X1 U4876 ( .A(n3956), .ZN(n5556) );
  AOI21_X1 U4877 ( .B1(n6804), .B2(n6795), .A(n5556), .ZN(n3957) );
  AND2_X1 U4878 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6199) );
  INV_X1 U4879 ( .A(n6199), .ZN(n3958) );
  NAND2_X1 U4880 ( .A1(n6750), .A2(n3958), .ZN(n3959) );
  AND2_X1 U4881 ( .A1(n6214), .A2(n3959), .ZN(n6178) );
  NAND2_X1 U4882 ( .A1(n6750), .A2(n3964), .ZN(n3960) );
  AND2_X1 U4883 ( .A1(n6178), .A2(n3960), .ZN(n5516) );
  NAND2_X1 U4884 ( .A1(n5516), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5542) );
  NOR2_X1 U4885 ( .A1(n3961), .A2(n6804), .ZN(n5110) );
  NAND2_X1 U4886 ( .A1(n3962), .A2(n5110), .ZN(n6240) );
  NAND2_X1 U4887 ( .A1(n6242), .A2(n6240), .ZN(n6375) );
  NAND3_X1 U4888 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n6375), .ZN(n6257) );
  INV_X1 U4889 ( .A(n6257), .ZN(n6247) );
  NAND2_X1 U4890 ( .A1(n5556), .A2(n6247), .ZN(n3963) );
  NOR2_X1 U4891 ( .A1(n5553), .A2(n3963), .ZN(n6197) );
  INV_X1 U4892 ( .A(n3964), .ZN(n3965) );
  NAND2_X1 U4893 ( .A1(n6188), .A2(n3965), .ZN(n5540) );
  INV_X1 U4894 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U4895 ( .A1(n5540), .A2(n5539), .ZN(n3966) );
  NAND2_X1 U4896 ( .A1(n5542), .A2(n3966), .ZN(n3967) );
  NAND2_X1 U4897 ( .A1(n6817), .A2(n3969), .ZN(n3970) );
  NAND2_X1 U4898 ( .A1(n3970), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3976) );
  INV_X1 U4899 ( .A(n3976), .ZN(n3978) );
  NAND2_X1 U4900 ( .A1(n3295), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4218) );
  NAND2_X1 U4901 ( .A1(n5510), .A2(EAX_REG_0__SCAN_IN), .ZN(n3974) );
  NAND2_X1 U4902 ( .A1(n6930), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3973)
         );
  OAI211_X1 U4903 ( .C1(n4218), .C2(n3272), .A(n3974), .B(n3973), .ZN(n3975)
         );
  AOI21_X1 U4904 ( .B1(n6995), .B2(n3972), .A(n3975), .ZN(n4122) );
  INV_X1 U4905 ( .A(n4122), .ZN(n3977) );
  OR2_X1 U4906 ( .A1(n3976), .A2(n4122), .ZN(n4124) );
  OAI21_X1 U4907 ( .B1(n3978), .B2(n3977), .A(n4124), .ZN(n4373) );
  INV_X1 U4908 ( .A(n7036), .ZN(n7033) );
  INV_X1 U4909 ( .A(n4016), .ZN(n4009) );
  INV_X1 U4910 ( .A(n4011), .ZN(n4015) );
  NAND3_X1 U4911 ( .A1(n3813), .A2(n7036), .A3(n4015), .ZN(n4006) );
  AND2_X1 U4912 ( .A1(n7028), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4075) );
  INV_X1 U4913 ( .A(n5499), .ZN(n5506) );
  NAND2_X1 U4914 ( .A1(n4075), .A2(n5506), .ZN(n7040) );
  NOR2_X1 U4915 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n7163) );
  NAND3_X1 U4916 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n7163), .ZN(n7031) );
  NAND2_X1 U4917 ( .A1(n7040), .A2(n7031), .ZN(n3979) );
  NOR2_X1 U4918 ( .A1(n6803), .A2(n3979), .ZN(n3980) );
  NAND2_X1 U4919 ( .A1(n3998), .A2(n3826), .ZN(n3985) );
  INV_X1 U4920 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5820) );
  INV_X1 U4921 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5134) );
  INV_X1 U4922 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6140) );
  INV_X1 U4923 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5977) );
  INV_X1 U4924 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6124) );
  INV_X1 U4925 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6111) );
  INV_X1 U4926 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6084) );
  INV_X1 U4927 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6077) );
  NOR2_X1 U4928 ( .A1(n5505), .A2(n6077), .ZN(n3982) );
  XNOR2_X1 U4929 ( .A(n3982), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5513)
         );
  NOR2_X1 U4930 ( .A1(n5513), .A2(n3983), .ZN(n3984) );
  NAND2_X1 U4931 ( .A1(n3985), .A2(n6515), .ZN(n6548) );
  INV_X1 U4932 ( .A(n6548), .ZN(n6528) );
  NOR2_X1 U4933 ( .A1(n4373), .A2(n6528), .ZN(n4005) );
  INV_X1 U4934 ( .A(n3465), .ZN(n4021) );
  NAND2_X1 U4935 ( .A1(n3998), .A2(n4021), .ZN(n6545) );
  INV_X1 U4936 ( .A(n6995), .ZN(n4523) );
  NOR2_X1 U4937 ( .A1(n6545), .A2(n4523), .ZN(n4004) );
  NOR2_X1 U4938 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3994) );
  NAND2_X1 U4939 ( .A1(n4097), .A2(n3994), .ZN(n3986) );
  NOR2_X1 U4940 ( .A1(n3987), .A2(n3986), .ZN(n3988) );
  NAND2_X1 U4941 ( .A1(n6507), .A2(n6504), .ZN(n5915) );
  AND2_X1 U4942 ( .A1(n5915), .A2(REIP_REG_0__SCAN_IN), .ZN(n4003) );
  OR2_X1 U4943 ( .A1(n3852), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3990)
         );
  NAND2_X1 U4944 ( .A1(n3990), .A2(n3989), .ZN(n4152) );
  INV_X1 U4945 ( .A(n3994), .ZN(n3991) );
  AND2_X1 U4946 ( .A1(n4097), .A2(n3991), .ZN(n3995) );
  NAND2_X1 U4947 ( .A1(EBX_REG_31__SCAN_IN), .A2(n3998), .ZN(n5923) );
  INV_X1 U4948 ( .A(n5923), .ZN(n3992) );
  AND2_X1 U4949 ( .A1(n3447), .A2(n3992), .ZN(n3993) );
  INV_X1 U4950 ( .A(n7060), .ZN(n4095) );
  NAND2_X1 U4951 ( .A1(n4095), .A2(n3994), .ZN(n7022) );
  NAND2_X1 U4952 ( .A1(n3596), .A2(n7022), .ZN(n5922) );
  INV_X1 U4953 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U4954 ( .A1(n3995), .A2(n6027), .ZN(n3996) );
  NAND2_X1 U4955 ( .A1(n5922), .A2(n3996), .ZN(n3997) );
  NAND2_X1 U4956 ( .A1(n6543), .A2(EBX_REG_0__SCAN_IN), .ZN(n4001) );
  AND2_X1 U4957 ( .A1(n5513), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3999) );
  OAI21_X1 U4958 ( .B1(n6525), .B2(n6518), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4000) );
  OAI211_X1 U4959 ( .C1(n4152), .C2(n6527), .A(n4001), .B(n4000), .ZN(n4002)
         );
  OR4_X1 U4960 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(U2827) );
  INV_X1 U4961 ( .A(n4006), .ZN(n4008) );
  INV_X1 U4962 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n5677) );
  NOR2_X2 U4963 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6923) );
  AND2_X1 U4964 ( .A1(n6923), .A2(n3983), .ZN(n4949) );
  INV_X1 U4965 ( .A(n4949), .ZN(n4007) );
  OAI211_X1 U4966 ( .C1(n4008), .C2(n5677), .A(n4007), .B(n6598), .ZN(U2788)
         );
  OR2_X1 U4967 ( .A1(n4061), .A2(n4040), .ZN(n4014) );
  INV_X1 U4968 ( .A(n4335), .ZN(n4010) );
  OR3_X1 U4969 ( .A1(n4077), .A2(n4010), .A3(n4009), .ZN(n4012) );
  AOI22_X1 U4970 ( .A1(n4012), .A2(n4040), .B1(n3813), .B2(n4011), .ZN(n4013)
         );
  AND2_X1 U4971 ( .A1(n4014), .A2(n4013), .ZN(n6990) );
  NAND2_X1 U4972 ( .A1(n3813), .A2(n4015), .ZN(n4017) );
  NAND2_X1 U4973 ( .A1(n4017), .A2(n4016), .ZN(n4020) );
  INV_X1 U4974 ( .A(n3826), .ZN(n4018) );
  NAND2_X1 U4975 ( .A1(n4040), .A2(n4018), .ZN(n4019) );
  NAND2_X1 U4976 ( .A1(n4020), .A2(n4019), .ZN(n6409) );
  OR2_X1 U4977 ( .A1(n3596), .A2(n4021), .ZN(n4026) );
  AOI21_X1 U4978 ( .B1(n4026), .B2(n7060), .A(READY_N), .ZN(n7161) );
  NOR2_X1 U4979 ( .A1(n6409), .A2(n7161), .ZN(n6987) );
  OR2_X1 U4980 ( .A1(n6987), .A2(n7033), .ZN(n4024) );
  INV_X1 U4981 ( .A(n4024), .ZN(n6416) );
  INV_X1 U4982 ( .A(MORE_REG_SCAN_IN), .ZN(n4022) );
  OR2_X1 U4983 ( .A1(n6416), .A2(n4022), .ZN(n4023) );
  OAI21_X1 U4984 ( .B1(n6990), .B2(n4024), .A(n4023), .ZN(U3471) );
  OAI21_X1 U4985 ( .B1(n4949), .B2(READREQUEST_REG_SCAN_IN), .A(n7157), .ZN(
        n4025) );
  OAI21_X1 U4986 ( .B1(n7157), .B2(n4026), .A(n4025), .ZN(U3474) );
  AND3_X1 U4987 ( .A1(n3761), .A2(n3940), .A3(n3939), .ZN(n4028) );
  AND2_X1 U4988 ( .A1(n3191), .A2(n4028), .ZN(n4031) );
  INV_X1 U4989 ( .A(n4029), .ZN(n4030) );
  NAND2_X1 U4990 ( .A1(n4031), .A2(n4030), .ZN(n6994) );
  NAND2_X1 U4991 ( .A1(n4027), .A2(n6994), .ZN(n4037) );
  INV_X1 U4992 ( .A(n4032), .ZN(n4069) );
  INV_X1 U4993 ( .A(n4033), .ZN(n4194) );
  NAND3_X1 U4994 ( .A1(n6996), .A2(n4069), .A3(n4194), .ZN(n4034) );
  OAI21_X1 U4995 ( .B1(n4182), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4034), 
        .ZN(n4035) );
  INV_X1 U4996 ( .A(n4035), .ZN(n4036) );
  NAND2_X1 U4997 ( .A1(n4037), .A2(n4036), .ZN(n7003) );
  INV_X1 U4998 ( .A(n7147), .ZN(n4072) );
  INV_X1 U4999 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4068) );
  NOR2_X1 U5000 ( .A1(n3983), .A2(n4068), .ZN(n4041) );
  INV_X1 U5001 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U5002 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4038), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6805), .ZN(n4067) );
  AOI222_X1 U5003 ( .A1(n7003), .A2(n4072), .B1(n4041), .B2(n4067), .C1(n4039), 
        .C2(n7026), .ZN(n4059) );
  NOR2_X1 U5004 ( .A1(n4144), .A2(n4095), .ZN(n4042) );
  OAI22_X1 U5005 ( .A1(n4182), .A2(n7060), .B1(n4042), .B2(n3761), .ZN(n4044)
         );
  INV_X1 U5006 ( .A(READY_N), .ZN(n4043) );
  NAND2_X1 U5007 ( .A1(n4044), .A2(n4043), .ZN(n4045) );
  NAND2_X1 U5008 ( .A1(n4045), .A2(n4335), .ZN(n4047) );
  NAND2_X1 U5009 ( .A1(n4047), .A2(n4046), .ZN(n4056) );
  INV_X1 U5010 ( .A(n4048), .ZN(n4049) );
  NOR2_X1 U5011 ( .A1(n3191), .A2(n4049), .ZN(n4331) );
  OAI21_X1 U5012 ( .B1(n3465), .B2(n3439), .A(n4050), .ZN(n4051) );
  NOR2_X1 U5013 ( .A1(n4331), .A2(n4051), .ZN(n4055) );
  INV_X1 U5014 ( .A(n4052), .ZN(n4053) );
  NAND2_X1 U5015 ( .A1(n4054), .A2(n4053), .ZN(n4141) );
  AND3_X1 U5016 ( .A1(n4056), .A2(n4055), .A3(n4141), .ZN(n4188) );
  INV_X1 U5017 ( .A(n4188), .ZN(n7002) );
  NAND2_X1 U5018 ( .A1(n7002), .A2(n7036), .ZN(n6403) );
  NAND2_X1 U5019 ( .A1(n7028), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U5020 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4202) );
  NOR2_X1 U5021 ( .A1(n7028), .A2(n4202), .ZN(n7043) );
  NAND2_X1 U5022 ( .A1(FLUSH_REG_SCAN_IN), .A2(n7043), .ZN(n4057) );
  NAND3_X1 U5023 ( .A1(n6403), .A2(n7137), .A3(n4057), .ZN(n7145) );
  INV_X1 U5024 ( .A(n7145), .ZN(n7140) );
  NOR2_X1 U5025 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6297), .ZN(n7141)
         );
  OAI21_X1 U5026 ( .B1(n7140), .B2(n7141), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4058) );
  OAI21_X1 U5027 ( .B1(n4059), .B2(n7140), .A(n4058), .ZN(U3460) );
  AOI21_X1 U5028 ( .B1(n7026), .B2(n4069), .A(n7140), .ZN(n4074) );
  NAND2_X1 U5029 ( .A1(n4060), .A2(n6994), .ZN(n4066) );
  NAND2_X1 U5030 ( .A1(n4061), .A2(n4335), .ZN(n4185) );
  XNOR2_X1 U5031 ( .A(n4032), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4064)
         );
  MUX2_X1 U5032 ( .A(n3743), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n4062) );
  OAI22_X1 U5033 ( .A1(n4182), .A2(n4062), .B1(n4180), .B2(n4064), .ZN(n4063)
         );
  AOI21_X1 U5034 ( .B1(n4185), .B2(n4064), .A(n4063), .ZN(n4065) );
  NAND2_X1 U5035 ( .A1(n4066), .A2(n4065), .ZN(n4189) );
  NOR3_X1 U5036 ( .A1(n3983), .A2(n4068), .A3(n4067), .ZN(n4071) );
  NOR3_X1 U5037 ( .A1(n4069), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6297), 
        .ZN(n4070) );
  AOI211_X1 U5038 ( .C1(n4189), .C2(n4072), .A(n4071), .B(n4070), .ZN(n4073)
         );
  OAI22_X1 U5039 ( .A1(n4074), .A2(n3187), .B1(n7140), .B2(n4073), .ZN(U3459)
         );
  NAND2_X1 U5040 ( .A1(n4075), .A2(STATEBS16_REG_SCAN_IN), .ZN(n7044) );
  XOR2_X1 U5041 ( .A(n4076), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n4091) );
  NAND2_X1 U5042 ( .A1(n4091), .A2(n6700), .ZN(n4085) );
  NAND2_X1 U5043 ( .A1(n7028), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4079) );
  INV_X1 U5044 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6414) );
  NAND2_X1 U5045 ( .A1(n6414), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4078) );
  AND2_X1 U5046 ( .A1(n4079), .A2(n4078), .ZN(n4227) );
  NAND2_X1 U5047 ( .A1(n6927), .A2(n4080), .ZN(n7159) );
  NAND2_X1 U5048 ( .A1(n7159), .A2(n7028), .ZN(n4081) );
  NAND2_X1 U5049 ( .A1(n4227), .A2(n6162), .ZN(n4083) );
  NAND2_X1 U5050 ( .A1(n6803), .A2(REIP_REG_0__SCAN_IN), .ZN(n4087) );
  INV_X1 U5051 ( .A(n4087), .ZN(n4082) );
  AOI21_X1 U5052 ( .B1(PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4083), .A(n4082), 
        .ZN(n4084) );
  OAI211_X1 U5053 ( .C1(n6679), .C2(n4373), .A(n4085), .B(n4084), .ZN(U2986)
         );
  OAI21_X1 U5054 ( .B1(n5258), .B2(n4086), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4088) );
  OAI211_X1 U5055 ( .C1(n6775), .C2(n4152), .A(n4088), .B(n4087), .ZN(n4090)
         );
  AOI211_X1 U5056 ( .C1(n6801), .C2(n4091), .A(n4090), .B(n4089), .ZN(n4092)
         );
  INV_X1 U5057 ( .A(n4092), .ZN(U3018) );
  INV_X1 U5058 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4099) );
  INV_X1 U5059 ( .A(n7023), .ZN(n4093) );
  INV_X1 U5060 ( .A(n4182), .ZN(n6999) );
  NAND2_X1 U5061 ( .A1(n6999), .A2(n4340), .ZN(n4094) );
  NAND2_X1 U5062 ( .A1(n6660), .A2(n4094), .ZN(n4096) );
  NAND2_X1 U5063 ( .A1(n6590), .A2(n4097), .ZN(n6565) );
  INV_X1 U5064 ( .A(n4202), .ZN(n4171) );
  NAND2_X1 U5065 ( .A1(n7028), .A2(n4171), .ZN(n6570) );
  INV_X1 U5066 ( .A(n6570), .ZN(n6578) );
  NOR2_X4 U5067 ( .A1(n6590), .A2(n7160), .ZN(n6594) );
  AOI22_X1 U5068 ( .A1(n6578), .A2(UWORD_REG_3__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4098) );
  OAI21_X1 U5069 ( .B1(n4099), .B2(n6565), .A(n4098), .ZN(U2904) );
  INV_X1 U5070 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6615) );
  AOI22_X1 U5071 ( .A1(n6578), .A2(UWORD_REG_11__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4100) );
  OAI21_X1 U5072 ( .B1(n6615), .B2(n6565), .A(n4100), .ZN(U2896) );
  INV_X1 U5073 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5074 ( .A1(n6578), .A2(UWORD_REG_7__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4101) );
  OAI21_X1 U5075 ( .B1(n4102), .B2(n6565), .A(n4101), .ZN(U2900) );
  INV_X1 U5076 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5665) );
  AOI22_X1 U5077 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6578), .B1(n6594), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4103) );
  OAI21_X1 U5078 ( .B1(n5665), .B2(n6565), .A(n4103), .ZN(U2907) );
  INV_X1 U5079 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5868) );
  AOI22_X1 U5080 ( .A1(n6578), .A2(UWORD_REG_5__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4104) );
  OAI21_X1 U5081 ( .B1(n5868), .B2(n6565), .A(n4104), .ZN(U2902) );
  INV_X1 U5082 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5083 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6578), .B1(n6594), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4105) );
  OAI21_X1 U5084 ( .B1(n4106), .B2(n6565), .A(n4105), .ZN(U2903) );
  INV_X1 U5085 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5681) );
  AOI22_X1 U5086 ( .A1(n6578), .A2(UWORD_REG_10__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4107) );
  OAI21_X1 U5087 ( .B1(n5681), .B2(n6565), .A(n4107), .ZN(U2897) );
  INV_X1 U5088 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5089 ( .A1(n6578), .A2(UWORD_REG_6__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4108) );
  OAI21_X1 U5090 ( .B1(n4109), .B2(n6565), .A(n4108), .ZN(U2901) );
  INV_X1 U5091 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5092 ( .A1(n6578), .A2(UWORD_REG_8__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4110) );
  OAI21_X1 U5093 ( .B1(n4111), .B2(n6565), .A(n4110), .ZN(U2899) );
  INV_X1 U5094 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6618) );
  AOI22_X1 U5095 ( .A1(n6578), .A2(UWORD_REG_12__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4112) );
  OAI21_X1 U5096 ( .B1(n6618), .B2(n6565), .A(n4112), .ZN(U2895) );
  INV_X1 U5097 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6611) );
  AOI22_X1 U5098 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6578), .B1(n6594), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4113) );
  OAI21_X1 U5099 ( .B1(n6611), .B2(n6565), .A(n4113), .ZN(U2898) );
  INV_X1 U5100 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5850) );
  AOI22_X1 U5101 ( .A1(n7160), .A2(UWORD_REG_2__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4114) );
  OAI21_X1 U5102 ( .B1(n5850), .B2(n6565), .A(n4114), .ZN(U2905) );
  INV_X1 U5103 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5104 ( .A1(n7160), .A2(UWORD_REG_13__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4115) );
  OAI21_X1 U5105 ( .B1(n4116), .B2(n6565), .A(n4115), .ZN(U2894) );
  NAND2_X1 U5106 ( .A1(n3196), .A2(n3972), .ZN(n4121) );
  NAND2_X1 U5107 ( .A1(n5501), .A2(EAX_REG_1__SCAN_IN), .ZN(n4118) );
  NAND2_X1 U5108 ( .A1(n6930), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4117)
         );
  OAI211_X1 U5109 ( .C1(n4218), .C2(n3743), .A(n4118), .B(n4117), .ZN(n4119)
         );
  INV_X1 U5110 ( .A(n4119), .ZN(n4120) );
  NAND2_X1 U5111 ( .A1(n4121), .A2(n4120), .ZN(n4166) );
  NAND2_X1 U5112 ( .A1(n4122), .A2(n5506), .ZN(n4123) );
  NAND2_X1 U5113 ( .A1(n4124), .A2(n4123), .ZN(n4165) );
  NAND2_X1 U5114 ( .A1(n4166), .A2(n4165), .ZN(n4164) );
  OAI21_X1 U5115 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4125), .ZN(n6703) );
  NAND2_X1 U5116 ( .A1(n6703), .A2(n5506), .ZN(n4127) );
  NAND2_X1 U5117 ( .A1(n5509), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4126)
         );
  NAND2_X1 U5118 ( .A1(n4127), .A2(n4126), .ZN(n4128) );
  AOI21_X1 U5119 ( .B1(n5501), .B2(EAX_REG_2__SCAN_IN), .A(n4128), .ZN(n4131)
         );
  INV_X1 U5120 ( .A(n4218), .ZN(n4129) );
  NAND2_X1 U5121 ( .A1(n4129), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4130) );
  AND2_X1 U5122 ( .A1(n4131), .A2(n4130), .ZN(n4133) );
  NAND2_X1 U5123 ( .A1(n4164), .A2(n4133), .ZN(n4139) );
  INV_X1 U5124 ( .A(n3972), .ZN(n4132) );
  INV_X1 U5125 ( .A(n5509), .ZN(n5366) );
  OAI21_X1 U5126 ( .B1(n6284), .B2(n4132), .A(n5366), .ZN(n4138) );
  NAND2_X1 U5127 ( .A1(n4139), .A2(n4138), .ZN(n4137) );
  INV_X1 U5128 ( .A(n4164), .ZN(n4135) );
  INV_X1 U5129 ( .A(n4133), .ZN(n4134) );
  NAND2_X1 U5130 ( .A1(n4135), .A2(n4134), .ZN(n4136) );
  NAND2_X1 U5131 ( .A1(n4137), .A2(n4136), .ZN(n4245) );
  NOR2_X1 U5132 ( .A1(n4139), .A2(n4138), .ZN(n4140) );
  NOR2_X1 U5133 ( .A1(n4245), .A2(n4140), .ZN(n6699) );
  INV_X1 U5134 ( .A(n6699), .ZN(n4641) );
  AND2_X1 U5135 ( .A1(n3476), .A2(n4333), .ZN(n4146) );
  INV_X1 U5136 ( .A(n4142), .ZN(n4145) );
  NOR2_X1 U5137 ( .A1(n3444), .A2(n4143), .ZN(n4332) );
  NAND4_X1 U5138 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4332), .ZN(n4147)
         );
  INV_X2 U5139 ( .A(n6055), .ZN(n6063) );
  AND2_X1 U5140 ( .A1(n6063), .A2(n3444), .ZN(n4592) );
  INV_X2 U5141 ( .A(n4592), .ZN(n6058) );
  AND2_X1 U5142 ( .A1(n6063), .A2(n4149), .ZN(n6056) );
  INV_X2 U5143 ( .A(n6056), .ZN(n6060) );
  INV_X1 U5144 ( .A(n4248), .ZN(n4150) );
  XNOR2_X1 U5145 ( .A(n4249), .B(n4150), .ZN(n6798) );
  INV_X1 U5146 ( .A(n6798), .ZN(n4151) );
  INV_X1 U5147 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5816) );
  OAI222_X1 U5148 ( .A1(n4641), .A2(n6058), .B1(n6060), .B2(n4151), .C1(n6063), 
        .C2(n5816), .ZN(U2857) );
  OAI222_X1 U5149 ( .A1(n4373), .A2(n6058), .B1(n6063), .B2(n3835), .C1(n4152), 
        .C2(n6060), .ZN(U2859) );
  XOR2_X1 U5150 ( .A(n4154), .B(n4153), .Z(n4226) );
  INV_X1 U5151 ( .A(n4226), .ZN(n4163) );
  INV_X1 U5152 ( .A(n6745), .ZN(n4159) );
  INV_X1 U5153 ( .A(REIP_REG_1__SCAN_IN), .ZN(n7074) );
  NOR2_X1 U5154 ( .A1(n6774), .A2(n7074), .ZN(n4230) );
  INV_X1 U5155 ( .A(n5029), .ZN(n4157) );
  INV_X1 U5156 ( .A(n4155), .ZN(n4156) );
  AOI21_X1 U5157 ( .B1(n4157), .B2(n5526), .A(n4156), .ZN(n4168) );
  NOR2_X1 U5158 ( .A1(n6775), .A2(n4168), .ZN(n4158) );
  AOI211_X1 U5159 ( .C1(INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n4159), .A(n4230), 
        .B(n4158), .ZN(n4162) );
  NAND3_X1 U5160 ( .A1(n6750), .A2(n6805), .A3(n4160), .ZN(n4161) );
  OAI211_X1 U5161 ( .C1(n4163), .C2(n6773), .A(n4162), .B(n4161), .ZN(U3017)
         );
  OAI21_X1 U5162 ( .B1(n4166), .B2(n4165), .A(n4164), .ZN(n5038) );
  OAI22_X1 U5163 ( .A1(n6060), .A2(n4168), .B1(n4167), .B2(n6063), .ZN(n4169)
         );
  INV_X1 U5164 ( .A(n4169), .ZN(n4170) );
  OAI21_X1 U5165 ( .B1(n5038), .B2(n6058), .A(n4170), .ZN(U2858) );
  INV_X1 U5166 ( .A(n4600), .ZN(n4382) );
  NOR2_X1 U5167 ( .A1(n3983), .A2(FLUSH_REG_SCAN_IN), .ZN(n4197) );
  INV_X1 U5168 ( .A(n4197), .ZN(n4193) );
  INV_X1 U5169 ( .A(n4172), .ZN(n4192) );
  NAND2_X1 U5170 ( .A1(n4173), .A2(n6994), .ZN(n4187) );
  MUX2_X1 U5171 ( .A(n4174), .B(n6301), .S(n4032), .Z(n4175) );
  NOR2_X1 U5172 ( .A1(n4175), .A2(n4172), .ZN(n4184) );
  NAND2_X1 U5173 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4177) );
  INV_X1 U5174 ( .A(n4177), .ZN(n4176) );
  MUX2_X1 U5175 ( .A(n4177), .B(n4176), .S(n6301), .Z(n4181) );
  NAND2_X1 U5176 ( .A1(n4032), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4178) );
  NAND2_X1 U5177 ( .A1(n4178), .A2(n3298), .ZN(n4179) );
  NAND2_X1 U5178 ( .A1(n3581), .A2(n4179), .ZN(n6298) );
  OAI22_X1 U5179 ( .A1(n4182), .A2(n4181), .B1(n4180), .B2(n6298), .ZN(n4183)
         );
  AOI21_X1 U5180 ( .B1(n4185), .B2(n4184), .A(n4183), .ZN(n4186) );
  NAND2_X1 U5181 ( .A1(n4187), .A2(n4186), .ZN(n6296) );
  MUX2_X1 U5182 ( .A(n6296), .B(n6301), .S(n4188), .Z(n7017) );
  MUX2_X1 U5183 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4189), .S(n7002), 
        .Z(n7011) );
  NAND3_X1 U5184 ( .A1(n7017), .A2(n3983), .A3(n7011), .ZN(n4191) );
  OAI21_X1 U5185 ( .B1(n4193), .B2(n4192), .A(n4191), .ZN(n6992) );
  NAND2_X1 U5186 ( .A1(n6992), .A2(n4194), .ZN(n4200) );
  NOR2_X1 U5187 ( .A1(n4195), .A2(n3283), .ZN(n4196) );
  XNOR2_X1 U5188 ( .A(n4196), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6402)
         );
  OAI22_X1 U5189 ( .A1(n6402), .A2(n3191), .B1(n6407), .B2(n7002), .ZN(n4199)
         );
  AND2_X1 U5190 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4197), .ZN(n4198)
         );
  AOI21_X1 U5191 ( .B1(n4199), .B2(n3983), .A(n4198), .ZN(n6991) );
  NAND2_X1 U5192 ( .A1(n4200), .A2(n6991), .ZN(n4203) );
  OAI21_X1 U5193 ( .B1(n4203), .B2(FLUSH_REG_SCAN_IN), .A(n7043), .ZN(n4201)
         );
  NAND2_X1 U5194 ( .A1(n4600), .A2(n4201), .ZN(n6810) );
  NOR2_X1 U5195 ( .A1(n4203), .A2(n4202), .ZN(n7027) );
  AND2_X1 U5196 ( .A1(n3454), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6292) );
  OAI22_X1 U5197 ( .A1(n6817), .A2(n6927), .B1(n4523), .B2(n6292), .ZN(n4204)
         );
  OAI21_X1 U5198 ( .B1(n7027), .B2(n4204), .A(n6810), .ZN(n4205) );
  OAI21_X1 U5199 ( .B1(n6810), .B2(n7000), .A(n4205), .ZN(U3465) );
  AND2_X1 U5200 ( .A1(n4250), .A2(n4206), .ZN(n4207) );
  OR2_X1 U5201 ( .A1(n4207), .A2(n4234), .ZN(n6776) );
  INV_X1 U5202 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U5203 ( .A1(n4208), .A2(n3972), .ZN(n4214) );
  OAI21_X1 U5204 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4209), .A(n4219), 
        .ZN(n6693) );
  AOI22_X1 U5205 ( .A1(n6693), .A2(n5506), .B1(n5509), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4211) );
  NAND2_X1 U5206 ( .A1(n5501), .A2(EAX_REG_3__SCAN_IN), .ZN(n4210) );
  OAI211_X1 U5207 ( .C1(n4218), .C2(n3298), .A(n4211), .B(n4210), .ZN(n4212)
         );
  INV_X1 U5208 ( .A(n4212), .ZN(n4213) );
  NAND2_X1 U5209 ( .A1(n4214), .A2(n4213), .ZN(n4246) );
  NAND2_X1 U5210 ( .A1(n4215), .A2(n3972), .ZN(n4223) );
  NAND2_X1 U5211 ( .A1(n6930), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4217)
         );
  NAND2_X1 U5212 ( .A1(n5501), .A2(EAX_REG_4__SCAN_IN), .ZN(n4216) );
  OAI211_X1 U5213 ( .C1(n4218), .C2(n6407), .A(n4217), .B(n4216), .ZN(n4221)
         );
  AOI21_X1 U5214 ( .B1(n4219), .B2(n5013), .A(n4237), .ZN(n5007) );
  NOR2_X1 U5215 ( .A1(n5007), .A2(n5499), .ZN(n4220) );
  AOI21_X1 U5216 ( .B1(n4221), .B2(n5499), .A(n4220), .ZN(n4222) );
  NAND2_X1 U5217 ( .A1(n4223), .A2(n4222), .ZN(n4224) );
  AND3_X2 U5218 ( .A1(n4245), .A2(n4246), .A3(n4224), .ZN(n4329) );
  AOI21_X1 U5219 ( .B1(n4245), .B2(n4246), .A(n4224), .ZN(n4225) );
  OR2_X1 U5220 ( .A1(n4329), .A2(n4225), .ZN(n4371) );
  OAI222_X1 U5221 ( .A1(n6776), .A2(n6060), .B1(n6063), .B2(n5832), .C1(n6058), 
        .C2(n4371), .ZN(U2855) );
  NAND2_X1 U5222 ( .A1(n4226), .A2(n6700), .ZN(n4232) );
  INV_X1 U5223 ( .A(n4227), .ZN(n4228) );
  NOR2_X1 U5224 ( .A1(n6704), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4229)
         );
  AOI211_X1 U5225 ( .C1(n6694), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4230), 
        .B(n4229), .ZN(n4231) );
  OAI211_X1 U5226 ( .C1(n6679), .C2(n5038), .A(n4232), .B(n4231), .ZN(U2985)
         );
  OR2_X1 U5227 ( .A1(n4234), .A2(n4233), .ZN(n4235) );
  NAND2_X1 U5228 ( .A1(n4316), .A2(n4235), .ZN(n6765) );
  NAND2_X1 U5229 ( .A1(n4236), .A2(n3972), .ZN(n4243) );
  INV_X1 U5230 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4240) );
  OAI21_X1 U5231 ( .B1(n4237), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4320), 
        .ZN(n6685) );
  NAND2_X1 U5232 ( .A1(n6685), .A2(n5506), .ZN(n4239) );
  NAND2_X1 U5233 ( .A1(n5509), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4238)
         );
  OAI211_X1 U5234 ( .C1(n5369), .C2(n4240), .A(n4239), .B(n4238), .ZN(n4241)
         );
  INV_X1 U5235 ( .A(n4241), .ZN(n4242) );
  XNOR2_X1 U5236 ( .A(n4329), .B(n4328), .ZN(n6680) );
  INV_X1 U5237 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4244) );
  OAI222_X1 U5238 ( .A1(n6765), .A2(n6060), .B1(n6058), .B2(n6680), .C1(n6063), 
        .C2(n4244), .ZN(U2854) );
  XOR2_X1 U5239 ( .A(n4246), .B(n4245), .Z(n6690) );
  INV_X1 U5240 ( .A(n6690), .ZN(n4372) );
  OAI21_X1 U5241 ( .B1(n4249), .B2(n4248), .A(n4247), .ZN(n4251) );
  AND2_X1 U5242 ( .A1(n4251), .A2(n4250), .ZN(n6786) );
  AOI22_X1 U5243 ( .A1(n6056), .A2(n6786), .B1(n6055), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4252) );
  OAI21_X1 U5244 ( .B1(n4372), .B2(n6058), .A(n4252), .ZN(U2856) );
  OAI21_X1 U5245 ( .B1(n4255), .B2(n4254), .A(n4253), .ZN(n6772) );
  INV_X1 U5246 ( .A(n4371), .ZN(n5016) );
  INV_X2 U5247 ( .A(n6679), .ZN(n6698) );
  INV_X1 U5248 ( .A(n5007), .ZN(n4257) );
  AOI22_X1 U5249 ( .A1(n6694), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6785), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4256) );
  OAI21_X1 U5250 ( .B1(n4257), .B2(n6704), .A(n4256), .ZN(n4258) );
  AOI21_X1 U5251 ( .B1(n5016), .B2(n6698), .A(n4258), .ZN(n4259) );
  OAI21_X1 U5252 ( .B1(n6681), .B2(n6772), .A(n4259), .ZN(U2982) );
  INV_X1 U5253 ( .A(n4027), .ZN(n6281) );
  INV_X1 U5254 ( .A(n4842), .ZN(n4260) );
  NOR2_X1 U5255 ( .A1(n4260), .A2(n6927), .ZN(n4850) );
  INV_X1 U5256 ( .A(n4173), .ZN(n6546) );
  INV_X1 U5257 ( .A(n4261), .ZN(n4596) );
  INV_X1 U5258 ( .A(n4595), .ZN(n5062) );
  NOR2_X1 U5259 ( .A1(n4596), .A2(n5062), .ZN(n4760) );
  AND2_X1 U5260 ( .A1(n4262), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4849) );
  AOI22_X1 U5261 ( .A1(n4850), .A2(n6546), .B1(n4760), .B2(n4849), .ZN(n4301)
         );
  INV_X1 U5262 ( .A(DATAI_2_), .ZN(n6626) );
  NOR2_X1 U5263 ( .A1(n6626), .A2(n4600), .ZN(n6946) );
  INV_X1 U5264 ( .A(n6946), .ZN(n4877) );
  NAND3_X1 U5265 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7016), .A3(n7005), .ZN(n6819) );
  OR2_X1 U5266 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6819), .ZN(n4296)
         );
  NOR2_X1 U5267 ( .A1(n4262), .A2(n6930), .ZN(n4594) );
  OAI21_X1 U5268 ( .B1(n4760), .B2(n6930), .A(n4382), .ZN(n4756) );
  AOI211_X1 U5269 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4296), .A(n4594), .B(
        n4756), .ZN(n4267) );
  AND2_X1 U5270 ( .A1(n6923), .A2(n6414), .ZN(n4806) );
  INV_X1 U5271 ( .A(n4208), .ZN(n6294) );
  AND3_X1 U5272 ( .A1(n6284), .A2(n4836), .A3(n3196), .ZN(n4264) );
  NAND2_X1 U5273 ( .A1(n6294), .A2(n4264), .ZN(n4554) );
  NOR2_X1 U5274 ( .A1(n6284), .A2(n4376), .ZN(n6291) );
  NAND2_X1 U5275 ( .A1(n6291), .A2(n4751), .ZN(n6818) );
  OR2_X1 U5276 ( .A1(n6818), .A2(n6414), .ZN(n4265) );
  NAND2_X1 U5277 ( .A1(n4842), .A2(n3283), .ZN(n6812) );
  OAI211_X1 U5278 ( .C1(n4806), .C2(n4554), .A(n6811), .B(n6812), .ZN(n4266)
         );
  NAND2_X1 U5279 ( .A1(n4267), .A2(n4266), .ZN(n4293) );
  NAND2_X1 U5280 ( .A1(n4293), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4272) );
  NAND2_X1 U5281 ( .A1(n6698), .A2(DATAI_26_), .ZN(n6949) );
  INV_X1 U5282 ( .A(n6949), .ZN(n6872) );
  INV_X1 U5283 ( .A(n7137), .ZN(n4269) );
  NAND2_X1 U5284 ( .A1(n4295), .A2(n3439), .ZN(n4816) );
  NAND2_X1 U5285 ( .A1(n6698), .A2(DATAI_18_), .ZN(n6875) );
  OR2_X1 U5286 ( .A1(n6818), .A2(n4836), .ZN(n6822) );
  OAI22_X1 U5287 ( .A1(n4816), .A2(n4296), .B1(n6875), .B2(n6822), .ZN(n4270)
         );
  AOI21_X1 U5288 ( .B1(n6872), .B2(n4298), .A(n4270), .ZN(n4271) );
  OAI211_X1 U5289 ( .C1(n4301), .C2(n4877), .A(n4272), .B(n4271), .ZN(U3054)
         );
  INV_X1 U5290 ( .A(DATAI_1_), .ZN(n6624) );
  NOR2_X1 U5291 ( .A1(n6624), .A2(n4600), .ZN(n6940) );
  INV_X1 U5292 ( .A(n6940), .ZN(n4857) );
  NAND2_X1 U5293 ( .A1(n4293), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U5294 ( .A1(n6698), .A2(DATAI_25_), .ZN(n6943) );
  INV_X1 U5295 ( .A(n6943), .ZN(n6868) );
  NAND2_X1 U5296 ( .A1(n4295), .A2(n3447), .ZN(n4802) );
  NAND2_X1 U5297 ( .A1(n6698), .A2(DATAI_17_), .ZN(n6871) );
  OAI22_X1 U5298 ( .A1(n4802), .A2(n4296), .B1(n6871), .B2(n6822), .ZN(n4273)
         );
  AOI21_X1 U5299 ( .B1(n6868), .B2(n4298), .A(n4273), .ZN(n4274) );
  OAI211_X1 U5300 ( .C1(n4301), .C2(n4857), .A(n4275), .B(n4274), .ZN(U3053)
         );
  INV_X1 U5301 ( .A(DATAI_0_), .ZN(n6622) );
  NOR2_X1 U5302 ( .A1(n6622), .A2(n4600), .ZN(n6934) );
  INV_X1 U5303 ( .A(n6934), .ZN(n4852) );
  NAND2_X1 U5304 ( .A1(n4293), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4278) );
  NAND2_X1 U5305 ( .A1(n6698), .A2(DATAI_24_), .ZN(n6937) );
  INV_X1 U5306 ( .A(n6937), .ZN(n6864) );
  NAND2_X1 U5307 ( .A1(n4295), .A2(n4097), .ZN(n4812) );
  NAND2_X1 U5308 ( .A1(n6698), .A2(DATAI_16_), .ZN(n6867) );
  OAI22_X1 U5309 ( .A1(n4812), .A2(n4296), .B1(n6867), .B2(n6822), .ZN(n4276)
         );
  AOI21_X1 U5310 ( .B1(n6864), .B2(n4298), .A(n4276), .ZN(n4277) );
  OAI211_X1 U5311 ( .C1(n4301), .C2(n4852), .A(n4278), .B(n4277), .ZN(U3052)
         );
  INV_X1 U5312 ( .A(DATAI_5_), .ZN(n6632) );
  NOR2_X1 U5313 ( .A1(n6632), .A2(n4600), .ZN(n6964) );
  INV_X1 U5314 ( .A(n6964), .ZN(n4889) );
  NAND2_X1 U5315 ( .A1(n4293), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4282) );
  NAND2_X1 U5316 ( .A1(n6698), .A2(DATAI_29_), .ZN(n6967) );
  INV_X1 U5317 ( .A(n6967), .ZN(n6880) );
  NAND2_X1 U5318 ( .A1(n4295), .A2(n4279), .ZN(n4820) );
  NAND2_X1 U5319 ( .A1(n6698), .A2(DATAI_21_), .ZN(n6883) );
  OAI22_X1 U5320 ( .A1(n4820), .A2(n4296), .B1(n6883), .B2(n6822), .ZN(n4280)
         );
  AOI21_X1 U5321 ( .B1(n6880), .B2(n4298), .A(n4280), .ZN(n4281) );
  OAI211_X1 U5322 ( .C1(n4301), .C2(n4889), .A(n4282), .B(n4281), .ZN(U3057)
         );
  INV_X1 U5323 ( .A(DATAI_6_), .ZN(n6634) );
  NOR2_X1 U5324 ( .A1(n6634), .A2(n4600), .ZN(n6971) );
  INV_X1 U5325 ( .A(n6971), .ZN(n4913) );
  NAND2_X1 U5326 ( .A1(n4293), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4285) );
  INV_X1 U5327 ( .A(DATAI_30_), .ZN(n5896) );
  NAND2_X1 U5328 ( .A1(n4295), .A2(n3184), .ZN(n4905) );
  NAND2_X1 U5329 ( .A1(n6698), .A2(DATAI_22_), .ZN(n6975) );
  OAI22_X1 U5330 ( .A1(n4905), .A2(n4296), .B1(n6975), .B2(n6822), .ZN(n4283)
         );
  AOI21_X1 U5331 ( .B1(n6968), .B2(n4298), .A(n4283), .ZN(n4284) );
  OAI211_X1 U5332 ( .C1(n4301), .C2(n4913), .A(n4285), .B(n4284), .ZN(U3058)
         );
  INV_X1 U5333 ( .A(DATAI_7_), .ZN(n6636) );
  NOR2_X1 U5334 ( .A1(n6636), .A2(n4600), .ZN(n6981) );
  INV_X1 U5335 ( .A(n6981), .ZN(n4867) );
  NAND2_X1 U5336 ( .A1(n4293), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4288) );
  NAND2_X1 U5337 ( .A1(n6698), .A2(DATAI_31_), .ZN(n6986) );
  INV_X1 U5338 ( .A(n6986), .ZN(n6889) );
  NAND2_X1 U5339 ( .A1(n4295), .A2(n3444), .ZN(n4824) );
  NAND2_X1 U5340 ( .A1(n6698), .A2(DATAI_23_), .ZN(n6893) );
  OAI22_X1 U5341 ( .A1(n4824), .A2(n4296), .B1(n6893), .B2(n6822), .ZN(n4286)
         );
  AOI21_X1 U5342 ( .B1(n6889), .B2(n4298), .A(n4286), .ZN(n4287) );
  OAI211_X1 U5343 ( .C1(n4301), .C2(n4867), .A(n4288), .B(n4287), .ZN(U3059)
         );
  INV_X1 U5344 ( .A(DATAI_3_), .ZN(n6628) );
  NOR2_X1 U5345 ( .A1(n6628), .A2(n4600), .ZN(n6952) );
  INV_X1 U5346 ( .A(n6952), .ZN(n4862) );
  NAND2_X1 U5347 ( .A1(n4293), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4292) );
  NAND2_X1 U5348 ( .A1(n6698), .A2(DATAI_27_), .ZN(n6904) );
  INV_X1 U5349 ( .A(n6904), .ZN(n6950) );
  NAND2_X1 U5350 ( .A1(n4295), .A2(n4289), .ZN(n4828) );
  NAND2_X1 U5351 ( .A1(n6698), .A2(DATAI_19_), .ZN(n6955) );
  OAI22_X1 U5352 ( .A1(n4828), .A2(n4296), .B1(n6955), .B2(n6822), .ZN(n4290)
         );
  AOI21_X1 U5353 ( .B1(n6950), .B2(n4298), .A(n4290), .ZN(n4291) );
  OAI211_X1 U5354 ( .C1(n4301), .C2(n4862), .A(n4292), .B(n4291), .ZN(U3055)
         );
  INV_X1 U5355 ( .A(DATAI_4_), .ZN(n6630) );
  NOR2_X1 U5356 ( .A1(n6630), .A2(n4600), .ZN(n6958) );
  INV_X1 U5357 ( .A(n6958), .ZN(n4872) );
  NAND2_X1 U5358 ( .A1(n4293), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4300) );
  NAND2_X1 U5359 ( .A1(n6698), .A2(DATAI_28_), .ZN(n6908) );
  INV_X1 U5360 ( .A(n6908), .ZN(n6956) );
  NAND2_X1 U5361 ( .A1(n4295), .A2(n4294), .ZN(n4832) );
  NAND2_X1 U5362 ( .A1(n6698), .A2(DATAI_20_), .ZN(n6961) );
  OAI22_X1 U5363 ( .A1(n4832), .A2(n4296), .B1(n6961), .B2(n6822), .ZN(n4297)
         );
  AOI21_X1 U5364 ( .B1(n6956), .B2(n4298), .A(n4297), .ZN(n4299) );
  OAI211_X1 U5365 ( .C1(n4301), .C2(n4872), .A(n4300), .B(n4299), .ZN(U3056)
         );
  OR2_X1 U5366 ( .A1(n6291), .A2(n6927), .ZN(n4302) );
  NAND2_X1 U5367 ( .A1(n3196), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6288) );
  NAND2_X1 U5368 ( .A1(n6288), .A2(n6923), .ZN(n6921) );
  NAND2_X1 U5369 ( .A1(n4302), .A2(n6921), .ZN(n4307) );
  AND2_X1 U5370 ( .A1(n4060), .A2(n4027), .ZN(n4798) );
  AND2_X1 U5371 ( .A1(n4798), .A2(n3283), .ZN(n6857) );
  INV_X1 U5372 ( .A(n4309), .ZN(n6912) );
  AOI21_X1 U5373 ( .B1(n6857), .B2(n6995), .A(n6912), .ZN(n4306) );
  INV_X1 U5374 ( .A(n4306), .ZN(n4303) );
  NAND2_X1 U5375 ( .A1(n4307), .A2(n4303), .ZN(n4305) );
  NAND2_X1 U5376 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6855), .ZN(n4304) );
  NAND2_X1 U5377 ( .A1(n4305), .A2(n4304), .ZN(n6913) );
  INV_X1 U5378 ( .A(n6913), .ZN(n4314) );
  AOI21_X1 U5379 ( .B1(n7000), .B2(STATE2_REG_3__SCAN_IN), .A(n4600), .ZN(
        n6814) );
  NAND2_X1 U5380 ( .A1(n4307), .A2(n4306), .ZN(n4308) );
  OAI211_X1 U5381 ( .C1(n6855), .C2(n6923), .A(n6814), .B(n4308), .ZN(n6914)
         );
  NAND2_X1 U5382 ( .A1(n6914), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4313) );
  INV_X1 U5383 ( .A(n6917), .ZN(n4311) );
  NAND3_X1 U5384 ( .A1(n6291), .A2(n4836), .A3(n3196), .ZN(n6894) );
  OAI22_X1 U5385 ( .A1(n4905), .A2(n4309), .B1(n6975), .B2(n6894), .ZN(n4310)
         );
  AOI21_X1 U5386 ( .B1(n6968), .B2(n4311), .A(n4310), .ZN(n4312) );
  OAI211_X1 U5387 ( .C1(n4314), .C2(n4913), .A(n4313), .B(n4312), .ZN(U3082)
         );
  NAND2_X1 U5388 ( .A1(n4316), .A2(n4315), .ZN(n4317) );
  NAND2_X1 U5389 ( .A1(n4447), .A2(n4317), .ZN(n6752) );
  INV_X1 U5390 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U5391 ( .A1(n4318), .A2(n3972), .ZN(n4326) );
  AOI21_X1 U5392 ( .B1(n4320), .B2(n4319), .A(n4414), .ZN(n6519) );
  NAND2_X1 U5393 ( .A1(n6519), .A2(n5506), .ZN(n4324) );
  INV_X1 U5394 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4322) );
  OAI21_X1 U5395 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6414), .A(n6930), 
        .ZN(n4321) );
  OAI21_X1 U5396 ( .B1(n5369), .B2(n4322), .A(n4321), .ZN(n4323) );
  NAND2_X1 U5397 ( .A1(n4324), .A2(n4323), .ZN(n4325) );
  NAND2_X1 U5398 ( .A1(n4326), .A2(n4325), .ZN(n4327) );
  AOI21_X1 U5399 ( .B1(n4329), .B2(n4328), .A(n4327), .ZN(n4330) );
  OR2_X1 U5400 ( .A1(n4503), .A2(n4330), .ZN(n6516) );
  OAI222_X1 U5401 ( .A1(n6752), .A2(n6060), .B1(n6063), .B2(n6523), .C1(n6058), 
        .C2(n6516), .ZN(U2853) );
  NAND2_X1 U5402 ( .A1(n4331), .A2(n7036), .ZN(n4342) );
  NAND3_X1 U5403 ( .A1(n4333), .A2(n4332), .A3(n3184), .ZN(n4334) );
  OAI22_X1 U5404 ( .A1(n4336), .A2(n4335), .B1(n3939), .B2(n4334), .ZN(n4337)
         );
  INV_X1 U5405 ( .A(n4337), .ZN(n4341) );
  NOR2_X1 U5406 ( .A1(n4338), .A2(n5526), .ZN(n4339) );
  NAND2_X2 U5407 ( .A1(n4340), .A2(n4339), .ZN(n6656) );
  NAND2_X1 U5408 ( .A1(n3452), .A2(n3444), .ZN(n4343) );
  AND2_X1 U5409 ( .A1(n6064), .A2(n3295), .ZN(n6558) );
  AND2_X1 U5410 ( .A1(n3430), .A2(n3444), .ZN(n4344) );
  AOI22_X1 U5411 ( .A1(n5004), .A2(DATAI_2_), .B1(EAX_REG_2__SCAN_IN), .B2(
        n6561), .ZN(n4345) );
  OAI21_X1 U5412 ( .B1(n4641), .B2(n6345), .A(n4345), .ZN(U2889) );
  NOR2_X1 U5413 ( .A1(n3196), .A2(n6414), .ZN(n4346) );
  AOI21_X1 U5414 ( .B1(n4838), .B2(n4346), .A(n6927), .ZN(n4348) );
  AND2_X1 U5415 ( .A1(n4173), .A2(n6995), .ZN(n4799) );
  NAND3_X1 U5416 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n7010), .A3(n7005), .ZN(n4598) );
  NOR2_X1 U5417 ( .A1(n7000), .A2(n4598), .ZN(n4368) );
  AOI21_X1 U5418 ( .B1(n4799), .B2(n3293), .A(n4368), .ZN(n4350) );
  AOI22_X1 U5419 ( .A1(n4348), .A2(n4350), .B1(n6927), .B2(n4598), .ZN(n4347)
         );
  NAND2_X1 U5420 ( .A1(n6814), .A2(n4347), .ZN(n4367) );
  INV_X1 U5421 ( .A(n4348), .ZN(n4349) );
  OAI22_X1 U5422 ( .A1(n4350), .A2(n4349), .B1(n6930), .B2(n4598), .ZN(n4366)
         );
  AOI22_X1 U5423 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4367), .B1(n6934), 
        .B2(n4366), .ZN(n4353) );
  NAND2_X1 U5424 ( .A1(n4351), .A2(n4836), .ZN(n4450) );
  INV_X1 U5425 ( .A(n6867), .ZN(n6919) );
  AOI22_X1 U5426 ( .A1(n6920), .A2(n4368), .B1(n4482), .B2(n6919), .ZN(n4352)
         );
  OAI211_X1 U5427 ( .C1(n6937), .C2(n4632), .A(n4353), .B(n4352), .ZN(U3092)
         );
  AOI22_X1 U5428 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4367), .B1(n6981), 
        .B2(n4366), .ZN(n4355) );
  INV_X1 U5429 ( .A(n6893), .ZN(n6977) );
  AOI22_X1 U5430 ( .A1(n6979), .A2(n4368), .B1(n4482), .B2(n6977), .ZN(n4354)
         );
  OAI211_X1 U5431 ( .C1(n6986), .C2(n4632), .A(n4355), .B(n4354), .ZN(U3099)
         );
  AOI22_X1 U5432 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4367), .B1(n6946), 
        .B2(n4366), .ZN(n4357) );
  INV_X1 U5433 ( .A(n6875), .ZN(n6944) );
  AOI22_X1 U5434 ( .A1(n6945), .A2(n4368), .B1(n4482), .B2(n6944), .ZN(n4356)
         );
  OAI211_X1 U5435 ( .C1(n6949), .C2(n4632), .A(n4357), .B(n4356), .ZN(U3094)
         );
  AOI22_X1 U5436 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4367), .B1(n6940), 
        .B2(n4366), .ZN(n4359) );
  INV_X1 U5437 ( .A(n6871), .ZN(n6938) );
  AOI22_X1 U5438 ( .A1(n6939), .A2(n4368), .B1(n4482), .B2(n6938), .ZN(n4358)
         );
  OAI211_X1 U5439 ( .C1(n6943), .C2(n4632), .A(n4359), .B(n4358), .ZN(U3093)
         );
  AOI22_X1 U5440 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4367), .B1(n6952), 
        .B2(n4366), .ZN(n4361) );
  INV_X1 U5441 ( .A(n6955), .ZN(n6901) );
  AOI22_X1 U5442 ( .A1(n6951), .A2(n4368), .B1(n4482), .B2(n6901), .ZN(n4360)
         );
  OAI211_X1 U5443 ( .C1(n6904), .C2(n4632), .A(n4361), .B(n4360), .ZN(U3095)
         );
  AOI22_X1 U5444 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4367), .B1(n6964), 
        .B2(n4366), .ZN(n4363) );
  INV_X1 U5445 ( .A(n6883), .ZN(n6962) );
  AOI22_X1 U5446 ( .A1(n6963), .A2(n4368), .B1(n4482), .B2(n6962), .ZN(n4362)
         );
  OAI211_X1 U5447 ( .C1(n6967), .C2(n4632), .A(n4363), .B(n4362), .ZN(U3097)
         );
  AOI22_X1 U5448 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4367), .B1(n6958), 
        .B2(n4366), .ZN(n4365) );
  INV_X1 U5449 ( .A(n6961), .ZN(n6905) );
  AOI22_X1 U5450 ( .A1(n6957), .A2(n4368), .B1(n4482), .B2(n6905), .ZN(n4364)
         );
  OAI211_X1 U5451 ( .C1(n6908), .C2(n4632), .A(n4365), .B(n4364), .ZN(U3096)
         );
  INV_X1 U5452 ( .A(n6968), .ZN(n4932) );
  AOI22_X1 U5453 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4367), .B1(n6971), 
        .B2(n4366), .ZN(n4370) );
  INV_X1 U5454 ( .A(n6975), .ZN(n6841) );
  AOI22_X1 U5455 ( .A1(n6970), .A2(n4368), .B1(n4482), .B2(n6841), .ZN(n4369)
         );
  OAI211_X1 U5456 ( .C1(n4932), .C2(n4632), .A(n4370), .B(n4369), .ZN(U3098)
         );
  INV_X1 U5457 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6593) );
  OAI222_X1 U5458 ( .A1(n5038), .A2(n6345), .B1(n5048), .B2(n6624), .C1(n6064), 
        .C2(n6593), .ZN(U2890) );
  INV_X1 U5459 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6587) );
  OAI222_X1 U5460 ( .A1(n4371), .A2(n6345), .B1(n5048), .B2(n6630), .C1(n6064), 
        .C2(n6587), .ZN(U2887) );
  INV_X1 U5461 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6589) );
  OAI222_X1 U5462 ( .A1(n4372), .A2(n6345), .B1(n5048), .B2(n6628), .C1(n6064), 
        .C2(n6589), .ZN(U2888) );
  INV_X1 U5463 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6597) );
  OAI222_X1 U5464 ( .A1(n4373), .A2(n6345), .B1(n5048), .B2(n6622), .C1(n6064), 
        .C2(n6597), .ZN(U2891) );
  OAI222_X1 U5465 ( .A1(n6516), .A2(n6345), .B1(n5048), .B2(n6634), .C1(n6064), 
        .C2(n4322), .ZN(U2885) );
  NAND2_X1 U5466 ( .A1(n4798), .A2(n6923), .ZN(n6854) );
  INV_X1 U5467 ( .A(n6854), .ZN(n4374) );
  NOR2_X1 U5468 ( .A1(n4595), .A2(n7016), .ZN(n4452) );
  AOI22_X1 U5469 ( .A1(n4374), .A2(n4173), .B1(n4849), .B2(n4452), .ZN(n4412)
         );
  INV_X1 U5470 ( .A(n4809), .ZN(n4375) );
  NOR2_X1 U5471 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4375), .ZN(n4385)
         );
  INV_X1 U5472 ( .A(n4798), .ZN(n4380) );
  INV_X1 U5473 ( .A(n4376), .ZN(n4377) );
  INV_X1 U5474 ( .A(n4445), .ZN(n4378) );
  OAI21_X1 U5475 ( .B1(n4378), .B2(n4909), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4379) );
  NAND3_X1 U5476 ( .A1(n4380), .A2(n6923), .A3(n4379), .ZN(n4384) );
  NAND2_X1 U5477 ( .A1(n4595), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4381) );
  NAND2_X1 U5478 ( .A1(n4382), .A2(n4381), .ZN(n6863) );
  NOR3_X1 U5479 ( .A1(n6863), .A2(n7016), .A3(n4594), .ZN(n4383) );
  OAI211_X1 U5480 ( .C1(n3454), .C2(n4385), .A(n4384), .B(n4383), .ZN(n4407)
         );
  NAND2_X1 U5481 ( .A1(n4407), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4388)
         );
  INV_X1 U5482 ( .A(n4385), .ZN(n4408) );
  OAI22_X1 U5483 ( .A1(n4812), .A2(n4408), .B1(n6937), .B2(n4445), .ZN(n4386)
         );
  AOI21_X1 U5484 ( .B1(n6919), .B2(n4909), .A(n4386), .ZN(n4387) );
  OAI211_X1 U5485 ( .C1(n4412), .C2(n4852), .A(n4388), .B(n4387), .ZN(U3132)
         );
  NAND2_X1 U5486 ( .A1(n4407), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4391)
         );
  OAI22_X1 U5487 ( .A1(n4824), .A2(n4408), .B1(n6986), .B2(n4445), .ZN(n4389)
         );
  AOI21_X1 U5488 ( .B1(n6977), .B2(n4909), .A(n4389), .ZN(n4390) );
  OAI211_X1 U5489 ( .C1(n4412), .C2(n4867), .A(n4391), .B(n4390), .ZN(U3139)
         );
  NAND2_X1 U5490 ( .A1(n4407), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4394)
         );
  OAI22_X1 U5491 ( .A1(n4816), .A2(n4408), .B1(n6949), .B2(n4445), .ZN(n4392)
         );
  AOI21_X1 U5492 ( .B1(n6944), .B2(n4909), .A(n4392), .ZN(n4393) );
  OAI211_X1 U5493 ( .C1(n4412), .C2(n4877), .A(n4394), .B(n4393), .ZN(U3134)
         );
  NAND2_X1 U5494 ( .A1(n4407), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4397)
         );
  OAI22_X1 U5495 ( .A1(n4802), .A2(n4408), .B1(n6943), .B2(n4445), .ZN(n4395)
         );
  AOI21_X1 U5496 ( .B1(n6938), .B2(n4909), .A(n4395), .ZN(n4396) );
  OAI211_X1 U5497 ( .C1(n4412), .C2(n4857), .A(n4397), .B(n4396), .ZN(U3133)
         );
  NAND2_X1 U5498 ( .A1(n4407), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4400)
         );
  OAI22_X1 U5499 ( .A1(n4832), .A2(n4408), .B1(n6908), .B2(n4445), .ZN(n4398)
         );
  AOI21_X1 U5500 ( .B1(n6905), .B2(n4909), .A(n4398), .ZN(n4399) );
  OAI211_X1 U5501 ( .C1(n4412), .C2(n4872), .A(n4400), .B(n4399), .ZN(U3136)
         );
  NAND2_X1 U5502 ( .A1(n4407), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4403)
         );
  OAI22_X1 U5503 ( .A1(n4820), .A2(n4408), .B1(n6967), .B2(n4445), .ZN(n4401)
         );
  AOI21_X1 U5504 ( .B1(n6962), .B2(n4909), .A(n4401), .ZN(n4402) );
  OAI211_X1 U5505 ( .C1(n4412), .C2(n4889), .A(n4403), .B(n4402), .ZN(U3137)
         );
  NAND2_X1 U5506 ( .A1(n4407), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4406)
         );
  OAI22_X1 U5507 ( .A1(n4905), .A2(n4408), .B1(n4932), .B2(n4445), .ZN(n4404)
         );
  AOI21_X1 U5508 ( .B1(n6841), .B2(n4909), .A(n4404), .ZN(n4405) );
  OAI211_X1 U5509 ( .C1(n4412), .C2(n4913), .A(n4406), .B(n4405), .ZN(U3138)
         );
  NAND2_X1 U5510 ( .A1(n4407), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4411)
         );
  OAI22_X1 U5511 ( .A1(n4828), .A2(n4408), .B1(n6904), .B2(n4445), .ZN(n4409)
         );
  AOI21_X1 U5512 ( .B1(n6901), .B2(n4909), .A(n4409), .ZN(n4410) );
  OAI211_X1 U5513 ( .C1(n4412), .C2(n4862), .A(n4411), .B(n4410), .ZN(U3135)
         );
  NAND2_X1 U5514 ( .A1(n4413), .A2(n3972), .ZN(n4419) );
  OAI21_X1 U5515 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n4414), .A(n4486), 
        .ZN(n6675) );
  INV_X1 U5516 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4416) );
  INV_X1 U5517 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4415) );
  OAI22_X1 U5518 ( .A1(n5369), .A2(n4416), .B1(n5366), .B2(n4415), .ZN(n4417)
         );
  AOI21_X1 U5519 ( .B1(n6675), .B2(n5506), .A(n4417), .ZN(n4418) );
  INV_X1 U5520 ( .A(n4502), .ZN(n4420) );
  XNOR2_X1 U5521 ( .A(n4420), .B(n4503), .ZN(n6672) );
  INV_X1 U5522 ( .A(n6672), .ZN(n4449) );
  OAI222_X1 U5523 ( .A1(n6345), .A2(n4449), .B1(n6064), .B2(n4416), .C1(n6636), 
        .C2(n5048), .ZN(U2884) );
  OAI222_X1 U5524 ( .A1(n6345), .A2(n6680), .B1(n6064), .B2(n4240), .C1(n6632), 
        .C2(n5048), .ZN(U2886) );
  NOR3_X1 U5525 ( .A1(n7010), .A2(n7016), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4422) );
  INV_X1 U5526 ( .A(n4422), .ZN(n4843) );
  NOR2_X1 U5527 ( .A1(n7000), .A2(n4843), .ZN(n4442) );
  AOI21_X1 U5528 ( .B1(n4799), .B2(n4842), .A(n4442), .ZN(n4424) );
  NAND2_X1 U5529 ( .A1(n4425), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4519) );
  NAND3_X1 U5530 ( .A1(n6923), .A2(n4424), .A3(n4519), .ZN(n4421) );
  OAI211_X1 U5531 ( .C1(n6923), .C2(n4422), .A(n6814), .B(n4421), .ZN(n4441)
         );
  NAND2_X1 U5532 ( .A1(n6923), .A2(n4519), .ZN(n4423) );
  OAI22_X1 U5533 ( .A1(n4424), .A2(n4423), .B1(n6930), .B2(n4843), .ZN(n4440)
         );
  AOI22_X1 U5534 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4441), .B1(n6958), 
        .B2(n4440), .ZN(n4427) );
  AOI22_X1 U5535 ( .A1(n6957), .A2(n4442), .B1(n6956), .B2(n4885), .ZN(n4426)
         );
  OAI211_X1 U5536 ( .C1(n6961), .C2(n4445), .A(n4427), .B(n4426), .ZN(U3128)
         );
  AOI22_X1 U5537 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4441), .B1(n6952), 
        .B2(n4440), .ZN(n4429) );
  AOI22_X1 U5538 ( .A1(n6951), .A2(n4442), .B1(n6950), .B2(n4885), .ZN(n4428)
         );
  OAI211_X1 U5539 ( .C1(n6955), .C2(n4445), .A(n4429), .B(n4428), .ZN(U3127)
         );
  AOI22_X1 U5540 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4441), .B1(n6934), 
        .B2(n4440), .ZN(n4431) );
  AOI22_X1 U5541 ( .A1(n6920), .A2(n4442), .B1(n6864), .B2(n4885), .ZN(n4430)
         );
  OAI211_X1 U5542 ( .C1(n6867), .C2(n4445), .A(n4431), .B(n4430), .ZN(U3124)
         );
  AOI22_X1 U5543 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4441), .B1(n6971), 
        .B2(n4440), .ZN(n4433) );
  AOI22_X1 U5544 ( .A1(n6970), .A2(n4442), .B1(n6968), .B2(n4885), .ZN(n4432)
         );
  OAI211_X1 U5545 ( .C1(n6975), .C2(n4445), .A(n4433), .B(n4432), .ZN(U3130)
         );
  AOI22_X1 U5546 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4441), .B1(n6946), 
        .B2(n4440), .ZN(n4435) );
  AOI22_X1 U5547 ( .A1(n6945), .A2(n4442), .B1(n6872), .B2(n4885), .ZN(n4434)
         );
  OAI211_X1 U5548 ( .C1(n6875), .C2(n4445), .A(n4435), .B(n4434), .ZN(U3126)
         );
  AOI22_X1 U5549 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4441), .B1(n6940), 
        .B2(n4440), .ZN(n4437) );
  AOI22_X1 U5550 ( .A1(n6939), .A2(n4442), .B1(n6868), .B2(n4885), .ZN(n4436)
         );
  OAI211_X1 U5551 ( .C1(n6871), .C2(n4445), .A(n4437), .B(n4436), .ZN(U3125)
         );
  AOI22_X1 U5552 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4441), .B1(n6981), 
        .B2(n4440), .ZN(n4439) );
  AOI22_X1 U5553 ( .A1(n6979), .A2(n4442), .B1(n6889), .B2(n4885), .ZN(n4438)
         );
  OAI211_X1 U5554 ( .C1(n6893), .C2(n4445), .A(n4439), .B(n4438), .ZN(U3131)
         );
  AOI22_X1 U5555 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4441), .B1(n6964), 
        .B2(n4440), .ZN(n4444) );
  AOI22_X1 U5556 ( .A1(n6963), .A2(n4442), .B1(n6880), .B2(n4885), .ZN(n4443)
         );
  OAI211_X1 U5557 ( .C1(n6883), .C2(n4445), .A(n4444), .B(n4443), .ZN(U3129)
         );
  AND2_X1 U5558 ( .A1(n4447), .A2(n4446), .ZN(n4448) );
  OR2_X1 U5559 ( .A1(n4448), .A2(n4509), .ZN(n6735) );
  INV_X1 U5560 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5760) );
  OAI222_X1 U5561 ( .A1(n6735), .A2(n6060), .B1(n6063), .B2(n5760), .C1(n6058), 
        .C2(n4449), .ZN(U2852) );
  NAND2_X1 U5562 ( .A1(n4450), .A2(n6985), .ZN(n4451) );
  AOI21_X1 U5563 ( .B1(n4451), .B2(STATEBS16_REG_SCAN_IN), .A(n6927), .ZN(
        n4455) );
  NOR2_X1 U5564 ( .A1(n6281), .A2(n4060), .ZN(n4522) );
  AND2_X1 U5565 ( .A1(n4522), .A2(n4173), .ZN(n6925) );
  AOI22_X1 U5566 ( .A1(n4455), .A2(n6925), .B1(n4452), .B2(n4594), .ZN(n4485)
         );
  NOR2_X1 U5567 ( .A1(n4849), .A2(n6863), .ZN(n5059) );
  INV_X1 U5568 ( .A(n6925), .ZN(n4454) );
  NAND3_X1 U5569 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7010), .ZN(n6931) );
  NOR2_X1 U5570 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6931), .ZN(n4457)
         );
  NOR2_X1 U5571 ( .A1(n3454), .A2(n4457), .ZN(n4453) );
  AOI21_X1 U5572 ( .B1(n4455), .B2(n4454), .A(n4453), .ZN(n4456) );
  OAI211_X1 U5573 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6930), .A(n5059), .B(n4456), .ZN(n4479) );
  NAND2_X1 U5574 ( .A1(n4479), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4460)
         );
  INV_X1 U5575 ( .A(n4457), .ZN(n4480) );
  OAI22_X1 U5576 ( .A1(n4816), .A2(n4480), .B1(n6985), .B2(n6875), .ZN(n4458)
         );
  AOI21_X1 U5577 ( .B1(n4482), .B2(n6872), .A(n4458), .ZN(n4459) );
  OAI211_X1 U5578 ( .C1(n4485), .C2(n4877), .A(n4460), .B(n4459), .ZN(U3102)
         );
  NAND2_X1 U5579 ( .A1(n4479), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4463)
         );
  OAI22_X1 U5580 ( .A1(n4824), .A2(n4480), .B1(n6985), .B2(n6893), .ZN(n4461)
         );
  AOI21_X1 U5581 ( .B1(n4482), .B2(n6889), .A(n4461), .ZN(n4462) );
  OAI211_X1 U5582 ( .C1(n4485), .C2(n4867), .A(n4463), .B(n4462), .ZN(U3107)
         );
  NAND2_X1 U5583 ( .A1(n4479), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4466)
         );
  OAI22_X1 U5584 ( .A1(n4820), .A2(n4480), .B1(n6985), .B2(n6883), .ZN(n4464)
         );
  AOI21_X1 U5585 ( .B1(n4482), .B2(n6880), .A(n4464), .ZN(n4465) );
  OAI211_X1 U5586 ( .C1(n4485), .C2(n4889), .A(n4466), .B(n4465), .ZN(U3105)
         );
  NAND2_X1 U5587 ( .A1(n4479), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4469)
         );
  OAI22_X1 U5588 ( .A1(n4828), .A2(n4480), .B1(n6985), .B2(n6955), .ZN(n4467)
         );
  AOI21_X1 U5589 ( .B1(n4482), .B2(n6950), .A(n4467), .ZN(n4468) );
  OAI211_X1 U5590 ( .C1(n4485), .C2(n4862), .A(n4469), .B(n4468), .ZN(U3103)
         );
  NAND2_X1 U5591 ( .A1(n4479), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4472)
         );
  OAI22_X1 U5592 ( .A1(n4905), .A2(n4480), .B1(n6985), .B2(n6975), .ZN(n4470)
         );
  AOI21_X1 U5593 ( .B1(n4482), .B2(n6968), .A(n4470), .ZN(n4471) );
  OAI211_X1 U5594 ( .C1(n4485), .C2(n4913), .A(n4472), .B(n4471), .ZN(U3106)
         );
  NAND2_X1 U5595 ( .A1(n4479), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4475)
         );
  OAI22_X1 U5596 ( .A1(n4802), .A2(n4480), .B1(n6985), .B2(n6871), .ZN(n4473)
         );
  AOI21_X1 U5597 ( .B1(n4482), .B2(n6868), .A(n4473), .ZN(n4474) );
  OAI211_X1 U5598 ( .C1(n4485), .C2(n4857), .A(n4475), .B(n4474), .ZN(U3101)
         );
  NAND2_X1 U5599 ( .A1(n4479), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4478)
         );
  OAI22_X1 U5600 ( .A1(n4832), .A2(n4480), .B1(n6985), .B2(n6961), .ZN(n4476)
         );
  AOI21_X1 U5601 ( .B1(n4482), .B2(n6956), .A(n4476), .ZN(n4477) );
  OAI211_X1 U5602 ( .C1(n4485), .C2(n4872), .A(n4478), .B(n4477), .ZN(U3104)
         );
  NAND2_X1 U5603 ( .A1(n4479), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4484)
         );
  OAI22_X1 U5604 ( .A1(n4812), .A2(n4480), .B1(n6985), .B2(n6867), .ZN(n4481)
         );
  AOI21_X1 U5605 ( .B1(n4482), .B2(n6864), .A(n4481), .ZN(n4483) );
  OAI211_X1 U5606 ( .C1(n4485), .C2(n4852), .A(n4484), .B(n4483), .ZN(U3100)
         );
  XNOR2_X1 U5607 ( .A(n4487), .B(n4486), .ZN(n5145) );
  AOI22_X1 U5608 ( .A1(n5307), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5460), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4491) );
  AOI22_X1 U5609 ( .A1(n5478), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4490) );
  AOI22_X1 U5610 ( .A1(n5338), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4489) );
  AOI22_X1 U5611 ( .A1(n5221), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4488) );
  NAND4_X1 U5612 ( .A1(n4491), .A2(n4490), .A3(n4489), .A4(n4488), .ZN(n4497)
         );
  AOI22_X1 U5613 ( .A1(n5332), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5614 ( .A1(n5333), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4494) );
  AOI22_X1 U5615 ( .A1(n5475), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4493) );
  AOI22_X1 U5616 ( .A1(n5486), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4492) );
  NAND4_X1 U5617 ( .A1(n4495), .A2(n4494), .A3(n4493), .A4(n4492), .ZN(n4496)
         );
  OAI21_X1 U5618 ( .B1(n4497), .B2(n4496), .A(n3972), .ZN(n4500) );
  NAND2_X1 U5619 ( .A1(n5501), .A2(EAX_REG_8__SCAN_IN), .ZN(n4499) );
  NAND2_X1 U5620 ( .A1(n5509), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4498)
         );
  NAND3_X1 U5621 ( .A1(n4500), .A2(n4499), .A3(n4498), .ZN(n4501) );
  AOI21_X1 U5622 ( .B1(n5145), .B2(n5506), .A(n4501), .ZN(n4507) );
  INV_X1 U5623 ( .A(n4576), .ZN(n4505) );
  AOI21_X1 U5624 ( .B1(n4507), .B2(n4506), .A(n4505), .ZN(n4586) );
  NOR2_X1 U5625 ( .A1(n4509), .A2(n4508), .ZN(n4510) );
  OR2_X1 U5626 ( .A1(n4589), .A2(n4510), .ZN(n6729) );
  OAI22_X1 U5627 ( .A1(n6729), .A2(n6060), .B1(n5146), .B2(n6063), .ZN(n4511)
         );
  AOI21_X1 U5628 ( .B1(n4586), .B2(n4592), .A(n4511), .ZN(n4512) );
  INV_X1 U5629 ( .A(n4512), .ZN(U2851) );
  OAI21_X1 U5630 ( .B1(n3188), .B2(n4515), .A(n4514), .ZN(n6756) );
  NAND2_X1 U5631 ( .A1(n6803), .A2(REIP_REG_6__SCAN_IN), .ZN(n6753) );
  OAI21_X1 U5632 ( .B1(n6162), .B2(n4319), .A(n6753), .ZN(n4517) );
  NOR2_X1 U5633 ( .A1(n6516), .A2(n6679), .ZN(n4516) );
  AOI211_X1 U5634 ( .C1(n6663), .C2(n6519), .A(n4517), .B(n4516), .ZN(n4518)
         );
  OAI21_X1 U5635 ( .B1(n6681), .B2(n6756), .A(n4518), .ZN(U2980) );
  INV_X1 U5636 ( .A(n4838), .ZN(n6924) );
  NAND2_X1 U5637 ( .A1(n4519), .A2(n6924), .ZN(n6289) );
  INV_X1 U5638 ( .A(n6284), .ZN(n4520) );
  NOR3_X1 U5639 ( .A1(n6289), .A2(n4520), .A3(n6288), .ZN(n4521) );
  NOR2_X1 U5640 ( .A1(n4521), .A2(n6927), .ZN(n4530) );
  NAND2_X1 U5641 ( .A1(n4522), .A2(n6546), .ZN(n5063) );
  OR2_X1 U5642 ( .A1(n5063), .A2(n4523), .ZN(n4525) );
  INV_X1 U5643 ( .A(n6918), .ZN(n4524) );
  NAND2_X1 U5644 ( .A1(n4524), .A2(n7016), .ZN(n4555) );
  NAND2_X1 U5645 ( .A1(n4525), .A2(n4555), .ZN(n4532) );
  NAND3_X1 U5646 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7016), .A3(n7010), .ZN(n5057) );
  INV_X1 U5647 ( .A(n5057), .ZN(n4526) );
  AOI22_X1 U5648 ( .A1(n4530), .A2(n4532), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4526), .ZN(n4560) );
  AND2_X1 U5649 ( .A1(n4527), .A2(n6284), .ZN(n4528) );
  OAI22_X1 U5650 ( .A1(n4812), .A2(n4555), .B1(n6867), .B2(n4554), .ZN(n4529)
         );
  AOI21_X1 U5651 ( .B1(n6864), .B2(n5085), .A(n4529), .ZN(n4535) );
  INV_X1 U5652 ( .A(n4530), .ZN(n4533) );
  INV_X1 U5653 ( .A(n6814), .ZN(n6926) );
  AOI21_X1 U5654 ( .B1(n6927), .B2(n5057), .A(n6926), .ZN(n4531) );
  OAI21_X1 U5655 ( .B1(n4533), .B2(n4532), .A(n4531), .ZN(n4557) );
  NAND2_X1 U5656 ( .A1(n4557), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4534) );
  OAI211_X1 U5657 ( .C1(n4560), .C2(n4852), .A(n4535), .B(n4534), .ZN(U3044)
         );
  OAI22_X1 U5658 ( .A1(n4824), .A2(n4555), .B1(n6893), .B2(n4554), .ZN(n4536)
         );
  AOI21_X1 U5659 ( .B1(n6889), .B2(n5085), .A(n4536), .ZN(n4538) );
  NAND2_X1 U5660 ( .A1(n4557), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4537) );
  OAI211_X1 U5661 ( .C1(n4560), .C2(n4867), .A(n4538), .B(n4537), .ZN(U3051)
         );
  OAI22_X1 U5662 ( .A1(n4828), .A2(n4555), .B1(n6955), .B2(n4554), .ZN(n4539)
         );
  AOI21_X1 U5663 ( .B1(n6950), .B2(n5085), .A(n4539), .ZN(n4541) );
  NAND2_X1 U5664 ( .A1(n4557), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4540) );
  OAI211_X1 U5665 ( .C1(n4560), .C2(n4862), .A(n4541), .B(n4540), .ZN(U3047)
         );
  OAI22_X1 U5666 ( .A1(n4820), .A2(n4555), .B1(n6883), .B2(n4554), .ZN(n4542)
         );
  AOI21_X1 U5667 ( .B1(n6880), .B2(n5085), .A(n4542), .ZN(n4544) );
  NAND2_X1 U5668 ( .A1(n4557), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4543) );
  OAI211_X1 U5669 ( .C1(n4560), .C2(n4889), .A(n4544), .B(n4543), .ZN(U3049)
         );
  OAI22_X1 U5670 ( .A1(n4905), .A2(n4555), .B1(n6975), .B2(n4554), .ZN(n4545)
         );
  AOI21_X1 U5671 ( .B1(n6968), .B2(n5085), .A(n4545), .ZN(n4547) );
  NAND2_X1 U5672 ( .A1(n4557), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4546) );
  OAI211_X1 U5673 ( .C1(n4560), .C2(n4913), .A(n4547), .B(n4546), .ZN(U3050)
         );
  OAI22_X1 U5674 ( .A1(n4802), .A2(n4555), .B1(n6871), .B2(n4554), .ZN(n4548)
         );
  AOI21_X1 U5675 ( .B1(n6868), .B2(n5085), .A(n4548), .ZN(n4550) );
  NAND2_X1 U5676 ( .A1(n4557), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4549) );
  OAI211_X1 U5677 ( .C1(n4560), .C2(n4857), .A(n4550), .B(n4549), .ZN(U3045)
         );
  OAI22_X1 U5678 ( .A1(n4816), .A2(n4555), .B1(n6875), .B2(n4554), .ZN(n4551)
         );
  AOI21_X1 U5679 ( .B1(n6872), .B2(n5085), .A(n4551), .ZN(n4553) );
  NAND2_X1 U5680 ( .A1(n4557), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4552) );
  OAI211_X1 U5681 ( .C1(n4560), .C2(n4877), .A(n4553), .B(n4552), .ZN(U3046)
         );
  OAI22_X1 U5682 ( .A1(n4832), .A2(n4555), .B1(n6961), .B2(n4554), .ZN(n4556)
         );
  AOI21_X1 U5683 ( .B1(n6956), .B2(n5085), .A(n4556), .ZN(n4559) );
  NAND2_X1 U5684 ( .A1(n4557), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4558) );
  OAI211_X1 U5685 ( .C1(n4560), .C2(n4872), .A(n4559), .B(n4558), .ZN(U3048)
         );
  INV_X1 U5686 ( .A(n4586), .ZN(n5155) );
  INV_X1 U5687 ( .A(DATAI_8_), .ZN(n6638) );
  INV_X1 U5688 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6582) );
  OAI222_X1 U5689 ( .A1(n5155), .A2(n6345), .B1(n5048), .B2(n6638), .C1(n6064), 
        .C2(n6582), .ZN(U2883) );
  INV_X1 U5690 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4561) );
  XNOR2_X1 U5691 ( .A(n4562), .B(n4561), .ZN(n6491) );
  OR2_X1 U5692 ( .A1(n6491), .A2(n5499), .ZN(n4575) );
  AOI22_X1 U5693 ( .A1(n5510), .A2(EAX_REG_9__SCAN_IN), .B1(n5509), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5694 ( .A1(n5486), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4566) );
  AOI22_X1 U5695 ( .A1(n5460), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U5696 ( .A1(n5338), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4564) );
  AOI22_X1 U5697 ( .A1(n5480), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4563) );
  NAND4_X1 U5698 ( .A1(n4566), .A2(n4565), .A3(n4564), .A4(n4563), .ZN(n4572)
         );
  AOI22_X1 U5699 ( .A1(n5332), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U5700 ( .A1(n5478), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U5701 ( .A1(n5333), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5702 ( .A1(n5307), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4567) );
  NAND4_X1 U5703 ( .A1(n4570), .A2(n4569), .A3(n4568), .A4(n4567), .ZN(n4571)
         );
  OAI21_X1 U5704 ( .B1(n4572), .B2(n4571), .A(n3972), .ZN(n4573) );
  AOI21_X1 U5705 ( .B1(n4577), .B2(n4576), .A(n4898), .ZN(n6488) );
  INV_X1 U5706 ( .A(n6488), .ZN(n4579) );
  AOI22_X1 U5707 ( .A1(n5004), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6561), .ZN(n4578) );
  OAI21_X1 U5708 ( .B1(n4579), .B2(n6345), .A(n4578), .ZN(U2882) );
  OR2_X1 U5709 ( .A1(n4581), .A2(n4580), .ZN(n4582) );
  NAND2_X1 U5710 ( .A1(n4583), .A2(n4582), .ZN(n6728) );
  AOI22_X1 U5711 ( .A1(n6694), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6785), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4584) );
  OAI21_X1 U5712 ( .B1(n6704), .B2(n5145), .A(n4584), .ZN(n4585) );
  AOI21_X1 U5713 ( .B1(n4586), .B2(n6698), .A(n4585), .ZN(n4587) );
  OAI21_X1 U5714 ( .B1(n6728), .B2(n6681), .A(n4587), .ZN(U2978) );
  OR2_X1 U5715 ( .A1(n4589), .A2(n4588), .ZN(n4590) );
  NAND2_X1 U5716 ( .A1(n4895), .A2(n4590), .ZN(n6717) );
  OAI22_X1 U5717 ( .A1(n6717), .A2(n6060), .B1(n6494), .B2(n6063), .ZN(n4591)
         );
  AOI21_X1 U5718 ( .B1(n6488), .B2(n4592), .A(n4591), .ZN(n4593) );
  INV_X1 U5719 ( .A(n4593), .ZN(U2850) );
  AND2_X1 U5720 ( .A1(n3293), .A2(n4173), .ZN(n4602) );
  INV_X1 U5721 ( .A(n4602), .ZN(n4597) );
  INV_X1 U5722 ( .A(n4594), .ZN(n6860) );
  NAND2_X1 U5723 ( .A1(n4596), .A2(n4595), .ZN(n4847) );
  OAI22_X1 U5724 ( .A1(n4597), .A2(n6927), .B1(n6860), .B2(n4847), .ZN(n4628)
         );
  NOR2_X1 U5725 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4598), .ZN(n4601)
         );
  INV_X1 U5726 ( .A(n4601), .ZN(n4626) );
  OAI22_X1 U5727 ( .A1(n4824), .A2(n4626), .B1(n6986), .B2(n6894), .ZN(n4599)
         );
  AOI21_X1 U5728 ( .B1(n6981), .B2(n4628), .A(n4599), .ZN(n4607) );
  INV_X1 U5729 ( .A(n4849), .ZN(n6852) );
  AOI21_X1 U5730 ( .B1(n4847), .B2(STATE2_REG_2__SCAN_IN), .A(n4600), .ZN(
        n4844) );
  OAI211_X1 U5731 ( .C1(n3454), .C2(n4601), .A(n6852), .B(n4844), .ZN(n4605)
         );
  NAND3_X1 U5732 ( .A1(n4632), .A2(n6923), .A3(n6894), .ZN(n4603) );
  INV_X1 U5733 ( .A(n4806), .ZN(n6858) );
  AOI21_X1 U5734 ( .B1(n4603), .B2(n6858), .A(n4602), .ZN(n4604) );
  NAND2_X1 U5735 ( .A1(n4629), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4606) );
  OAI211_X1 U5736 ( .C1(n4632), .C2(n6893), .A(n4607), .B(n4606), .ZN(U3091)
         );
  OAI22_X1 U5737 ( .A1(n4812), .A2(n4626), .B1(n6937), .B2(n6894), .ZN(n4608)
         );
  AOI21_X1 U5738 ( .B1(n6934), .B2(n4628), .A(n4608), .ZN(n4610) );
  NAND2_X1 U5739 ( .A1(n4629), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4609) );
  OAI211_X1 U5740 ( .C1(n4632), .C2(n6867), .A(n4610), .B(n4609), .ZN(U3084)
         );
  OAI22_X1 U5741 ( .A1(n4802), .A2(n4626), .B1(n6943), .B2(n6894), .ZN(n4611)
         );
  AOI21_X1 U5742 ( .B1(n6940), .B2(n4628), .A(n4611), .ZN(n4613) );
  NAND2_X1 U5743 ( .A1(n4629), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4612) );
  OAI211_X1 U5744 ( .C1(n4632), .C2(n6871), .A(n4613), .B(n4612), .ZN(U3085)
         );
  OAI22_X1 U5745 ( .A1(n4905), .A2(n4626), .B1(n4932), .B2(n6894), .ZN(n4614)
         );
  AOI21_X1 U5746 ( .B1(n6971), .B2(n4628), .A(n4614), .ZN(n4616) );
  NAND2_X1 U5747 ( .A1(n4629), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4615) );
  OAI211_X1 U5748 ( .C1(n4632), .C2(n6975), .A(n4616), .B(n4615), .ZN(U3090)
         );
  OAI22_X1 U5749 ( .A1(n4816), .A2(n4626), .B1(n6949), .B2(n6894), .ZN(n4617)
         );
  AOI21_X1 U5750 ( .B1(n6946), .B2(n4628), .A(n4617), .ZN(n4619) );
  NAND2_X1 U5751 ( .A1(n4629), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4618) );
  OAI211_X1 U5752 ( .C1(n4632), .C2(n6875), .A(n4619), .B(n4618), .ZN(U3086)
         );
  OAI22_X1 U5753 ( .A1(n4828), .A2(n4626), .B1(n6904), .B2(n6894), .ZN(n4620)
         );
  AOI21_X1 U5754 ( .B1(n6952), .B2(n4628), .A(n4620), .ZN(n4622) );
  NAND2_X1 U5755 ( .A1(n4629), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4621) );
  OAI211_X1 U5756 ( .C1(n4632), .C2(n6955), .A(n4622), .B(n4621), .ZN(U3087)
         );
  OAI22_X1 U5757 ( .A1(n4820), .A2(n4626), .B1(n6967), .B2(n6894), .ZN(n4623)
         );
  AOI21_X1 U5758 ( .B1(n6964), .B2(n4628), .A(n4623), .ZN(n4625) );
  NAND2_X1 U5759 ( .A1(n4629), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4624) );
  OAI211_X1 U5760 ( .C1(n4632), .C2(n6883), .A(n4625), .B(n4624), .ZN(U3089)
         );
  OAI22_X1 U5761 ( .A1(n4832), .A2(n4626), .B1(n6908), .B2(n6894), .ZN(n4627)
         );
  AOI21_X1 U5762 ( .B1(n6958), .B2(n4628), .A(n4627), .ZN(n4631) );
  NAND2_X1 U5763 ( .A1(n4629), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4630) );
  OAI211_X1 U5764 ( .C1(n4632), .C2(n6961), .A(n4631), .B(n4630), .ZN(U3088)
         );
  INV_X1 U5765 ( .A(n6545), .ZN(n5036) );
  INV_X1 U5766 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6537) );
  AND2_X1 U5767 ( .A1(n6537), .A2(REIP_REG_1__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U5768 ( .A1(n6532), .A2(n4633), .B1(n6543), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4638) );
  OR2_X1 U5769 ( .A1(n6507), .A2(REIP_REG_1__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U5770 ( .A1(n5033), .A2(n6504), .ZN(n6538) );
  NAND2_X1 U5771 ( .A1(n6538), .A2(REIP_REG_2__SCAN_IN), .ZN(n4637) );
  INV_X1 U5772 ( .A(n6703), .ZN(n4634) );
  AOI22_X1 U5773 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6525), .B1(n6518), 
        .B2(n4634), .ZN(n4636) );
  NAND2_X1 U5774 ( .A1(n6798), .A2(n6539), .ZN(n4635) );
  NAND4_X1 U5775 ( .A1(n4638), .A2(n4637), .A3(n4636), .A4(n4635), .ZN(n4639)
         );
  AOI21_X1 U5776 ( .B1(n5036), .B2(n4060), .A(n4639), .ZN(n4640) );
  OAI21_X1 U5777 ( .B1(n4641), .B2(n6528), .A(n4640), .ZN(U2825) );
  XOR2_X1 U5778 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4642), .Z(n6444) );
  AOI22_X1 U5779 ( .A1(n5333), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4646) );
  AOI22_X1 U5780 ( .A1(n5307), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4645) );
  AOI22_X1 U5781 ( .A1(n5486), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4644) );
  AOI22_X1 U5782 ( .A1(n5478), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4643) );
  NAND4_X1 U5783 ( .A1(n4646), .A2(n4645), .A3(n4644), .A4(n4643), .ZN(n4652)
         );
  AOI22_X1 U5784 ( .A1(n5332), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4650) );
  AOI22_X1 U5785 ( .A1(n5475), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5460), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4649) );
  AOI22_X1 U5786 ( .A1(n5221), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4648) );
  AOI22_X1 U5787 ( .A1(n5338), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4647) );
  NAND4_X1 U5788 ( .A1(n4650), .A2(n4649), .A3(n4648), .A4(n4647), .ZN(n4651)
         );
  OR2_X1 U5789 ( .A1(n4652), .A2(n4651), .ZN(n4653) );
  AOI22_X1 U5790 ( .A1(n3972), .A2(n4653), .B1(n5509), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4655) );
  NAND2_X1 U5791 ( .A1(n5501), .A2(EAX_REG_14__SCAN_IN), .ZN(n4654) );
  OAI211_X1 U5792 ( .C1(n6444), .C2(n5499), .A(n4655), .B(n4654), .ZN(n4901)
         );
  XNOR2_X1 U5793 ( .A(n4656), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6457)
         );
  AOI22_X1 U5794 ( .A1(n5332), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4660) );
  AOI22_X1 U5795 ( .A1(n5307), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5796 ( .A1(n5221), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5797 ( .A1(n5338), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4657) );
  NAND4_X1 U5798 ( .A1(n4660), .A2(n4659), .A3(n4658), .A4(n4657), .ZN(n4666)
         );
  AOI22_X1 U5799 ( .A1(n5333), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4664) );
  AOI22_X1 U5800 ( .A1(n5460), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4663) );
  AOI22_X1 U5801 ( .A1(n5486), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4662) );
  AOI22_X1 U5802 ( .A1(n5476), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4661) );
  NAND4_X1 U5803 ( .A1(n4664), .A2(n4663), .A3(n4662), .A4(n4661), .ZN(n4665)
         );
  OAI21_X1 U5804 ( .B1(n4666), .B2(n4665), .A(n3972), .ZN(n4669) );
  NAND2_X1 U5805 ( .A1(n5501), .A2(EAX_REG_13__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U5806 ( .A1(n5509), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4667)
         );
  NAND3_X1 U5807 ( .A1(n4669), .A2(n4668), .A3(n4667), .ZN(n4670) );
  AOI21_X1 U5808 ( .B1(n6457), .B2(n5506), .A(n4670), .ZN(n5044) );
  XOR2_X1 U5809 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n4671), .Z(n6662) );
  INV_X1 U5810 ( .A(n6662), .ZN(n4686) );
  AOI22_X1 U5811 ( .A1(n5307), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5333), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4675) );
  AOI22_X1 U5812 ( .A1(n5486), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5813 ( .A1(n5332), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5814 ( .A1(n5480), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4672) );
  NAND4_X1 U5815 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(n4672), .ZN(n4681)
         );
  AOI22_X1 U5816 ( .A1(n5485), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4679) );
  AOI22_X1 U5817 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5475), .B1(n5476), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5818 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5460), .B1(n5221), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4677) );
  AOI22_X1 U5819 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n5338), .B1(n5487), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4676) );
  NAND4_X1 U5820 ( .A1(n4679), .A2(n4678), .A3(n4677), .A4(n4676), .ZN(n4680)
         );
  OAI21_X1 U5821 ( .B1(n4681), .B2(n4680), .A(n3972), .ZN(n4684) );
  NAND2_X1 U5822 ( .A1(n5501), .A2(EAX_REG_12__SCAN_IN), .ZN(n4683) );
  NAND2_X1 U5823 ( .A1(n5509), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4682)
         );
  NAND3_X1 U5824 ( .A1(n4684), .A2(n4683), .A3(n4682), .ZN(n4685) );
  AOI21_X1 U5825 ( .B1(n4686), .B2(n5506), .A(n4685), .ZN(n5002) );
  XNOR2_X1 U5826 ( .A(n4687), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5101)
         );
  AOI22_X1 U5827 ( .A1(n5333), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4691) );
  AOI22_X1 U5828 ( .A1(n5460), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4690) );
  AOI22_X1 U5829 ( .A1(n5478), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4689) );
  AOI22_X1 U5830 ( .A1(n5486), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4688) );
  NAND4_X1 U5831 ( .A1(n4691), .A2(n4690), .A3(n4689), .A4(n4688), .ZN(n4697)
         );
  AOI22_X1 U5832 ( .A1(n5332), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4695) );
  AOI22_X1 U5833 ( .A1(n5307), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4694) );
  AOI22_X1 U5834 ( .A1(n5480), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4693) );
  AOI22_X1 U5835 ( .A1(n5221), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5338), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4692) );
  NAND4_X1 U5836 ( .A1(n4695), .A2(n4694), .A3(n4693), .A4(n4692), .ZN(n4696)
         );
  OAI21_X1 U5837 ( .B1(n4697), .B2(n4696), .A(n3972), .ZN(n4700) );
  NAND2_X1 U5838 ( .A1(n5501), .A2(EAX_REG_11__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U5839 ( .A1(n5509), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4698)
         );
  NAND3_X1 U5840 ( .A1(n4700), .A2(n4699), .A3(n4698), .ZN(n4701) );
  AOI21_X1 U5841 ( .B1(n5101), .B2(n5506), .A(n4701), .ZN(n4955) );
  OR2_X1 U5842 ( .A1(n5002), .A2(n4955), .ZN(n4998) );
  NOR2_X1 U5843 ( .A1(n5044), .A2(n4998), .ZN(n4899) );
  AND2_X1 U5844 ( .A1(n4901), .A2(n4899), .ZN(n4716) );
  XOR2_X1 U5845 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n4702), .Z(n6477) );
  AOI22_X1 U5846 ( .A1(n5485), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4706) );
  AOI22_X1 U5847 ( .A1(n5486), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5848 ( .A1(n5460), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5849 ( .A1(n5221), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5338), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4703) );
  NAND4_X1 U5850 ( .A1(n4706), .A2(n4705), .A3(n4704), .A4(n4703), .ZN(n4712)
         );
  AOI22_X1 U5851 ( .A1(n5478), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4710) );
  AOI22_X1 U5852 ( .A1(n5307), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5333), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4709) );
  AOI22_X1 U5853 ( .A1(n5332), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4708) );
  AOI22_X1 U5854 ( .A1(n3525), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4707) );
  NAND4_X1 U5855 ( .A1(n4710), .A2(n4709), .A3(n4708), .A4(n4707), .ZN(n4711)
         );
  OR2_X1 U5856 ( .A1(n4712), .A2(n4711), .ZN(n4713) );
  AOI22_X1 U5857 ( .A1(n3972), .A2(n4713), .B1(n5509), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U5858 ( .A1(n5501), .A2(EAX_REG_10__SCAN_IN), .ZN(n4714) );
  OAI211_X1 U5859 ( .C1(n6477), .C2(n5499), .A(n4715), .B(n4714), .ZN(n4897)
         );
  NAND2_X1 U5860 ( .A1(n4898), .A2(n4735), .ZN(n4903) );
  INV_X1 U5861 ( .A(n4903), .ZN(n4738) );
  NAND2_X1 U5862 ( .A1(n4717), .A2(n5820), .ZN(n4719) );
  INV_X1 U5863 ( .A(n4981), .ZN(n4718) );
  NAND2_X1 U5864 ( .A1(n4719), .A2(n4718), .ZN(n6173) );
  AOI22_X1 U5865 ( .A1(n5485), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4723) );
  AOI22_X1 U5866 ( .A1(n5476), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5460), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4722) );
  AOI22_X1 U5867 ( .A1(n3525), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4721) );
  AOI22_X1 U5868 ( .A1(n5480), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4720) );
  NAND4_X1 U5869 ( .A1(n4723), .A2(n4722), .A3(n4721), .A4(n4720), .ZN(n4729)
         );
  AOI22_X1 U5870 ( .A1(n5307), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5486), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4727) );
  AOI22_X1 U5871 ( .A1(n5333), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4726) );
  AOI22_X1 U5872 ( .A1(n5332), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4725) );
  AOI22_X1 U5873 ( .A1(n5338), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4724) );
  NAND4_X1 U5874 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4728)
         );
  OAI21_X1 U5875 ( .B1(n4729), .B2(n4728), .A(n3972), .ZN(n4732) );
  NAND2_X1 U5876 ( .A1(n5501), .A2(EAX_REG_15__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U5877 ( .A1(n5509), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4730)
         );
  NAND3_X1 U5878 ( .A1(n4732), .A2(n4731), .A3(n4730), .ZN(n4733) );
  AOI21_X1 U5879 ( .B1(n6173), .B2(n5506), .A(n4733), .ZN(n4734) );
  INV_X1 U5880 ( .A(n4734), .ZN(n4737) );
  OAI21_X1 U5881 ( .B1(n4738), .B2(n4737), .A(n4986), .ZN(n6177) );
  AOI22_X1 U5882 ( .A1(n5004), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6561), .ZN(n4739) );
  OAI21_X1 U5883 ( .B1(n6177), .B2(n6345), .A(n4739), .ZN(U2876) );
  INV_X1 U5884 ( .A(EBX_REG_15__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U5885 ( .A1(n3211), .A2(n4740), .ZN(n4741) );
  NAND2_X1 U5886 ( .A1(n3201), .A2(n4741), .ZN(n4945) );
  OAI222_X1 U5887 ( .A1(n6177), .A2(n6058), .B1(n6063), .B2(n4742), .C1(n6060), 
        .C2(n4945), .ZN(U2844) );
  OAI21_X1 U5888 ( .B1(n4745), .B2(n4744), .A(n4743), .ZN(n6719) );
  INV_X1 U5889 ( .A(n6491), .ZN(n4747) );
  NAND2_X1 U5890 ( .A1(n6803), .A2(REIP_REG_9__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U5891 ( .A1(n6694), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4746)
         );
  OAI211_X1 U5892 ( .C1(n6704), .C2(n4747), .A(n6716), .B(n4746), .ZN(n4748)
         );
  AOI21_X1 U5893 ( .B1(n6488), .B2(n6698), .A(n4748), .ZN(n4749) );
  OAI21_X1 U5894 ( .B1(n6719), .B2(n6681), .A(n4749), .ZN(U2977) );
  INV_X1 U5895 ( .A(n4804), .ZN(n4750) );
  NOR3_X2 U5896 ( .A1(n4750), .A2(n4751), .A3(n6817), .ZN(n4801) );
  AND2_X1 U5897 ( .A1(n4751), .A2(n6284), .ZN(n4752) );
  NAND2_X1 U5898 ( .A1(n6294), .A2(n4752), .ZN(n4923) );
  INV_X1 U5899 ( .A(n4923), .ZN(n4753) );
  INV_X1 U5900 ( .A(n4944), .ZN(n4754) );
  NOR3_X1 U5901 ( .A1(n4801), .A2(n4754), .A3(n6927), .ZN(n4755) );
  NAND2_X1 U5902 ( .A1(n6546), .A2(n3293), .ZN(n4915) );
  OAI21_X1 U5903 ( .B1(n4755), .B2(n4806), .A(n4915), .ZN(n4759) );
  NAND3_X1 U5904 ( .A1(n7016), .A2(n7010), .A3(n7005), .ZN(n4920) );
  NOR2_X1 U5905 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4920), .ZN(n4789)
         );
  INV_X1 U5906 ( .A(n4789), .ZN(n4757) );
  AOI211_X1 U5907 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4757), .A(n4849), .B(
        n4756), .ZN(n4758) );
  INV_X1 U5908 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4765) );
  INV_X1 U5909 ( .A(n4760), .ZN(n4761) );
  OAI22_X1 U5910 ( .A1(n4915), .A2(n6927), .B1(n6860), .B2(n4761), .ZN(n4792)
         );
  AOI22_X1 U5911 ( .A1(n6939), .A2(n4789), .B1(n4801), .B2(n6868), .ZN(n4762)
         );
  OAI21_X1 U5912 ( .B1(n6871), .B2(n4944), .A(n4762), .ZN(n4763) );
  AOI21_X1 U5913 ( .B1(n6940), .B2(n4792), .A(n4763), .ZN(n4764) );
  OAI21_X1 U5914 ( .B1(n4795), .B2(n4765), .A(n4764), .ZN(U3021) );
  AOI22_X1 U5915 ( .A1(n6979), .A2(n4789), .B1(n4801), .B2(n6889), .ZN(n4766)
         );
  OAI21_X1 U5916 ( .B1(n6893), .B2(n4944), .A(n4766), .ZN(n4767) );
  AOI21_X1 U5917 ( .B1(n6981), .B2(n4792), .A(n4767), .ZN(n4768) );
  OAI21_X1 U5918 ( .B1(n4795), .B2(n4769), .A(n4768), .ZN(U3027) );
  AOI22_X1 U5919 ( .A1(n6957), .A2(n4789), .B1(n4801), .B2(n6956), .ZN(n4770)
         );
  OAI21_X1 U5920 ( .B1(n6961), .B2(n4944), .A(n4770), .ZN(n4771) );
  AOI21_X1 U5921 ( .B1(n6958), .B2(n4792), .A(n4771), .ZN(n4772) );
  OAI21_X1 U5922 ( .B1(n4795), .B2(n5893), .A(n4772), .ZN(U3024) );
  INV_X1 U5923 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4776) );
  AOI22_X1 U5924 ( .A1(n6951), .A2(n4789), .B1(n4801), .B2(n6950), .ZN(n4773)
         );
  OAI21_X1 U5925 ( .B1(n6955), .B2(n4944), .A(n4773), .ZN(n4774) );
  AOI21_X1 U5926 ( .B1(n6952), .B2(n4792), .A(n4774), .ZN(n4775) );
  OAI21_X1 U5927 ( .B1(n4795), .B2(n4776), .A(n4775), .ZN(U3023) );
  AOI22_X1 U5928 ( .A1(n6945), .A2(n4789), .B1(n4801), .B2(n6872), .ZN(n4777)
         );
  OAI21_X1 U5929 ( .B1(n6875), .B2(n4944), .A(n4777), .ZN(n4778) );
  AOI21_X1 U5930 ( .B1(n6946), .B2(n4792), .A(n4778), .ZN(n4779) );
  OAI21_X1 U5931 ( .B1(n4795), .B2(n4780), .A(n4779), .ZN(U3022) );
  AOI22_X1 U5932 ( .A1(n6920), .A2(n4789), .B1(n4801), .B2(n6864), .ZN(n4781)
         );
  OAI21_X1 U5933 ( .B1(n6867), .B2(n4944), .A(n4781), .ZN(n4782) );
  AOI21_X1 U5934 ( .B1(n6934), .B2(n4792), .A(n4782), .ZN(n4783) );
  OAI21_X1 U5935 ( .B1(n4795), .B2(n4784), .A(n4783), .ZN(U3020) );
  AOI22_X1 U5936 ( .A1(n6963), .A2(n4789), .B1(n4801), .B2(n6880), .ZN(n4785)
         );
  OAI21_X1 U5937 ( .B1(n6883), .B2(n4944), .A(n4785), .ZN(n4786) );
  AOI21_X1 U5938 ( .B1(n6964), .B2(n4792), .A(n4786), .ZN(n4787) );
  OAI21_X1 U5939 ( .B1(n4795), .B2(n4788), .A(n4787), .ZN(U3025) );
  AOI22_X1 U5940 ( .A1(n6970), .A2(n4789), .B1(n4801), .B2(n6968), .ZN(n4790)
         );
  OAI21_X1 U5941 ( .B1(n6975), .B2(n4944), .A(n4790), .ZN(n4791) );
  AOI21_X1 U5942 ( .B1(n6971), .B2(n4792), .A(n4791), .ZN(n4793) );
  OAI21_X1 U5943 ( .B1(n4795), .B2(n4794), .A(n4793), .ZN(U3026) );
  NAND2_X1 U5944 ( .A1(n4898), .A2(n4897), .ZN(n4999) );
  OAI21_X1 U5945 ( .B1(n4898), .B2(n4897), .A(n4999), .ZN(n6476) );
  INV_X1 U5946 ( .A(DATAI_10_), .ZN(n6643) );
  INV_X1 U5947 ( .A(EAX_REG_10__SCAN_IN), .ZN(n4796) );
  OAI222_X1 U5948 ( .A1(n6476), .A2(n6345), .B1(n5048), .B2(n6643), .C1(n6064), 
        .C2(n4796), .ZN(U2881) );
  INV_X1 U5949 ( .A(n4906), .ZN(n4797) );
  AOI21_X1 U5950 ( .B1(n4799), .B2(n4798), .A(n4797), .ZN(n4805) );
  INV_X1 U5951 ( .A(n4805), .ZN(n4800) );
  AOI22_X1 U5952 ( .A1(n4800), .A2(n6923), .B1(n4809), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n4914) );
  INV_X1 U5953 ( .A(n4801), .ZN(n4907) );
  OAI22_X1 U5954 ( .A1(n4907), .A2(n6871), .B1(n4906), .B2(n4802), .ZN(n4803)
         );
  AOI21_X1 U5955 ( .B1(n6868), .B2(n4909), .A(n4803), .ZN(n4811) );
  AOI21_X1 U5956 ( .B1(n4804), .B2(n3196), .A(n6679), .ZN(n4807) );
  OAI21_X1 U5957 ( .B1(n4807), .B2(n4806), .A(n4805), .ZN(n4808) );
  OAI211_X1 U5958 ( .C1(n4809), .C2(n6923), .A(n6814), .B(n4808), .ZN(n4910)
         );
  NAND2_X1 U5959 ( .A1(n4910), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4810)
         );
  OAI211_X1 U5960 ( .C1(n4914), .C2(n4857), .A(n4811), .B(n4810), .ZN(U3141)
         );
  OAI22_X1 U5961 ( .A1(n4907), .A2(n6867), .B1(n4906), .B2(n4812), .ZN(n4813)
         );
  AOI21_X1 U5962 ( .B1(n6864), .B2(n4909), .A(n4813), .ZN(n4815) );
  NAND2_X1 U5963 ( .A1(n4910), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4814)
         );
  OAI211_X1 U5964 ( .C1(n4914), .C2(n4852), .A(n4815), .B(n4814), .ZN(U3140)
         );
  OAI22_X1 U5965 ( .A1(n4907), .A2(n6875), .B1(n4906), .B2(n4816), .ZN(n4817)
         );
  AOI21_X1 U5966 ( .B1(n6872), .B2(n4909), .A(n4817), .ZN(n4819) );
  NAND2_X1 U5967 ( .A1(n4910), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4818)
         );
  OAI211_X1 U5968 ( .C1(n4914), .C2(n4877), .A(n4819), .B(n4818), .ZN(U3142)
         );
  OAI22_X1 U5969 ( .A1(n4907), .A2(n6883), .B1(n4906), .B2(n4820), .ZN(n4821)
         );
  AOI21_X1 U5970 ( .B1(n6880), .B2(n4909), .A(n4821), .ZN(n4823) );
  NAND2_X1 U5971 ( .A1(n4910), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4822)
         );
  OAI211_X1 U5972 ( .C1(n4914), .C2(n4889), .A(n4823), .B(n4822), .ZN(U3145)
         );
  OAI22_X1 U5973 ( .A1(n4907), .A2(n6893), .B1(n4906), .B2(n4824), .ZN(n4825)
         );
  AOI21_X1 U5974 ( .B1(n6889), .B2(n4909), .A(n4825), .ZN(n4827) );
  NAND2_X1 U5975 ( .A1(n4910), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4826)
         );
  OAI211_X1 U5976 ( .C1(n4914), .C2(n4867), .A(n4827), .B(n4826), .ZN(U3147)
         );
  OAI22_X1 U5977 ( .A1(n4907), .A2(n6955), .B1(n4906), .B2(n4828), .ZN(n4829)
         );
  AOI21_X1 U5978 ( .B1(n6950), .B2(n4909), .A(n4829), .ZN(n4831) );
  NAND2_X1 U5979 ( .A1(n4910), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4830)
         );
  OAI211_X1 U5980 ( .C1(n4914), .C2(n4862), .A(n4831), .B(n4830), .ZN(U3143)
         );
  OAI22_X1 U5981 ( .A1(n4907), .A2(n6961), .B1(n4906), .B2(n4832), .ZN(n4833)
         );
  AOI21_X1 U5982 ( .B1(n6956), .B2(n4909), .A(n4833), .ZN(n4835) );
  NAND2_X1 U5983 ( .A1(n4910), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4834)
         );
  OAI211_X1 U5984 ( .C1(n4914), .C2(n4872), .A(n4835), .B(n4834), .ZN(U3144)
         );
  INV_X1 U5985 ( .A(n4885), .ZN(n4839) );
  AND2_X1 U5986 ( .A1(n3196), .A2(n4836), .ZN(n4837) );
  NAND2_X1 U5987 ( .A1(n4838), .A2(n4837), .ZN(n6974) );
  AOI21_X1 U5988 ( .B1(n4839), .B2(n6974), .A(n6414), .ZN(n4840) );
  AOI211_X1 U5989 ( .C1(n4842), .C2(n4841), .A(n6927), .B(n4840), .ZN(n4846)
         );
  NOR2_X1 U5990 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4843), .ZN(n4886)
         );
  OAI211_X1 U5991 ( .C1(n3454), .C2(n4886), .A(n6860), .B(n4844), .ZN(n4845)
         );
  INV_X1 U5992 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4855) );
  INV_X1 U5993 ( .A(n4847), .ZN(n4848) );
  AOI22_X1 U5994 ( .A1(n4850), .A2(n4173), .B1(n4849), .B2(n4848), .ZN(n4888)
         );
  AOI22_X1 U5995 ( .A1(n6920), .A2(n4886), .B1(n6919), .B2(n4885), .ZN(n4851)
         );
  OAI21_X1 U5996 ( .B1(n4852), .B2(n4888), .A(n4851), .ZN(n4853) );
  AOI21_X1 U5997 ( .B1(n6864), .B2(n6976), .A(n4853), .ZN(n4854) );
  OAI21_X1 U5998 ( .B1(n4893), .B2(n4855), .A(n4854), .ZN(U3116) );
  INV_X1 U5999 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4860) );
  AOI22_X1 U6000 ( .A1(n6939), .A2(n4886), .B1(n6938), .B2(n4885), .ZN(n4856)
         );
  OAI21_X1 U6001 ( .B1(n4857), .B2(n4888), .A(n4856), .ZN(n4858) );
  AOI21_X1 U6002 ( .B1(n6868), .B2(n6976), .A(n4858), .ZN(n4859) );
  OAI21_X1 U6003 ( .B1(n4893), .B2(n4860), .A(n4859), .ZN(U3117) );
  INV_X1 U6004 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4865) );
  AOI22_X1 U6005 ( .A1(n6951), .A2(n4886), .B1(n6901), .B2(n4885), .ZN(n4861)
         );
  OAI21_X1 U6006 ( .B1(n4862), .B2(n4888), .A(n4861), .ZN(n4863) );
  AOI21_X1 U6007 ( .B1(n6950), .B2(n6976), .A(n4863), .ZN(n4864) );
  OAI21_X1 U6008 ( .B1(n4893), .B2(n4865), .A(n4864), .ZN(U3119) );
  INV_X1 U6009 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4870) );
  AOI22_X1 U6010 ( .A1(n6979), .A2(n4886), .B1(n6977), .B2(n4885), .ZN(n4866)
         );
  OAI21_X1 U6011 ( .B1(n4867), .B2(n4888), .A(n4866), .ZN(n4868) );
  AOI21_X1 U6012 ( .B1(n6889), .B2(n6976), .A(n4868), .ZN(n4869) );
  OAI21_X1 U6013 ( .B1(n4893), .B2(n4870), .A(n4869), .ZN(U3123) );
  INV_X1 U6014 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4875) );
  AOI22_X1 U6015 ( .A1(n6957), .A2(n4886), .B1(n6905), .B2(n4885), .ZN(n4871)
         );
  OAI21_X1 U6016 ( .B1(n4872), .B2(n4888), .A(n4871), .ZN(n4873) );
  AOI21_X1 U6017 ( .B1(n6956), .B2(n6976), .A(n4873), .ZN(n4874) );
  OAI21_X1 U6018 ( .B1(n4893), .B2(n4875), .A(n4874), .ZN(U3120) );
  INV_X1 U6019 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4880) );
  AOI22_X1 U6020 ( .A1(n6945), .A2(n4886), .B1(n6944), .B2(n4885), .ZN(n4876)
         );
  OAI21_X1 U6021 ( .B1(n4877), .B2(n4888), .A(n4876), .ZN(n4878) );
  AOI21_X1 U6022 ( .B1(n6872), .B2(n6976), .A(n4878), .ZN(n4879) );
  OAI21_X1 U6023 ( .B1(n4893), .B2(n4880), .A(n4879), .ZN(U3118) );
  INV_X1 U6024 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4884) );
  AOI22_X1 U6025 ( .A1(n6970), .A2(n4886), .B1(n6841), .B2(n4885), .ZN(n4881)
         );
  OAI21_X1 U6026 ( .B1(n4913), .B2(n4888), .A(n4881), .ZN(n4882) );
  AOI21_X1 U6027 ( .B1(n6968), .B2(n6976), .A(n4882), .ZN(n4883) );
  OAI21_X1 U6028 ( .B1(n4893), .B2(n4884), .A(n4883), .ZN(U3122) );
  INV_X1 U6029 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4892) );
  AOI22_X1 U6030 ( .A1(n6963), .A2(n4886), .B1(n6962), .B2(n4885), .ZN(n4887)
         );
  OAI21_X1 U6031 ( .B1(n4889), .B2(n4888), .A(n4887), .ZN(n4890) );
  AOI21_X1 U6032 ( .B1(n6880), .B2(n6976), .A(n4890), .ZN(n4891) );
  OAI21_X1 U6033 ( .B1(n4893), .B2(n4892), .A(n4891), .ZN(U3121) );
  NAND2_X1 U6034 ( .A1(n4895), .A2(n4894), .ZN(n4896) );
  NAND2_X1 U6035 ( .A1(n4956), .A2(n4896), .ZN(n6474) );
  INV_X1 U6036 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5678) );
  OAI222_X1 U6037 ( .A1(n6474), .A2(n6060), .B1(n6063), .B2(n5678), .C1(n6058), 
        .C2(n6476), .ZN(U2849) );
  AND2_X1 U6038 ( .A1(n4898), .A2(n4897), .ZN(n4900) );
  OR2_X1 U6039 ( .A1(n5046), .A2(n4901), .ZN(n4902) );
  NAND2_X1 U6040 ( .A1(n4903), .A2(n4902), .ZN(n6446) );
  AOI22_X1 U6041 ( .A1(n5004), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6561), .ZN(n4904) );
  OAI21_X1 U6042 ( .B1(n6446), .B2(n6345), .A(n4904), .ZN(U2877) );
  OAI22_X1 U6043 ( .A1(n4907), .A2(n6975), .B1(n4906), .B2(n4905), .ZN(n4908)
         );
  AOI21_X1 U6044 ( .B1(n6968), .B2(n4909), .A(n4908), .ZN(n4912) );
  NAND2_X1 U6045 ( .A1(n4910), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4911)
         );
  OAI211_X1 U6046 ( .C1(n4914), .C2(n4913), .A(n4912), .B(n4911), .ZN(U3146)
         );
  INV_X1 U6047 ( .A(n4915), .ZN(n4916) );
  NOR2_X1 U6048 ( .A1(n7000), .A2(n4920), .ZN(n4941) );
  AOI21_X1 U6049 ( .B1(n4916), .B2(n6995), .A(n4941), .ZN(n4921) );
  OR2_X1 U6050 ( .A1(n4923), .A2(n6414), .ZN(n4917) );
  AOI22_X1 U6051 ( .A1(n4921), .A2(n4919), .B1(n6927), .B2(n4920), .ZN(n4918)
         );
  NAND2_X1 U6052 ( .A1(n6814), .A2(n4918), .ZN(n4940) );
  INV_X1 U6053 ( .A(n4919), .ZN(n4922) );
  OAI22_X1 U6054 ( .A1(n4922), .A2(n4921), .B1(n6930), .B2(n4920), .ZN(n4939)
         );
  AOI22_X1 U6055 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4940), .B1(n6934), 
        .B2(n4939), .ZN(n4925) );
  NOR2_X2 U6056 ( .A1(n4923), .A2(n6817), .ZN(n5087) );
  AOI22_X1 U6057 ( .A1(n6920), .A2(n4941), .B1(n6919), .B2(n5087), .ZN(n4924)
         );
  OAI211_X1 U6058 ( .C1(n6937), .C2(n4944), .A(n4925), .B(n4924), .ZN(U3028)
         );
  AOI22_X1 U6059 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4940), .B1(n6981), 
        .B2(n4939), .ZN(n4927) );
  AOI22_X1 U6060 ( .A1(n6979), .A2(n4941), .B1(n6977), .B2(n5087), .ZN(n4926)
         );
  OAI211_X1 U6061 ( .C1(n6986), .C2(n4944), .A(n4927), .B(n4926), .ZN(U3035)
         );
  AOI22_X1 U6062 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4940), .B1(n6946), 
        .B2(n4939), .ZN(n4929) );
  AOI22_X1 U6063 ( .A1(n6945), .A2(n4941), .B1(n6944), .B2(n5087), .ZN(n4928)
         );
  OAI211_X1 U6064 ( .C1(n6949), .C2(n4944), .A(n4929), .B(n4928), .ZN(U3030)
         );
  AOI22_X1 U6065 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4940), .B1(n6971), 
        .B2(n4939), .ZN(n4931) );
  AOI22_X1 U6066 ( .A1(n6970), .A2(n4941), .B1(n6841), .B2(n5087), .ZN(n4930)
         );
  OAI211_X1 U6067 ( .C1(n4932), .C2(n4944), .A(n4931), .B(n4930), .ZN(U3034)
         );
  AOI22_X1 U6068 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4940), .B1(n6958), 
        .B2(n4939), .ZN(n4934) );
  AOI22_X1 U6069 ( .A1(n6957), .A2(n4941), .B1(n6905), .B2(n5087), .ZN(n4933)
         );
  OAI211_X1 U6070 ( .C1(n6908), .C2(n4944), .A(n4934), .B(n4933), .ZN(U3032)
         );
  AOI22_X1 U6071 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4940), .B1(n6940), 
        .B2(n4939), .ZN(n4936) );
  AOI22_X1 U6072 ( .A1(n6939), .A2(n4941), .B1(n6938), .B2(n5087), .ZN(n4935)
         );
  OAI211_X1 U6073 ( .C1(n6943), .C2(n4944), .A(n4936), .B(n4935), .ZN(U3029)
         );
  AOI22_X1 U6074 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4940), .B1(n6952), 
        .B2(n4939), .ZN(n4938) );
  AOI22_X1 U6075 ( .A1(n6951), .A2(n4941), .B1(n6901), .B2(n5087), .ZN(n4937)
         );
  OAI211_X1 U6076 ( .C1(n6904), .C2(n4944), .A(n4938), .B(n4937), .ZN(U3031)
         );
  AOI22_X1 U6077 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4940), .B1(n6964), 
        .B2(n4939), .ZN(n4943) );
  AOI22_X1 U6078 ( .A1(n6963), .A2(n4941), .B1(n6962), .B2(n5087), .ZN(n4942)
         );
  OAI211_X1 U6079 ( .C1(n6967), .C2(n4944), .A(n4943), .B(n4942), .ZN(U3033)
         );
  INV_X1 U6080 ( .A(n4945), .ZN(n6396) );
  INV_X1 U6081 ( .A(REIP_REG_10__SCAN_IN), .ZN(n7089) );
  INV_X1 U6082 ( .A(REIP_REG_8__SCAN_IN), .ZN(n7085) );
  INV_X1 U6083 ( .A(REIP_REG_6__SCAN_IN), .ZN(n7082) );
  INV_X1 U6084 ( .A(REIP_REG_4__SCAN_IN), .ZN(n7079) );
  NAND3_X1 U6085 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5012) );
  NOR2_X1 U6086 ( .A1(n7079), .A2(n5012), .ZN(n6531) );
  NAND2_X1 U6087 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6531), .ZN(n6506) );
  NOR2_X1 U6088 ( .A1(n7082), .A2(n6506), .ZN(n6495) );
  NAND2_X1 U6089 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6495), .ZN(n5151) );
  NOR2_X1 U6090 ( .A1(n7085), .A2(n5151), .ZN(n5144) );
  NAND2_X1 U6091 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5144), .ZN(n6472) );
  NOR2_X1 U6092 ( .A1(n7089), .A2(n6472), .ZN(n4958) );
  NAND2_X1 U6093 ( .A1(REIP_REG_11__SCAN_IN), .A2(n4958), .ZN(n4960) );
  NOR2_X1 U6094 ( .A1(n6507), .A2(n4960), .ZN(n6452) );
  INV_X1 U6095 ( .A(n6452), .ZN(n6440) );
  NAND3_X1 U6096 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n4947) );
  NOR2_X1 U6097 ( .A1(n6440), .A2(n4947), .ZN(n4991) );
  INV_X1 U6098 ( .A(n4991), .ZN(n4946) );
  OAI22_X1 U6099 ( .A1(n4946), .A2(REIP_REG_15__SCAN_IN), .B1(n6173), .B2(
        n6541), .ZN(n4952) );
  INV_X1 U6100 ( .A(n6525), .ZN(n5990) );
  NOR2_X1 U6101 ( .A1(n4960), .A2(n4947), .ZN(n5910) );
  OR2_X1 U6102 ( .A1(n6507), .A2(n5910), .ZN(n4948) );
  AND2_X1 U6103 ( .A1(n4948), .A2(n6504), .ZN(n6450) );
  INV_X1 U6104 ( .A(n6450), .ZN(n4990) );
  AOI22_X1 U6105 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6543), .B1(
        REIP_REG_15__SCAN_IN), .B2(n4990), .ZN(n4950) );
  NAND2_X1 U6106 ( .A1(n6504), .A2(n4949), .ZN(n6511) );
  OAI211_X1 U6107 ( .C1(n5990), .C2(n5820), .A(n4950), .B(n6511), .ZN(n4951)
         );
  AOI211_X1 U6108 ( .C1(n6396), .C2(n6539), .A(n4952), .B(n4951), .ZN(n4953)
         );
  OAI21_X1 U6109 ( .B1(n6177), .B2(n6515), .A(n4953), .ZN(U2812) );
  OR2_X1 U6110 ( .A1(n4999), .A2(n4955), .ZN(n5001) );
  INV_X1 U6111 ( .A(n5001), .ZN(n4954) );
  AOI21_X1 U6112 ( .B1(n4955), .B2(n4999), .A(n4954), .ZN(n5103) );
  INV_X1 U6113 ( .A(n5103), .ZN(n4967) );
  AOI21_X1 U6114 ( .B1(n4957), .B2(n4956), .A(n5053), .ZN(n6707) );
  NAND3_X1 U6115 ( .A1(n6532), .A2(n4960), .A3(n4958), .ZN(n4959) );
  OAI21_X1 U6116 ( .B1(n6541), .B2(n5101), .A(n4959), .ZN(n4963) );
  INV_X1 U6117 ( .A(n6504), .ZN(n5030) );
  OAI21_X1 U6118 ( .B1(n5030), .B2(n4960), .A(n5915), .ZN(n6465) );
  INV_X1 U6119 ( .A(REIP_REG_11__SCAN_IN), .ZN(n7087) );
  AOI22_X1 U6120 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6543), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n6525), .ZN(n4961) );
  OAI211_X1 U6121 ( .C1(n6465), .C2(n7087), .A(n4961), .B(n6511), .ZN(n4962)
         );
  AOI211_X1 U6122 ( .C1(n6707), .C2(n6539), .A(n4963), .B(n4962), .ZN(n4964)
         );
  OAI21_X1 U6123 ( .B1(n4967), .B2(n6515), .A(n4964), .ZN(U2816) );
  AOI22_X1 U6124 ( .A1(n6707), .A2(n6056), .B1(EBX_REG_11__SCAN_IN), .B2(n6055), .ZN(n4965) );
  OAI21_X1 U6125 ( .B1(n4967), .B2(n6058), .A(n4965), .ZN(U2848) );
  AOI22_X1 U6126 ( .A1(n5004), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6561), .ZN(n4966) );
  OAI21_X1 U6127 ( .B1(n4967), .B2(n6345), .A(n4966), .ZN(U2880) );
  OR2_X1 U6128 ( .A1(n5055), .A2(n4968), .ZN(n4969) );
  NAND2_X1 U6129 ( .A1(n3211), .A2(n4969), .ZN(n6442) );
  INV_X1 U6130 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6441) );
  OAI222_X1 U6131 ( .A1(n6442), .A2(n6060), .B1(n6063), .B2(n6441), .C1(n6058), 
        .C2(n6446), .ZN(U2845) );
  AOI22_X1 U6132 ( .A1(n5485), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4974) );
  AOI22_X1 U6133 ( .A1(n5333), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4973) );
  AOI22_X1 U6134 ( .A1(n5307), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4972) );
  AOI22_X1 U6135 ( .A1(n5480), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4971) );
  NAND4_X1 U6136 ( .A1(n4974), .A2(n4973), .A3(n4972), .A4(n4971), .ZN(n4980)
         );
  AOI22_X1 U6137 ( .A1(n5476), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5460), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4978) );
  AOI22_X1 U6138 ( .A1(n5486), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4977) );
  AOI22_X1 U6139 ( .A1(n5332), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4976) );
  AOI22_X1 U6140 ( .A1(n5221), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4975) );
  NAND4_X1 U6141 ( .A1(n4978), .A2(n4977), .A3(n4976), .A4(n4975), .ZN(n4979)
         );
  OR2_X1 U6142 ( .A1(n4980), .A2(n4979), .ZN(n4984) );
  XNOR2_X1 U6143 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4981), .ZN(n6168)
         );
  AOI22_X1 U6144 ( .A1(n5509), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n5506), 
        .B2(n6168), .ZN(n4982) );
  OAI21_X1 U6145 ( .B1(n5369), .B2(n5665), .A(n4982), .ZN(n4983) );
  AOI21_X1 U6146 ( .B1(n5467), .B2(n4984), .A(n4983), .ZN(n4985) );
  AND2_X1 U6147 ( .A1(n4986), .A2(n4985), .ZN(n4987) );
  NOR2_X1 U6148 ( .A1(n5140), .A2(n4987), .ZN(n6560) );
  INV_X1 U6149 ( .A(n6560), .ZN(n5116) );
  NAND2_X1 U6150 ( .A1(n3201), .A2(n4988), .ZN(n4989) );
  NAND2_X1 U6151 ( .A1(n5119), .A2(n4989), .ZN(n6385) );
  INV_X1 U6152 ( .A(n6385), .ZN(n4996) );
  INV_X1 U6153 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5117) );
  OAI22_X1 U6154 ( .A1(n6522), .A2(n5117), .B1(n6168), .B2(n6541), .ZN(n4995)
         );
  NAND2_X1 U6155 ( .A1(REIP_REG_15__SCAN_IN), .A2(n4991), .ZN(n5208) );
  INV_X1 U6156 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7099) );
  INV_X1 U6157 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7097) );
  AOI21_X1 U6158 ( .B1(n4991), .B2(n7097), .A(n4990), .ZN(n4993) );
  AOI21_X1 U6159 ( .B1(n6525), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6524), 
        .ZN(n4992) );
  OAI221_X1 U6160 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5208), .C1(n7099), .C2(
        n4993), .A(n4992), .ZN(n4994) );
  AOI211_X1 U6161 ( .C1(n4996), .C2(n6539), .A(n4995), .B(n4994), .ZN(n4997)
         );
  OAI21_X1 U6162 ( .B1(n5116), .B2(n6515), .A(n4997), .ZN(U2811) );
  OR2_X1 U6163 ( .A1(n4999), .A2(n4998), .ZN(n5045) );
  INV_X1 U6164 ( .A(n5045), .ZN(n5000) );
  AOI21_X1 U6165 ( .B1(n5002), .B2(n5001), .A(n5000), .ZN(n6664) );
  INV_X1 U6166 ( .A(n6664), .ZN(n5006) );
  XNOR2_X1 U6167 ( .A(n5053), .B(n5049), .ZN(n6467) );
  AOI22_X1 U6168 ( .A1(n6467), .A2(n6056), .B1(n6055), .B2(EBX_REG_12__SCAN_IN), .ZN(n5003) );
  OAI21_X1 U6169 ( .B1(n5006), .B2(n6058), .A(n5003), .ZN(U2847) );
  AOI22_X1 U6170 ( .A1(n5004), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n6561), .ZN(n5005) );
  OAI21_X1 U6171 ( .B1(n5006), .B2(n6345), .A(n5005), .ZN(U2879) );
  NAND2_X1 U6172 ( .A1(n6518), .A2(n5007), .ZN(n5008) );
  OAI211_X1 U6173 ( .C1(n6527), .C2(n6776), .A(n5008), .B(n6511), .ZN(n5010)
         );
  NOR3_X1 U6174 ( .A1(n6507), .A2(REIP_REG_4__SCAN_IN), .A3(n5012), .ZN(n5009)
         );
  AOI211_X1 U6175 ( .C1(n6543), .C2(EBX_REG_4__SCAN_IN), .A(n5010), .B(n5009), 
        .ZN(n5011) );
  OAI21_X1 U6176 ( .B1(n6545), .B2(n6402), .A(n5011), .ZN(n5015) );
  OAI21_X1 U6177 ( .B1(n5030), .B2(n5012), .A(n5915), .ZN(n6551) );
  OAI22_X1 U6178 ( .A1(n6551), .A2(n7079), .B1(n5013), .B2(n5990), .ZN(n5014)
         );
  AOI211_X1 U6179 ( .C1(n5016), .C2(n6548), .A(n5015), .B(n5014), .ZN(n5017)
         );
  INV_X1 U6180 ( .A(n5017), .ZN(U2823) );
  INV_X1 U6181 ( .A(n5094), .ZN(n5021) );
  AOI21_X1 U6182 ( .B1(n5019), .B2(n5093), .A(n5018), .ZN(n5020) );
  AOI21_X1 U6183 ( .B1(n5021), .B2(n5093), .A(n5020), .ZN(n5039) );
  INV_X1 U6184 ( .A(n5039), .ZN(n5028) );
  INV_X1 U6185 ( .A(n6750), .ZN(n6383) );
  AOI22_X1 U6186 ( .A1(n6241), .A2(n5023), .B1(n6743), .B2(n5022), .ZN(n6742)
         );
  OAI21_X1 U6187 ( .B1(n6727), .B2(n6383), .A(n6742), .ZN(n6715) );
  NOR2_X1 U6188 ( .A1(n6474), .A2(n6775), .ZN(n5026) );
  NOR2_X1 U6189 ( .A1(n6744), .A2(n6804), .ZN(n6763) );
  NOR2_X1 U6190 ( .A1(n6746), .A2(n6763), .ZN(n6779) );
  NOR3_X1 U6191 ( .A1(n6779), .A2(n6749), .A3(n6751), .ZN(n6758) );
  NAND2_X1 U6192 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6758), .ZN(n6726)
         );
  INV_X1 U6193 ( .A(n6726), .ZN(n6738) );
  AND2_X1 U6194 ( .A1(n6727), .A2(n6738), .ZN(n6720) );
  OAI221_X1 U6195 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n6724), .C2(n5891), .A(n6720), 
        .ZN(n5024) );
  OAI21_X1 U6196 ( .B1(n6774), .B2(n7089), .A(n5024), .ZN(n5025) );
  AOI211_X1 U6197 ( .C1(n6715), .C2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5026), .B(n5025), .ZN(n5027) );
  OAI21_X1 U6198 ( .B1(n5028), .B2(n6773), .A(n5027), .ZN(U3008) );
  AOI22_X1 U6199 ( .A1(n5030), .A2(REIP_REG_1__SCAN_IN), .B1(n6539), .B2(n5029), .ZN(n5031) );
  OAI21_X1 U6200 ( .B1(n6541), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5031), 
        .ZN(n5032) );
  AOI21_X1 U6201 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6525), .A(n5032), 
        .ZN(n5034) );
  OAI211_X1 U6202 ( .C1(n6522), .C2(n4167), .A(n5034), .B(n5033), .ZN(n5035)
         );
  AOI21_X1 U6203 ( .B1(n4027), .B2(n5036), .A(n5035), .ZN(n5037) );
  OAI21_X1 U6204 ( .B1(n5038), .B2(n6528), .A(n5037), .ZN(U2826) );
  NAND2_X1 U6205 ( .A1(n5039), .A2(n6700), .ZN(n5043) );
  INV_X1 U6206 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5040) );
  OAI22_X1 U6207 ( .A1(n6162), .A2(n5040), .B1(n6774), .B2(n7089), .ZN(n5041)
         );
  AOI21_X1 U6208 ( .B1(n6663), .B2(n6477), .A(n5041), .ZN(n5042) );
  OAI211_X1 U6209 ( .C1(n6679), .C2(n6476), .A(n5043), .B(n5042), .ZN(U2976)
         );
  AND2_X1 U6210 ( .A1(n5045), .A2(n5044), .ZN(n5047) );
  INV_X1 U6211 ( .A(DATAI_13_), .ZN(n6652) );
  INV_X1 U6212 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6575) );
  OAI222_X1 U6213 ( .A1(n6458), .A2(n6345), .B1(n5048), .B2(n6652), .C1(n6064), 
        .C2(n6575), .ZN(U2878) );
  INV_X1 U6214 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5056) );
  INV_X1 U6215 ( .A(n5049), .ZN(n5052) );
  INV_X1 U6216 ( .A(n5050), .ZN(n5051) );
  AOI21_X1 U6217 ( .B1(n5053), .B2(n5052), .A(n5051), .ZN(n5054) );
  OR2_X1 U6218 ( .A1(n5055), .A2(n5054), .ZN(n6275) );
  OAI222_X1 U6219 ( .A1(n6458), .A2(n6058), .B1(n6063), .B2(n5056), .C1(n6275), 
        .C2(n6060), .ZN(U2846) );
  NOR2_X1 U6220 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5057), .ZN(n5086)
         );
  OAI21_X1 U6221 ( .B1(n5087), .B2(n5085), .A(n6858), .ZN(n5058) );
  NAND2_X1 U6222 ( .A1(n5058), .A2(n5063), .ZN(n5060) );
  OAI221_X1 U6223 ( .B1(n5086), .B2(n3454), .C1(n5086), .C2(n5060), .A(n5059), 
        .ZN(n5061) );
  INV_X1 U6224 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5066) );
  AOI22_X1 U6225 ( .A1(n6939), .A2(n5086), .B1(n6938), .B2(n5085), .ZN(n5065)
         );
  NAND2_X1 U6226 ( .A1(n5062), .A2(n7016), .ZN(n6853) );
  OAI22_X1 U6227 ( .A1(n5063), .A2(n6927), .B1(n6860), .B2(n6853), .ZN(n5088)
         );
  AOI22_X1 U6228 ( .A1(n6940), .A2(n5088), .B1(n6868), .B2(n5087), .ZN(n5064)
         );
  OAI211_X1 U6229 ( .C1(n5092), .C2(n5066), .A(n5065), .B(n5064), .ZN(U3037)
         );
  INV_X1 U6230 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5069) );
  AOI22_X1 U6231 ( .A1(n6920), .A2(n5086), .B1(n6919), .B2(n5085), .ZN(n5068)
         );
  AOI22_X1 U6232 ( .A1(n6934), .A2(n5088), .B1(n6864), .B2(n5087), .ZN(n5067)
         );
  OAI211_X1 U6233 ( .C1(n5092), .C2(n5069), .A(n5068), .B(n5067), .ZN(U3036)
         );
  INV_X1 U6234 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5072) );
  AOI22_X1 U6235 ( .A1(n6979), .A2(n5086), .B1(n6977), .B2(n5085), .ZN(n5071)
         );
  AOI22_X1 U6236 ( .A1(n6981), .A2(n5088), .B1(n6889), .B2(n5087), .ZN(n5070)
         );
  OAI211_X1 U6237 ( .C1(n5092), .C2(n5072), .A(n5071), .B(n5070), .ZN(U3043)
         );
  INV_X1 U6238 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5075) );
  AOI22_X1 U6239 ( .A1(n6951), .A2(n5086), .B1(n6901), .B2(n5085), .ZN(n5074)
         );
  AOI22_X1 U6240 ( .A1(n6952), .A2(n5088), .B1(n6950), .B2(n5087), .ZN(n5073)
         );
  OAI211_X1 U6241 ( .C1(n5092), .C2(n5075), .A(n5074), .B(n5073), .ZN(U3039)
         );
  INV_X1 U6242 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5078) );
  AOI22_X1 U6243 ( .A1(n6945), .A2(n5086), .B1(n6944), .B2(n5085), .ZN(n5077)
         );
  AOI22_X1 U6244 ( .A1(n6946), .A2(n5088), .B1(n6872), .B2(n5087), .ZN(n5076)
         );
  OAI211_X1 U6245 ( .C1(n5092), .C2(n5078), .A(n5077), .B(n5076), .ZN(U3038)
         );
  INV_X1 U6246 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5081) );
  AOI22_X1 U6247 ( .A1(n6963), .A2(n5086), .B1(n6962), .B2(n5085), .ZN(n5080)
         );
  AOI22_X1 U6248 ( .A1(n6964), .A2(n5088), .B1(n6880), .B2(n5087), .ZN(n5079)
         );
  OAI211_X1 U6249 ( .C1(n5092), .C2(n5081), .A(n5080), .B(n5079), .ZN(U3041)
         );
  INV_X1 U6250 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5084) );
  AOI22_X1 U6251 ( .A1(n6970), .A2(n5086), .B1(n6841), .B2(n5085), .ZN(n5083)
         );
  AOI22_X1 U6252 ( .A1(n6971), .A2(n5088), .B1(n6968), .B2(n5087), .ZN(n5082)
         );
  OAI211_X1 U6253 ( .C1(n5092), .C2(n5084), .A(n5083), .B(n5082), .ZN(U3042)
         );
  INV_X1 U6254 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5091) );
  AOI22_X1 U6255 ( .A1(n6957), .A2(n5086), .B1(n6905), .B2(n5085), .ZN(n5090)
         );
  AOI22_X1 U6256 ( .A1(n6958), .A2(n5088), .B1(n6956), .B2(n5087), .ZN(n5089)
         );
  OAI211_X1 U6257 ( .C1(n5092), .C2(n5091), .A(n5090), .B(n5089), .ZN(U3040)
         );
  AND2_X1 U6258 ( .A1(n5094), .A2(n5093), .ZN(n5099) );
  INV_X1 U6259 ( .A(n5095), .ZN(n5097) );
  NAND2_X1 U6260 ( .A1(n5097), .A2(n5096), .ZN(n5098) );
  XNOR2_X1 U6261 ( .A(n5099), .B(n5098), .ZN(n6708) );
  NAND2_X1 U6262 ( .A1(n6803), .A2(REIP_REG_11__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U6263 ( .A1(n6694), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5100)
         );
  OAI211_X1 U6264 ( .C1(n6704), .C2(n5101), .A(n6705), .B(n5100), .ZN(n5102)
         );
  AOI21_X1 U6265 ( .B1(n5103), .B2(n6698), .A(n5102), .ZN(n5104) );
  OAI21_X1 U6266 ( .B1(n6708), .B2(n6681), .A(n5104), .ZN(U2975) );
  XNOR2_X1 U6267 ( .A(n6262), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5106)
         );
  XNOR2_X1 U6268 ( .A(n5105), .B(n5106), .ZN(n6667) );
  INV_X1 U6269 ( .A(n5262), .ZN(n5109) );
  INV_X1 U6270 ( .A(n5107), .ZN(n5108) );
  AOI21_X1 U6271 ( .B1(n5109), .B2(n6241), .A(n5108), .ZN(n6709) );
  NOR2_X1 U6272 ( .A1(n5262), .A2(n5110), .ZN(n6390) );
  INV_X1 U6273 ( .A(n6390), .ZN(n6272) );
  NAND2_X1 U6274 ( .A1(n5256), .A2(n6272), .ZN(n6712) );
  AOI21_X1 U6275 ( .B1(n6709), .B2(n6712), .A(n5841), .ZN(n5114) );
  INV_X1 U6276 ( .A(REIP_REG_12__SCAN_IN), .ZN(n7092) );
  NAND3_X1 U6277 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5841), .A3(n6272), .ZN(n5112) );
  NAND2_X1 U6278 ( .A1(n6467), .A2(n6799), .ZN(n5111) );
  OAI211_X1 U6279 ( .C1(n7092), .C2(n6774), .A(n5112), .B(n5111), .ZN(n5113)
         );
  NOR2_X1 U6280 ( .A1(n5114), .A2(n5113), .ZN(n5115) );
  OAI21_X1 U6281 ( .B1(n6667), .B2(n6773), .A(n5115), .ZN(U3006) );
  OAI222_X1 U6282 ( .A1(n5117), .A2(n6063), .B1(n6060), .B2(n6385), .C1(n5116), 
        .C2(n6058), .ZN(U2843) );
  AND2_X1 U6283 ( .A1(n5119), .A2(n5118), .ZN(n5120) );
  OR2_X1 U6284 ( .A1(n5120), .A2(n5159), .ZN(n6431) );
  INV_X1 U6285 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6286 ( .A1(n5503), .A2(n5499), .ZN(n5283) );
  AOI22_X1 U6287 ( .A1(n5478), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6288 ( .A1(n5476), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6289 ( .A1(n5338), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5121) );
  AND3_X1 U6290 ( .A1(n5122), .A2(n5499), .A3(n5121), .ZN(n5125) );
  AOI22_X1 U6291 ( .A1(n5475), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5124) );
  AOI22_X1 U6292 ( .A1(n5438), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5123) );
  NAND4_X1 U6293 ( .A1(n5126), .A2(n5125), .A3(n5124), .A4(n5123), .ZN(n5132)
         );
  AOI22_X1 U6294 ( .A1(n5332), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5307), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n5130) );
  AOI22_X1 U6295 ( .A1(n5485), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5486), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n5129) );
  AOI22_X1 U6296 ( .A1(n5333), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5128) );
  AOI22_X1 U6297 ( .A1(n5221), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5127) );
  NAND4_X1 U6298 ( .A1(n5130), .A2(n5129), .A3(n5128), .A4(n5127), .ZN(n5131)
         );
  OR2_X1 U6299 ( .A1(n5132), .A2(n5131), .ZN(n5133) );
  NAND2_X1 U6300 ( .A1(n5283), .A2(n5133), .ZN(n5139) );
  NOR2_X1 U6301 ( .A1(n5134), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5135) );
  AOI21_X1 U6302 ( .B1(n5501), .B2(EAX_REG_17__SCAN_IN), .A(n5135), .ZN(n5138)
         );
  XNOR2_X1 U6303 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .B(n5136), .ZN(n6430)
         );
  AND2_X1 U6304 ( .A1(n6430), .A2(n5506), .ZN(n5137) );
  AOI21_X1 U6305 ( .B1(n5139), .B2(n5138), .A(n5137), .ZN(n5141) );
  AND2_X2 U6306 ( .A1(n5140), .A2(n5141), .ZN(n5179) );
  NOR2_X1 U6307 ( .A1(n5140), .A2(n5141), .ZN(n5142) );
  OR2_X1 U6308 ( .A1(n5179), .A2(n5142), .ZN(n6432) );
  OAI222_X1 U6309 ( .A1(n6060), .A2(n6431), .B1(n6063), .B2(n5143), .C1(n6058), 
        .C2(n6432), .ZN(U2842) );
  INV_X1 U6310 ( .A(n5144), .ZN(n6479) );
  NAND2_X1 U6311 ( .A1(n6532), .A2(n6479), .ZN(n5150) );
  NAND2_X1 U6312 ( .A1(n5150), .A2(n6504), .ZN(n6485) );
  NOR2_X1 U6313 ( .A1(n6729), .A2(n6527), .ZN(n5153) );
  OAI21_X1 U6314 ( .B1(n6541), .B2(n5145), .A(n6511), .ZN(n5148) );
  NOR2_X1 U6315 ( .A1(n6522), .A2(n5146), .ZN(n5147) );
  AOI211_X1 U6316 ( .C1(n6525), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5148), 
        .B(n5147), .ZN(n5149) );
  OAI21_X1 U6317 ( .B1(n5151), .B2(n5150), .A(n5149), .ZN(n5152) );
  AOI211_X1 U6318 ( .C1(REIP_REG_8__SCAN_IN), .C2(n6485), .A(n5153), .B(n5152), 
        .ZN(n5154) );
  OAI21_X1 U6319 ( .B1(n5155), .B2(n6515), .A(n5154), .ZN(U2819) );
  MUX2_X1 U6320 ( .A(n5243), .B(n5156), .S(n5537), .Z(n5157) );
  INV_X1 U6321 ( .A(n5157), .ZN(n5158) );
  NAND2_X1 U6322 ( .A1(n5159), .A2(n5158), .ZN(n5205) );
  OR2_X1 U6323 ( .A1(n5159), .A2(n5158), .ZN(n5160) );
  AND2_X1 U6324 ( .A1(n5205), .A2(n5160), .ZN(n6377) );
  INV_X1 U6325 ( .A(n6377), .ZN(n5183) );
  AOI22_X1 U6326 ( .A1(n5478), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n5164) );
  AOI22_X1 U6327 ( .A1(n5333), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5163) );
  AOI22_X1 U6328 ( .A1(n5486), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5162) );
  AOI22_X1 U6329 ( .A1(n5485), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5161) );
  NAND4_X1 U6330 ( .A1(n5164), .A2(n5163), .A3(n5162), .A4(n5161), .ZN(n5170)
         );
  AOI22_X1 U6331 ( .A1(n5332), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5168) );
  AOI22_X1 U6332 ( .A1(n5307), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5460), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5167) );
  AOI22_X1 U6333 ( .A1(n5221), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5166) );
  AOI22_X1 U6334 ( .A1(n5338), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5165) );
  NAND4_X1 U6335 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n5169)
         );
  NOR2_X1 U6336 ( .A1(n5170), .A2(n5169), .ZN(n5174) );
  OAI21_X1 U6337 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6414), .A(n6930), 
        .ZN(n5171) );
  INV_X1 U6338 ( .A(n5171), .ZN(n5172) );
  AOI21_X1 U6339 ( .B1(n5501), .B2(EAX_REG_18__SCAN_IN), .A(n5172), .ZN(n5173)
         );
  OAI21_X1 U6340 ( .B1(n5503), .B2(n5174), .A(n5173), .ZN(n5177) );
  OAI21_X1 U6341 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5175), .A(n5198), 
        .ZN(n6362) );
  OR2_X1 U6342 ( .A1(n5499), .A2(n6362), .ZN(n5176) );
  OR2_X1 U6343 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  AND2_X1 U6344 ( .A1(n5203), .A2(n5180), .ZN(n6552) );
  INV_X1 U6345 ( .A(n6552), .ZN(n5181) );
  OAI222_X1 U6346 ( .A1(n6060), .A2(n5183), .B1(n6063), .B2(n5182), .C1(n6058), 
        .C2(n5181), .ZN(U2841) );
  AOI22_X1 U6347 ( .A1(n5307), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5187) );
  AOI22_X1 U6348 ( .A1(n5478), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5186) );
  AOI22_X1 U6349 ( .A1(n5333), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5185) );
  AOI22_X1 U6350 ( .A1(n5476), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5184) );
  NAND4_X1 U6351 ( .A1(n5187), .A2(n5186), .A3(n5185), .A4(n5184), .ZN(n5195)
         );
  AOI22_X1 U6352 ( .A1(n3488), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5460), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5193) );
  AOI22_X1 U6353 ( .A1(n5486), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6354 ( .A1(n5485), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U6355 ( .A1(n5338), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5188) );
  AND3_X1 U6356 ( .A1(n5189), .A2(n5499), .A3(n5188), .ZN(n5191) );
  AOI22_X1 U6357 ( .A1(n5480), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5190) );
  NAND4_X1 U6358 ( .A1(n5193), .A2(n5192), .A3(n5191), .A4(n5190), .ZN(n5194)
         );
  OAI21_X1 U6359 ( .B1(n5195), .B2(n5194), .A(n5283), .ZN(n5197) );
  AOI22_X1 U6360 ( .A1(n5510), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6930), .ZN(n5196) );
  NAND2_X1 U6361 ( .A1(n5197), .A2(n5196), .ZN(n5200) );
  XNOR2_X1 U6362 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n5198), .ZN(n6159)
         );
  NAND2_X1 U6363 ( .A1(n6159), .A2(n5506), .ZN(n5199) );
  NAND2_X1 U6364 ( .A1(n5200), .A2(n5199), .ZN(n5202) );
  INV_X1 U6365 ( .A(n5240), .ZN(n5201) );
  AOI21_X1 U6366 ( .B1(n5203), .B2(n5202), .A(n5201), .ZN(n6353) );
  INV_X1 U6367 ( .A(n6353), .ZN(n5214) );
  XNOR2_X1 U6368 ( .A(n5205), .B(n5204), .ZN(n6254) );
  AOI22_X1 U6369 ( .A1(n6254), .A2(n6056), .B1(n6055), .B2(EBX_REG_19__SCAN_IN), .ZN(n5206) );
  OAI21_X1 U6370 ( .B1(n5214), .B2(n6058), .A(n5206), .ZN(U2840) );
  INV_X1 U6371 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6161) );
  AOI22_X1 U6372 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6543), .B1(n6159), .B2(n6518), .ZN(n5207) );
  OAI211_X1 U6373 ( .C1(n5990), .C2(n6161), .A(n5207), .B(n6511), .ZN(n5210)
         );
  INV_X1 U6374 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7101) );
  NOR2_X1 U6375 ( .A1(n7099), .A2(n5208), .ZN(n6435) );
  NAND2_X1 U6376 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6435), .ZN(n6321) );
  NOR3_X1 U6377 ( .A1(REIP_REG_19__SCAN_IN), .A2(n7101), .A3(n6321), .ZN(n5209) );
  AOI211_X1 U6378 ( .C1(n6539), .C2(n6254), .A(n5210), .B(n5209), .ZN(n5213)
         );
  NOR2_X1 U6379 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6321), .ZN(n6021) );
  NAND3_X1 U6380 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5913) );
  INV_X1 U6381 ( .A(n5913), .ZN(n5211) );
  OAI21_X1 U6382 ( .B1(n5211), .B2(n6507), .A(n6450), .ZN(n6434) );
  OAI21_X1 U6383 ( .B1(n6021), .B2(n6434), .A(REIP_REG_19__SCAN_IN), .ZN(n5212) );
  OAI211_X1 U6384 ( .C1(n5214), .C2(n6515), .A(n5213), .B(n5212), .ZN(U2808)
         );
  AOI21_X1 U6385 ( .B1(n5216), .B2(n5215), .A(n3179), .ZN(n6280) );
  INV_X1 U6386 ( .A(n6458), .ZN(n5219) );
  NAND2_X1 U6387 ( .A1(n6785), .A2(REIP_REG_13__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U6388 ( .A1(n6694), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5217)
         );
  OAI211_X1 U6389 ( .C1(n6704), .C2(n6457), .A(n6276), .B(n5217), .ZN(n5218)
         );
  AOI21_X1 U6390 ( .B1(n5219), .B2(n6698), .A(n5218), .ZN(n5220) );
  OAI21_X1 U6391 ( .B1(n6280), .B2(n6681), .A(n5220), .ZN(U2973) );
  AOI22_X1 U6392 ( .A1(n3488), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5225) );
  AOI22_X1 U6393 ( .A1(n5478), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5224) );
  AOI22_X1 U6394 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5480), .B1(n5460), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5223) );
  AOI22_X1 U6395 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5221), .B1(n3421), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5222) );
  NAND4_X1 U6396 ( .A1(n5225), .A2(n5224), .A3(n5223), .A4(n5222), .ZN(n5231)
         );
  AOI22_X1 U6397 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5307), .B1(n5475), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5229) );
  AOI22_X1 U6398 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n5333), .B1(n5477), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5228) );
  AOI22_X1 U6399 ( .A1(n5486), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5227) );
  AOI22_X1 U6400 ( .A1(n3525), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5226) );
  NAND4_X1 U6401 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n5230)
         );
  NOR2_X1 U6402 ( .A1(n5231), .A2(n5230), .ZN(n5235) );
  NAND2_X1 U6403 ( .A1(n6930), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5232)
         );
  NAND2_X1 U6404 ( .A1(n5499), .A2(n5232), .ZN(n5233) );
  AOI21_X1 U6405 ( .B1(n5501), .B2(EAX_REG_20__SCAN_IN), .A(n5233), .ZN(n5234)
         );
  OAI21_X1 U6406 ( .B1(n5503), .B2(n5235), .A(n5234), .ZN(n5238) );
  OAI21_X1 U6407 ( .B1(n5236), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5285), 
        .ZN(n6330) );
  OR2_X1 U6408 ( .A1(n6330), .A2(n5499), .ZN(n5237) );
  NAND2_X1 U6409 ( .A1(n5238), .A2(n5237), .ZN(n5239) );
  AND2_X1 U6410 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  OR2_X1 U6411 ( .A1(n5241), .A2(n5290), .ZN(n6155) );
  MUX2_X1 U6412 ( .A(n5243), .B(n3913), .S(n5242), .Z(n5245) );
  XNOR2_X1 U6413 ( .A(n5245), .B(n5244), .ZN(n6324) );
  OAI222_X1 U6414 ( .A1(n6058), .A2(n6155), .B1(n6063), .B2(n5246), .C1(n6324), 
        .C2(n6060), .ZN(U2839) );
  NAND2_X1 U6415 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  XNOR2_X1 U6416 ( .A(n3190), .B(n5249), .ZN(n5269) );
  INV_X1 U6417 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6418 ( .A1(n6803), .A2(REIP_REG_14__SCAN_IN), .ZN(n5255) );
  OAI21_X1 U6419 ( .B1(n6162), .B2(n5251), .A(n5255), .ZN(n5253) );
  NOR2_X1 U6420 ( .A1(n6446), .A2(n6679), .ZN(n5252) );
  AOI211_X1 U6421 ( .C1(n6663), .C2(n6444), .A(n5253), .B(n5252), .ZN(n5254)
         );
  OAI21_X1 U6422 ( .B1(n5269), .B2(n6681), .A(n5254), .ZN(U2972) );
  NOR2_X1 U6423 ( .A1(n6390), .A2(n6389), .ZN(n5267) );
  OAI21_X1 U6424 ( .B1(n6442), .B2(n6775), .A(n5255), .ZN(n5266) );
  NOR2_X1 U6425 ( .A1(n5256), .A2(n5841), .ZN(n5260) );
  AND2_X1 U6426 ( .A1(n5257), .A2(n5260), .ZN(n6273) );
  NAND2_X1 U6427 ( .A1(n5258), .A2(n6389), .ZN(n5259) );
  OAI211_X1 U6428 ( .C1(n5261), .C2(n5260), .A(n6709), .B(n5259), .ZN(n6274)
         );
  AOI221_X1 U6429 ( .B1(n5263), .B2(n6273), .C1(n5262), .C2(n6273), .A(n6274), 
        .ZN(n5264) );
  NOR2_X1 U6430 ( .A1(n5264), .A2(n6388), .ZN(n5265) );
  AOI211_X1 U6431 ( .C1(n5267), .C2(n6388), .A(n5266), .B(n5265), .ZN(n5268)
         );
  OAI21_X1 U6432 ( .B1(n5269), .B2(n6773), .A(n5268), .ZN(U3004) );
  AOI22_X1 U6433 ( .A1(n5438), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6434 ( .A1(n5485), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6435 ( .A1(n3421), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5270) );
  AND3_X1 U6436 ( .A1(n5271), .A2(n5499), .A3(n5270), .ZN(n5274) );
  AOI22_X1 U6437 ( .A1(n5477), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5273) );
  AOI22_X1 U6438 ( .A1(n5480), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5272) );
  NAND4_X1 U6439 ( .A1(n5275), .A2(n5274), .A3(n5273), .A4(n5272), .ZN(n5281)
         );
  AOI22_X1 U6440 ( .A1(n3488), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5279) );
  AOI22_X1 U6441 ( .A1(n5307), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5278) );
  AOI22_X1 U6442 ( .A1(n5486), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5277) );
  AOI22_X1 U6443 ( .A1(n5333), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3525), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5276) );
  NAND4_X1 U6444 ( .A1(n5279), .A2(n5278), .A3(n5277), .A4(n5276), .ZN(n5280)
         );
  OR2_X1 U6445 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  NAND2_X1 U6446 ( .A1(n5283), .A2(n5282), .ZN(n5288) );
  NOR2_X1 U6447 ( .A1(n6140), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5284) );
  AOI21_X1 U6448 ( .B1(n5501), .B2(EAX_REG_21__SCAN_IN), .A(n5284), .ZN(n5287)
         );
  XNOR2_X1 U6449 ( .A(n5285), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6142)
         );
  AND2_X1 U6450 ( .A1(n6142), .A2(n5506), .ZN(n5286) );
  AOI21_X1 U6451 ( .B1(n5288), .B2(n5287), .A(n5286), .ZN(n5291) );
  AND2_X2 U6452 ( .A1(n5290), .A2(n5291), .ZN(n6003) );
  INV_X1 U6453 ( .A(n6003), .ZN(n5289) );
  OAI21_X1 U6454 ( .B1(n5291), .B2(n5290), .A(n5289), .ZN(n6145) );
  AOI22_X1 U6455 ( .A1(n6558), .A2(DATAI_21_), .B1(n6561), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6456 ( .A1(n6562), .A2(DATAI_5_), .ZN(n5292) );
  OAI211_X1 U6457 ( .C1(n6145), .C2(n6345), .A(n5293), .B(n5292), .ZN(U2870)
         );
  NAND3_X1 U6458 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5912) );
  NOR2_X1 U6459 ( .A1(n5912), .A2(n6321), .ZN(n6011) );
  INV_X1 U6460 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U6461 ( .A1(n6011), .A2(n7107), .ZN(n6006) );
  AND2_X1 U6462 ( .A1(n3209), .A2(n5294), .ZN(n5295) );
  NOR2_X1 U6463 ( .A1(n6008), .A2(n5295), .ZN(n6366) );
  AOI21_X1 U6464 ( .B1(n6532), .B2(n5912), .A(n6434), .ZN(n6325) );
  NOR2_X1 U6465 ( .A1(n6325), .A2(n7107), .ZN(n5298) );
  INV_X1 U6466 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6062) );
  AOI22_X1 U6467 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6525), .B1(n6518), 
        .B2(n6142), .ZN(n5296) );
  OAI21_X1 U6468 ( .B1(n6522), .B2(n6062), .A(n5296), .ZN(n5297) );
  AOI211_X1 U6469 ( .C1(n6366), .C2(n6539), .A(n5298), .B(n5297), .ZN(n5299)
         );
  OAI211_X1 U6470 ( .C1(n6145), .C2(n6515), .A(n6006), .B(n5299), .ZN(U2806)
         );
  AND2_X1 U6471 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5518) );
  AOI22_X1 U6472 ( .A1(n5485), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5306) );
  AOI22_X1 U6473 ( .A1(n5333), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5305) );
  AOI22_X1 U6474 ( .A1(n5475), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5304) );
  AOI22_X1 U6475 ( .A1(n3421), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5303) );
  NAND4_X1 U6476 ( .A1(n5306), .A2(n5305), .A3(n5304), .A4(n5303), .ZN(n5313)
         );
  AOI22_X1 U6477 ( .A1(n5307), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5460), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5311) );
  AOI22_X1 U6478 ( .A1(n5486), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5310) );
  AOI22_X1 U6479 ( .A1(n5332), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5309) );
  AOI22_X1 U6480 ( .A1(n3525), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5308) );
  NAND4_X1 U6481 ( .A1(n5311), .A2(n5310), .A3(n5309), .A4(n5308), .ZN(n5312)
         );
  NOR2_X1 U6482 ( .A1(n5313), .A2(n5312), .ZN(n5317) );
  NAND2_X1 U6483 ( .A1(n6930), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5314)
         );
  NAND2_X1 U6484 ( .A1(n5499), .A2(n5314), .ZN(n5315) );
  AOI21_X1 U6485 ( .B1(n5501), .B2(EAX_REG_22__SCAN_IN), .A(n5315), .ZN(n5316)
         );
  OAI21_X1 U6486 ( .B1(n5503), .B2(n5317), .A(n5316), .ZN(n5321) );
  OR2_X1 U6487 ( .A1(n5318), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5319)
         );
  AND2_X1 U6488 ( .A1(n5364), .A2(n5319), .ZN(n6136) );
  NAND2_X1 U6489 ( .A1(n6136), .A2(n5506), .ZN(n5320) );
  AOI22_X1 U6490 ( .A1(n5485), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5325) );
  AOI22_X1 U6491 ( .A1(n5333), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5324) );
  AOI22_X1 U6492 ( .A1(n5307), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5323) );
  AOI22_X1 U6493 ( .A1(n5332), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5322) );
  NAND4_X1 U6494 ( .A1(n5325), .A2(n5324), .A3(n5323), .A4(n5322), .ZN(n5331)
         );
  AOI22_X1 U6495 ( .A1(n3525), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5329) );
  AOI22_X1 U6496 ( .A1(n5486), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5328) );
  AOI22_X1 U6497 ( .A1(n5438), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5327) );
  AOI22_X1 U6498 ( .A1(n5338), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5326) );
  NAND4_X1 U6499 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), .ZN(n5330)
         );
  NOR2_X1 U6500 ( .A1(n5331), .A2(n5330), .ZN(n5352) );
  AOI22_X1 U6501 ( .A1(n5332), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n5337) );
  AOI22_X1 U6502 ( .A1(n5333), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n5336) );
  AOI22_X1 U6503 ( .A1(n5438), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5335) );
  AOI22_X1 U6504 ( .A1(n3525), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5334) );
  NAND4_X1 U6505 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n5344)
         );
  AOI22_X1 U6506 ( .A1(n5307), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5342) );
  AOI22_X1 U6507 ( .A1(n5478), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n5341) );
  AOI22_X1 U6508 ( .A1(n5221), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5338), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5340) );
  AOI22_X1 U6509 ( .A1(n5486), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5339) );
  NAND4_X1 U6510 ( .A1(n5342), .A2(n5341), .A3(n5340), .A4(n5339), .ZN(n5343)
         );
  NOR2_X1 U6511 ( .A1(n5344), .A2(n5343), .ZN(n5351) );
  XOR2_X1 U6512 ( .A(n5352), .B(n5351), .Z(n5345) );
  NAND2_X1 U6513 ( .A1(n5345), .A2(n5467), .ZN(n5348) );
  OAI21_X1 U6514 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6124), .A(n5499), .ZN(
        n5346) );
  AOI21_X1 U6515 ( .B1(n5501), .B2(EAX_REG_23__SCAN_IN), .A(n5346), .ZN(n5347)
         );
  NAND2_X1 U6516 ( .A1(n5348), .A2(n5347), .ZN(n5350) );
  XNOR2_X1 U6517 ( .A(n5364), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6126)
         );
  NAND2_X1 U6518 ( .A1(n6126), .A2(n5506), .ZN(n5349) );
  NAND2_X1 U6519 ( .A1(n5350), .A2(n5349), .ZN(n5988) );
  NOR2_X1 U6520 ( .A1(n5352), .A2(n5351), .ZN(n5383) );
  AOI22_X1 U6521 ( .A1(n5485), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5356) );
  AOI22_X1 U6522 ( .A1(n5333), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5355) );
  AOI22_X1 U6523 ( .A1(n5307), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n5354) );
  AOI22_X1 U6524 ( .A1(n5332), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n5353) );
  NAND4_X1 U6525 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), .ZN(n5362)
         );
  AOI22_X1 U6526 ( .A1(n3525), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5360) );
  AOI22_X1 U6527 ( .A1(n5486), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5221), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5359) );
  AOI22_X1 U6528 ( .A1(n5438), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5358) );
  AOI22_X1 U6529 ( .A1(n3421), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5357) );
  NAND4_X1 U6530 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), .ZN(n5361)
         );
  OR2_X1 U6531 ( .A1(n5362), .A2(n5361), .ZN(n5382) );
  INV_X1 U6532 ( .A(n5382), .ZN(n5363) );
  XNOR2_X1 U6533 ( .A(n5383), .B(n5363), .ZN(n5371) );
  OAI21_X1 U6534 ( .B1(n5364), .B2(n6124), .A(n5977), .ZN(n5365) );
  NAND2_X1 U6535 ( .A1(n5365), .A2(n5388), .ZN(n5978) );
  NOR2_X1 U6536 ( .A1(n5366), .A2(n5977), .ZN(n5367) );
  AOI21_X1 U6537 ( .B1(n5978), .B2(n5506), .A(n5367), .ZN(n5368) );
  OAI21_X1 U6538 ( .B1(n5369), .B2(n4111), .A(n5368), .ZN(n5370) );
  AOI21_X1 U6539 ( .B1(n5371), .B2(n5467), .A(n5370), .ZN(n5559) );
  AOI22_X1 U6540 ( .A1(n5485), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5375) );
  AOI22_X1 U6541 ( .A1(n5486), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5374) );
  AOI22_X1 U6542 ( .A1(n5332), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n5373) );
  AOI22_X1 U6543 ( .A1(n3365), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5372) );
  NAND4_X1 U6544 ( .A1(n5375), .A2(n5374), .A3(n5373), .A4(n5372), .ZN(n5381)
         );
  AOI22_X1 U6545 ( .A1(n5478), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5379) );
  AOI22_X1 U6546 ( .A1(n5333), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5460), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5378) );
  AOI22_X1 U6547 ( .A1(n3525), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5377) );
  AOI22_X1 U6548 ( .A1(n5338), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5376) );
  NAND4_X1 U6549 ( .A1(n5379), .A2(n5378), .A3(n5377), .A4(n5376), .ZN(n5380)
         );
  NOR2_X1 U6550 ( .A1(n5381), .A2(n5380), .ZN(n5393) );
  NAND2_X1 U6551 ( .A1(n5383), .A2(n5382), .ZN(n5392) );
  XOR2_X1 U6552 ( .A(n5393), .B(n5392), .Z(n5386) );
  NAND2_X1 U6553 ( .A1(n5501), .A2(EAX_REG_25__SCAN_IN), .ZN(n5384) );
  OAI211_X1 U6554 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6111), .A(n5384), .B(
        n5499), .ZN(n5385) );
  AOI21_X1 U6555 ( .B1(n5386), .B2(n5467), .A(n5385), .ZN(n5387) );
  INV_X1 U6556 ( .A(n5387), .ZN(n5391) );
  AND2_X1 U6557 ( .A1(n5388), .A2(n6111), .ZN(n5389) );
  NOR2_X1 U6558 ( .A1(n5409), .A2(n5389), .ZN(n6113) );
  NAND2_X1 U6559 ( .A1(n6113), .A2(n5506), .ZN(n5390) );
  NAND2_X1 U6560 ( .A1(n5391), .A2(n5390), .ZN(n5964) );
  NOR2_X1 U6561 ( .A1(n5393), .A2(n5392), .ZN(n5415) );
  AOI22_X1 U6562 ( .A1(n5485), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5397) );
  AOI22_X1 U6563 ( .A1(n5333), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5396) );
  AOI22_X1 U6564 ( .A1(n3365), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5395) );
  AOI22_X1 U6565 ( .A1(n3488), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n5394) );
  NAND4_X1 U6566 ( .A1(n5397), .A2(n5396), .A3(n5395), .A4(n5394), .ZN(n5404)
         );
  AOI22_X1 U6567 ( .A1(n3525), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5402) );
  AOI22_X1 U6568 ( .A1(n5398), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5401) );
  AOI22_X1 U6569 ( .A1(n5438), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5400) );
  AOI22_X1 U6570 ( .A1(n5338), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5399) );
  NAND4_X1 U6571 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n5403)
         );
  OR2_X1 U6572 ( .A1(n5404), .A2(n5403), .ZN(n5414) );
  INV_X1 U6573 ( .A(n5414), .ZN(n5405) );
  XNOR2_X1 U6574 ( .A(n5415), .B(n5405), .ZN(n5406) );
  NAND2_X1 U6575 ( .A1(n5406), .A2(n5467), .ZN(n5413) );
  NAND2_X1 U6576 ( .A1(n6930), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5407)
         );
  NAND2_X1 U6577 ( .A1(n5499), .A2(n5407), .ZN(n5408) );
  AOI21_X1 U6578 ( .B1(n5501), .B2(EAX_REG_26__SCAN_IN), .A(n5408), .ZN(n5412)
         );
  NOR2_X1 U6579 ( .A1(n5409), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5410)
         );
  OR2_X1 U6580 ( .A1(n5428), .A2(n5410), .ZN(n6315) );
  NOR2_X1 U6581 ( .A1(n6315), .A2(n5499), .ZN(n5411) );
  AOI21_X1 U6582 ( .B1(n5413), .B2(n5412), .A(n5411), .ZN(n6045) );
  AND2_X2 U6583 ( .A1(n6044), .A2(n6045), .ZN(n5950) );
  NAND2_X1 U6584 ( .A1(n5415), .A2(n5414), .ZN(n5432) );
  AOI22_X1 U6585 ( .A1(n3488), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n5419) );
  AOI22_X1 U6586 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5460), .B1(n5475), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n5418) );
  AOI22_X1 U6587 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n5486), .B1(n3400), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5417) );
  AOI22_X1 U6588 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n5338), .B1(n5487), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5416) );
  NAND4_X1 U6589 ( .A1(n5419), .A2(n5418), .A3(n5417), .A4(n5416), .ZN(n5425)
         );
  AOI22_X1 U6590 ( .A1(n5333), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5423) );
  AOI22_X1 U6591 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n5480), .B1(n3525), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5422) );
  AOI22_X1 U6592 ( .A1(n5478), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5421) );
  AOI22_X1 U6593 ( .A1(n5307), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5420) );
  NAND4_X1 U6594 ( .A1(n5423), .A2(n5422), .A3(n5421), .A4(n5420), .ZN(n5424)
         );
  NOR2_X1 U6595 ( .A1(n5425), .A2(n5424), .ZN(n5433) );
  XOR2_X1 U6596 ( .A(n5432), .B(n5433), .Z(n5426) );
  NAND2_X1 U6597 ( .A1(n5426), .A2(n5467), .ZN(n5431) );
  INV_X1 U6598 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6101) );
  OAI21_X1 U6599 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6101), .A(n5499), .ZN(
        n5427) );
  AOI21_X1 U6600 ( .B1(n5501), .B2(EAX_REG_27__SCAN_IN), .A(n5427), .ZN(n5430)
         );
  XNOR2_X1 U6601 ( .A(n5428), .B(n6101), .ZN(n6105) );
  AND2_X1 U6602 ( .A1(n6105), .A2(n5506), .ZN(n5429) );
  AOI21_X1 U6603 ( .B1(n5431), .B2(n5430), .A(n5429), .ZN(n5953) );
  AND2_X2 U6604 ( .A1(n5950), .A2(n5953), .ZN(n5951) );
  NOR2_X1 U6605 ( .A1(n5433), .A2(n5432), .ZN(n5455) );
  AOI22_X1 U6606 ( .A1(n5485), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5478), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5437) );
  AOI22_X1 U6607 ( .A1(n5333), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5436) );
  AOI22_X1 U6608 ( .A1(n3365), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5435) );
  AOI22_X1 U6609 ( .A1(n3488), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5434) );
  NAND4_X1 U6610 ( .A1(n5437), .A2(n5436), .A3(n5435), .A4(n5434), .ZN(n5444)
         );
  AOI22_X1 U6611 ( .A1(n3525), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5442) );
  AOI22_X1 U6612 ( .A1(n5486), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5441) );
  AOI22_X1 U6613 ( .A1(n5438), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5440) );
  AOI22_X1 U6614 ( .A1(n5338), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5439) );
  NAND4_X1 U6615 ( .A1(n5442), .A2(n5441), .A3(n5440), .A4(n5439), .ZN(n5443)
         );
  OR2_X1 U6616 ( .A1(n5444), .A2(n5443), .ZN(n5454) );
  INV_X1 U6617 ( .A(n5454), .ZN(n5445) );
  XNOR2_X1 U6618 ( .A(n5455), .B(n5445), .ZN(n5446) );
  NAND2_X1 U6619 ( .A1(n5446), .A2(n5467), .ZN(n5453) );
  NAND2_X1 U6620 ( .A1(n6930), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5447)
         );
  NAND2_X1 U6621 ( .A1(n5499), .A2(n5447), .ZN(n5448) );
  AOI21_X1 U6622 ( .B1(n5501), .B2(EAX_REG_28__SCAN_IN), .A(n5448), .ZN(n5452)
         );
  OR2_X1 U6623 ( .A1(n5449), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5450)
         );
  NAND2_X1 U6624 ( .A1(n5472), .A2(n5450), .ZN(n6095) );
  NOR2_X1 U6625 ( .A1(n6095), .A2(n5499), .ZN(n5451) );
  AOI21_X1 U6626 ( .B1(n5453), .B2(n5452), .A(n5451), .ZN(n5940) );
  NAND2_X1 U6627 ( .A1(n5455), .A2(n5454), .ZN(n5494) );
  AOI22_X1 U6628 ( .A1(n5478), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5459) );
  AOI22_X1 U6629 ( .A1(n3488), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5458) );
  AOI22_X1 U6630 ( .A1(n5338), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5457) );
  AOI22_X1 U6631 ( .A1(n5307), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5456) );
  NAND4_X1 U6632 ( .A1(n5459), .A2(n5458), .A3(n5457), .A4(n5456), .ZN(n5466)
         );
  AOI22_X1 U6633 ( .A1(n5485), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5476), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5464) );
  AOI22_X1 U6634 ( .A1(n5333), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5460), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5463) );
  AOI22_X1 U6635 ( .A1(n3525), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5480), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5462) );
  AOI22_X1 U6636 ( .A1(n5486), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5461) );
  NAND4_X1 U6637 ( .A1(n5464), .A2(n5463), .A3(n5462), .A4(n5461), .ZN(n5465)
         );
  NOR2_X1 U6638 ( .A1(n5466), .A2(n5465), .ZN(n5495) );
  XOR2_X1 U6639 ( .A(n5494), .B(n5495), .Z(n5468) );
  NAND2_X1 U6640 ( .A1(n5468), .A2(n5467), .ZN(n5471) );
  OAI21_X1 U6641 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6084), .A(n5499), .ZN(
        n5469) );
  AOI21_X1 U6642 ( .B1(n5501), .B2(EAX_REG_29__SCAN_IN), .A(n5469), .ZN(n5470)
         );
  NAND2_X1 U6643 ( .A1(n5471), .A2(n5470), .ZN(n5474) );
  XNOR2_X1 U6644 ( .A(n5472), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6087)
         );
  NAND2_X1 U6645 ( .A1(n6087), .A2(n5506), .ZN(n5473) );
  NAND2_X1 U6646 ( .A1(n5474), .A2(n5473), .ZN(n5932) );
  OR2_X2 U6647 ( .A1(n5939), .A2(n5932), .ZN(n6030) );
  AOI22_X1 U6648 ( .A1(n5476), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5475), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5484) );
  AOI22_X1 U6649 ( .A1(n3525), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5483) );
  AOI22_X1 U6650 ( .A1(n5478), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5477), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5482) );
  AOI22_X1 U6651 ( .A1(n5480), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5479), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5481) );
  NAND4_X1 U6652 ( .A1(n5484), .A2(n5483), .A3(n5482), .A4(n5481), .ZN(n5493)
         );
  AOI22_X1 U6653 ( .A1(n3488), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5485), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n5491) );
  AOI22_X1 U6654 ( .A1(n5307), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5333), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5490) );
  AOI22_X1 U6655 ( .A1(n5486), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5438), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5489) );
  AOI22_X1 U6656 ( .A1(n5338), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5487), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5488) );
  NAND4_X1 U6657 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n5492)
         );
  NOR2_X1 U6658 ( .A1(n5493), .A2(n5492), .ZN(n5497) );
  NOR2_X1 U6659 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  XOR2_X1 U6660 ( .A(n5497), .B(n5496), .Z(n5504) );
  NAND2_X1 U6661 ( .A1(n6930), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5498)
         );
  NAND2_X1 U6662 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  AOI21_X1 U6663 ( .B1(n5501), .B2(EAX_REG_30__SCAN_IN), .A(n5500), .ZN(n5502)
         );
  OAI21_X1 U6664 ( .B1(n5504), .B2(n5503), .A(n5502), .ZN(n5508) );
  XNOR2_X1 U6665 ( .A(n5505), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6302)
         );
  NAND2_X1 U6666 ( .A1(n6302), .A2(n5506), .ZN(n5507) );
  NAND2_X1 U6667 ( .A1(n5508), .A2(n5507), .ZN(n6031) );
  NOR2_X2 U6668 ( .A1(n6030), .A2(n6031), .ZN(n6029) );
  AOI22_X1 U6669 ( .A1(n5510), .A2(EAX_REG_31__SCAN_IN), .B1(n5509), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5511) );
  XNOR2_X1 U6670 ( .A(n6029), .B(n5511), .ZN(n6065) );
  NAND2_X1 U6671 ( .A1(n6803), .A2(REIP_REG_31__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U6672 ( .A1(n6694), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5512)
         );
  OAI211_X1 U6673 ( .C1(n6704), .C2(n5513), .A(n5517), .B(n5512), .ZN(n5514)
         );
  AOI21_X1 U6674 ( .B1(n6065), .B2(n6698), .A(n5514), .ZN(n5515) );
  OAI21_X1 U6675 ( .B1(n3202), .B2(n6681), .A(n5515), .ZN(U2955) );
  OAI21_X1 U6676 ( .B1(n6383), .B2(n5518), .A(n5516), .ZN(n5522) );
  INV_X1 U6677 ( .A(n5517), .ZN(n5521) );
  INV_X1 U6678 ( .A(n5518), .ZN(n5519) );
  NOR3_X1 U6679 ( .A1(n5540), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5519), 
        .ZN(n5520) );
  AOI211_X1 U6680 ( .C1(n5522), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5521), .B(n5520), .ZN(n5530) );
  AND2_X1 U6681 ( .A1(n5526), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5523)
         );
  AOI21_X1 U6682 ( .B1(n3852), .B2(EBX_REG_30__SCAN_IN), .A(n5523), .ZN(n5534)
         );
  AOI21_X1 U6683 ( .B1(n5534), .B2(n5525), .A(n5533), .ZN(n5528) );
  AOI22_X1 U6684 ( .A1(n3852), .A2(EBX_REG_31__SCAN_IN), .B1(n5526), .B2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5527) );
  XNOR2_X1 U6685 ( .A(n5528), .B(n5527), .ZN(n6026) );
  NAND2_X1 U6686 ( .A1(n6026), .A2(n6799), .ZN(n5529) );
  OAI211_X1 U6687 ( .C1(n3202), .C2(n6773), .A(n5530), .B(n5529), .ZN(U2987)
         );
  INV_X1 U6688 ( .A(n5534), .ZN(n5536) );
  AOI211_X1 U6689 ( .C1(n5537), .C2(n5945), .A(n5536), .B(n5535), .ZN(n5538)
         );
  INV_X1 U6690 ( .A(REIP_REG_30__SCAN_IN), .ZN(n7128) );
  NOR2_X1 U6691 ( .A1(n6774), .A2(n7128), .ZN(n6079) );
  NOR3_X1 U6692 ( .A1(n5540), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5539), 
        .ZN(n5541) );
  INV_X1 U6693 ( .A(n6214), .ZN(n5543) );
  OAI211_X1 U6694 ( .C1(n6750), .C2(n5543), .A(n5542), .B(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5544) );
  OAI211_X1 U6695 ( .C1(n6082), .C2(n6773), .A(n5545), .B(n5544), .ZN(U2988)
         );
  INV_X1 U6696 ( .A(n5546), .ZN(n6213) );
  NAND2_X1 U6697 ( .A1(n6264), .A2(n6213), .ZN(n5547) );
  NAND2_X1 U6698 ( .A1(n5547), .A2(n6262), .ZN(n5548) );
  NAND2_X1 U6699 ( .A1(n5548), .A2(n6165), .ZN(n5549) );
  XNOR2_X1 U6700 ( .A(n6262), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6138)
         );
  NOR3_X1 U6701 ( .A1(n6147), .A2(n6131), .A3(n5553), .ZN(n6120) );
  NAND2_X1 U6702 ( .A1(n5986), .A2(n5559), .ZN(n5560) );
  NAND2_X1 U6703 ( .A1(n5963), .A2(n5560), .ZN(n6340) );
  NOR2_X1 U6704 ( .A1(n6340), .A2(n6679), .ZN(n5563) );
  NAND2_X1 U6705 ( .A1(n6803), .A2(REIP_REG_24__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U6706 ( .A1(n6694), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5561)
         );
  OAI211_X1 U6707 ( .C1(n6704), .C2(n5978), .A(n6217), .B(n5561), .ZN(n5562)
         );
  AOI22_X1 U6708 ( .A1(EBX_REG_24__SCAN_IN), .A2(keyinput166), .B1(
        INSTQUEUE_REG_2__1__SCAN_IN), .B2(keyinput222), .ZN(n5564) );
  OAI221_X1 U6709 ( .B1(EBX_REG_24__SCAN_IN), .B2(keyinput166), .C1(
        INSTQUEUE_REG_2__1__SCAN_IN), .C2(keyinput222), .A(n5564), .ZN(n5571)
         );
  AOI22_X1 U6710 ( .A1(DATAI_23_), .A2(keyinput224), .B1(
        INSTQUEUE_REG_4__2__SCAN_IN), .B2(keyinput135), .ZN(n5565) );
  OAI221_X1 U6711 ( .B1(DATAI_23_), .B2(keyinput224), .C1(
        INSTQUEUE_REG_4__2__SCAN_IN), .C2(keyinput135), .A(n5565), .ZN(n5570)
         );
  AOI22_X1 U6712 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(keyinput242), .B1(
        INSTQUEUE_REG_5__4__SCAN_IN), .B2(keyinput216), .ZN(n5566) );
  OAI221_X1 U6713 ( .B1(DATAWIDTH_REG_27__SCAN_IN), .B2(keyinput242), .C1(
        INSTQUEUE_REG_5__4__SCAN_IN), .C2(keyinput216), .A(n5566), .ZN(n5569)
         );
  AOI22_X1 U6714 ( .A1(UWORD_REG_1__SCAN_IN), .A2(keyinput189), .B1(
        INSTADDRPOINTER_REG_16__SCAN_IN), .B2(keyinput195), .ZN(n5567) );
  OAI221_X1 U6715 ( .B1(UWORD_REG_1__SCAN_IN), .B2(keyinput189), .C1(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C2(keyinput195), .A(n5567), .ZN(
        n5568) );
  NOR4_X1 U6716 ( .A1(n5571), .A2(n5570), .A3(n5569), .A4(n5568), .ZN(n5599)
         );
  AOI22_X1 U6717 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(keyinput149), 
        .B1(INSTQUEUE_REG_4__1__SCAN_IN), .B2(keyinput156), .ZN(n5572) );
  OAI221_X1 U6718 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput149), 
        .C1(INSTQUEUE_REG_4__1__SCAN_IN), .C2(keyinput156), .A(n5572), .ZN(
        n5579) );
  AOI22_X1 U6719 ( .A1(DATAI_0_), .A2(keyinput133), .B1(
        INSTADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput191), .ZN(n5573) );
  OAI221_X1 U6720 ( .B1(DATAI_0_), .B2(keyinput133), .C1(
        INSTADDRPOINTER_REG_5__SCAN_IN), .C2(keyinput191), .A(n5573), .ZN(
        n5578) );
  AOI22_X1 U6721 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(keyinput150), .B1(
        EBX_REG_7__SCAN_IN), .B2(keyinput255), .ZN(n5574) );
  OAI221_X1 U6722 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput150), 
        .C1(EBX_REG_7__SCAN_IN), .C2(keyinput255), .A(n5574), .ZN(n5577) );
  AOI22_X1 U6723 ( .A1(REIP_REG_14__SCAN_IN), .A2(keyinput131), .B1(
        INSTADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput225), .ZN(n5575) );
  OAI221_X1 U6724 ( .B1(REIP_REG_14__SCAN_IN), .B2(keyinput131), .C1(
        INSTADDRPOINTER_REG_22__SCAN_IN), .C2(keyinput225), .A(n5575), .ZN(
        n5576) );
  NOR4_X1 U6725 ( .A1(n5579), .A2(n5578), .A3(n5577), .A4(n5576), .ZN(n5598)
         );
  AOI22_X1 U6726 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(keyinput192), .B1(n6301), .B2(keyinput212), .ZN(n5580) );
  OAI221_X1 U6727 ( .B1(DATAWIDTH_REG_29__SCAN_IN), .B2(keyinput192), .C1(
        n6301), .C2(keyinput212), .A(n5580), .ZN(n5587) );
  AOI22_X1 U6728 ( .A1(DATAI_30_), .A2(keyinput157), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput221), .ZN(n5581) );
  OAI221_X1 U6729 ( .B1(DATAI_30_), .B2(keyinput157), .C1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .C2(keyinput221), .A(n5581), .ZN(
        n5586) );
  AOI22_X1 U6730 ( .A1(ADDRESS_REG_9__SCAN_IN), .A2(keyinput144), .B1(
        UWORD_REG_0__SCAN_IN), .B2(keyinput139), .ZN(n5582) );
  OAI221_X1 U6731 ( .B1(ADDRESS_REG_9__SCAN_IN), .B2(keyinput144), .C1(
        UWORD_REG_0__SCAN_IN), .C2(keyinput139), .A(n5582), .ZN(n5585) );
  AOI22_X1 U6732 ( .A1(DATAI_2_), .A2(keyinput240), .B1(DATAI_27_), .B2(
        keyinput138), .ZN(n5583) );
  OAI221_X1 U6733 ( .B1(DATAI_2_), .B2(keyinput240), .C1(DATAI_27_), .C2(
        keyinput138), .A(n5583), .ZN(n5584) );
  NOR4_X1 U6734 ( .A1(n5587), .A2(n5586), .A3(n5585), .A4(n5584), .ZN(n5597)
         );
  AOI22_X1 U6735 ( .A1(UWORD_REG_9__SCAN_IN), .A2(keyinput129), .B1(DATAI_8_), 
        .B2(keyinput244), .ZN(n5588) );
  OAI221_X1 U6736 ( .B1(UWORD_REG_9__SCAN_IN), .B2(keyinput129), .C1(DATAI_8_), 
        .C2(keyinput244), .A(n5588), .ZN(n5595) );
  AOI22_X1 U6737 ( .A1(DATAO_REG_2__SCAN_IN), .A2(keyinput213), .B1(
        INSTQUEUE_REG_1__4__SCAN_IN), .B2(keyinput145), .ZN(n5589) );
  OAI221_X1 U6738 ( .B1(DATAO_REG_2__SCAN_IN), .B2(keyinput213), .C1(
        INSTQUEUE_REG_1__4__SCAN_IN), .C2(keyinput145), .A(n5589), .ZN(n5594)
         );
  AOI22_X1 U6739 ( .A1(EBX_REG_21__SCAN_IN), .A2(keyinput210), .B1(
        INSTQUEUE_REG_4__5__SCAN_IN), .B2(keyinput163), .ZN(n5590) );
  OAI221_X1 U6740 ( .B1(EBX_REG_21__SCAN_IN), .B2(keyinput210), .C1(
        INSTQUEUE_REG_4__5__SCAN_IN), .C2(keyinput163), .A(n5590), .ZN(n5593)
         );
  AOI22_X1 U6741 ( .A1(EAX_REG_10__SCAN_IN), .A2(keyinput248), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput187), .ZN(n5591) );
  OAI221_X1 U6742 ( .B1(EAX_REG_10__SCAN_IN), .B2(keyinput248), .C1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(keyinput187), .A(n5591), .ZN(
        n5592) );
  NOR4_X1 U6743 ( .A1(n5595), .A2(n5594), .A3(n5593), .A4(n5592), .ZN(n5596)
         );
  NAND4_X1 U6744 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n5722)
         );
  AOI22_X1 U6745 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput153), .B1(
        INSTQUEUE_REG_2__4__SCAN_IN), .B2(keyinput215), .ZN(n5600) );
  OAI221_X1 U6746 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput153), .C1(
        INSTQUEUE_REG_2__4__SCAN_IN), .C2(keyinput215), .A(n5600), .ZN(n5607)
         );
  AOI22_X1 U6747 ( .A1(DATAI_13_), .A2(keyinput176), .B1(EBX_REG_27__SCAN_IN), 
        .B2(keyinput188), .ZN(n5601) );
  OAI221_X1 U6748 ( .B1(DATAI_13_), .B2(keyinput176), .C1(EBX_REG_27__SCAN_IN), 
        .C2(keyinput188), .A(n5601), .ZN(n5606) );
  AOI22_X1 U6749 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(keyinput167), 
        .B1(INSTQUEUE_REG_5__0__SCAN_IN), .B2(keyinput245), .ZN(n5602) );
  OAI221_X1 U6750 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(keyinput167), 
        .C1(INSTQUEUE_REG_5__0__SCAN_IN), .C2(keyinput245), .A(n5602), .ZN(
        n5605) );
  AOI22_X1 U6751 ( .A1(ADDRESS_REG_13__SCAN_IN), .A2(keyinput207), .B1(
        INSTQUEUE_REG_8__5__SCAN_IN), .B2(keyinput134), .ZN(n5603) );
  OAI221_X1 U6752 ( .B1(ADDRESS_REG_13__SCAN_IN), .B2(keyinput207), .C1(
        INSTQUEUE_REG_8__5__SCAN_IN), .C2(keyinput134), .A(n5603), .ZN(n5604)
         );
  NOR4_X1 U6753 ( .A1(n5607), .A2(n5606), .A3(n5605), .A4(n5604), .ZN(n5635)
         );
  AOI22_X1 U6754 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(keyinput209), .B1(
        INSTQUEUE_REG_9__1__SCAN_IN), .B2(keyinput130), .ZN(n5608) );
  OAI221_X1 U6755 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput209), 
        .C1(INSTQUEUE_REG_9__1__SCAN_IN), .C2(keyinput130), .A(n5608), .ZN(
        n5615) );
  AOI22_X1 U6756 ( .A1(EAX_REG_18__SCAN_IN), .A2(keyinput233), .B1(
        STATE2_REG_2__SCAN_IN), .B2(keyinput185), .ZN(n5609) );
  OAI221_X1 U6757 ( .B1(EAX_REG_18__SCAN_IN), .B2(keyinput233), .C1(
        STATE2_REG_2__SCAN_IN), .C2(keyinput185), .A(n5609), .ZN(n5614) );
  AOI22_X1 U6758 ( .A1(ADDRESS_REG_28__SCAN_IN), .A2(keyinput232), .B1(
        INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput249), .ZN(n5610) );
  OAI221_X1 U6759 ( .B1(ADDRESS_REG_28__SCAN_IN), .B2(keyinput232), .C1(
        INSTADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput249), .A(n5610), .ZN(
        n5613) );
  AOI22_X1 U6760 ( .A1(ADS_N_REG_SCAN_IN), .A2(keyinput141), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput140), .ZN(n5611) );
  OAI221_X1 U6761 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput141), .C1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .C2(keyinput140), .A(n5611), .ZN(
        n5612) );
  NOR4_X1 U6762 ( .A1(n5615), .A2(n5614), .A3(n5613), .A4(n5612), .ZN(n5634)
         );
  AOI22_X1 U6763 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(keyinput206), .B1(
        INSTQUEUE_REG_0__4__SCAN_IN), .B2(keyinput247), .ZN(n5616) );
  OAI221_X1 U6764 ( .B1(INSTQUEUE_REG_6__6__SCAN_IN), .B2(keyinput206), .C1(
        INSTQUEUE_REG_0__4__SCAN_IN), .C2(keyinput247), .A(n5616), .ZN(n5623)
         );
  AOI22_X1 U6765 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(keyinput170), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput154), .ZN(n5617) );
  OAI221_X1 U6766 ( .B1(DATAWIDTH_REG_28__SCAN_IN), .B2(keyinput170), .C1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .C2(keyinput154), .A(n5617), .ZN(n5622) );
  AOI22_X1 U6767 ( .A1(DATAO_REG_14__SCAN_IN), .A2(keyinput128), .B1(
        EBX_REG_26__SCAN_IN), .B2(keyinput142), .ZN(n5618) );
  OAI221_X1 U6768 ( .B1(DATAO_REG_14__SCAN_IN), .B2(keyinput128), .C1(
        EBX_REG_26__SCAN_IN), .C2(keyinput142), .A(n5618), .ZN(n5621) );
  AOI22_X1 U6769 ( .A1(UWORD_REG_4__SCAN_IN), .A2(keyinput203), .B1(
        INSTQUEUE_REG_11__2__SCAN_IN), .B2(keyinput204), .ZN(n5619) );
  OAI221_X1 U6770 ( .B1(UWORD_REG_4__SCAN_IN), .B2(keyinput203), .C1(
        INSTQUEUE_REG_11__2__SCAN_IN), .C2(keyinput204), .A(n5619), .ZN(n5620)
         );
  NOR4_X1 U6771 ( .A1(n5623), .A2(n5622), .A3(n5621), .A4(n5620), .ZN(n5633)
         );
  AOI22_X1 U6772 ( .A1(HOLD), .A2(keyinput186), .B1(
        INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput196), .ZN(n5624) );
  OAI221_X1 U6773 ( .B1(HOLD), .B2(keyinput186), .C1(
        INSTQUEUE_REG_14__4__SCAN_IN), .C2(keyinput196), .A(n5624), .ZN(n5631)
         );
  AOI22_X1 U6774 ( .A1(DATAO_REG_31__SCAN_IN), .A2(keyinput246), .B1(
        EAX_REG_21__SCAN_IN), .B2(keyinput169), .ZN(n5625) );
  OAI221_X1 U6775 ( .B1(DATAO_REG_31__SCAN_IN), .B2(keyinput246), .C1(
        EAX_REG_21__SCAN_IN), .C2(keyinput169), .A(n5625), .ZN(n5630) );
  AOI22_X1 U6776 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(keyinput218), 
        .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(keyinput241), .ZN(n5626) );
  OAI221_X1 U6777 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(keyinput218), 
        .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(keyinput241), .A(n5626), 
        .ZN(n5629) );
  AOI22_X1 U6778 ( .A1(EBX_REG_2__SCAN_IN), .A2(keyinput243), .B1(
        INSTQUEUE_REG_15__1__SCAN_IN), .B2(keyinput250), .ZN(n5627) );
  OAI221_X1 U6779 ( .B1(EBX_REG_2__SCAN_IN), .B2(keyinput243), .C1(
        INSTQUEUE_REG_15__1__SCAN_IN), .C2(keyinput250), .A(n5627), .ZN(n5628)
         );
  NOR4_X1 U6780 ( .A1(n5631), .A2(n5630), .A3(n5629), .A4(n5628), .ZN(n5632)
         );
  NAND4_X1 U6781 ( .A1(n5635), .A2(n5634), .A3(n5633), .A4(n5632), .ZN(n5721)
         );
  AOI22_X1 U6782 ( .A1(EAX_REG_28__SCAN_IN), .A2(keyinput205), .B1(
        PHYADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput239), .ZN(n5636) );
  OAI221_X1 U6783 ( .B1(EAX_REG_28__SCAN_IN), .B2(keyinput205), .C1(
        PHYADDRPOINTER_REG_15__SCAN_IN), .C2(keyinput239), .A(n5636), .ZN(
        n5644) );
  AOI22_X1 U6784 ( .A1(EBX_REG_4__SCAN_IN), .A2(keyinput147), .B1(
        INSTQUEUE_REG_6__3__SCAN_IN), .B2(keyinput177), .ZN(n5637) );
  OAI221_X1 U6785 ( .B1(EBX_REG_4__SCAN_IN), .B2(keyinput147), .C1(
        INSTQUEUE_REG_6__3__SCAN_IN), .C2(keyinput177), .A(n5637), .ZN(n5643)
         );
  INV_X1 U6786 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7116) );
  AOI22_X1 U6787 ( .A1(keyinput220), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n7116), .B2(keyinput183), .ZN(n5638) );
  OAI221_X1 U6788 ( .B1(keyinput220), .B2(INSTQUEUE_REG_4__0__SCAN_IN), .C1(
        n7116), .C2(keyinput183), .A(n5638), .ZN(n5642) );
  INV_X1 U6789 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5640) );
  AOI22_X1 U6790 ( .A1(n6597), .A2(keyinput152), .B1(n5640), .B2(keyinput236), 
        .ZN(n5639) );
  OAI221_X1 U6791 ( .B1(n6597), .B2(keyinput152), .C1(n5640), .C2(keyinput236), 
        .A(n5639), .ZN(n5641) );
  NOR4_X1 U6792 ( .A1(n5644), .A2(n5643), .A3(n5642), .A4(n5641), .ZN(n5675)
         );
  INV_X1 U6793 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5881) );
  INV_X1 U6794 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n7156) );
  AOI22_X1 U6795 ( .A1(n5881), .A2(keyinput136), .B1(keyinput237), .B2(n7156), 
        .ZN(n5645) );
  OAI221_X1 U6796 ( .B1(n5881), .B2(keyinput136), .C1(n7156), .C2(keyinput237), 
        .A(n5645), .ZN(n5652) );
  INV_X1 U6797 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5763) );
  AOI22_X1 U6798 ( .A1(n4855), .A2(keyinput174), .B1(keyinput197), .B2(n5763), 
        .ZN(n5646) );
  OAI221_X1 U6799 ( .B1(n4855), .B2(keyinput174), .C1(n5763), .C2(keyinput197), 
        .A(n5646), .ZN(n5651) );
  INV_X1 U6800 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n6567) );
  INV_X1 U6801 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n5854) );
  AOI22_X1 U6802 ( .A1(n6567), .A2(keyinput132), .B1(keyinput168), .B2(n5854), 
        .ZN(n5647) );
  OAI221_X1 U6803 ( .B1(n6567), .B2(keyinput132), .C1(n5854), .C2(keyinput168), 
        .A(n5647), .ZN(n5650) );
  INV_X1 U6804 ( .A(DATAI_14_), .ZN(n6655) );
  INV_X1 U6805 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n5827) );
  AOI22_X1 U6806 ( .A1(n6655), .A2(keyinput175), .B1(keyinput200), .B2(n5827), 
        .ZN(n5648) );
  OAI221_X1 U6807 ( .B1(n6655), .B2(keyinput175), .C1(n5827), .C2(keyinput200), 
        .A(n5648), .ZN(n5649) );
  NOR4_X1 U6808 ( .A1(n5652), .A2(n5651), .A3(n5650), .A4(n5649), .ZN(n5674)
         );
  INV_X1 U6809 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n7096) );
  AOI22_X1 U6810 ( .A1(n7096), .A2(keyinput253), .B1(n5853), .B2(keyinput178), 
        .ZN(n5653) );
  OAI221_X1 U6811 ( .B1(n7096), .B2(keyinput253), .C1(n5853), .C2(keyinput178), 
        .A(n5653), .ZN(n5661) );
  INV_X1 U6812 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5843) );
  INV_X1 U6813 ( .A(NA_N), .ZN(n7066) );
  AOI22_X1 U6814 ( .A1(n5843), .A2(keyinput171), .B1(keyinput182), .B2(n7066), 
        .ZN(n5654) );
  OAI221_X1 U6815 ( .B1(n5843), .B2(keyinput171), .C1(n7066), .C2(keyinput182), 
        .A(n5654), .ZN(n5660) );
  INV_X1 U6816 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n6834) );
  AOI22_X1 U6817 ( .A1(n6035), .A2(keyinput226), .B1(n6834), .B2(keyinput194), 
        .ZN(n5655) );
  OAI221_X1 U6818 ( .B1(n6035), .B2(keyinput226), .C1(n6834), .C2(keyinput194), 
        .A(n5655), .ZN(n5659) );
  INV_X1 U6819 ( .A(DATAI_19_), .ZN(n5657) );
  INV_X1 U6820 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7124) );
  AOI22_X1 U6821 ( .A1(n5657), .A2(keyinput160), .B1(keyinput161), .B2(n7124), 
        .ZN(n5656) );
  OAI221_X1 U6822 ( .B1(n5657), .B2(keyinput160), .C1(n7124), .C2(keyinput161), 
        .A(n5656), .ZN(n5658) );
  NOR4_X1 U6823 ( .A1(n5661), .A2(n5660), .A3(n5659), .A4(n5658), .ZN(n5673)
         );
  INV_X1 U6824 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7118) );
  INV_X1 U6825 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n5897) );
  AOI22_X1 U6826 ( .A1(n7118), .A2(keyinput164), .B1(keyinput173), .B2(n5897), 
        .ZN(n5662) );
  OAI221_X1 U6827 ( .B1(n7118), .B2(keyinput164), .C1(n5897), .C2(keyinput173), 
        .A(n5662), .ZN(n5671) );
  INV_X1 U6828 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6374) );
  INV_X1 U6829 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7108) );
  AOI22_X1 U6830 ( .A1(n6374), .A2(keyinput219), .B1(keyinput143), .B2(n7108), 
        .ZN(n5663) );
  OAI221_X1 U6831 ( .B1(n6374), .B2(keyinput219), .C1(n7108), .C2(keyinput143), 
        .A(n5663), .ZN(n5670) );
  INV_X1 U6832 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n5834) );
  AOI22_X1 U6833 ( .A1(n5665), .A2(keyinput254), .B1(keyinput208), .B2(n5834), 
        .ZN(n5664) );
  OAI221_X1 U6834 ( .B1(n5665), .B2(keyinput254), .C1(n5834), .C2(keyinput208), 
        .A(n5664), .ZN(n5669) );
  INV_X1 U6835 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5667) );
  INV_X1 U6836 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5869) );
  AOI22_X1 U6837 ( .A1(n5667), .A2(keyinput162), .B1(keyinput227), .B2(n5869), 
        .ZN(n5666) );
  OAI221_X1 U6838 ( .B1(n5667), .B2(keyinput162), .C1(n5869), .C2(keyinput227), 
        .A(n5666), .ZN(n5668) );
  NOR4_X1 U6839 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(n5672)
         );
  NAND4_X1 U6840 ( .A1(n5675), .A2(n5674), .A3(n5673), .A4(n5672), .ZN(n5720)
         );
  AOI22_X1 U6841 ( .A1(n5678), .A2(keyinput155), .B1(keyinput180), .B2(n5677), 
        .ZN(n5676) );
  OAI221_X1 U6842 ( .B1(n5678), .B2(keyinput155), .C1(n5677), .C2(keyinput180), 
        .A(n5676), .ZN(n5686) );
  INV_X1 U6843 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7050) );
  INV_X1 U6844 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6415) );
  AOI22_X1 U6845 ( .A1(n7050), .A2(keyinput229), .B1(keyinput238), .B2(n6415), 
        .ZN(n5679) );
  OAI221_X1 U6846 ( .B1(n7050), .B2(keyinput229), .C1(n6415), .C2(keyinput238), 
        .A(n5679), .ZN(n5685) );
  INV_X1 U6847 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6828) );
  AOI22_X1 U6848 ( .A1(n5681), .A2(keyinput137), .B1(n6828), .B2(keyinput228), 
        .ZN(n5680) );
  OAI221_X1 U6849 ( .B1(n5681), .B2(keyinput137), .C1(n6828), .C2(keyinput228), 
        .A(n5680), .ZN(n5684) );
  INV_X1 U6850 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n5883) );
  INV_X1 U6851 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n7048) );
  AOI22_X1 U6852 ( .A1(n5883), .A2(keyinput193), .B1(keyinput223), .B2(n7048), 
        .ZN(n5682) );
  OAI221_X1 U6853 ( .B1(n5883), .B2(keyinput193), .C1(n7048), .C2(keyinput223), 
        .A(n5682), .ZN(n5683) );
  NOR4_X1 U6854 ( .A1(n5686), .A2(n5685), .A3(n5684), .A4(n5683), .ZN(n5718)
         );
  INV_X1 U6855 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5688) );
  INV_X1 U6856 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n7117) );
  AOI22_X1 U6857 ( .A1(n5688), .A2(keyinput198), .B1(keyinput230), .B2(n7117), 
        .ZN(n5687) );
  OAI221_X1 U6858 ( .B1(n5688), .B2(keyinput198), .C1(n7117), .C2(keyinput230), 
        .A(n5687), .ZN(n5696) );
  INV_X1 U6859 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7134) );
  INV_X1 U6860 ( .A(DATAI_22_), .ZN(n5757) );
  AOI22_X1 U6861 ( .A1(n7134), .A2(keyinput151), .B1(keyinput201), .B2(n5757), 
        .ZN(n5689) );
  OAI221_X1 U6862 ( .B1(n7134), .B2(keyinput151), .C1(n5757), .C2(keyinput201), 
        .A(n5689), .ZN(n5695) );
  INV_X1 U6863 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n7052) );
  AOI22_X1 U6864 ( .A1(n7052), .A2(keyinput235), .B1(n5818), .B2(keyinput214), 
        .ZN(n5690) );
  OAI221_X1 U6865 ( .B1(n7052), .B2(keyinput235), .C1(n5818), .C2(keyinput214), 
        .A(n5690), .ZN(n5694) );
  INV_X1 U6866 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5692) );
  INV_X1 U6867 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7119) );
  AOI22_X1 U6868 ( .A1(n5692), .A2(keyinput148), .B1(keyinput181), .B2(n7119), 
        .ZN(n5691) );
  OAI221_X1 U6869 ( .B1(n5692), .B2(keyinput148), .C1(n7119), .C2(keyinput181), 
        .A(n5691), .ZN(n5693) );
  NOR4_X1 U6870 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5693), .ZN(n5717)
         );
  INV_X1 U6871 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n5733) );
  INV_X1 U6872 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7109) );
  AOI22_X1 U6873 ( .A1(n5733), .A2(keyinput179), .B1(keyinput172), .B2(n7109), 
        .ZN(n5697) );
  OAI221_X1 U6874 ( .B1(n5733), .B2(keyinput179), .C1(n7109), .C2(keyinput172), 
        .A(n5697), .ZN(n5706) );
  INV_X1 U6875 ( .A(REIP_REG_24__SCAN_IN), .ZN(n5976) );
  INV_X1 U6876 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5699) );
  AOI22_X1 U6877 ( .A1(n5976), .A2(keyinput217), .B1(n5699), .B2(keyinput158), 
        .ZN(n5698) );
  OAI221_X1 U6878 ( .B1(n5976), .B2(keyinput217), .C1(n5699), .C2(keyinput158), 
        .A(n5698), .ZN(n5705) );
  INV_X1 U6879 ( .A(DATAWIDTH_REG_26__SCAN_IN), .ZN(n7047) );
  AOI22_X1 U6880 ( .A1(n7047), .A2(keyinput146), .B1(n5841), .B2(keyinput234), 
        .ZN(n5700) );
  OAI221_X1 U6881 ( .B1(n7047), .B2(keyinput146), .C1(n5841), .C2(keyinput234), 
        .A(n5700), .ZN(n5704) );
  INV_X1 U6882 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5702) );
  INV_X1 U6883 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n5788) );
  AOI22_X1 U6884 ( .A1(n5702), .A2(keyinput199), .B1(keyinput190), .B2(n5788), 
        .ZN(n5701) );
  OAI221_X1 U6885 ( .B1(n5702), .B2(keyinput199), .C1(n5788), .C2(keyinput190), 
        .A(n5701), .ZN(n5703) );
  NOR4_X1 U6886 ( .A1(n5706), .A2(n5705), .A3(n5704), .A4(n5703), .ZN(n5716)
         );
  INV_X1 U6887 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n7049) );
  AOI22_X1 U6888 ( .A1(n6589), .A2(keyinput202), .B1(keyinput165), .B2(n7049), 
        .ZN(n5707) );
  OAI221_X1 U6889 ( .B1(n6589), .B2(keyinput202), .C1(n7049), .C2(keyinput165), 
        .A(n5707), .ZN(n5714) );
  AOI22_X1 U6890 ( .A1(n6624), .A2(keyinput211), .B1(n5977), .B2(keyinput231), 
        .ZN(n5708) );
  OAI221_X1 U6891 ( .B1(n6624), .B2(keyinput211), .C1(n5977), .C2(keyinput231), 
        .A(n5708), .ZN(n5713) );
  INV_X1 U6892 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6840) );
  AOI22_X1 U6893 ( .A1(n6840), .A2(keyinput251), .B1(keyinput159), .B2(n6441), 
        .ZN(n5709) );
  OAI221_X1 U6894 ( .B1(n6840), .B2(keyinput251), .C1(n6441), .C2(keyinput159), 
        .A(n5709), .ZN(n5712) );
  INV_X1 U6895 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n7051) );
  AOI22_X1 U6896 ( .A1(n7051), .A2(keyinput184), .B1(keyinput252), .B2(n7082), 
        .ZN(n5710) );
  OAI221_X1 U6897 ( .B1(n7051), .B2(keyinput184), .C1(n7082), .C2(keyinput252), 
        .A(n5710), .ZN(n5711) );
  NOR4_X1 U6898 ( .A1(n5714), .A2(n5713), .A3(n5712), .A4(n5711), .ZN(n5715)
         );
  NAND4_X1 U6899 ( .A1(n5718), .A2(n5717), .A3(n5716), .A4(n5715), .ZN(n5719)
         );
  NOR4_X1 U6900 ( .A1(n5722), .A2(n5721), .A3(n5720), .A4(n5719), .ZN(n5908)
         );
  OAI22_X1 U6901 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput15), .B1(keyinput83), 
        .B2(DATAI_1_), .ZN(n5723) );
  AOI221_X1 U6902 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput15), .C1(DATAI_1_), 
        .C2(keyinput83), .A(n5723), .ZN(n5730) );
  OAI22_X1 U6903 ( .A1(EAX_REG_10__SCAN_IN), .A2(keyinput120), .B1(
        DATAWIDTH_REG_28__SCAN_IN), .B2(keyinput42), .ZN(n5724) );
  AOI221_X1 U6904 ( .B1(EAX_REG_10__SCAN_IN), .B2(keyinput120), .C1(keyinput42), .C2(DATAWIDTH_REG_28__SCAN_IN), .A(n5724), .ZN(n5729) );
  OAI22_X1 U6905 ( .A1(EBX_REG_26__SCAN_IN), .A2(keyinput14), .B1(keyinput10), 
        .B2(DATAI_27_), .ZN(n5725) );
  AOI221_X1 U6906 ( .B1(EBX_REG_26__SCAN_IN), .B2(keyinput14), .C1(DATAI_27_), 
        .C2(keyinput10), .A(n5725), .ZN(n5728) );
  OAI22_X1 U6907 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(keyinput94), .B1(
        DATAWIDTH_REG_27__SCAN_IN), .B2(keyinput114), .ZN(n5726) );
  AOI221_X1 U6908 ( .B1(INSTQUEUE_REG_2__1__SCAN_IN), .B2(keyinput94), .C1(
        keyinput114), .C2(DATAWIDTH_REG_27__SCAN_IN), .A(n5726), .ZN(n5727) );
  NAND4_X1 U6909 ( .A1(n5730), .A2(n5729), .A3(n5728), .A4(n5727), .ZN(n5736)
         );
  AOI22_X1 U6910 ( .A1(n7119), .A2(keyinput53), .B1(keyinput124), .B2(n7082), 
        .ZN(n5731) );
  OAI221_X1 U6911 ( .B1(n7119), .B2(keyinput53), .C1(n7082), .C2(keyinput124), 
        .A(n5731), .ZN(n5735) );
  AOI22_X1 U6912 ( .A1(n7047), .A2(keyinput18), .B1(n5733), .B2(keyinput51), 
        .ZN(n5732) );
  OAI221_X1 U6913 ( .B1(n7047), .B2(keyinput18), .C1(n5733), .C2(keyinput51), 
        .A(n5732), .ZN(n5734) );
  OR3_X1 U6914 ( .A1(n5736), .A2(n5735), .A3(n5734), .ZN(n5755) );
  OAI22_X1 U6915 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(keyinput91), .B1(
        MEMORYFETCH_REG_SCAN_IN), .B2(keyinput52), .ZN(n5737) );
  AOI221_X1 U6916 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput91), 
        .C1(keyinput52), .C2(MEMORYFETCH_REG_SCAN_IN), .A(n5737), .ZN(n5744)
         );
  OAI22_X1 U6917 ( .A1(EBX_REG_10__SCAN_IN), .A2(keyinput27), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(keyinput44), .ZN(n5738) );
  AOI221_X1 U6918 ( .B1(EBX_REG_10__SCAN_IN), .B2(keyinput27), .C1(keyinput44), 
        .C2(ADDRESS_REG_21__SCAN_IN), .A(n5738), .ZN(n5743) );
  OAI22_X1 U6919 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(keyinput22), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(keyinput79), .ZN(n5739) );
  AOI221_X1 U6920 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput22), .C1(
        keyinput79), .C2(ADDRESS_REG_13__SCAN_IN), .A(n5739), .ZN(n5742) );
  OAI22_X1 U6921 ( .A1(UWORD_REG_14__SCAN_IN), .A2(keyinput4), .B1(keyinput47), 
        .B2(DATAI_14_), .ZN(n5740) );
  AOI221_X1 U6922 ( .B1(UWORD_REG_14__SCAN_IN), .B2(keyinput4), .C1(DATAI_14_), 
        .C2(keyinput47), .A(n5740), .ZN(n5741) );
  NAND4_X1 U6923 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n5741), .ZN(n5754)
         );
  OAI22_X1 U6924 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(keyinput90), .B1(
        INSTQUEUE_REG_6__6__SCAN_IN), .B2(keyinput78), .ZN(n5745) );
  AOI221_X1 U6925 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(keyinput90), 
        .C1(keyinput78), .C2(INSTQUEUE_REG_6__6__SCAN_IN), .A(n5745), .ZN(
        n5752) );
  OAI22_X1 U6926 ( .A1(EBX_REG_14__SCAN_IN), .A2(keyinput31), .B1(DATAI_8_), 
        .B2(keyinput116), .ZN(n5746) );
  AOI221_X1 U6927 ( .B1(EBX_REG_14__SCAN_IN), .B2(keyinput31), .C1(keyinput116), .C2(DATAI_8_), .A(n5746), .ZN(n5751) );
  OAI22_X1 U6928 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(keyinput97), .B1(
        keyinput9), .B2(EAX_REG_26__SCAN_IN), .ZN(n5747) );
  AOI221_X1 U6929 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput97), 
        .C1(EAX_REG_26__SCAN_IN), .C2(keyinput9), .A(n5747), .ZN(n5750) );
  OAI22_X1 U6930 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(keyinput100), .B1(
        keyinput74), .B2(EAX_REG_3__SCAN_IN), .ZN(n5748) );
  AOI221_X1 U6931 ( .B1(INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput100), .C1(
        EAX_REG_3__SCAN_IN), .C2(keyinput74), .A(n5748), .ZN(n5749) );
  NAND4_X1 U6932 ( .A1(n5752), .A2(n5751), .A3(n5750), .A4(n5749), .ZN(n5753)
         );
  NOR3_X1 U6933 ( .A1(n5755), .A2(n5754), .A3(n5753), .ZN(n5814) );
  OAI22_X1 U6934 ( .A1(n7050), .A2(keyinput101), .B1(n5757), .B2(keyinput73), 
        .ZN(n5756) );
  AOI221_X1 U6935 ( .B1(n7050), .B2(keyinput101), .C1(keyinput73), .C2(n5757), 
        .A(n5756), .ZN(n5767) );
  OAI22_X1 U6936 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput109), .B1(
        keyinput23), .B2(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5758) );
  AOI221_X1 U6937 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput109), .C1(
        DATAWIDTH_REG_1__SCAN_IN), .C2(keyinput23), .A(n5758), .ZN(n5766) );
  OAI22_X1 U6938 ( .A1(n6751), .A2(keyinput63), .B1(n5760), .B2(keyinput127), 
        .ZN(n5759) );
  AOI221_X1 U6939 ( .B1(n6751), .B2(keyinput63), .C1(keyinput127), .C2(n5760), 
        .A(n5759), .ZN(n5765) );
  INV_X1 U6940 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5762) );
  OAI22_X1 U6941 ( .A1(n5763), .A2(keyinput69), .B1(n5762), .B2(keyinput28), 
        .ZN(n5761) );
  AOI221_X1 U6942 ( .B1(n5763), .B2(keyinput69), .C1(keyinput28), .C2(n5762), 
        .A(n5761), .ZN(n5764) );
  NAND4_X1 U6943 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n5777)
         );
  OAI22_X1 U6944 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput30), .B1(
        keyinput13), .B2(ADS_N_REG_SCAN_IN), .ZN(n5768) );
  AOI221_X1 U6945 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput30), .C1(
        ADS_N_REG_SCAN_IN), .C2(keyinput13), .A(n5768), .ZN(n5775) );
  OAI22_X1 U6946 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(keyinput70), .B1(
        DATAO_REG_31__SCAN_IN), .B2(keyinput118), .ZN(n5769) );
  AOI221_X1 U6947 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput70), .C1(
        keyinput118), .C2(DATAO_REG_31__SCAN_IN), .A(n5769), .ZN(n5774) );
  OAI22_X1 U6948 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(keyinput21), .B1(
        keyinput26), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5770) );
  AOI221_X1 U6949 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput21), 
        .C1(PHYADDRPOINTER_REG_6__SCAN_IN), .C2(keyinput26), .A(n5770), .ZN(
        n5773) );
  OAI22_X1 U6950 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(keyinput87), .B1(
        DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput37), .ZN(n5771) );
  AOI221_X1 U6951 ( .B1(INSTQUEUE_REG_2__4__SCAN_IN), .B2(keyinput87), .C1(
        keyinput37), .C2(DATAWIDTH_REG_16__SCAN_IN), .A(n5771), .ZN(n5772) );
  NAND4_X1 U6952 ( .A1(n5775), .A2(n5774), .A3(n5773), .A4(n5772), .ZN(n5776)
         );
  NOR2_X1 U6953 ( .A1(n5777), .A2(n5776), .ZN(n5813) );
  OAI22_X1 U6954 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(keyinput20), .B1(
        keyinput77), .B2(EAX_REG_28__SCAN_IN), .ZN(n5778) );
  AOI221_X1 U6955 ( .B1(INSTQUEUE_REG_6__1__SCAN_IN), .B2(keyinput20), .C1(
        EAX_REG_28__SCAN_IN), .C2(keyinput77), .A(n5778), .ZN(n5785) );
  OAI22_X1 U6956 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(keyinput93), .B1(
        keyinput32), .B2(DATAI_19_), .ZN(n5779) );
  AOI221_X1 U6957 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput93), .C1(
        DATAI_19_), .C2(keyinput32), .A(n5779), .ZN(n5784) );
  OAI22_X1 U6958 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput25), .B1(
        UWORD_REG_0__SCAN_IN), .B2(keyinput11), .ZN(n5780) );
  AOI221_X1 U6959 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput25), .C1(keyinput11), .C2(UWORD_REG_0__SCAN_IN), .A(n5780), .ZN(n5783) );
  OAI22_X1 U6960 ( .A1(EBX_REG_27__SCAN_IN), .A2(keyinput60), .B1(
        UWORD_REG_4__SCAN_IN), .B2(keyinput75), .ZN(n5781) );
  AOI221_X1 U6961 ( .B1(EBX_REG_27__SCAN_IN), .B2(keyinput60), .C1(keyinput75), 
        .C2(UWORD_REG_4__SCAN_IN), .A(n5781), .ZN(n5782) );
  NAND4_X1 U6962 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n5792)
         );
  INV_X1 U6963 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5787) );
  AOI22_X1 U6964 ( .A1(n5787), .A2(keyinput122), .B1(keyinput12), .B2(n6111), 
        .ZN(n5786) );
  OAI221_X1 U6965 ( .B1(n5787), .B2(keyinput122), .C1(n6111), .C2(keyinput12), 
        .A(n5786), .ZN(n5791) );
  XNOR2_X1 U6966 ( .A(n3298), .B(keyinput84), .ZN(n5790) );
  XNOR2_X1 U6967 ( .A(keyinput62), .B(n5788), .ZN(n5789) );
  NOR4_X1 U6968 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n5812)
         );
  OAI22_X1 U6969 ( .A1(NA_N), .A2(keyinput54), .B1(ADDRESS_REG_25__SCAN_IN), 
        .B2(keyinput102), .ZN(n5793) );
  AOI221_X1 U6970 ( .B1(NA_N), .B2(keyinput54), .C1(keyinput102), .C2(
        ADDRESS_REG_25__SCAN_IN), .A(n5793), .ZN(n5800) );
  OAI22_X1 U6971 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(keyinput49), .B1(
        keyinput126), .B2(EAX_REG_16__SCAN_IN), .ZN(n5794) );
  AOI221_X1 U6972 ( .B1(INSTQUEUE_REG_6__3__SCAN_IN), .B2(keyinput49), .C1(
        EAX_REG_16__SCAN_IN), .C2(keyinput126), .A(n5794), .ZN(n5799) );
  OAI22_X1 U6973 ( .A1(STATE2_REG_2__SCAN_IN), .A2(keyinput57), .B1(
        INSTQUEUE_REG_4__5__SCAN_IN), .B2(keyinput35), .ZN(n5795) );
  AOI221_X1 U6974 ( .B1(STATE2_REG_2__SCAN_IN), .B2(keyinput57), .C1(
        keyinput35), .C2(INSTQUEUE_REG_4__5__SCAN_IN), .A(n5795), .ZN(n5798)
         );
  OAI22_X1 U6975 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(keyinput108), .B1(
        keyinput125), .B2(ADDRESS_REG_14__SCAN_IN), .ZN(n5796) );
  AOI221_X1 U6976 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput108), 
        .C1(ADDRESS_REG_14__SCAN_IN), .C2(keyinput125), .A(n5796), .ZN(n5797)
         );
  NAND4_X1 U6977 ( .A1(n5800), .A2(n5799), .A3(n5798), .A4(n5797), .ZN(n5810)
         );
  OAI22_X1 U6978 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(keyinput2), .B1(
        UWORD_REG_9__SCAN_IN), .B2(keyinput1), .ZN(n5801) );
  AOI221_X1 U6979 ( .B1(INSTQUEUE_REG_9__1__SCAN_IN), .B2(keyinput2), .C1(
        keyinput1), .C2(UWORD_REG_9__SCAN_IN), .A(n5801), .ZN(n5808) );
  OAI22_X1 U6980 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(keyinput59), .B1(
        keyinput7), .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5802) );
  AOI221_X1 U6981 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput59), 
        .C1(INSTQUEUE_REG_4__2__SCAN_IN), .C2(keyinput7), .A(n5802), .ZN(n5807) );
  OAI22_X1 U6982 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(keyinput67), .B1(
        keyinput0), .B2(DATAO_REG_14__SCAN_IN), .ZN(n5803) );
  AOI221_X1 U6983 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(keyinput67), 
        .C1(DATAO_REG_14__SCAN_IN), .C2(keyinput0), .A(n5803), .ZN(n5806) );
  OAI22_X1 U6984 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(keyinput71), .B1(
        INSTQUEUE_REG_14__3__SCAN_IN), .B2(keyinput34), .ZN(n5804) );
  AOI221_X1 U6985 ( .B1(INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput71), .C1(
        keyinput34), .C2(INSTQUEUE_REG_14__3__SCAN_IN), .A(n5804), .ZN(n5805)
         );
  NAND4_X1 U6986 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n5805), .ZN(n5809)
         );
  NOR2_X1 U6987 ( .A1(n5810), .A2(n5809), .ZN(n5811) );
  NAND4_X1 U6988 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n5866)
         );
  AOI22_X1 U6989 ( .A1(n5816), .A2(keyinput115), .B1(keyinput103), .B2(n5977), 
        .ZN(n5815) );
  OAI221_X1 U6990 ( .B1(n5816), .B2(keyinput115), .C1(n5977), .C2(keyinput103), 
        .A(n5815), .ZN(n5825) );
  AOI22_X1 U6991 ( .A1(n7124), .A2(keyinput33), .B1(n5818), .B2(keyinput86), 
        .ZN(n5817) );
  OAI221_X1 U6992 ( .B1(n7124), .B2(keyinput33), .C1(n5818), .C2(keyinput86), 
        .A(n5817), .ZN(n5824) );
  AOI22_X1 U6993 ( .A1(n5820), .A2(keyinput111), .B1(keyinput95), .B2(n7048), 
        .ZN(n5819) );
  OAI221_X1 U6994 ( .B1(n5820), .B2(keyinput111), .C1(n7048), .C2(keyinput95), 
        .A(n5819), .ZN(n5823) );
  INV_X1 U6995 ( .A(REIP_REG_14__SCAN_IN), .ZN(n7094) );
  AOI22_X1 U6996 ( .A1(n6791), .A2(keyinput81), .B1(keyinput3), .B2(n7094), 
        .ZN(n5821) );
  OAI221_X1 U6997 ( .B1(n6791), .B2(keyinput81), .C1(n7094), .C2(keyinput3), 
        .A(n5821), .ZN(n5822) );
  NOR4_X1 U6998 ( .A1(n5825), .A2(n5824), .A3(n5823), .A4(n5822), .ZN(n5864)
         );
  INV_X1 U6999 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n5828) );
  AOI22_X1 U7000 ( .A1(n5828), .A2(keyinput85), .B1(keyinput72), .B2(n5827), 
        .ZN(n5826) );
  OAI221_X1 U7001 ( .B1(n5828), .B2(keyinput85), .C1(n5827), .C2(keyinput72), 
        .A(n5826), .ZN(n5838) );
  INV_X1 U7002 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6571) );
  AOI22_X1 U7003 ( .A1(n6571), .A2(keyinput61), .B1(n4855), .B2(keyinput46), 
        .ZN(n5829) );
  OAI221_X1 U7004 ( .B1(n6571), .B2(keyinput61), .C1(n4855), .C2(keyinput46), 
        .A(n5829), .ZN(n5837) );
  INV_X1 U7005 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5831) );
  AOI22_X1 U7006 ( .A1(n5832), .A2(keyinput19), .B1(n5831), .B2(keyinput76), 
        .ZN(n5830) );
  OAI221_X1 U7007 ( .B1(n5832), .B2(keyinput19), .C1(n5831), .C2(keyinput76), 
        .A(n5830), .ZN(n5836) );
  INV_X1 U7008 ( .A(HOLD), .ZN(n7054) );
  AOI22_X1 U7009 ( .A1(n7054), .A2(keyinput58), .B1(keyinput80), .B2(n5834), 
        .ZN(n5833) );
  OAI221_X1 U7010 ( .B1(n7054), .B2(keyinput58), .C1(n5834), .C2(keyinput80), 
        .A(n5833), .ZN(n5835) );
  NOR4_X1 U7011 ( .A1(n5838), .A2(n5837), .A3(n5836), .A4(n5835), .ZN(n5863)
         );
  INV_X1 U7012 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6381) );
  AOI22_X1 U7013 ( .A1(n7116), .A2(keyinput55), .B1(n6381), .B2(keyinput121), 
        .ZN(n5839) );
  OAI221_X1 U7014 ( .B1(n7116), .B2(keyinput55), .C1(n6381), .C2(keyinput121), 
        .A(n5839), .ZN(n5848) );
  AOI22_X1 U7015 ( .A1(n7052), .A2(keyinput107), .B1(n5841), .B2(keyinput106), 
        .ZN(n5840) );
  OAI221_X1 U7016 ( .B1(n7052), .B2(keyinput107), .C1(n5841), .C2(keyinput106), 
        .A(n5840), .ZN(n5847) );
  AOI22_X1 U7017 ( .A1(n5843), .A2(keyinput43), .B1(n6840), .B2(keyinput123), 
        .ZN(n5842) );
  OAI221_X1 U7018 ( .B1(n5843), .B2(keyinput43), .C1(n6840), .C2(keyinput123), 
        .A(n5842), .ZN(n5846) );
  AOI22_X1 U7019 ( .A1(n5976), .A2(keyinput89), .B1(keyinput112), .B2(n6626), 
        .ZN(n5844) );
  OAI221_X1 U7020 ( .B1(n5976), .B2(keyinput89), .C1(n6626), .C2(keyinput112), 
        .A(n5844), .ZN(n5845) );
  NOR4_X1 U7021 ( .A1(n5848), .A2(n5847), .A3(n5846), .A4(n5845), .ZN(n5862)
         );
  AOI22_X1 U7022 ( .A1(n5850), .A2(keyinput105), .B1(n6062), .B2(keyinput82), 
        .ZN(n5849) );
  OAI221_X1 U7023 ( .B1(n5850), .B2(keyinput105), .C1(n6062), .C2(keyinput82), 
        .A(n5849), .ZN(n5860) );
  INV_X1 U7024 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n7046) );
  AOI22_X1 U7025 ( .A1(n7046), .A2(keyinput64), .B1(keyinput36), .B2(n7118), 
        .ZN(n5851) );
  OAI221_X1 U7026 ( .B1(n7046), .B2(keyinput64), .C1(n7118), .C2(keyinput36), 
        .A(n5851), .ZN(n5859) );
  AOI22_X1 U7027 ( .A1(n5854), .A2(keyinput40), .B1(n5853), .B2(keyinput50), 
        .ZN(n5852) );
  OAI221_X1 U7028 ( .B1(n5854), .B2(keyinput40), .C1(n5853), .C2(keyinput50), 
        .A(n5852), .ZN(n5858) );
  INV_X1 U7029 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6837) );
  INV_X1 U7030 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5856) );
  AOI22_X1 U7031 ( .A1(n6837), .A2(keyinput88), .B1(n5856), .B2(keyinput17), 
        .ZN(n5855) );
  OAI221_X1 U7032 ( .B1(n6837), .B2(keyinput88), .C1(n5856), .C2(keyinput17), 
        .A(n5855), .ZN(n5857) );
  NOR4_X1 U7033 ( .A1(n5860), .A2(n5859), .A3(n5858), .A4(n5857), .ZN(n5861)
         );
  NAND4_X1 U7034 ( .A1(n5864), .A2(n5863), .A3(n5862), .A4(n5861), .ZN(n5865)
         );
  NOR2_X1 U7035 ( .A1(n5866), .A2(n5865), .ZN(n5906) );
  AOI22_X1 U7036 ( .A1(n5869), .A2(keyinput99), .B1(keyinput41), .B2(n5868), 
        .ZN(n5867) );
  OAI221_X1 U7037 ( .B1(n5869), .B2(keyinput99), .C1(n5868), .C2(keyinput41), 
        .A(n5867), .ZN(n5878) );
  AOI22_X1 U7038 ( .A1(n6415), .A2(keyinput110), .B1(n7005), .B2(keyinput113), 
        .ZN(n5870) );
  OAI221_X1 U7039 ( .B1(n6415), .B2(keyinput110), .C1(n7005), .C2(keyinput113), 
        .A(n5870), .ZN(n5877) );
  INV_X1 U7040 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5873) );
  INV_X1 U7041 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5872) );
  AOI22_X1 U7042 ( .A1(n5873), .A2(keyinput6), .B1(n5872), .B2(keyinput92), 
        .ZN(n5871) );
  OAI221_X1 U7043 ( .B1(n5873), .B2(keyinput6), .C1(n5872), .C2(keyinput92), 
        .A(n5871), .ZN(n5876) );
  INV_X1 U7044 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6054) );
  AOI22_X1 U7045 ( .A1(n6597), .A2(keyinput24), .B1(n6054), .B2(keyinput38), 
        .ZN(n5874) );
  OAI221_X1 U7046 ( .B1(n6597), .B2(keyinput24), .C1(n6054), .C2(keyinput38), 
        .A(n5874), .ZN(n5875) );
  NOR4_X1 U7047 ( .A1(n5878), .A2(n5877), .A3(n5876), .A4(n5875), .ZN(n5905)
         );
  AOI22_X1 U7048 ( .A1(n6652), .A2(keyinput48), .B1(keyinput56), .B2(n7051), 
        .ZN(n5879) );
  OAI221_X1 U7049 ( .B1(n6652), .B2(keyinput48), .C1(n7051), .C2(keyinput56), 
        .A(n5879), .ZN(n5889) );
  AOI22_X1 U7050 ( .A1(n5881), .A2(keyinput8), .B1(keyinput98), .B2(n6035), 
        .ZN(n5880) );
  OAI221_X1 U7051 ( .B1(n5881), .B2(keyinput8), .C1(n6035), .C2(keyinput98), 
        .A(n5880), .ZN(n5888) );
  INV_X1 U7052 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5884) );
  AOI22_X1 U7053 ( .A1(n5884), .A2(keyinput68), .B1(keyinput65), .B2(n5883), 
        .ZN(n5882) );
  OAI221_X1 U7054 ( .B1(n5884), .B2(keyinput68), .C1(n5883), .C2(keyinput65), 
        .A(n5882), .ZN(n5887) );
  INV_X1 U7055 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6825) );
  AOI22_X1 U7056 ( .A1(n6834), .A2(keyinput66), .B1(n6825), .B2(keyinput117), 
        .ZN(n5885) );
  OAI221_X1 U7057 ( .B1(n6834), .B2(keyinput66), .C1(n6825), .C2(keyinput117), 
        .A(n5885), .ZN(n5886) );
  NOR4_X1 U7058 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(n5904)
         );
  AOI22_X1 U7059 ( .A1(n5891), .A2(keyinput39), .B1(keyinput5), .B2(n6622), 
        .ZN(n5890) );
  OAI221_X1 U7060 ( .B1(n5891), .B2(keyinput39), .C1(n6622), .C2(keyinput5), 
        .A(n5890), .ZN(n5902) );
  INV_X1 U7061 ( .A(DATAI_23_), .ZN(n5894) );
  AOI22_X1 U7062 ( .A1(n5894), .A2(keyinput96), .B1(n5893), .B2(keyinput119), 
        .ZN(n5892) );
  OAI221_X1 U7063 ( .B1(n5894), .B2(keyinput96), .C1(n5893), .C2(keyinput119), 
        .A(n5892), .ZN(n5901) );
  AOI22_X1 U7064 ( .A1(n5897), .A2(keyinput45), .B1(n5896), .B2(keyinput29), 
        .ZN(n5895) );
  OAI221_X1 U7065 ( .B1(n5897), .B2(keyinput45), .C1(n5896), .C2(keyinput29), 
        .A(n5895), .ZN(n5900) );
  INV_X1 U7066 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7088) );
  INV_X1 U7067 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7123) );
  AOI22_X1 U7068 ( .A1(n7088), .A2(keyinput16), .B1(keyinput104), .B2(n7123), 
        .ZN(n5898) );
  OAI221_X1 U7069 ( .B1(n7088), .B2(keyinput16), .C1(n7123), .C2(keyinput104), 
        .A(n5898), .ZN(n5899) );
  NOR4_X1 U7070 ( .A1(n5902), .A2(n5901), .A3(n5900), .A4(n5899), .ZN(n5903)
         );
  NAND4_X1 U7071 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n5907)
         );
  NOR2_X1 U7072 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  INV_X1 U7073 ( .A(n6065), .ZN(n5931) );
  NAND2_X1 U7074 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n6305) );
  INV_X1 U7075 ( .A(n6305), .ZN(n5921) );
  NAND3_X1 U7076 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        n5910), .ZN(n5911) );
  NOR3_X1 U7077 ( .A1(n5913), .A2(n5912), .A3(n5911), .ZN(n5989) );
  AND2_X1 U7078 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5989), .ZN(n5925) );
  NAND2_X1 U7079 ( .A1(n6504), .A2(n5925), .ZN(n5914) );
  NAND2_X1 U7080 ( .A1(n5915), .A2(n5914), .ZN(n5991) );
  OR2_X1 U7081 ( .A1(n6507), .A2(REIP_REG_24__SCAN_IN), .ZN(n5916) );
  AND2_X1 U7082 ( .A1(n5991), .A2(n5916), .ZN(n5972) );
  INV_X1 U7083 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7115) );
  NOR2_X1 U7084 ( .A1(n7115), .A2(n7116), .ZN(n5917) );
  OR2_X1 U7085 ( .A1(n6507), .A2(n5917), .ZN(n5918) );
  AND2_X1 U7086 ( .A1(n5972), .A2(n5918), .ZN(n6311) );
  INV_X1 U7087 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7121) );
  NOR2_X1 U7088 ( .A1(n7118), .A2(n7121), .ZN(n5919) );
  OR2_X1 U7089 ( .A1(n6507), .A2(n5919), .ZN(n5920) );
  NAND2_X1 U7090 ( .A1(n6311), .A2(n5920), .ZN(n6303) );
  INV_X1 U7091 ( .A(n6303), .ZN(n5946) );
  OAI21_X1 U7092 ( .B1(n6507), .B2(n5921), .A(n5946), .ZN(n5928) );
  INV_X1 U7093 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5924) );
  OAI22_X1 U7094 ( .A1(n5990), .A2(n5924), .B1(n5923), .B2(n5922), .ZN(n5927)
         );
  NAND2_X1 U7095 ( .A1(n6532), .A2(n5925), .ZN(n5982) );
  NOR2_X1 U7096 ( .A1(n5982), .A2(n5976), .ZN(n5968) );
  NAND2_X1 U7097 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5968), .ZN(n6312) );
  NOR2_X1 U7098 ( .A1(n7116), .A2(n6312), .ZN(n5961) );
  NAND3_X1 U7099 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .A3(
        n5961), .ZN(n5934) );
  NOR3_X1 U7100 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6305), .A3(n5934), .ZN(n5926) );
  AOI211_X1 U7101 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5928), .A(n5927), .B(n5926), .ZN(n5930) );
  NAND2_X1 U7102 ( .A1(n6026), .A2(n6539), .ZN(n5929) );
  OAI211_X1 U7103 ( .C1(n5931), .C2(n6515), .A(n5930), .B(n5929), .ZN(U2796)
         );
  NAND2_X1 U7104 ( .A1(n5939), .A2(n5932), .ZN(n5933) );
  AOI22_X1 U7105 ( .A1(n6087), .A2(n6518), .B1(REIP_REG_29__SCAN_IN), .B2(
        n6303), .ZN(n5936) );
  INV_X1 U7106 ( .A(n5934), .ZN(n6306) );
  AOI22_X1 U7107 ( .A1(EBX_REG_29__SCAN_IN), .A2(n6543), .B1(n6306), .B2(n7124), .ZN(n5935) );
  OAI211_X1 U7108 ( .C1(n6084), .C2(n5990), .A(n5936), .B(n5935), .ZN(n5937)
         );
  AOI21_X1 U7109 ( .B1(n6034), .B2(n6539), .A(n5937), .ZN(n5938) );
  OAI21_X1 U7110 ( .B1(n6085), .B2(n6515), .A(n5938), .ZN(U2798) );
  OAI21_X1 U7111 ( .B1(n5951), .B2(n5940), .A(n5939), .ZN(n6093) );
  AND3_X1 U7112 ( .A1(n7121), .A2(REIP_REG_27__SCAN_IN), .A3(n5961), .ZN(n5942) );
  OAI22_X1 U7113 ( .A1(n6037), .A2(n6522), .B1(n6095), .B2(n6541), .ZN(n5941)
         );
  AOI211_X1 U7114 ( .C1(n6525), .C2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5942), 
        .B(n5941), .ZN(n5949) );
  NAND2_X1 U7115 ( .A1(n5956), .A2(n5943), .ZN(n5944) );
  NAND2_X1 U7116 ( .A1(n5945), .A2(n5944), .ZN(n6183) );
  OAI22_X1 U7117 ( .A1(n6183), .A2(n6527), .B1(n5946), .B2(n7121), .ZN(n5947)
         );
  INV_X1 U7118 ( .A(n5947), .ZN(n5948) );
  OAI211_X1 U7119 ( .C1(n6093), .C2(n6515), .A(n5949), .B(n5948), .ZN(U2799)
         );
  INV_X1 U7120 ( .A(n5951), .ZN(n5952) );
  OAI21_X1 U7121 ( .B1(n5953), .B2(n5950), .A(n5952), .ZN(n6102) );
  OR2_X1 U7122 ( .A1(n6049), .A2(n5954), .ZN(n5955) );
  NAND2_X1 U7123 ( .A1(n5956), .A2(n5955), .ZN(n6191) );
  OAI22_X1 U7124 ( .A1(n6040), .A2(n6522), .B1(n6101), .B2(n5990), .ZN(n5958)
         );
  NOR2_X1 U7125 ( .A1(n6311), .A2(n7118), .ZN(n5957) );
  AOI211_X1 U7126 ( .C1(n6105), .C2(n6518), .A(n5958), .B(n5957), .ZN(n5959)
         );
  OAI21_X1 U7127 ( .B1(n6191), .B2(n6527), .A(n5959), .ZN(n5960) );
  AOI21_X1 U7128 ( .B1(n5961), .B2(n7118), .A(n5960), .ZN(n5962) );
  OAI21_X1 U7129 ( .B1(n6102), .B2(n6515), .A(n5962), .ZN(U2800) );
  AOI21_X1 U7130 ( .B1(n5964), .B2(n5963), .A(n6044), .ZN(n5965) );
  INV_X1 U7131 ( .A(n5965), .ZN(n6119) );
  OAI21_X1 U7132 ( .B1(n5996), .B2(n5975), .A(n5966), .ZN(n5967) );
  AND2_X1 U7133 ( .A1(n5967), .A2(n6047), .ZN(n6209) );
  NAND2_X1 U7134 ( .A1(n5968), .A2(n7115), .ZN(n5971) );
  INV_X1 U7135 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6053) );
  OAI22_X1 U7136 ( .A1(n6053), .A2(n6522), .B1(n6111), .B2(n5990), .ZN(n5969)
         );
  AOI21_X1 U7137 ( .B1(n6518), .B2(n6113), .A(n5969), .ZN(n5970) );
  OAI211_X1 U7138 ( .C1(n5972), .C2(n7115), .A(n5971), .B(n5970), .ZN(n5973)
         );
  AOI21_X1 U7139 ( .B1(n6209), .B2(n6539), .A(n5973), .ZN(n5974) );
  OAI21_X1 U7140 ( .B1(n6119), .B2(n6515), .A(n5974), .ZN(U2802) );
  XNOR2_X1 U7141 ( .A(n5996), .B(n5975), .ZN(n6218) );
  INV_X1 U7142 ( .A(n6218), .ZN(n5984) );
  OAI22_X1 U7143 ( .A1(n5977), .A2(n5990), .B1(n5976), .B2(n5991), .ZN(n5980)
         );
  NOR2_X1 U7144 ( .A1(n6541), .A2(n5978), .ZN(n5979) );
  AOI211_X1 U7145 ( .C1(n6543), .C2(EBX_REG_24__SCAN_IN), .A(n5980), .B(n5979), 
        .ZN(n5981) );
  OAI21_X1 U7146 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5982), .A(n5981), .ZN(n5983) );
  AOI21_X1 U7147 ( .B1(n5984), .B2(n6539), .A(n5983), .ZN(n5985) );
  OAI21_X1 U7148 ( .B1(n6340), .B2(n6515), .A(n5985), .ZN(U2803) );
  INV_X1 U7149 ( .A(n5986), .ZN(n5987) );
  AOI21_X1 U7150 ( .B1(n5988), .B2(n6005), .A(n5987), .ZN(n6127) );
  INV_X1 U7151 ( .A(n6127), .ZN(n6076) );
  AOI21_X1 U7152 ( .B1(n6532), .B2(n5989), .A(REIP_REG_23__SCAN_IN), .ZN(n5992) );
  OAI22_X1 U7153 ( .A1(n5992), .A2(n5991), .B1(n6124), .B2(n5990), .ZN(n5995)
         );
  INV_X1 U7154 ( .A(n6126), .ZN(n5993) );
  NOR2_X1 U7155 ( .A1(n6541), .A2(n5993), .ZN(n5994) );
  AOI211_X1 U7156 ( .C1(EBX_REG_23__SCAN_IN), .C2(n6543), .A(n5995), .B(n5994), 
        .ZN(n6001) );
  INV_X1 U7157 ( .A(n6010), .ZN(n5998) );
  INV_X1 U7158 ( .A(n5996), .ZN(n5997) );
  AOI21_X1 U7159 ( .B1(n5999), .B2(n5998), .A(n5997), .ZN(n6226) );
  NAND2_X1 U7160 ( .A1(n6226), .A2(n6539), .ZN(n6000) );
  OAI211_X1 U7161 ( .C1(n6076), .C2(n6515), .A(n6001), .B(n6000), .ZN(U2804)
         );
  OR2_X1 U7162 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  NAND2_X1 U7163 ( .A1(n6005), .A2(n6004), .ZN(n6346) );
  AOI21_X1 U7164 ( .B1(n6006), .B2(n6325), .A(n7108), .ZN(n6017) );
  NOR2_X1 U7165 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  OR2_X1 U7166 ( .A1(n6010), .A2(n6009), .ZN(n6236) );
  NAND3_X1 U7167 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6011), .A3(n7108), .ZN(
        n6015) );
  AOI22_X1 U7168 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6543), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6525), .ZN(n6012) );
  INV_X1 U7169 ( .A(n6012), .ZN(n6013) );
  AOI21_X1 U7170 ( .B1(n6518), .B2(n6136), .A(n6013), .ZN(n6014) );
  OAI211_X1 U7171 ( .C1(n6236), .C2(n6527), .A(n6015), .B(n6014), .ZN(n6016)
         );
  NOR2_X1 U7172 ( .A1(n6017), .A2(n6016), .ZN(n6018) );
  OAI21_X1 U7173 ( .B1(n6346), .B2(n6515), .A(n6018), .ZN(U2805) );
  NAND2_X1 U7174 ( .A1(n6552), .A2(n6503), .ZN(n6025) );
  AOI22_X1 U7175 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6543), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6434), .ZN(n6024) );
  AOI21_X1 U7176 ( .B1(n6525), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6524), 
        .ZN(n6019) );
  OAI21_X1 U7177 ( .B1(n6541), .B2(n6362), .A(n6019), .ZN(n6020) );
  AOI21_X1 U7178 ( .B1(n6377), .B2(n6539), .A(n6020), .ZN(n6023) );
  INV_X1 U7179 ( .A(n6021), .ZN(n6022) );
  NAND4_X1 U7180 ( .A1(n6025), .A2(n6024), .A3(n6023), .A4(n6022), .ZN(U2809)
         );
  INV_X1 U7181 ( .A(n6026), .ZN(n6028) );
  OAI22_X1 U7182 ( .A1(n6028), .A2(n6060), .B1(n6027), .B2(n6063), .ZN(U2828)
         );
  INV_X1 U7183 ( .A(n6331), .ZN(n6033) );
  AOI22_X1 U7184 ( .A1(n6304), .A2(n6056), .B1(EBX_REG_30__SCAN_IN), .B2(n6055), .ZN(n6032) );
  OAI21_X1 U7185 ( .B1(n6033), .B2(n6058), .A(n6032), .ZN(U2829) );
  INV_X1 U7186 ( .A(n6034), .ZN(n6036) );
  OAI222_X1 U7187 ( .A1(n6060), .A2(n6036), .B1(n6063), .B2(n6035), .C1(n6058), 
        .C2(n6085), .ZN(U2830) );
  OAI22_X1 U7188 ( .A1(n6183), .A2(n6060), .B1(n6037), .B2(n6063), .ZN(n6038)
         );
  INV_X1 U7189 ( .A(n6038), .ZN(n6039) );
  OAI21_X1 U7190 ( .B1(n6093), .B2(n6058), .A(n6039), .ZN(U2831) );
  OAI22_X1 U7191 ( .A1(n6191), .A2(n6060), .B1(n6040), .B2(n6063), .ZN(n6041)
         );
  INV_X1 U7192 ( .A(n6041), .ZN(n6042) );
  OAI21_X1 U7193 ( .B1(n6102), .B2(n6058), .A(n6042), .ZN(U2832) );
  INV_X1 U7194 ( .A(n5950), .ZN(n6043) );
  OAI21_X1 U7195 ( .B1(n6045), .B2(n6044), .A(n6043), .ZN(n6314) );
  AND2_X1 U7196 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  NOR2_X1 U7197 ( .A1(n6049), .A2(n6048), .ZN(n6316) );
  NOR2_X1 U7198 ( .A1(n6063), .A2(n6320), .ZN(n6050) );
  AOI21_X1 U7199 ( .B1(n6316), .B2(n6056), .A(n6050), .ZN(n6051) );
  OAI21_X1 U7200 ( .B1(n6314), .B2(n6058), .A(n6051), .ZN(U2833) );
  INV_X1 U7201 ( .A(n6209), .ZN(n6052) );
  OAI222_X1 U7202 ( .A1(n6058), .A2(n6119), .B1(n6063), .B2(n6053), .C1(n6052), 
        .C2(n6060), .ZN(U2834) );
  OAI222_X1 U7203 ( .A1(n6058), .A2(n6340), .B1(n6060), .B2(n6218), .C1(n6063), 
        .C2(n6054), .ZN(U2835) );
  AOI22_X1 U7204 ( .A1(n6226), .A2(n6056), .B1(n6055), .B2(EBX_REG_23__SCAN_IN), .ZN(n6057) );
  OAI21_X1 U7205 ( .B1(n6076), .B2(n6058), .A(n6057), .ZN(U2836) );
  OAI222_X1 U7206 ( .A1(n6060), .A2(n6236), .B1(n6063), .B2(n6059), .C1(n6058), 
        .C2(n6346), .ZN(U2837) );
  INV_X1 U7207 ( .A(n6366), .ZN(n6061) );
  OAI222_X1 U7208 ( .A1(n6058), .A2(n6145), .B1(n6063), .B2(n6062), .C1(n6061), 
        .C2(n6060), .ZN(U2838) );
  NAND3_X1 U7209 ( .A1(n6065), .A2(n4149), .A3(n6064), .ZN(n6067) );
  AOI22_X1 U7210 ( .A1(n6558), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6561), .ZN(n6066) );
  NAND2_X1 U7211 ( .A1(n6067), .A2(n6066), .ZN(U2860) );
  AOI22_X1 U7212 ( .A1(n6558), .A2(DATAI_29_), .B1(n6561), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7213 ( .A1(n6562), .A2(DATAI_13_), .ZN(n6068) );
  OAI211_X1 U7214 ( .C1(n6085), .C2(n6345), .A(n6069), .B(n6068), .ZN(U2862)
         );
  AOI22_X1 U7215 ( .A1(n6558), .A2(DATAI_27_), .B1(n6561), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7216 ( .A1(n6562), .A2(DATAI_11_), .ZN(n6070) );
  OAI211_X1 U7217 ( .C1(n6102), .C2(n6345), .A(n6071), .B(n6070), .ZN(U2864)
         );
  AOI22_X1 U7218 ( .A1(n6558), .A2(DATAI_25_), .B1(n6561), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7219 ( .A1(n6562), .A2(DATAI_9_), .ZN(n6072) );
  OAI211_X1 U7220 ( .C1(n6119), .C2(n6345), .A(n6073), .B(n6072), .ZN(U2866)
         );
  AOI22_X1 U7221 ( .A1(n6558), .A2(DATAI_23_), .B1(n6561), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7222 ( .A1(n6562), .A2(DATAI_7_), .ZN(n6074) );
  OAI211_X1 U7223 ( .C1(n6076), .C2(n6345), .A(n6075), .B(n6074), .ZN(U2868)
         );
  NAND2_X1 U7224 ( .A1(n6331), .A2(n6698), .ZN(n6081) );
  NOR2_X1 U7225 ( .A1(n6162), .A2(n6077), .ZN(n6078) );
  AOI211_X1 U7226 ( .C1(n6302), .C2(n6663), .A(n6079), .B(n6078), .ZN(n6080)
         );
  OAI211_X1 U7227 ( .C1(n6082), .C2(n6681), .A(n6081), .B(n6080), .ZN(U2956)
         );
  OAI21_X1 U7228 ( .B1(n6162), .B2(n6084), .A(n6083), .ZN(n6086) );
  NAND3_X1 U7229 ( .A1(n6089), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n6263), .ZN(n6091) );
  NOR2_X1 U7230 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6198) );
  NAND3_X1 U7231 ( .A1(n6116), .A2(n6131), .A3(n6198), .ZN(n6098) );
  AOI22_X1 U7232 ( .A1(n6091), .A2(n6098), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6204), .ZN(n6092) );
  XNOR2_X1 U7233 ( .A(n6092), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6186)
         );
  INV_X1 U7234 ( .A(n6093), .ZN(n6334) );
  NAND2_X1 U7235 ( .A1(n6803), .A2(REIP_REG_28__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7236 ( .A1(n6694), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6094)
         );
  OAI211_X1 U7237 ( .C1(n6704), .C2(n6095), .A(n6182), .B(n6094), .ZN(n6096)
         );
  AOI21_X1 U7238 ( .B1(n6334), .B2(n6698), .A(n6096), .ZN(n6097) );
  OAI21_X1 U7239 ( .B1(n6186), .B2(n6681), .A(n6097), .ZN(U2958) );
  NAND2_X1 U7240 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  XNOR2_X1 U7241 ( .A(n6100), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6195)
         );
  NAND2_X1 U7242 ( .A1(n6803), .A2(REIP_REG_27__SCAN_IN), .ZN(n6190) );
  OAI21_X1 U7243 ( .B1(n6162), .B2(n6101), .A(n6190), .ZN(n6104) );
  NOR2_X1 U7244 ( .A1(n6102), .A2(n6679), .ZN(n6103) );
  AOI211_X1 U7245 ( .C1(n6663), .C2(n6105), .A(n6104), .B(n6103), .ZN(n6106)
         );
  OAI21_X1 U7246 ( .B1(n6195), .B2(n6681), .A(n6106), .ZN(U2959) );
  XNOR2_X1 U7247 ( .A(n6262), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6107)
         );
  XNOR2_X1 U7248 ( .A(n3740), .B(n6107), .ZN(n6196) );
  NAND2_X1 U7249 ( .A1(n6196), .A2(n6700), .ZN(n6110) );
  NOR2_X1 U7250 ( .A1(n6774), .A2(n7116), .ZN(n6201) );
  NOR2_X1 U7251 ( .A1(n6704), .A2(n6315), .ZN(n6108) );
  AOI211_X1 U7252 ( .C1(n6694), .C2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6201), 
        .B(n6108), .ZN(n6109) );
  OAI211_X1 U7253 ( .C1(n6679), .C2(n6314), .A(n6110), .B(n6109), .ZN(U2960)
         );
  NAND2_X1 U7254 ( .A1(n6803), .A2(REIP_REG_25__SCAN_IN), .ZN(n6206) );
  OAI21_X1 U7255 ( .B1(n6162), .B2(n6111), .A(n6206), .ZN(n6112) );
  AOI21_X1 U7256 ( .B1(n6663), .B2(n6113), .A(n6112), .ZN(n6118) );
  OAI21_X1 U7257 ( .B1(n6116), .B2(n6115), .A(n6114), .ZN(n6205) );
  NAND2_X1 U7258 ( .A1(n6205), .A2(n6700), .ZN(n6117) );
  OAI211_X1 U7259 ( .C1(n6119), .C2(n6679), .A(n6118), .B(n6117), .ZN(U2961)
         );
  NOR2_X1 U7260 ( .A1(n6121), .A2(n6120), .ZN(n6123) );
  XNOR2_X1 U7261 ( .A(n6123), .B(n6122), .ZN(n6230) );
  INV_X1 U7262 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7111) );
  NOR2_X1 U7263 ( .A1(n6774), .A2(n7111), .ZN(n6225) );
  NOR2_X1 U7264 ( .A1(n6162), .A2(n6124), .ZN(n6125) );
  AOI211_X1 U7265 ( .C1(n6663), .C2(n6126), .A(n6225), .B(n6125), .ZN(n6129)
         );
  NAND2_X1 U7266 ( .A1(n6127), .A2(n6698), .ZN(n6128) );
  OAI211_X1 U7267 ( .C1(n6230), .C2(n6681), .A(n6129), .B(n6128), .ZN(U2963)
         );
  OAI21_X1 U7268 ( .B1(n6131), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6130), 
        .ZN(n6133) );
  XNOR2_X1 U7269 ( .A(n6131), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6132)
         );
  XNOR2_X1 U7270 ( .A(n6133), .B(n6132), .ZN(n6239) );
  NAND2_X1 U7271 ( .A1(n6785), .A2(REIP_REG_22__SCAN_IN), .ZN(n6235) );
  OAI21_X1 U7272 ( .B1(n6162), .B2(n5640), .A(n6235), .ZN(n6135) );
  NOR2_X1 U7273 ( .A1(n6346), .A2(n6679), .ZN(n6134) );
  AOI211_X1 U7274 ( .C1(n6663), .C2(n6136), .A(n6135), .B(n6134), .ZN(n6137)
         );
  OAI21_X1 U7275 ( .B1(n6239), .B2(n6681), .A(n6137), .ZN(U2964) );
  OAI21_X1 U7276 ( .B1(n6139), .B2(n6138), .A(n6130), .ZN(n6367) );
  NAND2_X1 U7277 ( .A1(n6367), .A2(n6700), .ZN(n6144) );
  OAI22_X1 U7278 ( .A1(n6162), .A2(n6140), .B1(n6774), .B2(n7107), .ZN(n6141)
         );
  AOI21_X1 U7279 ( .B1(n6663), .B2(n6142), .A(n6141), .ZN(n6143) );
  OAI211_X1 U7280 ( .C1(n6679), .C2(n6145), .A(n6144), .B(n6143), .ZN(U2965)
         );
  OR2_X1 U7281 ( .A1(n6146), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6150)
         );
  INV_X1 U7282 ( .A(n6147), .ZN(n6148) );
  NAND2_X1 U7283 ( .A1(n6148), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6149) );
  MUX2_X1 U7284 ( .A(n6150), .B(n6149), .S(n6263), .Z(n6151) );
  XOR2_X1 U7285 ( .A(n6151), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n6253) );
  INV_X1 U7286 ( .A(n6330), .ZN(n6154) );
  INV_X1 U7287 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7288 ( .A1(n6785), .A2(REIP_REG_20__SCAN_IN), .ZN(n6250) );
  OAI21_X1 U7289 ( .B1(n6162), .B2(n6152), .A(n6250), .ZN(n6153) );
  AOI21_X1 U7290 ( .B1(n6663), .B2(n6154), .A(n6153), .ZN(n6157) );
  NAND2_X1 U7291 ( .A1(n6350), .A2(n6698), .ZN(n6156) );
  OAI211_X1 U7292 ( .C1(n6253), .C2(n6681), .A(n6157), .B(n6156), .ZN(U2966)
         );
  XNOR2_X1 U7293 ( .A(n6262), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6158)
         );
  XNOR2_X1 U7294 ( .A(n6146), .B(n6158), .ZN(n6261) );
  NAND2_X1 U7295 ( .A1(n6663), .A2(n6159), .ZN(n6160) );
  NAND2_X1 U7296 ( .A1(n6785), .A2(REIP_REG_19__SCAN_IN), .ZN(n6255) );
  OAI211_X1 U7297 ( .C1(n6162), .C2(n6161), .A(n6160), .B(n6255), .ZN(n6163)
         );
  AOI21_X1 U7298 ( .B1(n6353), .B2(n6698), .A(n6163), .ZN(n6164) );
  OAI21_X1 U7299 ( .B1(n6261), .B2(n6681), .A(n6164), .ZN(U2967) );
  OAI21_X1 U7300 ( .B1(n6263), .B2(n6391), .A(n6165), .ZN(n6166) );
  XOR2_X1 U7301 ( .A(n6166), .B(n6264), .Z(n6386) );
  AOI22_X1 U7302 ( .A1(n6694), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6785), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n6167) );
  OAI21_X1 U7303 ( .B1(n6704), .B2(n6168), .A(n6167), .ZN(n6169) );
  AOI21_X1 U7304 ( .B1(n6560), .B2(n6698), .A(n6169), .ZN(n6170) );
  OAI21_X1 U7305 ( .B1(n6386), .B2(n6681), .A(n6170), .ZN(U2970) );
  XNOR2_X1 U7306 ( .A(n6262), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6171)
         );
  XNOR2_X1 U7307 ( .A(n6172), .B(n6171), .ZN(n6398) );
  NAND2_X1 U7308 ( .A1(n6398), .A2(n6700), .ZN(n6176) );
  AND2_X1 U7309 ( .A1(n6785), .A2(REIP_REG_15__SCAN_IN), .ZN(n6395) );
  NOR2_X1 U7310 ( .A1(n6173), .A2(n6704), .ZN(n6174) );
  AOI211_X1 U7311 ( .C1(n6694), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6395), 
        .B(n6174), .ZN(n6175) );
  OAI211_X1 U7312 ( .C1(n6679), .C2(n6177), .A(n6176), .B(n6175), .ZN(U2971)
         );
  INV_X1 U7313 ( .A(n6178), .ZN(n6193) );
  XNOR2_X1 U7314 ( .A(n6179), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6180)
         );
  NAND2_X1 U7315 ( .A1(n6188), .A2(n6180), .ZN(n6181) );
  OAI211_X1 U7316 ( .C1(n6183), .C2(n6775), .A(n6182), .B(n6181), .ZN(n6184)
         );
  AOI21_X1 U7317 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n6193), .A(n6184), 
        .ZN(n6185) );
  OAI21_X1 U7318 ( .B1(n6186), .B2(n6773), .A(n6185), .ZN(U2990) );
  INV_X1 U7319 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7320 ( .A1(n6188), .A2(n6187), .ZN(n6189) );
  OAI211_X1 U7321 ( .C1(n6191), .C2(n6775), .A(n6190), .B(n6189), .ZN(n6192)
         );
  AOI21_X1 U7322 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6193), .A(n6192), 
        .ZN(n6194) );
  OAI21_X1 U7323 ( .B1(n6195), .B2(n6773), .A(n6194), .ZN(U2991) );
  NAND2_X1 U7324 ( .A1(n6196), .A2(n6801), .ZN(n6203) );
  INV_X1 U7325 ( .A(n6197), .ZN(n6207) );
  NOR3_X1 U7326 ( .A1(n6207), .A2(n6199), .A3(n6198), .ZN(n6200) );
  AOI211_X1 U7327 ( .C1(n6316), .C2(n6799), .A(n6201), .B(n6200), .ZN(n6202)
         );
  OAI211_X1 U7328 ( .C1(n6214), .C2(n6204), .A(n6203), .B(n6202), .ZN(U2992)
         );
  NAND2_X1 U7329 ( .A1(n6205), .A2(n6801), .ZN(n6211) );
  OAI21_X1 U7330 ( .B1(n6207), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6206), 
        .ZN(n6208) );
  AOI21_X1 U7331 ( .B1(n6209), .B2(n6799), .A(n6208), .ZN(n6210) );
  OAI211_X1 U7332 ( .C1(n6214), .C2(n6212), .A(n6211), .B(n6210), .ZN(U2993)
         );
  NAND2_X1 U7333 ( .A1(n6213), .A2(n6375), .ZN(n6233) );
  INV_X1 U7334 ( .A(n6233), .ZN(n6371) );
  NAND3_X1 U7335 ( .A1(n6371), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n6231), .ZN(n6215) );
  AOI21_X1 U7336 ( .B1(n6216), .B2(n6215), .A(n6214), .ZN(n6220) );
  OAI21_X1 U7337 ( .B1(n6218), .B2(n6775), .A(n6217), .ZN(n6219) );
  AOI211_X1 U7338 ( .C1(n6221), .C2(n6801), .A(n6220), .B(n6219), .ZN(n6222)
         );
  INV_X1 U7339 ( .A(n6222), .ZN(U2994) );
  NOR3_X1 U7340 ( .A1(n6233), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n6223), 
        .ZN(n6224) );
  AOI211_X1 U7341 ( .C1(n6226), .C2(n6799), .A(n6225), .B(n6224), .ZN(n6229)
         );
  NAND2_X1 U7342 ( .A1(n6227), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6228) );
  OAI211_X1 U7343 ( .C1(n6230), .C2(n6773), .A(n6229), .B(n6228), .ZN(U2995)
         );
  OR3_X1 U7344 ( .A1(n6233), .A2(n6232), .A3(n6231), .ZN(n6234) );
  OAI211_X1 U7345 ( .C1(n6236), .C2(n6775), .A(n6235), .B(n6234), .ZN(n6237)
         );
  AOI21_X1 U7346 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6369), .A(n6237), 
        .ZN(n6238) );
  OAI21_X1 U7347 ( .B1(n6239), .B2(n6773), .A(n6238), .ZN(U2996) );
  INV_X1 U7348 ( .A(n6240), .ZN(n6245) );
  OAI21_X1 U7349 ( .B1(n6374), .B2(n6242), .A(n6241), .ZN(n6243) );
  NAND2_X1 U7350 ( .A1(n6244), .A2(n6243), .ZN(n6267) );
  AOI21_X1 U7351 ( .B1(n6245), .B2(n6374), .A(n6267), .ZN(n6382) );
  OAI21_X1 U7352 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6383), .A(n6382), 
        .ZN(n6259) );
  XNOR2_X1 U7353 ( .A(n6246), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6248)
         );
  NAND2_X1 U7354 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  OAI211_X1 U7355 ( .C1(n6324), .C2(n6775), .A(n6250), .B(n6249), .ZN(n6251)
         );
  AOI21_X1 U7356 ( .B1(n6259), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n6251), 
        .ZN(n6252) );
  OAI21_X1 U7357 ( .B1(n6253), .B2(n6773), .A(n6252), .ZN(U2998) );
  NAND2_X1 U7358 ( .A1(n6254), .A2(n6799), .ZN(n6256) );
  OAI211_X1 U7359 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6257), .A(n6256), .B(n6255), .ZN(n6258) );
  AOI21_X1 U7360 ( .B1(n6259), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6258), 
        .ZN(n6260) );
  OAI21_X1 U7361 ( .B1(n6261), .B2(n6773), .A(n6260), .ZN(U2999) );
  NOR3_X1 U7362 ( .A1(n6264), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6262), 
        .ZN(n6358) );
  NAND3_X1 U7363 ( .A1(n6264), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6263), .ZN(n6356) );
  INV_X1 U7364 ( .A(n6356), .ZN(n6265) );
  NOR2_X1 U7365 ( .A1(n6358), .A2(n6265), .ZN(n6266) );
  XNOR2_X1 U7366 ( .A(n6266), .B(n6374), .ZN(n6365) );
  AOI22_X1 U7367 ( .A1(n6803), .A2(REIP_REG_17__SCAN_IN), .B1(n6375), .B2(
        n6374), .ZN(n6269) );
  NAND2_X1 U7368 ( .A1(n6267), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6268) );
  OAI211_X1 U7369 ( .C1(n6431), .C2(n6775), .A(n6269), .B(n6268), .ZN(n6270)
         );
  INV_X1 U7370 ( .A(n6270), .ZN(n6271) );
  OAI21_X1 U7371 ( .B1(n6365), .B2(n6773), .A(n6271), .ZN(U3001) );
  AOI22_X1 U7372 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6274), .B1(n6273), .B2(n6272), .ZN(n6279) );
  INV_X1 U7373 ( .A(n6275), .ZN(n6454) );
  INV_X1 U7374 ( .A(n6276), .ZN(n6277) );
  AOI21_X1 U7375 ( .B1(n6454), .B2(n6799), .A(n6277), .ZN(n6278) );
  OAI211_X1 U7376 ( .C1(n6280), .C2(n6773), .A(n6279), .B(n6278), .ZN(U3005)
         );
  NOR2_X1 U7377 ( .A1(n3196), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6282) );
  OAI22_X1 U7378 ( .A1(n6921), .A2(n6282), .B1(n6281), .B2(n6292), .ZN(n6283)
         );
  MUX2_X1 U7379 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6283), .S(n6810), 
        .Z(U3464) );
  XNOR2_X1 U7380 ( .A(n6288), .B(n6284), .ZN(n6286) );
  INV_X1 U7381 ( .A(n4060), .ZN(n6285) );
  OAI22_X1 U7382 ( .A1(n6286), .A2(n6927), .B1(n6285), .B2(n6292), .ZN(n6287)
         );
  MUX2_X1 U7383 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6287), .S(n6810), 
        .Z(U3463) );
  INV_X1 U7384 ( .A(n6288), .ZN(n6290) );
  AOI21_X1 U7385 ( .B1(n6291), .B2(n6290), .A(n6289), .ZN(n6293) );
  OAI222_X1 U7386 ( .A1(n6858), .A2(n6294), .B1(n6927), .B2(n6293), .C1(n6292), 
        .C2(n6546), .ZN(n6295) );
  MUX2_X1 U7387 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6295), .S(n6810), 
        .Z(U3462) );
  INV_X1 U7388 ( .A(n6296), .ZN(n6299) );
  OAI22_X1 U7389 ( .A1(n6299), .A2(n7147), .B1(n6298), .B2(n6297), .ZN(n6300)
         );
  MUX2_X1 U7390 ( .A(n6301), .B(n6300), .S(n7145), .Z(U3456) );
  AND2_X1 U7391 ( .A1(DATAO_REG_31__SCAN_IN), .A2(n6594), .ZN(U2892) );
  AOI22_X1 U7392 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6303), .B1(n6302), .B2(
        n6518), .ZN(n6310) );
  AOI22_X1 U7393 ( .A1(EBX_REG_30__SCAN_IN), .A2(n6543), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6525), .ZN(n6309) );
  AOI22_X1 U7394 ( .A1(n6331), .A2(n6503), .B1(n6304), .B2(n6539), .ZN(n6308)
         );
  OAI211_X1 U7395 ( .C1(REIP_REG_30__SCAN_IN), .C2(REIP_REG_29__SCAN_IN), .A(
        n6306), .B(n6305), .ZN(n6307) );
  AOI21_X1 U7396 ( .B1(n7116), .B2(n6312), .A(n6311), .ZN(n6313) );
  AOI21_X1 U7397 ( .B1(n6525), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6313), 
        .ZN(n6319) );
  INV_X1 U7398 ( .A(n6314), .ZN(n6337) );
  INV_X1 U7399 ( .A(n6315), .ZN(n6317) );
  AOI222_X1 U7400 ( .A1(n6337), .A2(n6503), .B1(n6317), .B2(n6518), .C1(n6316), 
        .C2(n6539), .ZN(n6318) );
  OAI211_X1 U7401 ( .C1(n6320), .C2(n6522), .A(n6319), .B(n6318), .ZN(U2801)
         );
  AOI22_X1 U7402 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6543), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6525), .ZN(n6329) );
  INV_X1 U7403 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7104) );
  NOR2_X1 U7404 ( .A1(n7104), .A2(n7101), .ZN(n6323) );
  INV_X1 U7405 ( .A(n6321), .ZN(n6322) );
  AOI21_X1 U7406 ( .B1(n6323), .B2(n6322), .A(REIP_REG_20__SCAN_IN), .ZN(n6326) );
  OAI22_X1 U7407 ( .A1(n6326), .A2(n6325), .B1(n6324), .B2(n6527), .ZN(n6327)
         );
  AOI21_X1 U7408 ( .B1(n6350), .B2(n6503), .A(n6327), .ZN(n6328) );
  OAI211_X1 U7409 ( .C1(n6330), .C2(n6541), .A(n6329), .B(n6328), .ZN(U2807)
         );
  AOI22_X1 U7410 ( .A1(n6331), .A2(n6559), .B1(n6558), .B2(DATAI_30_), .ZN(
        n6333) );
  AOI22_X1 U7411 ( .A1(n6562), .A2(DATAI_14_), .B1(n6561), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7412 ( .A1(n6333), .A2(n6332), .ZN(U2861) );
  AOI22_X1 U7413 ( .A1(n6334), .A2(n6559), .B1(n6558), .B2(DATAI_28_), .ZN(
        n6336) );
  AOI22_X1 U7414 ( .A1(n6562), .A2(DATAI_12_), .B1(n6561), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7415 ( .A1(n6336), .A2(n6335), .ZN(U2863) );
  AOI22_X1 U7416 ( .A1(n6337), .A2(n6559), .B1(n6558), .B2(DATAI_26_), .ZN(
        n6339) );
  AOI22_X1 U7417 ( .A1(n6562), .A2(DATAI_10_), .B1(n6561), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U7418 ( .A1(n6339), .A2(n6338), .ZN(U2865) );
  INV_X1 U7419 ( .A(n6340), .ZN(n6341) );
  AOI22_X1 U7420 ( .A1(n6341), .A2(n6559), .B1(n6558), .B2(DATAI_24_), .ZN(
        n6343) );
  AOI22_X1 U7421 ( .A1(n6562), .A2(DATAI_8_), .B1(n6561), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U7422 ( .A1(n6343), .A2(n6342), .ZN(U2867) );
  INV_X1 U7423 ( .A(n6558), .ZN(n6344) );
  OAI22_X1 U7424 ( .A1(n6346), .A2(n6345), .B1(n6344), .B2(n5757), .ZN(n6347)
         );
  INV_X1 U7425 ( .A(n6347), .ZN(n6349) );
  AOI22_X1 U7426 ( .A1(n6562), .A2(DATAI_6_), .B1(n6561), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U7427 ( .A1(n6349), .A2(n6348), .ZN(U2869) );
  AOI22_X1 U7428 ( .A1(n6350), .A2(n6559), .B1(n6558), .B2(DATAI_20_), .ZN(
        n6352) );
  AOI22_X1 U7429 ( .A1(n6562), .A2(DATAI_4_), .B1(n6561), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U7430 ( .A1(n6352), .A2(n6351), .ZN(U2871) );
  AOI22_X1 U7431 ( .A1(n6353), .A2(n6559), .B1(n6558), .B2(DATAI_19_), .ZN(
        n6355) );
  AOI22_X1 U7432 ( .A1(n6562), .A2(DATAI_3_), .B1(n6561), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U7433 ( .A1(n6355), .A2(n6354), .ZN(U2872) );
  AOI22_X1 U7434 ( .A1(n6803), .A2(REIP_REG_18__SCAN_IN), .B1(n6694), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6361) );
  NOR2_X1 U7435 ( .A1(n6356), .A2(n6374), .ZN(n6357) );
  AOI21_X1 U7436 ( .B1(n6358), .B2(n6374), .A(n6357), .ZN(n6359) );
  XNOR2_X1 U7437 ( .A(n6359), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6378)
         );
  AOI22_X1 U7438 ( .A1(n6378), .A2(n6700), .B1(n6698), .B2(n6552), .ZN(n6360)
         );
  OAI211_X1 U7439 ( .C1(n6704), .C2(n6362), .A(n6361), .B(n6360), .ZN(U2968)
         );
  AOI22_X1 U7440 ( .A1(n6785), .A2(REIP_REG_17__SCAN_IN), .B1(n6694), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6364) );
  INV_X1 U7441 ( .A(n6432), .ZN(n6555) );
  AOI22_X1 U7442 ( .A1(n6555), .A2(n6698), .B1(n6663), .B2(n6430), .ZN(n6363)
         );
  OAI211_X1 U7443 ( .C1(n6365), .C2(n6681), .A(n6364), .B(n6363), .ZN(U2969)
         );
  AOI22_X1 U7444 ( .A1(n6367), .A2(n6801), .B1(n6799), .B2(n6366), .ZN(n6373)
         );
  INV_X1 U7445 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6370) );
  NOR2_X1 U7446 ( .A1(n6774), .A2(n7107), .ZN(n6368) );
  AOI221_X1 U7447 ( .B1(n6371), .B2(n6370), .C1(n6369), .C2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6368), .ZN(n6372) );
  NAND2_X1 U7448 ( .A1(n6373), .A2(n6372), .ZN(U2997) );
  NOR2_X1 U7449 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6374), .ZN(n6376)
         );
  AOI22_X1 U7450 ( .A1(n6803), .A2(REIP_REG_18__SCAN_IN), .B1(n6376), .B2(
        n6375), .ZN(n6380) );
  AOI22_X1 U7451 ( .A1(n6378), .A2(n6801), .B1(n6799), .B2(n6377), .ZN(n6379)
         );
  OAI211_X1 U7452 ( .C1(n6382), .C2(n6381), .A(n6380), .B(n6379), .ZN(U3000)
         );
  OAI21_X1 U7453 ( .B1(n6384), .B2(n6383), .A(n6709), .ZN(n6394) );
  OAI22_X1 U7454 ( .A1(n6386), .A2(n6773), .B1(n6775), .B2(n6385), .ZN(n6387)
         );
  AOI21_X1 U7455 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n6394), .A(n6387), 
        .ZN(n6393) );
  NOR3_X1 U7456 ( .A1(n6390), .A2(n6389), .A3(n6388), .ZN(n6397) );
  OAI221_X1 U7457 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n3732), .C2(n6391), .A(n6397), 
        .ZN(n6392) );
  OAI211_X1 U7458 ( .C1(n7099), .C2(n6774), .A(n6393), .B(n6392), .ZN(U3002)
         );
  INV_X1 U7459 ( .A(n6394), .ZN(n6401) );
  AOI21_X1 U7460 ( .B1(n6396), .B2(n6799), .A(n6395), .ZN(n6400) );
  AOI22_X1 U7461 ( .A1(n6398), .A2(n6801), .B1(n3732), .B2(n6397), .ZN(n6399)
         );
  OAI211_X1 U7462 ( .C1(n6401), .C2(n3732), .A(n6400), .B(n6399), .ZN(U3003)
         );
  INV_X1 U7463 ( .A(n6402), .ZN(n6405) );
  NOR3_X1 U7464 ( .A1(n7147), .A2(n6403), .A3(n3191), .ZN(n6404) );
  NAND2_X1 U7465 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  OAI21_X1 U7466 ( .B1(n7145), .B2(n6407), .A(n6406), .ZN(U3455) );
  INV_X1 U7467 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7072) );
  AOI21_X1 U7468 ( .B1(STATE_REG_1__SCAN_IN), .B2(n7072), .A(n7063), .ZN(n6412) );
  INV_X1 U7469 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6408) );
  AND2_X1 U7470 ( .A1(n7063), .A2(STATE_REG_1__SCAN_IN), .ZN(n7130) );
  AOI21_X1 U7471 ( .B1(n6412), .B2(n6408), .A(n7130), .ZN(U2789) );
  OAI21_X1 U7472 ( .B1(n6409), .B2(n7033), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6410) );
  OAI21_X1 U7473 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7035), .A(n6410), .ZN(
        U2790) );
  INV_X2 U7474 ( .A(n7130), .ZN(n7168) );
  NOR2_X1 U7475 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6413) );
  OAI21_X1 U7476 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6413), .A(n7168), .ZN(n6411)
         );
  OAI21_X1 U7477 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n7168), .A(n6411), .ZN(
        U2791) );
  NOR2_X1 U7478 ( .A1(n7130), .A2(n6412), .ZN(n7135) );
  OAI21_X1 U7479 ( .B1(BS16_N), .B2(n6413), .A(n7135), .ZN(n7133) );
  OAI21_X1 U7480 ( .B1(n7135), .B2(n6414), .A(n7133), .ZN(U2792) );
  OAI21_X1 U7481 ( .B1(n6416), .B2(n6415), .A(n6681), .ZN(U2793) );
  NOR4_X1 U7482 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6426) );
  AOI211_X1 U7483 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_28__SCAN_IN), .B(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6425) );
  NOR4_X1 U7484 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n6417) );
  NAND3_X1 U7485 ( .A1(n6417), .A2(n7046), .A3(n7047), .ZN(n6423) );
  NOR4_X1 U7486 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6421) );
  NOR4_X1 U7487 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6420)
         );
  NOR4_X1 U7488 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6419) );
  NOR4_X1 U7489 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6418) );
  NAND4_X1 U7490 ( .A1(n6421), .A2(n6420), .A3(n6419), .A4(n6418), .ZN(n6422)
         );
  NOR4_X1 U7491 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), 
        .A3(n6423), .A4(n6422), .ZN(n6424) );
  NAND3_X1 U7492 ( .A1(n6426), .A2(n6425), .A3(n6424), .ZN(n7151) );
  INV_X1 U7493 ( .A(n7151), .ZN(n7153) );
  NAND2_X1 U7494 ( .A1(n7153), .A2(n7074), .ZN(n7154) );
  OAI21_X1 U7495 ( .B1(n7153), .B2(BYTEENABLE_REG_1__SCAN_IN), .A(n7154), .ZN(
        n6427) );
  OR4_X1 U7496 ( .A1(n7151), .A2(DATAWIDTH_REG_1__SCAN_IN), .A3(
        REIP_REG_0__SCAN_IN), .A4(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U7497 ( .A1(n6427), .A2(n6428), .ZN(U2794) );
  NAND2_X1 U7498 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n7151), .ZN(n6429) );
  OAI211_X1 U7499 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(n7154), .A(n6429), .B(
        n6428), .ZN(U2795) );
  AOI22_X1 U7500 ( .A1(EBX_REG_17__SCAN_IN), .A2(n6543), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6525), .ZN(n6439) );
  AOI21_X1 U7501 ( .B1(n6518), .B2(n6430), .A(n6524), .ZN(n6438) );
  OAI22_X1 U7502 ( .A1(n6432), .A2(n6515), .B1(n6431), .B2(n6527), .ZN(n6433)
         );
  INV_X1 U7503 ( .A(n6433), .ZN(n6437) );
  OAI21_X1 U7504 ( .B1(REIP_REG_17__SCAN_IN), .B2(n6435), .A(n6434), .ZN(n6436) );
  NAND4_X1 U7505 ( .A1(n6439), .A2(n6438), .A3(n6437), .A4(n6436), .ZN(U2810)
         );
  NOR2_X1 U7506 ( .A1(n6440), .A2(n7092), .ZN(n6456) );
  AOI21_X1 U7507 ( .B1(REIP_REG_13__SCAN_IN), .B2(n6456), .A(
        REIP_REG_14__SCAN_IN), .ZN(n6451) );
  OAI22_X1 U7508 ( .A1(n6442), .A2(n6527), .B1(n6441), .B2(n6522), .ZN(n6443)
         );
  AOI211_X1 U7509 ( .C1(n6525), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6524), 
        .B(n6443), .ZN(n6449) );
  INV_X1 U7510 ( .A(n6444), .ZN(n6445) );
  OAI22_X1 U7511 ( .A1(n6446), .A2(n6515), .B1(n6445), .B2(n6541), .ZN(n6447)
         );
  INV_X1 U7512 ( .A(n6447), .ZN(n6448) );
  OAI211_X1 U7513 ( .C1(n6451), .C2(n6450), .A(n6449), .B(n6448), .ZN(U2813)
         );
  NAND2_X1 U7514 ( .A1(n6452), .A2(n7092), .ZN(n6469) );
  NAND2_X1 U7515 ( .A1(n6465), .A2(n6469), .ZN(n6453) );
  AOI22_X1 U7516 ( .A1(n6454), .A2(n6539), .B1(REIP_REG_13__SCAN_IN), .B2(
        n6453), .ZN(n6463) );
  AOI22_X1 U7517 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6543), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n6525), .ZN(n6462) );
  INV_X1 U7518 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6455) );
  AOI21_X1 U7519 ( .B1(n6456), .B2(n6455), .A(n6524), .ZN(n6461) );
  OAI22_X1 U7520 ( .A1(n6458), .A2(n6515), .B1(n6457), .B2(n6541), .ZN(n6459)
         );
  INV_X1 U7521 ( .A(n6459), .ZN(n6460) );
  NAND4_X1 U7522 ( .A1(n6463), .A2(n6462), .A3(n6461), .A4(n6460), .ZN(U2814)
         );
  OAI22_X1 U7523 ( .A1(n6465), .A2(n7092), .B1(n6464), .B2(n6522), .ZN(n6466)
         );
  AOI211_X1 U7524 ( .C1(n6525), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6524), 
        .B(n6466), .ZN(n6471) );
  AOI22_X1 U7525 ( .A1(n6664), .A2(n6503), .B1(n6518), .B2(n6662), .ZN(n6470)
         );
  NAND2_X1 U7526 ( .A1(n6467), .A2(n6539), .ZN(n6468) );
  NAND4_X1 U7527 ( .A1(n6471), .A2(n6470), .A3(n6469), .A4(n6468), .ZN(U2815)
         );
  NOR3_X1 U7528 ( .A1(n6507), .A2(REIP_REG_10__SCAN_IN), .A3(n6472), .ZN(n6473) );
  AOI211_X1 U7529 ( .C1(n6525), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6524), 
        .B(n6473), .ZN(n6483) );
  INV_X1 U7530 ( .A(n6474), .ZN(n6475) );
  AOI22_X1 U7531 ( .A1(n6475), .A2(n6539), .B1(EBX_REG_10__SCAN_IN), .B2(n6543), .ZN(n6482) );
  INV_X1 U7532 ( .A(n6476), .ZN(n6478) );
  AOI22_X1 U7533 ( .A1(n6478), .A2(n6503), .B1(n6518), .B2(n6477), .ZN(n6481)
         );
  NOR3_X1 U7534 ( .A1(n6507), .A2(REIP_REG_9__SCAN_IN), .A3(n6479), .ZN(n6484)
         );
  OAI21_X1 U7535 ( .B1(n6484), .B2(n6485), .A(REIP_REG_10__SCAN_IN), .ZN(n6480) );
  NAND4_X1 U7536 ( .A1(n6483), .A2(n6482), .A3(n6481), .A4(n6480), .ZN(U2817)
         );
  AOI21_X1 U7537 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6485), .A(n6484), .ZN(n6493)
         );
  NAND2_X1 U7538 ( .A1(n6525), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6486)
         );
  OAI211_X1 U7539 ( .C1(n6717), .C2(n6527), .A(n6511), .B(n6486), .ZN(n6487)
         );
  AOI21_X1 U7540 ( .B1(n6488), .B2(n6503), .A(n6487), .ZN(n6489) );
  INV_X1 U7541 ( .A(n6489), .ZN(n6490) );
  AOI21_X1 U7542 ( .B1(n6491), .B2(n6518), .A(n6490), .ZN(n6492) );
  OAI211_X1 U7543 ( .C1(n6494), .C2(n6522), .A(n6493), .B(n6492), .ZN(U2818)
         );
  INV_X1 U7544 ( .A(n6495), .ZN(n6496) );
  NOR2_X1 U7545 ( .A1(n6496), .A2(REIP_REG_7__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U7546 ( .A1(n6525), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6497)
         );
  NAND2_X1 U7547 ( .A1(n6497), .A2(n6511), .ZN(n6498) );
  AOI21_X1 U7548 ( .B1(n6532), .B2(n6499), .A(n6498), .ZN(n6501) );
  NAND2_X1 U7549 ( .A1(n6543), .A2(EBX_REG_7__SCAN_IN), .ZN(n6500) );
  OAI211_X1 U7550 ( .C1(n6735), .C2(n6527), .A(n6501), .B(n6500), .ZN(n6502)
         );
  AOI21_X1 U7551 ( .B1(n6672), .B2(n6503), .A(n6502), .ZN(n6509) );
  INV_X1 U7552 ( .A(n6506), .ZN(n6505) );
  OAI21_X1 U7553 ( .B1(n6507), .B2(n6505), .A(n6504), .ZN(n6533) );
  NOR3_X1 U7554 ( .A1(n6507), .A2(REIP_REG_6__SCAN_IN), .A3(n6506), .ZN(n6510)
         );
  OAI21_X1 U7555 ( .B1(n6533), .B2(n6510), .A(REIP_REG_7__SCAN_IN), .ZN(n6508)
         );
  OAI211_X1 U7556 ( .C1(n6541), .C2(n6675), .A(n6509), .B(n6508), .ZN(U2820)
         );
  AOI21_X1 U7557 ( .B1(n6533), .B2(REIP_REG_6__SCAN_IN), .A(n6510), .ZN(n6521)
         );
  NAND2_X1 U7558 ( .A1(n6525), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6512)
         );
  OAI211_X1 U7559 ( .C1(n6752), .C2(n6527), .A(n6512), .B(n6511), .ZN(n6513)
         );
  INV_X1 U7560 ( .A(n6513), .ZN(n6514) );
  OAI21_X1 U7561 ( .B1(n6516), .B2(n6515), .A(n6514), .ZN(n6517) );
  AOI21_X1 U7562 ( .B1(n6519), .B2(n6518), .A(n6517), .ZN(n6520) );
  OAI211_X1 U7563 ( .C1(n6523), .C2(n6522), .A(n6521), .B(n6520), .ZN(U2821)
         );
  AOI21_X1 U7564 ( .B1(n6525), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6524), 
        .ZN(n6526) );
  OAI21_X1 U7565 ( .B1(n6527), .B2(n6765), .A(n6526), .ZN(n6530) );
  NOR2_X1 U7566 ( .A1(n6680), .A2(n6528), .ZN(n6529) );
  AOI211_X1 U7567 ( .C1(n6543), .C2(EBX_REG_5__SCAN_IN), .A(n6530), .B(n6529), 
        .ZN(n6536) );
  AND2_X1 U7568 ( .A1(n6532), .A2(n6531), .ZN(n6534) );
  OAI21_X1 U7569 ( .B1(n6534), .B2(REIP_REG_5__SCAN_IN), .A(n6533), .ZN(n6535)
         );
  OAI211_X1 U7570 ( .C1(n6541), .C2(n6685), .A(n6536), .B(n6535), .ZN(U2822)
         );
  INV_X1 U7571 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7077) );
  OR2_X1 U7572 ( .A1(n6538), .A2(n6537), .ZN(n6550) );
  AOI22_X1 U7573 ( .A1(n6525), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6539), 
        .B2(n6786), .ZN(n6540) );
  OAI21_X1 U7574 ( .B1(n6541), .B2(n6693), .A(n6540), .ZN(n6542) );
  AOI21_X1 U7575 ( .B1(n6543), .B2(EBX_REG_3__SCAN_IN), .A(n6542), .ZN(n6544)
         );
  OAI21_X1 U7576 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(n6547) );
  AOI21_X1 U7577 ( .B1(n6690), .B2(n6548), .A(n6547), .ZN(n6549) );
  OAI221_X1 U7578 ( .B1(n6551), .B2(n7077), .C1(n6551), .C2(n6550), .A(n6549), 
        .ZN(U2824) );
  AOI22_X1 U7579 ( .A1(n6552), .A2(n6559), .B1(n6558), .B2(DATAI_18_), .ZN(
        n6554) );
  AOI22_X1 U7580 ( .A1(n6562), .A2(DATAI_2_), .B1(n6561), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U7581 ( .A1(n6554), .A2(n6553), .ZN(U2873) );
  AOI22_X1 U7582 ( .A1(n6555), .A2(n6559), .B1(n6558), .B2(DATAI_17_), .ZN(
        n6557) );
  AOI22_X1 U7583 ( .A1(n6562), .A2(DATAI_1_), .B1(n6561), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U7584 ( .A1(n6557), .A2(n6556), .ZN(U2874) );
  AOI22_X1 U7585 ( .A1(n6560), .A2(n6559), .B1(n6558), .B2(DATAI_16_), .ZN(
        n6564) );
  AOI22_X1 U7586 ( .A1(n6562), .A2(DATAI_0_), .B1(n6561), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U7587 ( .A1(n6564), .A2(n6563), .ZN(U2875) );
  INV_X1 U7588 ( .A(n6565), .ZN(n6568) );
  AOI22_X1 U7589 ( .A1(n6594), .A2(DATAO_REG_30__SCAN_IN), .B1(n6568), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6566) );
  OAI21_X1 U7590 ( .B1(n6567), .B2(n6570), .A(n6566), .ZN(U2893) );
  AOI22_X1 U7591 ( .A1(n6594), .A2(DATAO_REG_17__SCAN_IN), .B1(n6568), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6569) );
  OAI21_X1 U7592 ( .B1(n6571), .B2(n6570), .A(n6569), .ZN(U2906) );
  INV_X1 U7593 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6661) );
  AOI22_X1 U7594 ( .A1(n7160), .A2(LWORD_REG_15__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6572) );
  OAI21_X1 U7595 ( .B1(n6661), .B2(n6596), .A(n6572), .ZN(U2908) );
  AOI222_X1 U7596 ( .A1(n6578), .A2(LWORD_REG_14__SCAN_IN), .B1(n6590), .B2(
        EAX_REG_14__SCAN_IN), .C1(DATAO_REG_14__SCAN_IN), .C2(n6594), .ZN(
        n6573) );
  INV_X1 U7597 ( .A(n6573), .ZN(U2909) );
  AOI22_X1 U7598 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6578), .B1(n6594), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6574) );
  OAI21_X1 U7599 ( .B1(n6575), .B2(n6596), .A(n6574), .ZN(U2910) );
  INV_X1 U7600 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6650) );
  AOI22_X1 U7601 ( .A1(n7160), .A2(LWORD_REG_12__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6576) );
  OAI21_X1 U7602 ( .B1(n6650), .B2(n6596), .A(n6576), .ZN(U2911) );
  INV_X1 U7603 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6646) );
  AOI22_X1 U7604 ( .A1(n7160), .A2(LWORD_REG_11__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6577) );
  OAI21_X1 U7605 ( .B1(n6646), .B2(n6596), .A(n6577), .ZN(U2912) );
  AOI222_X1 U7606 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6578), .B1(n6590), .B2(
        EAX_REG_10__SCAN_IN), .C1(n6594), .C2(DATAO_REG_10__SCAN_IN), .ZN(
        n6579) );
  INV_X1 U7607 ( .A(n6579), .ZN(U2913) );
  INV_X1 U7608 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U7609 ( .A1(n7160), .A2(LWORD_REG_9__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6580) );
  OAI21_X1 U7610 ( .B1(n6641), .B2(n6596), .A(n6580), .ZN(U2914) );
  AOI22_X1 U7611 ( .A1(n7160), .A2(LWORD_REG_8__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6581) );
  OAI21_X1 U7612 ( .B1(n6582), .B2(n6596), .A(n6581), .ZN(U2915) );
  AOI22_X1 U7613 ( .A1(n7160), .A2(LWORD_REG_7__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6583) );
  OAI21_X1 U7614 ( .B1(n4416), .B2(n6596), .A(n6583), .ZN(U2916) );
  AOI22_X1 U7615 ( .A1(n7160), .A2(LWORD_REG_6__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6584) );
  OAI21_X1 U7616 ( .B1(n4322), .B2(n6596), .A(n6584), .ZN(U2917) );
  AOI22_X1 U7617 ( .A1(n7160), .A2(LWORD_REG_5__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6585) );
  OAI21_X1 U7618 ( .B1(n4240), .B2(n6596), .A(n6585), .ZN(U2918) );
  AOI22_X1 U7619 ( .A1(n7160), .A2(LWORD_REG_4__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6586) );
  OAI21_X1 U7620 ( .B1(n6587), .B2(n6596), .A(n6586), .ZN(U2919) );
  AOI22_X1 U7621 ( .A1(n7160), .A2(LWORD_REG_3__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6588) );
  OAI21_X1 U7622 ( .B1(n6589), .B2(n6596), .A(n6588), .ZN(U2920) );
  AOI222_X1 U7623 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n7160), .B1(n6590), .B2(
        EAX_REG_2__SCAN_IN), .C1(n6594), .C2(DATAO_REG_2__SCAN_IN), .ZN(n6591)
         );
  INV_X1 U7624 ( .A(n6591), .ZN(U2921) );
  AOI22_X1 U7625 ( .A1(n7160), .A2(LWORD_REG_1__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6592) );
  OAI21_X1 U7626 ( .B1(n6593), .B2(n6596), .A(n6592), .ZN(U2922) );
  AOI22_X1 U7627 ( .A1(n7160), .A2(LWORD_REG_0__SCAN_IN), .B1(n6594), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6595) );
  OAI21_X1 U7628 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(U2923) );
  INV_X1 U7629 ( .A(n6598), .ZN(n6599) );
  OAI21_X1 U7630 ( .B1(n3596), .B2(n4043), .A(n6599), .ZN(n6648) );
  AOI22_X1 U7631 ( .A1(n6658), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6653), .ZN(n6600) );
  OAI21_X1 U7632 ( .B1(n6622), .B2(n6656), .A(n6600), .ZN(U2924) );
  AOI22_X1 U7633 ( .A1(n6658), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6653), .ZN(n6601) );
  OAI21_X1 U7634 ( .B1(n6624), .B2(n6656), .A(n6601), .ZN(U2925) );
  AOI22_X1 U7635 ( .A1(n6658), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6653), .ZN(n6602) );
  OAI21_X1 U7636 ( .B1(n6626), .B2(n6656), .A(n6602), .ZN(U2926) );
  AOI22_X1 U7637 ( .A1(n6658), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6653), .ZN(n6603) );
  OAI21_X1 U7638 ( .B1(n6656), .B2(n6628), .A(n6603), .ZN(U2927) );
  AOI22_X1 U7639 ( .A1(n6658), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6653), .ZN(n6604) );
  OAI21_X1 U7640 ( .B1(n6656), .B2(n6630), .A(n6604), .ZN(U2928) );
  AOI22_X1 U7641 ( .A1(n6658), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6653), .ZN(n6605) );
  OAI21_X1 U7642 ( .B1(n6656), .B2(n6632), .A(n6605), .ZN(U2929) );
  AOI22_X1 U7643 ( .A1(n6658), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6653), .ZN(n6606) );
  OAI21_X1 U7644 ( .B1(n6656), .B2(n6634), .A(n6606), .ZN(U2930) );
  AOI22_X1 U7645 ( .A1(n6658), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6653), .ZN(n6607) );
  OAI21_X1 U7646 ( .B1(n6656), .B2(n6636), .A(n6607), .ZN(U2931) );
  AOI22_X1 U7647 ( .A1(n6658), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6653), .ZN(n6608) );
  OAI21_X1 U7648 ( .B1(n6638), .B2(n6656), .A(n6608), .ZN(U2932) );
  INV_X1 U7649 ( .A(DATAI_9_), .ZN(n6609) );
  NOR2_X1 U7650 ( .A1(n6656), .A2(n6609), .ZN(n6639) );
  AOI21_X1 U7651 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6648), .A(n6639), .ZN(n6610) );
  OAI21_X1 U7652 ( .B1(n6611), .B2(n6660), .A(n6610), .ZN(U2933) );
  AOI22_X1 U7653 ( .A1(n6658), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n6653), .ZN(n6612) );
  OAI21_X1 U7654 ( .B1(n6656), .B2(n6643), .A(n6612), .ZN(U2934) );
  INV_X1 U7655 ( .A(DATAI_11_), .ZN(n6613) );
  NOR2_X1 U7656 ( .A1(n6656), .A2(n6613), .ZN(n6644) );
  AOI21_X1 U7657 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6658), .A(n6644), .ZN(
        n6614) );
  OAI21_X1 U7658 ( .B1(n6615), .B2(n6660), .A(n6614), .ZN(U2935) );
  INV_X1 U7659 ( .A(DATAI_12_), .ZN(n6616) );
  NOR2_X1 U7660 ( .A1(n6656), .A2(n6616), .ZN(n6647) );
  AOI21_X1 U7661 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6648), .A(n6647), .ZN(
        n6617) );
  OAI21_X1 U7662 ( .B1(n6618), .B2(n6660), .A(n6617), .ZN(U2936) );
  AOI22_X1 U7663 ( .A1(n6658), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6653), .ZN(n6619) );
  OAI21_X1 U7664 ( .B1(n6652), .B2(n6656), .A(n6619), .ZN(U2937) );
  AOI22_X1 U7665 ( .A1(n6658), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n6653), .ZN(n6620) );
  OAI21_X1 U7666 ( .B1(n6655), .B2(n6656), .A(n6620), .ZN(U2938) );
  AOI22_X1 U7667 ( .A1(n6658), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6653), .ZN(n6621) );
  OAI21_X1 U7668 ( .B1(n6622), .B2(n6656), .A(n6621), .ZN(U2939) );
  AOI22_X1 U7669 ( .A1(n6658), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6653), .ZN(n6623) );
  OAI21_X1 U7670 ( .B1(n6624), .B2(n6656), .A(n6623), .ZN(U2940) );
  AOI22_X1 U7671 ( .A1(n6658), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6653), .ZN(n6625) );
  OAI21_X1 U7672 ( .B1(n6626), .B2(n6656), .A(n6625), .ZN(U2941) );
  AOI22_X1 U7673 ( .A1(n6658), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6653), .ZN(n6627) );
  OAI21_X1 U7674 ( .B1(n6656), .B2(n6628), .A(n6627), .ZN(U2942) );
  AOI22_X1 U7675 ( .A1(n6658), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6653), .ZN(n6629) );
  OAI21_X1 U7676 ( .B1(n6656), .B2(n6630), .A(n6629), .ZN(U2943) );
  AOI22_X1 U7677 ( .A1(n6658), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6653), .ZN(n6631) );
  OAI21_X1 U7678 ( .B1(n6656), .B2(n6632), .A(n6631), .ZN(U2944) );
  AOI22_X1 U7679 ( .A1(n6658), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6653), .ZN(n6633) );
  OAI21_X1 U7680 ( .B1(n6656), .B2(n6634), .A(n6633), .ZN(U2945) );
  AOI22_X1 U7681 ( .A1(n6658), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6653), .ZN(n6635) );
  OAI21_X1 U7682 ( .B1(n6656), .B2(n6636), .A(n6635), .ZN(U2946) );
  AOI22_X1 U7683 ( .A1(n6658), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6653), .ZN(n6637) );
  OAI21_X1 U7684 ( .B1(n6638), .B2(n6656), .A(n6637), .ZN(U2947) );
  AOI21_X1 U7685 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6648), .A(n6639), .ZN(n6640) );
  OAI21_X1 U7686 ( .B1(n6641), .B2(n6660), .A(n6640), .ZN(U2948) );
  AOI22_X1 U7687 ( .A1(n6658), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6653), .ZN(n6642) );
  OAI21_X1 U7688 ( .B1(n6656), .B2(n6643), .A(n6642), .ZN(U2949) );
  AOI21_X1 U7689 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6648), .A(n6644), .ZN(
        n6645) );
  OAI21_X1 U7690 ( .B1(n6646), .B2(n6660), .A(n6645), .ZN(U2950) );
  AOI21_X1 U7691 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6648), .A(n6647), .ZN(
        n6649) );
  OAI21_X1 U7692 ( .B1(n6650), .B2(n6660), .A(n6649), .ZN(U2951) );
  AOI22_X1 U7693 ( .A1(n6658), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6653), .ZN(n6651) );
  OAI21_X1 U7694 ( .B1(n6652), .B2(n6656), .A(n6651), .ZN(U2952) );
  AOI22_X1 U7695 ( .A1(n6658), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6653), .ZN(n6654) );
  OAI21_X1 U7696 ( .B1(n6655), .B2(n6656), .A(n6654), .ZN(U2953) );
  INV_X1 U7697 ( .A(n6656), .ZN(n6657) );
  AOI22_X1 U7698 ( .A1(n6658), .A2(LWORD_REG_15__SCAN_IN), .B1(n6657), .B2(
        DATAI_15_), .ZN(n6659) );
  OAI21_X1 U7699 ( .B1(n6661), .B2(n6660), .A(n6659), .ZN(U2954) );
  AOI22_X1 U7700 ( .A1(n6803), .A2(REIP_REG_12__SCAN_IN), .B1(n6694), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6666) );
  AOI22_X1 U7701 ( .A1(n6664), .A2(n6698), .B1(n6663), .B2(n6662), .ZN(n6665)
         );
  OAI211_X1 U7702 ( .C1(n6667), .C2(n6681), .A(n6666), .B(n6665), .ZN(U2974)
         );
  AOI22_X1 U7703 ( .A1(n6803), .A2(REIP_REG_7__SCAN_IN), .B1(n6694), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6674) );
  OAI21_X1 U7704 ( .B1(n6668), .B2(n6670), .A(n6669), .ZN(n6671) );
  INV_X1 U7705 ( .A(n6671), .ZN(n6737) );
  AOI22_X1 U7706 ( .A1(n6737), .A2(n6700), .B1(n6698), .B2(n6672), .ZN(n6673)
         );
  OAI211_X1 U7707 ( .C1(n6704), .C2(n6675), .A(n6674), .B(n6673), .ZN(U2979)
         );
  AOI22_X1 U7708 ( .A1(n6803), .A2(REIP_REG_5__SCAN_IN), .B1(n6694), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6684) );
  OAI21_X1 U7709 ( .B1(n3192), .B2(n6677), .A(n6676), .ZN(n6766) );
  OAI22_X1 U7710 ( .A1(n6766), .A2(n6681), .B1(n6680), .B2(n6679), .ZN(n6682)
         );
  INV_X1 U7711 ( .A(n6682), .ZN(n6683) );
  OAI211_X1 U7712 ( .C1(n6704), .C2(n6685), .A(n6684), .B(n6683), .ZN(U2981)
         );
  AOI22_X1 U7713 ( .A1(n6803), .A2(REIP_REG_3__SCAN_IN), .B1(n6694), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U7714 ( .A1(n6686), .A2(n6687), .ZN(n6688) );
  AND2_X1 U7715 ( .A1(n6689), .A2(n6688), .ZN(n6787) );
  AOI22_X1 U7716 ( .A1(n6690), .A2(n6698), .B1(n6700), .B2(n6787), .ZN(n6691)
         );
  OAI211_X1 U7717 ( .C1(n6704), .C2(n6693), .A(n6692), .B(n6691), .ZN(U2983)
         );
  AOI22_X1 U7718 ( .A1(n6803), .A2(REIP_REG_2__SCAN_IN), .B1(n6694), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6702) );
  XOR2_X1 U7719 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .B(n6695), .Z(n6696) );
  XNOR2_X1 U7720 ( .A(n6697), .B(n6696), .ZN(n6802) );
  AOI22_X1 U7721 ( .A1(n6802), .A2(n6700), .B1(n6699), .B2(n6698), .ZN(n6701)
         );
  OAI211_X1 U7722 ( .C1(n6704), .C2(n6703), .A(n6702), .B(n6701), .ZN(U2984)
         );
  INV_X1 U7723 ( .A(n6705), .ZN(n6706) );
  AOI21_X1 U7724 ( .B1(n6707), .B2(n6799), .A(n6706), .ZN(n6714) );
  INV_X1 U7725 ( .A(n6708), .ZN(n6711) );
  INV_X1 U7726 ( .A(n6709), .ZN(n6710) );
  AOI22_X1 U7727 ( .A1(n6711), .A2(n6801), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6710), .ZN(n6713) );
  NAND3_X1 U7728 ( .A1(n6714), .A2(n6713), .A3(n6712), .ZN(U3007) );
  INV_X1 U7729 ( .A(n6715), .ZN(n6725) );
  OAI21_X1 U7730 ( .B1(n6717), .B2(n6775), .A(n6716), .ZN(n6718) );
  INV_X1 U7731 ( .A(n6718), .ZN(n6723) );
  INV_X1 U7732 ( .A(n6719), .ZN(n6721) );
  AOI22_X1 U7733 ( .A1(n6721), .A2(n6801), .B1(n6720), .B2(n6724), .ZN(n6722)
         );
  OAI211_X1 U7734 ( .C1(n6725), .C2(n6724), .A(n6723), .B(n6722), .ZN(U3009)
         );
  AOI211_X1 U7735 ( .C1(n6741), .C2(n6734), .A(n6727), .B(n6726), .ZN(n6732)
         );
  NOR2_X1 U7736 ( .A1(n6728), .A2(n6773), .ZN(n6731) );
  OAI22_X1 U7737 ( .A1(n6729), .A2(n6775), .B1(n7085), .B2(n6774), .ZN(n6730)
         );
  NOR3_X1 U7738 ( .A1(n6732), .A2(n6731), .A3(n6730), .ZN(n6733) );
  OAI21_X1 U7739 ( .B1(n6742), .B2(n6734), .A(n6733), .ZN(U3010) );
  INV_X1 U7740 ( .A(n6735), .ZN(n6736) );
  AOI22_X1 U7741 ( .A1(n6736), .A2(n6799), .B1(n6785), .B2(REIP_REG_7__SCAN_IN), .ZN(n6740) );
  AOI22_X1 U7742 ( .A1(n6738), .A2(n6741), .B1(n6737), .B2(n6801), .ZN(n6739)
         );
  OAI211_X1 U7743 ( .C1(n6742), .C2(n6741), .A(n6740), .B(n6739), .ZN(U3011)
         );
  INV_X1 U7744 ( .A(n6743), .ZN(n6748) );
  INV_X1 U7745 ( .A(n6744), .ZN(n6747) );
  OAI22_X1 U7746 ( .A1(n6748), .A2(n6747), .B1(n6746), .B2(n6745), .ZN(n6800)
         );
  AOI221_X1 U7747 ( .B1(n6751), .B2(n6750), .C1(n6749), .C2(n6750), .A(n6800), 
        .ZN(n6771) );
  INV_X1 U7748 ( .A(n6752), .ZN(n6755) );
  INV_X1 U7749 ( .A(n6753), .ZN(n6754) );
  AOI21_X1 U7750 ( .B1(n6755), .B2(n6799), .A(n6754), .ZN(n6760) );
  INV_X1 U7751 ( .A(n6756), .ZN(n6757) );
  AOI22_X1 U7752 ( .A1(n6758), .A2(n6761), .B1(n6757), .B2(n6801), .ZN(n6759)
         );
  OAI211_X1 U7753 ( .C1(n6771), .C2(n6761), .A(n6760), .B(n6759), .ZN(U3012)
         );
  AOI211_X1 U7754 ( .C1(n6764), .C2(n6763), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .B(n6762), .ZN(n6770) );
  OAI22_X1 U7755 ( .A1(n6766), .A2(n6773), .B1(n6775), .B2(n6765), .ZN(n6767)
         );
  INV_X1 U7756 ( .A(n6767), .ZN(n6769) );
  NAND2_X1 U7757 ( .A1(n6803), .A2(REIP_REG_5__SCAN_IN), .ZN(n6768) );
  OAI211_X1 U7758 ( .C1(n6771), .C2(n6770), .A(n6769), .B(n6768), .ZN(U3013)
         );
  NOR2_X1 U7759 ( .A1(n6795), .A2(n6778), .ZN(n6796) );
  NOR2_X1 U7760 ( .A1(n6796), .A2(n6800), .ZN(n6792) );
  OAI222_X1 U7761 ( .A1(n6776), .A2(n6775), .B1(n6774), .B2(n7079), .C1(n6773), 
        .C2(n6772), .ZN(n6777) );
  INV_X1 U7762 ( .A(n6777), .ZN(n6783) );
  INV_X1 U7763 ( .A(n6778), .ZN(n6780) );
  NOR2_X1 U7764 ( .A1(n6780), .A2(n6779), .ZN(n6788) );
  OAI211_X1 U7765 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6788), .B(n6781), .ZN(n6782) );
  OAI211_X1 U7766 ( .C1(n6792), .C2(n6784), .A(n6783), .B(n6782), .ZN(U3014)
         );
  AOI22_X1 U7767 ( .A1(n6799), .A2(n6786), .B1(n6785), .B2(REIP_REG_3__SCAN_IN), .ZN(n6790) );
  AOI22_X1 U7768 ( .A1(n6788), .A2(n6791), .B1(n6787), .B2(n6801), .ZN(n6789)
         );
  OAI211_X1 U7769 ( .C1(n6792), .C2(n6791), .A(n6790), .B(n6789), .ZN(U3015)
         );
  NOR3_X1 U7770 ( .A1(n6795), .A2(n6794), .A3(n6793), .ZN(n6797) );
  AOI211_X1 U7771 ( .C1(n6799), .C2(n6798), .A(n6797), .B(n6796), .ZN(n6809)
         );
  AOI22_X1 U7772 ( .A1(n6802), .A2(n6801), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6800), .ZN(n6808) );
  NAND2_X1 U7773 ( .A1(n6803), .A2(REIP_REG_2__SCAN_IN), .ZN(n6807) );
  OR3_X1 U7774 ( .A1(n6805), .A2(n6804), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6806) );
  NAND4_X1 U7775 ( .A1(n6809), .A2(n6808), .A3(n6807), .A4(n6806), .ZN(U3016)
         );
  NOR2_X1 U7776 ( .A1(n7014), .A2(n6810), .ZN(U3019) );
  INV_X1 U7777 ( .A(n6811), .ZN(n6821) );
  INV_X1 U7778 ( .A(n6812), .ZN(n6813) );
  NOR2_X1 U7779 ( .A1(n7000), .A2(n6819), .ZN(n6845) );
  AOI21_X1 U7780 ( .B1(n6813), .B2(n6995), .A(n6845), .ZN(n6820) );
  INV_X1 U7781 ( .A(n6820), .ZN(n6815) );
  OAI21_X1 U7782 ( .B1(n6821), .B2(n6815), .A(n6814), .ZN(n6816) );
  AOI21_X1 U7783 ( .B1(n6927), .B2(n6819), .A(n6816), .ZN(n6851) );
  OR2_X1 U7784 ( .A1(n6818), .A2(n6817), .ZN(n6856) );
  AOI22_X1 U7785 ( .A1(n6920), .A2(n6845), .B1(n6919), .B2(n6888), .ZN(n6824)
         );
  OAI22_X1 U7786 ( .A1(n6821), .A2(n6820), .B1(n6819), .B2(n6930), .ZN(n6847)
         );
  AOI22_X1 U7787 ( .A1(n6847), .A2(n6934), .B1(n6864), .B2(n6846), .ZN(n6823)
         );
  OAI211_X1 U7788 ( .C1(n6851), .C2(n6825), .A(n6824), .B(n6823), .ZN(U3060)
         );
  AOI22_X1 U7789 ( .A1(n6939), .A2(n6845), .B1(n6938), .B2(n6888), .ZN(n6827)
         );
  AOI22_X1 U7790 ( .A1(n6847), .A2(n6940), .B1(n6868), .B2(n6846), .ZN(n6826)
         );
  OAI211_X1 U7791 ( .C1(n6851), .C2(n6828), .A(n6827), .B(n6826), .ZN(U3061)
         );
  INV_X1 U7792 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6831) );
  AOI22_X1 U7793 ( .A1(n6945), .A2(n6845), .B1(n6944), .B2(n6888), .ZN(n6830)
         );
  AOI22_X1 U7794 ( .A1(n6847), .A2(n6946), .B1(n6872), .B2(n6846), .ZN(n6829)
         );
  OAI211_X1 U7795 ( .C1(n6851), .C2(n6831), .A(n6830), .B(n6829), .ZN(U3062)
         );
  AOI22_X1 U7796 ( .A1(n6951), .A2(n6845), .B1(n6901), .B2(n6888), .ZN(n6833)
         );
  AOI22_X1 U7797 ( .A1(n6847), .A2(n6952), .B1(n6950), .B2(n6846), .ZN(n6832)
         );
  OAI211_X1 U7798 ( .C1(n6851), .C2(n6834), .A(n6833), .B(n6832), .ZN(U3063)
         );
  AOI22_X1 U7799 ( .A1(n6957), .A2(n6845), .B1(n6905), .B2(n6888), .ZN(n6836)
         );
  AOI22_X1 U7800 ( .A1(n6847), .A2(n6958), .B1(n6956), .B2(n6846), .ZN(n6835)
         );
  OAI211_X1 U7801 ( .C1(n6851), .C2(n6837), .A(n6836), .B(n6835), .ZN(U3064)
         );
  AOI22_X1 U7802 ( .A1(n6963), .A2(n6845), .B1(n6962), .B2(n6888), .ZN(n6839)
         );
  AOI22_X1 U7803 ( .A1(n6847), .A2(n6964), .B1(n6880), .B2(n6846), .ZN(n6838)
         );
  OAI211_X1 U7804 ( .C1(n6851), .C2(n6840), .A(n6839), .B(n6838), .ZN(U3065)
         );
  INV_X1 U7805 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6844) );
  AOI22_X1 U7806 ( .A1(n6970), .A2(n6845), .B1(n6841), .B2(n6888), .ZN(n6843)
         );
  AOI22_X1 U7807 ( .A1(n6847), .A2(n6971), .B1(n6968), .B2(n6846), .ZN(n6842)
         );
  OAI211_X1 U7808 ( .C1(n6851), .C2(n6844), .A(n6843), .B(n6842), .ZN(U3066)
         );
  INV_X1 U7809 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6850) );
  AOI22_X1 U7810 ( .A1(n6979), .A2(n6845), .B1(n6977), .B2(n6888), .ZN(n6849)
         );
  AOI22_X1 U7811 ( .A1(n6847), .A2(n6981), .B1(n6889), .B2(n6846), .ZN(n6848)
         );
  OAI211_X1 U7812 ( .C1(n6851), .C2(n6850), .A(n6849), .B(n6848), .ZN(U3067)
         );
  OAI22_X1 U7813 ( .A1(n6854), .A2(n4173), .B1(n6853), .B2(n6852), .ZN(n6887)
         );
  AND2_X1 U7814 ( .A1(n7000), .A2(n6855), .ZN(n6886) );
  AOI22_X1 U7815 ( .A1(n6934), .A2(n6887), .B1(n6920), .B2(n6886), .ZN(n6866)
         );
  NAND3_X1 U7816 ( .A1(n6856), .A2(n6923), .A3(n6917), .ZN(n6859) );
  AOI21_X1 U7817 ( .B1(n6859), .B2(n6858), .A(n6857), .ZN(n6862) );
  OAI211_X1 U7818 ( .C1(n3454), .C2(n6886), .A(n6860), .B(n7016), .ZN(n6861)
         );
  AOI22_X1 U7819 ( .A1(n6890), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6864), 
        .B2(n6888), .ZN(n6865) );
  OAI211_X1 U7820 ( .C1(n6867), .C2(n6917), .A(n6866), .B(n6865), .ZN(U3068)
         );
  AOI22_X1 U7821 ( .A1(n6940), .A2(n6887), .B1(n6939), .B2(n6886), .ZN(n6870)
         );
  AOI22_X1 U7822 ( .A1(n6890), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6868), 
        .B2(n6888), .ZN(n6869) );
  OAI211_X1 U7823 ( .C1(n6871), .C2(n6917), .A(n6870), .B(n6869), .ZN(U3069)
         );
  AOI22_X1 U7824 ( .A1(n6946), .A2(n6887), .B1(n6945), .B2(n6886), .ZN(n6874)
         );
  AOI22_X1 U7825 ( .A1(n6890), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6872), 
        .B2(n6888), .ZN(n6873) );
  OAI211_X1 U7826 ( .C1(n6875), .C2(n6917), .A(n6874), .B(n6873), .ZN(U3070)
         );
  AOI22_X1 U7827 ( .A1(n6952), .A2(n6887), .B1(n6951), .B2(n6886), .ZN(n6877)
         );
  AOI22_X1 U7828 ( .A1(n6890), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6950), 
        .B2(n6888), .ZN(n6876) );
  OAI211_X1 U7829 ( .C1(n6955), .C2(n6917), .A(n6877), .B(n6876), .ZN(U3071)
         );
  AOI22_X1 U7830 ( .A1(n6958), .A2(n6887), .B1(n6957), .B2(n6886), .ZN(n6879)
         );
  AOI22_X1 U7831 ( .A1(n6890), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6956), 
        .B2(n6888), .ZN(n6878) );
  OAI211_X1 U7832 ( .C1(n6961), .C2(n6917), .A(n6879), .B(n6878), .ZN(U3072)
         );
  AOI22_X1 U7833 ( .A1(n6964), .A2(n6887), .B1(n6963), .B2(n6886), .ZN(n6882)
         );
  AOI22_X1 U7834 ( .A1(n6890), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6880), 
        .B2(n6888), .ZN(n6881) );
  OAI211_X1 U7835 ( .C1(n6883), .C2(n6917), .A(n6882), .B(n6881), .ZN(U3073)
         );
  AOI22_X1 U7836 ( .A1(n6971), .A2(n6887), .B1(n6970), .B2(n6886), .ZN(n6885)
         );
  AOI22_X1 U7837 ( .A1(n6890), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6968), 
        .B2(n6888), .ZN(n6884) );
  OAI211_X1 U7838 ( .C1(n6975), .C2(n6917), .A(n6885), .B(n6884), .ZN(U3074)
         );
  AOI22_X1 U7839 ( .A1(n6981), .A2(n6887), .B1(n6979), .B2(n6886), .ZN(n6892)
         );
  AOI22_X1 U7840 ( .A1(n6890), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6889), 
        .B2(n6888), .ZN(n6891) );
  OAI211_X1 U7841 ( .C1(n6893), .C2(n6917), .A(n6892), .B(n6891), .ZN(U3075)
         );
  INV_X1 U7842 ( .A(n6894), .ZN(n6911) );
  AOI22_X1 U7843 ( .A1(n6920), .A2(n6912), .B1(n6919), .B2(n6911), .ZN(n6896)
         );
  AOI22_X1 U7844 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6914), .B1(n6934), 
        .B2(n6913), .ZN(n6895) );
  OAI211_X1 U7845 ( .C1(n6937), .C2(n6917), .A(n6896), .B(n6895), .ZN(U3076)
         );
  AOI22_X1 U7846 ( .A1(n6939), .A2(n6912), .B1(n6938), .B2(n6911), .ZN(n6898)
         );
  AOI22_X1 U7847 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6914), .B1(n6940), 
        .B2(n6913), .ZN(n6897) );
  OAI211_X1 U7848 ( .C1(n6943), .C2(n6917), .A(n6898), .B(n6897), .ZN(U3077)
         );
  AOI22_X1 U7849 ( .A1(n6945), .A2(n6912), .B1(n6944), .B2(n6911), .ZN(n6900)
         );
  AOI22_X1 U7850 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6914), .B1(n6946), 
        .B2(n6913), .ZN(n6899) );
  OAI211_X1 U7851 ( .C1(n6949), .C2(n6917), .A(n6900), .B(n6899), .ZN(U3078)
         );
  AOI22_X1 U7852 ( .A1(n6951), .A2(n6912), .B1(n6901), .B2(n6911), .ZN(n6903)
         );
  AOI22_X1 U7853 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6914), .B1(n6952), 
        .B2(n6913), .ZN(n6902) );
  OAI211_X1 U7854 ( .C1(n6904), .C2(n6917), .A(n6903), .B(n6902), .ZN(U3079)
         );
  AOI22_X1 U7855 ( .A1(n6957), .A2(n6912), .B1(n6905), .B2(n6911), .ZN(n6907)
         );
  AOI22_X1 U7856 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6914), .B1(n6958), 
        .B2(n6913), .ZN(n6906) );
  OAI211_X1 U7857 ( .C1(n6908), .C2(n6917), .A(n6907), .B(n6906), .ZN(U3080)
         );
  AOI22_X1 U7858 ( .A1(n6963), .A2(n6912), .B1(n6962), .B2(n6911), .ZN(n6910)
         );
  AOI22_X1 U7859 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6914), .B1(n6964), 
        .B2(n6913), .ZN(n6909) );
  OAI211_X1 U7860 ( .C1(n6967), .C2(n6917), .A(n6910), .B(n6909), .ZN(U3081)
         );
  AOI22_X1 U7861 ( .A1(n6979), .A2(n6912), .B1(n6977), .B2(n6911), .ZN(n6916)
         );
  AOI22_X1 U7862 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6914), .B1(n6981), 
        .B2(n6913), .ZN(n6915) );
  OAI211_X1 U7863 ( .C1(n6986), .C2(n6917), .A(n6916), .B(n6915), .ZN(U3083)
         );
  NOR2_X1 U7864 ( .A1(n6918), .A2(n7016), .ZN(n6978) );
  AOI22_X1 U7865 ( .A1(n6920), .A2(n6978), .B1(n6919), .B2(n6976), .ZN(n6936)
         );
  INV_X1 U7866 ( .A(n6921), .ZN(n6922) );
  AOI21_X1 U7867 ( .B1(n6924), .B2(n6923), .A(n6922), .ZN(n6933) );
  AOI21_X1 U7868 ( .B1(n6925), .B2(n6995), .A(n6978), .ZN(n6932) );
  INV_X1 U7869 ( .A(n6932), .ZN(n6929) );
  AOI21_X1 U7870 ( .B1(n6927), .B2(n6931), .A(n6926), .ZN(n6928) );
  OAI21_X1 U7871 ( .B1(n6933), .B2(n6929), .A(n6928), .ZN(n6982) );
  OAI22_X1 U7872 ( .A1(n6933), .A2(n6932), .B1(n6931), .B2(n6930), .ZN(n6980)
         );
  AOI22_X1 U7873 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6982), .B1(n6934), 
        .B2(n6980), .ZN(n6935) );
  OAI211_X1 U7874 ( .C1(n6937), .C2(n6985), .A(n6936), .B(n6935), .ZN(U3108)
         );
  AOI22_X1 U7875 ( .A1(n6939), .A2(n6978), .B1(n6938), .B2(n6976), .ZN(n6942)
         );
  AOI22_X1 U7876 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6982), .B1(n6940), 
        .B2(n6980), .ZN(n6941) );
  OAI211_X1 U7877 ( .C1(n6943), .C2(n6985), .A(n6942), .B(n6941), .ZN(U3109)
         );
  AOI22_X1 U7878 ( .A1(n6945), .A2(n6978), .B1(n6944), .B2(n6976), .ZN(n6948)
         );
  AOI22_X1 U7879 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6982), .B1(n6946), 
        .B2(n6980), .ZN(n6947) );
  OAI211_X1 U7880 ( .C1(n6949), .C2(n6985), .A(n6948), .B(n6947), .ZN(U3110)
         );
  INV_X1 U7881 ( .A(n6985), .ZN(n6969) );
  AOI22_X1 U7882 ( .A1(n6951), .A2(n6978), .B1(n6969), .B2(n6950), .ZN(n6954)
         );
  AOI22_X1 U7883 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6982), .B1(n6952), 
        .B2(n6980), .ZN(n6953) );
  OAI211_X1 U7884 ( .C1(n6955), .C2(n6974), .A(n6954), .B(n6953), .ZN(U3111)
         );
  AOI22_X1 U7885 ( .A1(n6957), .A2(n6978), .B1(n6969), .B2(n6956), .ZN(n6960)
         );
  AOI22_X1 U7886 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6982), .B1(n6958), 
        .B2(n6980), .ZN(n6959) );
  OAI211_X1 U7887 ( .C1(n6961), .C2(n6974), .A(n6960), .B(n6959), .ZN(U3112)
         );
  AOI22_X1 U7888 ( .A1(n6963), .A2(n6978), .B1(n6962), .B2(n6976), .ZN(n6966)
         );
  AOI22_X1 U7889 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6982), .B1(n6964), 
        .B2(n6980), .ZN(n6965) );
  OAI211_X1 U7890 ( .C1(n6967), .C2(n6985), .A(n6966), .B(n6965), .ZN(U3113)
         );
  AOI22_X1 U7891 ( .A1(n6970), .A2(n6978), .B1(n6969), .B2(n6968), .ZN(n6973)
         );
  AOI22_X1 U7892 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6982), .B1(n6971), 
        .B2(n6980), .ZN(n6972) );
  OAI211_X1 U7893 ( .C1(n6975), .C2(n6974), .A(n6973), .B(n6972), .ZN(U3114)
         );
  AOI22_X1 U7894 ( .A1(n6979), .A2(n6978), .B1(n6977), .B2(n6976), .ZN(n6984)
         );
  AOI22_X1 U7895 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6982), .B1(n6981), 
        .B2(n6980), .ZN(n6983) );
  OAI211_X1 U7896 ( .C1(n6986), .C2(n6985), .A(n6984), .B(n6983), .ZN(U3115)
         );
  OAI21_X1 U7897 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6987), 
        .ZN(n6988) );
  NAND4_X1 U7898 ( .A1(n6991), .A2(n6990), .A3(n6989), .A4(n6988), .ZN(n6993)
         );
  NOR2_X1 U7899 ( .A1(n6993), .A2(n6992), .ZN(n7019) );
  NAND2_X1 U7900 ( .A1(n6995), .A2(n6994), .ZN(n6998) );
  NAND2_X1 U7901 ( .A1(n6996), .A2(n3272), .ZN(n6997) );
  NAND2_X1 U7902 ( .A1(n6998), .A2(n6997), .ZN(n7139) );
  NAND2_X1 U7903 ( .A1(n6999), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n7148) );
  INV_X1 U7904 ( .A(n7148), .ZN(n7001) );
  OR3_X1 U7905 ( .A1(n7139), .A2(n7001), .A3(n7000), .ZN(n7004) );
  INV_X1 U7906 ( .A(n7004), .ZN(n7008) );
  NAND2_X1 U7907 ( .A1(n7011), .A2(n7010), .ZN(n7007) );
  OAI211_X1 U7908 ( .C1(n7005), .C2(n7004), .A(n7003), .B(n7002), .ZN(n7006)
         );
  OAI211_X1 U7909 ( .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n7008), .A(n7007), .B(n7006), .ZN(n7009) );
  OAI21_X1 U7910 ( .B1(n7011), .B2(n7010), .A(n7009), .ZN(n7013) );
  NAND2_X1 U7911 ( .A1(n7017), .A2(n7016), .ZN(n7012) );
  NAND2_X1 U7912 ( .A1(n7013), .A2(n7012), .ZN(n7015) );
  OAI211_X1 U7913 ( .C1(n7017), .C2(n7016), .A(n7015), .B(n7014), .ZN(n7018)
         );
  AND2_X1 U7914 ( .A1(n7019), .A2(n7018), .ZN(n7034) );
  NAND2_X1 U7916 ( .A1(n7034), .A2(n7036), .ZN(n7021) );
  NAND2_X1 U7917 ( .A1(n7160), .A2(READY_N), .ZN(n7020) );
  NAND2_X1 U7918 ( .A1(n7021), .A2(n7020), .ZN(n7025) );
  OR2_X1 U7919 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  AOI21_X1 U7920 ( .B1(n7026), .B2(n7163), .A(n7042), .ZN(n7029) );
  INV_X1 U7921 ( .A(n7042), .ZN(n7138) );
  OAI21_X1 U7922 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4043), .A(n7138), .ZN(
        n7038) );
  OAI33_X1 U7923 ( .A1(1'b0), .A2(n7029), .A3(STATE2_REG_0__SCAN_IN), .B1(
        n7028), .B2(n7027), .B3(n7038), .ZN(n7032) );
  OAI211_X1 U7924 ( .C1(n7034), .C2(n7033), .A(n7032), .B(n7031), .ZN(U3148)
         );
  INV_X1 U7925 ( .A(n7035), .ZN(n7037) );
  AOI21_X1 U7926 ( .B1(n7037), .B2(n4043), .A(n7036), .ZN(n7041) );
  OAI211_X1 U7927 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n7038), .ZN(n7039) );
  OAI211_X1 U7928 ( .C1(n7042), .C2(n7041), .A(n7040), .B(n7039), .ZN(U3149)
         );
  INV_X1 U7929 ( .A(n7043), .ZN(n7136) );
  OAI221_X1 U7930 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n4043), .A(n7136), .ZN(n7045) );
  OAI21_X1 U7931 ( .B1(n7163), .B2(n7045), .A(n7044), .ZN(U3150) );
  INV_X1 U7932 ( .A(n7135), .ZN(n7053) );
  AND2_X1 U7933 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n7053), .ZN(U3151) );
  AND2_X1 U7934 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n7053), .ZN(U3152) );
  NOR2_X1 U7935 ( .A1(n7135), .A2(n7046), .ZN(U3153) );
  AND2_X1 U7936 ( .A1(n7053), .A2(DATAWIDTH_REG_28__SCAN_IN), .ZN(U3154) );
  AND2_X1 U7937 ( .A1(n7053), .A2(DATAWIDTH_REG_27__SCAN_IN), .ZN(U3155) );
  NOR2_X1 U7938 ( .A1(n7135), .A2(n7047), .ZN(U3156) );
  AND2_X1 U7939 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n7053), .ZN(U3157) );
  AND2_X1 U7940 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n7053), .ZN(U3158) );
  AND2_X1 U7941 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n7053), .ZN(U3159) );
  AND2_X1 U7942 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n7053), .ZN(U3160) );
  NOR2_X1 U7943 ( .A1(n7135), .A2(n7048), .ZN(U3161) );
  AND2_X1 U7944 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n7053), .ZN(U3162) );
  AND2_X1 U7945 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n7053), .ZN(U3163) );
  AND2_X1 U7946 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n7053), .ZN(U3164) );
  AND2_X1 U7947 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n7053), .ZN(U3165) );
  NOR2_X1 U7948 ( .A1(n7135), .A2(n7049), .ZN(U3166) );
  AND2_X1 U7949 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n7053), .ZN(U3167) );
  AND2_X1 U7950 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n7053), .ZN(U3168) );
  AND2_X1 U7951 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n7053), .ZN(U3169) );
  NOR2_X1 U7952 ( .A1(n7135), .A2(n7050), .ZN(U3170) );
  AND2_X1 U7953 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n7053), .ZN(U3171) );
  AND2_X1 U7954 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n7053), .ZN(U3172) );
  AND2_X1 U7955 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n7053), .ZN(U3173) );
  NOR2_X1 U7956 ( .A1(n7135), .A2(n7051), .ZN(U3174) );
  AND2_X1 U7957 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n7053), .ZN(U3175) );
  AND2_X1 U7958 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n7053), .ZN(U3176) );
  AND2_X1 U7959 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n7053), .ZN(U3177) );
  AND2_X1 U7960 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n7053), .ZN(U3178) );
  NOR2_X1 U7961 ( .A1(n7135), .A2(n7052), .ZN(U3179) );
  AND2_X1 U7962 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n7053), .ZN(U3180) );
  NOR2_X1 U7963 ( .A1(n7072), .A2(n7055), .ZN(n7065) );
  NOR2_X1 U7964 ( .A1(n7072), .A2(n7054), .ZN(n7062) );
  AOI21_X1 U7965 ( .B1(STATE_REG_1__SCAN_IN), .B2(READY_N), .A(n7062), .ZN(
        n7069) );
  NOR2_X1 U7966 ( .A1(n7055), .A2(n7054), .ZN(n7058) );
  INV_X1 U7967 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7057) );
  AOI211_X1 U7968 ( .C1(STATE_REG_2__SCAN_IN), .C2(n7066), .A(
        STATE_REG_0__SCAN_IN), .B(n7065), .ZN(n7071) );
  AOI221_X1 U7969 ( .B1(n7058), .B2(n7168), .C1(n7057), .C2(n7168), .A(n7071), 
        .ZN(n7056) );
  OAI21_X1 U7970 ( .B1(n7065), .B2(n7069), .A(n7056), .ZN(U3181) );
  NOR2_X1 U7971 ( .A1(n7063), .A2(n7057), .ZN(n7067) );
  NOR2_X1 U7972 ( .A1(n7067), .A2(n7058), .ZN(n7061) );
  NAND2_X1 U7973 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n7059) );
  OAI211_X1 U7974 ( .C1(n7062), .C2(n7061), .A(n7060), .B(n7059), .ZN(U3182)
         );
  AOI221_X1 U7975 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4043), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7064) );
  AOI221_X1 U7976 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n7064), .C2(HOLD), .A(n7063), .ZN(n7070) );
  AOI21_X1 U7977 ( .B1(n7067), .B2(n7066), .A(n7065), .ZN(n7068) );
  OAI22_X1 U7978 ( .A1(n7071), .A2(n7070), .B1(n7069), .B2(n7068), .ZN(U3183)
         );
  NOR2_X1 U7979 ( .A1(n7072), .A2(n7168), .ZN(n7112) );
  INV_X1 U7980 ( .A(n7112), .ZN(n7127) );
  NAND2_X1 U7981 ( .A1(n7072), .A2(n7130), .ZN(n7122) );
  INV_X1 U7982 ( .A(n7122), .ZN(n7125) );
  AOI22_X1 U7983 ( .A1(REIP_REG_2__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n7168), .ZN(n7073) );
  OAI21_X1 U7984 ( .B1(n7074), .B2(n7127), .A(n7073), .ZN(U3184) );
  AOI22_X1 U7985 ( .A1(REIP_REG_2__SCAN_IN), .A2(n7112), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n7168), .ZN(n7075) );
  OAI21_X1 U7986 ( .B1(n7077), .B2(n7122), .A(n7075), .ZN(U3185) );
  AOI22_X1 U7987 ( .A1(REIP_REG_4__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n7168), .ZN(n7076) );
  OAI21_X1 U7988 ( .B1(n7077), .B2(n7127), .A(n7076), .ZN(U3186) );
  AOI22_X1 U7989 ( .A1(REIP_REG_5__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n7168), .ZN(n7078) );
  OAI21_X1 U7990 ( .B1(n7079), .B2(n7127), .A(n7078), .ZN(U3187) );
  AOI22_X1 U7991 ( .A1(REIP_REG_5__SCAN_IN), .A2(n7112), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n7168), .ZN(n7080) );
  OAI21_X1 U7992 ( .B1(n7082), .B2(n7122), .A(n7080), .ZN(U3188) );
  AOI22_X1 U7993 ( .A1(REIP_REG_7__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n7168), .ZN(n7081) );
  OAI21_X1 U7994 ( .B1(n7082), .B2(n7127), .A(n7081), .ZN(U3189) );
  AOI22_X1 U7995 ( .A1(REIP_REG_7__SCAN_IN), .A2(n7112), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n7168), .ZN(n7083) );
  OAI21_X1 U7996 ( .B1(n7085), .B2(n7122), .A(n7083), .ZN(U3190) );
  AOI22_X1 U7997 ( .A1(REIP_REG_9__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n7168), .ZN(n7084) );
  OAI21_X1 U7998 ( .B1(n7085), .B2(n7127), .A(n7084), .ZN(U3191) );
  AOI22_X1 U7999 ( .A1(REIP_REG_9__SCAN_IN), .A2(n7112), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n7168), .ZN(n7086) );
  OAI21_X1 U8000 ( .B1(n7089), .B2(n7122), .A(n7086), .ZN(U3192) );
  OAI222_X1 U8001 ( .A1(n7127), .A2(n7089), .B1(n7088), .B2(n7130), .C1(n7087), 
        .C2(n7122), .ZN(U3193) );
  AOI22_X1 U8002 ( .A1(REIP_REG_11__SCAN_IN), .A2(n7112), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n7168), .ZN(n7090) );
  OAI21_X1 U8003 ( .B1(n7092), .B2(n7122), .A(n7090), .ZN(U3194) );
  AOI22_X1 U8004 ( .A1(REIP_REG_13__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n7168), .ZN(n7091) );
  OAI21_X1 U8005 ( .B1(n7092), .B2(n7127), .A(n7091), .ZN(U3195) );
  AOI22_X1 U8006 ( .A1(REIP_REG_13__SCAN_IN), .A2(n7112), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n7168), .ZN(n7093) );
  OAI21_X1 U8007 ( .B1(n7094), .B2(n7122), .A(n7093), .ZN(U3196) );
  AOI222_X1 U8008 ( .A1(n7125), .A2(REIP_REG_15__SCAN_IN), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n7168), .C1(REIP_REG_14__SCAN_IN), .C2(
        n7112), .ZN(n7095) );
  INV_X1 U8009 ( .A(n7095), .ZN(U3197) );
  OAI222_X1 U8010 ( .A1(n7127), .A2(n7097), .B1(n7096), .B2(n7130), .C1(n7099), 
        .C2(n7122), .ZN(U3198) );
  AOI22_X1 U8011 ( .A1(REIP_REG_17__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n7168), .ZN(n7098) );
  OAI21_X1 U8012 ( .B1(n7099), .B2(n7127), .A(n7098), .ZN(U3199) );
  AOI22_X1 U8013 ( .A1(REIP_REG_17__SCAN_IN), .A2(n7112), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n7168), .ZN(n7100) );
  OAI21_X1 U8014 ( .B1(n7101), .B2(n7122), .A(n7100), .ZN(U3200) );
  AOI22_X1 U8015 ( .A1(REIP_REG_18__SCAN_IN), .A2(n7112), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n7168), .ZN(n7102) );
  OAI21_X1 U8016 ( .B1(n7104), .B2(n7122), .A(n7102), .ZN(U3201) );
  AOI22_X1 U8017 ( .A1(REIP_REG_20__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n7168), .ZN(n7103) );
  OAI21_X1 U8018 ( .B1(n7104), .B2(n7127), .A(n7103), .ZN(U3202) );
  AOI22_X1 U8019 ( .A1(REIP_REG_20__SCAN_IN), .A2(n7112), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n7168), .ZN(n7105) );
  OAI21_X1 U8020 ( .B1(n7107), .B2(n7122), .A(n7105), .ZN(U3203) );
  AOI22_X1 U8021 ( .A1(REIP_REG_22__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n7168), .ZN(n7106) );
  OAI21_X1 U8022 ( .B1(n7107), .B2(n7127), .A(n7106), .ZN(U3204) );
  OAI222_X1 U8023 ( .A1(n7122), .A2(n7111), .B1(n7109), .B2(n7130), .C1(n7108), 
        .C2(n7127), .ZN(U3205) );
  AOI22_X1 U8024 ( .A1(REIP_REG_24__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n7168), .ZN(n7110) );
  OAI21_X1 U8025 ( .B1(n7111), .B2(n7127), .A(n7110), .ZN(U3206) );
  AOI22_X1 U8026 ( .A1(REIP_REG_24__SCAN_IN), .A2(n7112), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n7168), .ZN(n7113) );
  OAI21_X1 U8027 ( .B1(n7115), .B2(n7122), .A(n7113), .ZN(U3207) );
  AOI22_X1 U8028 ( .A1(REIP_REG_26__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n7168), .ZN(n7114) );
  OAI21_X1 U8029 ( .B1(n7115), .B2(n7127), .A(n7114), .ZN(U3208) );
  OAI222_X1 U8030 ( .A1(n7122), .A2(n7118), .B1(n7117), .B2(n7130), .C1(n7116), 
        .C2(n7127), .ZN(U3209) );
  OAI222_X1 U8031 ( .A1(n7122), .A2(n7121), .B1(n7119), .B2(n7130), .C1(n7118), 
        .C2(n7127), .ZN(U3210) );
  AOI22_X1 U8032 ( .A1(REIP_REG_29__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n7168), .ZN(n7120) );
  OAI21_X1 U8033 ( .B1(n7121), .B2(n7127), .A(n7120), .ZN(U3211) );
  OAI222_X1 U8034 ( .A1(n7127), .A2(n7124), .B1(n7123), .B2(n7130), .C1(n7128), 
        .C2(n7122), .ZN(U3212) );
  AOI22_X1 U8035 ( .A1(REIP_REG_31__SCAN_IN), .A2(n7125), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n7168), .ZN(n7126) );
  OAI21_X1 U8036 ( .B1(n7128), .B2(n7127), .A(n7126), .ZN(U3213) );
  MUX2_X1 U8037 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n7168), .Z(U3445) );
  OAI22_X1 U8038 ( .A1(n7168), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        BE_N_REG_2__SCAN_IN), .B2(n7130), .ZN(n7129) );
  INV_X1 U8039 ( .A(n7129), .ZN(U3446) );
  OAI22_X1 U8040 ( .A1(n7168), .A2(BYTEENABLE_REG_1__SCAN_IN), .B1(
        BE_N_REG_1__SCAN_IN), .B2(n7130), .ZN(n7131) );
  INV_X1 U8041 ( .A(n7131), .ZN(U3447) );
  MUX2_X1 U8042 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n7168), .Z(U3448) );
  OAI21_X1 U8043 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n7135), .A(n7133), .ZN(
        n7132) );
  INV_X1 U8044 ( .A(n7132), .ZN(U3451) );
  OAI21_X1 U8045 ( .B1(n7135), .B2(n7134), .A(n7133), .ZN(U3452) );
  OAI211_X1 U8046 ( .C1(n3454), .C2(n7138), .A(n7137), .B(n7136), .ZN(U3453)
         );
  INV_X1 U8047 ( .A(n7139), .ZN(n7143) );
  AOI211_X1 U8048 ( .C1(n4068), .C2(STATE2_REG_1__SCAN_IN), .A(n7141), .B(
        n7140), .ZN(n7142) );
  OAI21_X1 U8049 ( .B1(n7143), .B2(n7147), .A(n7142), .ZN(n7144) );
  OAI21_X1 U8050 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7145), .A(n7144), 
        .ZN(n7146) );
  OAI21_X1 U8051 ( .B1(n7148), .B2(n7147), .A(n7146), .ZN(U3461) );
  NAND2_X1 U8052 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n7152) );
  AOI211_X1 U8053 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(n7154), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7149) );
  AOI21_X1 U8054 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n7151), .A(n7149), .ZN(
        n7150) );
  OAI21_X1 U8055 ( .B1(n7152), .B2(n7151), .A(n7150), .ZN(U3468) );
  OAI22_X1 U8056 ( .A1(n7154), .A2(REIP_REG_0__SCAN_IN), .B1(
        BYTEENABLE_REG_0__SCAN_IN), .B2(n7153), .ZN(n7155) );
  INV_X1 U8057 ( .A(n7155), .ZN(U3469) );
  MUX2_X1 U8058 ( .A(n7156), .B(W_R_N_REG_SCAN_IN), .S(n7168), .Z(U3470) );
  INV_X1 U8059 ( .A(n7157), .ZN(n7158) );
  AOI211_X1 U8060 ( .C1(n7160), .C2(n4043), .A(n7159), .B(n7158), .ZN(n7167)
         );
  OAI211_X1 U8061 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n7162), .A(n7161), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n7164) );
  AOI21_X1 U8062 ( .B1(n7164), .B2(STATE2_REG_0__SCAN_IN), .A(n7163), .ZN(
        n7166) );
  NAND2_X1 U8063 ( .A1(n7167), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n7165) );
  OAI21_X1 U8064 ( .B1(n7167), .B2(n7166), .A(n7165), .ZN(U3472) );
  MUX2_X1 U8065 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n7168), .Z(U3473) );
  OR2_X1 U3738 ( .A1(n3182), .A2(n3195), .ZN(n3181) );
  CLKBUF_X1 U3637 ( .A(n3400), .Z(n5221) );
  NAND2_X1 U3653 ( .A1(n4142), .A2(n3518), .ZN(n3443) );
  XNOR2_X1 U3654 ( .A(n3639), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6686)
         );
  NAND2_X1 U3693 ( .A1(n3624), .A2(n3623), .ZN(n6817) );
endmodule

