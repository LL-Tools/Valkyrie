

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput127, keyinput126,
         keyinput125, keyinput124, keyinput123, keyinput122, keyinput121,
         keyinput120, keyinput119, keyinput118, keyinput117, keyinput116,
         keyinput115, keyinput114, keyinput113, keyinput112, keyinput111,
         keyinput110, keyinput109, keyinput108, keyinput107, keyinput106,
         keyinput105, keyinput104, keyinput103, keyinput102, keyinput101,
         keyinput100, keyinput99, keyinput98, keyinput97, keyinput96,
         keyinput95, keyinput94, keyinput93, keyinput92, keyinput91,
         keyinput90, keyinput89, keyinput88, keyinput87, keyinput86,
         keyinput85, keyinput84, keyinput83, keyinput82, keyinput81,
         keyinput80, keyinput79, keyinput78, keyinput77, keyinput76,
         keyinput75, keyinput74, keyinput73, keyinput72, keyinput71,
         keyinput70, keyinput69, keyinput68, keyinput67, keyinput66,
         keyinput65, keyinput64, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752;

  NAND2_X1 U3527 ( .A1(n4644), .A2(n4643), .ZN(n4642) );
  CLKBUF_X1 U3528 ( .A(n3889), .Z(n4144) );
  CLKBUF_X2 U3529 ( .A(n3313), .Z(n4772) );
  CLKBUF_X2 U3530 ( .A(n3191), .Z(n3081) );
  CLKBUF_X2 U3531 ( .A(n3314), .Z(n3797) );
  CLKBUF_X2 U3532 ( .A(n3306), .Z(n4782) );
  CLKBUF_X2 U3533 ( .A(n3288), .Z(n4775) );
  CLKBUF_X2 U3534 ( .A(n3192), .Z(n3080) );
  CLKBUF_X1 U3535 ( .A(n3207), .Z(n4446) );
  AND2_X2 U3536 ( .A1(n3115), .A2(n4681), .ZN(n3447) );
  AND2_X2 U3537 ( .A1(n3117), .A2(n4362), .ZN(n3306) );
  CLKBUF_X1 U3538 ( .A(n4746), .Z(n3079) );
  NOR2_X1 U3539 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4746) );
  AND2_X1 U3540 ( .A1(n4248), .A2(n4362), .ZN(n3288) );
  CLKBUF_X2 U3541 ( .A(n3307), .Z(n4783) );
  CLKBUF_X2 U3542 ( .A(n3164), .Z(n4774) );
  AOI22_X1 U3543 ( .A1(n6633), .A2(keyinput34), .B1(keyinput72), .B2(n6632), 
        .ZN(n6631) );
  AOI21_X1 U3544 ( .B1(n6633), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3684) );
  OR2_X1 U3545 ( .A1(n4077), .A2(n4076), .ZN(n4078) );
  OAI221_X1 U3546 ( .B1(n6633), .B2(keyinput34), .C1(n6632), .C2(keyinput72), 
        .A(n6631), .ZN(n6642) );
  OR2_X1 U3547 ( .A1(n4692), .A2(n4987), .ZN(n4154) );
  INV_X1 U3548 ( .A(n3093), .ZN(n4987) );
  INV_X1 U3549 ( .A(n5513), .ZN(n5487) );
  NAND2_X1 U3550 ( .A1(n5136), .A2(n5135), .ZN(n5138) );
  INV_X2 U3551 ( .A(n4178), .ZN(n5054) );
  CLKBUF_X2 U3552 ( .A(n3175), .Z(n4773) );
  INV_X2 U3553 ( .A(n4159), .ZN(n4390) );
  NOR4_X1 U3554 ( .A1(n5094), .A2(REIP_REG_31__SCAN_IN), .A3(n6374), .A4(n6370), .ZN(n4900) );
  INV_X1 U3555 ( .A(n5452), .ZN(n5465) );
  AND2_X1 U3556 ( .A1(n4923), .A2(n4922), .ZN(n5207) );
  AND2_X2 U3557 ( .A1(n4977), .A2(n4967), .ZN(n4151) );
  OR2_X1 U3558 ( .A1(n4935), .A2(n5150), .ZN(n5152) );
  AND2_X1 U3559 ( .A1(n3347), .A2(n3346), .ZN(n5802) );
  INV_X1 U3560 ( .A(n5520), .ZN(n5512) );
  INV_X1 U3561 ( .A(n5679), .ZN(n5371) );
  AND3_X2 U3562 ( .A1(n3230), .A2(n3229), .A3(n3228), .ZN(n4126) );
  NAND2_X2 U3563 ( .A1(n3303), .A2(n3302), .ZN(n5805) );
  INV_X1 U3564 ( .A(n3470), .ZN(n3852) );
  OR2_X4 U3565 ( .A1(n3123), .A2(n3122), .ZN(n3996) );
  CLKBUF_X3 U3566 ( .A(n4002), .Z(n4263) );
  XNOR2_X2 U3567 ( .A(n3267), .B(n3266), .ZN(n3363) );
  OAI22_X2 U3568 ( .A1(n4267), .A2(STATE2_REG_0__SCAN_IN), .B1(n4004), .B2(
        n3263), .ZN(n3267) );
  AND2_X4 U3569 ( .A1(n4686), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3115)
         );
  OR2_X2 U3570 ( .A1(n4009), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5664)
         );
  OAI21_X2 U3571 ( .B1(n3815), .B2(n3814), .A(n4972), .ZN(n4854) );
  NAND2_X1 U3572 ( .A1(n4151), .A2(n4874), .ZN(n4692) );
  NOR2_X1 U3573 ( .A1(n5487), .A2(n3975), .ZN(n4954) );
  NAND2_X1 U3574 ( .A1(n5314), .A2(n5313), .ZN(n4935) );
  CLKBUF_X2 U3575 ( .A(n4936), .Z(n3093) );
  BUF_X1 U3576 ( .A(n5364), .Z(n3095) );
  OR2_X1 U3577 ( .A1(n3372), .A2(n6303), .ZN(n3470) );
  NAND2_X1 U3578 ( .A1(n3990), .A2(n3878), .ZN(n4936) );
  NOR2_X1 U3579 ( .A1(n3882), .A2(n3878), .ZN(n5364) );
  INV_X2 U3580 ( .A(n3996), .ZN(n3231) );
  OR2_X2 U3581 ( .A1(n3153), .A2(n3152), .ZN(n4159) );
  NOR2_X4 U3582 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4248) );
  INV_X2 U3583 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4686) );
  AOI22_X1 U3584 ( .A1(n5679), .A2(n5307), .B1(n5348), .B2(
        REIP_REG_18__SCAN_IN), .ZN(n4819) );
  AOI21_X1 U3585 ( .B1(n5207), .B2(n5669), .A(n5206), .ZN(n5208) );
  AOI21_X1 U3586 ( .B1(n5224), .B2(n5288), .A(n5211), .ZN(n5021) );
  AND2_X1 U3587 ( .A1(n5260), .A2(n5679), .ZN(n5206) );
  XNOR2_X1 U3588 ( .A(n4893), .B(n4892), .ZN(n4917) );
  AND2_X1 U3589 ( .A1(n4843), .A2(n4842), .ZN(n5189) );
  OAI21_X1 U3590 ( .B1(n4081), .B2(n4080), .A(n4079), .ZN(n5205) );
  NOR2_X1 U3591 ( .A1(n4966), .A2(n4870), .ZN(n4889) );
  XNOR2_X1 U3592 ( .A(n4621), .B(n3570), .ZN(n4671) );
  NAND2_X1 U3593 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  NAND2_X1 U3594 ( .A1(n4154), .A2(n4153), .ZN(n4880) );
  INV_X1 U3595 ( .A(n4692), .ZN(n4694) );
  NOR2_X1 U3596 ( .A1(n5124), .A2(n5125), .ZN(n5118) );
  AND2_X2 U3597 ( .A1(n4057), .A2(n4056), .ZN(n4178) );
  AND3_X1 U3598 ( .A1(n4055), .A2(STATE2_REG_0__SCAN_IN), .A3(n4054), .ZN(
        n4056) );
  OR2_X1 U3599 ( .A1(n3360), .A2(n4221), .ZN(n4288) );
  AND2_X1 U3600 ( .A1(n4219), .A2(n4218), .ZN(n4221) );
  NAND2_X1 U3601 ( .A1(n3341), .A2(n3340), .ZN(n4219) );
  NAND2_X1 U3603 ( .A1(n3384), .A2(n3383), .ZN(n4379) );
  OR2_X2 U3604 ( .A1(n4642), .A2(n3930), .ZN(n4827) );
  CLKBUF_X1 U3605 ( .A(n4349), .Z(n6017) );
  NAND2_X2 U3606 ( .A1(n5604), .A2(n5603), .ZN(n5661) );
  AND2_X1 U3607 ( .A1(n5604), .A2(n5363), .ZN(n6430) );
  NAND2_X1 U3608 ( .A1(n3329), .A2(n3101), .ZN(n3335) );
  AND2_X1 U3609 ( .A1(n6282), .A2(n6293), .ZN(n5604) );
  OR2_X2 U3610 ( .A1(n3862), .A2(n3861), .ZN(n6282) );
  NAND2_X1 U3611 ( .A1(n3301), .A2(n3300), .ZN(n3302) );
  AND3_X1 U3612 ( .A1(n4111), .A2(n3224), .A3(n3223), .ZN(n3300) );
  NAND2_X1 U3613 ( .A1(n3884), .A2(n3883), .ZN(n3888) );
  NOR2_X1 U3614 ( .A1(n3222), .A2(n3208), .ZN(n3209) );
  NAND2_X1 U3615 ( .A1(n4243), .A2(n3205), .ZN(n3220) );
  OR2_X1 U3616 ( .A1(n4241), .A2(n4299), .ZN(n4160) );
  NAND2_X1 U3617 ( .A1(n4222), .A2(n4987), .ZN(n3959) );
  OR2_X1 U3618 ( .A1(n4222), .A2(n3967), .ZN(n3961) );
  INV_X1 U3619 ( .A(n4091), .ZN(n3230) );
  BUF_X1 U3620 ( .A(n3890), .Z(n3967) );
  OR2_X1 U3621 ( .A1(n3834), .A2(n4936), .ZN(n4243) );
  AND2_X1 U3622 ( .A1(n3372), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3858) );
  BUF_X2 U3623 ( .A(n3894), .Z(n4156) );
  AND2_X2 U3624 ( .A1(n4279), .A2(n3882), .ZN(n5605) );
  NAND2_X1 U3625 ( .A1(n4485), .A2(n4301), .ZN(n4120) );
  OR2_X1 U3626 ( .A1(n3295), .A2(n3294), .ZN(n4055) );
  INV_X1 U3627 ( .A(n3882), .ZN(n4334) );
  OR2_X2 U3628 ( .A1(n3174), .A2(n3173), .ZN(n3990) );
  OR2_X2 U3629 ( .A1(n3143), .A2(n3142), .ZN(n4301) );
  AND2_X2 U3630 ( .A1(n3996), .A2(n3878), .ZN(n4046) );
  OR2_X1 U3631 ( .A1(n3163), .A2(n3162), .ZN(n4116) );
  BUF_X2 U3632 ( .A(n3283), .Z(n4780) );
  BUF_X2 U3633 ( .A(n3312), .Z(n3289) );
  AND2_X2 U3634 ( .A1(n3115), .A2(n4681), .ZN(n3098) );
  BUF_X2 U3635 ( .A(n3315), .Z(n3082) );
  AND2_X2 U3636 ( .A1(n3115), .A2(n4248), .ZN(n3192) );
  CLKBUF_X2 U3637 ( .A(n5593), .Z(n6421) );
  BUF_X2 U3638 ( .A(n3425), .Z(n3772) );
  AOI22_X1 U3639 ( .A1(n6572), .A2(keyinput118), .B1(keyinput46), .B2(n6571), 
        .ZN(n6570) );
  AND2_X2 U3640 ( .A1(n3237), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4252)
         );
  INV_X2 U3641 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3109) );
  INV_X1 U3642 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3237) );
  NAND2_X1 U3643 ( .A1(n3396), .A2(n3395), .ZN(n3438) );
  OR2_X1 U3644 ( .A1(n3360), .A2(n4221), .ZN(n3083) );
  INV_X1 U3645 ( .A(n3996), .ZN(n3084) );
  INV_X1 U3646 ( .A(n3305), .ZN(n3085) );
  INV_X1 U3647 ( .A(n3085), .ZN(n3086) );
  AND2_X2 U3648 ( .A1(n4252), .A2(n4362), .ZN(n3305) );
  AND2_X1 U3649 ( .A1(n5138), .A2(n5137), .ZN(n5215) );
  NAND2_X1 U3650 ( .A1(n4263), .A2(n3090), .ZN(n3087) );
  NAND2_X1 U3651 ( .A1(n3087), .A2(n3088), .ZN(n5663) );
  OR2_X1 U3652 ( .A1(n3089), .A2(n4007), .ZN(n3088) );
  INV_X1 U3653 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3089) );
  AND2_X1 U3654 ( .A1(n4046), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3090)
         );
  INV_X1 U3655 ( .A(n5363), .ZN(n3091) );
  NAND2_X1 U3656 ( .A1(n4061), .A2(n4060), .ZN(n4519) );
  NAND2_X1 U3657 ( .A1(n3227), .A2(n3882), .ZN(n6274) );
  XNOR2_X1 U3658 ( .A(n3364), .B(n4268), .ZN(n4349) );
  NAND2_X1 U3659 ( .A1(n4428), .A2(n4456), .ZN(n4455) );
  CLKBUF_X3 U3660 ( .A(n4936), .Z(n3094) );
  NAND2_X2 U3661 ( .A1(n4126), .A2(n3095), .ZN(n4370) );
  NAND2_X1 U3662 ( .A1(n3214), .A2(n3213), .ZN(n3299) );
  INV_X1 U3663 ( .A(n4242), .ZN(n3227) );
  AND2_X2 U3664 ( .A1(n3114), .A2(n4681), .ZN(n3175) );
  AND2_X1 U3665 ( .A1(n4248), .A2(n4362), .ZN(n3092) );
  NOR2_X4 U3666 ( .A1(n4827), .A2(n5331), .ZN(n5332) );
  AND2_X2 U3667 ( .A1(n4681), .A2(n4362), .ZN(n3307) );
  NAND2_X2 U3668 ( .A1(n3362), .A2(n3361), .ZN(n4258) );
  OR2_X2 U3669 ( .A1(n4255), .A2(n4256), .ZN(n4317) );
  AND2_X2 U3670 ( .A1(n3115), .A2(n4252), .ZN(n3191) );
  AND2_X2 U3671 ( .A1(n3117), .A2(n3116), .ZN(n3315) );
  NOR2_X2 U3672 ( .A1(n5152), .A2(n3949), .ZN(n5131) );
  OAI21_X2 U3673 ( .B1(n4321), .B2(n4320), .A(n4015), .ZN(n4326) );
  OAI21_X2 U3674 ( .B1(n4519), .B2(n4063), .A(n4062), .ZN(n4530) );
  OAI21_X2 U3675 ( .B1(n4671), .B2(n4672), .A(n3571), .ZN(n4822) );
  OAI21_X2 U3676 ( .B1(n4530), .B2(n4526), .A(n4527), .ZN(n4627) );
  XNOR2_X1 U3677 ( .A(n3337), .B(n3336), .ZN(n3993) );
  AOI21_X4 U3678 ( .B1(n5056), .B2(n4811), .A(n4810), .ZN(n5227) );
  NAND2_X2 U3679 ( .A1(n4808), .A2(n4807), .ZN(n5056) );
  AND2_X2 U3680 ( .A1(n3115), .A2(n4681), .ZN(n3097) );
  NOR2_X4 U3681 ( .A1(n4613), .A2(n4612), .ZN(n4644) );
  AOI211_X2 U3682 ( .C1(n5083), .C2(n5754), .A(n4705), .B(n4699), .ZN(n4702)
         );
  NAND2_X1 U3683 ( .A1(n3230), .A2(n3226), .ZN(n4242) );
  AND2_X1 U3684 ( .A1(n4807), .A2(n4068), .ZN(n4176) );
  AND2_X1 U3685 ( .A1(n5044), .A2(n5047), .ZN(n4811) );
  OR2_X1 U3686 ( .A1(n4247), .A2(n4123), .ZN(n4127) );
  OR2_X1 U3687 ( .A1(n4120), .A2(n3572), .ZN(n4088) );
  NAND2_X1 U3688 ( .A1(n3852), .A2(n4046), .ZN(n3859) );
  OR3_X1 U3689 ( .A1(READY_N), .A2(n4295), .A3(n4294), .ZN(n5609) );
  NAND2_X1 U3690 ( .A1(n4102), .A2(n4101), .ZN(n4162) );
  NAND2_X1 U3691 ( .A1(n4237), .A2(n4236), .ZN(n6266) );
  OR2_X1 U3692 ( .A1(n3096), .A2(n5777), .ZN(n6121) );
  OR2_X1 U3693 ( .A1(n6298), .A2(n3871), .ZN(n3872) );
  OAI21_X1 U3694 ( .B1(n3470), .B2(n3409), .A(n3408), .ZN(n3436) );
  NOR2_X1 U3695 ( .A1(n3095), .A2(n3826), .ZN(n3850) );
  NAND2_X1 U3696 ( .A1(n6261), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4767) );
  NOR2_X2 U3697 ( .A1(n3332), .A2(n6550), .ZN(n3615) );
  NOR2_X1 U3698 ( .A1(n4159), .A2(n6303), .ZN(n3326) );
  NOR2_X1 U3699 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4278), .ZN(n5841) );
  AND2_X1 U3700 ( .A1(n4095), .A2(n6276), .ZN(n5362) );
  AND2_X1 U3701 ( .A1(n3410), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3441)
         );
  NOR2_X1 U3702 ( .A1(n4127), .A2(n4125), .ZN(n6278) );
  INV_X1 U3703 ( .A(n3557), .ZN(n4890) );
  NAND2_X1 U3704 ( .A1(n4752), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4751)
         );
  NAND2_X1 U3705 ( .A1(n3771), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3874)
         );
  NAND2_X1 U3706 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3704), .ZN(n3724)
         );
  NAND2_X1 U3707 ( .A1(n4822), .A2(n3639), .ZN(n5232) );
  NAND2_X1 U3708 ( .A1(n3441), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3463)
         );
  AOI21_X1 U3709 ( .B1(n5777), .B2(n3348), .A(n6550), .ZN(n4306) );
  NAND2_X1 U3710 ( .A1(n5224), .A2(n4082), .ZN(n4083) );
  INV_X1 U3711 ( .A(n4809), .ZN(n4810) );
  NAND2_X1 U3712 ( .A1(n3365), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3214) );
  CLKBUF_X1 U3713 ( .A(n4267), .Z(n5774) );
  INV_X1 U3714 ( .A(n5773), .ZN(n6087) );
  OR2_X1 U3715 ( .A1(n6121), .A2(n6159), .ZN(n6165) );
  AOI21_X1 U3716 ( .B1(n3858), .B2(n3869), .A(n3857), .ZN(n3862) );
  AND2_X1 U3717 ( .A1(n4372), .A2(n4371), .ZN(n6286) );
  INV_X1 U3718 ( .A(n6305), .ZN(n6293) );
  NAND2_X1 U3719 ( .A1(n5362), .A2(n6293), .ZN(n6435) );
  NAND2_X1 U3720 ( .A1(n5486), .A2(n3877), .ZN(n5452) );
  AND2_X1 U3721 ( .A1(n4895), .A2(n3881), .ZN(n5517) );
  AND2_X1 U3722 ( .A1(n5566), .A2(n4300), .ZN(n5556) );
  AND2_X1 U3723 ( .A1(n5566), .A2(n4302), .ZN(n5559) );
  AND2_X1 U3724 ( .A1(n5566), .A2(n4298), .ZN(n5563) );
  INV_X1 U3725 ( .A(n5566), .ZN(n5558) );
  INV_X1 U3726 ( .A(n4198), .ZN(n4202) );
  NAND2_X1 U3727 ( .A1(n5371), .A2(n4188), .ZN(n5676) );
  XNOR2_X1 U3728 ( .A(n4180), .B(n5065), .ZN(n5269) );
  XNOR2_X1 U3729 ( .A(n5021), .B(n4840), .ZN(n5278) );
  NOR2_X1 U3730 ( .A1(n5302), .A2(n4163), .ZN(n5285) );
  AND2_X1 U3731 ( .A1(n4162), .A2(n4161), .ZN(n5754) );
  XNOR2_X1 U3732 ( .A(n3335), .B(n3334), .ZN(n3336) );
  AOI22_X1 U3733 ( .A1(n3164), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3155) );
  CLKBUF_X2 U3734 ( .A(n3086), .Z(n4781) );
  NOR2_X1 U3735 ( .A1(n3438), .A2(n3437), .ZN(n3472) );
  NOR2_X2 U3736 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3116) );
  AND2_X2 U3737 ( .A1(n6260), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3117)
         );
  AND2_X1 U3738 ( .A1(n4390), .A2(n4301), .ZN(n3204) );
  OR2_X1 U3739 ( .A1(n3382), .A2(n3381), .ZN(n4018) );
  NAND2_X1 U3740 ( .A1(n3882), .A2(n4159), .ZN(n3372) );
  NOR2_X1 U3741 ( .A1(n3820), .A2(n3827), .ZN(n3821) );
  NOR2_X1 U3742 ( .A1(n3724), .A2(n3723), .ZN(n3759) );
  INV_X1 U3743 ( .A(n4455), .ZN(n3511) );
  XNOR2_X1 U3744 ( .A(n3438), .B(n3436), .ZN(n4016) );
  AND2_X1 U3745 ( .A1(n3106), .A2(n5045), .ZN(n4809) );
  OR2_X1 U3746 ( .A1(n3280), .A2(n3279), .ZN(n3995) );
  OR3_X1 U3747 ( .A1(n4380), .A2(n3096), .A3(n4263), .ZN(n5804) );
  AND2_X1 U3748 ( .A1(n6018), .A2(n6017), .ZN(n6052) );
  INV_X1 U3749 ( .A(n4116), .ZN(n3207) );
  AOI21_X1 U3750 ( .B1(n6311), .B2(n5074), .A(n4680), .ZN(n4278) );
  AND2_X2 U3751 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4362) );
  AND2_X1 U3752 ( .A1(n4090), .A2(n4089), .ZN(n4105) );
  OAI21_X1 U3753 ( .B1(n3859), .B2(n3867), .A(n3856), .ZN(n3857) );
  INV_X1 U3754 ( .A(n3386), .ZN(n3387) );
  NAND2_X1 U3755 ( .A1(n3387), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3412)
         );
  AND2_X1 U3756 ( .A1(n5604), .A2(n5076), .ZN(n5583) );
  NOR2_X1 U3757 ( .A1(n3874), .A2(n3873), .ZN(n4706) );
  NAND2_X1 U3758 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n4706), .ZN(n4745)
         );
  AND2_X1 U3759 ( .A1(n3809), .A2(n3808), .ZN(n3814) );
  AND2_X1 U3760 ( .A1(n3790), .A2(n3789), .ZN(n4920) );
  AND2_X1 U3761 ( .A1(n3759), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3770)
         );
  AND2_X1 U3762 ( .A1(n3706), .A2(n3705), .ZN(n5135) );
  NOR2_X1 U3763 ( .A1(n6633), .A2(n3687), .ZN(n3704) );
  NAND2_X1 U3764 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3687)
         );
  AND2_X1 U3765 ( .A1(n3605), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3589)
         );
  NAND2_X1 U3766 ( .A1(n3589), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3657)
         );
  INV_X1 U3767 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6571) );
  AND2_X1 U3768 ( .A1(n3622), .A2(n3621), .ZN(n5007) );
  OR2_X1 U3769 ( .A1(n5006), .A2(n5007), .ZN(n5004) );
  NOR2_X1 U3770 ( .A1(n3588), .A2(n3587), .ZN(n3633) );
  NAND2_X1 U3771 ( .A1(n3556), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3588)
         );
  NOR2_X1 U3772 ( .A1(n3542), .A2(n3541), .ZN(n3556) );
  INV_X1 U3773 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3541) );
  NAND2_X1 U3774 ( .A1(n3536), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3542)
         );
  AND3_X1 U3775 ( .A1(n3525), .A2(n3524), .A3(n3523), .ZN(n4600) );
  NAND2_X1 U3777 ( .A1(n3493), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3494)
         );
  NOR2_X1 U3778 ( .A1(n6638), .A2(n3494), .ZN(n3536) );
  CLKBUF_X1 U3779 ( .A(n4513), .Z(n4599) );
  NAND2_X1 U3780 ( .A1(n3474), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3492)
         );
  NOR2_X1 U3781 ( .A1(n6711), .A2(n3463), .ZN(n3474) );
  AOI21_X1 U3782 ( .B1(n3446), .B2(n3615), .A(n3445), .ZN(n4309) );
  NAND2_X1 U3783 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3386) );
  NAND2_X1 U3784 ( .A1(n4078), .A2(n5224), .ZN(n4079) );
  AND2_X1 U3785 ( .A1(n3963), .A2(n3962), .ZN(n4207) );
  AND2_X1 U3786 ( .A1(n3954), .A2(n3953), .ZN(n4982) );
  INV_X1 U3787 ( .A(n4981), .ZN(n5114) );
  INV_X1 U3788 ( .A(n4170), .ZN(n4171) );
  AND2_X1 U3789 ( .A1(n3933), .A2(n3932), .ZN(n5331) );
  AND2_X1 U3790 ( .A1(n3929), .A2(n3928), .ZN(n4824) );
  NAND2_X1 U3791 ( .A1(n4169), .A2(n4638), .ZN(n4662) );
  AND2_X1 U3792 ( .A1(n3923), .A2(n3922), .ZN(n4643) );
  AND2_X1 U3793 ( .A1(n3916), .A2(n3915), .ZN(n4545) );
  NAND2_X1 U3794 ( .A1(n4162), .A2(n6278), .ZN(n5741) );
  AOI21_X1 U3795 ( .B1(n4223), .B2(n4222), .A(n3888), .ZN(n5515) );
  INV_X1 U3796 ( .A(n5768), .ZN(n4136) );
  NOR2_X1 U3797 ( .A1(n6396), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4187) );
  OR2_X1 U3798 ( .A1(n4242), .A2(n4156), .ZN(n4294) );
  NAND2_X1 U3799 ( .A1(n3304), .A2(n6303), .ZN(n3329) );
  INV_X1 U3800 ( .A(n3300), .ZN(n3225) );
  NAND2_X1 U3801 ( .A1(n3236), .A2(n3108), .ZN(n3268) );
  INV_X1 U3802 ( .A(n4088), .ZN(n6261) );
  INV_X1 U3803 ( .A(n3248), .ZN(n3249) );
  NAND2_X1 U3804 ( .A1(n3343), .A2(n3342), .ZN(n3347) );
  INV_X1 U3805 ( .A(n3345), .ZN(n3342) );
  INV_X1 U3806 ( .A(n5804), .ZN(n5803) );
  INV_X1 U3807 ( .A(n4263), .ZN(n4414) );
  INV_X1 U3808 ( .A(n5954), .ZN(n6082) );
  INV_X1 U3809 ( .A(n6159), .ZN(n6198) );
  AND2_X1 U3810 ( .A1(n3096), .A2(n5802), .ZN(n6046) );
  OR2_X1 U3811 ( .A1(n6382), .A2(n4278), .ZN(n4587) );
  OAI21_X1 U3812 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6384), .A(n5841), 
        .ZN(n6202) );
  AND2_X1 U3813 ( .A1(n4361), .A2(n4360), .ZN(n6271) );
  OR2_X1 U3814 ( .A1(n4242), .A2(n6423), .ZN(n6296) );
  INV_X1 U3815 ( .A(n6430), .ZN(n3870) );
  NAND2_X1 U3816 ( .A1(n3980), .A2(n5105), .ZN(n3987) );
  INV_X1 U3817 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6638) );
  AND2_X1 U3818 ( .A1(n5486), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5519) );
  AND2_X2 U3819 ( .A1(n4895), .A2(n3974), .ZN(n5513) );
  INV_X1 U3820 ( .A(n5555), .ZN(n5550) );
  AND2_X1 U3821 ( .A1(n5554), .A2(n4916), .ZN(n5549) );
  AND2_X1 U3822 ( .A1(n4217), .A2(n6293), .ZN(n5554) );
  OR2_X1 U3823 ( .A1(n5556), .A2(n5559), .ZN(n5562) );
  OAI21_X1 U3824 ( .B1(n4293), .B2(n4292), .A(n6293), .ZN(n4296) );
  INV_X1 U3825 ( .A(n5562), .ZN(n5008) );
  INV_X1 U3826 ( .A(n5563), .ZN(n5178) );
  NOR2_X1 U3828 ( .A1(n4751), .A2(n4703), .ZN(n3876) );
  INV_X1 U3829 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6633) );
  NOR2_X1 U3830 ( .A1(n5721), .A2(n4647), .ZN(n4536) );
  OR2_X1 U3831 ( .A1(n5241), .A2(n5252), .ZN(n4883) );
  NAND2_X1 U3832 ( .A1(n5197), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5013) );
  AND2_X1 U3833 ( .A1(n5238), .A2(n5237), .ZN(n5247) );
  NOR2_X1 U3834 ( .A1(n5272), .A2(n4164), .ZN(n5263) );
  NAND2_X1 U3835 ( .A1(n4817), .A2(n4816), .ZN(n4818) );
  NAND2_X1 U3836 ( .A1(n4815), .A2(n5224), .ZN(n4816) );
  NAND2_X1 U3837 ( .A1(n4813), .A2(n4178), .ZN(n4817) );
  NOR2_X1 U3838 ( .A1(n5336), .A2(n5324), .ZN(n5318) );
  NOR2_X1 U3839 ( .A1(n5741), .A2(n4648), .ZN(n5347) );
  NOR2_X1 U3840 ( .A1(n5752), .A2(n4646), .ZN(n4651) );
  INV_X1 U3841 ( .A(n5764), .ZN(n5733) );
  INV_X1 U3842 ( .A(n4536), .ZN(n5757) );
  INV_X1 U3843 ( .A(n5754), .ZN(n5771) );
  AND2_X1 U3844 ( .A1(n4162), .A2(n6264), .ZN(n5768) );
  INV_X1 U3845 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6113) );
  NOR2_X2 U3846 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6432) );
  INV_X1 U3847 ( .A(n6432), .ZN(n6203) );
  INV_X1 U3848 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U3849 ( .A1(n4374), .A2(n5961), .ZN(n6403) );
  INV_X1 U3850 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U3851 ( .A1(n6384), .A2(n6431), .ZN(n6396) );
  INV_X1 U3852 ( .A(n6394), .ZN(n6389) );
  INV_X1 U3853 ( .A(n5828), .ZN(n5830) );
  CLKBUF_X1 U3854 ( .A(n4580), .Z(n5873) );
  NOR2_X1 U3855 ( .A1(n6113), .A2(n5930), .ZN(n5949) );
  INV_X1 U3856 ( .A(n5982), .ZN(n5973) );
  AND2_X1 U3857 ( .A1(n5922), .A2(n6046), .ZN(n5982) );
  INV_X1 U3858 ( .A(n6081), .ZN(n6062) );
  OR2_X1 U3859 ( .A1(n6049), .A2(n6158), .ZN(n6081) );
  OR2_X1 U3860 ( .A1(n6092), .A2(n6170), .ZN(n6110) );
  OAI21_X1 U3861 ( .B1(n6187), .B2(n6384), .A(n6171), .ZN(n6189) );
  INV_X1 U3862 ( .A(n6165), .ZN(n6188) );
  INV_X1 U3863 ( .A(n6208), .ZN(n6253) );
  NAND2_X1 U3864 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6282), .ZN(n6386) );
  OR2_X1 U3865 ( .A1(n3863), .A2(n6303), .ZN(n6305) );
  AND2_X1 U3866 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6326), .ZN(n6429) );
  AOI211_X1 U3867 ( .C1(n5531), .C2(n5517), .A(n4901), .B(n4900), .ZN(n4905)
         );
  OAI21_X1 U3868 ( .B1(n5067), .B2(n5449), .A(n4210), .ZN(n4211) );
  INV_X1 U3869 ( .A(n4928), .ZN(n4210) );
  NAND2_X1 U3870 ( .A1(n5269), .A2(n5679), .ZN(n4197) );
  AOI21_X1 U3871 ( .B1(n3104), .B2(n5669), .A(n4195), .ZN(n4196) );
  NAND2_X1 U3872 ( .A1(n4194), .A2(n4193), .ZN(n4195) );
  INV_X1 U3873 ( .A(n5278), .ZN(n4848) );
  AND2_X1 U3874 ( .A1(n5267), .A2(n5754), .ZN(n5268) );
  OR2_X2 U3875 ( .A1(n4926), .A2(n3971), .ZN(n3099) );
  NOR2_X1 U3876 ( .A1(n5159), .A2(n5158), .ZN(n3100) );
  AND2_X1 U3877 ( .A1(n3328), .A2(n3327), .ZN(n3101) );
  INV_X1 U3878 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U3879 ( .A1(n5554), .A2(n4301), .ZN(n5555) );
  AND2_X1 U3880 ( .A1(n4279), .A2(n4301), .ZN(n3102) );
  NAND2_X1 U3881 ( .A1(n5224), .A2(n5299), .ZN(n3103) );
  AND2_X1 U3882 ( .A1(n4198), .A2(n4185), .ZN(n3104) );
  INV_X1 U3883 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4082) );
  NOR2_X1 U3884 ( .A1(n4963), .A2(n4750), .ZN(n3105) );
  INV_X1 U3885 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6586) );
  NAND2_X1 U3886 ( .A1(n5224), .A2(n5340), .ZN(n3106) );
  NAND2_X1 U3887 ( .A1(n4297), .A2(n4159), .ZN(n3107) );
  INV_X1 U3888 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6734) );
  INV_X1 U3889 ( .A(n5673), .ZN(n5233) );
  OR2_X1 U3890 ( .A1(n3238), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3108)
         );
  AND2_X1 U3891 ( .A1(n3228), .A2(n3102), .ZN(n3189) );
  AND2_X1 U3892 ( .A1(n3858), .A2(n3866), .ZN(n3845) );
  OR2_X1 U3893 ( .A1(n3262), .A2(n3261), .ZN(n3264) );
  AND2_X1 U3894 ( .A1(n6113), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3830)
         );
  INV_X1 U3895 ( .A(n3264), .ZN(n4004) );
  INV_X1 U3896 ( .A(n5273), .ZN(n4075) );
  XNOR2_X1 U3897 ( .A(n3109), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3827)
         );
  NOR2_X1 U3898 ( .A1(n3457), .A2(n3456), .ZN(n4044) );
  AND2_X1 U3899 ( .A1(n4379), .A2(n3394), .ZN(n3396) );
  NOR2_X1 U3900 ( .A1(n4301), .A2(n6550), .ZN(n3349) );
  NAND2_X1 U3901 ( .A1(n3472), .A2(n3471), .ZN(n4054) );
  INV_X1 U3902 ( .A(n3212), .ZN(n3213) );
  AOI21_X1 U3903 ( .B1(n3365), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3246), 
        .ZN(n3248) );
  INV_X1 U3904 ( .A(n3994), .ZN(n3324) );
  AOI21_X1 U3905 ( .B1(n6734), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3821), 
        .ZN(n3822) );
  NAND2_X1 U3906 ( .A1(n4222), .A2(n3094), .ZN(n3889) );
  INV_X1 U3907 ( .A(n4316), .ZN(n3419) );
  INV_X1 U3908 ( .A(n4745), .ZN(n3875) );
  INV_X1 U3909 ( .A(n3492), .ZN(n3493) );
  OR2_X1 U3910 ( .A1(n3431), .A2(n3430), .ZN(n4035) );
  INV_X1 U3911 ( .A(n3349), .ZN(n4723) );
  INV_X1 U3912 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5011) );
  AND2_X1 U3913 ( .A1(n4071), .A2(n4811), .ZN(n4170) );
  OR2_X1 U3914 ( .A1(n3321), .A2(n3320), .ZN(n3994) );
  NAND2_X1 U3915 ( .A1(n3371), .A2(n3370), .ZN(n4268) );
  AND2_X1 U3916 ( .A1(n6048), .A2(n3245), .ZN(n4421) );
  NAND2_X1 U3917 ( .A1(n3204), .A2(n4214), .ZN(n4091) );
  OR2_X1 U3918 ( .A1(n6630), .A2(n3823), .ZN(n3867) );
  NOR2_X1 U3919 ( .A1(n6622), .A2(n5388), .ZN(n5161) );
  INV_X1 U3920 ( .A(n4723), .ZN(n4797) );
  INV_X1 U3921 ( .A(n5113), .ZN(n3958) );
  INV_X1 U3922 ( .A(n3810), .ZN(n3769) );
  OR2_X1 U3923 ( .A1(n4621), .A2(n3570), .ZN(n3571) );
  AND2_X1 U3924 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n3875), .ZN(n4752)
         );
  INV_X1 U3925 ( .A(n5110), .ZN(n4192) );
  AND2_X1 U3926 ( .A1(n3638), .A2(n4946), .ZN(n3639) );
  INV_X1 U3927 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3587) );
  INV_X1 U3928 ( .A(n4514), .ZN(n3510) );
  NAND2_X1 U3929 ( .A1(n3440), .A2(n3439), .ZN(n4029) );
  NAND2_X1 U3930 ( .A1(n5196), .A2(n5011), .ZN(n5012) );
  AND2_X1 U3931 ( .A1(n4176), .A2(n4069), .ZN(n4172) );
  INV_X2 U3932 ( .A(n4178), .ZN(n5224) );
  AND2_X1 U3933 ( .A1(n3897), .A2(n3896), .ZN(n4256) );
  INV_X1 U3934 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6260) );
  OR2_X1 U3935 ( .A1(n3096), .A2(n6164), .ZN(n5986) );
  INV_X1 U3936 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6667) );
  OR2_X2 U3937 ( .A1(n3185), .A2(n3184), .ZN(n3878) );
  AND2_X1 U3938 ( .A1(n3869), .A2(n3860), .ZN(n3861) );
  NOR2_X1 U3939 ( .A1(n5505), .A2(n4855), .ZN(n3984) );
  INV_X1 U3940 ( .A(n3982), .ZN(n3985) );
  NOR2_X1 U3941 ( .A1(n6571), .A2(n3606), .ZN(n3605) );
  NAND2_X1 U3942 ( .A1(n3633), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3606)
         );
  INV_X1 U3943 ( .A(n3412), .ZN(n3410) );
  AND2_X1 U3944 ( .A1(n3920), .A2(n3919), .ZN(n4612) );
  INV_X1 U3945 ( .A(n3079), .ZN(n4795) );
  NAND2_X1 U3946 ( .A1(n5233), .A2(n4192), .ZN(n4193) );
  NOR2_X1 U3947 ( .A1(n3657), .A2(n3656), .ZN(n3658) );
  AND2_X1 U3948 ( .A1(n4949), .A2(n4948), .ZN(n5230) );
  NAND2_X1 U3949 ( .A1(n3511), .A2(n3510), .ZN(n4513) );
  INV_X1 U3950 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6711) );
  INV_X1 U3951 ( .A(n5262), .ZN(n4139) );
  NAND2_X1 U3952 ( .A1(n5013), .A2(n5012), .ZN(n5015) );
  AND2_X1 U3953 ( .A1(n3970), .A2(n3969), .ZN(n3971) );
  AOI21_X1 U3954 ( .B1(n4808), .B2(n4172), .A(n4171), .ZN(n5220) );
  AND2_X1 U3955 ( .A1(n3902), .A2(n3901), .ZN(n4406) );
  AOI21_X1 U3956 ( .B1(n5802), .B2(n4046), .A(n3991), .ZN(n5675) );
  NAND2_X1 U3957 ( .A1(n3345), .A2(n3344), .ZN(n3346) );
  INV_X1 U3958 ( .A(n5889), .ZN(n4488) );
  AND2_X1 U3959 ( .A1(n4263), .A2(n4264), .ZN(n5922) );
  INV_X2 U3960 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6550) );
  INV_X1 U3961 ( .A(n5605), .ZN(n6423) );
  NOR2_X1 U3962 ( .A1(n3985), .A2(n3984), .ZN(n3986) );
  NOR2_X1 U3963 ( .A1(n5162), .A2(n5154), .ZN(n5145) );
  OR2_X1 U3964 ( .A1(n6434), .A2(n3872), .ZN(n5486) );
  AND2_X1 U3965 ( .A1(n5486), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4895) );
  INV_X1 U3966 ( .A(n5505), .ZN(n5518) );
  AND2_X1 U3967 ( .A1(n5486), .A2(n3981), .ZN(n5520) );
  INV_X1 U3968 ( .A(n5554), .ZN(n5535) );
  INV_X1 U3969 ( .A(n4199), .ZN(n4201) );
  CLKBUF_X1 U3971 ( .A(n4260), .Z(n4315) );
  INV_X1 U3972 ( .A(n5609), .ZN(n5645) );
  OAI21_X1 U3973 ( .B1(n5605), .B2(n6420), .A(n6430), .ZN(n5658) );
  INV_X1 U3974 ( .A(n5107), .ZN(n5199) );
  AND2_X1 U3975 ( .A1(n3770), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3771)
         );
  AND2_X1 U3976 ( .A1(n3689), .A2(n3688), .ZN(n4992) );
  INV_X1 U3977 ( .A(n5676), .ZN(n5662) );
  AND2_X1 U3978 ( .A1(n5604), .A2(n4181), .ZN(n5679) );
  XNOR2_X1 U3979 ( .A(n5015), .B(n5014), .ZN(n5243) );
  OR2_X1 U3980 ( .A1(n5266), .A2(n4138), .ZN(n5262) );
  XNOR2_X1 U3981 ( .A(n4818), .B(n3941), .ZN(n5307) );
  NOR2_X1 U3982 ( .A1(n5690), .A2(n4664), .ZN(n5350) );
  INV_X1 U3983 ( .A(n5741), .ZN(n5721) );
  NAND2_X1 U3984 ( .A1(n4136), .A2(n4132), .ZN(n4647) );
  AND2_X1 U3985 ( .A1(n4162), .A2(n4107), .ZN(n5764) );
  INV_X1 U3986 ( .A(n5841), .ZN(n5961) );
  INV_X1 U3987 ( .A(n6386), .ZN(n4680) );
  OAI21_X1 U3988 ( .B1(n5782), .B2(n5781), .A(n5780), .ZN(n5799) );
  INV_X1 U3989 ( .A(n5802), .ZN(n5777) );
  OAI21_X1 U3990 ( .B1(n5842), .B2(n5858), .A(n6021), .ZN(n5859) );
  INV_X1 U3991 ( .A(n5884), .ZN(n4590) );
  AND2_X1 U3992 ( .A1(n5922), .A2(n6082), .ZN(n5889) );
  AND2_X1 U3993 ( .A1(n5922), .A2(n4281), .ZN(n5918) );
  AND2_X1 U3994 ( .A1(n5922), .A2(n5895), .ZN(n5948) );
  OR2_X1 U3995 ( .A1(n3096), .A2(n5802), .ZN(n5954) );
  OAI21_X1 U3996 ( .B1(n6025), .B2(n6024), .A(n6023), .ZN(n6041) );
  NAND2_X1 U3997 ( .A1(n4414), .A2(n4380), .ZN(n6049) );
  INV_X1 U3998 ( .A(n6065), .ZN(n6109) );
  INV_X1 U3999 ( .A(n6120), .ZN(n6153) );
  AND2_X1 U4000 ( .A1(n6303), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4186) );
  INV_X1 U4001 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6617) );
  NAND2_X1 U4002 ( .A1(n3870), .A2(n6435), .ZN(n6434) );
  NAND2_X1 U4003 ( .A1(n3987), .A2(n3986), .ZN(n3988) );
  INV_X1 U4004 ( .A(n5519), .ZN(n5499) );
  INV_X1 U4005 ( .A(n5517), .ZN(n5449) );
  OAI21_X1 U4006 ( .B1(n4894), .B2(n3983), .A(n4895), .ZN(n5505) );
  OR2_X1 U4007 ( .A1(n4974), .A2(n4973), .ZN(n5107) );
  INV_X1 U4008 ( .A(n5549), .ZN(n5553) );
  NAND2_X1 U4009 ( .A1(n4296), .A2(n5609), .ZN(n5566) );
  INV_X1 U4010 ( .A(n5583), .ZN(n5602) );
  AOI21_X1 U4011 ( .B1(n5233), .B2(n4939), .A(n4820), .ZN(n4821) );
  NAND2_X1 U4012 ( .A1(n5676), .A2(n4191), .ZN(n5673) );
  AOI21_X1 U4013 ( .B1(n5269), .B2(n5764), .A(n5268), .ZN(n5270) );
  INV_X1 U4014 ( .A(n5348), .ZN(n5740) );
  NOR2_X1 U4015 ( .A1(n5347), .A2(n4651), .ZN(n5690) );
  NAND2_X1 U4016 ( .A1(n4647), .A2(n5758), .ZN(n5752) );
  INV_X1 U4017 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U4018 ( .A1(n5803), .A2(n5802), .ZN(n5862) );
  NAND3_X1 U4019 ( .A1(n4415), .A2(n4414), .A3(n6046), .ZN(n5884) );
  INV_X1 U4020 ( .A(n5881), .ZN(n4500) );
  INV_X1 U4021 ( .A(n5918), .ZN(n5898) );
  INV_X1 U4022 ( .A(n5948), .ZN(n5947) );
  OR2_X1 U4023 ( .A1(n6049), .A2(n5954), .ZN(n6004) );
  OR2_X1 U4024 ( .A1(n6049), .A2(n6121), .ZN(n6045) );
  OR2_X1 U4025 ( .A1(n6049), .A2(n6047), .ZN(n6065) );
  NAND2_X1 U4026 ( .A1(n6198), .A2(n6082), .ZN(n6156) );
  OR2_X1 U4027 ( .A1(n6159), .A2(n6158), .ZN(n6208) );
  NAND2_X1 U4028 ( .A1(n6198), .A2(n6046), .ZN(n6258) );
  INV_X1 U4029 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6384) );
  INV_X1 U4030 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6322) );
  INV_X1 U4031 ( .A(n6429), .ZN(n6375) );
  NAND2_X1 U4032 ( .A1(n4197), .A2(n4196), .ZN(U2963) );
  AND2_X2 U4033 ( .A1(n4252), .A2(n3116), .ZN(n3283) );
  AOI22_X1 U4034 ( .A1(n3191), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U4035 ( .A1(n3192), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3112) );
  AND2_X2 U4036 ( .A1(n3109), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3114)
         );
  AND2_X4 U4037 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4681) );
  AND2_X2 U4038 ( .A1(n3114), .A2(n4248), .ZN(n3164) );
  AOI22_X1 U4039 ( .A1(n3175), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3164), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3111) );
  AND2_X2 U4040 ( .A1(n3116), .A2(n4681), .ZN(n3252) );
  AOI22_X1 U4041 ( .A1(n3097), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3110) );
  NAND4_X1 U4042 ( .A1(n3113), .A2(n3112), .A3(n3111), .A4(n3110), .ZN(n3123)
         );
  AND2_X4 U4043 ( .A1(n3114), .A2(n4252), .ZN(n3312) );
  AND2_X4 U4044 ( .A1(n3114), .A2(n3117), .ZN(n3313) );
  AOI22_X1 U4045 ( .A1(n3312), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3121) );
  AOI22_X1 U4046 ( .A1(n3306), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3120) );
  AND2_X2 U4047 ( .A1(n3115), .A2(n3117), .ZN(n3314) );
  AND2_X2 U4048 ( .A1(n3116), .A2(n4248), .ZN(n3425) );
  AOI22_X1 U4049 ( .A1(n3314), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U4050 ( .A1(n3315), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3118) );
  NAND4_X1 U4051 ( .A1(n3121), .A2(n3120), .A3(n3119), .A4(n3118), .ZN(n3122)
         );
  AOI22_X1 U4052 ( .A1(n3191), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U4053 ( .A1(n3314), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U4054 ( .A1(n3098), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U4055 ( .A1(n3312), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3124) );
  NAND4_X1 U4056 ( .A1(n3127), .A2(n3126), .A3(n3125), .A4(n3124), .ZN(n3133)
         );
  AOI22_X1 U4057 ( .A1(n3164), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U4058 ( .A1(n3192), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U4059 ( .A1(n3306), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U4060 ( .A1(n3313), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3128) );
  NAND4_X1 U4061 ( .A1(n3131), .A2(n3130), .A3(n3129), .A4(n3128), .ZN(n3132)
         );
  OR2_X2 U4062 ( .A1(n3133), .A2(n3132), .ZN(n3332) );
  NAND2_X2 U4063 ( .A1(n3231), .A2(n3332), .ZN(n4214) );
  INV_X2 U4064 ( .A(n3332), .ZN(n4485) );
  AOI22_X1 U4065 ( .A1(n3175), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3164), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U4066 ( .A1(n3283), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3136) );
  AOI22_X1 U4067 ( .A1(n3312), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U4068 ( .A1(n3425), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3092), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3134) );
  NAND4_X1 U4069 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3143)
         );
  AOI22_X1 U4070 ( .A1(n3191), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U4071 ( .A1(n3314), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U4072 ( .A1(n3447), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4073 ( .A1(n3313), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3138) );
  NAND4_X1 U4074 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n3142)
         );
  AOI22_X1 U4075 ( .A1(n3175), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3164), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4076 ( .A1(n3191), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4077 ( .A1(n3192), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4078 ( .A1(n3447), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3144) );
  NAND4_X1 U4079 ( .A1(n3147), .A2(n3146), .A3(n3145), .A4(n3144), .ZN(n3153)
         );
  AOI22_X1 U4080 ( .A1(n3312), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4081 ( .A1(n3306), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U4082 ( .A1(n3314), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U4083 ( .A1(n3315), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3148) );
  NAND4_X1 U4084 ( .A1(n3151), .A2(n3150), .A3(n3149), .A4(n3148), .ZN(n3152)
         );
  AND3_X1 U4085 ( .A1(n4214), .A2(n4120), .A3(n4390), .ZN(n3190) );
  AOI22_X1 U4086 ( .A1(n3191), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4087 ( .A1(n3312), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4088 ( .A1(n3305), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3092), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3154) );
  NAND4_X1 U4089 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n3163)
         );
  AOI22_X1 U4090 ( .A1(n3098), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4091 ( .A1(n3192), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4092 ( .A1(n3314), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4093 ( .A1(n3315), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3158) );
  NAND4_X1 U4094 ( .A1(n3161), .A2(n3160), .A3(n3159), .A4(n3158), .ZN(n3162)
         );
  NAND2_X2 U4095 ( .A1(n4485), .A2(n3996), .ZN(n4297) );
  AOI22_X1 U4096 ( .A1(n3175), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3164), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4097 ( .A1(n3191), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U4098 ( .A1(n3192), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4099 ( .A1(n3098), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3165) );
  NAND4_X1 U4100 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3174)
         );
  AOI22_X1 U4101 ( .A1(n3312), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4102 ( .A1(n3306), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3092), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4103 ( .A1(n3314), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4104 ( .A1(n3315), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3169) );
  NAND4_X1 U4105 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3173)
         );
  NAND2_X1 U4106 ( .A1(n4297), .A2(n3990), .ZN(n3228) );
  AOI22_X1 U4107 ( .A1(n3175), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3164), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4108 ( .A1(n3191), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4109 ( .A1(n3192), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4110 ( .A1(n3447), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3176) );
  NAND4_X1 U4111 ( .A1(n3179), .A2(n3178), .A3(n3177), .A4(n3176), .ZN(n3185)
         );
  AOI22_X1 U4112 ( .A1(n3312), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4113 ( .A1(n3306), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4114 ( .A1(n3314), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4115 ( .A1(n3315), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3180) );
  NAND4_X1 U4116 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3184)
         );
  INV_X2 U4117 ( .A(n3878), .ZN(n4279) );
  OAI21_X1 U4118 ( .B1(n4390), .B2(n3332), .A(n4214), .ZN(n3186) );
  INV_X1 U4119 ( .A(n3186), .ZN(n3187) );
  NAND2_X1 U4120 ( .A1(n3187), .A2(n4446), .ZN(n3188) );
  OAI211_X1 U4121 ( .C1(n3190), .C2(n4446), .A(n3189), .B(n3188), .ZN(n3203)
         );
  AOI22_X1 U4122 ( .A1(n3447), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3164), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4123 ( .A1(n3191), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3195) );
  AOI22_X1 U4124 ( .A1(n3313), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4125 ( .A1(n3192), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3193) );
  NAND4_X1 U4126 ( .A1(n3196), .A2(n3195), .A3(n3194), .A4(n3193), .ZN(n3202)
         );
  AOI22_X1 U4127 ( .A1(n3314), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4128 ( .A1(n3283), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4129 ( .A1(n3086), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3092), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U4130 ( .A1(n3312), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3197) );
  NAND4_X1 U4131 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n3197), .ZN(n3201)
         );
  OR2_X4 U4132 ( .A1(n3202), .A2(n3201), .ZN(n3882) );
  NAND2_X1 U4133 ( .A1(n3203), .A2(n4334), .ZN(n3215) );
  NAND2_X1 U4134 ( .A1(n4390), .A2(n3996), .ZN(n3834) );
  NAND2_X1 U4135 ( .A1(n4091), .A2(n5605), .ZN(n3205) );
  INV_X1 U4136 ( .A(n3220), .ZN(n3210) );
  OAI211_X2 U4137 ( .C1(n4297), .C2(n4159), .A(n4301), .B(n4214), .ZN(n4087)
         );
  INV_X1 U4138 ( .A(n4087), .ZN(n3206) );
  NAND2_X1 U4139 ( .A1(n3206), .A2(n3107), .ZN(n3222) );
  NOR2_X1 U4140 ( .A1(n6617), .A2(n6322), .ZN(n6323) );
  AOI21_X1 U4141 ( .B1(n6322), .B2(n6617), .A(n6323), .ZN(n3973) );
  NOR2_X1 U4142 ( .A1(n3878), .A2(n3973), .ZN(n3232) );
  AND2_X2 U4143 ( .A1(n3207), .A2(n3990), .ZN(n3997) );
  OAI21_X1 U4144 ( .B1(n3232), .B2(n3996), .A(n3997), .ZN(n3208) );
  NAND3_X1 U4145 ( .A1(n3215), .A2(n3210), .A3(n3209), .ZN(n3211) );
  AND2_X2 U4146 ( .A1(n3211), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3365) );
  NAND2_X1 U4147 ( .A1(n6431), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3863) );
  MUX2_X1 U4148 ( .A(n3863), .B(n4187), .S(n6113), .Z(n3212) );
  INV_X1 U4149 ( .A(n3215), .ZN(n3216) );
  NAND2_X1 U4150 ( .A1(n4046), .A2(n4390), .ZN(n4117) );
  NAND2_X1 U4151 ( .A1(n3216), .A2(n4117), .ZN(n4111) );
  NOR2_X1 U4152 ( .A1(n3990), .A2(n4116), .ZN(n4213) );
  NAND2_X1 U4153 ( .A1(n4213), .A2(n4334), .ZN(n4112) );
  NAND2_X1 U4154 ( .A1(n3997), .A2(n4297), .ZN(n3217) );
  OAI211_X1 U4155 ( .C1(n4279), .C2(n4116), .A(n3217), .B(n3882), .ZN(n3219)
         );
  OR2_X1 U4156 ( .A1(n6396), .A2(n6303), .ZN(n6306) );
  INV_X1 U4157 ( .A(n6306), .ZN(n3218) );
  OAI211_X1 U4158 ( .C1(n4112), .C2(n4120), .A(n3219), .B(n3218), .ZN(n3221)
         );
  NOR2_X1 U4159 ( .A1(n3221), .A2(n3220), .ZN(n3224) );
  INV_X1 U4160 ( .A(n3990), .ZN(n4586) );
  OAI21_X1 U4161 ( .B1(n3222), .B2(n4586), .A(n3878), .ZN(n3223) );
  NAND2_X2 U4162 ( .A1(n3299), .A2(n3225), .ZN(n3303) );
  INV_X1 U4163 ( .A(n3997), .ZN(n4114) );
  NOR2_X1 U4164 ( .A1(n4114), .A2(n3996), .ZN(n3226) );
  AND2_X1 U4165 ( .A1(n4120), .A2(n4116), .ZN(n3229) );
  NAND3_X1 U4166 ( .A1(n4213), .A2(n5364), .A3(n3231), .ZN(n4241) );
  NAND2_X1 U4167 ( .A1(n3332), .A2(n4301), .ZN(n4299) );
  OAI211_X1 U4168 ( .C1(n6274), .C2(n3232), .A(n4370), .B(n4160), .ZN(n3233)
         );
  NAND2_X1 U4169 ( .A1(n3233), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3239) );
  INV_X1 U4170 ( .A(n3239), .ZN(n3236) );
  XNOR2_X1 U4171 ( .A(n6113), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6160)
         );
  NAND2_X1 U4172 ( .A1(n4187), .A2(n6160), .ZN(n3235) );
  NAND2_X1 U4173 ( .A1(n3863), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4174 ( .A1(n3235), .A2(n3234), .ZN(n3238) );
  NAND2_X1 U4175 ( .A1(n3303), .A2(n3268), .ZN(n3242) );
  INV_X1 U4176 ( .A(n3365), .ZN(n3241) );
  INV_X1 U4177 ( .A(n3238), .ZN(n3240) );
  OAI211_X2 U4178 ( .C1(n3241), .C2(n3237), .A(n3240), .B(n3239), .ZN(n3269)
         );
  NAND2_X1 U4179 ( .A1(n3242), .A2(n3269), .ZN(n3247) );
  AND2_X1 U4180 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3243) );
  NAND2_X1 U4181 ( .A1(n3243), .A2(n6405), .ZN(n6048) );
  INV_X1 U4182 ( .A(n3243), .ZN(n3244) );
  NAND2_X1 U4183 ( .A1(n3244), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3245) );
  INV_X1 U4184 ( .A(n4187), .ZN(n3368) );
  INV_X1 U4185 ( .A(n3863), .ZN(n3367) );
  OAI22_X1 U4186 ( .A1(n4421), .A2(n3368), .B1(n3367), .B2(n6405), .ZN(n3246)
         );
  NAND2_X1 U4187 ( .A1(n3247), .A2(n3248), .ZN(n3251) );
  INV_X1 U4188 ( .A(n3247), .ZN(n3250) );
  NAND2_X2 U4189 ( .A1(n3250), .A2(n3249), .ZN(n3364) );
  NAND2_X1 U4190 ( .A1(n3251), .A2(n3364), .ZN(n4267) );
  AOI22_X1 U4191 ( .A1(n4773), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4192 ( .A1(n3081), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4193 ( .A1(n3080), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3254) );
  BUF_X2 U4194 ( .A(n3252), .Z(n3725) );
  AOI22_X1 U4195 ( .A1(n3098), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3253) );
  NAND4_X1 U4196 ( .A1(n3256), .A2(n3255), .A3(n3254), .A4(n3253), .ZN(n3262)
         );
  AOI22_X1 U4197 ( .A1(n3289), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4198 ( .A1(n4782), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4199 ( .A1(n3797), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4200 ( .A1(n3082), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3257) );
  NAND4_X1 U4201 ( .A1(n3260), .A2(n3259), .A3(n3258), .A4(n3257), .ZN(n3261)
         );
  INV_X1 U4202 ( .A(n3326), .ZN(n3263) );
  INV_X1 U4203 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6552) );
  NOR2_X1 U4204 ( .A1(n3882), .A2(n6303), .ZN(n3282) );
  NAND2_X1 U4205 ( .A1(n3282), .A2(n3264), .ZN(n3265) );
  OAI21_X1 U4206 ( .B1(n3470), .B2(n6552), .A(n3265), .ZN(n3266) );
  NAND2_X1 U4207 ( .A1(n3269), .A2(n3268), .ZN(n3270) );
  XNOR2_X2 U4208 ( .A(n3303), .B(n3270), .ZN(n4239) );
  AOI22_X1 U4209 ( .A1(n3081), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4210 ( .A1(n3080), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4782), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4211 ( .A1(n3289), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4212 ( .A1(n3797), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3271) );
  NAND4_X1 U4213 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3280)
         );
  AOI22_X1 U4214 ( .A1(n4773), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4215 ( .A1(n4774), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4216 ( .A1(n4781), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4217 ( .A1(n3772), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3275) );
  NAND4_X1 U4218 ( .A1(n3278), .A2(n3277), .A3(n3276), .A4(n3275), .ZN(n3279)
         );
  NAND2_X1 U4219 ( .A1(n3326), .A2(n3995), .ZN(n3281) );
  INV_X1 U4221 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3298) );
  NAND2_X1 U4222 ( .A1(n3282), .A2(n3995), .ZN(n3297) );
  AOI22_X1 U4223 ( .A1(n4773), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4224 ( .A1(n4780), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4225 ( .A1(n4772), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4226 ( .A1(n3797), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3284) );
  NAND4_X1 U4227 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3295)
         );
  AOI22_X1 U4228 ( .A1(n3081), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3080), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4229 ( .A1(n3447), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4230 ( .A1(n4782), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4231 ( .A1(n3289), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3290) );
  NAND4_X1 U4232 ( .A1(n3293), .A2(n3292), .A3(n3291), .A4(n3290), .ZN(n3294)
         );
  INV_X1 U4233 ( .A(n4055), .ZN(n4045) );
  NAND2_X1 U4234 ( .A1(n3326), .A2(n4045), .ZN(n3296) );
  OAI211_X1 U4235 ( .C1(n3470), .C2(n3298), .A(n3297), .B(n3296), .ZN(n3334)
         );
  INV_X1 U4236 ( .A(n3299), .ZN(n3301) );
  INV_X1 U4237 ( .A(n5805), .ZN(n3304) );
  AOI22_X1 U4238 ( .A1(n3098), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4239 ( .A1(n3081), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4773), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4240 ( .A1(n4781), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4782), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4241 ( .A1(n3772), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3308) );
  NAND4_X1 U4242 ( .A1(n3311), .A2(n3310), .A3(n3309), .A4(n3308), .ZN(n3321)
         );
  AOI22_X1 U4243 ( .A1(n3289), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4244 ( .A1(n3797), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4245 ( .A1(n4780), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4246 ( .A1(n3080), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3316) );
  NAND4_X1 U4247 ( .A1(n3319), .A2(n3318), .A3(n3317), .A4(n3316), .ZN(n3320)
         );
  NAND2_X1 U4248 ( .A1(n4390), .A2(n4055), .ZN(n3322) );
  OAI211_X1 U4249 ( .C1(n3324), .C2(n3882), .A(n3322), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n3323) );
  AOI21_X1 U4250 ( .B1(n3852), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n3323), 
        .ZN(n3345) );
  XNOR2_X1 U4251 ( .A(n3324), .B(n4055), .ZN(n3325) );
  NAND2_X1 U4252 ( .A1(n3325), .A2(n3326), .ZN(n3344) );
  OR2_X1 U4253 ( .A1(n3345), .A2(n3344), .ZN(n3328) );
  NAND2_X1 U4254 ( .A1(n3326), .A2(n4055), .ZN(n3327) );
  OAI21_X1 U4255 ( .B1(n3337), .B2(n3334), .A(n3335), .ZN(n3331) );
  NAND2_X1 U4256 ( .A1(n3337), .A2(n3334), .ZN(n3330) );
  NAND2_X1 U4257 ( .A1(n3331), .A2(n3330), .ZN(n3394) );
  XNOR2_X1 U4258 ( .A(n3363), .B(n3394), .ZN(n4002) );
  NAND2_X1 U4259 ( .A1(n4002), .A2(n3615), .ZN(n3333) );
  NAND2_X1 U4260 ( .A1(n6550), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3557) );
  NAND2_X1 U4261 ( .A1(n3333), .A2(n3557), .ZN(n3360) );
  NAND2_X1 U4262 ( .A1(n3993), .A2(n3615), .ZN(n3341) );
  AOI22_X1 U4263 ( .A1(n3349), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6550), .ZN(n3339) );
  NOR2_X1 U4264 ( .A1(n4299), .A2(n6550), .ZN(n3413) );
  NAND2_X1 U4265 ( .A1(n3413), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3338) );
  AND2_X1 U4266 ( .A1(n3339), .A2(n3338), .ZN(n3340) );
  OAI21_X1 U4267 ( .B1(n5805), .B2(STATE2_REG_0__SCAN_IN), .A(n3344), .ZN(
        n3343) );
  INV_X1 U4268 ( .A(n4120), .ZN(n3348) );
  INV_X1 U4269 ( .A(n3615), .ZN(n3637) );
  OR2_X1 U4270 ( .A1(n5805), .A2(n3637), .ZN(n3354) );
  INV_X1 U4271 ( .A(n3413), .ZN(n3390) );
  NAND2_X1 U4272 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6550), .ZN(n3351)
         );
  NAND2_X1 U4273 ( .A1(n3349), .A2(EAX_REG_0__SCAN_IN), .ZN(n3350) );
  OAI211_X1 U4274 ( .C1(n3390), .C2(n6260), .A(n3351), .B(n3350), .ZN(n3352)
         );
  INV_X1 U4275 ( .A(n3352), .ZN(n3353) );
  NAND2_X1 U4276 ( .A1(n3354), .A2(n3353), .ZN(n4305) );
  NAND2_X1 U4277 ( .A1(n4306), .A2(n4305), .ZN(n4304) );
  INV_X1 U4278 ( .A(n4305), .ZN(n3355) );
  NAND2_X1 U4279 ( .A1(n3355), .A2(n3079), .ZN(n3356) );
  NAND2_X1 U4280 ( .A1(n4304), .A2(n3356), .ZN(n4218) );
  INV_X1 U4281 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3359) );
  NAND2_X1 U4282 ( .A1(n3413), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3358) );
  OAI21_X1 U4283 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3386), .ZN(n5672) );
  AOI22_X1 U4284 ( .A1(n3079), .A2(n5672), .B1(n4890), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3357) );
  OAI211_X1 U4285 ( .C1(n4723), .C2(n3359), .A(n3358), .B(n3357), .ZN(n4287)
         );
  NAND2_X1 U4286 ( .A1(n4288), .A2(n4287), .ZN(n3362) );
  NAND2_X1 U4287 ( .A1(n3360), .A2(n4221), .ZN(n3361) );
  INV_X1 U4288 ( .A(n3363), .ZN(n3395) );
  NAND2_X1 U4289 ( .A1(n3395), .A2(n3394), .ZN(n3385) );
  NAND2_X1 U4290 ( .A1(n3365), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3371) );
  NAND3_X1 U4291 ( .A1(n6734), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5930) );
  OR2_X1 U4292 ( .A1(n5949), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3366)
         );
  NAND3_X1 U4293 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6204) );
  NOR2_X1 U4294 ( .A1(n6113), .A2(n6204), .ZN(n6252) );
  INV_X1 U4295 ( .A(n6252), .ZN(n6192) );
  NAND2_X1 U4296 ( .A1(n3366), .A2(n6192), .ZN(n5955) );
  OAI22_X1 U4297 ( .A1(n5955), .A2(n3368), .B1(n3367), .B2(n6734), .ZN(n3369)
         );
  INV_X1 U4298 ( .A(n3369), .ZN(n3370) );
  NAND2_X1 U4299 ( .A1(n4349), .A2(n6303), .ZN(n3384) );
  AOI22_X1 U4300 ( .A1(n4773), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4301 ( .A1(n3081), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4302 ( .A1(n3080), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4303 ( .A1(n3098), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3373) );
  NAND4_X1 U4304 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3382)
         );
  AOI22_X1 U4305 ( .A1(n3289), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4306 ( .A1(n4782), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4307 ( .A1(n3797), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4308 ( .A1(n3082), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3377) );
  NAND4_X1 U4309 ( .A1(n3380), .A2(n3379), .A3(n3378), .A4(n3377), .ZN(n3381)
         );
  AOI22_X1 U4310 ( .A1(n3852), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3858), 
        .B2(n4018), .ZN(n3383) );
  XNOR2_X2 U4311 ( .A(n3385), .B(n4379), .ZN(n4380) );
  NAND2_X1 U4312 ( .A1(n4380), .A2(n3615), .ZN(n3393) );
  OAI21_X1 U4313 ( .B1(n3387), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3412), 
        .ZN(n5511) );
  AOI22_X1 U4314 ( .A1(n5511), .A2(n3079), .B1(n4890), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3389) );
  NAND2_X1 U4315 ( .A1(n4797), .A2(EAX_REG_3__SCAN_IN), .ZN(n3388) );
  OAI211_X1 U4316 ( .C1(n3390), .C2(n3109), .A(n3389), .B(n3388), .ZN(n3391)
         );
  INV_X1 U4317 ( .A(n3391), .ZN(n3392) );
  NAND2_X1 U4318 ( .A1(n3393), .A2(n3392), .ZN(n4259) );
  NAND2_X1 U4319 ( .A1(n4258), .A2(n4259), .ZN(n4260) );
  INV_X1 U4320 ( .A(n4260), .ZN(n3420) );
  INV_X1 U4321 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4322 ( .A1(n3097), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4323 ( .A1(n4773), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4324 ( .A1(n3080), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        INSTQUEUE_REG_13__4__SCAN_IN), .B2(n4775), .ZN(n3398) );
  AOI22_X1 U4325 ( .A1(n4782), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        INSTQUEUE_REG_0__4__SCAN_IN), .B2(n4783), .ZN(n3397) );
  NAND4_X1 U4326 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3406)
         );
  AOI22_X1 U4327 ( .A1(n3725), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3081), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4328 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3797), .B1(n4781), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4329 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3082), .B1(
        INSTQUEUE_REG_1__4__SCAN_IN), .B2(n3772), .ZN(n3402) );
  AOI22_X1 U4330 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4772), .B1(n3289), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3401) );
  NAND4_X1 U4331 ( .A1(n3404), .A2(n3403), .A3(n3402), .A4(n3401), .ZN(n3405)
         );
  NOR2_X1 U4332 ( .A1(n3406), .A2(n3405), .ZN(n4026) );
  INV_X1 U4333 ( .A(n4026), .ZN(n3407) );
  NAND2_X1 U4334 ( .A1(n3858), .A2(n3407), .ZN(n3408) );
  INV_X1 U4335 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3411) );
  AOI21_X1 U4336 ( .B1(n3412), .B2(n3411), .A(n3441), .ZN(n4328) );
  AOI22_X1 U4337 ( .A1(n4797), .A2(EAX_REG_4__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6550), .ZN(n3415) );
  NAND2_X1 U4338 ( .A1(n3413), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3414) );
  NAND2_X1 U4339 ( .A1(n3415), .A2(n3414), .ZN(n3416) );
  NAND2_X1 U4340 ( .A1(n3416), .A2(n4795), .ZN(n3417) );
  OAI21_X1 U4341 ( .B1(n4328), .B2(n4795), .A(n3417), .ZN(n3418) );
  AOI21_X1 U4342 ( .B1(n4016), .B2(n3615), .A(n3418), .ZN(n4316) );
  NAND2_X1 U4343 ( .A1(n3420), .A2(n3419), .ZN(n4308) );
  INV_X1 U4344 ( .A(n3438), .ZN(n3433) );
  INV_X1 U4345 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6481) );
  AOI22_X1 U4346 ( .A1(n4773), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4347 ( .A1(n3081), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4348 ( .A1(n3080), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4349 ( .A1(n3447), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3421) );
  NAND4_X1 U4350 ( .A1(n3424), .A2(n3423), .A3(n3422), .A4(n3421), .ZN(n3431)
         );
  AOI22_X1 U4351 ( .A1(n3289), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4352 ( .A1(n4782), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4353 ( .A1(n3797), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4354 ( .A1(n3082), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3426) );
  NAND4_X1 U4355 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n3430)
         );
  NAND2_X1 U4356 ( .A1(n3858), .A2(n4035), .ZN(n3432) );
  OAI21_X1 U4357 ( .B1(n3470), .B2(n6481), .A(n3432), .ZN(n3435) );
  AOI21_X1 U4358 ( .B1(n3433), .B2(n3436), .A(n3435), .ZN(n3434) );
  INV_X1 U4359 ( .A(n3434), .ZN(n3440) );
  NAND2_X1 U4360 ( .A1(n3436), .A2(n3435), .ZN(n3437) );
  INV_X1 U4361 ( .A(n3472), .ZN(n3439) );
  INV_X1 U4362 ( .A(n4029), .ZN(n3446) );
  INV_X1 U4363 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3444) );
  OAI21_X1 U4364 ( .B1(n3441), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3463), 
        .ZN(n5481) );
  NAND2_X1 U4365 ( .A1(n5481), .A2(n3079), .ZN(n3443) );
  NAND2_X1 U4366 ( .A1(n4890), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3442)
         );
  OAI211_X1 U4367 ( .C1(n4723), .C2(n3444), .A(n3443), .B(n3442), .ZN(n3445)
         );
  NOR2_X2 U4368 ( .A1(n4308), .A2(n4309), .ZN(n4310) );
  INV_X1 U4369 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4370 ( .A1(n3097), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4371 ( .A1(n4773), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4372 ( .A1(n4781), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4373 ( .A1(n3772), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4374 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3457)
         );
  AOI22_X1 U4375 ( .A1(n3725), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3081), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4376 ( .A1(n3080), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4377 ( .A1(n4782), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4378 ( .A1(n4783), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4379 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3456)
         );
  INV_X1 U4380 ( .A(n4044), .ZN(n3458) );
  NAND2_X1 U4381 ( .A1(n3858), .A2(n3458), .ZN(n3459) );
  OAI21_X1 U4382 ( .B1(n3470), .B2(n3460), .A(n3459), .ZN(n3471) );
  OR2_X1 U4383 ( .A1(n3472), .A2(n3471), .ZN(n4034) );
  NAND2_X1 U4384 ( .A1(n4034), .A2(n3615), .ZN(n3467) );
  INV_X1 U4385 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3462) );
  INV_X1 U4386 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6164) );
  OAI21_X1 U4387 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6164), .A(n6550), 
        .ZN(n3461) );
  OAI21_X1 U4388 ( .B1(n4723), .B2(n3462), .A(n3461), .ZN(n3465) );
  AOI21_X1 U4389 ( .B1(n6711), .B2(n3463), .A(n3474), .ZN(n5464) );
  NAND2_X1 U4390 ( .A1(n5464), .A2(n3079), .ZN(n3464) );
  NAND2_X1 U4391 ( .A1(n3465), .A2(n3464), .ZN(n3466) );
  NAND2_X1 U4392 ( .A1(n3467), .A2(n3466), .ZN(n4404) );
  AND2_X2 U4393 ( .A1(n4310), .A2(n4404), .ZN(n4403) );
  INV_X1 U4394 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U4395 ( .A1(n3858), .A2(n4055), .ZN(n3468) );
  OAI21_X1 U4396 ( .B1(n3470), .B2(n3469), .A(n3468), .ZN(n3473) );
  XNOR2_X1 U4397 ( .A(n3473), .B(n4054), .ZN(n4047) );
  NAND2_X1 U4398 ( .A1(n4047), .A2(n3615), .ZN(n3478) );
  OAI21_X1 U4399 ( .B1(n3474), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3492), 
        .ZN(n5451) );
  NAND2_X1 U4400 ( .A1(n5451), .A2(n3079), .ZN(n3476) );
  AOI22_X1 U4401 ( .A1(n4797), .A2(EAX_REG_7__SCAN_IN), .B1(n4890), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3475) );
  AND2_X1 U4402 ( .A1(n3476), .A2(n3475), .ZN(n3477) );
  NAND2_X1 U4403 ( .A1(n3478), .A2(n3477), .ZN(n4429) );
  AND2_X2 U4404 ( .A1(n4403), .A2(n4429), .ZN(n4428) );
  XNOR2_X1 U4405 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3492), .ZN(n5441) );
  AOI22_X1 U4406 ( .A1(n3081), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4407 ( .A1(n3080), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4408 ( .A1(n4772), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4409 ( .A1(n3797), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3479) );
  NAND4_X1 U4410 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3488)
         );
  AOI22_X1 U4411 ( .A1(n4773), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4412 ( .A1(n3098), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4413 ( .A1(n4782), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4414 ( .A1(n3289), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3483) );
  NAND4_X1 U4415 ( .A1(n3486), .A2(n3485), .A3(n3484), .A4(n3483), .ZN(n3487)
         );
  OR2_X1 U4416 ( .A1(n3488), .A2(n3487), .ZN(n3489) );
  AOI22_X1 U4417 ( .A1(n3615), .A2(n3489), .B1(n4890), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3491) );
  NAND2_X1 U4418 ( .A1(n4797), .A2(EAX_REG_8__SCAN_IN), .ZN(n3490) );
  OAI211_X1 U4419 ( .C1(n5441), .C2(n4795), .A(n3491), .B(n3490), .ZN(n4456)
         );
  NAND2_X1 U4420 ( .A1(n3494), .A2(n6638), .ZN(n3496) );
  INV_X1 U4421 ( .A(n3536), .ZN(n3495) );
  NAND2_X1 U4422 ( .A1(n3496), .A2(n3495), .ZN(n5434) );
  AOI22_X1 U4423 ( .A1(n4773), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4424 ( .A1(n3080), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4425 ( .A1(n4772), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4426 ( .A1(n3772), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4427 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3506)
         );
  AOI22_X1 U4428 ( .A1(n3081), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4429 ( .A1(n3797), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4782), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4430 ( .A1(n3447), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U4431 ( .A1(n3289), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3501) );
  NAND4_X1 U4432 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3505)
         );
  OAI21_X1 U4433 ( .B1(n3506), .B2(n3505), .A(n3615), .ZN(n3508) );
  NAND2_X1 U4434 ( .A1(n4797), .A2(EAX_REG_9__SCAN_IN), .ZN(n3507) );
  OAI211_X1 U4435 ( .C1(n3557), .C2(n6638), .A(n3508), .B(n3507), .ZN(n3509)
         );
  AOI21_X1 U4436 ( .B1(n5434), .B2(n3079), .A(n3509), .ZN(n4514) );
  AOI22_X1 U4437 ( .A1(n4773), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4438 ( .A1(n3080), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4439 ( .A1(n3097), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4440 ( .A1(n3797), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3512) );
  NAND4_X1 U4441 ( .A1(n3515), .A2(n3514), .A3(n3513), .A4(n3512), .ZN(n3521)
         );
  AOI22_X1 U4442 ( .A1(n3289), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4443 ( .A1(n3081), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4444 ( .A1(n4782), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4445 ( .A1(n3082), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3516) );
  NAND4_X1 U4446 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3520)
         );
  OAI21_X1 U4447 ( .B1(n3521), .B2(n3520), .A(n3615), .ZN(n3525) );
  NAND2_X1 U4448 ( .A1(n4797), .A2(EAX_REG_10__SCAN_IN), .ZN(n3524) );
  XOR2_X1 U4449 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3536), .Z(n5428) );
  INV_X1 U4450 ( .A(n5428), .ZN(n3522) );
  AOI22_X1 U4451 ( .A1(n4890), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n3079), 
        .B2(n3522), .ZN(n3523) );
  NOR2_X2 U4452 ( .A1(n4513), .A2(n4600), .ZN(n4598) );
  AOI22_X1 U4453 ( .A1(n3081), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4773), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4454 ( .A1(n3080), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4455 ( .A1(n3797), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4456 ( .A1(n3289), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3526) );
  NAND4_X1 U4457 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(n3535)
         );
  AOI22_X1 U4458 ( .A1(n4774), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4459 ( .A1(n3447), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4460 ( .A1(n4772), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4461 ( .A1(n4782), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3530) );
  NAND4_X1 U4462 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(n3534)
         );
  NOR2_X1 U4463 ( .A1(n3535), .A2(n3534), .ZN(n3540) );
  INV_X1 U4464 ( .A(n3542), .ZN(n3537) );
  XNOR2_X1 U4465 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3537), .ZN(n4632)
         );
  AOI22_X1 U4466 ( .A1(n3079), .A2(n4632), .B1(n4890), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3539) );
  NAND2_X1 U4467 ( .A1(n4797), .A2(EAX_REG_11__SCAN_IN), .ZN(n3538) );
  OAI211_X1 U4468 ( .C1(n3637), .C2(n3540), .A(n3539), .B(n3538), .ZN(n4608)
         );
  AND2_X2 U4469 ( .A1(n4598), .A2(n4608), .ZN(n4623) );
  XOR2_X1 U4470 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3556), .Z(n5417) );
  AOI22_X1 U4471 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3289), .B1(n4772), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4472 ( .A1(n4773), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4473 ( .A1(n3080), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4474 ( .A1(n4782), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3543) );
  NAND4_X1 U4475 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3552)
         );
  AOI22_X1 U4476 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3081), .B1(n3797), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4477 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4780), .B1(n4774), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4478 ( .A1(n3097), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4479 ( .A1(n3082), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3547) );
  NAND4_X1 U4480 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(n3551)
         );
  OR2_X1 U4481 ( .A1(n3552), .A2(n3551), .ZN(n3553) );
  AOI22_X1 U4482 ( .A1(n3615), .A2(n3553), .B1(n4890), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3555) );
  NAND2_X1 U4483 ( .A1(n4797), .A2(EAX_REG_12__SCAN_IN), .ZN(n3554) );
  OAI211_X1 U4484 ( .C1(n5417), .C2(n4795), .A(n3555), .B(n3554), .ZN(n4622)
         );
  XNOR2_X1 U4485 ( .A(n3588), .B(n3587), .ZN(n5407) );
  INV_X1 U4486 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6562) );
  OAI22_X1 U4487 ( .A1(n4723), .A2(n6562), .B1(n3557), .B2(n3587), .ZN(n3558)
         );
  AOI21_X1 U4488 ( .B1(n5407), .B2(n3079), .A(n3558), .ZN(n3570) );
  AOI22_X1 U4489 ( .A1(n4773), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4490 ( .A1(n3081), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4491 ( .A1(n3080), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4492 ( .A1(n3098), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3559) );
  NAND4_X1 U4493 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3568)
         );
  AOI22_X1 U4494 ( .A1(n3289), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4495 ( .A1(n4782), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4496 ( .A1(n3797), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4497 ( .A1(n3082), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4498 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3567)
         );
  OR2_X1 U4499 ( .A1(n3568), .A2(n3567), .ZN(n3569) );
  NAND2_X1 U4500 ( .A1(n3615), .A2(n3569), .ZN(n4672) );
  NAND2_X1 U4501 ( .A1(n4159), .A2(n3996), .ZN(n3572) );
  AOI22_X1 U4502 ( .A1(n3447), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4503 ( .A1(n3312), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4504 ( .A1(n4773), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3080), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4505 ( .A1(n3772), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3573) );
  NAND4_X1 U4506 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3582)
         );
  AOI22_X1 U4507 ( .A1(n3081), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4508 ( .A1(n3797), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4509 ( .A1(n4780), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4510 ( .A1(n4782), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3577) );
  NAND4_X1 U4511 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3581)
         );
  NOR2_X1 U4512 ( .A1(n3582), .A2(n3581), .ZN(n3586) );
  OAI21_X1 U4513 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6164), .A(n6550), 
        .ZN(n3583) );
  INV_X1 U4514 ( .A(n3583), .ZN(n3584) );
  AOI21_X1 U4515 ( .B1(n4797), .B2(EAX_REG_17__SCAN_IN), .A(n3584), .ZN(n3585)
         );
  OAI21_X1 U4516 ( .B1(n4767), .B2(n3586), .A(n3585), .ZN(n3591) );
  OAI21_X1 U4517 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3589), .A(n3657), 
        .ZN(n5392) );
  OR2_X1 U4518 ( .A1(n4795), .A2(n5392), .ZN(n3590) );
  AND2_X1 U4519 ( .A1(n3591), .A2(n3590), .ZN(n5229) );
  XNOR2_X1 U4520 ( .A(n3605), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5040)
         );
  AOI22_X1 U4521 ( .A1(n3098), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4522 ( .A1(n4781), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4782), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4523 ( .A1(n3797), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4524 ( .A1(n4772), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3592) );
  NAND4_X1 U4525 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3601)
         );
  AOI22_X1 U4526 ( .A1(n3081), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4773), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4527 ( .A1(n4774), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4528 ( .A1(n3289), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4529 ( .A1(n3080), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3596) );
  NAND4_X1 U4530 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3600)
         );
  NOR2_X1 U4531 ( .A1(n3601), .A2(n3600), .ZN(n3603) );
  AOI22_X1 U4532 ( .A1(n4797), .A2(EAX_REG_16__SCAN_IN), .B1(n4890), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3602) );
  OAI21_X1 U4533 ( .B1(n4767), .B2(n3603), .A(n3602), .ZN(n3604) );
  AOI21_X1 U4534 ( .B1(n5040), .B2(n3079), .A(n3604), .ZN(n4950) );
  AOI21_X1 U4535 ( .B1(n6571), .B2(n3606), .A(n3605), .ZN(n5402) );
  OR2_X1 U4536 ( .A1(n5402), .A2(n4795), .ZN(n3622) );
  AOI22_X1 U4537 ( .A1(n3081), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4782), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4538 ( .A1(n3289), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4539 ( .A1(n3797), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4540 ( .A1(n4773), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3607) );
  NAND4_X1 U4541 ( .A1(n3610), .A2(n3609), .A3(n3608), .A4(n3607), .ZN(n3617)
         );
  AOI22_X1 U4542 ( .A1(n3097), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4543 ( .A1(n4780), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4544 ( .A1(n3080), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4545 ( .A1(n3772), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3611) );
  NAND4_X1 U4546 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(n3616)
         );
  OAI21_X1 U4547 ( .B1(n3617), .B2(n3616), .A(n3615), .ZN(n3620) );
  NAND2_X1 U4548 ( .A1(n3349), .A2(EAX_REG_15__SCAN_IN), .ZN(n3619) );
  NAND2_X1 U4549 ( .A1(n4890), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3618)
         );
  AND3_X1 U4550 ( .A1(n3620), .A2(n3619), .A3(n3618), .ZN(n3621) );
  NOR2_X1 U4551 ( .A1(n4950), .A2(n5007), .ZN(n4948) );
  AND2_X1 U4552 ( .A1(n5229), .A2(n4948), .ZN(n3638) );
  AOI22_X1 U4553 ( .A1(n4774), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4554 ( .A1(n4781), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4782), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4555 ( .A1(n3289), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4556 ( .A1(n3797), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3623) );
  NAND4_X1 U4557 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3632)
         );
  AOI22_X1 U4558 ( .A1(n3081), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4773), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4559 ( .A1(n3097), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4560 ( .A1(n3080), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4561 ( .A1(n3772), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3627) );
  NAND4_X1 U4562 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3631)
         );
  NOR2_X1 U4563 ( .A1(n3632), .A2(n3631), .ZN(n3636) );
  XNOR2_X1 U4564 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3633), .ZN(n5059)
         );
  AOI22_X1 U4565 ( .A1(n3079), .A2(n5059), .B1(n4890), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3635) );
  NAND2_X1 U4566 ( .A1(n3349), .A2(EAX_REG_14__SCAN_IN), .ZN(n3634) );
  OAI211_X1 U4567 ( .C1(n3637), .C2(n3636), .A(n3635), .B(n3634), .ZN(n4946)
         );
  AOI22_X1 U4568 ( .A1(n3081), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4569 ( .A1(n3289), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4570 ( .A1(n3097), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4571 ( .A1(n3082), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3640) );
  NAND4_X1 U4572 ( .A1(n3643), .A2(n3642), .A3(n3641), .A4(n3640), .ZN(n3649)
         );
  AOI22_X1 U4573 ( .A1(n4780), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4574 ( .A1(n4773), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4575 ( .A1(n3080), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4576 ( .A1(n4782), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3644) );
  NAND4_X1 U4577 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3648)
         );
  NOR2_X1 U4578 ( .A1(n3649), .A2(n3648), .ZN(n3653) );
  NAND2_X1 U4579 ( .A1(n6550), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3650)
         );
  NAND2_X1 U4580 ( .A1(n4795), .A2(n3650), .ZN(n3651) );
  AOI21_X1 U4581 ( .B1(n4797), .B2(EAX_REG_18__SCAN_IN), .A(n3651), .ZN(n3652)
         );
  OAI21_X1 U4582 ( .B1(n4767), .B2(n3653), .A(n3652), .ZN(n3655) );
  XNOR2_X1 U4583 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3657), .ZN(n4939)
         );
  NAND2_X1 U4584 ( .A1(n3079), .A2(n4939), .ZN(n3654) );
  NAND2_X1 U4585 ( .A1(n3655), .A2(n3654), .ZN(n4804) );
  OR2_X2 U4586 ( .A1(n5232), .A2(n4804), .ZN(n5157) );
  INV_X1 U4587 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3656) );
  OR2_X1 U4588 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3659)
         );
  NAND2_X1 U4589 ( .A1(n3659), .A2(n3687), .ZN(n5223) );
  AOI22_X1 U4590 ( .A1(n3081), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4591 ( .A1(n3289), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4592 ( .A1(n3797), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4782), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4593 ( .A1(n4774), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3660) );
  NAND4_X1 U4594 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3669)
         );
  AOI22_X1 U4595 ( .A1(n3097), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4773), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4596 ( .A1(n3080), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4597 ( .A1(n3772), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4598 ( .A1(n3082), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3664) );
  NAND4_X1 U4599 ( .A1(n3667), .A2(n3666), .A3(n3665), .A4(n3664), .ZN(n3668)
         );
  NOR2_X1 U4600 ( .A1(n3669), .A2(n3668), .ZN(n3672) );
  OAI21_X1 U4601 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6164), .A(n6550), 
        .ZN(n3671) );
  NAND2_X1 U4602 ( .A1(n3349), .A2(EAX_REG_19__SCAN_IN), .ZN(n3670) );
  OAI211_X1 U4603 ( .C1(n4767), .C2(n3672), .A(n3671), .B(n3670), .ZN(n3673)
         );
  OAI21_X1 U4604 ( .B1(n5223), .B2(n4795), .A(n3673), .ZN(n5156) );
  NOR2_X4 U4605 ( .A1(n5157), .A2(n5156), .ZN(n5158) );
  AOI22_X1 U4606 ( .A1(n4773), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4607 ( .A1(n3081), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4608 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3080), .B1(n4781), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4609 ( .A1(n3447), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3674) );
  NAND4_X1 U4610 ( .A1(n3677), .A2(n3676), .A3(n3675), .A4(n3674), .ZN(n3683)
         );
  AOI22_X1 U4611 ( .A1(n3312), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4612 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4782), .B1(n4775), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4613 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3797), .B1(n3772), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4614 ( .A1(n3082), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3678) );
  NAND4_X1 U4615 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3682)
         );
  NOR2_X1 U4616 ( .A1(n3683), .A2(n3682), .ZN(n3686) );
  AOI21_X1 U4617 ( .B1(n4797), .B2(EAX_REG_20__SCAN_IN), .A(n3684), .ZN(n3685)
         );
  OAI21_X1 U4618 ( .B1(n4767), .B2(n3686), .A(n3685), .ZN(n3689) );
  AOI21_X1 U4619 ( .B1(n6633), .B2(n3687), .A(n3704), .ZN(n5141) );
  NAND2_X1 U4620 ( .A1(n5141), .A2(n3079), .ZN(n3688) );
  AOI22_X1 U4622 ( .A1(n3797), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4623 ( .A1(n4773), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4624 ( .A1(n3097), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4625 ( .A1(n4782), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3690) );
  NAND4_X1 U4626 ( .A1(n3693), .A2(n3692), .A3(n3691), .A4(n3690), .ZN(n3699)
         );
  AOI22_X1 U4627 ( .A1(n3081), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4628 ( .A1(n3080), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4629 ( .A1(n3082), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4630 ( .A1(n3289), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3694) );
  NAND4_X1 U4631 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3698)
         );
  NOR2_X1 U4632 ( .A1(n3699), .A2(n3698), .ZN(n3703) );
  NAND2_X1 U4633 ( .A1(n6550), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3700)
         );
  NAND2_X1 U4634 ( .A1(n4795), .A2(n3700), .ZN(n3701) );
  AOI21_X1 U4635 ( .B1(n4797), .B2(EAX_REG_21__SCAN_IN), .A(n3701), .ZN(n3702)
         );
  OAI21_X1 U4636 ( .B1(n4767), .B2(n3703), .A(n3702), .ZN(n3706) );
  OAI21_X1 U4637 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n3704), .A(n3724), 
        .ZN(n5214) );
  OR2_X1 U4638 ( .A1(n4795), .A2(n5214), .ZN(n3705) );
  AOI22_X1 U4639 ( .A1(n3080), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4640 ( .A1(n4772), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4641 ( .A1(n3081), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4642 ( .A1(n3797), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3707) );
  NAND4_X1 U4643 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3716)
         );
  AOI22_X1 U4644 ( .A1(n3447), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4645 ( .A1(n4773), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4646 ( .A1(n4782), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4647 ( .A1(n3312), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3711) );
  NAND4_X1 U4648 ( .A1(n3714), .A2(n3713), .A3(n3712), .A4(n3711), .ZN(n3715)
         );
  NOR2_X1 U4649 ( .A1(n3716), .A2(n3715), .ZN(n3720) );
  NAND2_X1 U4650 ( .A1(n6550), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3717)
         );
  NAND2_X1 U4651 ( .A1(n4795), .A2(n3717), .ZN(n3718) );
  AOI21_X1 U4652 ( .B1(n4797), .B2(EAX_REG_22__SCAN_IN), .A(n3718), .ZN(n3719)
         );
  OAI21_X1 U4653 ( .B1(n4767), .B2(n3720), .A(n3719), .ZN(n3722) );
  XNOR2_X1 U4654 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .B(n3724), .ZN(n5122)
         );
  NAND2_X1 U4655 ( .A1(n5122), .A2(n3079), .ZN(n3721) );
  NAND2_X1 U4656 ( .A1(n3722), .A2(n3721), .ZN(n4841) );
  NOR2_X2 U4657 ( .A1(n5138), .A2(n4841), .ZN(n4182) );
  INV_X1 U4658 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3723) );
  XNOR2_X1 U4659 ( .A(n3770), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5027)
         );
  AOI22_X1 U4660 ( .A1(n4773), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4661 ( .A1(n3289), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4662 ( .A1(n3098), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4663 ( .A1(n3081), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3726) );
  NAND4_X1 U4664 ( .A1(n3729), .A2(n3728), .A3(n3727), .A4(n3726), .ZN(n3735)
         );
  AOI22_X1 U4665 ( .A1(n4780), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4666 ( .A1(n3797), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4782), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4667 ( .A1(n3080), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4668 ( .A1(n4772), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3730) );
  NAND4_X1 U4669 ( .A1(n3733), .A2(n3732), .A3(n3731), .A4(n3730), .ZN(n3734)
         );
  NOR2_X1 U4670 ( .A1(n3735), .A2(n3734), .ZN(n3762) );
  AOI22_X1 U4671 ( .A1(n4773), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4672 ( .A1(n3081), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3080), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4673 ( .A1(n4774), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4674 ( .A1(n4782), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4675 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3745)
         );
  AOI22_X1 U4676 ( .A1(n3289), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4677 ( .A1(n3447), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4678 ( .A1(n3797), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4679 ( .A1(n3082), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3740) );
  NAND4_X1 U4680 ( .A1(n3743), .A2(n3742), .A3(n3741), .A4(n3740), .ZN(n3744)
         );
  NOR2_X1 U4681 ( .A1(n3745), .A2(n3744), .ZN(n3763) );
  NOR2_X1 U4682 ( .A1(n3762), .A2(n3763), .ZN(n3784) );
  AOI22_X1 U4683 ( .A1(n4773), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4684 ( .A1(n3081), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4685 ( .A1(n3080), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4686 ( .A1(n3447), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3746) );
  NAND4_X1 U4687 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3755)
         );
  AOI22_X1 U4688 ( .A1(n3289), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4689 ( .A1(n4782), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4690 ( .A1(n3797), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4691 ( .A1(n3082), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4692 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3754)
         );
  OR2_X1 U4693 ( .A1(n3755), .A2(n3754), .ZN(n3783) );
  XNOR2_X1 U4694 ( .A(n3784), .B(n3783), .ZN(n3757) );
  AOI22_X1 U4695 ( .A1(n3349), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4890), .ZN(n3756) );
  OAI21_X1 U4696 ( .B1(n3757), .B2(n4767), .A(n3756), .ZN(n3758) );
  AOI21_X1 U4697 ( .B1(n5027), .B2(n3079), .A(n3758), .ZN(n4199) );
  INV_X1 U4698 ( .A(n3770), .ZN(n3761) );
  OR2_X1 U4699 ( .A1(n3759), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3760)
         );
  NAND2_X1 U4700 ( .A1(n3761), .A2(n3760), .ZN(n5110) );
  XNOR2_X1 U4701 ( .A(n3763), .B(n3762), .ZN(n3764) );
  NOR2_X1 U4702 ( .A1(n4767), .A2(n3764), .ZN(n3768) );
  INV_X1 U4703 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3766) );
  NAND2_X1 U4704 ( .A1(n6550), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3765)
         );
  OAI211_X1 U4705 ( .C1(n4723), .C2(n3766), .A(n4795), .B(n3765), .ZN(n3767)
         );
  OAI22_X1 U4706 ( .A1(n5110), .A2(n4795), .B1(n3768), .B2(n3767), .ZN(n4184)
         );
  OR2_X1 U4707 ( .A1(n4199), .A2(n4184), .ZN(n3810) );
  AND2_X2 U4708 ( .A1(n4182), .A2(n3769), .ZN(n4921) );
  OAI21_X1 U4709 ( .B1(n3771), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n3874), 
        .ZN(n5210) );
  OR2_X1 U4710 ( .A1(n5210), .A2(n4795), .ZN(n3790) );
  AOI22_X1 U4711 ( .A1(n3081), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4712 ( .A1(n4773), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4713 ( .A1(n3772), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4714 ( .A1(n4772), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3773) );
  NAND4_X1 U4715 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3782)
         );
  AOI22_X1 U4716 ( .A1(n3098), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4717 ( .A1(n4780), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3080), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4718 ( .A1(n3797), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4782), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4719 ( .A1(n3312), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3082), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4720 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3781)
         );
  NOR2_X1 U4721 ( .A1(n3782), .A2(n3781), .ZN(n3792) );
  NAND2_X1 U4722 ( .A1(n3784), .A2(n3783), .ZN(n3791) );
  XNOR2_X1 U4723 ( .A(n3792), .B(n3791), .ZN(n3788) );
  NAND2_X1 U4724 ( .A1(n6550), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3785)
         );
  NAND2_X1 U4725 ( .A1(n4795), .A2(n3785), .ZN(n3786) );
  AOI21_X1 U4726 ( .B1(n4797), .B2(EAX_REG_25__SCAN_IN), .A(n3786), .ZN(n3787)
         );
  OAI21_X1 U4727 ( .B1(n3788), .B2(n4767), .A(n3787), .ZN(n3789) );
  NAND2_X1 U4728 ( .A1(n4921), .A2(n4920), .ZN(n4922) );
  INV_X1 U4729 ( .A(n4922), .ZN(n3815) );
  NOR2_X1 U4730 ( .A1(n3792), .A2(n3791), .ZN(n4719) );
  AOI22_X1 U4731 ( .A1(n4773), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4732 ( .A1(n3081), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4733 ( .A1(n3080), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4734 ( .A1(n3098), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3793) );
  NAND4_X1 U4735 ( .A1(n3796), .A2(n3795), .A3(n3794), .A4(n3793), .ZN(n3803)
         );
  AOI22_X1 U4736 ( .A1(n3312), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4737 ( .A1(n4782), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4738 ( .A1(n3797), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4739 ( .A1(n3082), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3798) );
  NAND4_X1 U4740 ( .A1(n3801), .A2(n3800), .A3(n3799), .A4(n3798), .ZN(n3802)
         );
  OR2_X1 U4741 ( .A1(n3803), .A2(n3802), .ZN(n4718) );
  XNOR2_X1 U4742 ( .A(n4719), .B(n4718), .ZN(n3807) );
  NAND2_X1 U4743 ( .A1(n6550), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3804)
         );
  NAND2_X1 U4744 ( .A1(n4795), .A2(n3804), .ZN(n3805) );
  AOI21_X1 U4745 ( .B1(n4797), .B2(EAX_REG_26__SCAN_IN), .A(n3805), .ZN(n3806)
         );
  OAI21_X1 U4746 ( .B1(n3807), .B2(n4767), .A(n3806), .ZN(n3809) );
  XNOR2_X1 U4747 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n3874), .ZN(n4863)
         );
  NAND2_X1 U4748 ( .A1(n4863), .A2(n3079), .ZN(n3808) );
  AND2_X1 U4749 ( .A1(n5136), .A2(n5135), .ZN(n3813) );
  OR2_X1 U4750 ( .A1(n3810), .A2(n4841), .ZN(n3812) );
  NAND2_X1 U4751 ( .A1(n3814), .A2(n4920), .ZN(n3811) );
  NOR2_X1 U4752 ( .A1(n3812), .A2(n3811), .ZN(n4726) );
  NAND2_X1 U4753 ( .A1(n3813), .A2(n4726), .ZN(n4972) );
  XNOR2_X1 U4754 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3831) );
  NAND2_X1 U4755 ( .A1(n3831), .A2(n3830), .ZN(n3829) );
  NAND2_X1 U4756 ( .A1(n6667), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3816) );
  NAND2_X1 U4757 ( .A1(n3829), .A2(n3816), .ZN(n3825) );
  XNOR2_X1 U4758 ( .A(n4686), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3824)
         );
  INV_X1 U4759 ( .A(n3824), .ZN(n3817) );
  NAND2_X1 U4760 ( .A1(n3825), .A2(n3817), .ZN(n3819) );
  NAND2_X1 U4761 ( .A1(n6405), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U4762 ( .A1(n3819), .A2(n3818), .ZN(n3828) );
  INV_X1 U4763 ( .A(n3828), .ZN(n3820) );
  OAI222_X1 U4764 ( .A1(n6586), .A2(n3822), .B1(n6586), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3822), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3869) );
  NAND2_X1 U4765 ( .A1(n3822), .A2(n6586), .ZN(n3823) );
  XNOR2_X1 U4766 ( .A(n3825), .B(n3824), .ZN(n3866) );
  INV_X1 U4767 ( .A(n3845), .ZN(n3851) );
  AND2_X1 U4768 ( .A1(n4279), .A2(n3996), .ZN(n3826) );
  INV_X1 U4769 ( .A(n4046), .ZN(n4028) );
  XNOR2_X1 U4770 ( .A(n3828), .B(n3827), .ZN(n3864) );
  INV_X1 U4771 ( .A(n3858), .ZN(n3832) );
  OAI21_X1 U4772 ( .B1(n3832), .B2(n4279), .A(n3996), .ZN(n3840) );
  OAI21_X1 U4773 ( .B1(n3831), .B2(n3830), .A(n3829), .ZN(n3841) );
  INV_X1 U4774 ( .A(n3841), .ZN(n3865) );
  XNOR2_X1 U4775 ( .A(n6260), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3835)
         );
  NOR2_X1 U4776 ( .A1(n3832), .A2(n3835), .ZN(n3833) );
  OAI21_X1 U4777 ( .B1(n3840), .B2(n3865), .A(n3833), .ZN(n3839) );
  INV_X1 U4778 ( .A(n3834), .ZN(n4104) );
  OAI21_X1 U4779 ( .B1(n4104), .B2(n3835), .A(n3882), .ZN(n3836) );
  OAI211_X1 U4780 ( .C1(n3859), .C2(n3865), .A(n3850), .B(n3836), .ZN(n3837)
         );
  INV_X1 U4781 ( .A(n3837), .ZN(n3838) );
  AOI21_X1 U4782 ( .B1(n3859), .B2(n3839), .A(n3838), .ZN(n3844) );
  INV_X1 U4783 ( .A(n3840), .ZN(n3842) );
  NOR3_X1 U4784 ( .A1(n3842), .A2(n6303), .A3(n3841), .ZN(n3843) );
  NOR2_X1 U4785 ( .A1(n3844), .A2(n3843), .ZN(n3849) );
  INV_X1 U4786 ( .A(n3866), .ZN(n3847) );
  INV_X1 U4787 ( .A(n3850), .ZN(n3846) );
  AOI211_X1 U4788 ( .C1(n3852), .C2(n3847), .A(n3846), .B(n3845), .ZN(n3848)
         );
  OAI222_X1 U4789 ( .A1(n3851), .A2(n3850), .B1(n4028), .B2(n3864), .C1(n3849), 
        .C2(n3848), .ZN(n3855) );
  AOI21_X1 U4790 ( .B1(n3867), .B2(n3864), .A(n3852), .ZN(n3853) );
  INV_X1 U4791 ( .A(n3853), .ZN(n3854) );
  AOI22_X1 U4792 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6303), .B1(n3855), .B2(n3854), .ZN(n3856) );
  INV_X1 U4793 ( .A(n3859), .ZN(n3860) );
  INV_X1 U4794 ( .A(n6274), .ZN(n5363) );
  AND3_X1 U4795 ( .A1(n3866), .A2(n3865), .A3(n3864), .ZN(n3868) );
  OAI21_X1 U4796 ( .B1(n3869), .B2(n3868), .A(n3867), .ZN(n4095) );
  NAND2_X1 U4797 ( .A1(n4126), .A2(n4334), .ZN(n4093) );
  INV_X1 U4798 ( .A(n4093), .ZN(n6276) );
  NAND2_X1 U4799 ( .A1(n6550), .A2(n6431), .ZN(n6311) );
  NOR3_X1 U4800 ( .A1(n6303), .A2(n6384), .A3(n6311), .ZN(n6298) );
  AND2_X2 U4801 ( .A1(n4187), .A2(n6550), .ZN(n5348) );
  AND2_X1 U4802 ( .A1(n4186), .A2(n3079), .ZN(n6307) );
  OR2_X1 U4803 ( .A1(n5348), .A2(n6307), .ZN(n3871) );
  INV_X1 U4804 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3873) );
  INV_X1 U4805 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4703) );
  XNOR2_X1 U4806 ( .A(n3876), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4909)
         );
  NOR2_X1 U4807 ( .A1(n4909), .A2(n6431), .ZN(n3877) );
  NAND2_X1 U4808 ( .A1(n3882), .A2(n3878), .ZN(n3894) );
  NOR2_X1 U4809 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n6291) );
  INV_X1 U4810 ( .A(EBX_REG_31__SCAN_IN), .ZN(n3879) );
  OR2_X1 U4811 ( .A1(n6291), .A2(n3879), .ZN(n3880) );
  NOR2_X1 U4812 ( .A1(n4156), .A2(n3880), .ZN(n3881) );
  NAND2_X1 U4813 ( .A1(n4586), .A2(n3882), .ZN(n3890) );
  AND2_X2 U4814 ( .A1(n3890), .A2(n3094), .ZN(n4155) );
  INV_X1 U4815 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U4816 ( .A1(n4155), .A2(n5759), .ZN(n3884) );
  INV_X4 U4817 ( .A(n3894), .ZN(n4222) );
  MUX2_X1 U4818 ( .A(n3889), .B(n3094), .S(EBX_REG_1__SCAN_IN), .Z(n3883) );
  INV_X1 U4819 ( .A(EBX_REG_0__SCAN_IN), .ZN(n3885) );
  OR2_X1 U4820 ( .A1(n3890), .A2(n3885), .ZN(n3887) );
  NAND2_X1 U4821 ( .A1(n4987), .A2(n3885), .ZN(n3886) );
  NAND2_X1 U4822 ( .A1(n3887), .A2(n3886), .ZN(n4552) );
  XNOR2_X1 U4823 ( .A(n3888), .B(n4552), .ZN(n4223) );
  OR2_X1 U4824 ( .A1(n4144), .A2(EBX_REG_2__SCAN_IN), .ZN(n3893) );
  NAND2_X1 U4825 ( .A1(n3093), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3891)
         );
  OAI211_X1 U4826 ( .C1(n4156), .C2(EBX_REG_2__SCAN_IN), .A(n3967), .B(n3891), 
        .ZN(n3892) );
  AND2_X1 U4827 ( .A1(n3893), .A2(n3892), .ZN(n5514) );
  NAND2_X1 U4828 ( .A1(n5515), .A2(n5514), .ZN(n4255) );
  MUX2_X1 U4829 ( .A(n3959), .B(n3967), .S(EBX_REG_3__SCAN_IN), .Z(n3897) );
  NAND2_X1 U4830 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4156), .ZN(n3895)
         );
  AND2_X1 U4831 ( .A1(n3961), .A2(n3895), .ZN(n3896) );
  INV_X1 U4832 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U4833 ( .A1(n4155), .A2(n5731), .ZN(n3899) );
  MUX2_X1 U4834 ( .A(n4144), .B(n3093), .S(EBX_REG_4__SCAN_IN), .Z(n3898) );
  NAND2_X1 U4835 ( .A1(n3899), .A2(n3898), .ZN(n4318) );
  NOR2_X4 U4836 ( .A1(n4317), .A2(n4318), .ZN(n4410) );
  MUX2_X1 U4837 ( .A(n3959), .B(n3967), .S(EBX_REG_5__SCAN_IN), .Z(n3902) );
  NAND2_X1 U4838 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4156), .ZN(n3900)
         );
  AND2_X1 U4839 ( .A1(n3961), .A2(n3900), .ZN(n3901) );
  INV_X1 U4840 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U4841 ( .A1(n4155), .A2(n5719), .ZN(n3904) );
  MUX2_X1 U4842 ( .A(n4144), .B(n3094), .S(EBX_REG_6__SCAN_IN), .Z(n3903) );
  NAND2_X1 U4843 ( .A1(n3904), .A2(n3903), .ZN(n4407) );
  NOR2_X1 U4844 ( .A1(n4406), .A2(n4407), .ZN(n3905) );
  AND2_X2 U4845 ( .A1(n4410), .A2(n3905), .ZN(n4433) );
  INV_X1 U4846 ( .A(n3959), .ZN(n4152) );
  INV_X1 U4847 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U4848 ( .A1(n4152), .A2(n5459), .ZN(n3908) );
  INV_X1 U4849 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U4850 ( .A1(n3967), .A2(n6517), .ZN(n3906) );
  OAI211_X1 U4851 ( .C1(n4156), .C2(EBX_REG_7__SCAN_IN), .A(n3906), .B(n3093), 
        .ZN(n3907) );
  NAND2_X1 U4852 ( .A1(n3908), .A2(n3907), .ZN(n4432) );
  NAND2_X1 U4853 ( .A1(n4433), .A2(n4432), .ZN(n4431) );
  INV_X1 U4854 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U4855 ( .A1(n4155), .A2(n5697), .ZN(n3910) );
  MUX2_X1 U4856 ( .A(n4144), .B(n3094), .S(EBX_REG_8__SCAN_IN), .Z(n3909) );
  NAND2_X1 U4857 ( .A1(n3910), .A2(n3909), .ZN(n4457) );
  OR2_X2 U4858 ( .A1(n4431), .A2(n4457), .ZN(n4516) );
  MUX2_X1 U4859 ( .A(n3959), .B(n3967), .S(EBX_REG_9__SCAN_IN), .Z(n3913) );
  NAND2_X1 U4860 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n4156), .ZN(n3911)
         );
  AND2_X1 U4861 ( .A1(n3961), .A2(n3911), .ZN(n3912) );
  NAND2_X1 U4862 ( .A1(n3913), .A2(n3912), .ZN(n4546) );
  OR2_X1 U4863 ( .A1(n4144), .A2(EBX_REG_10__SCAN_IN), .ZN(n3916) );
  NAND2_X1 U4864 ( .A1(n3093), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3914) );
  OAI211_X1 U4865 ( .C1(n4156), .C2(EBX_REG_10__SCAN_IN), .A(n3967), .B(n3914), 
        .ZN(n3915) );
  NAND2_X1 U4866 ( .A1(n4546), .A2(n4545), .ZN(n3917) );
  OR2_X2 U4867 ( .A1(n4516), .A2(n3917), .ZN(n4613) );
  MUX2_X1 U4868 ( .A(n3959), .B(n3967), .S(EBX_REG_11__SCAN_IN), .Z(n3920) );
  NAND2_X1 U4869 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n4156), .ZN(n3918) );
  AND2_X1 U4870 ( .A1(n3961), .A2(n3918), .ZN(n3919) );
  OR2_X1 U4871 ( .A1(n4144), .A2(EBX_REG_12__SCAN_IN), .ZN(n3923) );
  NAND2_X1 U4872 ( .A1(n3094), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3921) );
  OAI211_X1 U4873 ( .C1(n4156), .C2(EBX_REG_12__SCAN_IN), .A(n3967), .B(n3921), 
        .ZN(n3922) );
  MUX2_X1 U4874 ( .A(n3959), .B(n3967), .S(EBX_REG_13__SCAN_IN), .Z(n3926) );
  NAND2_X1 U4875 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4156), .ZN(n3924) );
  AND2_X1 U4876 ( .A1(n3961), .A2(n3924), .ZN(n3925) );
  NAND2_X1 U4877 ( .A1(n3926), .A2(n3925), .ZN(n4825) );
  OR2_X1 U4878 ( .A1(n4144), .A2(EBX_REG_14__SCAN_IN), .ZN(n3929) );
  NAND2_X1 U4879 ( .A1(n3093), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3927) );
  OAI211_X1 U4880 ( .C1(n4156), .C2(EBX_REG_14__SCAN_IN), .A(n3967), .B(n3927), 
        .ZN(n3928) );
  NAND2_X1 U4881 ( .A1(n4825), .A2(n4824), .ZN(n3930) );
  MUX2_X1 U4882 ( .A(n3959), .B(n3967), .S(EBX_REG_15__SCAN_IN), .Z(n3933) );
  NAND2_X1 U4883 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n4156), .ZN(n3931) );
  AND2_X1 U4884 ( .A1(n3961), .A2(n3931), .ZN(n3932) );
  INV_X1 U4885 ( .A(EBX_REG_16__SCAN_IN), .ZN(n3934) );
  INV_X1 U4886 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6682) );
  OAI22_X1 U4887 ( .A1(n4155), .A2(n3934), .B1(n4222), .B2(n6682), .ZN(n3935)
         );
  XNOR2_X1 U4888 ( .A(n3935), .B(n3094), .ZN(n4951) );
  AND2_X2 U4889 ( .A1(n5332), .A2(n4951), .ZN(n5314) );
  MUX2_X1 U4890 ( .A(n3959), .B(n3967), .S(EBX_REG_17__SCAN_IN), .Z(n3938) );
  NAND2_X1 U4891 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n4156), .ZN(n3936) );
  AND2_X1 U4892 ( .A1(n3961), .A2(n3936), .ZN(n3937) );
  NAND2_X1 U4893 ( .A1(n3938), .A2(n3937), .ZN(n5313) );
  INV_X1 U4894 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U4895 ( .A1(n4155), .A2(n6701), .ZN(n3940) );
  MUX2_X1 U4896 ( .A(n4144), .B(n3093), .S(EBX_REG_19__SCAN_IN), .Z(n3939) );
  NAND2_X1 U4897 ( .A1(n3940), .A2(n3939), .ZN(n5150) );
  INV_X1 U4898 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3941) );
  NAND2_X1 U4899 ( .A1(n4155), .A2(n3941), .ZN(n3943) );
  INV_X1 U4900 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U4901 ( .A1(n4222), .A2(n4994), .ZN(n3942) );
  NAND2_X1 U4902 ( .A1(n3943), .A2(n3942), .ZN(n4937) );
  INV_X1 U4903 ( .A(n4937), .ZN(n4988) );
  INV_X1 U4904 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U4905 ( .A1(n4155), .A2(n5299), .ZN(n3946) );
  INV_X1 U4906 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3944) );
  NAND2_X1 U4907 ( .A1(n4222), .A2(n3944), .ZN(n3945) );
  NAND2_X1 U4908 ( .A1(n3946), .A2(n3945), .ZN(n4989) );
  NAND2_X1 U4909 ( .A1(n4937), .A2(n3944), .ZN(n3947) );
  OAI21_X1 U4910 ( .B1(n4989), .B2(n4987), .A(n3947), .ZN(n3948) );
  OAI21_X1 U4911 ( .B1(n4987), .B2(n4988), .A(n3948), .ZN(n3949) );
  INV_X1 U4912 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U4913 ( .A1(n4155), .A2(n5288), .ZN(n3951) );
  MUX2_X1 U4914 ( .A(n4144), .B(n3093), .S(EBX_REG_21__SCAN_IN), .Z(n3950) );
  AND2_X1 U4915 ( .A1(n3951), .A2(n3950), .ZN(n5130) );
  NAND2_X1 U4916 ( .A1(n5131), .A2(n5130), .ZN(n4983) );
  MUX2_X1 U4917 ( .A(n3959), .B(n3967), .S(EBX_REG_22__SCAN_IN), .Z(n3954) );
  INV_X1 U4918 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5281) );
  OAI21_X1 U4919 ( .B1(n4222), .B2(n5281), .A(n3961), .ZN(n3952) );
  INV_X1 U4920 ( .A(n3952), .ZN(n3953) );
  NOR2_X2 U4921 ( .A1(n4983), .A2(n4982), .ZN(n4981) );
  OR2_X1 U4922 ( .A1(n4144), .A2(EBX_REG_23__SCAN_IN), .ZN(n3957) );
  NAND2_X1 U4923 ( .A1(n3094), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3955) );
  OAI211_X1 U4924 ( .C1(n4156), .C2(EBX_REG_23__SCAN_IN), .A(n3967), .B(n3955), 
        .ZN(n3956) );
  NAND2_X1 U4925 ( .A1(n3957), .A2(n3956), .ZN(n5113) );
  NAND2_X1 U4926 ( .A1(n4981), .A2(n3958), .ZN(n5116) );
  MUX2_X1 U4927 ( .A(n3959), .B(n3967), .S(EBX_REG_24__SCAN_IN), .Z(n3963) );
  NAND2_X1 U4928 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n4156), .ZN(n3960) );
  AND2_X1 U4929 ( .A1(n3961), .A2(n3960), .ZN(n3962) );
  NOR2_X2 U4930 ( .A1(n5116), .A2(n4207), .ZN(n4208) );
  OR2_X1 U4931 ( .A1(n4144), .A2(EBX_REG_25__SCAN_IN), .ZN(n3966) );
  NAND2_X1 U4932 ( .A1(n3093), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3964) );
  OAI211_X1 U4933 ( .C1(n4156), .C2(EBX_REG_25__SCAN_IN), .A(n3967), .B(n3964), 
        .ZN(n3965) );
  AND2_X1 U4934 ( .A1(n3966), .A2(n3965), .ZN(n4925) );
  NAND2_X1 U4935 ( .A1(n4208), .A2(n4925), .ZN(n4926) );
  INV_X1 U4936 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4855) );
  NAND2_X1 U4937 ( .A1(n4152), .A2(n4855), .ZN(n3970) );
  INV_X1 U4938 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U4939 ( .A1(n3967), .A2(n5253), .ZN(n3968) );
  OAI211_X1 U4940 ( .C1(n4156), .C2(EBX_REG_26__SCAN_IN), .A(n3968), .B(n3094), 
        .ZN(n3969) );
  NAND2_X1 U4941 ( .A1(n4926), .A2(n3971), .ZN(n3972) );
  NAND2_X1 U4942 ( .A1(n3099), .A2(n3972), .ZN(n5258) );
  OAI22_X1 U4943 ( .A1(n4854), .A2(n5452), .B1(n5449), .B2(n5258), .ZN(n3989)
         );
  INV_X1 U4944 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6504) );
  INV_X1 U4945 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6583) );
  INV_X1 U4946 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5162) );
  INV_X1 U4947 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6622) );
  INV_X1 U4948 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U4949 ( .A1(n3973), .A2(n6326), .ZN(n6321) );
  NAND2_X1 U4950 ( .A1(n4279), .A2(n6321), .ZN(n4099) );
  AND3_X1 U4951 ( .A1(n4099), .A2(n6291), .A3(n3882), .ZN(n3974) );
  INV_X1 U4952 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6348) );
  INV_X1 U4953 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6345) );
  INV_X1 U4954 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6407) );
  INV_X1 U4955 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6335) );
  INV_X1 U4956 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6333) );
  NOR3_X1 U4957 ( .A1(n6407), .A2(n6335), .A3(n6333), .ZN(n5488) );
  NAND3_X1 U4958 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .A3(
        n5488), .ZN(n5423) );
  NAND3_X1 U4959 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U4960 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5421) );
  NOR4_X1 U4961 ( .A1(n6345), .A2(n5423), .A3(n5422), .A4(n5421), .ZN(n5409)
         );
  NAND2_X1 U4962 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5409), .ZN(n5405) );
  NOR2_X1 U4963 ( .A1(n6348), .A2(n5405), .ZN(n4831) );
  NAND2_X1 U4964 ( .A1(REIP_REG_14__SCAN_IN), .A2(n4831), .ZN(n3975) );
  NAND3_X1 U4965 ( .A1(n4954), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U4966 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5161), .ZN(n5154) );
  NAND2_X1 U4967 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5145), .ZN(n5124) );
  NAND2_X1 U4968 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5125) );
  NAND2_X1 U4969 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5118), .ZN(n4899) );
  OR2_X1 U4970 ( .A1(n6583), .A2(n4899), .ZN(n4924) );
  INV_X1 U4971 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6639) );
  OAI21_X1 U4972 ( .B1(n6504), .B2(n4924), .A(n6639), .ZN(n3980) );
  NAND3_X1 U4973 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4898) );
  NAND2_X1 U4974 ( .A1(n5487), .A2(n5486), .ZN(n4558) );
  INV_X1 U4975 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6361) );
  INV_X1 U4976 ( .A(n4558), .ZN(n5424) );
  INV_X1 U4977 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6357) );
  INV_X1 U4978 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6487) );
  NOR3_X1 U4979 ( .A1(n6357), .A2(n5162), .A3(n6487), .ZN(n3977) );
  INV_X1 U4980 ( .A(n5486), .ZN(n5507) );
  NOR2_X1 U4981 ( .A1(n5507), .A2(n3975), .ZN(n4832) );
  NAND4_X1 U4982 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(n4832), .ZN(n3976) );
  NAND2_X1 U4983 ( .A1(n4558), .A2(n3976), .ZN(n5387) );
  OAI21_X1 U4984 ( .B1(n5424), .B2(n3977), .A(n5387), .ZN(n5146) );
  AOI221_X1 U4985 ( .B1(n6361), .B2(n4558), .C1(n5125), .C2(n4558), .A(n5146), 
        .ZN(n3978) );
  INV_X1 U4986 ( .A(n3978), .ZN(n5117) );
  AOI21_X1 U4987 ( .B1(n4898), .B2(n4558), .A(n5117), .ZN(n3979) );
  INV_X1 U4988 ( .A(n3979), .ZN(n5105) );
  AND2_X1 U4989 ( .A1(n4909), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4990 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n5519), .B1(n4863), 
        .B2(n5520), .ZN(n3982) );
  INV_X1 U4991 ( .A(n6321), .ZN(n6292) );
  AOI21_X1 U4992 ( .B1(n6292), .B2(n6291), .A(n6423), .ZN(n4894) );
  NOR3_X1 U4993 ( .A1(n4334), .A2(EBX_REG_31__SCAN_IN), .A3(n6291), .ZN(n3983)
         );
  OR2_X1 U4994 ( .A1(n3989), .A2(n3988), .ZN(U2801) );
  NAND2_X1 U4995 ( .A1(n4334), .A2(n3990), .ZN(n4118) );
  OAI21_X1 U4996 ( .B1(n6423), .B2(n3994), .A(n4118), .ZN(n3991) );
  INV_X1 U4997 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6679) );
  NOR2_X1 U4998 ( .A1(n5675), .A2(n6679), .ZN(n5674) );
  NAND2_X1 U4999 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5742) );
  OR2_X1 U5000 ( .A1(n5675), .A2(n5742), .ZN(n4001) );
  OAI21_X1 U5001 ( .B1(n5674), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4001), 
        .ZN(n3992) );
  INV_X1 U5002 ( .A(n3992), .ZN(n4386) );
  NAND2_X1 U5003 ( .A1(n3096), .A2(n4046), .ZN(n4000) );
  NAND2_X1 U5004 ( .A1(n3995), .A2(n3994), .ZN(n4003) );
  OAI211_X1 U5005 ( .C1(n3995), .C2(n3994), .A(n5605), .B(n4003), .ZN(n3998)
         );
  AND3_X1 U5006 ( .A1(n3998), .A2(n3997), .A3(n3996), .ZN(n3999) );
  NAND2_X1 U5007 ( .A1(n4000), .A2(n3999), .ZN(n4385) );
  NAND2_X1 U5008 ( .A1(n4386), .A2(n4385), .ZN(n4384) );
  NAND2_X1 U5009 ( .A1(n4384), .A2(n4001), .ZN(n5667) );
  NAND2_X1 U5010 ( .A1(n4263), .A2(n4046), .ZN(n4008) );
  NAND2_X1 U5011 ( .A1(n4003), .A2(n4004), .ZN(n4017) );
  OAI21_X1 U5012 ( .B1(n4004), .B2(n4003), .A(n4017), .ZN(n4006) );
  INV_X1 U5013 ( .A(n4118), .ZN(n4005) );
  AOI21_X1 U5014 ( .B1(n4006), .B2(n5605), .A(n4005), .ZN(n4007) );
  NAND2_X1 U5015 ( .A1(n4008), .A2(n4007), .ZN(n4009) );
  OAI21_X1 U5016 ( .B1(n5667), .B2(n5663), .A(n5664), .ZN(n4321) );
  NAND2_X1 U5017 ( .A1(n4380), .A2(n4046), .ZN(n4013) );
  INV_X1 U5018 ( .A(n4018), .ZN(n4010) );
  XNOR2_X1 U5019 ( .A(n4017), .B(n4010), .ZN(n4011) );
  NAND2_X1 U5020 ( .A1(n4011), .A2(n5605), .ZN(n4012) );
  NAND2_X1 U5021 ( .A1(n4013), .A2(n4012), .ZN(n4014) );
  XNOR2_X1 U5022 ( .A(n4014), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4320)
         );
  NAND2_X1 U5023 ( .A1(n4014), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4015)
         );
  NAND2_X1 U5024 ( .A1(n4016), .A2(n4046), .ZN(n4021) );
  NAND2_X1 U5025 ( .A1(n4018), .A2(n4017), .ZN(n4025) );
  XOR2_X1 U5026 ( .A(n4026), .B(n4025), .Z(n4019) );
  NAND2_X1 U5027 ( .A1(n4019), .A2(n5605), .ZN(n4020) );
  NAND2_X1 U5028 ( .A1(n4021), .A2(n4020), .ZN(n4022) );
  XNOR2_X1 U5029 ( .A(n4022), .B(n5731), .ZN(n4327) );
  NAND2_X1 U5030 ( .A1(n4326), .A2(n4327), .ZN(n4024) );
  NAND2_X1 U5031 ( .A1(n4022), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4023)
         );
  NAND2_X1 U5032 ( .A1(n4024), .A2(n4023), .ZN(n4397) );
  NOR2_X1 U5033 ( .A1(n4026), .A2(n4025), .ZN(n4036) );
  XNOR2_X1 U5034 ( .A(n4036), .B(n4035), .ZN(n4027) );
  OAI22_X1 U5035 ( .A1(n4029), .A2(n4028), .B1(n4027), .B2(n6423), .ZN(n4030)
         );
  INV_X1 U5036 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4130) );
  XNOR2_X1 U5037 ( .A(n4030), .B(n4130), .ZN(n4398) );
  NAND2_X1 U5038 ( .A1(n4397), .A2(n4398), .ZN(n4032) );
  NAND2_X1 U5039 ( .A1(n4030), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4031)
         );
  NAND2_X1 U5040 ( .A1(n4032), .A2(n4031), .ZN(n4507) );
  AND2_X1 U5041 ( .A1(n4046), .A2(n4054), .ZN(n4033) );
  NAND2_X1 U5042 ( .A1(n4034), .A2(n4033), .ZN(n4039) );
  NAND2_X1 U5043 ( .A1(n4036), .A2(n4035), .ZN(n4043) );
  XOR2_X1 U5044 ( .A(n4044), .B(n4043), .Z(n4037) );
  NAND2_X1 U5045 ( .A1(n4037), .A2(n5605), .ZN(n4038) );
  NAND2_X1 U5046 ( .A1(n4039), .A2(n4038), .ZN(n4040) );
  XNOR2_X1 U5047 ( .A(n4040), .B(n5719), .ZN(n4508) );
  NAND2_X1 U5048 ( .A1(n4507), .A2(n4508), .ZN(n4042) );
  NAND2_X1 U5049 ( .A1(n4040), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4041)
         );
  NAND2_X1 U5050 ( .A1(n4042), .A2(n4041), .ZN(n4501) );
  NOR2_X1 U5051 ( .A1(n4044), .A2(n4043), .ZN(n4053) );
  XOR2_X1 U5052 ( .A(n4045), .B(n4053), .Z(n4049) );
  NAND2_X1 U5053 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  OAI21_X1 U5054 ( .B1(n4049), .B2(n6423), .A(n4048), .ZN(n4050) );
  XNOR2_X1 U5055 ( .A(n4050), .B(n6517), .ZN(n4502) );
  NAND2_X1 U5056 ( .A1(n4501), .A2(n4502), .ZN(n4052) );
  NAND2_X1 U5057 ( .A1(n4050), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4051)
         );
  NAND2_X1 U5058 ( .A1(n4052), .A2(n4051), .ZN(n4562) );
  NAND2_X1 U5059 ( .A1(n4053), .A2(n4055), .ZN(n4058) );
  INV_X1 U5060 ( .A(n4117), .ZN(n4057) );
  OAI21_X1 U5061 ( .B1(n4058), .B2(n6423), .A(n5054), .ZN(n4059) );
  XNOR2_X1 U5062 ( .A(n4059), .B(n5697), .ZN(n4563) );
  NAND2_X1 U5063 ( .A1(n4562), .A2(n4563), .ZN(n4061) );
  NAND2_X1 U5064 ( .A1(n4059), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4060)
         );
  INV_X1 U5065 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4542) );
  NOR2_X1 U5066 ( .A1(n5054), .A2(n4542), .ZN(n4063) );
  NAND2_X1 U5067 ( .A1(n5224), .A2(n4542), .ZN(n4062) );
  INV_X1 U5068 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4541) );
  AND2_X1 U5069 ( .A1(n5224), .A2(n4541), .ZN(n4526) );
  NAND2_X1 U5070 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4527) );
  INV_X1 U5071 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U5072 ( .A1(n5224), .A2(n6579), .ZN(n4628) );
  NAND2_X1 U5073 ( .A1(n4627), .A2(n4628), .ZN(n4064) );
  NAND2_X1 U5074 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4629) );
  NAND2_X1 U5075 ( .A1(n4064), .A2(n4629), .ZN(n4637) );
  INV_X1 U5076 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4065) );
  NOR2_X1 U5077 ( .A1(n5054), .A2(n4065), .ZN(n4640) );
  OR2_X2 U5078 ( .A1(n4637), .A2(n4640), .ZN(n4169) );
  NAND2_X1 U5079 ( .A1(n5224), .A2(n4065), .ZN(n4638) );
  INV_X1 U5080 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4066) );
  NAND2_X1 U5081 ( .A1(n5224), .A2(n4066), .ZN(n4807) );
  NAND2_X1 U5082 ( .A1(n5224), .A2(n6682), .ZN(n4067) );
  INV_X1 U5083 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5340) );
  INV_X1 U5084 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U5085 ( .A1(n5224), .A2(n5354), .ZN(n5045) );
  AND2_X1 U5086 ( .A1(n4067), .A2(n4809), .ZN(n4068) );
  NAND2_X1 U5087 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4129) );
  NAND2_X1 U5088 ( .A1(n5224), .A2(n4129), .ZN(n4069) );
  AND2_X1 U5089 ( .A1(n4638), .A2(n4172), .ZN(n4074) );
  INV_X1 U5090 ( .A(n4172), .ZN(n4070) );
  XNOR2_X1 U5091 ( .A(n5054), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4661)
         );
  OR2_X1 U5092 ( .A1(n4070), .A2(n4661), .ZN(n4072) );
  INV_X1 U5093 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U5094 ( .A1(n6682), .A2(n5321), .ZN(n4812) );
  OAI21_X1 U5095 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n4812), .A(n4178), 
        .ZN(n4071) );
  NAND2_X1 U5096 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U5097 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U5098 ( .A1(n4072), .A2(n4170), .ZN(n4073) );
  AOI21_X2 U5099 ( .B1(n4169), .B2(n4074), .A(n4073), .ZN(n4077) );
  INV_X1 U5100 ( .A(n4077), .ZN(n4081) );
  NOR2_X1 U5101 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5292) );
  NOR2_X1 U5102 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5275) );
  INV_X1 U5103 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5064) );
  INV_X1 U5104 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5065) );
  NAND4_X1 U5105 ( .A1(n5292), .A2(n5275), .A3(n5064), .A4(n5065), .ZN(n4080)
         );
  AND2_X1 U5106 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4137) );
  INV_X1 U5107 ( .A(n4137), .ZN(n4164) );
  AND2_X1 U5108 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5293) );
  INV_X1 U5109 ( .A(n5293), .ZN(n4163) );
  NAND2_X1 U5110 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5273) );
  NAND3_X1 U5111 ( .A1(n4137), .A2(n5293), .A3(n4075), .ZN(n4076) );
  XNOR2_X1 U5112 ( .A(n5054), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5204)
         );
  NAND2_X2 U5113 ( .A1(n5205), .A2(n5204), .ZN(n5203) );
  NAND2_X2 U5114 ( .A1(n5203), .A2(n4083), .ZN(n4867) );
  NAND2_X1 U5115 ( .A1(n5224), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4860) );
  NOR2_X2 U5116 ( .A1(n4867), .A2(n4860), .ZN(n5197) );
  NAND3_X1 U5117 ( .A1(n5197), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4688) );
  NAND2_X1 U5118 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4165) );
  NAND2_X1 U5119 ( .A1(n4178), .A2(n5253), .ZN(n5010) );
  INV_X1 U5120 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U5121 ( .A1(n5014), .A2(n5011), .ZN(n5239) );
  NOR3_X1 U5122 ( .A1(n5010), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5239), 
        .ZN(n4689) );
  INV_X1 U5123 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6731) );
  NAND2_X1 U5124 ( .A1(n4689), .A2(n6731), .ZN(n4084) );
  OAI22_X1 U5125 ( .A1(n4688), .A2(n4165), .B1(n5203), .B2(n4084), .ZN(n4085)
         );
  XNOR2_X1 U5126 ( .A(n4085), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4912)
         );
  INV_X1 U5127 ( .A(n6282), .ZN(n4086) );
  NOR2_X1 U5128 ( .A1(n4088), .A2(n4279), .ZN(n4124) );
  NAND2_X1 U5129 ( .A1(n4086), .A2(n4124), .ZN(n4231) );
  NOR2_X1 U5130 ( .A1(n4087), .A2(n4114), .ZN(n4090) );
  NAND2_X1 U5131 ( .A1(n4088), .A2(n4334), .ZN(n4089) );
  NAND2_X1 U5132 ( .A1(n4091), .A2(n3882), .ZN(n4092) );
  MUX2_X1 U5133 ( .A(n6423), .B(n4092), .S(n4297), .Z(n4109) );
  NAND2_X1 U5134 ( .A1(n4105), .A2(n4109), .ZN(n4094) );
  NAND2_X1 U5135 ( .A1(n4094), .A2(n4093), .ZN(n4233) );
  NAND2_X1 U5136 ( .A1(n3878), .A2(n6321), .ZN(n4096) );
  INV_X1 U5137 ( .A(n4095), .ZN(n6277) );
  NOR2_X1 U5138 ( .A1(n6277), .A2(READY_N), .ZN(n4225) );
  NAND3_X1 U5139 ( .A1(n4096), .A2(n4225), .A3(n4116), .ZN(n4097) );
  NAND3_X1 U5140 ( .A1(n4231), .A2(n4233), .A3(n4097), .ZN(n4098) );
  NAND2_X1 U5141 ( .A1(n4098), .A2(n6293), .ZN(n4102) );
  INV_X1 U5142 ( .A(READY_N), .ZN(n6420) );
  NAND2_X1 U5143 ( .A1(n4099), .A2(n6420), .ZN(n4229) );
  OAI211_X1 U5144 ( .C1(n4242), .C2(n4229), .A(n3882), .B(n4299), .ZN(n4100)
         );
  NAND3_X1 U5145 ( .A1(n5604), .A2(n4446), .A3(n4100), .ZN(n4101) );
  OAI211_X1 U5146 ( .C1(n4390), .C2(n4160), .A(n4370), .B(n4294), .ZN(n4103)
         );
  INV_X1 U5147 ( .A(n4103), .ZN(n4106) );
  NAND2_X1 U5148 ( .A1(n4105), .A2(n4104), .ZN(n6284) );
  NAND2_X1 U5149 ( .A1(n4105), .A2(n3095), .ZN(n6275) );
  NAND3_X1 U5150 ( .A1(n4106), .A2(n6284), .A3(n6275), .ZN(n4107) );
  INV_X1 U5151 ( .A(n4165), .ZN(n4140) );
  NAND2_X1 U5152 ( .A1(n4087), .A2(n4987), .ZN(n4108) );
  AND2_X1 U5153 ( .A1(n4109), .A2(n4108), .ZN(n4110) );
  NAND2_X1 U5154 ( .A1(n4111), .A2(n4110), .ZN(n4247) );
  INV_X1 U5155 ( .A(n4112), .ZN(n4113) );
  NAND2_X1 U5156 ( .A1(n4113), .A2(n6261), .ZN(n4353) );
  NAND2_X1 U5157 ( .A1(n4334), .A2(n3878), .ZN(n5369) );
  OR2_X1 U5158 ( .A1(n5369), .A2(n4116), .ZN(n4232) );
  NAND2_X1 U5159 ( .A1(n4155), .A2(n4232), .ZN(n4115) );
  NAND2_X1 U5160 ( .A1(n4115), .A2(n4114), .ZN(n4244) );
  OAI21_X1 U5161 ( .B1(n4299), .B2(n3882), .A(n4116), .ZN(n4240) );
  OAI21_X1 U5162 ( .B1(n4118), .B2(n4117), .A(n4240), .ZN(n4119) );
  INV_X1 U5163 ( .A(n4119), .ZN(n4122) );
  OR2_X1 U5164 ( .A1(n4241), .A2(n4120), .ZN(n4121) );
  NAND4_X1 U5165 ( .A1(n4353), .A2(n4244), .A3(n4122), .A4(n4121), .ZN(n4123)
         );
  INV_X1 U5166 ( .A(n4124), .ZN(n4125) );
  INV_X1 U5167 ( .A(n5369), .ZN(n4464) );
  NAND2_X1 U5168 ( .A1(n4126), .A2(n4464), .ZN(n5075) );
  INV_X1 U5169 ( .A(n5075), .ZN(n6264) );
  NAND2_X1 U5170 ( .A1(n4162), .A2(n4127), .ZN(n4132) );
  NAND2_X1 U5171 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5241) );
  AOI21_X1 U5172 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n5723) );
  NAND2_X1 U5173 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5722) );
  NOR2_X1 U5174 ( .A1(n5723), .A2(n5722), .ZN(n4468) );
  NAND2_X1 U5175 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4468), .ZN(n4537)
         );
  NOR2_X1 U5176 ( .A1(n5719), .A2(n4537), .ZN(n4533) );
  NAND2_X1 U5177 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U5178 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4543) );
  NOR2_X1 U5179 ( .A1(n5702), .A2(n4543), .ZN(n4131) );
  NAND2_X1 U5180 ( .A1(n4533), .A2(n4131), .ZN(n4648) );
  INV_X1 U5181 ( .A(n4648), .ZN(n4128) );
  NAND2_X1 U5182 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5324) );
  NOR2_X1 U5183 ( .A1(n6579), .A2(n4065), .ZN(n4666) );
  NAND2_X1 U5184 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4666), .ZN(n4664) );
  OR2_X1 U5185 ( .A1(n5354), .A2(n4664), .ZN(n5323) );
  NOR2_X1 U5186 ( .A1(n5324), .A2(n5323), .ZN(n4133) );
  NAND2_X1 U5187 ( .A1(n4128), .A2(n4133), .ZN(n5291) );
  OR2_X1 U5188 ( .A1(n4163), .A2(n4129), .ZN(n4177) );
  INV_X1 U5189 ( .A(n4647), .ZN(n4532) );
  NAND4_X1 U5190 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4474) );
  NOR3_X1 U5191 ( .A1(n4130), .A2(n5719), .A3(n4474), .ZN(n4531) );
  NAND2_X1 U5192 ( .A1(n4131), .A2(n4531), .ZN(n4646) );
  INV_X1 U5193 ( .A(n4646), .ZN(n4134) );
  INV_X1 U5194 ( .A(n4132), .ZN(n5345) );
  NOR2_X1 U5195 ( .A1(n5721), .A2(n5345), .ZN(n5765) );
  OAI22_X1 U5196 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5765), .B1(n5348), 
        .B2(n4162), .ZN(n5767) );
  NAND2_X1 U5197 ( .A1(n5741), .A2(n5767), .ZN(n4649) );
  OAI221_X1 U5198 ( .B1(n4532), .B2(n4134), .C1(n4532), .C2(n4133), .A(n4649), 
        .ZN(n5290) );
  AOI221_X1 U5199 ( .B1(n5291), .B2(n5757), .C1(n4177), .C2(n5757), .A(n5290), 
        .ZN(n5289) );
  OR2_X1 U5200 ( .A1(n4536), .A2(n4075), .ZN(n4135) );
  NAND2_X1 U5201 ( .A1(n5289), .A2(n4135), .ZN(n5266) );
  NAND2_X1 U5202 ( .A1(n6679), .A2(n4136), .ZN(n5758) );
  AOI21_X1 U5203 ( .B1(n5752), .B2(n5741), .A(n4137), .ZN(n4138) );
  NAND3_X1 U5204 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n4139), .ZN(n5237) );
  NAND2_X1 U5205 ( .A1(n4139), .A2(n4536), .ZN(n5238) );
  OAI21_X1 U5206 ( .B1(n5241), .B2(n5237), .A(n5238), .ZN(n4700) );
  OAI21_X1 U5207 ( .B1(n4140), .B2(n4536), .A(n4700), .ZN(n4141) );
  NAND2_X1 U5208 ( .A1(n4141), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4168) );
  INV_X1 U5209 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4914) );
  OR2_X1 U5210 ( .A1(n4155), .A2(n4914), .ZN(n4143) );
  NAND2_X1 U5211 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4142) );
  AND2_X1 U5212 ( .A1(n4143), .A2(n4142), .ZN(n4693) );
  NAND2_X1 U5213 ( .A1(n4155), .A2(n5011), .ZN(n4146) );
  MUX2_X1 U5214 ( .A(n4144), .B(n3094), .S(EBX_REG_27__SCAN_IN), .Z(n4145) );
  NAND2_X1 U5215 ( .A1(n4146), .A2(n4145), .ZN(n4975) );
  NOR2_X4 U5216 ( .A1(n3099), .A2(n4975), .ZN(n4977) );
  INV_X1 U5217 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U5218 ( .A1(n4152), .A2(n6528), .ZN(n4149) );
  NAND2_X1 U5219 ( .A1(n3967), .A2(n5014), .ZN(n4147) );
  OAI211_X1 U5220 ( .C1(n4156), .C2(EBX_REG_28__SCAN_IN), .A(n4147), .B(n3093), 
        .ZN(n4148) );
  NAND2_X1 U5221 ( .A1(n4149), .A2(n4148), .ZN(n4967) );
  INV_X1 U5222 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6515) );
  NOR2_X1 U5223 ( .A1(n4156), .A2(EBX_REG_29__SCAN_IN), .ZN(n4150) );
  AOI21_X1 U5224 ( .B1(n4155), .B2(n6515), .A(n4150), .ZN(n4874) );
  INV_X1 U5225 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4961) );
  AND2_X1 U5226 ( .A1(n4152), .A2(n4961), .ZN(n4875) );
  NAND2_X1 U5227 ( .A1(n4151), .A2(n4875), .ZN(n4153) );
  NOR2_X1 U5228 ( .A1(n4694), .A2(n4987), .ZN(n4691) );
  AOI21_X1 U5229 ( .B1(n4693), .B2(n4880), .A(n4691), .ZN(n4158) );
  INV_X1 U5230 ( .A(n4155), .ZN(n4554) );
  OAI22_X1 U5231 ( .A1(n4554), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4156), .ZN(n4157) );
  XNOR2_X1 U5232 ( .A(n4158), .B(n4157), .ZN(n5531) );
  OAI21_X1 U5233 ( .B1(n4160), .B2(n4159), .A(n6296), .ZN(n4161) );
  INV_X1 U5234 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6684) );
  NOR2_X1 U5235 ( .A1(n5740), .A2(n6684), .ZN(n4907) );
  NAND2_X1 U5236 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5350), .ZN(n5336) );
  NAND3_X1 U5237 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5318), .ZN(n5302) );
  NAND2_X1 U5238 ( .A1(n5285), .A2(n4075), .ZN(n5272) );
  NAND3_X1 U5239 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n5263), .ZN(n5252) );
  NOR3_X1 U5240 ( .A1(n4165), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4883), 
        .ZN(n4166) );
  AOI211_X1 U5241 ( .C1(n5531), .C2(n5754), .A(n4907), .B(n4166), .ZN(n4167)
         );
  OAI211_X1 U5242 ( .C1(n4912), .C2(n5733), .A(n4168), .B(n4167), .ZN(U2987)
         );
  NAND2_X2 U5243 ( .A1(n4662), .A2(n4661), .ZN(n4808) );
  XNOR2_X1 U5244 ( .A(n5054), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5219)
         );
  NAND2_X1 U5245 ( .A1(n5220), .A2(n5219), .ZN(n5032) );
  NAND2_X1 U5246 ( .A1(n5224), .A2(n6701), .ZN(n5031) );
  AND2_X1 U5247 ( .A1(n5031), .A2(n3103), .ZN(n4173) );
  NAND2_X1 U5248 ( .A1(n5032), .A2(n4173), .ZN(n4175) );
  OR2_X1 U5249 ( .A1(n5224), .A2(n5299), .ZN(n4174) );
  NAND2_X1 U5250 ( .A1(n4175), .A2(n4174), .ZN(n5212) );
  XNOR2_X1 U5251 ( .A(n5054), .B(n5288), .ZN(n5213) );
  NOR2_X2 U5252 ( .A1(n5212), .A2(n5213), .ZN(n5211) );
  NOR2_X1 U5253 ( .A1(n5054), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4839)
         );
  NAND2_X1 U5254 ( .A1(n5211), .A2(n4839), .ZN(n5023) );
  NAND2_X1 U5255 ( .A1(n4808), .A2(n4176), .ZN(n4814) );
  OR4_X1 U5256 ( .A1(n4178), .A2(n4814), .A3(n5273), .A4(n4177), .ZN(n4179) );
  NAND2_X1 U5257 ( .A1(n5023), .A2(n4179), .ZN(n4180) );
  INV_X1 U5258 ( .A(n6284), .ZN(n4181) );
  INV_X1 U5259 ( .A(n4182), .ZN(n4843) );
  INV_X1 U5260 ( .A(n4184), .ZN(n4183) );
  NAND2_X1 U5261 ( .A1(n4182), .A2(n4183), .ZN(n4198) );
  NAND2_X1 U5262 ( .A1(n4843), .A2(n4184), .ZN(n4185) );
  NAND2_X1 U5263 ( .A1(n4186), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6314) );
  OR2_X2 U5264 ( .A1(n6314), .A2(n6203), .ZN(n5682) );
  INV_X1 U5265 ( .A(n5682), .ZN(n5669) );
  OR2_X1 U5266 ( .A1(n4187), .A2(n6432), .ZN(n6419) );
  NAND2_X1 U5267 ( .A1(n6419), .A2(n6303), .ZN(n4188) );
  AOI22_X1 U5268 ( .A1(n5348), .A2(REIP_REG_23__SCAN_IN), .B1(n5662), .B2(
        PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4194) );
  NAND2_X1 U5269 ( .A1(n6303), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4190) );
  NAND2_X1 U5270 ( .A1(n6164), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4189) );
  AND2_X1 U5271 ( .A1(n4190), .A2(n4189), .ZN(n5677) );
  INV_X1 U5272 ( .A(n5677), .ZN(n4191) );
  INV_X1 U5273 ( .A(n4921), .ZN(n4200) );
  OAI21_X2 U5274 ( .B1(n4202), .B2(n4201), .A(n4200), .ZN(n5025) );
  INV_X1 U5275 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4203) );
  OAI22_X1 U5276 ( .A1(n4203), .A2(n5499), .B1(n5512), .B2(n5027), .ZN(n4204)
         );
  AOI21_X1 U5277 ( .B1(n5518), .B2(EBX_REG_24__SCAN_IN), .A(n4204), .ZN(n4206)
         );
  NAND2_X1 U5278 ( .A1(n5117), .A2(REIP_REG_24__SCAN_IN), .ZN(n4205) );
  OAI211_X1 U5279 ( .C1(n5025), .C2(n5452), .A(n4206), .B(n4205), .ZN(n4212)
         );
  AND2_X1 U5280 ( .A1(n5116), .A2(n4207), .ZN(n4209) );
  OR2_X1 U5281 ( .A1(n4209), .A2(n4208), .ZN(n5067) );
  NOR2_X1 U5282 ( .A1(REIP_REG_24__SCAN_IN), .A2(n4899), .ZN(n4928) );
  OR2_X1 U5283 ( .A1(n4212), .A2(n4211), .ZN(U2803) );
  INV_X1 U5284 ( .A(n6278), .ZN(n4216) );
  INV_X1 U5285 ( .A(n4301), .ZN(n4916) );
  NAND3_X1 U5286 ( .A1(n4213), .A2(n4390), .A3(n4916), .ZN(n4215) );
  OR2_X1 U5287 ( .A1(n4215), .A2(n4214), .ZN(n4291) );
  OAI22_X1 U5288 ( .A1(n6282), .A2(n4216), .B1(n4156), .B2(n4291), .ZN(n4217)
         );
  NOR2_X1 U5289 ( .A1(n4219), .A2(n4218), .ZN(n4220) );
  OR2_X1 U5290 ( .A1(n4221), .A2(n4220), .ZN(n4467) );
  XNOR2_X1 U5291 ( .A(n4223), .B(n4222), .ZN(n5753) );
  AOI22_X1 U5292 ( .A1(n5549), .A2(n5753), .B1(n5535), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4224) );
  OAI21_X1 U5293 ( .B1(n5555), .B2(n4467), .A(n4224), .ZN(U2858) );
  INV_X1 U5294 ( .A(n6275), .ZN(n4339) );
  NAND2_X1 U5295 ( .A1(n6282), .A2(n4339), .ZN(n4228) );
  INV_X1 U5296 ( .A(n4225), .ZN(n4226) );
  OR2_X1 U5297 ( .A1(n4370), .A2(n4226), .ZN(n4227) );
  NAND2_X1 U5298 ( .A1(n4228), .A2(n4227), .ZN(n4293) );
  INV_X1 U5299 ( .A(n4293), .ZN(n4237) );
  OR2_X1 U5300 ( .A1(n5075), .A2(n6321), .ZN(n4230) );
  AOI21_X1 U5301 ( .B1(n4230), .B2(n3091), .A(n4229), .ZN(n4235) );
  NAND3_X1 U5302 ( .A1(n4233), .A2(n4232), .A3(n4231), .ZN(n4234) );
  AOI21_X1 U5303 ( .B1(n6282), .B2(n4235), .A(n4234), .ZN(n4236) );
  NAND2_X1 U5304 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n5074) );
  NOR2_X1 U5305 ( .A1(n6303), .A2(n5074), .ZN(n6312) );
  AOI22_X1 U5306 ( .A1(n6293), .A2(n6266), .B1(FLUSH_REG_SCAN_IN), .B2(n6312), 
        .ZN(n5356) );
  NAND2_X1 U5307 ( .A1(n6303), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U5308 ( .A1(n5356), .A2(n6382), .ZN(n6394) );
  OAI21_X1 U5309 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6386), .A(n6394), 
        .ZN(n6392) );
  INV_X1 U5310 ( .A(n6392), .ZN(n4254) );
  INV_X1 U5311 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4238) );
  AOI22_X1 U5312 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4238), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5759), .ZN(n4679) );
  NOR2_X1 U5313 ( .A1(n6431), .A2(n6679), .ZN(n4251) );
  AND4_X1 U5314 ( .A1(n4243), .A2(n4242), .A3(n4241), .A4(n4240), .ZN(n4245)
         );
  NAND3_X1 U5315 ( .A1(n4370), .A2(n4245), .A3(n4244), .ZN(n4246) );
  OR2_X1 U5316 ( .A1(n4247), .A2(n4246), .ZN(n6262) );
  INV_X1 U5317 ( .A(n6262), .ZN(n4347) );
  NOR2_X1 U5318 ( .A1(n5075), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4342)
         );
  INV_X1 U5319 ( .A(n4342), .ZN(n4250) );
  INV_X1 U5320 ( .A(n4681), .ZN(n4678) );
  INV_X1 U5321 ( .A(n4248), .ZN(n4365) );
  NAND3_X1 U5322 ( .A1(n6261), .A2(n4678), .A3(n4365), .ZN(n4249) );
  OAI211_X1 U5323 ( .C1(n4239), .C2(n4347), .A(n4250), .B(n4249), .ZN(n6265)
         );
  INV_X1 U5324 ( .A(n6396), .ZN(n5357) );
  AOI222_X1 U5325 ( .A1(n4680), .A2(n4252), .B1(n4679), .B2(n4251), .C1(n6265), 
        .C2(n5357), .ZN(n4253) );
  OAI22_X1 U5326 ( .A1(n4254), .A2(n3237), .B1(n6389), .B2(n4253), .ZN(U3460)
         );
  NAND2_X1 U5327 ( .A1(n4255), .A2(n4256), .ZN(n4257) );
  AND2_X1 U5328 ( .A1(n4317), .A2(n4257), .ZN(n5737) );
  INV_X1 U5329 ( .A(n5737), .ZN(n4262) );
  INV_X1 U5330 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6499) );
  OR2_X1 U5331 ( .A1(n4258), .A2(n4259), .ZN(n4261) );
  NAND2_X1 U5332 ( .A1(n4261), .A2(n4315), .ZN(n5501) );
  OAI222_X1 U5333 ( .A1(n4262), .A2(n5553), .B1(n5554), .B2(n6499), .C1(n5501), 
        .C2(n5555), .ZN(U2856) );
  INV_X1 U5334 ( .A(n4379), .ZN(n4264) );
  INV_X1 U5335 ( .A(n5986), .ZN(n4265) );
  NAND2_X1 U5336 ( .A1(n5922), .A2(n4265), .ZN(n4266) );
  NAND2_X1 U5337 ( .A1(n4266), .A2(n6432), .ZN(n4276) );
  INV_X1 U5338 ( .A(n4239), .ZN(n5896) );
  NOR2_X1 U5339 ( .A1(n5774), .A2(n5896), .ZN(n6114) );
  INV_X1 U5340 ( .A(n4268), .ZN(n4368) );
  NAND2_X1 U5341 ( .A1(n6114), .A2(n4368), .ZN(n4418) );
  OR2_X1 U5342 ( .A1(n4418), .A2(n5805), .ZN(n4270) );
  NAND3_X1 U5343 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6734), .A3(n6667), .ZN(n4413) );
  NOR2_X1 U5344 ( .A1(n6113), .A2(n4413), .ZN(n5890) );
  INV_X1 U5345 ( .A(n5890), .ZN(n4269) );
  NAND2_X1 U5346 ( .A1(n4270), .A2(n4269), .ZN(n4277) );
  INV_X1 U5347 ( .A(n4277), .ZN(n4271) );
  OR2_X1 U5348 ( .A1(n4276), .A2(n4271), .ZN(n4274) );
  INV_X1 U5349 ( .A(n4413), .ZN(n4272) );
  NAND2_X1 U5350 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4272), .ZN(n4273) );
  NAND2_X1 U5351 ( .A1(n4274), .A2(n4273), .ZN(n5891) );
  INV_X1 U5352 ( .A(n5891), .ZN(n4493) );
  INV_X1 U5353 ( .A(DATAI_1_), .ZN(n4307) );
  NOR2_X2 U5354 ( .A1(n4307), .A2(n5961), .ZN(n6213) );
  INV_X1 U5355 ( .A(n6213), .ZN(n4286) );
  AOI21_X1 U5356 ( .B1(n4413), .B2(n6203), .A(n6202), .ZN(n4275) );
  OAI21_X1 U5357 ( .B1(n4277), .B2(n4276), .A(n4275), .ZN(n5892) );
  NAND2_X1 U5358 ( .A1(n5892), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4285) );
  NOR2_X2 U5359 ( .A1(n4587), .A2(n4279), .ZN(n6214) );
  INV_X1 U5360 ( .A(DATAI_17_), .ZN(n4280) );
  NOR2_X1 U5361 ( .A1(n5682), .A2(n4280), .ZN(n6126) );
  INV_X1 U5362 ( .A(n6126), .ZN(n6218) );
  INV_X1 U5363 ( .A(n6121), .ZN(n4281) );
  INV_X1 U5364 ( .A(DATAI_25_), .ZN(n4282) );
  NOR2_X1 U5365 ( .A1(n5682), .A2(n4282), .ZN(n6215) );
  INV_X1 U5366 ( .A(n6215), .ZN(n6129) );
  OAI22_X1 U5367 ( .A1(n6218), .A2(n5898), .B1(n4488), .B2(n6129), .ZN(n4283)
         );
  AOI21_X1 U5368 ( .B1(n6214), .B2(n5890), .A(n4283), .ZN(n4284) );
  OAI211_X1 U5369 ( .C1(n4493), .C2(n4286), .A(n4285), .B(n4284), .ZN(U3061)
         );
  NOR2_X1 U5370 ( .A1(n3083), .A2(n4287), .ZN(n4289) );
  NOR2_X1 U5371 ( .A1(n4258), .A2(n4289), .ZN(n5668) );
  INV_X1 U5372 ( .A(n5668), .ZN(n4303) );
  INV_X1 U5373 ( .A(n3095), .ZN(n4290) );
  NOR2_X1 U5374 ( .A1(n4291), .A2(n4290), .ZN(n4292) );
  INV_X1 U5375 ( .A(n5604), .ZN(n4295) );
  NAND2_X1 U5376 ( .A1(n4297), .A2(n4301), .ZN(n4298) );
  INV_X1 U5377 ( .A(n4299), .ZN(n4300) );
  AND2_X1 U5378 ( .A1(n3084), .A2(n4301), .ZN(n4302) );
  INV_X1 U5379 ( .A(DATAI_2_), .ZN(n6616) );
  OAI222_X1 U5380 ( .A1(n4303), .A2(n5178), .B1(n5008), .B2(n6616), .C1(n5566), 
        .C2(n3359), .ZN(U2889) );
  INV_X1 U5381 ( .A(DATAI_3_), .ZN(n4585) );
  INV_X1 U5382 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5638) );
  OAI222_X1 U5383 ( .A1(n5501), .A2(n5178), .B1(n5008), .B2(n4585), .C1(n5566), 
        .C2(n5638), .ZN(U2888) );
  OAI21_X1 U5384 ( .B1(n4306), .B2(n4305), .A(n4304), .ZN(n5683) );
  INV_X1 U5385 ( .A(DATAI_0_), .ZN(n4333) );
  INV_X1 U5386 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5633) );
  OAI222_X1 U5387 ( .A1(n5683), .A2(n5178), .B1(n5008), .B2(n4333), .C1(n5566), 
        .C2(n5633), .ZN(U2891) );
  INV_X1 U5388 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5635) );
  OAI222_X1 U5389 ( .A1(n4467), .A2(n5178), .B1(n5008), .B2(n4307), .C1(n5566), 
        .C2(n5635), .ZN(U2890) );
  AND2_X1 U5390 ( .A1(n4308), .A2(n4309), .ZN(n4312) );
  CLKBUF_X1 U5391 ( .A(n4310), .Z(n4311) );
  OR2_X1 U5392 ( .A1(n4312), .A2(n4311), .ZN(n5470) );
  XNOR2_X1 U5393 ( .A(n4410), .B(n4406), .ZN(n5471) );
  AOI22_X1 U5394 ( .A1(n5549), .A2(n5471), .B1(n5535), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4313) );
  OAI21_X1 U5395 ( .B1(n5470), .B2(n5555), .A(n4313), .ZN(U2854) );
  INV_X1 U5396 ( .A(n4308), .ZN(n4314) );
  AOI21_X1 U5397 ( .B1(n4316), .B2(n4315), .A(n4314), .ZN(n5492) );
  INV_X1 U5398 ( .A(n5492), .ZN(n4332) );
  AOI21_X1 U5399 ( .B1(n4318), .B2(n4317), .A(n4410), .ZN(n5729) );
  AOI22_X1 U5400 ( .A1(n5549), .A2(n5729), .B1(n5535), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4319) );
  OAI21_X1 U5401 ( .B1(n4332), .B2(n5555), .A(n4319), .ZN(U2855) );
  XNOR2_X1 U5402 ( .A(n4321), .B(n4320), .ZN(n5734) );
  NOR2_X1 U5403 ( .A1(n5740), .A2(n6335), .ZN(n5736) );
  AOI21_X1 U5404 ( .B1(n5662), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5736), 
        .ZN(n4323) );
  OR2_X1 U5405 ( .A1(n5673), .A2(n5511), .ZN(n4322) );
  OAI211_X1 U5406 ( .C1(n5501), .C2(n5682), .A(n4323), .B(n4322), .ZN(n4324)
         );
  INV_X1 U5407 ( .A(n4324), .ZN(n4325) );
  OAI21_X1 U5408 ( .B1(n5734), .B2(n5371), .A(n4325), .ZN(U2983) );
  XNOR2_X1 U5409 ( .A(n4326), .B(n4327), .ZN(n5726) );
  INV_X1 U5410 ( .A(n4328), .ZN(n5485) );
  AOI22_X1 U5411 ( .A1(n5662), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n5348), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4329) );
  OAI21_X1 U5412 ( .B1(n5485), .B2(n5673), .A(n4329), .ZN(n4330) );
  AOI21_X1 U5413 ( .B1(n5492), .B2(n5669), .A(n4330), .ZN(n4331) );
  OAI21_X1 U5414 ( .B1(n5726), .B2(n5371), .A(n4331), .ZN(U2982) );
  INV_X1 U5415 ( .A(DATAI_4_), .ZN(n6678) );
  INV_X1 U5416 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5640) );
  OAI222_X1 U5417 ( .A1(n4332), .A2(n5178), .B1(n5008), .B2(n6678), .C1(n5566), 
        .C2(n5640), .ZN(U2887) );
  INV_X1 U5418 ( .A(DATAI_5_), .ZN(n4479) );
  OAI222_X1 U5419 ( .A1(n5470), .A2(n5178), .B1(n5008), .B2(n4479), .C1(n5566), 
        .C2(n3444), .ZN(U2886) );
  INV_X1 U5420 ( .A(n5892), .ZN(n4396) );
  INV_X1 U5421 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4338) );
  NOR2_X2 U5422 ( .A1(n4333), .A2(n5961), .ZN(n6196) );
  INV_X1 U5423 ( .A(DATAI_16_), .ZN(n6597) );
  NOR2_X1 U5424 ( .A1(n5682), .A2(n6597), .ZN(n6122) );
  INV_X1 U5425 ( .A(n6122), .ZN(n6212) );
  INV_X1 U5426 ( .A(DATAI_24_), .ZN(n4850) );
  NOR2_X1 U5427 ( .A1(n5682), .A2(n4850), .ZN(n6209) );
  NOR2_X2 U5428 ( .A1(n4334), .A2(n4587), .ZN(n6197) );
  AOI22_X1 U5429 ( .A1(n5889), .A2(n6209), .B1(n6197), .B2(n5890), .ZN(n4335)
         );
  OAI21_X1 U5430 ( .B1(n5898), .B2(n6212), .A(n4335), .ZN(n4336) );
  AOI21_X1 U5431 ( .B1(n6196), .B2(n5891), .A(n4336), .ZN(n4337) );
  OAI21_X1 U5432 ( .B1(n4396), .B2(n4338), .A(n4337), .ZN(U3060) );
  OR2_X1 U5433 ( .A1(n6278), .A2(n4339), .ZN(n4357) );
  INV_X1 U5434 ( .A(n4353), .ZN(n4341) );
  MUX2_X1 U5435 ( .A(n4357), .B(n4341), .S(n4681), .Z(n4340) );
  AOI21_X1 U5436 ( .B1(n6264), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4340), 
        .ZN(n4345) );
  MUX2_X1 U5437 ( .A(n4341), .B(n4357), .S(n4681), .Z(n4343) );
  NOR2_X1 U5438 ( .A1(n4343), .A2(n4342), .ZN(n4344) );
  MUX2_X1 U5439 ( .A(n4345), .B(n4344), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n4346) );
  OAI21_X1 U5440 ( .B1(n4347), .B2(n5774), .A(n4346), .ZN(n4684) );
  INV_X1 U5441 ( .A(n6266), .ZN(n4348) );
  MUX2_X1 U5442 ( .A(n4684), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(n4348), 
        .Z(n6270) );
  NAND2_X1 U5443 ( .A1(n6431), .A2(n6270), .ZN(n4364) );
  OR2_X1 U5444 ( .A1(n6266), .A2(n3109), .ZN(n4361) );
  NAND2_X1 U5445 ( .A1(n6017), .A2(n6262), .ZN(n4359) );
  NOR2_X1 U5446 ( .A1(n4681), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4350)
         );
  XNOR2_X1 U5447 ( .A(n4350), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4356)
         );
  NAND2_X1 U5448 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4351) );
  XOR2_X1 U5449 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n4351), .Z(n4354) );
  AOI21_X1 U5450 ( .B1(n4681), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3109), 
        .ZN(n4352) );
  NOR2_X1 U5451 ( .A1(n4773), .A2(n4352), .ZN(n6387) );
  OAI22_X1 U5452 ( .A1(n5075), .A2(n4354), .B1(n6387), .B2(n4353), .ZN(n4355)
         );
  AOI21_X1 U5453 ( .B1(n4357), .B2(n4356), .A(n4355), .ZN(n4358) );
  NAND2_X1 U5454 ( .A1(n4359), .A2(n4358), .ZN(n6385) );
  NAND2_X1 U5455 ( .A1(n6266), .A2(n6385), .ZN(n4360) );
  INV_X1 U5456 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5372) );
  NAND2_X1 U5457 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5372), .ZN(n4366) );
  INV_X1 U5458 ( .A(n4362), .ZN(n4363) );
  OAI22_X1 U5459 ( .A1(n4364), .A2(n6271), .B1(n4366), .B2(n4363), .ZN(n6288)
         );
  NAND2_X1 U5460 ( .A1(n6288), .A2(n4365), .ZN(n4376) );
  OAI21_X1 U5461 ( .B1(n6266), .B2(STATE2_REG_1__SCAN_IN), .A(n4366), .ZN(
        n4367) );
  NAND2_X1 U5462 ( .A1(n4367), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4372) );
  NOR2_X1 U5463 ( .A1(n3364), .A2(n4368), .ZN(n4369) );
  XNOR2_X1 U5464 ( .A(n4369), .B(n6586), .ZN(n5482) );
  INV_X1 U5465 ( .A(n4370), .ZN(n5358) );
  NAND3_X1 U5466 ( .A1(n5482), .A2(n5358), .A3(n6431), .ZN(n4371) );
  NAND3_X1 U5467 ( .A1(n4376), .A2(n6286), .A3(n5372), .ZN(n4373) );
  NAND2_X1 U5468 ( .A1(n4373), .A2(n6312), .ZN(n4374) );
  INV_X1 U5469 ( .A(n5074), .ZN(n4375) );
  AND3_X1 U5470 ( .A1(n4376), .A2(n6286), .A3(n4375), .ZN(n6299) );
  NOR2_X1 U5471 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6431), .ZN(n6399) );
  OAI22_X1 U5472 ( .A1(n5777), .A2(n6203), .B1(n5805), .B2(n6399), .ZN(n4377)
         );
  OAI21_X1 U5473 ( .B1(n6299), .B2(n4377), .A(n6403), .ZN(n4378) );
  OAI21_X1 U5474 ( .B1(n6403), .B2(n6113), .A(n4378), .ZN(U3465) );
  NAND2_X1 U5475 ( .A1(n4263), .A2(n4379), .ZN(n6159) );
  OR2_X1 U5476 ( .A1(n5986), .A2(n6159), .ZN(n6116) );
  AND2_X1 U5477 ( .A1(n6116), .A2(n6049), .ZN(n4570) );
  NAND2_X1 U5478 ( .A1(n3096), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6398) );
  INV_X1 U5479 ( .A(n6398), .ZN(n6050) );
  NAND2_X1 U5480 ( .A1(n5922), .A2(n6050), .ZN(n5923) );
  AOI21_X1 U5481 ( .B1(n4570), .B2(n5923), .A(n6203), .ZN(n4382) );
  INV_X1 U5482 ( .A(n4380), .ZN(n4415) );
  NAND2_X1 U5483 ( .A1(n6432), .A2(n6164), .ZN(n6199) );
  INV_X1 U5484 ( .A(n6017), .ZN(n5924) );
  OAI22_X1 U5485 ( .A1(n4415), .A2(n6199), .B1(n5924), .B2(n6399), .ZN(n4381)
         );
  OAI21_X1 U5486 ( .B1(n4382), .B2(n4381), .A(n6403), .ZN(n4383) );
  OAI21_X1 U5487 ( .B1(n6403), .B2(n6734), .A(n4383), .ZN(U3462) );
  OAI21_X1 U5488 ( .B1(n4386), .B2(n4385), .A(n4384), .ZN(n5755) );
  INV_X1 U5489 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4463) );
  NOR2_X1 U5490 ( .A1(n4467), .A2(n5682), .ZN(n4388) );
  OAI22_X1 U5491 ( .A1(n5676), .A2(n4463), .B1(n5740), .B2(n6407), .ZN(n4387)
         );
  AOI211_X1 U5492 ( .C1(n5233), .C2(n4463), .A(n4388), .B(n4387), .ZN(n4389)
         );
  OAI21_X1 U5493 ( .B1(n5755), .B2(n5371), .A(n4389), .ZN(U2985) );
  INV_X1 U5494 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4395) );
  NOR2_X2 U5495 ( .A1(n4587), .A2(n4390), .ZN(n6232) );
  INV_X1 U5496 ( .A(DATAI_20_), .ZN(n4391) );
  NOR2_X1 U5497 ( .A1(n5682), .A2(n4391), .ZN(n6138) );
  INV_X1 U5498 ( .A(n6138), .ZN(n6236) );
  INV_X1 U5499 ( .A(DATAI_28_), .ZN(n5176) );
  NOR2_X1 U5500 ( .A1(n5682), .A2(n5176), .ZN(n6233) );
  INV_X1 U5501 ( .A(n6233), .ZN(n6141) );
  OAI22_X1 U5502 ( .A1(n6236), .A2(n5898), .B1(n4488), .B2(n6141), .ZN(n4392)
         );
  AOI21_X1 U5503 ( .B1(n6232), .B2(n5890), .A(n4392), .ZN(n4394) );
  NOR2_X2 U5504 ( .A1(n6678), .A2(n5961), .ZN(n6231) );
  NAND2_X1 U5505 ( .A1(n5891), .A2(n6231), .ZN(n4393) );
  OAI211_X1 U5506 ( .C1(n4396), .C2(n4395), .A(n4394), .B(n4393), .ZN(U3064)
         );
  XNOR2_X1 U5507 ( .A(n4397), .B(n4398), .ZN(n4471) );
  INV_X1 U5508 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6339) );
  NOR2_X1 U5509 ( .A1(n5740), .A2(n6339), .ZN(n4473) );
  AOI21_X1 U5510 ( .B1(n5662), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4473), 
        .ZN(n4400) );
  OR2_X1 U5511 ( .A1(n5673), .A2(n5481), .ZN(n4399) );
  OAI211_X1 U5512 ( .C1(n5470), .C2(n5682), .A(n4400), .B(n4399), .ZN(n4401)
         );
  INV_X1 U5513 ( .A(n4401), .ZN(n4402) );
  OAI21_X1 U5514 ( .B1(n4471), .B2(n5371), .A(n4402), .ZN(U2981) );
  NOR2_X1 U5515 ( .A1(n4311), .A2(n4404), .ZN(n4405) );
  OR2_X1 U5516 ( .A1(n4403), .A2(n4405), .ZN(n5463) );
  INV_X1 U5517 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4412) );
  INV_X1 U5518 ( .A(n4406), .ZN(n4409) );
  INV_X1 U5519 ( .A(n4407), .ZN(n4408) );
  AOI21_X1 U5520 ( .B1(n4410), .B2(n4409), .A(n4408), .ZN(n4411) );
  OR2_X1 U5521 ( .A1(n4433), .A2(n4411), .ZN(n5460) );
  OAI222_X1 U5522 ( .A1(n5463), .A2(n5555), .B1(n4412), .B2(n5554), .C1(n5553), 
        .C2(n5460), .ZN(U2853) );
  INV_X1 U5523 ( .A(DATAI_6_), .ZN(n6645) );
  OAI222_X1 U5524 ( .A1(n5463), .A2(n5178), .B1(n5008), .B2(n6645), .C1(n5566), 
        .C2(n3462), .ZN(U2885) );
  NOR2_X1 U5525 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4413), .ZN(n5880)
         );
  NAND3_X1 U5526 ( .A1(n4488), .A2(n6432), .A3(n5884), .ZN(n4416) );
  NAND2_X1 U5527 ( .A1(n4416), .A2(n6199), .ZN(n4419) );
  INV_X1 U5528 ( .A(n4421), .ZN(n4417) );
  NOR2_X1 U5529 ( .A1(n4417), .A2(n6550), .ZN(n6170) );
  INV_X1 U5530 ( .A(n6160), .ZN(n5956) );
  AND2_X1 U5531 ( .A1(n5955), .A2(n5956), .ZN(n5775) );
  OAI21_X1 U5532 ( .B1(n5775), .B2(n6550), .A(n5841), .ZN(n5778) );
  AOI211_X1 U5533 ( .C1(n4419), .C2(n4418), .A(n6170), .B(n5778), .ZN(n4420)
         );
  OAI21_X1 U5534 ( .B1(n5880), .B2(n6384), .A(n4420), .ZN(n5881) );
  INV_X1 U5535 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4427) );
  INV_X1 U5536 ( .A(n6209), .ZN(n6125) );
  NOR2_X1 U5537 ( .A1(n6017), .A2(n6203), .ZN(n5773) );
  NAND2_X1 U5538 ( .A1(n5773), .A2(n6114), .ZN(n4423) );
  NOR2_X1 U5539 ( .A1(n4421), .A2(n6550), .ZN(n6161) );
  NAND2_X1 U5540 ( .A1(n5775), .A2(n6161), .ZN(n4422) );
  NAND2_X1 U5541 ( .A1(n4423), .A2(n4422), .ZN(n5879) );
  AOI22_X1 U5542 ( .A1(n5879), .A2(n6196), .B1(n6197), .B2(n5880), .ZN(n4424)
         );
  OAI21_X1 U5543 ( .B1(n5884), .B2(n6125), .A(n4424), .ZN(n4425) );
  AOI21_X1 U5544 ( .B1(n5889), .B2(n6122), .A(n4425), .ZN(n4426) );
  OAI21_X1 U5545 ( .B1(n4500), .B2(n4427), .A(n4426), .ZN(U3052) );
  NOR2_X1 U5546 ( .A1(n4403), .A2(n4429), .ZN(n4430) );
  OR2_X1 U5547 ( .A1(n4428), .A2(n4430), .ZN(n5453) );
  OR2_X1 U5548 ( .A1(n4433), .A2(n4432), .ZN(n4434) );
  NAND2_X1 U5549 ( .A1(n4431), .A2(n4434), .ZN(n5712) );
  INV_X1 U5550 ( .A(n5712), .ZN(n4435) );
  AOI22_X1 U5551 ( .A1(n5549), .A2(n4435), .B1(n5535), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4436) );
  OAI21_X1 U5552 ( .B1(n5453), .B2(n5555), .A(n4436), .ZN(U2852) );
  INV_X1 U5553 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4441) );
  INV_X1 U5554 ( .A(DATAI_31_), .ZN(n4437) );
  NOR2_X1 U5555 ( .A1(n5682), .A2(n4437), .ZN(n6254) );
  INV_X1 U5556 ( .A(DATAI_7_), .ZN(n4454) );
  NOR2_X2 U5557 ( .A1(n4454), .A2(n5961), .ZN(n6250) );
  AOI22_X1 U5558 ( .A1(n4590), .A2(n6254), .B1(n6250), .B2(n5879), .ZN(n4440)
         );
  NOR2_X2 U5559 ( .A1(n4587), .A2(n4916), .ZN(n6251) );
  INV_X1 U5560 ( .A(DATAI_23_), .ZN(n4438) );
  NOR2_X1 U5561 ( .A1(n5682), .A2(n4438), .ZN(n6152) );
  AOI22_X1 U5562 ( .A1(n6251), .A2(n5880), .B1(n5889), .B2(n6152), .ZN(n4439)
         );
  OAI211_X1 U5563 ( .C1(n4500), .C2(n4441), .A(n4440), .B(n4439), .ZN(U3059)
         );
  INV_X1 U5564 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4444) );
  AOI22_X1 U5565 ( .A1(n4590), .A2(n6233), .B1(n6231), .B2(n5879), .ZN(n4443)
         );
  AOI22_X1 U5566 ( .A1(n6232), .A2(n5880), .B1(n5889), .B2(n6138), .ZN(n4442)
         );
  OAI211_X1 U5567 ( .C1(n4500), .C2(n4444), .A(n4443), .B(n4442), .ZN(U3056)
         );
  INV_X1 U5568 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4450) );
  INV_X1 U5569 ( .A(DATAI_26_), .ZN(n4445) );
  NOR2_X1 U5570 ( .A1(n5682), .A2(n4445), .ZN(n6221) );
  NOR2_X2 U5571 ( .A1(n6616), .A2(n5961), .ZN(n6219) );
  AOI22_X1 U5572 ( .A1(n4590), .A2(n6221), .B1(n6219), .B2(n5879), .ZN(n4449)
         );
  NOR2_X2 U5573 ( .A1(n4587), .A2(n4446), .ZN(n6220) );
  INV_X1 U5574 ( .A(DATAI_18_), .ZN(n4447) );
  NOR2_X1 U5575 ( .A1(n5682), .A2(n4447), .ZN(n6130) );
  AOI22_X1 U5576 ( .A1(n6220), .A2(n5880), .B1(n5889), .B2(n6130), .ZN(n4448)
         );
  OAI211_X1 U5577 ( .C1(n4500), .C2(n4450), .A(n4449), .B(n4448), .ZN(U3054)
         );
  INV_X1 U5578 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4453) );
  AOI22_X1 U5579 ( .A1(n4590), .A2(n6215), .B1(n6213), .B2(n5879), .ZN(n4452)
         );
  AOI22_X1 U5580 ( .A1(n6214), .A2(n5880), .B1(n5889), .B2(n6126), .ZN(n4451)
         );
  OAI211_X1 U5581 ( .C1(n4500), .C2(n4453), .A(n4452), .B(n4451), .ZN(U3053)
         );
  INV_X1 U5582 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5644) );
  OAI222_X1 U5583 ( .A1(n5453), .A2(n5178), .B1(n5008), .B2(n4454), .C1(n5566), 
        .C2(n5644), .ZN(U2884) );
  OAI21_X1 U5584 ( .B1(n4428), .B2(n4456), .A(n4455), .ZN(n5440) );
  INV_X1 U5585 ( .A(n4516), .ZN(n4547) );
  AOI21_X1 U5586 ( .B1(n4457), .B2(n4431), .A(n4547), .ZN(n5701) );
  AOI22_X1 U5587 ( .A1(n5549), .A2(n5701), .B1(n5535), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4458) );
  OAI21_X1 U5588 ( .B1(n5440), .B2(n5555), .A(n4458), .ZN(U2851) );
  AOI22_X1 U5589 ( .A1(n5562), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n5558), .ZN(n4459) );
  OAI21_X1 U5590 ( .B1(n5440), .B2(n5178), .A(n4459), .ZN(U2883) );
  NAND2_X1 U5591 ( .A1(n4895), .A2(n3095), .ZN(n4460) );
  NAND2_X1 U5592 ( .A1(n4460), .A2(n5452), .ZN(n5523) );
  INV_X1 U5593 ( .A(n5523), .ZN(n4561) );
  AOI22_X1 U5594 ( .A1(EBX_REG_1__SCAN_IN), .A2(n5518), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5519), .ZN(n4461) );
  OAI221_X1 U5595 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5487), .C1(n6407), .C2(
        n5486), .A(n4461), .ZN(n4462) );
  AOI21_X1 U5596 ( .B1(n5520), .B2(n4463), .A(n4462), .ZN(n4466) );
  AND2_X1 U5597 ( .A1(n4895), .A2(n4464), .ZN(n5522) );
  AOI22_X1 U5598 ( .A1(n5896), .A2(n5522), .B1(n5517), .B2(n5753), .ZN(n4465)
         );
  OAI211_X1 U5599 ( .C1(n4561), .C2(n4467), .A(n4466), .B(n4465), .ZN(U2826)
         );
  AOI21_X1 U5600 ( .B1(n5721), .B2(n4468), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n4470) );
  NAND2_X1 U5601 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4538) );
  INV_X1 U5602 ( .A(n4649), .ZN(n4535) );
  AOI21_X1 U5603 ( .B1(n4647), .B2(n4538), .A(n4535), .ZN(n4469) );
  INV_X1 U5604 ( .A(n4469), .ZN(n5748) );
  AOI21_X1 U5605 ( .B1(n4537), .B2(n5757), .A(n5748), .ZN(n5720) );
  OAI22_X1 U5606 ( .A1(n4471), .A2(n5733), .B1(n4470), .B2(n5720), .ZN(n4472)
         );
  AOI211_X1 U5607 ( .C1(n5754), .C2(n5471), .A(n4473), .B(n4472), .ZN(n4478)
         );
  INV_X1 U5608 ( .A(n5752), .ZN(n4476) );
  INV_X1 U5609 ( .A(n4474), .ZN(n4475) );
  NAND3_X1 U5610 ( .A1(n4476), .A2(n4130), .A3(n4475), .ZN(n4477) );
  NAND2_X1 U5611 ( .A1(n4478), .A2(n4477), .ZN(U3013) );
  NOR2_X2 U5612 ( .A1(n4479), .A2(n5961), .ZN(n6237) );
  INV_X1 U5613 ( .A(n6237), .ZN(n4484) );
  NAND2_X1 U5614 ( .A1(n5892), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4483) );
  NOR2_X2 U5615 ( .A1(n4587), .A2(n3084), .ZN(n6238) );
  INV_X1 U5616 ( .A(DATAI_21_), .ZN(n6663) );
  NOR2_X1 U5617 ( .A1(n5682), .A2(n6663), .ZN(n6142) );
  INV_X1 U5618 ( .A(n6142), .ZN(n6242) );
  INV_X1 U5619 ( .A(DATAI_29_), .ZN(n4480) );
  NOR2_X1 U5620 ( .A1(n5682), .A2(n4480), .ZN(n6239) );
  INV_X1 U5621 ( .A(n6239), .ZN(n6145) );
  OAI22_X1 U5622 ( .A1(n6242), .A2(n5898), .B1(n4488), .B2(n6145), .ZN(n4481)
         );
  AOI21_X1 U5623 ( .B1(n6238), .B2(n5890), .A(n4481), .ZN(n4482) );
  OAI211_X1 U5624 ( .C1(n4493), .C2(n4484), .A(n4483), .B(n4482), .ZN(U3065)
         );
  NOR2_X2 U5625 ( .A1(n6645), .A2(n5961), .ZN(n6243) );
  INV_X1 U5626 ( .A(n6243), .ZN(n4492) );
  NAND2_X1 U5627 ( .A1(n5892), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4491) );
  NOR2_X2 U5628 ( .A1(n4587), .A2(n4485), .ZN(n6244) );
  INV_X1 U5629 ( .A(DATAI_22_), .ZN(n4486) );
  NOR2_X1 U5630 ( .A1(n5682), .A2(n4486), .ZN(n6146) );
  INV_X1 U5631 ( .A(n6146), .ZN(n6248) );
  INV_X1 U5632 ( .A(DATAI_30_), .ZN(n4487) );
  NOR2_X1 U5633 ( .A1(n5682), .A2(n4487), .ZN(n6245) );
  INV_X1 U5634 ( .A(n6245), .ZN(n6149) );
  OAI22_X1 U5635 ( .A1(n6248), .A2(n5898), .B1(n4488), .B2(n6149), .ZN(n4489)
         );
  AOI21_X1 U5636 ( .B1(n6244), .B2(n5890), .A(n4489), .ZN(n4490) );
  OAI211_X1 U5637 ( .C1(n4493), .C2(n4492), .A(n4491), .B(n4490), .ZN(U3066)
         );
  INV_X1 U5638 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4496) );
  AOI22_X1 U5639 ( .A1(n4590), .A2(n6245), .B1(n6243), .B2(n5879), .ZN(n4495)
         );
  AOI22_X1 U5640 ( .A1(n6244), .A2(n5880), .B1(n5889), .B2(n6146), .ZN(n4494)
         );
  OAI211_X1 U5641 ( .C1(n4500), .C2(n4496), .A(n4495), .B(n4494), .ZN(U3058)
         );
  INV_X1 U5642 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4499) );
  AOI22_X1 U5643 ( .A1(n4590), .A2(n6239), .B1(n6237), .B2(n5879), .ZN(n4498)
         );
  AOI22_X1 U5644 ( .A1(n6238), .A2(n5880), .B1(n5889), .B2(n6142), .ZN(n4497)
         );
  OAI211_X1 U5645 ( .C1(n4500), .C2(n4499), .A(n4498), .B(n4497), .ZN(U3057)
         );
  XNOR2_X1 U5646 ( .A(n4501), .B(n4502), .ZN(n5706) );
  INV_X1 U5647 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6340) );
  NOR2_X1 U5648 ( .A1(n5740), .A2(n6340), .ZN(n5709) );
  AOI21_X1 U5649 ( .B1(n5662), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5709), 
        .ZN(n4504) );
  OR2_X1 U5650 ( .A1(n5673), .A2(n5451), .ZN(n4503) );
  OAI211_X1 U5651 ( .C1(n5453), .C2(n5682), .A(n4504), .B(n4503), .ZN(n4505)
         );
  INV_X1 U5652 ( .A(n4505), .ZN(n4506) );
  OAI21_X1 U5653 ( .B1(n5706), .B2(n5371), .A(n4506), .ZN(U2979) );
  XNOR2_X1 U5654 ( .A(n4507), .B(n4508), .ZN(n5714) );
  INV_X1 U5655 ( .A(REIP_REG_6__SCAN_IN), .ZN(n4509) );
  OAI22_X1 U5656 ( .A1(n5676), .A2(n6711), .B1(n5740), .B2(n4509), .ZN(n4511)
         );
  NOR2_X1 U5657 ( .A1(n5463), .A2(n5682), .ZN(n4510) );
  AOI211_X1 U5658 ( .C1(n5233), .C2(n5464), .A(n4511), .B(n4510), .ZN(n4512)
         );
  OAI21_X1 U5659 ( .B1(n5714), .B2(n5371), .A(n4512), .ZN(U2980) );
  NAND2_X1 U5660 ( .A1(n4455), .A2(n4514), .ZN(n4515) );
  NAND2_X1 U5661 ( .A1(n4599), .A2(n4515), .ZN(n5435) );
  XNOR2_X1 U5662 ( .A(n4516), .B(n4546), .ZN(n5691) );
  AOI22_X1 U5663 ( .A1(n5549), .A2(n5691), .B1(n5535), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n4517) );
  OAI21_X1 U5664 ( .B1(n5435), .B2(n5555), .A(n4517), .ZN(U2850) );
  INV_X1 U5665 ( .A(DATAI_9_), .ZN(n4518) );
  INV_X1 U5666 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6568) );
  OAI222_X1 U5667 ( .A1(n5435), .A2(n5178), .B1(n5008), .B2(n4518), .C1(n5566), 
        .C2(n6568), .ZN(U2882) );
  XNOR2_X1 U5668 ( .A(n5054), .B(n4542), .ZN(n4520) );
  XNOR2_X1 U5669 ( .A(n4519), .B(n4520), .ZN(n5693) );
  NAND2_X1 U5670 ( .A1(n5693), .A2(n5679), .ZN(n4525) );
  INV_X1 U5671 ( .A(n5434), .ZN(n4523) );
  INV_X1 U5672 ( .A(REIP_REG_9__SCAN_IN), .ZN(n4521) );
  OAI22_X1 U5673 ( .A1(n5676), .A2(n6638), .B1(n5740), .B2(n4521), .ZN(n4522)
         );
  AOI21_X1 U5674 ( .B1(n5233), .B2(n4523), .A(n4522), .ZN(n4524) );
  OAI211_X1 U5675 ( .C1(n5682), .C2(n5435), .A(n4525), .B(n4524), .ZN(U2977)
         );
  INV_X1 U5676 ( .A(n4526), .ZN(n4528) );
  NAND2_X1 U5677 ( .A1(n4528), .A2(n4527), .ZN(n4529) );
  XNOR2_X1 U5678 ( .A(n4530), .B(n4529), .ZN(n4607) );
  INV_X1 U5679 ( .A(n5702), .ZN(n4540) );
  OAI22_X1 U5680 ( .A1(n4533), .A2(n5741), .B1(n4532), .B2(n4531), .ZN(n4534)
         );
  NOR2_X1 U5681 ( .A1(n4535), .A2(n4534), .ZN(n5705) );
  OAI21_X1 U5682 ( .B1(n4540), .B2(n4536), .A(n5705), .ZN(n5692) );
  INV_X1 U5683 ( .A(n4537), .ZN(n4539) );
  OAI21_X1 U5684 ( .B1(n5752), .B2(n4538), .A(n5741), .ZN(n5724) );
  NAND2_X1 U5685 ( .A1(n4539), .A2(n5724), .ZN(n5713) );
  NOR2_X1 U5686 ( .A1(n5719), .A2(n5713), .ZN(n5708) );
  NAND2_X1 U5687 ( .A1(n4540), .A2(n5708), .ZN(n5696) );
  AOI21_X1 U5688 ( .B1(n4542), .B2(n4541), .A(n5696), .ZN(n4544) );
  AOI22_X1 U5689 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5692), .B1(n4544), .B2(n4543), .ZN(n4551) );
  AOI21_X1 U5690 ( .B1(n4547), .B2(n4546), .A(n4545), .ZN(n4549) );
  INV_X1 U5691 ( .A(n4613), .ZN(n4548) );
  NOR2_X1 U5692 ( .A1(n4549), .A2(n4548), .ZN(n5545) );
  AND2_X1 U5693 ( .A1(n5348), .A2(REIP_REG_10__SCAN_IN), .ZN(n4604) );
  AOI21_X1 U5694 ( .B1(n5754), .B2(n5545), .A(n4604), .ZN(n4550) );
  OAI211_X1 U5695 ( .C1(n4607), .C2(n5733), .A(n4551), .B(n4550), .ZN(U3008)
         );
  INV_X1 U5696 ( .A(n5805), .ZN(n6263) );
  INV_X1 U5697 ( .A(n4552), .ZN(n4553) );
  OAI21_X1 U5698 ( .B1(n4554), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4553), 
        .ZN(n5772) );
  OAI22_X1 U5699 ( .A1(n3885), .A2(n5505), .B1(n5449), .B2(n5772), .ZN(n4557)
         );
  INV_X1 U5700 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4555) );
  AOI21_X1 U5701 ( .B1(n5499), .B2(n5512), .A(n4555), .ZN(n4556) );
  AOI211_X1 U5702 ( .C1(n5522), .C2(n6263), .A(n4557), .B(n4556), .ZN(n4560)
         );
  NAND2_X1 U5703 ( .A1(n4558), .A2(REIP_REG_0__SCAN_IN), .ZN(n4559) );
  OAI211_X1 U5704 ( .C1(n4561), .C2(n5683), .A(n4560), .B(n4559), .ZN(U2827)
         );
  XNOR2_X1 U5705 ( .A(n4562), .B(n4563), .ZN(n5698) );
  INV_X1 U5706 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4565) );
  INV_X1 U5707 ( .A(REIP_REG_8__SCAN_IN), .ZN(n4564) );
  OAI22_X1 U5708 ( .A1(n5676), .A2(n4565), .B1(n5740), .B2(n4564), .ZN(n4567)
         );
  NOR2_X1 U5709 ( .A1(n5440), .A2(n5682), .ZN(n4566) );
  AOI211_X1 U5710 ( .C1(n5233), .C2(n5441), .A(n4567), .B(n4566), .ZN(n4568)
         );
  OAI21_X1 U5711 ( .B1(n5698), .B2(n5371), .A(n4568), .ZN(U2978) );
  NOR2_X1 U5712 ( .A1(n4263), .A2(n6398), .ZN(n4569) );
  AOI21_X1 U5713 ( .B1(n4570), .B2(n4569), .A(n6203), .ZN(n4576) );
  NAND2_X1 U5714 ( .A1(n5774), .A2(n5896), .ZN(n6016) );
  NOR2_X1 U5715 ( .A1(n6017), .A2(n6016), .ZN(n5836) );
  NAND2_X1 U5716 ( .A1(n5836), .A2(n6263), .ZN(n4572) );
  INV_X1 U5717 ( .A(n6048), .ZN(n4571) );
  NAND2_X1 U5718 ( .A1(n4571), .A2(n6734), .ZN(n4592) );
  NAND2_X1 U5719 ( .A1(n4572), .A2(n4592), .ZN(n4578) );
  NAND2_X1 U5720 ( .A1(n4576), .A2(n4578), .ZN(n4575) );
  NAND3_X1 U5721 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6734), .A3(n6405), .ZN(n5835) );
  INV_X1 U5722 ( .A(n5835), .ZN(n4573) );
  NAND2_X1 U5723 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4573), .ZN(n4574) );
  NAND2_X1 U5724 ( .A1(n4575), .A2(n4574), .ZN(n5875) );
  INV_X1 U5725 ( .A(n5875), .ZN(n4597) );
  INV_X1 U5726 ( .A(n6196), .ZN(n4584) );
  INV_X1 U5727 ( .A(n4576), .ZN(n4579) );
  AOI21_X1 U5728 ( .B1(n5835), .B2(n6203), .A(n6202), .ZN(n4577) );
  OAI21_X1 U5729 ( .B1(n4579), .B2(n4578), .A(n4577), .ZN(n5876) );
  NAND2_X1 U5730 ( .A1(n3096), .A2(n5777), .ZN(n6158) );
  NOR3_X1 U5731 ( .A1(n4380), .A2(n4263), .A3(n6158), .ZN(n4580) );
  INV_X1 U5732 ( .A(n4592), .ZN(n5874) );
  AOI22_X1 U5733 ( .A1(n5873), .A2(n6209), .B1(n6197), .B2(n5874), .ZN(n4581)
         );
  OAI21_X1 U5734 ( .B1(n6212), .B2(n5884), .A(n4581), .ZN(n4582) );
  AOI21_X1 U5735 ( .B1(n5876), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4582), 
        .ZN(n4583) );
  OAI21_X1 U5736 ( .B1(n4597), .B2(n4584), .A(n4583), .ZN(U3044) );
  NOR2_X2 U5737 ( .A1(n4585), .A2(n5961), .ZN(n6225) );
  INV_X1 U5738 ( .A(n6225), .ZN(n4596) );
  NOR2_X2 U5739 ( .A1(n4587), .A2(n4586), .ZN(n6226) );
  INV_X1 U5740 ( .A(n6226), .ZN(n4593) );
  INV_X1 U5741 ( .A(DATAI_19_), .ZN(n4588) );
  NOR2_X1 U5742 ( .A1(n5682), .A2(n4588), .ZN(n6134) );
  INV_X1 U5743 ( .A(DATAI_27_), .ZN(n4589) );
  NOR2_X1 U5744 ( .A1(n5682), .A2(n4589), .ZN(n6227) );
  AOI22_X1 U5745 ( .A1(n6134), .A2(n4590), .B1(n5873), .B2(n6227), .ZN(n4591)
         );
  OAI21_X1 U5746 ( .B1(n4593), .B2(n4592), .A(n4591), .ZN(n4594) );
  AOI21_X1 U5747 ( .B1(n5876), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4594), 
        .ZN(n4595) );
  OAI21_X1 U5748 ( .B1(n4597), .B2(n4596), .A(n4595), .ZN(U3047) );
  AOI21_X1 U5749 ( .B1(n4600), .B2(n4599), .A(n4609), .ZN(n5546) );
  INV_X1 U5750 ( .A(n5546), .ZN(n4602) );
  AOI22_X1 U5751 ( .A1(n5562), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5558), .ZN(n4601) );
  OAI21_X1 U5752 ( .B1(n4602), .B2(n5178), .A(n4601), .ZN(U2881) );
  AND2_X1 U5753 ( .A1(n5662), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4603)
         );
  AOI211_X1 U5754 ( .C1(n5233), .C2(n5428), .A(n4604), .B(n4603), .ZN(n4606)
         );
  NAND2_X1 U5755 ( .A1(n5546), .A2(n5669), .ZN(n4605) );
  OAI211_X1 U5756 ( .C1(n4607), .C2(n5371), .A(n4606), .B(n4605), .ZN(U2976)
         );
  INV_X1 U5757 ( .A(n4608), .ZN(n4611) );
  INV_X1 U5758 ( .A(n4609), .ZN(n4610) );
  AOI21_X1 U5759 ( .B1(n4611), .B2(n4610), .A(n4623), .ZN(n4634) );
  INV_X1 U5760 ( .A(n4634), .ZN(n4625) );
  INV_X1 U5761 ( .A(n4632), .ZN(n4619) );
  AND2_X1 U5762 ( .A1(n4613), .A2(n4612), .ZN(n4614) );
  OR2_X1 U5763 ( .A1(n4614), .A2(n4644), .ZN(n5685) );
  NOR3_X2 U5764 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5507), .A3(n6203), .ZN(
        n5483) );
  AOI21_X1 U5765 ( .B1(n5519), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5483), 
        .ZN(n4616) );
  OAI21_X1 U5766 ( .B1(n5409), .B2(n5487), .A(n5486), .ZN(n5416) );
  AOI22_X1 U5767 ( .A1(EBX_REG_11__SCAN_IN), .A2(n5518), .B1(
        REIP_REG_11__SCAN_IN), .B2(n5416), .ZN(n4615) );
  OAI211_X1 U5768 ( .C1(n5449), .C2(n5685), .A(n4616), .B(n4615), .ZN(n4618)
         );
  NAND2_X1 U5769 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5455) );
  NAND4_X1 U5770 ( .A1(n5513), .A2(REIP_REG_4__SCAN_IN), .A3(
        REIP_REG_5__SCAN_IN), .A4(n5488), .ZN(n5469) );
  NOR2_X1 U5771 ( .A1(n5455), .A2(n5469), .ZN(n5444) );
  NAND2_X1 U5772 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5444), .ZN(n5439) );
  NOR3_X1 U5773 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5421), .A3(n5439), .ZN(n4617) );
  AOI211_X1 U5774 ( .C1(n5520), .C2(n4619), .A(n4618), .B(n4617), .ZN(n4620)
         );
  OAI21_X1 U5775 ( .B1(n4625), .B2(n5452), .A(n4620), .ZN(U2816) );
  INV_X1 U5776 ( .A(DATAI_11_), .ZN(n6648) );
  INV_X1 U5777 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6596) );
  OAI222_X1 U5778 ( .A1(n4625), .A2(n5178), .B1(n5008), .B2(n6648), .C1(n5566), 
        .C2(n6596), .ZN(U2880) );
  OAI21_X1 U5779 ( .B1(n4623), .B2(n4622), .A(n4621), .ZN(n4657) );
  AOI22_X1 U5780 ( .A1(n5562), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n5558), .ZN(n4624) );
  OAI21_X1 U5781 ( .B1(n4657), .B2(n5178), .A(n4624), .ZN(U2879) );
  INV_X1 U5782 ( .A(EBX_REG_11__SCAN_IN), .ZN(n4626) );
  OAI222_X1 U5783 ( .A1(n5685), .A2(n5553), .B1(n5554), .B2(n4626), .C1(n4625), 
        .C2(n5555), .ZN(U2848) );
  NAND2_X1 U5784 ( .A1(n4629), .A2(n4628), .ZN(n4630) );
  XNOR2_X1 U5785 ( .A(n4627), .B(n4630), .ZN(n5687) );
  INV_X1 U5786 ( .A(n5687), .ZN(n4636) );
  AOI22_X1 U5787 ( .A1(n5662), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n5348), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n4631) );
  OAI21_X1 U5788 ( .B1(n4632), .B2(n5673), .A(n4631), .ZN(n4633) );
  AOI21_X1 U5789 ( .B1(n4634), .B2(n5669), .A(n4633), .ZN(n4635) );
  OAI21_X1 U5790 ( .B1(n4636), .B2(n5371), .A(n4635), .ZN(U2975) );
  INV_X1 U5791 ( .A(n4638), .ZN(n4639) );
  NOR2_X1 U5792 ( .A1(n4640), .A2(n4639), .ZN(n4641) );
  XNOR2_X1 U5793 ( .A(n4637), .B(n4641), .ZN(n4660) );
  OAI21_X1 U5794 ( .B1(n4644), .B2(n4643), .A(n4642), .ZN(n4645) );
  INV_X1 U5795 ( .A(n4645), .ZN(n5541) );
  AND2_X1 U5796 ( .A1(n5348), .A2(REIP_REG_12__SCAN_IN), .ZN(n4656) );
  INV_X1 U5797 ( .A(n4666), .ZN(n4667) );
  AOI22_X1 U5798 ( .A1(n5721), .A2(n4648), .B1(n4647), .B2(n4646), .ZN(n4650)
         );
  NAND2_X1 U5799 ( .A1(n4650), .A2(n4649), .ZN(n5684) );
  AOI221_X1 U5800 ( .B1(n5721), .B2(n4667), .C1(n4651), .C2(n4667), .A(n5684), 
        .ZN(n4652) );
  AOI221_X1 U5801 ( .B1(n5690), .B2(n4065), .C1(n6579), .C2(n4065), .A(n4652), 
        .ZN(n4653) );
  AOI211_X1 U5802 ( .C1(n5754), .C2(n5541), .A(n4656), .B(n4653), .ZN(n4654)
         );
  OAI21_X1 U5803 ( .B1(n4660), .B2(n5733), .A(n4654), .ZN(U3006) );
  AND2_X1 U5804 ( .A1(n5662), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4655)
         );
  AOI211_X1 U5805 ( .C1(n5233), .C2(n5417), .A(n4656), .B(n4655), .ZN(n4659)
         );
  INV_X1 U5806 ( .A(n4657), .ZN(n5542) );
  NAND2_X1 U5807 ( .A1(n5542), .A2(n5669), .ZN(n4658) );
  OAI211_X1 U5808 ( .C1(n4660), .C2(n5371), .A(n4659), .B(n4658), .ZN(U2974)
         );
  OAI21_X1 U5809 ( .B1(n4662), .B2(n4661), .A(n4808), .ZN(n4663) );
  INV_X1 U5810 ( .A(n4663), .ZN(n4677) );
  AOI21_X1 U5811 ( .B1(n5768), .B2(n4664), .A(n5684), .ZN(n4665) );
  OAI21_X1 U5812 ( .B1(n4666), .B2(n5765), .A(n4665), .ZN(n5344) );
  NOR2_X1 U5813 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4667), .ZN(n5346)
         );
  INV_X1 U5814 ( .A(n5690), .ZN(n4668) );
  AOI22_X1 U5815 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5344), .B1(n5346), .B2(n4668), .ZN(n4670) );
  XNOR2_X1 U5816 ( .A(n4642), .B(n4825), .ZN(n5539) );
  AND2_X1 U5817 ( .A1(n5348), .A2(REIP_REG_13__SCAN_IN), .ZN(n4673) );
  AOI21_X1 U5818 ( .B1(n5754), .B2(n5539), .A(n4673), .ZN(n4669) );
  OAI211_X1 U5819 ( .C1(n4677), .C2(n5733), .A(n4670), .B(n4669), .ZN(U3005)
         );
  XOR2_X1 U5820 ( .A(n4672), .B(n4671), .Z(n5564) );
  AOI21_X1 U5821 ( .B1(n5662), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n4673), 
        .ZN(n4674) );
  OAI21_X1 U5822 ( .B1(n5407), .B2(n5673), .A(n4674), .ZN(n4675) );
  AOI21_X1 U5823 ( .B1(n5564), .B2(n5669), .A(n4675), .ZN(n4676) );
  OAI21_X1 U5824 ( .B1(n4677), .B2(n5371), .A(n4676), .ZN(U2973) );
  AOI21_X1 U5825 ( .B1(n4678), .B2(n4680), .A(n6389), .ZN(n4687) );
  NOR3_X1 U5826 ( .A1(n6431), .A2(n6679), .A3(n4679), .ZN(n4683) );
  AND3_X1 U5827 ( .A1(n4681), .A2(n4686), .A3(n4680), .ZN(n4682) );
  AOI211_X1 U5828 ( .C1(n4684), .C2(n5357), .A(n4683), .B(n4682), .ZN(n4685)
         );
  OAI22_X1 U5829 ( .A1(n4687), .A2(n4686), .B1(n6389), .B2(n4685), .ZN(U3459)
         );
  INV_X1 U5830 ( .A(n4688), .ZN(n4866) );
  OAI22_X1 U5831 ( .A1(n4866), .A2(n4689), .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n4867), .ZN(n4690) );
  XNOR2_X1 U5832 ( .A(n4690), .B(n6731), .ZN(n4803) );
  AOI211_X1 U5833 ( .C1(n4151), .C2(n4692), .A(n4693), .B(n4691), .ZN(n4698)
         );
  INV_X1 U5834 ( .A(n4151), .ZN(n4696) );
  INV_X1 U5835 ( .A(n4693), .ZN(n4695) );
  AOI211_X1 U5836 ( .C1(n4987), .C2(n4696), .A(n4695), .B(n4694), .ZN(n4697)
         );
  NOR2_X1 U5837 ( .A1(n4698), .A2(n4697), .ZN(n5083) );
  INV_X1 U5838 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6374) );
  NOR2_X1 U5839 ( .A1(n5740), .A2(n6374), .ZN(n4705) );
  NOR3_X1 U5840 ( .A1(n6515), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4883), 
        .ZN(n4699) );
  INV_X1 U5841 ( .A(n4700), .ZN(n4885) );
  OAI211_X1 U5842 ( .C1(n4885), .C2(n6515), .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5238), .ZN(n4701) );
  OAI211_X1 U5843 ( .C1(n4803), .C2(n5733), .A(n4702), .B(n4701), .ZN(U2988)
         );
  XNOR2_X1 U5844 ( .A(n4751), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5080)
         );
  NOR2_X1 U5845 ( .A1(n5676), .A2(n4703), .ZN(n4704) );
  AOI211_X1 U5846 ( .C1(n5080), .C2(n5233), .A(n4705), .B(n4704), .ZN(n4802)
         );
  OR2_X1 U5847 ( .A1(n4706), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4707)
         );
  NAND2_X1 U5848 ( .A1(n4707), .A2(n4745), .ZN(n5202) );
  AOI22_X1 U5849 ( .A1(n3081), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4711) );
  AOI22_X1 U5850 ( .A1(n4773), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4710) );
  AOI22_X1 U5851 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4772), .B1(n3772), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4709) );
  AOI22_X1 U5852 ( .A1(n4782), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4708) );
  NAND4_X1 U5853 ( .A1(n4711), .A2(n4710), .A3(n4709), .A4(n4708), .ZN(n4717)
         );
  AOI22_X1 U5854 ( .A1(n3098), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4715) );
  AOI22_X1 U5855 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4781), .B1(n3080), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4714) );
  AOI22_X1 U5856 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3797), .B1(n3082), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5857 ( .A1(n3312), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4712) );
  NAND4_X1 U5858 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4716)
         );
  NOR2_X1 U5859 ( .A1(n4717), .A2(n4716), .ZN(n4730) );
  NAND2_X1 U5860 ( .A1(n4719), .A2(n4718), .ZN(n4729) );
  XNOR2_X1 U5861 ( .A(n4730), .B(n4729), .ZN(n4720) );
  NOR2_X1 U5862 ( .A1(n4720), .A2(n4767), .ZN(n4725) );
  INV_X1 U5863 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4722) );
  NAND2_X1 U5864 ( .A1(n6550), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4721)
         );
  OAI211_X1 U5865 ( .C1(n4723), .C2(n4722), .A(n4795), .B(n4721), .ZN(n4724)
         );
  OAI22_X1 U5866 ( .A1(n5202), .A2(n4795), .B1(n4725), .B2(n4724), .ZN(n4971)
         );
  INV_X1 U5867 ( .A(n4726), .ZN(n4727) );
  NOR2_X1 U5868 ( .A1(n4971), .A2(n4727), .ZN(n4728) );
  NAND2_X1 U5869 ( .A1(n5135), .A2(n4728), .ZN(n4963) );
  NOR2_X1 U5870 ( .A1(n4730), .A2(n4729), .ZN(n4764) );
  AOI22_X1 U5871 ( .A1(n4773), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4774), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5872 ( .A1(n3081), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5873 ( .A1(n3080), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U5874 ( .A1(n3097), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4731) );
  NAND4_X1 U5875 ( .A1(n4734), .A2(n4733), .A3(n4732), .A4(n4731), .ZN(n4740)
         );
  AOI22_X1 U5876 ( .A1(n3312), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4738) );
  AOI22_X1 U5877 ( .A1(n4782), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4737) );
  AOI22_X1 U5878 ( .A1(n3797), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4736) );
  AOI22_X1 U5879 ( .A1(n3082), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4735) );
  NAND4_X1 U5880 ( .A1(n4738), .A2(n4737), .A3(n4736), .A4(n4735), .ZN(n4739)
         );
  OR2_X1 U5881 ( .A1(n4740), .A2(n4739), .ZN(n4763) );
  INV_X1 U5882 ( .A(n4763), .ZN(n4741) );
  XNOR2_X1 U5883 ( .A(n4764), .B(n4741), .ZN(n4742) );
  INV_X1 U5884 ( .A(n4767), .ZN(n4792) );
  NAND2_X1 U5885 ( .A1(n4742), .A2(n4792), .ZN(n4749) );
  NAND2_X1 U5886 ( .A1(n6550), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4743)
         );
  NAND2_X1 U5887 ( .A1(n4795), .A2(n4743), .ZN(n4744) );
  AOI21_X1 U5888 ( .B1(n4797), .B2(EAX_REG_28__SCAN_IN), .A(n4744), .ZN(n4748)
         );
  XNOR2_X1 U5889 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .B(n4745), .ZN(n5097)
         );
  AND2_X1 U5890 ( .A1(n5097), .A2(n3079), .ZN(n4747) );
  AOI21_X1 U5891 ( .B1(n4749), .B2(n4748), .A(n4747), .ZN(n4964) );
  INV_X1 U5892 ( .A(n4964), .ZN(n4750) );
  NAND2_X1 U5893 ( .A1(n5136), .A2(n3105), .ZN(n4966) );
  OAI21_X1 U5894 ( .B1(n4752), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4751), 
        .ZN(n5088) );
  AOI22_X1 U5895 ( .A1(n3081), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4773), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4756) );
  AOI22_X1 U5896 ( .A1(n3312), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4755) );
  AOI22_X1 U5897 ( .A1(n3797), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4782), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4754) );
  AOI22_X1 U5898 ( .A1(n3082), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4753) );
  NAND4_X1 U5899 ( .A1(n4756), .A2(n4755), .A3(n4754), .A4(n4753), .ZN(n4762)
         );
  AOI22_X1 U5900 ( .A1(n4774), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4760) );
  AOI22_X1 U5901 ( .A1(n3080), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4759) );
  AOI22_X1 U5902 ( .A1(n3098), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4758) );
  AOI22_X1 U5903 ( .A1(n4775), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4757) );
  NAND4_X1 U5904 ( .A1(n4760), .A2(n4759), .A3(n4758), .A4(n4757), .ZN(n4761)
         );
  NOR2_X1 U5905 ( .A1(n4762), .A2(n4761), .ZN(n4771) );
  NAND2_X1 U5906 ( .A1(n4764), .A2(n4763), .ZN(n4770) );
  XNOR2_X1 U5907 ( .A(n4771), .B(n4770), .ZN(n4768) );
  AOI21_X1 U5908 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6550), .A(n3079), 
        .ZN(n4766) );
  NAND2_X1 U5909 ( .A1(n3349), .A2(EAX_REG_29__SCAN_IN), .ZN(n4765) );
  OAI211_X1 U5910 ( .C1(n4768), .C2(n4767), .A(n4766), .B(n4765), .ZN(n4769)
         );
  OAI21_X1 U5911 ( .B1(n4795), .B2(n5088), .A(n4769), .ZN(n4870) );
  NOR2_X1 U5912 ( .A1(n4771), .A2(n4770), .ZN(n4791) );
  AOI22_X1 U5913 ( .A1(n3289), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4772), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4779) );
  AOI22_X1 U5914 ( .A1(n3081), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4773), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4778) );
  AOI22_X1 U5915 ( .A1(n4774), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4777) );
  AOI22_X1 U5916 ( .A1(n3797), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4775), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4776) );
  NAND4_X1 U5917 ( .A1(n4779), .A2(n4778), .A3(n4777), .A4(n4776), .ZN(n4789)
         );
  AOI22_X1 U5918 ( .A1(n3447), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4780), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4787) );
  AOI22_X1 U5919 ( .A1(n3080), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4781), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4786) );
  AOI22_X1 U5920 ( .A1(n4782), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5921 ( .A1(n3082), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4783), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4784) );
  NAND4_X1 U5922 ( .A1(n4787), .A2(n4786), .A3(n4785), .A4(n4784), .ZN(n4788)
         );
  NOR2_X1 U5923 ( .A1(n4789), .A2(n4788), .ZN(n4790) );
  XNOR2_X1 U5924 ( .A(n4791), .B(n4790), .ZN(n4793) );
  NAND2_X1 U5925 ( .A1(n4793), .A2(n4792), .ZN(n4800) );
  NAND2_X1 U5926 ( .A1(n6550), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4794)
         );
  NAND2_X1 U5927 ( .A1(n4795), .A2(n4794), .ZN(n4796) );
  AOI21_X1 U5928 ( .B1(n4797), .B2(EAX_REG_30__SCAN_IN), .A(n4796), .ZN(n4799)
         );
  AND2_X1 U5929 ( .A1(n5080), .A2(n3079), .ZN(n4798) );
  AOI21_X1 U5930 ( .B1(n4800), .B2(n4799), .A(n4798), .ZN(n4888) );
  XNOR2_X1 U5931 ( .A(n4889), .B(n4888), .ZN(n4915) );
  INV_X1 U5932 ( .A(n4915), .ZN(n5170) );
  NAND2_X1 U5933 ( .A1(n5170), .A2(n5669), .ZN(n4801) );
  OAI211_X1 U5934 ( .C1(n4803), .C2(n5371), .A(n4802), .B(n4801), .ZN(U2956)
         );
  INV_X1 U5935 ( .A(n5232), .ZN(n4806) );
  INV_X1 U5936 ( .A(n4804), .ZN(n4805) );
  OAI21_X1 U5937 ( .B1(n4806), .B2(n4805), .A(n5157), .ZN(n5000) );
  NOR2_X1 U5938 ( .A1(n5227), .A2(n4812), .ZN(n4813) );
  NOR2_X1 U5939 ( .A1(n4814), .A2(n5321), .ZN(n4815) );
  OAI21_X1 U5940 ( .B1(n5676), .B2(n3656), .A(n4819), .ZN(n4820) );
  OAI21_X1 U5941 ( .B1(n5000), .B2(n5682), .A(n4821), .ZN(U2968) );
  NAND2_X1 U5942 ( .A1(n4947), .A2(n4946), .ZN(n5006) );
  OAI21_X1 U5943 ( .B1(n4947), .B2(n4946), .A(n5006), .ZN(n5057) );
  AOI22_X1 U5944 ( .A1(n5562), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5558), .ZN(n4823) );
  OAI21_X1 U5945 ( .B1(n5057), .B2(n5178), .A(n4823), .ZN(U2877) );
  INV_X1 U5946 ( .A(n4642), .ZN(n4826) );
  AOI21_X1 U5947 ( .B1(n4826), .B2(n4825), .A(n4824), .ZN(n4828) );
  INV_X1 U5948 ( .A(n4827), .ZN(n5335) );
  NOR2_X1 U5949 ( .A1(n4828), .A2(n5335), .ZN(n5349) );
  AOI22_X1 U5950 ( .A1(n5349), .A2(n5549), .B1(EBX_REG_14__SCAN_IN), .B2(n5535), .ZN(n4829) );
  OAI21_X1 U5951 ( .B1(n5057), .B2(n5555), .A(n4829), .ZN(U2845) );
  AOI21_X1 U5952 ( .B1(n5519), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5483), 
        .ZN(n4830) );
  OAI21_X1 U5953 ( .B1(n5512), .B2(n5059), .A(n4830), .ZN(n4837) );
  AOI21_X1 U5954 ( .B1(n5513), .B2(n4831), .A(REIP_REG_14__SCAN_IN), .ZN(n4835) );
  NOR2_X1 U5955 ( .A1(n5424), .A2(n4832), .ZN(n5398) );
  INV_X1 U5956 ( .A(n5398), .ZN(n4834) );
  INV_X1 U5957 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4833) );
  OAI22_X1 U5958 ( .A1(n4835), .A2(n4834), .B1(n4833), .B2(n5505), .ZN(n4836)
         );
  AOI211_X1 U5959 ( .C1(n5349), .C2(n5517), .A(n4837), .B(n4836), .ZN(n4838)
         );
  OAI21_X1 U5960 ( .B1(n5057), .B2(n5452), .A(n4838), .ZN(U2813) );
  AOI21_X1 U5961 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5054), .A(n4839), 
        .ZN(n4840) );
  NAND2_X1 U5962 ( .A1(n5138), .A2(n4841), .ZN(n4842) );
  INV_X1 U5963 ( .A(n5122), .ZN(n4845) );
  AOI22_X1 U5964 ( .A1(n5662), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .B1(n5348), 
        .B2(REIP_REG_22__SCAN_IN), .ZN(n4844) );
  OAI21_X1 U5965 ( .B1(n4845), .B2(n5673), .A(n4844), .ZN(n4846) );
  AOI21_X1 U5966 ( .B1(n5189), .B2(n5669), .A(n4846), .ZN(n4847) );
  OAI21_X1 U5967 ( .B1(n4848), .B2(n5371), .A(n4847), .ZN(U2964) );
  INV_X1 U5968 ( .A(n5556), .ZN(n5177) );
  NAND2_X1 U5969 ( .A1(EAX_REG_24__SCAN_IN), .A2(n5558), .ZN(n4849) );
  OAI21_X1 U5970 ( .B1(n5177), .B2(n4850), .A(n4849), .ZN(n4851) );
  AOI21_X1 U5971 ( .B1(n5559), .B2(DATAI_8_), .A(n4851), .ZN(n4852) );
  OAI21_X1 U5972 ( .B1(n5025), .B2(n5178), .A(n4852), .ZN(U2867) );
  INV_X1 U5973 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4853) );
  OAI222_X1 U5974 ( .A1(n5555), .A2(n5025), .B1(n5554), .B2(n4853), .C1(n5067), 
        .C2(n5553), .ZN(U2835) );
  OAI22_X1 U5975 ( .A1(n5258), .A2(n5553), .B1(n4855), .B2(n5554), .ZN(n4856)
         );
  INV_X1 U5976 ( .A(n4856), .ZN(n4857) );
  OAI21_X1 U5977 ( .B1(n4854), .B2(n5555), .A(n4857), .ZN(U2833) );
  AOI22_X1 U5978 ( .A1(n5559), .A2(DATAI_10_), .B1(n5558), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n4859) );
  NAND2_X1 U5979 ( .A1(n5556), .A2(DATAI_26_), .ZN(n4858) );
  OAI211_X1 U5980 ( .C1(n4854), .C2(n5178), .A(n4859), .B(n4858), .ZN(U2865)
         );
  NAND2_X1 U5981 ( .A1(n5010), .A2(n4860), .ZN(n4861) );
  XNOR2_X1 U5982 ( .A(n4867), .B(n4861), .ZN(n5255) );
  NAND2_X1 U5983 ( .A1(n5255), .A2(n5679), .ZN(n4865) );
  OAI22_X1 U5984 ( .A1(n5676), .A2(n3873), .B1(n5740), .B2(n6639), .ZN(n4862)
         );
  AOI21_X1 U5985 ( .B1(n5233), .B2(n4863), .A(n4862), .ZN(n4864) );
  OAI211_X1 U5986 ( .C1(n5682), .C2(n4854), .A(n4865), .B(n4864), .ZN(U2960)
         );
  NOR2_X1 U5987 ( .A1(n5010), .A2(n5239), .ZN(n4868) );
  AOI21_X1 U5988 ( .B1(n4868), .B2(n4867), .A(n4866), .ZN(n4869) );
  XNOR2_X1 U5989 ( .A(n4869), .B(n6515), .ZN(n4887) );
  AOI21_X1 U5990 ( .B1(n4870), .B2(n4966), .A(n4889), .ZN(n5173) );
  NAND2_X1 U5991 ( .A1(n5348), .A2(REIP_REG_29__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U5992 ( .A1(n5662), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4871)
         );
  OAI211_X1 U5993 ( .C1(n5673), .C2(n5088), .A(n4881), .B(n4871), .ZN(n4872)
         );
  AOI21_X1 U5994 ( .B1(n5173), .B2(n5669), .A(n4872), .ZN(n4873) );
  OAI21_X1 U5995 ( .B1(n4887), .B2(n5371), .A(n4873), .ZN(U2957) );
  NAND2_X1 U5996 ( .A1(n4874), .A2(n3093), .ZN(n4877) );
  INV_X1 U5997 ( .A(n4875), .ZN(n4876) );
  NAND2_X1 U5998 ( .A1(n4877), .A2(n4876), .ZN(n4878) );
  NOR2_X1 U5999 ( .A1(n4151), .A2(n4878), .ZN(n4879) );
  NOR2_X1 U6000 ( .A1(n4880), .A2(n4879), .ZN(n5091) );
  NAND2_X1 U6001 ( .A1(n5091), .A2(n5754), .ZN(n4882) );
  OAI211_X1 U6002 ( .C1(INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n4883), .A(n4882), .B(n4881), .ZN(n4884) );
  AOI21_X1 U6003 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n4885), .A(n4884), 
        .ZN(n4886) );
  OAI21_X1 U6004 ( .B1(n4887), .B2(n5733), .A(n4886), .ZN(U2989) );
  NAND2_X1 U6005 ( .A1(n4889), .A2(n4888), .ZN(n4893) );
  AOI22_X1 U6006 ( .A1(n3349), .A2(EAX_REG_31__SCAN_IN), .B1(n4890), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4891) );
  INV_X1 U6007 ( .A(n4891), .ZN(n4892) );
  INV_X1 U6008 ( .A(n4917), .ZN(n4906) );
  INV_X1 U6009 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4897) );
  NAND3_X1 U6010 ( .A1(n4895), .A2(EBX_REG_31__SCAN_IN), .A3(n4894), .ZN(n4896) );
  OAI21_X1 U6011 ( .B1(n5499), .B2(n4897), .A(n4896), .ZN(n4901) );
  NOR2_X1 U6012 ( .A1(n4899), .A2(n4898), .ZN(n5106) );
  NAND3_X1 U6013 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5106), .ZN(n5094) );
  INV_X1 U6014 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U6015 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4902) );
  AOI21_X1 U6016 ( .B1(n5513), .B2(n4902), .A(n5105), .ZN(n5095) );
  OAI21_X1 U6017 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5487), .A(n5095), .ZN(n5081) );
  NOR2_X1 U6018 ( .A1(n5487), .A2(REIP_REG_30__SCAN_IN), .ZN(n4903) );
  OAI21_X1 U6019 ( .B1(n5081), .B2(n4903), .A(REIP_REG_31__SCAN_IN), .ZN(n4904) );
  OAI211_X1 U6020 ( .C1(n4906), .C2(n5452), .A(n4905), .B(n4904), .ZN(U2796)
         );
  AOI21_X1 U6021 ( .B1(n5662), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4907), 
        .ZN(n4908) );
  OAI21_X1 U6022 ( .B1(n5673), .B2(n4909), .A(n4908), .ZN(n4910) );
  AOI21_X1 U6023 ( .B1(n4917), .B2(n5669), .A(n4910), .ZN(n4911) );
  OAI21_X1 U6024 ( .B1(n4912), .B2(n5371), .A(n4911), .ZN(U2955) );
  INV_X1 U6025 ( .A(n5083), .ZN(n4913) );
  OAI222_X1 U6026 ( .A1(n5555), .A2(n4915), .B1(n4914), .B2(n5554), .C1(n4913), 
        .C2(n5553), .ZN(U2829) );
  NAND3_X1 U6027 ( .A1(n4917), .A2(n4916), .A3(n5566), .ZN(n4919) );
  AOI22_X1 U6028 ( .A1(n5556), .A2(DATAI_31_), .B1(n5558), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U6029 ( .A1(n4919), .A2(n4918), .ZN(U2860) );
  OR2_X1 U6030 ( .A1(n4921), .A2(n4920), .ZN(n4923) );
  OAI22_X1 U6031 ( .A1(REIP_REG_25__SCAN_IN), .A2(n4924), .B1(n5210), .B2(
        n5512), .ZN(n4933) );
  OR2_X1 U6032 ( .A1(n4208), .A2(n4925), .ZN(n4927) );
  AND2_X1 U6033 ( .A1(n4927), .A2(n4926), .ZN(n5259) );
  INV_X1 U6034 ( .A(n5259), .ZN(n4931) );
  OAI21_X1 U6035 ( .B1(n4928), .B2(n5117), .A(REIP_REG_25__SCAN_IN), .ZN(n4930) );
  AOI22_X1 U6036 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5518), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5519), .ZN(n4929) );
  OAI211_X1 U6037 ( .C1(n5449), .C2(n4931), .A(n4930), .B(n4929), .ZN(n4932)
         );
  AOI211_X1 U6038 ( .C1(n5207), .C2(n5465), .A(n4933), .B(n4932), .ZN(n4934)
         );
  INV_X1 U6039 ( .A(n4934), .ZN(U2802) );
  MUX2_X1 U6040 ( .A(EBX_REG_18__SCAN_IN), .B(n4937), .S(n3094), .Z(n4938) );
  INV_X1 U6041 ( .A(n4938), .ZN(n5149) );
  XNOR2_X1 U6042 ( .A(n4935), .B(n5149), .ZN(n5308) );
  INV_X1 U6043 ( .A(n4939), .ZN(n4941) );
  AOI21_X1 U6044 ( .B1(n5519), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5483), 
        .ZN(n4940) );
  OAI21_X1 U6045 ( .B1(n5512), .B2(n4941), .A(n4940), .ZN(n4944) );
  AOI22_X1 U6046 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5518), .B1(n5161), .B2(n6487), .ZN(n4942) );
  OAI21_X1 U6047 ( .B1(n6487), .B2(n5387), .A(n4942), .ZN(n4943) );
  AOI211_X1 U6048 ( .C1(n5308), .C2(n5517), .A(n4944), .B(n4943), .ZN(n4945)
         );
  OAI21_X1 U6049 ( .B1(n5000), .B2(n5452), .A(n4945), .ZN(U2809) );
  AND2_X1 U6050 ( .A1(n4947), .A2(n4946), .ZN(n4949) );
  AOI21_X1 U6051 ( .B1(n4950), .B2(n5004), .A(n5230), .ZN(n5042) );
  INV_X1 U6052 ( .A(n5042), .ZN(n5003) );
  NOR2_X1 U6053 ( .A1(n5332), .A2(n4951), .ZN(n4952) );
  OR2_X1 U6054 ( .A1(n5314), .A2(n4952), .ZN(n4995) );
  INV_X1 U6055 ( .A(n4995), .ZN(n5327) );
  INV_X1 U6056 ( .A(n5483), .ZN(n5472) );
  NAND2_X1 U6057 ( .A1(n5519), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4953)
         );
  OAI211_X1 U6058 ( .C1(n5512), .C2(n5040), .A(n5472), .B(n4953), .ZN(n4958)
         );
  INV_X1 U6059 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6593) );
  AND2_X1 U6060 ( .A1(n6593), .A2(n4954), .ZN(n5397) );
  OAI21_X1 U6061 ( .B1(n5398), .B2(n5397), .A(REIP_REG_16__SCAN_IN), .ZN(n4956) );
  INV_X1 U6062 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6352) );
  NAND3_X1 U6063 ( .A1(REIP_REG_15__SCAN_IN), .A2(n4954), .A3(n6352), .ZN(
        n4955) );
  OAI211_X1 U6064 ( .C1(n5505), .C2(n3934), .A(n4956), .B(n4955), .ZN(n4957)
         );
  AOI211_X1 U6065 ( .C1(n5327), .C2(n5517), .A(n4958), .B(n4957), .ZN(n4959)
         );
  OAI21_X1 U6066 ( .B1(n5003), .B2(n5452), .A(n4959), .ZN(U2811) );
  INV_X1 U6067 ( .A(n5173), .ZN(n4962) );
  INV_X1 U6068 ( .A(n5091), .ZN(n4960) );
  OAI222_X1 U6069 ( .A1(n5555), .A2(n4962), .B1(n4961), .B2(n5554), .C1(n4960), 
        .C2(n5553), .ZN(U2830) );
  INV_X1 U6070 ( .A(n5136), .ZN(n4991) );
  NOR2_X1 U6071 ( .A1(n4991), .A2(n4963), .ZN(n4973) );
  OR2_X1 U6072 ( .A1(n4973), .A2(n4964), .ZN(n4965) );
  NAND2_X1 U6073 ( .A1(n4966), .A2(n4965), .ZN(n5179) );
  NOR2_X1 U6074 ( .A1(n4977), .A2(n4967), .ZN(n4968) );
  OR2_X1 U6075 ( .A1(n4151), .A2(n4968), .ZN(n5246) );
  OAI22_X1 U6076 ( .A1(n5246), .A2(n5553), .B1(n6528), .B2(n5554), .ZN(n4969)
         );
  INV_X1 U6077 ( .A(n4969), .ZN(n4970) );
  OAI21_X1 U6078 ( .B1(n5179), .B2(n5555), .A(n4970), .ZN(U2831) );
  AND2_X1 U6079 ( .A1(n4972), .A2(n4971), .ZN(n4974) );
  AND2_X1 U6080 ( .A1(n3099), .A2(n4975), .ZN(n4976) );
  NOR2_X1 U6081 ( .A1(n4977), .A2(n4976), .ZN(n5249) );
  AOI22_X1 U6082 ( .A1(n5249), .A2(n5549), .B1(EBX_REG_27__SCAN_IN), .B2(n5535), .ZN(n4978) );
  OAI21_X1 U6083 ( .B1(n5107), .B2(n5555), .A(n4978), .ZN(U2832) );
  INV_X1 U6084 ( .A(n5207), .ZN(n4980) );
  AOI22_X1 U6085 ( .A1(n5259), .A2(n5549), .B1(EBX_REG_25__SCAN_IN), .B2(n5535), .ZN(n4979) );
  OAI21_X1 U6086 ( .B1(n4980), .B2(n5555), .A(n4979), .ZN(U2834) );
  INV_X1 U6087 ( .A(n5189), .ZN(n4986) );
  INV_X1 U6088 ( .A(EBX_REG_22__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U6089 ( .A1(n4983), .A2(n4982), .ZN(n4984) );
  NAND2_X1 U6090 ( .A1(n5114), .A2(n4984), .ZN(n5276) );
  OAI222_X1 U6091 ( .A1(n5555), .A2(n4986), .B1(n5554), .B2(n4985), .C1(n5276), 
        .C2(n5553), .ZN(U2837) );
  MUX2_X1 U6092 ( .A(n4988), .B(n4987), .S(n5152), .Z(n4990) );
  XNOR2_X1 U6093 ( .A(n4990), .B(n4989), .ZN(n5295) );
  INV_X1 U6094 ( .A(n5295), .ZN(n5142) );
  OAI21_X1 U6095 ( .B1(n4992), .B2(n5158), .A(n4991), .ZN(n5143) );
  OAI222_X1 U6096 ( .A1(n5553), .A2(n5142), .B1(n3944), .B2(n5554), .C1(n5555), 
        .C2(n5143), .ZN(U2839) );
  INV_X1 U6097 ( .A(n5308), .ZN(n4993) );
  OAI222_X1 U6098 ( .A1(n5000), .A2(n5555), .B1(n4994), .B2(n5554), .C1(n5553), 
        .C2(n4993), .ZN(U2841) );
  OAI222_X1 U6099 ( .A1(n5003), .A2(n5555), .B1(n5554), .B2(n3934), .C1(n4995), 
        .C2(n5553), .ZN(U2843) );
  AOI22_X1 U6100 ( .A1(n5559), .A2(DATAI_4_), .B1(n5558), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U6101 ( .A1(n5556), .A2(DATAI_20_), .ZN(n4996) );
  OAI211_X1 U6102 ( .C1(n5143), .C2(n5178), .A(n4997), .B(n4996), .ZN(U2871)
         );
  AOI22_X1 U6103 ( .A1(n5556), .A2(DATAI_18_), .B1(n5558), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n4999) );
  NAND2_X1 U6104 ( .A1(n5559), .A2(DATAI_2_), .ZN(n4998) );
  OAI211_X1 U6105 ( .C1(n5000), .C2(n5178), .A(n4999), .B(n4998), .ZN(U2873)
         );
  AOI22_X1 U6106 ( .A1(n5556), .A2(DATAI_16_), .B1(n5558), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5002) );
  NAND2_X1 U6107 ( .A1(n5559), .A2(DATAI_0_), .ZN(n5001) );
  OAI211_X1 U6108 ( .C1(n5003), .C2(n5178), .A(n5002), .B(n5001), .ZN(U2875)
         );
  INV_X1 U6109 ( .A(n5004), .ZN(n5005) );
  AOI21_X1 U6110 ( .B1(n5007), .B2(n5006), .A(n5005), .ZN(n5536) );
  INV_X1 U6111 ( .A(n5536), .ZN(n5009) );
  INV_X1 U6112 ( .A(DATAI_15_), .ZN(n6527) );
  INV_X1 U6113 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6729) );
  OAI222_X1 U6114 ( .A1(n5009), .A2(n5178), .B1(n6527), .B2(n5008), .C1(n5566), 
        .C2(n6729), .ZN(U2876) );
  NOR2_X1 U6115 ( .A1(n5203), .A2(n5010), .ZN(n5196) );
  NAND2_X1 U6116 ( .A1(n5243), .A2(n5679), .ZN(n5020) );
  INV_X1 U6117 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5017) );
  INV_X1 U6118 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5016) );
  OAI22_X1 U6119 ( .A1(n5676), .A2(n5017), .B1(n5740), .B2(n5016), .ZN(n5018)
         );
  AOI21_X1 U6120 ( .B1(n5233), .B2(n5097), .A(n5018), .ZN(n5019) );
  OAI211_X1 U6121 ( .C1(n5682), .C2(n5179), .A(n5020), .B(n5019), .ZN(U2958)
         );
  NAND4_X1 U6122 ( .A1(n5021), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .A4(n5224), .ZN(n5022) );
  OAI21_X1 U6123 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5023), .A(n5022), 
        .ZN(n5024) );
  XNOR2_X1 U6124 ( .A(n5024), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5071)
         );
  INV_X1 U6125 ( .A(n5025), .ZN(n5029) );
  NAND2_X1 U6126 ( .A1(n5348), .A2(REIP_REG_24__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6127 ( .A1(n5662), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5026)
         );
  OAI211_X1 U6128 ( .C1(n5673), .C2(n5027), .A(n5066), .B(n5026), .ZN(n5028)
         );
  AOI21_X1 U6129 ( .B1(n5029), .B2(n5669), .A(n5028), .ZN(n5030) );
  OAI21_X1 U6130 ( .B1(n5071), .B2(n5371), .A(n5030), .ZN(U2962) );
  NAND2_X1 U6131 ( .A1(n5032), .A2(n5031), .ZN(n5034) );
  XNOR2_X1 U6132 ( .A(n5054), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5033)
         );
  XNOR2_X1 U6133 ( .A(n5034), .B(n5033), .ZN(n5296) );
  NAND2_X1 U6134 ( .A1(n5296), .A2(n5679), .ZN(n5037) );
  OAI22_X1 U6135 ( .A1(n5676), .A2(n6633), .B1(n5740), .B2(n6357), .ZN(n5035)
         );
  AOI21_X1 U6136 ( .B1(n5233), .B2(n5141), .A(n5035), .ZN(n5036) );
  OAI211_X1 U6137 ( .C1(n5682), .C2(n5143), .A(n5037), .B(n5036), .ZN(U2966)
         );
  XNOR2_X1 U6138 ( .A(n5054), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5038)
         );
  XNOR2_X1 U6139 ( .A(n5227), .B(n5038), .ZN(n5326) );
  AOI22_X1 U6140 ( .A1(n5662), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n5348), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5039) );
  OAI21_X1 U6141 ( .B1(n5040), .B2(n5673), .A(n5039), .ZN(n5041) );
  AOI21_X1 U6142 ( .B1(n5042), .B2(n5669), .A(n5041), .ZN(n5043) );
  OAI21_X1 U6143 ( .B1(n5326), .B2(n5371), .A(n5043), .ZN(U2970) );
  NAND2_X1 U6144 ( .A1(n5056), .A2(n5044), .ZN(n5046) );
  NAND2_X1 U6145 ( .A1(n5046), .A2(n5045), .ZN(n5049) );
  NAND2_X1 U6146 ( .A1(n3106), .A2(n5047), .ZN(n5048) );
  XNOR2_X1 U6147 ( .A(n5049), .B(n5048), .ZN(n5338) );
  INV_X1 U6148 ( .A(n5402), .ZN(n5051) );
  AOI22_X1 U6149 ( .A1(n5662), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n5348), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5050) );
  OAI21_X1 U6150 ( .B1(n5051), .B2(n5673), .A(n5050), .ZN(n5052) );
  AOI21_X1 U6151 ( .B1(n5536), .B2(n5669), .A(n5052), .ZN(n5053) );
  OAI21_X1 U6152 ( .B1(n5338), .B2(n5371), .A(n5053), .ZN(U2971) );
  XNOR2_X1 U6153 ( .A(n5054), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5055)
         );
  XNOR2_X1 U6154 ( .A(n5056), .B(n5055), .ZN(n5351) );
  INV_X1 U6155 ( .A(n5351), .ZN(n5063) );
  INV_X1 U6156 ( .A(n5057), .ZN(n5061) );
  AOI22_X1 U6157 ( .A1(n5662), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n5348), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5058) );
  OAI21_X1 U6158 ( .B1(n5059), .B2(n5673), .A(n5058), .ZN(n5060) );
  AOI21_X1 U6159 ( .B1(n5061), .B2(n5669), .A(n5060), .ZN(n5062) );
  OAI21_X1 U6160 ( .B1(n5063), .B2(n5371), .A(n5062), .ZN(U2972) );
  OAI21_X1 U6161 ( .B1(n5272), .B2(n5065), .A(n5064), .ZN(n5069) );
  OAI21_X1 U6162 ( .B1(n5067), .B2(n5771), .A(n5066), .ZN(n5068) );
  AOI21_X1 U6163 ( .B1(n5262), .B2(n5069), .A(n5068), .ZN(n5070) );
  OAI21_X1 U6164 ( .B1(n5071), .B2(n5733), .A(n5070), .ZN(U2994) );
  OAI211_X1 U6165 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3096), .A(n6398), .B(
        n6432), .ZN(n5072) );
  OAI21_X1 U6166 ( .B1(n4239), .B2(n6399), .A(n5072), .ZN(n5073) );
  MUX2_X1 U6167 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5073), .S(n6403), 
        .Z(U3464) );
  NOR2_X1 U6168 ( .A1(n5074), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5593) );
  AOI21_X1 U6169 ( .B1(n5075), .B2(n6296), .A(n6321), .ZN(n5076) );
  NOR2_X4 U6170 ( .A1(n6421), .A2(n5583), .ZN(n5597) );
  AND2_X1 U6171 ( .A1(n5597), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6172 ( .A(n6435), .ZN(n5079) );
  INV_X1 U6173 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n5078) );
  AOI21_X1 U6174 ( .B1(n6432), .B2(n6431), .A(n6430), .ZN(n5077) );
  OAI21_X1 U6175 ( .B1(n5079), .B2(n5078), .A(n5077), .ZN(U2788) );
  AOI22_X1 U6176 ( .A1(EBX_REG_30__SCAN_IN), .A2(n5518), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n5519), .ZN(n5087) );
  AOI22_X1 U6177 ( .A1(REIP_REG_30__SCAN_IN), .A2(n5081), .B1(n5080), .B2(
        n5520), .ZN(n5086) );
  NOR3_X1 U6178 ( .A1(n5094), .A2(REIP_REG_30__SCAN_IN), .A3(n6370), .ZN(n5082) );
  AOI21_X1 U6179 ( .B1(n5170), .B2(n5465), .A(n5082), .ZN(n5085) );
  NAND2_X1 U6180 ( .A1(n5083), .A2(n5517), .ZN(n5084) );
  NAND4_X1 U6181 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(U2797)
         );
  NOR2_X1 U6182 ( .A1(n5088), .A2(n5512), .ZN(n5090) );
  INV_X1 U6183 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6703) );
  OAI22_X1 U6184 ( .A1(n5095), .A2(n6370), .B1(n6703), .B2(n5499), .ZN(n5089)
         );
  AOI211_X1 U6185 ( .C1(n5518), .C2(EBX_REG_29__SCAN_IN), .A(n5090), .B(n5089), 
        .ZN(n5093) );
  AOI22_X1 U6186 ( .A1(n5173), .A2(n5465), .B1(n5091), .B2(n5517), .ZN(n5092)
         );
  OAI211_X1 U6187 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5094), .A(n5093), .B(n5092), .ZN(U2798) );
  AOI22_X1 U6188 ( .A1(EBX_REG_28__SCAN_IN), .A2(n5518), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5519), .ZN(n5102) );
  INV_X1 U6189 ( .A(n5095), .ZN(n5096) );
  AOI22_X1 U6190 ( .A1(n5097), .A2(n5520), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5096), .ZN(n5101) );
  OAI22_X1 U6191 ( .A1(n5179), .A2(n5452), .B1(n5449), .B2(n5246), .ZN(n5098)
         );
  INV_X1 U6192 ( .A(n5098), .ZN(n5100) );
  NAND3_X1 U6193 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5106), .A3(n5016), .ZN(
        n5099) );
  NAND4_X1 U6194 ( .A1(n5102), .A2(n5101), .A3(n5100), .A4(n5099), .ZN(U2799)
         );
  INV_X1 U6195 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6367) );
  AOI22_X1 U6196 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5518), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5519), .ZN(n5103) );
  OAI21_X1 U6197 ( .B1(n5202), .B2(n5512), .A(n5103), .ZN(n5104) );
  AOI221_X1 U6198 ( .B1(n5106), .B2(n6367), .C1(n5105), .C2(
        REIP_REG_27__SCAN_IN), .A(n5104), .ZN(n5109) );
  AOI22_X1 U6199 ( .A1(n5199), .A2(n5465), .B1(n5517), .B2(n5249), .ZN(n5108)
         );
  NAND2_X1 U6200 ( .A1(n5109), .A2(n5108), .ZN(U2800) );
  INV_X1 U6201 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5111) );
  OAI22_X1 U6202 ( .A1(n5111), .A2(n5499), .B1(n5110), .B2(n5512), .ZN(n5112)
         );
  AOI21_X1 U6203 ( .B1(EBX_REG_23__SCAN_IN), .B2(n5518), .A(n5112), .ZN(n5121)
         );
  NAND2_X1 U6204 ( .A1(n5114), .A2(n5113), .ZN(n5115) );
  AND2_X1 U6205 ( .A1(n5116), .A2(n5115), .ZN(n5267) );
  AOI22_X1 U6206 ( .A1(n3104), .A2(n5465), .B1(n5517), .B2(n5267), .ZN(n5120)
         );
  OAI21_X1 U6207 ( .B1(REIP_REG_23__SCAN_IN), .B2(n5118), .A(n5117), .ZN(n5119) );
  NAND3_X1 U6208 ( .A1(n5121), .A2(n5120), .A3(n5119), .ZN(U2804) );
  AOI22_X1 U6209 ( .A1(EBX_REG_22__SCAN_IN), .A2(n5518), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5519), .ZN(n5129) );
  AOI22_X1 U6210 ( .A1(n5122), .A2(n5520), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5146), .ZN(n5128) );
  NOR2_X1 U6211 ( .A1(n5276), .A2(n5449), .ZN(n5123) );
  AOI21_X1 U6212 ( .B1(n5189), .B2(n5465), .A(n5123), .ZN(n5127) );
  INV_X1 U6213 ( .A(n5124), .ZN(n5134) );
  OAI211_X1 U6214 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5134), .B(n5125), .ZN(n5126) );
  NAND4_X1 U6215 ( .A1(n5129), .A2(n5128), .A3(n5127), .A4(n5126), .ZN(U2805)
         );
  XNOR2_X1 U6216 ( .A(n5131), .B(n5130), .ZN(n5282) );
  INV_X1 U6217 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6359) );
  AOI22_X1 U6218 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5518), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5519), .ZN(n5132) );
  OAI21_X1 U6219 ( .B1(n5214), .B2(n5512), .A(n5132), .ZN(n5133) );
  AOI221_X1 U6220 ( .B1(n5134), .B2(n6359), .C1(n5146), .C2(
        REIP_REG_21__SCAN_IN), .A(n5133), .ZN(n5140) );
  OR2_X1 U6221 ( .A1(n5136), .A2(n5135), .ZN(n5137) );
  NAND2_X1 U6222 ( .A1(n5215), .A2(n5465), .ZN(n5139) );
  OAI211_X1 U6223 ( .C1(n5449), .C2(n5282), .A(n5140), .B(n5139), .ZN(U2806)
         );
  AOI22_X1 U6224 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n5519), .B1(n5141), 
        .B2(n5520), .ZN(n5148) );
  OAI22_X1 U6225 ( .A1(n5143), .A2(n5452), .B1(n5449), .B2(n5142), .ZN(n5144)
         );
  AOI221_X1 U6226 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5146), .C1(n5145), .C2(
        n5146), .A(n5144), .ZN(n5147) );
  OAI211_X1 U6227 ( .C1(n3944), .C2(n5505), .A(n5148), .B(n5147), .ZN(U2807)
         );
  OAI21_X1 U6228 ( .B1(n4935), .B2(n4938), .A(n5150), .ZN(n5151) );
  OAI21_X1 U6229 ( .B1(n5152), .B2(n4938), .A(n5151), .ZN(n5306) );
  INV_X1 U6230 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5153) );
  OAI22_X1 U6231 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5154), .B1(n5153), .B2(
        n5499), .ZN(n5155) );
  AOI211_X1 U6232 ( .C1(n5518), .C2(EBX_REG_19__SCAN_IN), .A(n5483), .B(n5155), 
        .ZN(n5166) );
  AND2_X1 U6233 ( .A1(n5157), .A2(n5156), .ZN(n5159) );
  INV_X1 U6234 ( .A(n5387), .ZN(n5160) );
  AOI21_X1 U6235 ( .B1(n5161), .B2(n6487), .A(n5160), .ZN(n5163) );
  OAI22_X1 U6236 ( .A1(n5163), .A2(n5162), .B1(n5223), .B2(n5512), .ZN(n5164)
         );
  AOI21_X1 U6237 ( .B1(n3100), .B2(n5465), .A(n5164), .ZN(n5165) );
  OAI211_X1 U6238 ( .C1(n5449), .C2(n5306), .A(n5166), .B(n5165), .ZN(U2808)
         );
  INV_X1 U6239 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6572) );
  AOI22_X1 U6240 ( .A1(n3104), .A2(n5550), .B1(n5549), .B2(n5267), .ZN(n5167)
         );
  OAI21_X1 U6241 ( .B1(n5554), .B2(n6572), .A(n5167), .ZN(U2836) );
  AOI22_X1 U6242 ( .A1(n5215), .A2(n5550), .B1(EBX_REG_21__SCAN_IN), .B2(n5535), .ZN(n5168) );
  OAI21_X1 U6243 ( .B1(n5282), .B2(n5553), .A(n5168), .ZN(U2838) );
  AOI22_X1 U6244 ( .A1(n3100), .A2(n5550), .B1(EBX_REG_19__SCAN_IN), .B2(n5535), .ZN(n5169) );
  OAI21_X1 U6245 ( .B1(n5553), .B2(n5306), .A(n5169), .ZN(U2840) );
  AOI22_X1 U6246 ( .A1(n5170), .A2(n5563), .B1(n5556), .B2(DATAI_30_), .ZN(
        n5172) );
  AOI22_X1 U6247 ( .A1(n5559), .A2(DATAI_14_), .B1(n5558), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6248 ( .A1(n5172), .A2(n5171), .ZN(U2861) );
  AOI22_X1 U6249 ( .A1(n5173), .A2(n5563), .B1(n5556), .B2(DATAI_29_), .ZN(
        n5175) );
  AOI22_X1 U6250 ( .A1(n5559), .A2(DATAI_13_), .B1(n5558), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6251 ( .A1(n5175), .A2(n5174), .ZN(U2862) );
  OAI22_X1 U6252 ( .A1(n5179), .A2(n5178), .B1(n5177), .B2(n5176), .ZN(n5180)
         );
  INV_X1 U6253 ( .A(n5180), .ZN(n5182) );
  AOI22_X1 U6254 ( .A1(n5559), .A2(DATAI_12_), .B1(n5558), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6255 ( .A1(n5182), .A2(n5181), .ZN(U2863) );
  AOI22_X1 U6256 ( .A1(n5199), .A2(n5563), .B1(n5556), .B2(DATAI_27_), .ZN(
        n5184) );
  AOI22_X1 U6257 ( .A1(n5559), .A2(DATAI_11_), .B1(n5558), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6258 ( .A1(n5184), .A2(n5183), .ZN(U2864) );
  AOI22_X1 U6259 ( .A1(n5207), .A2(n5563), .B1(n5556), .B2(DATAI_25_), .ZN(
        n5186) );
  AOI22_X1 U6260 ( .A1(n5559), .A2(DATAI_9_), .B1(n5558), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6261 ( .A1(n5186), .A2(n5185), .ZN(U2866) );
  AOI22_X1 U6262 ( .A1(n3104), .A2(n5563), .B1(n5556), .B2(DATAI_23_), .ZN(
        n5188) );
  AOI22_X1 U6263 ( .A1(n5559), .A2(DATAI_7_), .B1(n5558), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6264 ( .A1(n5188), .A2(n5187), .ZN(U2868) );
  AOI22_X1 U6265 ( .A1(n5189), .A2(n5563), .B1(n5556), .B2(DATAI_22_), .ZN(
        n5191) );
  AOI22_X1 U6266 ( .A1(n5559), .A2(DATAI_6_), .B1(n5558), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6267 ( .A1(n5191), .A2(n5190), .ZN(U2869) );
  AOI22_X1 U6268 ( .A1(n5215), .A2(n5563), .B1(n5556), .B2(DATAI_21_), .ZN(
        n5193) );
  AOI22_X1 U6269 ( .A1(n5559), .A2(DATAI_5_), .B1(n5558), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6270 ( .A1(n5193), .A2(n5192), .ZN(U2870) );
  AOI22_X1 U6271 ( .A1(n3100), .A2(n5563), .B1(n5556), .B2(DATAI_19_), .ZN(
        n5195) );
  AOI22_X1 U6272 ( .A1(n5559), .A2(DATAI_3_), .B1(n5558), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6273 ( .A1(n5195), .A2(n5194), .ZN(U2872) );
  AOI22_X1 U6274 ( .A1(n5348), .A2(REIP_REG_27__SCAN_IN), .B1(n5662), .B2(
        PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5201) );
  NOR2_X1 U6275 ( .A1(n5197), .A2(n5196), .ZN(n5198) );
  XNOR2_X1 U6276 ( .A(n5198), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5248)
         );
  AOI22_X1 U6277 ( .A1(n5248), .A2(n5679), .B1(n5669), .B2(n5199), .ZN(n5200)
         );
  OAI211_X1 U6278 ( .C1(n5673), .C2(n5202), .A(n5201), .B(n5200), .ZN(U2959)
         );
  AOI22_X1 U6279 ( .A1(n5348), .A2(REIP_REG_25__SCAN_IN), .B1(n5662), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5209) );
  OAI21_X1 U6280 ( .B1(n5205), .B2(n5204), .A(n5203), .ZN(n5260) );
  OAI211_X1 U6281 ( .C1(n5673), .C2(n5210), .A(n5209), .B(n5208), .ZN(U2961)
         );
  INV_X1 U6282 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6720) );
  AOI21_X1 U6283 ( .B1(n5213), .B2(n5212), .A(n5211), .ZN(n5283) );
  INV_X1 U6284 ( .A(n5283), .ZN(n5217) );
  INV_X1 U6285 ( .A(n5214), .ZN(n5216) );
  AOI222_X1 U6286 ( .A1(n5217), .A2(n5679), .B1(n5216), .B2(n5233), .C1(n5669), 
        .C2(n5215), .ZN(n5218) );
  NAND2_X1 U6287 ( .A1(n5348), .A2(REIP_REG_21__SCAN_IN), .ZN(n5286) );
  OAI211_X1 U6288 ( .C1(n6720), .C2(n5676), .A(n5218), .B(n5286), .ZN(U2965)
         );
  AOI22_X1 U6289 ( .A1(n5348), .A2(REIP_REG_19__SCAN_IN), .B1(n5662), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5222) );
  XNOR2_X1 U6290 ( .A(n5220), .B(n5219), .ZN(n5304) );
  AOI22_X1 U6291 ( .A1(n5304), .A2(n5679), .B1(n5669), .B2(n3100), .ZN(n5221)
         );
  OAI211_X1 U6292 ( .C1(n5673), .C2(n5223), .A(n5222), .B(n5221), .ZN(U2967)
         );
  INV_X1 U6293 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5396) );
  OR2_X1 U6294 ( .A1(n5224), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5226)
         );
  NAND3_X1 U6295 ( .A1(n5227), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5224), .ZN(n5225) );
  OAI21_X1 U6296 ( .B1(n5227), .B2(n5226), .A(n5225), .ZN(n5228) );
  XNOR2_X1 U6297 ( .A(n5228), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5316)
         );
  INV_X1 U6298 ( .A(n5316), .ZN(n5235) );
  INV_X1 U6299 ( .A(n5392), .ZN(n5234) );
  OR2_X1 U6300 ( .A1(n5230), .A2(n5229), .ZN(n5231) );
  AND2_X1 U6301 ( .A1(n5232), .A2(n5231), .ZN(n5557) );
  AOI222_X1 U6302 ( .A1(n5235), .A2(n5679), .B1(n5234), .B2(n5233), .C1(n5669), 
        .C2(n5557), .ZN(n5236) );
  NAND2_X1 U6303 ( .A1(n5348), .A2(REIP_REG_17__SCAN_IN), .ZN(n5319) );
  OAI211_X1 U6304 ( .C1(n5396), .C2(n5676), .A(n5236), .B(n5319), .ZN(U2969)
         );
  AOI22_X1 U6305 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n5247), .B1(n5348), .B2(REIP_REG_28__SCAN_IN), .ZN(n5245) );
  INV_X1 U6306 ( .A(n5239), .ZN(n5240) );
  NOR2_X1 U6307 ( .A1(n5240), .A2(n5252), .ZN(n5242) );
  AOI22_X1 U6308 ( .A1(n5764), .A2(n5243), .B1(n5242), .B2(n5241), .ZN(n5244)
         );
  OAI211_X1 U6309 ( .C1(n5771), .C2(n5246), .A(n5245), .B(n5244), .ZN(U2990)
         );
  AOI22_X1 U6310 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n5247), .B1(n5348), .B2(REIP_REG_27__SCAN_IN), .ZN(n5251) );
  AOI22_X1 U6311 ( .A1(n5754), .A2(n5249), .B1(n5764), .B2(n5248), .ZN(n5250)
         );
  OAI211_X1 U6312 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5252), .A(n5251), .B(n5250), .ZN(U2991) );
  AOI22_X1 U6313 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n5262), .B1(n5348), .B2(REIP_REG_26__SCAN_IN), .ZN(n5257) );
  AOI22_X1 U6314 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .B1(n4082), .B2(n5253), .ZN(n5254)
         );
  AOI22_X1 U6315 ( .A1(n5255), .A2(n5764), .B1(n5263), .B2(n5254), .ZN(n5256)
         );
  OAI211_X1 U6316 ( .C1(n5771), .C2(n5258), .A(n5257), .B(n5256), .ZN(U2992)
         );
  AOI22_X1 U6317 ( .A1(n5260), .A2(n5764), .B1(n5754), .B2(n5259), .ZN(n5265)
         );
  NOR2_X1 U6318 ( .A1(n5740), .A2(n6504), .ZN(n5261) );
  AOI221_X1 U6319 ( .B1(n5263), .B2(n4082), .C1(n5262), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5261), .ZN(n5264) );
  NAND2_X1 U6320 ( .A1(n5265), .A2(n5264), .ZN(U2993) );
  AOI22_X1 U6321 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n5266), .B1(n5348), .B2(REIP_REG_23__SCAN_IN), .ZN(n5271) );
  OAI211_X1 U6322 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5272), .A(n5271), .B(n5270), .ZN(U2995) );
  NAND2_X1 U6323 ( .A1(n5285), .A2(n5273), .ZN(n5274) );
  OAI22_X1 U6324 ( .A1(n5276), .A2(n5771), .B1(n5275), .B2(n5274), .ZN(n5277)
         );
  AOI21_X1 U6325 ( .B1(n5278), .B2(n5764), .A(n5277), .ZN(n5280) );
  NAND2_X1 U6326 ( .A1(n5348), .A2(REIP_REG_22__SCAN_IN), .ZN(n5279) );
  OAI211_X1 U6327 ( .C1(n5289), .C2(n5281), .A(n5280), .B(n5279), .ZN(U2996)
         );
  OAI22_X1 U6328 ( .A1(n5283), .A2(n5733), .B1(n5771), .B2(n5282), .ZN(n5284)
         );
  AOI21_X1 U6329 ( .B1(n5285), .B2(n5288), .A(n5284), .ZN(n5287) );
  OAI211_X1 U6330 ( .C1(n5289), .C2(n5288), .A(n5287), .B(n5286), .ZN(U2997)
         );
  AOI221_X1 U6331 ( .B1(n5321), .B2(n5721), .C1(n5291), .C2(n5721), .A(n5290), 
        .ZN(n5322) );
  OAI21_X1 U6332 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5752), .A(n5322), 
        .ZN(n5310) );
  AOI21_X1 U6333 ( .B1(n3941), .B2(n5757), .A(n5310), .ZN(n5301) );
  NOR3_X1 U6334 ( .A1(n5293), .A2(n5292), .A3(n5302), .ZN(n5294) );
  AOI21_X1 U6335 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5348), .A(n5294), .ZN(n5298) );
  AOI22_X1 U6336 ( .A1(n5296), .A2(n5764), .B1(n5754), .B2(n5295), .ZN(n5297)
         );
  OAI211_X1 U6337 ( .C1(n5299), .C2(n5301), .A(n5298), .B(n5297), .ZN(U2998)
         );
  NAND2_X1 U6338 ( .A1(n5348), .A2(REIP_REG_19__SCAN_IN), .ZN(n5300) );
  OAI221_X1 U6339 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5302), .C1(
        n6701), .C2(n5301), .A(n5300), .ZN(n5303) );
  AOI21_X1 U6340 ( .B1(n5304), .B2(n5764), .A(n5303), .ZN(n5305) );
  OAI21_X1 U6341 ( .B1(n5771), .B2(n5306), .A(n5305), .ZN(U2999) );
  AOI22_X1 U6342 ( .A1(n5754), .A2(n5308), .B1(n5764), .B2(n5307), .ZN(n5312)
         );
  NOR2_X1 U6343 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5321), .ZN(n5309)
         );
  AOI22_X1 U6344 ( .A1(n5310), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .B1(n5318), .B2(n5309), .ZN(n5311) );
  OAI211_X1 U6345 ( .C1(n6487), .C2(n5740), .A(n5312), .B(n5311), .ZN(U3000)
         );
  OR2_X1 U6346 ( .A1(n5314), .A2(n5313), .ZN(n5315) );
  NAND2_X1 U6347 ( .A1(n4935), .A2(n5315), .ZN(n5534) );
  OAI22_X1 U6348 ( .A1(n5316), .A2(n5733), .B1(n5771), .B2(n5534), .ZN(n5317)
         );
  AOI21_X1 U6349 ( .B1(n5318), .B2(n5321), .A(n5317), .ZN(n5320) );
  OAI211_X1 U6350 ( .C1(n5322), .C2(n5321), .A(n5320), .B(n5319), .ZN(U3001)
         );
  AOI21_X1 U6351 ( .B1(n5757), .B2(n5323), .A(n5684), .ZN(n5337) );
  AOI21_X1 U6352 ( .B1(n5340), .B2(n6682), .A(n5336), .ZN(n5325) );
  AOI22_X1 U6353 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5348), .B1(n5325), .B2(
        n5324), .ZN(n5330) );
  INV_X1 U6354 ( .A(n5326), .ZN(n5328) );
  AOI22_X1 U6355 ( .A1(n5328), .A2(n5764), .B1(n5754), .B2(n5327), .ZN(n5329)
         );
  OAI211_X1 U6356 ( .C1(n5337), .C2(n6682), .A(n5330), .B(n5329), .ZN(U3002)
         );
  INV_X1 U6357 ( .A(n5331), .ZN(n5334) );
  INV_X1 U6358 ( .A(n5332), .ZN(n5333) );
  OAI21_X1 U6359 ( .B1(n5335), .B2(n5334), .A(n5333), .ZN(n5538) );
  INV_X1 U6360 ( .A(n5336), .ZN(n5341) );
  OAI22_X1 U6361 ( .A1(n5338), .A2(n5733), .B1(n5337), .B2(n5340), .ZN(n5339)
         );
  AOI21_X1 U6362 ( .B1(n5341), .B2(n5340), .A(n5339), .ZN(n5343) );
  NAND2_X1 U6363 ( .A1(n5348), .A2(REIP_REG_15__SCAN_IN), .ZN(n5342) );
  OAI211_X1 U6364 ( .C1(n5771), .C2(n5538), .A(n5343), .B(n5342), .ZN(U3003)
         );
  AOI221_X1 U6365 ( .B1(n5347), .B2(n5346), .C1(n5345), .C2(n5346), .A(n5344), 
        .ZN(n5355) );
  AOI22_X1 U6366 ( .A1(n5754), .A2(n5349), .B1(n5348), .B2(
        REIP_REG_14__SCAN_IN), .ZN(n5353) );
  AOI22_X1 U6367 ( .A1(n5351), .A2(n5764), .B1(n5350), .B2(n5354), .ZN(n5352)
         );
  OAI211_X1 U6368 ( .C1(n5355), .C2(n5354), .A(n5353), .B(n5352), .ZN(U3004)
         );
  INV_X1 U6369 ( .A(n5356), .ZN(n5359) );
  NAND4_X1 U6370 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5482), .ZN(n5360)
         );
  OAI21_X1 U6371 ( .B1(n6394), .B2(n6586), .A(n5360), .ZN(U3455) );
  OAI21_X1 U6372 ( .B1(STATE_REG_2__SCAN_IN), .B2(n6322), .A(
        STATE_REG_0__SCAN_IN), .ZN(n5367) );
  NOR2_X1 U6373 ( .A1(ADS_N_REG_SCAN_IN), .A2(n5367), .ZN(n5361) );
  NOR2_X1 U6374 ( .A1(n6429), .A2(n5361), .ZN(U2789) );
  OAI22_X1 U6375 ( .A1(n6282), .A2(n3095), .B1(n5363), .B2(n5362), .ZN(n5370)
         );
  OAI21_X1 U6376 ( .B1(n6305), .B2(n5370), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5365) );
  OAI21_X1 U6377 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6306), .A(n5365), .ZN(
        U2790) );
  INV_X1 U6378 ( .A(n6429), .ZN(n6336) );
  NOR2_X1 U6379 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5368) );
  OAI21_X1 U6380 ( .B1(n5368), .B2(D_C_N_REG_SCAN_IN), .A(n6375), .ZN(n5366)
         );
  OAI21_X1 U6381 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6336), .A(n5366), .ZN(
        U2791) );
  NAND2_X1 U6382 ( .A1(n6336), .A2(n5367), .ZN(n6750) );
  INV_X1 U6383 ( .A(n6750), .ZN(n6380) );
  OAI21_X1 U6384 ( .B1(n5368), .B2(BS16_N), .A(n6380), .ZN(n6378) );
  OAI21_X1 U6385 ( .B1(n6380), .B2(n6164), .A(n6378), .ZN(U2792) );
  NAND2_X1 U6386 ( .A1(n6423), .A2(n5369), .ZN(n6433) );
  AOI21_X1 U6387 ( .B1(n6433), .B2(n6321), .A(READY_N), .ZN(n6422) );
  NOR2_X1 U6388 ( .A1(n6422), .A2(n5370), .ZN(n6273) );
  NOR2_X1 U6389 ( .A1(n6273), .A2(n6305), .ZN(n6418) );
  OAI21_X1 U6390 ( .B1(n6418), .B2(n5372), .A(n5371), .ZN(U2793) );
  NOR2_X1 U6391 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6446) );
  AOI211_X1 U6392 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_28__SCAN_IN), .B(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n5373) );
  INV_X1 U6393 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6518) );
  INV_X1 U6394 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6719) );
  NAND4_X1 U6395 ( .A1(n6446), .A2(n5373), .A3(n6518), .A4(n6719), .ZN(n5381)
         );
  OR4_X1 U6396 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n5380) );
  INV_X1 U6397 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6536) );
  INV_X1 U6398 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6629) );
  INV_X1 U6399 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6632) );
  INV_X1 U6400 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6553) );
  NAND4_X1 U6401 ( .A1(n6536), .A2(n6629), .A3(n6632), .A4(n6553), .ZN(n5379)
         );
  NOR4_X1 U6402 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5377) );
  NOR4_X1 U6403 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5376) );
  NOR4_X1 U6404 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n5375) );
  NOR4_X1 U6405 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n5374) );
  NAND4_X1 U6406 ( .A1(n5377), .A2(n5376), .A3(n5375), .A4(n5374), .ZN(n5378)
         );
  NOR4_X2 U6407 ( .A1(n5381), .A2(n5380), .A3(n5379), .A4(n5378), .ZN(n6414)
         );
  INV_X1 U6408 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5383) );
  NOR3_X1 U6409 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5384) );
  OAI21_X1 U6410 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5384), .A(n6414), .ZN(n5382)
         );
  OAI21_X1 U6411 ( .B1(n6414), .B2(n5383), .A(n5382), .ZN(U2794) );
  INV_X1 U6412 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6379) );
  AOI21_X1 U6413 ( .B1(n6407), .B2(n6379), .A(n5384), .ZN(n5386) );
  INV_X1 U6414 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5385) );
  INV_X1 U6415 ( .A(n6414), .ZN(n6409) );
  AOI22_X1 U6416 ( .A1(n6414), .A2(n5386), .B1(n5385), .B2(n6409), .ZN(U2795)
         );
  AOI21_X1 U6417 ( .B1(n6622), .B2(n5388), .A(n5387), .ZN(n5389) );
  AOI211_X1 U6418 ( .C1(n5518), .C2(EBX_REG_17__SCAN_IN), .A(n5483), .B(n5389), 
        .ZN(n5395) );
  INV_X1 U6419 ( .A(n5534), .ZN(n5390) );
  NAND2_X1 U6420 ( .A1(n5517), .A2(n5390), .ZN(n5391) );
  OAI21_X1 U6421 ( .B1(n5512), .B2(n5392), .A(n5391), .ZN(n5393) );
  AOI21_X1 U6422 ( .B1(n5557), .B2(n5465), .A(n5393), .ZN(n5394) );
  OAI211_X1 U6423 ( .C1(n5396), .C2(n5499), .A(n5395), .B(n5394), .ZN(U2810)
         );
  AOI211_X1 U6424 ( .C1(n5519), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5483), 
        .B(n5397), .ZN(n5400) );
  AOI22_X1 U6425 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5518), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5398), .ZN(n5399) );
  NAND2_X1 U6426 ( .A1(n5400), .A2(n5399), .ZN(n5401) );
  AOI21_X1 U6427 ( .B1(n5536), .B2(n5465), .A(n5401), .ZN(n5404) );
  NAND2_X1 U6428 ( .A1(n5402), .A2(n5520), .ZN(n5403) );
  OAI211_X1 U6429 ( .C1(n5538), .C2(n5449), .A(n5404), .B(n5403), .ZN(U2812)
         );
  AOI22_X1 U6430 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5518), .B1(n5517), .B2(n5539), .ZN(n5413) );
  NOR3_X1 U6431 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5487), .A3(n5405), .ZN(n5406) );
  AOI211_X1 U6432 ( .C1(n5519), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5483), 
        .B(n5406), .ZN(n5412) );
  INV_X1 U6433 ( .A(n5407), .ZN(n5408) );
  AOI22_X1 U6434 ( .A1(n5564), .A2(n5465), .B1(n5520), .B2(n5408), .ZN(n5411)
         );
  INV_X1 U6435 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6651) );
  AND3_X1 U6436 ( .A1(n6651), .A2(n5513), .A3(n5409), .ZN(n5415) );
  OAI21_X1 U6437 ( .B1(n5416), .B2(n5415), .A(REIP_REG_13__SCAN_IN), .ZN(n5410) );
  NAND4_X1 U6438 ( .A1(n5413), .A2(n5412), .A3(n5411), .A4(n5410), .ZN(U2814)
         );
  AOI22_X1 U6439 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n5519), .B1(n5517), 
        .B2(n5541), .ZN(n5420) );
  INV_X1 U6440 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5544) );
  NOR2_X1 U6441 ( .A1(n5544), .A2(n5505), .ZN(n5414) );
  AOI211_X1 U6442 ( .C1(n5416), .C2(REIP_REG_12__SCAN_IN), .A(n5415), .B(n5414), .ZN(n5419) );
  AOI22_X1 U6443 ( .A1(n5542), .A2(n5465), .B1(n5520), .B2(n5417), .ZN(n5418)
         );
  NAND4_X1 U6444 ( .A1(n5420), .A2(n5419), .A3(n5418), .A4(n5472), .ZN(U2815)
         );
  OAI21_X1 U6445 ( .B1(REIP_REG_10__SCAN_IN), .B2(REIP_REG_9__SCAN_IN), .A(
        n5421), .ZN(n5431) );
  INV_X1 U6446 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5548) );
  INV_X1 U6447 ( .A(n5422), .ZN(n5425) );
  AOI21_X1 U6448 ( .B1(n5513), .B2(n5423), .A(n5507), .ZN(n5475) );
  OAI21_X1 U6449 ( .B1(n5425), .B2(n5424), .A(n5475), .ZN(n5443) );
  AOI22_X1 U6450 ( .A1(n5517), .A2(n5545), .B1(REIP_REG_10__SCAN_IN), .B2(
        n5443), .ZN(n5426) );
  OAI21_X1 U6451 ( .B1(n5548), .B2(n5505), .A(n5426), .ZN(n5427) );
  AOI211_X1 U6452 ( .C1(n5519), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5483), 
        .B(n5427), .ZN(n5430) );
  AOI22_X1 U6453 ( .A1(n5546), .A2(n5465), .B1(n5520), .B2(n5428), .ZN(n5429)
         );
  OAI211_X1 U6454 ( .C1(n5439), .C2(n5431), .A(n5430), .B(n5429), .ZN(U2817)
         );
  AOI22_X1 U6455 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5518), .B1(n5517), .B2(n5691), 
        .ZN(n5432) );
  OAI211_X1 U6456 ( .C1(n5499), .C2(n6638), .A(n5432), .B(n5472), .ZN(n5433)
         );
  AOI21_X1 U6457 ( .B1(REIP_REG_9__SCAN_IN), .B2(n5443), .A(n5433), .ZN(n5438)
         );
  OAI22_X1 U6458 ( .A1(n5435), .A2(n5452), .B1(n5434), .B2(n5512), .ZN(n5436)
         );
  INV_X1 U6459 ( .A(n5436), .ZN(n5437) );
  OAI211_X1 U6460 ( .C1(REIP_REG_9__SCAN_IN), .C2(n5439), .A(n5438), .B(n5437), 
        .ZN(U2818) );
  AOI22_X1 U6461 ( .A1(EBX_REG_8__SCAN_IN), .A2(n5518), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n5519), .ZN(n5448) );
  AOI21_X1 U6462 ( .B1(n5517), .B2(n5701), .A(n5483), .ZN(n5447) );
  INV_X1 U6463 ( .A(n5440), .ZN(n5442) );
  AOI22_X1 U6464 ( .A1(n5442), .A2(n5465), .B1(n5520), .B2(n5441), .ZN(n5446)
         );
  OAI21_X1 U6465 ( .B1(REIP_REG_8__SCAN_IN), .B2(n5444), .A(n5443), .ZN(n5445)
         );
  NAND4_X1 U6466 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(U2819)
         );
  OAI22_X1 U6467 ( .A1(n5449), .A2(n5712), .B1(n6340), .B2(n5475), .ZN(n5450)
         );
  AOI211_X1 U6468 ( .C1(n5519), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5483), 
        .B(n5450), .ZN(n5458) );
  AOI21_X1 U6469 ( .B1(n6340), .B2(n4509), .A(n5469), .ZN(n5456) );
  OAI22_X1 U6470 ( .A1(n5453), .A2(n5452), .B1(n5451), .B2(n5512), .ZN(n5454)
         );
  AOI21_X1 U6471 ( .B1(n5456), .B2(n5455), .A(n5454), .ZN(n5457) );
  OAI211_X1 U6472 ( .C1(n5459), .C2(n5505), .A(n5458), .B(n5457), .ZN(U2820)
         );
  INV_X1 U6473 ( .A(n5460), .ZN(n5717) );
  AOI22_X1 U6474 ( .A1(EBX_REG_6__SCAN_IN), .A2(n5518), .B1(n5517), .B2(n5717), 
        .ZN(n5461) );
  OAI21_X1 U6475 ( .B1(n4509), .B2(n5475), .A(n5461), .ZN(n5462) );
  AOI211_X1 U6476 ( .C1(n5519), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5483), 
        .B(n5462), .ZN(n5468) );
  INV_X1 U6477 ( .A(n5463), .ZN(n5466) );
  AOI22_X1 U6478 ( .A1(n5466), .A2(n5465), .B1(n5464), .B2(n5520), .ZN(n5467)
         );
  OAI211_X1 U6479 ( .C1(REIP_REG_6__SCAN_IN), .C2(n5469), .A(n5468), .B(n5467), 
        .ZN(U2821) );
  INV_X1 U6480 ( .A(n5470), .ZN(n5479) );
  INV_X1 U6481 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5474) );
  AOI22_X1 U6482 ( .A1(EBX_REG_5__SCAN_IN), .A2(n5518), .B1(n5517), .B2(n5471), 
        .ZN(n5473) );
  OAI211_X1 U6483 ( .C1(n5499), .C2(n5474), .A(n5473), .B(n5472), .ZN(n5478)
         );
  NAND3_X1 U6484 ( .A1(n5513), .A2(REIP_REG_4__SCAN_IN), .A3(n5488), .ZN(n5476) );
  AOI21_X1 U6485 ( .B1(n6339), .B2(n5476), .A(n5475), .ZN(n5477) );
  AOI211_X1 U6486 ( .C1(n5479), .C2(n5523), .A(n5478), .B(n5477), .ZN(n5480)
         );
  OAI21_X1 U6487 ( .B1(n5481), .B2(n5512), .A(n5480), .ZN(U2822) );
  NAND2_X1 U6488 ( .A1(n5513), .A2(n5488), .ZN(n5495) );
  AOI22_X1 U6489 ( .A1(EBX_REG_4__SCAN_IN), .A2(n5518), .B1(n5482), .B2(n5522), 
        .ZN(n5494) );
  AOI21_X1 U6490 ( .B1(n5519), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5483), 
        .ZN(n5484) );
  OAI21_X1 U6491 ( .B1(n5512), .B2(n5485), .A(n5484), .ZN(n5491) );
  OAI21_X1 U6492 ( .B1(n5488), .B2(n5487), .A(n5486), .ZN(n5508) );
  AOI22_X1 U6493 ( .A1(n5517), .A2(n5729), .B1(REIP_REG_4__SCAN_IN), .B2(n5508), .ZN(n5489) );
  INV_X1 U6494 ( .A(n5489), .ZN(n5490) );
  AOI211_X1 U6495 ( .C1(n5492), .C2(n5523), .A(n5491), .B(n5490), .ZN(n5493)
         );
  OAI211_X1 U6496 ( .C1(REIP_REG_4__SCAN_IN), .C2(n5495), .A(n5494), .B(n5493), 
        .ZN(U2823) );
  INV_X1 U6497 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6498 ( .A1(n5517), .A2(n5737), .ZN(n5497) );
  NAND2_X1 U6499 ( .A1(n5522), .A2(n6017), .ZN(n5496) );
  OAI211_X1 U6500 ( .C1(n5499), .C2(n5498), .A(n5497), .B(n5496), .ZN(n5500)
         );
  INV_X1 U6501 ( .A(n5500), .ZN(n5504) );
  INV_X1 U6502 ( .A(n5501), .ZN(n5502) );
  NAND2_X1 U6503 ( .A1(n5523), .A2(n5502), .ZN(n5503) );
  OAI211_X1 U6504 ( .C1(n5505), .C2(n6499), .A(n5504), .B(n5503), .ZN(n5506)
         );
  INV_X1 U6505 ( .A(n5506), .ZN(n5510) );
  AOI211_X1 U6506 ( .C1(n5513), .C2(n6407), .A(n5507), .B(n6333), .ZN(n5530)
         );
  OAI21_X1 U6507 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5530), .A(n5508), .ZN(n5509)
         );
  OAI211_X1 U6508 ( .C1(n5512), .C2(n5511), .A(n5510), .B(n5509), .ZN(U2824)
         );
  AOI21_X1 U6509 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5513), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5529) );
  OAI21_X1 U6510 ( .B1(n5515), .B2(n5514), .A(n4255), .ZN(n5516) );
  INV_X1 U6511 ( .A(n5516), .ZN(n5746) );
  AOI22_X1 U6512 ( .A1(EBX_REG_2__SCAN_IN), .A2(n5518), .B1(n5517), .B2(n5746), 
        .ZN(n5527) );
  INV_X1 U6513 ( .A(n5672), .ZN(n5521) );
  AOI22_X1 U6514 ( .A1(n5521), .A2(n5520), .B1(n5519), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5526) );
  INV_X1 U6515 ( .A(n5774), .ZN(n6401) );
  NAND2_X1 U6516 ( .A1(n5522), .A2(n6401), .ZN(n5525) );
  NAND2_X1 U6517 ( .A1(n5523), .A2(n5668), .ZN(n5524) );
  AND4_X1 U6518 ( .A1(n5527), .A2(n5526), .A3(n5525), .A4(n5524), .ZN(n5528)
         );
  OAI21_X1 U6519 ( .B1(n5530), .B2(n5529), .A(n5528), .ZN(U2825) );
  AOI22_X1 U6520 ( .A1(n5535), .A2(EBX_REG_31__SCAN_IN), .B1(n5531), .B2(n5549), .ZN(n5532) );
  INV_X1 U6521 ( .A(n5532), .ZN(U2828) );
  AOI22_X1 U6522 ( .A1(n5557), .A2(n5550), .B1(EBX_REG_17__SCAN_IN), .B2(n5535), .ZN(n5533) );
  OAI21_X1 U6523 ( .B1(n5553), .B2(n5534), .A(n5533), .ZN(U2842) );
  AOI22_X1 U6524 ( .A1(n5536), .A2(n5550), .B1(EBX_REG_15__SCAN_IN), .B2(n5535), .ZN(n5537) );
  OAI21_X1 U6525 ( .B1(n5553), .B2(n5538), .A(n5537), .ZN(U2844) );
  INV_X1 U6526 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6530) );
  AOI22_X1 U6527 ( .A1(n5564), .A2(n5550), .B1(n5549), .B2(n5539), .ZN(n5540)
         );
  OAI21_X1 U6528 ( .B1(n5554), .B2(n6530), .A(n5540), .ZN(U2846) );
  AOI22_X1 U6529 ( .A1(n5542), .A2(n5550), .B1(n5549), .B2(n5541), .ZN(n5543)
         );
  OAI21_X1 U6530 ( .B1(n5554), .B2(n5544), .A(n5543), .ZN(U2847) );
  AOI22_X1 U6531 ( .A1(n5546), .A2(n5550), .B1(n5549), .B2(n5545), .ZN(n5547)
         );
  OAI21_X1 U6532 ( .B1(n5554), .B2(n5548), .A(n5547), .ZN(U2849) );
  INV_X1 U6533 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5552) );
  AOI22_X1 U6534 ( .A1(n5668), .A2(n5550), .B1(n5549), .B2(n5746), .ZN(n5551)
         );
  OAI21_X1 U6535 ( .B1(n5554), .B2(n5552), .A(n5551), .ZN(U2857) );
  OAI222_X1 U6536 ( .A1(n5683), .A2(n5555), .B1(n3885), .B2(n5554), .C1(n5553), 
        .C2(n5772), .ZN(U2859) );
  AOI22_X1 U6537 ( .A1(n5557), .A2(n5563), .B1(n5556), .B2(DATAI_17_), .ZN(
        n5561) );
  AOI22_X1 U6538 ( .A1(n5559), .A2(DATAI_1_), .B1(n5558), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U6539 ( .A1(n5561), .A2(n5560), .ZN(U2874) );
  AOI22_X1 U6540 ( .A1(n5564), .A2(n5563), .B1(DATAI_13_), .B2(n5562), .ZN(
        n5565) );
  OAI21_X1 U6541 ( .B1(n6562), .B2(n5566), .A(n5565), .ZN(U2878) );
  INV_X1 U6542 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U6543 ( .A1(n5583), .A2(n3882), .ZN(n5582) );
  AOI22_X1 U6544 ( .A1(n6421), .A2(UWORD_REG_14__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5567) );
  OAI21_X1 U6545 ( .B1(n5631), .B2(n5582), .A(n5567), .ZN(U2893) );
  INV_X1 U6546 ( .A(EAX_REG_29__SCAN_IN), .ZN(n5629) );
  AOI22_X1 U6547 ( .A1(n6421), .A2(UWORD_REG_13__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n5568) );
  OAI21_X1 U6548 ( .B1(n5629), .B2(n5582), .A(n5568), .ZN(U2894) );
  INV_X1 U6549 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6505) );
  AOI22_X1 U6550 ( .A1(n6421), .A2(UWORD_REG_12__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5569) );
  OAI21_X1 U6551 ( .B1(n6505), .B2(n5582), .A(n5569), .ZN(U2895) );
  AOI22_X1 U6552 ( .A1(n6421), .A2(UWORD_REG_11__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5570) );
  OAI21_X1 U6553 ( .B1(n4722), .B2(n5582), .A(n5570), .ZN(U2896) );
  INV_X1 U6554 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5625) );
  AOI22_X1 U6555 ( .A1(n6421), .A2(UWORD_REG_10__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5571) );
  OAI21_X1 U6556 ( .B1(n5625), .B2(n5582), .A(n5571), .ZN(U2897) );
  INV_X1 U6557 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5623) );
  AOI22_X1 U6558 ( .A1(n6421), .A2(UWORD_REG_9__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n5572) );
  OAI21_X1 U6559 ( .B1(n5623), .B2(n5582), .A(n5572), .ZN(U2898) );
  INV_X1 U6560 ( .A(EAX_REG_24__SCAN_IN), .ZN(n5621) );
  AOI22_X1 U6561 ( .A1(n6421), .A2(UWORD_REG_8__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5573) );
  OAI21_X1 U6562 ( .B1(n5621), .B2(n5582), .A(n5573), .ZN(U2899) );
  AOI22_X1 U6563 ( .A1(n6421), .A2(UWORD_REG_7__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5574) );
  OAI21_X1 U6564 ( .B1(n3766), .B2(n5582), .A(n5574), .ZN(U2900) );
  INV_X1 U6565 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5618) );
  AOI22_X1 U6566 ( .A1(n5593), .A2(UWORD_REG_6__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5575) );
  OAI21_X1 U6567 ( .B1(n5618), .B2(n5582), .A(n5575), .ZN(U2901) );
  INV_X1 U6568 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5616) );
  AOI22_X1 U6569 ( .A1(n5593), .A2(UWORD_REG_5__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5576) );
  OAI21_X1 U6570 ( .B1(n5616), .B2(n5582), .A(n5576), .ZN(U2902) );
  INV_X1 U6571 ( .A(EAX_REG_20__SCAN_IN), .ZN(n5614) );
  AOI22_X1 U6572 ( .A1(n5593), .A2(UWORD_REG_4__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5577) );
  OAI21_X1 U6573 ( .B1(n5614), .B2(n5582), .A(n5577), .ZN(U2903) );
  INV_X1 U6574 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5612) );
  AOI22_X1 U6575 ( .A1(n5593), .A2(UWORD_REG_3__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5578) );
  OAI21_X1 U6576 ( .B1(n5612), .B2(n5582), .A(n5578), .ZN(U2904) );
  INV_X1 U6577 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6613) );
  AOI22_X1 U6578 ( .A1(n5593), .A2(UWORD_REG_2__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5579) );
  OAI21_X1 U6579 ( .B1(n6613), .B2(n5582), .A(n5579), .ZN(U2905) );
  INV_X1 U6580 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5608) );
  AOI22_X1 U6581 ( .A1(n5593), .A2(UWORD_REG_1__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5580) );
  OAI21_X1 U6582 ( .B1(n5608), .B2(n5582), .A(n5580), .ZN(U2906) );
  INV_X1 U6583 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6700) );
  AOI22_X1 U6584 ( .A1(n5593), .A2(UWORD_REG_0__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5581) );
  OAI21_X1 U6585 ( .B1(n6700), .B2(n5582), .A(n5581), .ZN(U2907) );
  AOI22_X1 U6586 ( .A1(n5593), .A2(LWORD_REG_15__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5584) );
  OAI21_X1 U6587 ( .B1(n6729), .B2(n5602), .A(n5584), .ZN(U2908) );
  INV_X1 U6588 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5657) );
  AOI22_X1 U6589 ( .A1(n5593), .A2(LWORD_REG_14__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5585) );
  OAI21_X1 U6590 ( .B1(n5657), .B2(n5602), .A(n5585), .ZN(U2909) );
  AOI22_X1 U6591 ( .A1(n5593), .A2(LWORD_REG_13__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5586) );
  OAI21_X1 U6592 ( .B1(n6562), .B2(n5602), .A(n5586), .ZN(U2910) );
  INV_X1 U6593 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5654) );
  AOI22_X1 U6594 ( .A1(n6421), .A2(LWORD_REG_12__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5587) );
  OAI21_X1 U6595 ( .B1(n5654), .B2(n5602), .A(n5587), .ZN(U2911) );
  AOI22_X1 U6596 ( .A1(n6421), .A2(LWORD_REG_11__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5588) );
  OAI21_X1 U6597 ( .B1(n6596), .B2(n5602), .A(n5588), .ZN(U2912) );
  INV_X1 U6598 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5651) );
  AOI22_X1 U6599 ( .A1(n6421), .A2(LWORD_REG_10__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5589) );
  OAI21_X1 U6600 ( .B1(n5651), .B2(n5602), .A(n5589), .ZN(U2913) );
  AOI22_X1 U6601 ( .A1(n6421), .A2(LWORD_REG_9__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5590) );
  OAI21_X1 U6602 ( .B1(n6568), .B2(n5602), .A(n5590), .ZN(U2914) );
  INV_X1 U6603 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5647) );
  AOI22_X1 U6604 ( .A1(n6421), .A2(LWORD_REG_8__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5591) );
  OAI21_X1 U6605 ( .B1(n5647), .B2(n5602), .A(n5591), .ZN(U2915) );
  AOI22_X1 U6606 ( .A1(n6421), .A2(LWORD_REG_7__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5592) );
  OAI21_X1 U6607 ( .B1(n5644), .B2(n5602), .A(n5592), .ZN(U2916) );
  AOI22_X1 U6608 ( .A1(n5593), .A2(LWORD_REG_6__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5594) );
  OAI21_X1 U6609 ( .B1(n3462), .B2(n5602), .A(n5594), .ZN(U2917) );
  AOI22_X1 U6610 ( .A1(n6421), .A2(LWORD_REG_5__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5595) );
  OAI21_X1 U6611 ( .B1(n3444), .B2(n5602), .A(n5595), .ZN(U2918) );
  AOI22_X1 U6612 ( .A1(n6421), .A2(LWORD_REG_4__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5596) );
  OAI21_X1 U6613 ( .B1(n5640), .B2(n5602), .A(n5596), .ZN(U2919) );
  AOI22_X1 U6614 ( .A1(n6421), .A2(LWORD_REG_3__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5598) );
  OAI21_X1 U6615 ( .B1(n5638), .B2(n5602), .A(n5598), .ZN(U2920) );
  AOI22_X1 U6616 ( .A1(n6421), .A2(LWORD_REG_2__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5599) );
  OAI21_X1 U6617 ( .B1(n3359), .B2(n5602), .A(n5599), .ZN(U2921) );
  AOI22_X1 U6618 ( .A1(n6421), .A2(LWORD_REG_1__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5600) );
  OAI21_X1 U6619 ( .B1(n5635), .B2(n5602), .A(n5600), .ZN(U2922) );
  AOI22_X1 U6620 ( .A1(n6421), .A2(LWORD_REG_0__SCAN_IN), .B1(n5597), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5601) );
  OAI21_X1 U6621 ( .B1(n5633), .B2(n5602), .A(n5601), .ZN(U2923) );
  INV_X1 U6622 ( .A(n6296), .ZN(n5603) );
  AOI22_X1 U6623 ( .A1(n5645), .A2(DATAI_0_), .B1(UWORD_REG_0__SCAN_IN), .B2(
        n5648), .ZN(n5606) );
  OAI21_X1 U6624 ( .B1(n6700), .B2(n5661), .A(n5606), .ZN(U2924) );
  AOI22_X1 U6625 ( .A1(n5645), .A2(DATAI_1_), .B1(UWORD_REG_1__SCAN_IN), .B2(
        n5648), .ZN(n5607) );
  OAI21_X1 U6626 ( .B1(n5608), .B2(n5661), .A(n5607), .ZN(U2925) );
  INV_X1 U6627 ( .A(n5609), .ZN(n5659) );
  AOI22_X1 U6628 ( .A1(n5659), .A2(DATAI_2_), .B1(UWORD_REG_2__SCAN_IN), .B2(
        n5648), .ZN(n5610) );
  OAI21_X1 U6629 ( .B1(n6613), .B2(n5661), .A(n5610), .ZN(U2926) );
  AOI22_X1 U6630 ( .A1(n5645), .A2(DATAI_3_), .B1(UWORD_REG_3__SCAN_IN), .B2(
        n5648), .ZN(n5611) );
  OAI21_X1 U6631 ( .B1(n5612), .B2(n5661), .A(n5611), .ZN(U2927) );
  AOI22_X1 U6632 ( .A1(n5659), .A2(DATAI_4_), .B1(UWORD_REG_4__SCAN_IN), .B2(
        n5648), .ZN(n5613) );
  OAI21_X1 U6633 ( .B1(n5614), .B2(n5661), .A(n5613), .ZN(U2928) );
  AOI22_X1 U6634 ( .A1(n5645), .A2(DATAI_5_), .B1(UWORD_REG_5__SCAN_IN), .B2(
        n5648), .ZN(n5615) );
  OAI21_X1 U6635 ( .B1(n5616), .B2(n5661), .A(n5615), .ZN(U2929) );
  AOI22_X1 U6636 ( .A1(n5645), .A2(DATAI_6_), .B1(UWORD_REG_6__SCAN_IN), .B2(
        n5648), .ZN(n5617) );
  OAI21_X1 U6637 ( .B1(n5618), .B2(n5661), .A(n5617), .ZN(U2930) );
  AOI22_X1 U6638 ( .A1(n5659), .A2(DATAI_7_), .B1(UWORD_REG_7__SCAN_IN), .B2(
        n5648), .ZN(n5619) );
  OAI21_X1 U6639 ( .B1(n3766), .B2(n5661), .A(n5619), .ZN(U2931) );
  AOI22_X1 U6640 ( .A1(n5645), .A2(DATAI_8_), .B1(UWORD_REG_8__SCAN_IN), .B2(
        n5648), .ZN(n5620) );
  OAI21_X1 U6641 ( .B1(n5621), .B2(n5661), .A(n5620), .ZN(U2932) );
  AOI22_X1 U6642 ( .A1(n5659), .A2(DATAI_9_), .B1(UWORD_REG_9__SCAN_IN), .B2(
        n5648), .ZN(n5622) );
  OAI21_X1 U6643 ( .B1(n5623), .B2(n5661), .A(n5622), .ZN(U2933) );
  AOI22_X1 U6644 ( .A1(n5645), .A2(DATAI_10_), .B1(UWORD_REG_10__SCAN_IN), 
        .B2(n5648), .ZN(n5624) );
  OAI21_X1 U6645 ( .B1(n5625), .B2(n5661), .A(n5624), .ZN(U2934) );
  AOI22_X1 U6646 ( .A1(n5645), .A2(DATAI_11_), .B1(UWORD_REG_11__SCAN_IN), 
        .B2(n5648), .ZN(n5626) );
  OAI21_X1 U6647 ( .B1(n4722), .B2(n5661), .A(n5626), .ZN(U2935) );
  AOI22_X1 U6648 ( .A1(n5645), .A2(DATAI_12_), .B1(UWORD_REG_12__SCAN_IN), 
        .B2(n5658), .ZN(n5627) );
  OAI21_X1 U6649 ( .B1(n6505), .B2(n5661), .A(n5627), .ZN(U2936) );
  AOI22_X1 U6650 ( .A1(n5645), .A2(DATAI_13_), .B1(UWORD_REG_13__SCAN_IN), 
        .B2(n5658), .ZN(n5628) );
  OAI21_X1 U6651 ( .B1(n5629), .B2(n5661), .A(n5628), .ZN(U2937) );
  AOI22_X1 U6652 ( .A1(n5645), .A2(DATAI_14_), .B1(UWORD_REG_14__SCAN_IN), 
        .B2(n5658), .ZN(n5630) );
  OAI21_X1 U6653 ( .B1(n5631), .B2(n5661), .A(n5630), .ZN(U2938) );
  AOI22_X1 U6654 ( .A1(n5645), .A2(DATAI_0_), .B1(LWORD_REG_0__SCAN_IN), .B2(
        n5658), .ZN(n5632) );
  OAI21_X1 U6655 ( .B1(n5633), .B2(n5661), .A(n5632), .ZN(U2939) );
  AOI22_X1 U6656 ( .A1(n5645), .A2(DATAI_1_), .B1(LWORD_REG_1__SCAN_IN), .B2(
        n5648), .ZN(n5634) );
  OAI21_X1 U6657 ( .B1(n5635), .B2(n5661), .A(n5634), .ZN(U2940) );
  AOI22_X1 U6658 ( .A1(n5645), .A2(DATAI_2_), .B1(LWORD_REG_2__SCAN_IN), .B2(
        n5648), .ZN(n5636) );
  OAI21_X1 U6659 ( .B1(n3359), .B2(n5661), .A(n5636), .ZN(U2941) );
  AOI22_X1 U6660 ( .A1(n5645), .A2(DATAI_3_), .B1(LWORD_REG_3__SCAN_IN), .B2(
        n5648), .ZN(n5637) );
  OAI21_X1 U6661 ( .B1(n5638), .B2(n5661), .A(n5637), .ZN(U2942) );
  AOI22_X1 U6662 ( .A1(n5645), .A2(DATAI_4_), .B1(LWORD_REG_4__SCAN_IN), .B2(
        n5648), .ZN(n5639) );
  OAI21_X1 U6663 ( .B1(n5640), .B2(n5661), .A(n5639), .ZN(U2943) );
  AOI22_X1 U6664 ( .A1(n5645), .A2(DATAI_5_), .B1(LWORD_REG_5__SCAN_IN), .B2(
        n5648), .ZN(n5641) );
  OAI21_X1 U6665 ( .B1(n3444), .B2(n5661), .A(n5641), .ZN(U2944) );
  AOI22_X1 U6666 ( .A1(n5645), .A2(DATAI_6_), .B1(LWORD_REG_6__SCAN_IN), .B2(
        n5648), .ZN(n5642) );
  OAI21_X1 U6667 ( .B1(n3462), .B2(n5661), .A(n5642), .ZN(U2945) );
  AOI22_X1 U6668 ( .A1(n5645), .A2(DATAI_7_), .B1(LWORD_REG_7__SCAN_IN), .B2(
        n5648), .ZN(n5643) );
  OAI21_X1 U6669 ( .B1(n5644), .B2(n5661), .A(n5643), .ZN(U2946) );
  AOI22_X1 U6670 ( .A1(n5645), .A2(DATAI_8_), .B1(LWORD_REG_8__SCAN_IN), .B2(
        n5648), .ZN(n5646) );
  OAI21_X1 U6671 ( .B1(n5647), .B2(n5661), .A(n5646), .ZN(U2947) );
  AOI22_X1 U6672 ( .A1(n5659), .A2(DATAI_9_), .B1(LWORD_REG_9__SCAN_IN), .B2(
        n5648), .ZN(n5649) );
  OAI21_X1 U6673 ( .B1(n6568), .B2(n5661), .A(n5649), .ZN(U2948) );
  AOI22_X1 U6674 ( .A1(n5659), .A2(DATAI_10_), .B1(LWORD_REG_10__SCAN_IN), 
        .B2(n5658), .ZN(n5650) );
  OAI21_X1 U6675 ( .B1(n5651), .B2(n5661), .A(n5650), .ZN(U2949) );
  AOI22_X1 U6676 ( .A1(n5659), .A2(DATAI_11_), .B1(LWORD_REG_11__SCAN_IN), 
        .B2(n5658), .ZN(n5652) );
  OAI21_X1 U6677 ( .B1(n6596), .B2(n5661), .A(n5652), .ZN(U2950) );
  AOI22_X1 U6678 ( .A1(n5659), .A2(DATAI_12_), .B1(LWORD_REG_12__SCAN_IN), 
        .B2(n5658), .ZN(n5653) );
  OAI21_X1 U6679 ( .B1(n5654), .B2(n5661), .A(n5653), .ZN(U2951) );
  AOI22_X1 U6680 ( .A1(n5659), .A2(DATAI_13_), .B1(LWORD_REG_13__SCAN_IN), 
        .B2(n5658), .ZN(n5655) );
  OAI21_X1 U6681 ( .B1(n6562), .B2(n5661), .A(n5655), .ZN(U2952) );
  AOI22_X1 U6682 ( .A1(n5659), .A2(DATAI_14_), .B1(LWORD_REG_14__SCAN_IN), 
        .B2(n5658), .ZN(n5656) );
  OAI21_X1 U6683 ( .B1(n5657), .B2(n5661), .A(n5656), .ZN(U2953) );
  AOI22_X1 U6684 ( .A1(n5659), .A2(DATAI_15_), .B1(LWORD_REG_15__SCAN_IN), 
        .B2(n5658), .ZN(n5660) );
  OAI21_X1 U6685 ( .B1(n6729), .B2(n5661), .A(n5660), .ZN(U2954) );
  AOI22_X1 U6686 ( .A1(n5348), .A2(REIP_REG_2__SCAN_IN), .B1(n5662), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5671) );
  INV_X1 U6687 ( .A(n5663), .ZN(n5665) );
  NAND2_X1 U6688 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  XNOR2_X1 U6689 ( .A(n5667), .B(n5666), .ZN(n5747) );
  AOI22_X1 U6690 ( .A1(n5747), .A2(n5679), .B1(n5669), .B2(n5668), .ZN(n5670)
         );
  OAI211_X1 U6691 ( .C1(n5673), .C2(n5672), .A(n5671), .B(n5670), .ZN(U2984)
         );
  AOI21_X1 U6692 ( .B1(n5675), .B2(n6679), .A(n5674), .ZN(n5763) );
  NAND2_X1 U6693 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  AOI22_X1 U6694 ( .A1(n5679), .A2(n5763), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5678), .ZN(n5681) );
  NAND2_X1 U6695 ( .A1(n5348), .A2(REIP_REG_0__SCAN_IN), .ZN(n5680) );
  OAI211_X1 U6696 ( .C1(n5683), .C2(n5682), .A(n5681), .B(n5680), .ZN(U2986)
         );
  INV_X1 U6697 ( .A(n5684), .ZN(n5689) );
  OAI22_X1 U6698 ( .A1(n5771), .A2(n5685), .B1(n5740), .B2(n6345), .ZN(n5686)
         );
  AOI21_X1 U6699 ( .B1(n5764), .B2(n5687), .A(n5686), .ZN(n5688) );
  OAI221_X1 U6700 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5690), .C1(
        n6579), .C2(n5689), .A(n5688), .ZN(U3007) );
  AOI22_X1 U6701 ( .A1(n5754), .A2(n5691), .B1(n5348), .B2(REIP_REG_9__SCAN_IN), .ZN(n5695) );
  AOI22_X1 U6702 ( .A1(n5693), .A2(n5764), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n5692), .ZN(n5694) );
  OAI211_X1 U6703 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n5696), .A(n5695), 
        .B(n5694), .ZN(U3009) );
  NOR2_X1 U6704 ( .A1(n5740), .A2(n4564), .ZN(n5700) );
  OAI22_X1 U6705 ( .A1(n5698), .A2(n5733), .B1(n5705), .B2(n5697), .ZN(n5699)
         );
  AOI211_X1 U6706 ( .C1(n5754), .C2(n5701), .A(n5700), .B(n5699), .ZN(n5704)
         );
  OAI211_X1 U6707 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5708), .B(n5702), .ZN(n5703) );
  NAND2_X1 U6708 ( .A1(n5704), .A2(n5703), .ZN(U3010) );
  OAI22_X1 U6709 ( .A1(n5706), .A2(n5733), .B1(n5705), .B2(n6517), .ZN(n5707)
         );
  AOI21_X1 U6710 ( .B1(n5708), .B2(n6517), .A(n5707), .ZN(n5711) );
  INV_X1 U6711 ( .A(n5709), .ZN(n5710) );
  OAI211_X1 U6712 ( .C1(n5771), .C2(n5712), .A(n5711), .B(n5710), .ZN(U3011)
         );
  NOR2_X1 U6713 ( .A1(n5740), .A2(n4509), .ZN(n5716) );
  OAI22_X1 U6714 ( .A1(n5714), .A2(n5733), .B1(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .B2(n5713), .ZN(n5715) );
  AOI211_X1 U6715 ( .C1(n5754), .C2(n5717), .A(n5716), .B(n5715), .ZN(n5718)
         );
  OAI21_X1 U6716 ( .B1(n5720), .B2(n5719), .A(n5718), .ZN(U3012) );
  AOI21_X1 U6717 ( .B1(n5721), .B2(n5723), .A(n5748), .ZN(n5739) );
  INV_X1 U6718 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6501) );
  NOR2_X1 U6719 ( .A1(n5740), .A2(n6501), .ZN(n5728) );
  OAI21_X1 U6720 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5722), .ZN(n5725) );
  INV_X1 U6721 ( .A(n5723), .ZN(n5743) );
  NAND2_X1 U6722 ( .A1(n5724), .A2(n5743), .ZN(n5732) );
  OAI22_X1 U6723 ( .A1(n5726), .A2(n5733), .B1(n5725), .B2(n5732), .ZN(n5727)
         );
  AOI211_X1 U6724 ( .C1(n5754), .C2(n5729), .A(n5728), .B(n5727), .ZN(n5730)
         );
  OAI21_X1 U6725 ( .B1(n5739), .B2(n5731), .A(n5730), .ZN(U3014) );
  INV_X1 U6726 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6655) );
  OAI22_X1 U6727 ( .A1(n5734), .A2(n5733), .B1(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n5732), .ZN(n5735) );
  AOI211_X1 U6728 ( .C1(n5754), .C2(n5737), .A(n5736), .B(n5735), .ZN(n5738)
         );
  OAI21_X1 U6729 ( .B1(n5739), .B2(n6655), .A(n5738), .ZN(U3015) );
  NAND2_X1 U6730 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n3089), .ZN(n5751)
         );
  NOR2_X1 U6731 ( .A1(n5740), .A2(n6333), .ZN(n5745) );
  AOI221_X1 U6732 ( .B1(n3089), .B2(n5743), .C1(n5742), .C2(n5743), .A(n5741), 
        .ZN(n5744) );
  AOI211_X1 U6733 ( .C1(n5754), .C2(n5746), .A(n5745), .B(n5744), .ZN(n5750)
         );
  AOI22_X1 U6734 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n5748), .B1(n5764), 
        .B2(n5747), .ZN(n5749) );
  OAI211_X1 U6735 ( .C1(n5752), .C2(n5751), .A(n5750), .B(n5749), .ZN(U3016)
         );
  AOI22_X1 U6736 ( .A1(n5754), .A2(n5753), .B1(n5348), .B2(REIP_REG_1__SCAN_IN), .ZN(n5762) );
  INV_X1 U6737 ( .A(n5755), .ZN(n5756) );
  AOI22_X1 U6738 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5767), .B1(n5764), 
        .B2(n5756), .ZN(n5761) );
  NAND3_X1 U6739 ( .A1(n5759), .A2(n5758), .A3(n5757), .ZN(n5760) );
  NAND3_X1 U6740 ( .A1(n5762), .A2(n5761), .A3(n5760), .ZN(U3017) );
  AOI22_X1 U6741 ( .A1(n5764), .A2(n5763), .B1(n5348), .B2(REIP_REG_0__SCAN_IN), .ZN(n5770) );
  INV_X1 U6742 ( .A(n5765), .ZN(n5766) );
  OAI22_X1 U6743 ( .A1(n5768), .A2(n5767), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5766), .ZN(n5769) );
  OAI211_X1 U6744 ( .C1(n5772), .C2(n5771), .A(n5770), .B(n5769), .ZN(U3018)
         );
  NOR2_X1 U6745 ( .A1(n6630), .A2(n6403), .ZN(U3019) );
  NAND3_X1 U6746 ( .A1(n6734), .A2(n6405), .A3(n6667), .ZN(n5811) );
  NOR2_X1 U6747 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5811), .ZN(n5798)
         );
  AND2_X1 U6748 ( .A1(n4239), .A2(n5774), .ZN(n5987) );
  INV_X1 U6749 ( .A(n5987), .ZN(n5959) );
  INV_X1 U6750 ( .A(n5775), .ZN(n5776) );
  INV_X1 U6751 ( .A(n6170), .ZN(n5958) );
  OAI22_X1 U6752 ( .A1(n6087), .A2(n5959), .B1(n5776), .B2(n5958), .ZN(n5797)
         );
  AOI22_X1 U6753 ( .A1(n6197), .A2(n5798), .B1(n6196), .B2(n5797), .ZN(n5784)
         );
  NAND2_X1 U6754 ( .A1(n5803), .A2(n5777), .ZN(n5828) );
  AOI21_X1 U6755 ( .B1(n5828), .B2(n6258), .A(n6164), .ZN(n5782) );
  NAND2_X1 U6756 ( .A1(n5924), .A2(n5987), .ZN(n5806) );
  NAND2_X1 U6757 ( .A1(n5806), .A2(n6432), .ZN(n5781) );
  INV_X1 U6758 ( .A(n5798), .ZN(n5779) );
  AOI211_X1 U6759 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5779), .A(n6161), .B(
        n5778), .ZN(n5780) );
  AOI22_X1 U6760 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n5799), .B1(n6122), 
        .B2(n5830), .ZN(n5783) );
  OAI211_X1 U6761 ( .C1(n6125), .C2(n6258), .A(n5784), .B(n5783), .ZN(U3020)
         );
  AOI22_X1 U6762 ( .A1(n6214), .A2(n5798), .B1(n6213), .B2(n5797), .ZN(n5786)
         );
  AOI22_X1 U6763 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n5799), .B1(n6126), 
        .B2(n5830), .ZN(n5785) );
  OAI211_X1 U6764 ( .C1(n6129), .C2(n6258), .A(n5786), .B(n5785), .ZN(U3021)
         );
  INV_X1 U6765 ( .A(n6221), .ZN(n6133) );
  AOI22_X1 U6766 ( .A1(n6219), .A2(n5797), .B1(n6220), .B2(n5798), .ZN(n5788)
         );
  AOI22_X1 U6767 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n5799), .B1(n6130), 
        .B2(n5830), .ZN(n5787) );
  OAI211_X1 U6768 ( .C1(n6133), .C2(n6258), .A(n5788), .B(n5787), .ZN(U3022)
         );
  INV_X1 U6769 ( .A(n6227), .ZN(n6137) );
  AOI22_X1 U6770 ( .A1(n6226), .A2(n5798), .B1(n6225), .B2(n5797), .ZN(n5790)
         );
  AOI22_X1 U6771 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n5799), .B1(n6134), 
        .B2(n5830), .ZN(n5789) );
  OAI211_X1 U6772 ( .C1(n6137), .C2(n6258), .A(n5790), .B(n5789), .ZN(U3023)
         );
  AOI22_X1 U6773 ( .A1(n6232), .A2(n5798), .B1(n6231), .B2(n5797), .ZN(n5792)
         );
  AOI22_X1 U6774 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n5799), .B1(n6138), 
        .B2(n5830), .ZN(n5791) );
  OAI211_X1 U6775 ( .C1(n6141), .C2(n6258), .A(n5792), .B(n5791), .ZN(U3024)
         );
  AOI22_X1 U6776 ( .A1(n6238), .A2(n5798), .B1(n6237), .B2(n5797), .ZN(n5794)
         );
  AOI22_X1 U6777 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n5799), .B1(n6142), 
        .B2(n5830), .ZN(n5793) );
  OAI211_X1 U6778 ( .C1(n6145), .C2(n6258), .A(n5794), .B(n5793), .ZN(U3025)
         );
  AOI22_X1 U6779 ( .A1(n6244), .A2(n5798), .B1(n6243), .B2(n5797), .ZN(n5796)
         );
  AOI22_X1 U6780 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n5799), .B1(n6146), 
        .B2(n5830), .ZN(n5795) );
  OAI211_X1 U6781 ( .C1(n6149), .C2(n6258), .A(n5796), .B(n5795), .ZN(U3026)
         );
  INV_X1 U6782 ( .A(n6254), .ZN(n6157) );
  AOI22_X1 U6783 ( .A1(n6251), .A2(n5798), .B1(n6250), .B2(n5797), .ZN(n5801)
         );
  AOI22_X1 U6784 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n5799), .B1(n6152), 
        .B2(n5830), .ZN(n5800) );
  OAI211_X1 U6785 ( .C1(n6157), .C2(n6258), .A(n5801), .B(n5800), .ZN(U3027)
         );
  NOR2_X1 U6786 ( .A1(n6113), .A2(n5811), .ZN(n5829) );
  AOI22_X1 U6787 ( .A1(n6209), .A2(n5830), .B1(n6197), .B2(n5829), .ZN(n5815)
         );
  OAI21_X1 U6788 ( .B1(n5804), .B2(n6164), .A(n6432), .ZN(n5813) );
  OR2_X1 U6789 ( .A1(n5806), .A2(n5805), .ZN(n5808) );
  INV_X1 U6790 ( .A(n5829), .ZN(n5807) );
  AND2_X1 U6791 ( .A1(n5808), .A2(n5807), .ZN(n5812) );
  INV_X1 U6792 ( .A(n5812), .ZN(n5810) );
  AOI21_X1 U6793 ( .B1(n6203), .B2(n5811), .A(n6202), .ZN(n5809) );
  OAI21_X1 U6794 ( .B1(n5813), .B2(n5810), .A(n5809), .ZN(n5832) );
  OAI22_X1 U6795 ( .A1(n5813), .A2(n5812), .B1(n6550), .B2(n5811), .ZN(n5831)
         );
  AOI22_X1 U6796 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5832), .B1(n6196), 
        .B2(n5831), .ZN(n5814) );
  OAI211_X1 U6797 ( .C1(n5862), .C2(n6212), .A(n5815), .B(n5814), .ZN(U3028)
         );
  AOI22_X1 U6798 ( .A1(n6214), .A2(n5829), .B1(n5830), .B2(n6215), .ZN(n5817)
         );
  AOI22_X1 U6799 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5832), .B1(n6213), 
        .B2(n5831), .ZN(n5816) );
  OAI211_X1 U6800 ( .C1(n5862), .C2(n6218), .A(n5817), .B(n5816), .ZN(U3029)
         );
  INV_X1 U6801 ( .A(n5862), .ZN(n5838) );
  AOI22_X1 U6802 ( .A1(n5838), .A2(n6130), .B1(n6220), .B2(n5829), .ZN(n5819)
         );
  AOI22_X1 U6803 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5832), .B1(n6219), 
        .B2(n5831), .ZN(n5818) );
  OAI211_X1 U6804 ( .C1(n6133), .C2(n5828), .A(n5819), .B(n5818), .ZN(U3030)
         );
  AOI22_X1 U6805 ( .A1(n5838), .A2(n6134), .B1(n6226), .B2(n5829), .ZN(n5821)
         );
  AOI22_X1 U6806 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5832), .B1(n6225), 
        .B2(n5831), .ZN(n5820) );
  OAI211_X1 U6807 ( .C1(n6137), .C2(n5828), .A(n5821), .B(n5820), .ZN(U3031)
         );
  AOI22_X1 U6808 ( .A1(n6233), .A2(n5830), .B1(n6232), .B2(n5829), .ZN(n5823)
         );
  AOI22_X1 U6809 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5832), .B1(n6231), 
        .B2(n5831), .ZN(n5822) );
  OAI211_X1 U6810 ( .C1(n5862), .C2(n6236), .A(n5823), .B(n5822), .ZN(U3032)
         );
  AOI22_X1 U6811 ( .A1(n6238), .A2(n5829), .B1(n5830), .B2(n6239), .ZN(n5825)
         );
  AOI22_X1 U6812 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5832), .B1(n6237), 
        .B2(n5831), .ZN(n5824) );
  OAI211_X1 U6813 ( .C1(n5862), .C2(n6242), .A(n5825), .B(n5824), .ZN(U3033)
         );
  AOI22_X1 U6814 ( .A1(n6244), .A2(n5829), .B1(n5838), .B2(n6146), .ZN(n5827)
         );
  AOI22_X1 U6815 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5832), .B1(n6243), 
        .B2(n5831), .ZN(n5826) );
  OAI211_X1 U6816 ( .C1(n6149), .C2(n5828), .A(n5827), .B(n5826), .ZN(U3034)
         );
  INV_X1 U6817 ( .A(n6152), .ZN(n6259) );
  AOI22_X1 U6818 ( .A1(n6254), .A2(n5830), .B1(n6251), .B2(n5829), .ZN(n5834)
         );
  AOI22_X1 U6819 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5832), .B1(n6250), 
        .B2(n5831), .ZN(n5833) );
  OAI211_X1 U6820 ( .C1(n5862), .C2(n6259), .A(n5834), .B(n5833), .ZN(U3035)
         );
  NOR2_X1 U6821 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5835), .ZN(n5858)
         );
  INV_X1 U6822 ( .A(n5836), .ZN(n5839) );
  NAND3_X1 U6823 ( .A1(n6170), .A2(n6160), .A3(n6734), .ZN(n5837) );
  OAI21_X1 U6824 ( .B1(n5839), .B2(n6203), .A(n5837), .ZN(n5857) );
  AOI22_X1 U6825 ( .A1(n5858), .A2(n6197), .B1(n6196), .B2(n5857), .ZN(n5844)
         );
  OAI21_X1 U6826 ( .B1(n5838), .B2(n5873), .A(n6199), .ZN(n5840) );
  AOI21_X1 U6827 ( .B1(n5840), .B2(n5839), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5842) );
  OAI21_X1 U6828 ( .B1(n6160), .B2(n6550), .A(n5841), .ZN(n6168) );
  NOR2_X1 U6829 ( .A1(n6161), .A2(n6168), .ZN(n6021) );
  AOI22_X1 U6830 ( .A1(n5859), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6122), 
        .B2(n5873), .ZN(n5843) );
  OAI211_X1 U6831 ( .C1(n6125), .C2(n5862), .A(n5844), .B(n5843), .ZN(U3036)
         );
  AOI22_X1 U6832 ( .A1(n6214), .A2(n5858), .B1(n6213), .B2(n5857), .ZN(n5846)
         );
  AOI22_X1 U6833 ( .A1(n5859), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6126), 
        .B2(n5873), .ZN(n5845) );
  OAI211_X1 U6834 ( .C1(n5862), .C2(n6129), .A(n5846), .B(n5845), .ZN(U3037)
         );
  AOI22_X1 U6835 ( .A1(n5858), .A2(n6220), .B1(n6219), .B2(n5857), .ZN(n5848)
         );
  AOI22_X1 U6836 ( .A1(n5859), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6130), 
        .B2(n5873), .ZN(n5847) );
  OAI211_X1 U6837 ( .C1(n5862), .C2(n6133), .A(n5848), .B(n5847), .ZN(U3038)
         );
  AOI22_X1 U6838 ( .A1(n5858), .A2(n6226), .B1(n6225), .B2(n5857), .ZN(n5850)
         );
  AOI22_X1 U6839 ( .A1(n5859), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6134), 
        .B2(n5873), .ZN(n5849) );
  OAI211_X1 U6840 ( .C1(n5862), .C2(n6137), .A(n5850), .B(n5849), .ZN(U3039)
         );
  AOI22_X1 U6841 ( .A1(n5858), .A2(n6232), .B1(n6231), .B2(n5857), .ZN(n5852)
         );
  AOI22_X1 U6842 ( .A1(n5859), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6138), 
        .B2(n5873), .ZN(n5851) );
  OAI211_X1 U6843 ( .C1(n5862), .C2(n6141), .A(n5852), .B(n5851), .ZN(U3040)
         );
  AOI22_X1 U6844 ( .A1(n6238), .A2(n5858), .B1(n6237), .B2(n5857), .ZN(n5854)
         );
  AOI22_X1 U6845 ( .A1(n5859), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6142), 
        .B2(n5873), .ZN(n5853) );
  OAI211_X1 U6846 ( .C1(n5862), .C2(n6145), .A(n5854), .B(n5853), .ZN(U3041)
         );
  AOI22_X1 U6847 ( .A1(n6244), .A2(n5858), .B1(n6243), .B2(n5857), .ZN(n5856)
         );
  AOI22_X1 U6848 ( .A1(n5859), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6146), 
        .B2(n5873), .ZN(n5855) );
  OAI211_X1 U6849 ( .C1(n5862), .C2(n6149), .A(n5856), .B(n5855), .ZN(U3042)
         );
  AOI22_X1 U6850 ( .A1(n5858), .A2(n6251), .B1(n6250), .B2(n5857), .ZN(n5861)
         );
  AOI22_X1 U6851 ( .A1(n5859), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6152), 
        .B2(n5873), .ZN(n5860) );
  OAI211_X1 U6852 ( .C1(n5862), .C2(n6157), .A(n5861), .B(n5860), .ZN(U3043)
         );
  AOI22_X1 U6853 ( .A1(n6214), .A2(n5874), .B1(n6215), .B2(n5873), .ZN(n5864)
         );
  AOI22_X1 U6854 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n5876), .B1(n6213), 
        .B2(n5875), .ZN(n5863) );
  OAI211_X1 U6855 ( .C1(n6218), .C2(n5884), .A(n5864), .B(n5863), .ZN(U3045)
         );
  INV_X1 U6856 ( .A(n6130), .ZN(n6224) );
  AOI22_X1 U6857 ( .A1(n6220), .A2(n5874), .B1(n6221), .B2(n5873), .ZN(n5866)
         );
  AOI22_X1 U6858 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5876), .B1(n6219), 
        .B2(n5875), .ZN(n5865) );
  OAI211_X1 U6859 ( .C1(n6224), .C2(n5884), .A(n5866), .B(n5865), .ZN(U3046)
         );
  AOI22_X1 U6860 ( .A1(n6232), .A2(n5874), .B1(n6233), .B2(n5873), .ZN(n5868)
         );
  AOI22_X1 U6861 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5876), .B1(n6231), 
        .B2(n5875), .ZN(n5867) );
  OAI211_X1 U6862 ( .C1(n6236), .C2(n5884), .A(n5868), .B(n5867), .ZN(U3048)
         );
  AOI22_X1 U6863 ( .A1(n6238), .A2(n5874), .B1(n6239), .B2(n5873), .ZN(n5870)
         );
  AOI22_X1 U6864 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n5876), .B1(n6237), 
        .B2(n5875), .ZN(n5869) );
  OAI211_X1 U6865 ( .C1(n6242), .C2(n5884), .A(n5870), .B(n5869), .ZN(U3049)
         );
  AOI22_X1 U6866 ( .A1(n6244), .A2(n5874), .B1(n6245), .B2(n5873), .ZN(n5872)
         );
  AOI22_X1 U6867 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5876), .B1(n6243), 
        .B2(n5875), .ZN(n5871) );
  OAI211_X1 U6868 ( .C1(n6248), .C2(n5884), .A(n5872), .B(n5871), .ZN(U3050)
         );
  AOI22_X1 U6869 ( .A1(n6251), .A2(n5874), .B1(n6254), .B2(n5873), .ZN(n5878)
         );
  AOI22_X1 U6870 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5876), .B1(n6250), 
        .B2(n5875), .ZN(n5877) );
  OAI211_X1 U6871 ( .C1(n6259), .C2(n5884), .A(n5878), .B(n5877), .ZN(U3051)
         );
  AOI22_X1 U6872 ( .A1(n6226), .A2(n5880), .B1(n6225), .B2(n5879), .ZN(n5883)
         );
  AOI22_X1 U6873 ( .A1(n5881), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6134), 
        .B2(n5889), .ZN(n5882) );
  OAI211_X1 U6874 ( .C1(n6137), .C2(n5884), .A(n5883), .B(n5882), .ZN(U3055)
         );
  AOI22_X1 U6875 ( .A1(n6220), .A2(n5890), .B1(n5889), .B2(n6221), .ZN(n5886)
         );
  AOI22_X1 U6876 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5892), .B1(n6219), 
        .B2(n5891), .ZN(n5885) );
  OAI211_X1 U6877 ( .C1(n6224), .C2(n5898), .A(n5886), .B(n5885), .ZN(U3062)
         );
  INV_X1 U6878 ( .A(n6134), .ZN(n6230) );
  AOI22_X1 U6879 ( .A1(n6226), .A2(n5890), .B1(n5889), .B2(n6227), .ZN(n5888)
         );
  AOI22_X1 U6880 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5892), .B1(n6225), 
        .B2(n5891), .ZN(n5887) );
  OAI211_X1 U6881 ( .C1(n6230), .C2(n5898), .A(n5888), .B(n5887), .ZN(U3063)
         );
  AOI22_X1 U6882 ( .A1(n6251), .A2(n5890), .B1(n5889), .B2(n6254), .ZN(n5894)
         );
  AOI22_X1 U6883 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5892), .B1(n6250), 
        .B2(n5891), .ZN(n5893) );
  OAI211_X1 U6884 ( .C1(n6259), .C2(n5898), .A(n5894), .B(n5893), .ZN(U3067)
         );
  INV_X1 U6885 ( .A(n6158), .ZN(n5895) );
  NOR2_X1 U6886 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5930), .ZN(n5917)
         );
  NAND2_X1 U6887 ( .A1(n6401), .A2(n5896), .ZN(n6193) );
  NAND3_X1 U6888 ( .A1(n6161), .A2(n6160), .A3(n6734), .ZN(n5897) );
  OAI21_X1 U6889 ( .B1(n6087), .B2(n6193), .A(n5897), .ZN(n5916) );
  AOI22_X1 U6890 ( .A1(n6197), .A2(n5917), .B1(n6196), .B2(n5916), .ZN(n5903)
         );
  AOI21_X1 U6891 ( .B1(n5898), .B2(n5947), .A(n6164), .ZN(n5901) );
  NAND2_X1 U6892 ( .A1(n6193), .A2(n6432), .ZN(n6167) );
  INV_X1 U6893 ( .A(n5917), .ZN(n5899) );
  AOI211_X1 U6894 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5899), .A(n6170), .B(
        n6168), .ZN(n5900) );
  OAI211_X1 U6895 ( .C1(n5901), .C2(n6167), .A(n5900), .B(n6734), .ZN(n5919)
         );
  AOI22_X1 U6896 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n5919), .B1(n6209), 
        .B2(n5918), .ZN(n5902) );
  OAI211_X1 U6897 ( .C1(n6212), .C2(n5947), .A(n5903), .B(n5902), .ZN(U3068)
         );
  AOI22_X1 U6898 ( .A1(n6214), .A2(n5917), .B1(n6213), .B2(n5916), .ZN(n5905)
         );
  AOI22_X1 U6899 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n5919), .B1(n6215), 
        .B2(n5918), .ZN(n5904) );
  OAI211_X1 U6900 ( .C1(n6218), .C2(n5947), .A(n5905), .B(n5904), .ZN(U3069)
         );
  AOI22_X1 U6901 ( .A1(n6219), .A2(n5916), .B1(n6220), .B2(n5917), .ZN(n5907)
         );
  AOI22_X1 U6902 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n5919), .B1(n6221), 
        .B2(n5918), .ZN(n5906) );
  OAI211_X1 U6903 ( .C1(n6224), .C2(n5947), .A(n5907), .B(n5906), .ZN(U3070)
         );
  AOI22_X1 U6904 ( .A1(n6226), .A2(n5917), .B1(n6225), .B2(n5916), .ZN(n5909)
         );
  AOI22_X1 U6905 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n5919), .B1(n6227), 
        .B2(n5918), .ZN(n5908) );
  OAI211_X1 U6906 ( .C1(n6230), .C2(n5947), .A(n5909), .B(n5908), .ZN(U3071)
         );
  AOI22_X1 U6907 ( .A1(n6232), .A2(n5917), .B1(n6231), .B2(n5916), .ZN(n5911)
         );
  AOI22_X1 U6908 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n5919), .B1(n6233), 
        .B2(n5918), .ZN(n5910) );
  OAI211_X1 U6909 ( .C1(n6236), .C2(n5947), .A(n5911), .B(n5910), .ZN(U3072)
         );
  AOI22_X1 U6910 ( .A1(n6238), .A2(n5917), .B1(n6237), .B2(n5916), .ZN(n5913)
         );
  AOI22_X1 U6911 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n5919), .B1(n6239), 
        .B2(n5918), .ZN(n5912) );
  OAI211_X1 U6912 ( .C1(n6242), .C2(n5947), .A(n5913), .B(n5912), .ZN(U3073)
         );
  AOI22_X1 U6913 ( .A1(n6244), .A2(n5917), .B1(n6243), .B2(n5916), .ZN(n5915)
         );
  AOI22_X1 U6914 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n5919), .B1(n6245), 
        .B2(n5918), .ZN(n5914) );
  OAI211_X1 U6915 ( .C1(n6248), .C2(n5947), .A(n5915), .B(n5914), .ZN(U3074)
         );
  AOI22_X1 U6916 ( .A1(n6251), .A2(n5917), .B1(n6250), .B2(n5916), .ZN(n5921)
         );
  AOI22_X1 U6917 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n5919), .B1(n6254), 
        .B2(n5918), .ZN(n5920) );
  OAI211_X1 U6918 ( .C1(n6259), .C2(n5947), .A(n5921), .B(n5920), .ZN(U3075)
         );
  AOI22_X1 U6919 ( .A1(n5949), .A2(n6197), .B1(n6122), .B2(n5982), .ZN(n5934)
         );
  NAND2_X1 U6920 ( .A1(n6432), .A2(n5923), .ZN(n5931) );
  INV_X1 U6921 ( .A(n6193), .ZN(n5925) );
  NAND3_X1 U6922 ( .A1(n5925), .A2(n5924), .A3(n6263), .ZN(n5927) );
  INV_X1 U6923 ( .A(n5949), .ZN(n5926) );
  AND2_X1 U6924 ( .A1(n5927), .A2(n5926), .ZN(n5932) );
  INV_X1 U6925 ( .A(n5932), .ZN(n5929) );
  AOI21_X1 U6926 ( .B1(n5930), .B2(n6203), .A(n6202), .ZN(n5928) );
  OAI21_X1 U6927 ( .B1(n5931), .B2(n5929), .A(n5928), .ZN(n5951) );
  OAI22_X1 U6928 ( .A1(n5932), .A2(n5931), .B1(n6550), .B2(n5930), .ZN(n5950)
         );
  AOI22_X1 U6929 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5951), .B1(n6196), 
        .B2(n5950), .ZN(n5933) );
  OAI211_X1 U6930 ( .C1(n6125), .C2(n5947), .A(n5934), .B(n5933), .ZN(U3076)
         );
  AOI22_X1 U6931 ( .A1(n6214), .A2(n5949), .B1(n6215), .B2(n5948), .ZN(n5936)
         );
  AOI22_X1 U6932 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5951), .B1(n6213), 
        .B2(n5950), .ZN(n5935) );
  OAI211_X1 U6933 ( .C1(n6218), .C2(n5973), .A(n5936), .B(n5935), .ZN(U3077)
         );
  AOI22_X1 U6934 ( .A1(n5949), .A2(n6220), .B1(n6130), .B2(n5982), .ZN(n5938)
         );
  AOI22_X1 U6935 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5951), .B1(n6219), 
        .B2(n5950), .ZN(n5937) );
  OAI211_X1 U6936 ( .C1(n6133), .C2(n5947), .A(n5938), .B(n5937), .ZN(U3078)
         );
  AOI22_X1 U6937 ( .A1(n5949), .A2(n6226), .B1(n6134), .B2(n5982), .ZN(n5940)
         );
  AOI22_X1 U6938 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5951), .B1(n6225), 
        .B2(n5950), .ZN(n5939) );
  OAI211_X1 U6939 ( .C1(n6137), .C2(n5947), .A(n5940), .B(n5939), .ZN(U3079)
         );
  AOI22_X1 U6940 ( .A1(n5949), .A2(n6232), .B1(n6233), .B2(n5948), .ZN(n5942)
         );
  AOI22_X1 U6941 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5951), .B1(n6231), 
        .B2(n5950), .ZN(n5941) );
  OAI211_X1 U6942 ( .C1(n6236), .C2(n5973), .A(n5942), .B(n5941), .ZN(U3080)
         );
  AOI22_X1 U6943 ( .A1(n6238), .A2(n5949), .B1(n6142), .B2(n5982), .ZN(n5944)
         );
  AOI22_X1 U6944 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5951), .B1(n6237), 
        .B2(n5950), .ZN(n5943) );
  OAI211_X1 U6945 ( .C1(n6145), .C2(n5947), .A(n5944), .B(n5943), .ZN(U3081)
         );
  AOI22_X1 U6946 ( .A1(n6244), .A2(n5949), .B1(n6146), .B2(n5982), .ZN(n5946)
         );
  AOI22_X1 U6947 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5951), .B1(n6243), 
        .B2(n5950), .ZN(n5945) );
  OAI211_X1 U6948 ( .C1(n6149), .C2(n5947), .A(n5946), .B(n5945), .ZN(U3082)
         );
  AOI22_X1 U6949 ( .A1(n5949), .A2(n6251), .B1(n6254), .B2(n5948), .ZN(n5953)
         );
  AOI22_X1 U6950 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5951), .B1(n6250), 
        .B2(n5950), .ZN(n5952) );
  OAI211_X1 U6951 ( .C1(n6259), .C2(n5973), .A(n5953), .B(n5952), .ZN(U3083)
         );
  NAND3_X1 U6952 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6405), .A3(n6667), .ZN(n5990) );
  NOR2_X1 U6953 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5990), .ZN(n5981)
         );
  NAND2_X1 U6954 ( .A1(n6017), .A2(n6432), .ZN(n6163) );
  INV_X1 U6955 ( .A(n5955), .ZN(n5957) );
  NAND2_X1 U6956 ( .A1(n5957), .A2(n5956), .ZN(n6083) );
  OAI22_X1 U6957 ( .A1(n5959), .A2(n6163), .B1(n5958), .B2(n6083), .ZN(n5980)
         );
  AOI22_X1 U6958 ( .A1(n6197), .A2(n5981), .B1(n6196), .B2(n5980), .ZN(n5966)
         );
  OAI21_X1 U6959 ( .B1(n5987), .B2(n6203), .A(n6087), .ZN(n5960) );
  NAND3_X1 U6960 ( .A1(n5973), .A2(n6004), .A3(n5960), .ZN(n5964) );
  INV_X1 U6961 ( .A(n6161), .ZN(n6084) );
  AOI21_X1 U6962 ( .B1(n6083), .B2(STATE2_REG_2__SCAN_IN), .A(n5961), .ZN(
        n6090) );
  OAI211_X1 U6963 ( .C1(n6384), .C2(n5981), .A(n6084), .B(n6090), .ZN(n5962)
         );
  INV_X1 U6964 ( .A(n5962), .ZN(n5963) );
  OAI211_X1 U6965 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6087), .A(n5964), .B(
        n5963), .ZN(n5983) );
  AOI22_X1 U6966 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n5983), .B1(n6209), 
        .B2(n5982), .ZN(n5965) );
  OAI211_X1 U6967 ( .C1(n6212), .C2(n6004), .A(n5966), .B(n5965), .ZN(U3084)
         );
  AOI22_X1 U6968 ( .A1(n6214), .A2(n5981), .B1(n6213), .B2(n5980), .ZN(n5968)
         );
  AOI22_X1 U6969 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n5983), .B1(n6215), 
        .B2(n5982), .ZN(n5967) );
  OAI211_X1 U6970 ( .C1(n6218), .C2(n6004), .A(n5968), .B(n5967), .ZN(U3085)
         );
  AOI22_X1 U6971 ( .A1(n6219), .A2(n5980), .B1(n6220), .B2(n5981), .ZN(n5970)
         );
  AOI22_X1 U6972 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n5983), .B1(n6221), 
        .B2(n5982), .ZN(n5969) );
  OAI211_X1 U6973 ( .C1(n6224), .C2(n6004), .A(n5970), .B(n5969), .ZN(U3086)
         );
  AOI22_X1 U6974 ( .A1(n6226), .A2(n5981), .B1(n6225), .B2(n5980), .ZN(n5972)
         );
  INV_X1 U6975 ( .A(n6004), .ZN(n6010) );
  AOI22_X1 U6976 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(n5983), .B1(n6134), 
        .B2(n6010), .ZN(n5971) );
  OAI211_X1 U6977 ( .C1(n6137), .C2(n5973), .A(n5972), .B(n5971), .ZN(U3087)
         );
  AOI22_X1 U6978 ( .A1(n6232), .A2(n5981), .B1(n6231), .B2(n5980), .ZN(n5975)
         );
  AOI22_X1 U6979 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n5983), .B1(n6233), 
        .B2(n5982), .ZN(n5974) );
  OAI211_X1 U6980 ( .C1(n6236), .C2(n6004), .A(n5975), .B(n5974), .ZN(U3088)
         );
  AOI22_X1 U6981 ( .A1(n6238), .A2(n5981), .B1(n6237), .B2(n5980), .ZN(n5977)
         );
  AOI22_X1 U6982 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n5983), .B1(n6239), 
        .B2(n5982), .ZN(n5976) );
  OAI211_X1 U6983 ( .C1(n6242), .C2(n6004), .A(n5977), .B(n5976), .ZN(U3089)
         );
  AOI22_X1 U6984 ( .A1(n6244), .A2(n5981), .B1(n6243), .B2(n5980), .ZN(n5979)
         );
  AOI22_X1 U6985 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n5983), .B1(n6245), 
        .B2(n5982), .ZN(n5978) );
  OAI211_X1 U6986 ( .C1(n6248), .C2(n6004), .A(n5979), .B(n5978), .ZN(U3090)
         );
  AOI22_X1 U6987 ( .A1(n6251), .A2(n5981), .B1(n6250), .B2(n5980), .ZN(n5985)
         );
  AOI22_X1 U6988 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n5983), .B1(n6254), 
        .B2(n5982), .ZN(n5984) );
  OAI211_X1 U6989 ( .C1(n6259), .C2(n6004), .A(n5985), .B(n5984), .ZN(U3091)
         );
  INV_X1 U6990 ( .A(n6045), .ZN(n6001) );
  NOR2_X1 U6991 ( .A1(n6113), .A2(n5990), .ZN(n6009) );
  AOI22_X1 U6992 ( .A1(n6122), .A2(n6001), .B1(n6197), .B2(n6009), .ZN(n5994)
         );
  OAI21_X1 U6993 ( .B1(n6049), .B2(n5986), .A(n6432), .ZN(n5991) );
  NAND2_X1 U6994 ( .A1(n6017), .A2(n6263), .ZN(n6194) );
  INV_X1 U6995 ( .A(n6194), .ZN(n6115) );
  AOI21_X1 U6996 ( .B1(n6115), .B2(n5987), .A(n6009), .ZN(n5992) );
  INV_X1 U6997 ( .A(n5992), .ZN(n5989) );
  AOI21_X1 U6998 ( .B1(n6203), .B2(n5990), .A(n6202), .ZN(n5988) );
  OAI21_X1 U6999 ( .B1(n5991), .B2(n5989), .A(n5988), .ZN(n6012) );
  OAI22_X1 U7000 ( .A1(n5992), .A2(n5991), .B1(n6550), .B2(n5990), .ZN(n6011)
         );
  AOI22_X1 U7001 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6012), .B1(n6196), 
        .B2(n6011), .ZN(n5993) );
  OAI211_X1 U7002 ( .C1(n6125), .C2(n6004), .A(n5994), .B(n5993), .ZN(U3092)
         );
  AOI22_X1 U7003 ( .A1(n6214), .A2(n6009), .B1(n6126), .B2(n6001), .ZN(n5996)
         );
  AOI22_X1 U7004 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6012), .B1(n6213), 
        .B2(n6011), .ZN(n5995) );
  OAI211_X1 U7005 ( .C1(n6129), .C2(n6004), .A(n5996), .B(n5995), .ZN(U3093)
         );
  AOI22_X1 U7006 ( .A1(n6130), .A2(n6001), .B1(n6220), .B2(n6009), .ZN(n5998)
         );
  AOI22_X1 U7007 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6012), .B1(n6219), 
        .B2(n6011), .ZN(n5997) );
  OAI211_X1 U7008 ( .C1(n6133), .C2(n6004), .A(n5998), .B(n5997), .ZN(U3094)
         );
  AOI22_X1 U7009 ( .A1(n6134), .A2(n6001), .B1(n6226), .B2(n6009), .ZN(n6000)
         );
  AOI22_X1 U7010 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6012), .B1(n6225), 
        .B2(n6011), .ZN(n5999) );
  OAI211_X1 U7011 ( .C1(n6137), .C2(n6004), .A(n6000), .B(n5999), .ZN(U3095)
         );
  AOI22_X1 U7012 ( .A1(n6138), .A2(n6001), .B1(n6232), .B2(n6009), .ZN(n6003)
         );
  AOI22_X1 U7013 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6012), .B1(n6231), 
        .B2(n6011), .ZN(n6002) );
  OAI211_X1 U7014 ( .C1(n6141), .C2(n6004), .A(n6003), .B(n6002), .ZN(U3096)
         );
  AOI22_X1 U7015 ( .A1(n6238), .A2(n6009), .B1(n6239), .B2(n6010), .ZN(n6006)
         );
  AOI22_X1 U7016 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6012), .B1(n6237), 
        .B2(n6011), .ZN(n6005) );
  OAI211_X1 U7017 ( .C1(n6242), .C2(n6045), .A(n6006), .B(n6005), .ZN(U3097)
         );
  AOI22_X1 U7018 ( .A1(n6244), .A2(n6009), .B1(n6245), .B2(n6010), .ZN(n6008)
         );
  AOI22_X1 U7019 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6012), .B1(n6243), 
        .B2(n6011), .ZN(n6007) );
  OAI211_X1 U7020 ( .C1(n6248), .C2(n6045), .A(n6008), .B(n6007), .ZN(U3098)
         );
  AOI22_X1 U7021 ( .A1(n6254), .A2(n6010), .B1(n6251), .B2(n6009), .ZN(n6014)
         );
  AOI22_X1 U7022 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6012), .B1(n6250), 
        .B2(n6011), .ZN(n6013) );
  OAI211_X1 U7023 ( .C1(n6259), .C2(n6045), .A(n6014), .B(n6013), .ZN(U3099)
         );
  NAND3_X1 U7024 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6405), .ZN(n6057) );
  NOR2_X1 U7025 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6057), .ZN(n6040)
         );
  AOI22_X1 U7026 ( .A1(n6122), .A2(n6062), .B1(n6197), .B2(n6040), .ZN(n6027)
         );
  NAND2_X1 U7027 ( .A1(n6081), .A2(n6045), .ZN(n6015) );
  AOI21_X1 U7028 ( .B1(n6015), .B2(STATEBS16_REG_SCAN_IN), .A(n6203), .ZN(
        n6022) );
  INV_X1 U7029 ( .A(n6016), .ZN(n6018) );
  INV_X1 U7030 ( .A(n6052), .ZN(n6024) );
  INV_X1 U7031 ( .A(n6040), .ZN(n6019) );
  AOI22_X1 U7032 ( .A1(n6022), .A2(n6024), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n6019), .ZN(n6020) );
  OAI211_X1 U7033 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6550), .A(n6021), .B(n6020), .ZN(n6042) );
  INV_X1 U7034 ( .A(n6022), .ZN(n6025) );
  NAND3_X1 U7035 ( .A1(n6170), .A2(n6160), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6023) );
  AOI22_X1 U7036 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n6042), .B1(n6196), 
        .B2(n6041), .ZN(n6026) );
  OAI211_X1 U7037 ( .C1(n6125), .C2(n6045), .A(n6027), .B(n6026), .ZN(U3100)
         );
  AOI22_X1 U7038 ( .A1(n6214), .A2(n6040), .B1(n6126), .B2(n6062), .ZN(n6029)
         );
  AOI22_X1 U7039 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n6042), .B1(n6213), 
        .B2(n6041), .ZN(n6028) );
  OAI211_X1 U7040 ( .C1(n6129), .C2(n6045), .A(n6029), .B(n6028), .ZN(U3101)
         );
  AOI22_X1 U7041 ( .A1(n6130), .A2(n6062), .B1(n6220), .B2(n6040), .ZN(n6031)
         );
  AOI22_X1 U7042 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n6042), .B1(n6219), 
        .B2(n6041), .ZN(n6030) );
  OAI211_X1 U7043 ( .C1(n6133), .C2(n6045), .A(n6031), .B(n6030), .ZN(U3102)
         );
  AOI22_X1 U7044 ( .A1(n6134), .A2(n6062), .B1(n6226), .B2(n6040), .ZN(n6033)
         );
  AOI22_X1 U7045 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n6042), .B1(n6225), 
        .B2(n6041), .ZN(n6032) );
  OAI211_X1 U7046 ( .C1(n6137), .C2(n6045), .A(n6033), .B(n6032), .ZN(U3103)
         );
  AOI22_X1 U7047 ( .A1(n6138), .A2(n6062), .B1(n6232), .B2(n6040), .ZN(n6035)
         );
  AOI22_X1 U7048 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n6042), .B1(n6231), 
        .B2(n6041), .ZN(n6034) );
  OAI211_X1 U7049 ( .C1(n6141), .C2(n6045), .A(n6035), .B(n6034), .ZN(U3104)
         );
  AOI22_X1 U7050 ( .A1(n6238), .A2(n6040), .B1(n6142), .B2(n6062), .ZN(n6037)
         );
  AOI22_X1 U7051 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n6042), .B1(n6237), 
        .B2(n6041), .ZN(n6036) );
  OAI211_X1 U7052 ( .C1(n6145), .C2(n6045), .A(n6037), .B(n6036), .ZN(U3105)
         );
  AOI22_X1 U7053 ( .A1(n6244), .A2(n6040), .B1(n6146), .B2(n6062), .ZN(n6039)
         );
  AOI22_X1 U7054 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n6042), .B1(n6243), 
        .B2(n6041), .ZN(n6038) );
  OAI211_X1 U7055 ( .C1(n6149), .C2(n6045), .A(n6039), .B(n6038), .ZN(U3106)
         );
  AOI22_X1 U7056 ( .A1(n6152), .A2(n6062), .B1(n6251), .B2(n6040), .ZN(n6044)
         );
  AOI22_X1 U7057 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n6042), .B1(n6250), 
        .B2(n6041), .ZN(n6043) );
  OAI211_X1 U7058 ( .C1(n6157), .C2(n6045), .A(n6044), .B(n6043), .ZN(U3107)
         );
  INV_X1 U7059 ( .A(n6046), .ZN(n6047) );
  NOR2_X1 U7060 ( .A1(n6048), .A2(n6734), .ZN(n6076) );
  AOI22_X1 U7061 ( .A1(n6122), .A2(n6109), .B1(n6197), .B2(n6076), .ZN(n6061)
         );
  INV_X1 U7062 ( .A(n6057), .ZN(n6055) );
  INV_X1 U7063 ( .A(n6202), .ZN(n6054) );
  INV_X1 U7064 ( .A(n6049), .ZN(n6051) );
  AOI21_X1 U7065 ( .B1(n6051), .B2(n6050), .A(n6203), .ZN(n6056) );
  AOI21_X1 U7066 ( .B1(n6052), .B2(n6263), .A(n6076), .ZN(n6058) );
  NAND2_X1 U7067 ( .A1(n6056), .A2(n6058), .ZN(n6053) );
  OAI211_X1 U7068 ( .C1(n6432), .C2(n6055), .A(n6054), .B(n6053), .ZN(n6078)
         );
  INV_X1 U7069 ( .A(n6056), .ZN(n6059) );
  OAI22_X1 U7070 ( .A1(n6059), .A2(n6058), .B1(n6057), .B2(n6550), .ZN(n6077)
         );
  AOI22_X1 U7071 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6078), .B1(n6196), 
        .B2(n6077), .ZN(n6060) );
  OAI211_X1 U7072 ( .C1(n6125), .C2(n6081), .A(n6061), .B(n6060), .ZN(U3108)
         );
  AOI22_X1 U7073 ( .A1(n6214), .A2(n6076), .B1(n6215), .B2(n6062), .ZN(n6064)
         );
  AOI22_X1 U7074 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6078), .B1(n6213), 
        .B2(n6077), .ZN(n6063) );
  OAI211_X1 U7075 ( .C1(n6218), .C2(n6065), .A(n6064), .B(n6063), .ZN(U3109)
         );
  AOI22_X1 U7076 ( .A1(n6130), .A2(n6109), .B1(n6220), .B2(n6076), .ZN(n6067)
         );
  AOI22_X1 U7077 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6078), .B1(n6219), 
        .B2(n6077), .ZN(n6066) );
  OAI211_X1 U7078 ( .C1(n6133), .C2(n6081), .A(n6067), .B(n6066), .ZN(U3110)
         );
  AOI22_X1 U7079 ( .A1(n6134), .A2(n6109), .B1(n6226), .B2(n6076), .ZN(n6069)
         );
  AOI22_X1 U7080 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6078), .B1(n6225), 
        .B2(n6077), .ZN(n6068) );
  OAI211_X1 U7081 ( .C1(n6137), .C2(n6081), .A(n6069), .B(n6068), .ZN(U3111)
         );
  AOI22_X1 U7082 ( .A1(n6138), .A2(n6109), .B1(n6232), .B2(n6076), .ZN(n6071)
         );
  AOI22_X1 U7083 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6078), .B1(n6231), 
        .B2(n6077), .ZN(n6070) );
  OAI211_X1 U7084 ( .C1(n6141), .C2(n6081), .A(n6071), .B(n6070), .ZN(U3112)
         );
  AOI22_X1 U7085 ( .A1(n6238), .A2(n6076), .B1(n6142), .B2(n6109), .ZN(n6073)
         );
  AOI22_X1 U7086 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6078), .B1(n6237), 
        .B2(n6077), .ZN(n6072) );
  OAI211_X1 U7087 ( .C1(n6145), .C2(n6081), .A(n6073), .B(n6072), .ZN(U3113)
         );
  AOI22_X1 U7088 ( .A1(n6244), .A2(n6076), .B1(n6146), .B2(n6109), .ZN(n6075)
         );
  AOI22_X1 U7089 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6078), .B1(n6243), 
        .B2(n6077), .ZN(n6074) );
  OAI211_X1 U7090 ( .C1(n6149), .C2(n6081), .A(n6075), .B(n6074), .ZN(U3114)
         );
  AOI22_X1 U7091 ( .A1(n6152), .A2(n6109), .B1(n6251), .B2(n6076), .ZN(n6080)
         );
  AOI22_X1 U7092 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6078), .B1(n6250), 
        .B2(n6077), .ZN(n6079) );
  OAI211_X1 U7093 ( .C1(n6157), .C2(n6081), .A(n6080), .B(n6079), .ZN(U3115)
         );
  NAND3_X1 U7094 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6667), .ZN(n6119) );
  NOR2_X1 U7095 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6119), .ZN(n6108)
         );
  INV_X1 U7096 ( .A(n6114), .ZN(n6085) );
  OAI22_X1 U7097 ( .A1(n6085), .A2(n6163), .B1(n6084), .B2(n6083), .ZN(n6107)
         );
  AOI22_X1 U7098 ( .A1(n6197), .A2(n6108), .B1(n6196), .B2(n6107), .ZN(n6094)
         );
  INV_X1 U7099 ( .A(n6156), .ZN(n6086) );
  OAI21_X1 U7100 ( .B1(n6109), .B2(n6086), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6089) );
  OAI21_X1 U7101 ( .B1(n6114), .B2(n6203), .A(n6087), .ZN(n6088) );
  NAND2_X1 U7102 ( .A1(n6089), .A2(n6088), .ZN(n6091) );
  OAI211_X1 U7103 ( .C1(n6108), .C2(n6384), .A(n6091), .B(n6090), .ZN(n6092)
         );
  AOI22_X1 U7104 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n6110), .B1(n6209), 
        .B2(n6109), .ZN(n6093) );
  OAI211_X1 U7105 ( .C1(n6212), .C2(n6156), .A(n6094), .B(n6093), .ZN(U3116)
         );
  AOI22_X1 U7106 ( .A1(n6214), .A2(n6108), .B1(n6213), .B2(n6107), .ZN(n6096)
         );
  AOI22_X1 U7107 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n6110), .B1(n6215), 
        .B2(n6109), .ZN(n6095) );
  OAI211_X1 U7108 ( .C1(n6218), .C2(n6156), .A(n6096), .B(n6095), .ZN(U3117)
         );
  AOI22_X1 U7109 ( .A1(n6219), .A2(n6107), .B1(n6220), .B2(n6108), .ZN(n6098)
         );
  AOI22_X1 U7110 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n6110), .B1(n6221), 
        .B2(n6109), .ZN(n6097) );
  OAI211_X1 U7111 ( .C1(n6224), .C2(n6156), .A(n6098), .B(n6097), .ZN(U3118)
         );
  AOI22_X1 U7112 ( .A1(n6226), .A2(n6108), .B1(n6225), .B2(n6107), .ZN(n6100)
         );
  AOI22_X1 U7113 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(n6110), .B1(n6227), 
        .B2(n6109), .ZN(n6099) );
  OAI211_X1 U7114 ( .C1(n6230), .C2(n6156), .A(n6100), .B(n6099), .ZN(U3119)
         );
  AOI22_X1 U7115 ( .A1(n6232), .A2(n6108), .B1(n6231), .B2(n6107), .ZN(n6102)
         );
  AOI22_X1 U7116 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n6110), .B1(n6233), 
        .B2(n6109), .ZN(n6101) );
  OAI211_X1 U7117 ( .C1(n6236), .C2(n6156), .A(n6102), .B(n6101), .ZN(U3120)
         );
  AOI22_X1 U7118 ( .A1(n6238), .A2(n6108), .B1(n6237), .B2(n6107), .ZN(n6104)
         );
  AOI22_X1 U7119 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n6110), .B1(n6239), 
        .B2(n6109), .ZN(n6103) );
  OAI211_X1 U7120 ( .C1(n6242), .C2(n6156), .A(n6104), .B(n6103), .ZN(U3121)
         );
  AOI22_X1 U7121 ( .A1(n6244), .A2(n6108), .B1(n6243), .B2(n6107), .ZN(n6106)
         );
  AOI22_X1 U7122 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(n6110), .B1(n6245), 
        .B2(n6109), .ZN(n6105) );
  OAI211_X1 U7123 ( .C1(n6248), .C2(n6156), .A(n6106), .B(n6105), .ZN(U3122)
         );
  AOI22_X1 U7124 ( .A1(n6251), .A2(n6108), .B1(n6250), .B2(n6107), .ZN(n6112)
         );
  AOI22_X1 U7125 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n6110), .B1(n6254), 
        .B2(n6109), .ZN(n6111) );
  OAI211_X1 U7126 ( .C1(n6259), .C2(n6156), .A(n6112), .B(n6111), .ZN(U3123)
         );
  NOR2_X1 U7127 ( .A1(n6113), .A2(n6119), .ZN(n6151) );
  AOI21_X1 U7128 ( .B1(n6115), .B2(n6114), .A(n6151), .ZN(n6117) );
  OAI22_X1 U7129 ( .A1(n6117), .A2(n6203), .B1(n6119), .B2(n6550), .ZN(n6150)
         );
  AOI22_X1 U7130 ( .A1(n6197), .A2(n6151), .B1(n6196), .B2(n6150), .ZN(n6124)
         );
  AND2_X1 U7131 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  AOI221_X1 U7132 ( .B1(n6203), .B2(n6119), .C1(n6432), .C2(n6118), .A(n6202), 
        .ZN(n6120) );
  AOI22_X1 U7133 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6153), .B1(n6122), 
        .B2(n6188), .ZN(n6123) );
  OAI211_X1 U7134 ( .C1(n6125), .C2(n6156), .A(n6124), .B(n6123), .ZN(U3124)
         );
  AOI22_X1 U7135 ( .A1(n6214), .A2(n6151), .B1(n6213), .B2(n6150), .ZN(n6128)
         );
  AOI22_X1 U7136 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6153), .B1(n6126), 
        .B2(n6188), .ZN(n6127) );
  OAI211_X1 U7137 ( .C1(n6129), .C2(n6156), .A(n6128), .B(n6127), .ZN(U3125)
         );
  AOI22_X1 U7138 ( .A1(n6219), .A2(n6150), .B1(n6220), .B2(n6151), .ZN(n6132)
         );
  AOI22_X1 U7139 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6153), .B1(n6130), 
        .B2(n6188), .ZN(n6131) );
  OAI211_X1 U7140 ( .C1(n6133), .C2(n6156), .A(n6132), .B(n6131), .ZN(U3126)
         );
  AOI22_X1 U7141 ( .A1(n6226), .A2(n6151), .B1(n6225), .B2(n6150), .ZN(n6136)
         );
  AOI22_X1 U7142 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6153), .B1(n6134), 
        .B2(n6188), .ZN(n6135) );
  OAI211_X1 U7143 ( .C1(n6137), .C2(n6156), .A(n6136), .B(n6135), .ZN(U3127)
         );
  AOI22_X1 U7144 ( .A1(n6232), .A2(n6151), .B1(n6231), .B2(n6150), .ZN(n6140)
         );
  AOI22_X1 U7145 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6153), .B1(n6138), 
        .B2(n6188), .ZN(n6139) );
  OAI211_X1 U7146 ( .C1(n6141), .C2(n6156), .A(n6140), .B(n6139), .ZN(U3128)
         );
  AOI22_X1 U7147 ( .A1(n6238), .A2(n6151), .B1(n6237), .B2(n6150), .ZN(n6144)
         );
  AOI22_X1 U7148 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6153), .B1(n6142), 
        .B2(n6188), .ZN(n6143) );
  OAI211_X1 U7149 ( .C1(n6145), .C2(n6156), .A(n6144), .B(n6143), .ZN(U3129)
         );
  AOI22_X1 U7150 ( .A1(n6244), .A2(n6151), .B1(n6243), .B2(n6150), .ZN(n6148)
         );
  AOI22_X1 U7151 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6153), .B1(n6146), 
        .B2(n6188), .ZN(n6147) );
  OAI211_X1 U7152 ( .C1(n6149), .C2(n6156), .A(n6148), .B(n6147), .ZN(U3130)
         );
  AOI22_X1 U7153 ( .A1(n6251), .A2(n6151), .B1(n6250), .B2(n6150), .ZN(n6155)
         );
  AOI22_X1 U7154 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6153), .B1(n6152), 
        .B2(n6188), .ZN(n6154) );
  OAI211_X1 U7155 ( .C1(n6157), .C2(n6156), .A(n6155), .B(n6154), .ZN(U3131)
         );
  NOR2_X1 U7156 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6204), .ZN(n6187)
         );
  NAND3_X1 U7157 ( .A1(n6161), .A2(n6160), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6162) );
  OAI21_X1 U7158 ( .B1(n6163), .B2(n6193), .A(n6162), .ZN(n6186) );
  AOI22_X1 U7159 ( .A1(n6197), .A2(n6187), .B1(n6196), .B2(n6186), .ZN(n6173)
         );
  AOI21_X1 U7160 ( .B1(n6165), .B2(n6208), .A(n6164), .ZN(n6166) );
  NOR2_X1 U7161 ( .A1(n6167), .A2(n6166), .ZN(n6169) );
  NOR4_X1 U7162 ( .A1(n6734), .A2(n6170), .A3(n6169), .A4(n6168), .ZN(n6171)
         );
  AOI22_X1 U7163 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6189), .B1(n6209), 
        .B2(n6188), .ZN(n6172) );
  OAI211_X1 U7164 ( .C1(n6212), .C2(n6208), .A(n6173), .B(n6172), .ZN(U3132)
         );
  AOI22_X1 U7165 ( .A1(n6214), .A2(n6187), .B1(n6213), .B2(n6186), .ZN(n6175)
         );
  AOI22_X1 U7166 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6189), .B1(n6215), 
        .B2(n6188), .ZN(n6174) );
  OAI211_X1 U7167 ( .C1(n6218), .C2(n6208), .A(n6175), .B(n6174), .ZN(U3133)
         );
  AOI22_X1 U7168 ( .A1(n6219), .A2(n6186), .B1(n6220), .B2(n6187), .ZN(n6177)
         );
  AOI22_X1 U7169 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6189), .B1(n6221), 
        .B2(n6188), .ZN(n6176) );
  OAI211_X1 U7170 ( .C1(n6224), .C2(n6208), .A(n6177), .B(n6176), .ZN(U3134)
         );
  AOI22_X1 U7171 ( .A1(n6226), .A2(n6187), .B1(n6225), .B2(n6186), .ZN(n6179)
         );
  AOI22_X1 U7172 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6189), .B1(n6227), 
        .B2(n6188), .ZN(n6178) );
  OAI211_X1 U7173 ( .C1(n6230), .C2(n6208), .A(n6179), .B(n6178), .ZN(U3135)
         );
  AOI22_X1 U7174 ( .A1(n6232), .A2(n6187), .B1(n6231), .B2(n6186), .ZN(n6181)
         );
  AOI22_X1 U7175 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6189), .B1(n6233), 
        .B2(n6188), .ZN(n6180) );
  OAI211_X1 U7176 ( .C1(n6236), .C2(n6208), .A(n6181), .B(n6180), .ZN(U3136)
         );
  AOI22_X1 U7177 ( .A1(n6238), .A2(n6187), .B1(n6237), .B2(n6186), .ZN(n6183)
         );
  AOI22_X1 U7178 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6189), .B1(n6239), 
        .B2(n6188), .ZN(n6182) );
  OAI211_X1 U7179 ( .C1(n6242), .C2(n6208), .A(n6183), .B(n6182), .ZN(U3137)
         );
  AOI22_X1 U7180 ( .A1(n6244), .A2(n6187), .B1(n6243), .B2(n6186), .ZN(n6185)
         );
  AOI22_X1 U7181 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6189), .B1(n6245), 
        .B2(n6188), .ZN(n6184) );
  OAI211_X1 U7182 ( .C1(n6248), .C2(n6208), .A(n6185), .B(n6184), .ZN(U3138)
         );
  AOI22_X1 U7183 ( .A1(n6251), .A2(n6187), .B1(n6250), .B2(n6186), .ZN(n6191)
         );
  AOI22_X1 U7184 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6189), .B1(n6254), 
        .B2(n6188), .ZN(n6190) );
  OAI211_X1 U7185 ( .C1(n6259), .C2(n6208), .A(n6191), .B(n6190), .ZN(U3139)
         );
  OAI21_X1 U7186 ( .B1(n6194), .B2(n6193), .A(n6192), .ZN(n6206) );
  INV_X1 U7187 ( .A(n6206), .ZN(n6195) );
  OAI22_X1 U7188 ( .A1(n6195), .A2(n6203), .B1(n6204), .B2(n6550), .ZN(n6249)
         );
  AOI22_X1 U7189 ( .A1(n6252), .A2(n6197), .B1(n6196), .B2(n6249), .ZN(n6211)
         );
  AOI21_X1 U7190 ( .B1(n6198), .B2(n3096), .A(n5682), .ZN(n6201) );
  INV_X1 U7191 ( .A(n6199), .ZN(n6200) );
  NOR2_X1 U7192 ( .A1(n6201), .A2(n6200), .ZN(n6207) );
  AOI21_X1 U7193 ( .B1(n6204), .B2(n6203), .A(n6202), .ZN(n6205) );
  OAI21_X1 U7194 ( .B1(n6207), .B2(n6206), .A(n6205), .ZN(n6255) );
  AOI22_X1 U7195 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6255), .B1(n6209), 
        .B2(n6253), .ZN(n6210) );
  OAI211_X1 U7196 ( .C1(n6212), .C2(n6258), .A(n6211), .B(n6210), .ZN(U3140)
         );
  AOI22_X1 U7197 ( .A1(n6214), .A2(n6252), .B1(n6213), .B2(n6249), .ZN(n6217)
         );
  AOI22_X1 U7198 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6255), .B1(n6215), 
        .B2(n6253), .ZN(n6216) );
  OAI211_X1 U7199 ( .C1(n6218), .C2(n6258), .A(n6217), .B(n6216), .ZN(U3141)
         );
  AOI22_X1 U7200 ( .A1(n6252), .A2(n6220), .B1(n6219), .B2(n6249), .ZN(n6223)
         );
  AOI22_X1 U7201 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6255), .B1(n6221), 
        .B2(n6253), .ZN(n6222) );
  OAI211_X1 U7202 ( .C1(n6224), .C2(n6258), .A(n6223), .B(n6222), .ZN(U3142)
         );
  AOI22_X1 U7203 ( .A1(n6252), .A2(n6226), .B1(n6225), .B2(n6249), .ZN(n6229)
         );
  AOI22_X1 U7204 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6255), .B1(n6227), 
        .B2(n6253), .ZN(n6228) );
  OAI211_X1 U7205 ( .C1(n6230), .C2(n6258), .A(n6229), .B(n6228), .ZN(U3143)
         );
  AOI22_X1 U7206 ( .A1(n6252), .A2(n6232), .B1(n6231), .B2(n6249), .ZN(n6235)
         );
  AOI22_X1 U7207 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6255), .B1(n6233), 
        .B2(n6253), .ZN(n6234) );
  OAI211_X1 U7208 ( .C1(n6236), .C2(n6258), .A(n6235), .B(n6234), .ZN(U3144)
         );
  AOI22_X1 U7209 ( .A1(n6238), .A2(n6252), .B1(n6237), .B2(n6249), .ZN(n6241)
         );
  AOI22_X1 U7210 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6255), .B1(n6239), 
        .B2(n6253), .ZN(n6240) );
  OAI211_X1 U7211 ( .C1(n6242), .C2(n6258), .A(n6241), .B(n6240), .ZN(U3145)
         );
  AOI22_X1 U7212 ( .A1(n6244), .A2(n6252), .B1(n6243), .B2(n6249), .ZN(n6247)
         );
  AOI22_X1 U7213 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6255), .B1(n6245), 
        .B2(n6253), .ZN(n6246) );
  OAI211_X1 U7214 ( .C1(n6248), .C2(n6258), .A(n6247), .B(n6246), .ZN(U3146)
         );
  AOI22_X1 U7215 ( .A1(n6252), .A2(n6251), .B1(n6250), .B2(n6249), .ZN(n6257)
         );
  AOI22_X1 U7216 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6255), .B1(n6254), 
        .B2(n6253), .ZN(n6256) );
  OAI211_X1 U7217 ( .C1(n6259), .C2(n6258), .A(n6257), .B(n6256), .ZN(U3147)
         );
  AOI22_X1 U7218 ( .A1(n6263), .A2(n6262), .B1(n6261), .B2(n6260), .ZN(n6391)
         );
  NAND2_X1 U7219 ( .A1(n6264), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6397) );
  AND3_X1 U7220 ( .A1(n6391), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6397), 
        .ZN(n6268) );
  NAND2_X1 U7221 ( .A1(n6266), .A2(n6265), .ZN(n6267) );
  AOI222_X1 U7222 ( .A1(n6268), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n6268), .B2(n6267), .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6267), 
        .ZN(n6269) );
  AOI222_X1 U7223 ( .A1(n6405), .A2(n6270), .B1(n6405), .B2(n6269), .C1(n6270), 
        .C2(n6269), .ZN(n6272) );
  OAI21_X1 U7224 ( .B1(n6272), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6271), 
        .ZN(n6290) );
  AOI21_X1 U7225 ( .B1(n6272), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6289) );
  OAI21_X1 U7226 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6273), 
        .ZN(n6285) );
  AND3_X1 U7227 ( .A1(n6284), .A2(n6275), .A3(n3091), .ZN(n6281) );
  NAND2_X1 U7228 ( .A1(n6277), .A2(n6276), .ZN(n6280) );
  NAND2_X1 U7229 ( .A1(n6282), .A2(n6278), .ZN(n6279) );
  OAI211_X1 U7230 ( .C1(n6282), .C2(n6281), .A(n6280), .B(n6279), .ZN(n6283)
         );
  INV_X1 U7231 ( .A(n6283), .ZN(n6417) );
  NAND4_X1 U7232 ( .A1(n6286), .A2(n6285), .A3(n6417), .A4(n6284), .ZN(n6287)
         );
  AOI211_X1 U7233 ( .C1(n6290), .C2(n6289), .A(n6288), .B(n6287), .ZN(n6302)
         );
  NAND2_X1 U7234 ( .A1(n6292), .A2(n6291), .ZN(n6297) );
  AOI22_X1 U7235 ( .A1(n6293), .A2(n6302), .B1(READY_N), .B2(n6421), .ZN(n6294) );
  INV_X1 U7236 ( .A(n6294), .ZN(n6295) );
  OAI21_X1 U7237 ( .B1(n6297), .B2(n6296), .A(n6295), .ZN(n6383) );
  OAI21_X1 U7238 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6420), .A(n6383), .ZN(
        n6304) );
  AOI221_X1 U7239 ( .B1(n6299), .B2(STATE2_REG_0__SCAN_IN), .C1(n6304), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6298), .ZN(n6301) );
  OAI211_X1 U7240 ( .C1(n6311), .C2(n6386), .A(n6303), .B(n6383), .ZN(n6300)
         );
  OAI211_X1 U7241 ( .C1(n6302), .C2(n6305), .A(n6301), .B(n6300), .ZN(U3148)
         );
  NAND2_X1 U7242 ( .A1(n6303), .A2(n6550), .ZN(n6313) );
  NAND3_X1 U7243 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6313), .A3(n6304), .ZN(
        n6310) );
  OAI21_X1 U7244 ( .B1(READY_N), .B2(n6306), .A(n6305), .ZN(n6308) );
  AOI21_X1 U7245 ( .B1(n6308), .B2(n6383), .A(n6307), .ZN(n6309) );
  NAND2_X1 U7246 ( .A1(n6310), .A2(n6309), .ZN(U3149) );
  INV_X1 U7247 ( .A(n6311), .ZN(n6424) );
  INV_X1 U7248 ( .A(n6312), .ZN(n6381) );
  OAI211_X1 U7249 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6420), .A(n6381), .B(
        n6313), .ZN(n6315) );
  OAI21_X1 U7250 ( .B1(n6424), .B2(n6315), .A(n6314), .ZN(U3150) );
  NOR2_X1 U7251 ( .A1(n6380), .A2(n6719), .ZN(U3151) );
  AND2_X1 U7252 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6750), .ZN(U3152) );
  INV_X1 U7253 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6697) );
  NOR2_X1 U7254 ( .A1(n6380), .A2(n6697), .ZN(U3154) );
  NOR2_X1 U7255 ( .A1(n6380), .A2(n6536), .ZN(U3155) );
  INV_X1 U7256 ( .A(DATAWIDTH_REG_26__SCAN_IN), .ZN(n6512) );
  NOR2_X1 U7257 ( .A1(n6380), .A2(n6512), .ZN(U3156) );
  AND2_X1 U7258 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6750), .ZN(U3157) );
  AND2_X1 U7259 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6750), .ZN(U3158) );
  NOR2_X1 U7260 ( .A1(n6380), .A2(n6632), .ZN(U3159) );
  INV_X1 U7261 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6600) );
  NOR2_X1 U7262 ( .A1(n6380), .A2(n6600), .ZN(U3160) );
  AND2_X1 U7263 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6750), .ZN(U3161) );
  AND2_X1 U7264 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6750), .ZN(U3162) );
  NOR2_X1 U7265 ( .A1(n6380), .A2(n6518), .ZN(U3163) );
  AND2_X1 U7266 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6750), .ZN(U3164) );
  AND2_X1 U7267 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6750), .ZN(U3165) );
  AND2_X1 U7268 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6750), .ZN(U3166) );
  AND2_X1 U7269 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6750), .ZN(U3167) );
  NOR2_X1 U7270 ( .A1(n6380), .A2(n6629), .ZN(U3168) );
  AND2_X1 U7271 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6750), .ZN(U3169) );
  AND2_X1 U7272 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6750), .ZN(U3170) );
  AND2_X1 U7273 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6750), .ZN(U3171) );
  NOR2_X1 U7274 ( .A1(n6380), .A2(n6553), .ZN(U3172) );
  AND2_X1 U7275 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6750), .ZN(U3173) );
  AND2_X1 U7276 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6750), .ZN(U3174) );
  AND2_X1 U7277 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6750), .ZN(U3175) );
  AND2_X1 U7278 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6750), .ZN(U3176) );
  AND2_X1 U7279 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6750), .ZN(U3177) );
  AND2_X1 U7280 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6750), .ZN(U3178) );
  AND2_X1 U7281 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6750), .ZN(U3179) );
  AND2_X1 U7282 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6750), .ZN(U3180) );
  AOI22_X1 U7283 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6331) );
  AND2_X1 U7284 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6319) );
  INV_X1 U7285 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6317) );
  INV_X1 U7286 ( .A(NA_N), .ZN(n6324) );
  AOI221_X1 U7287 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6324), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6328) );
  AOI221_X1 U7288 ( .B1(n6319), .B2(n6375), .C1(n6317), .C2(n6336), .A(n6328), 
        .ZN(n6316) );
  OAI21_X1 U7289 ( .B1(n6323), .B2(n6331), .A(n6316), .ZN(U3181) );
  NOR2_X1 U7290 ( .A1(n6326), .A2(n6317), .ZN(n6325) );
  NAND2_X1 U7291 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6318) );
  OAI21_X1 U7292 ( .B1(n6325), .B2(n6319), .A(n6318), .ZN(n6320) );
  OAI211_X1 U7293 ( .C1(n6322), .C2(n6420), .A(n6321), .B(n6320), .ZN(U3182)
         );
  AOI21_X1 U7294 ( .B1(n6325), .B2(n6324), .A(n6323), .ZN(n6330) );
  AOI221_X1 U7295 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6420), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6327) );
  AOI221_X1 U7296 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6327), .C2(HOLD), .A(n6326), .ZN(n6329) );
  OAI22_X1 U7297 ( .A1(n6331), .A2(n6330), .B1(n6329), .B2(n6328), .ZN(U3183)
         );
  NAND2_X1 U7298 ( .A1(n6429), .A2(n6617), .ZN(n6369) );
  INV_X1 U7299 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U7300 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6429), .ZN(n6373) );
  OAI222_X1 U7301 ( .A1(n6369), .A2(n6333), .B1(n6732), .B2(n6429), .C1(n6407), 
        .C2(n6373), .ZN(U3184) );
  INV_X1 U7302 ( .A(n6369), .ZN(n6371) );
  AOI22_X1 U7303 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6336), .ZN(n6332) );
  OAI21_X1 U7304 ( .B1(n6333), .B2(n6373), .A(n6332), .ZN(U3185) );
  AOI22_X1 U7305 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6336), .ZN(n6334) );
  OAI21_X1 U7306 ( .B1(n6335), .B2(n6373), .A(n6334), .ZN(U3186) );
  AOI22_X1 U7307 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6336), .ZN(n6337) );
  OAI21_X1 U7308 ( .B1(n6501), .B2(n6373), .A(n6337), .ZN(U3187) );
  AOI22_X1 U7309 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6375), .ZN(n6338) );
  OAI21_X1 U7310 ( .B1(n6339), .B2(n6373), .A(n6338), .ZN(U3188) );
  INV_X1 U7311 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6486) );
  OAI222_X1 U7312 ( .A1(n6373), .A2(n4509), .B1(n6486), .B2(n6429), .C1(n6340), 
        .C2(n6369), .ZN(U3189) );
  INV_X1 U7313 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6496) );
  OAI222_X1 U7314 ( .A1(n6373), .A2(n6340), .B1(n6496), .B2(n6429), .C1(n4564), 
        .C2(n6369), .ZN(U3190) );
  AOI22_X1 U7315 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6375), .ZN(n6341) );
  OAI21_X1 U7316 ( .B1(n4564), .B2(n6373), .A(n6341), .ZN(U3191) );
  AOI22_X1 U7317 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6375), .ZN(n6342) );
  OAI21_X1 U7318 ( .B1(n4521), .B2(n6373), .A(n6342), .ZN(U3192) );
  INV_X1 U7319 ( .A(n6373), .ZN(n6364) );
  AOI22_X1 U7320 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6364), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6375), .ZN(n6343) );
  OAI21_X1 U7321 ( .B1(n6345), .B2(n6369), .A(n6343), .ZN(U3193) );
  AOI22_X1 U7322 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6375), .ZN(n6344) );
  OAI21_X1 U7323 ( .B1(n6345), .B2(n6373), .A(n6344), .ZN(U3194) );
  AOI22_X1 U7324 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6364), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6375), .ZN(n6346) );
  OAI21_X1 U7325 ( .B1(n6348), .B2(n6369), .A(n6346), .ZN(U3195) );
  AOI22_X1 U7326 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6375), .ZN(n6347) );
  OAI21_X1 U7327 ( .B1(n6348), .B2(n6373), .A(n6347), .ZN(U3196) );
  INV_X1 U7328 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6482) );
  INV_X1 U7329 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6349) );
  OAI222_X1 U7330 ( .A1(n6369), .A2(n6593), .B1(n6482), .B2(n6429), .C1(n6349), 
        .C2(n6373), .ZN(U3197) );
  AOI22_X1 U7331 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6375), .ZN(n6350) );
  OAI21_X1 U7332 ( .B1(n6593), .B2(n6373), .A(n6350), .ZN(U3198) );
  AOI22_X1 U7333 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6375), .ZN(n6351) );
  OAI21_X1 U7334 ( .B1(n6352), .B2(n6373), .A(n6351), .ZN(U3199) );
  AOI22_X1 U7335 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6364), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6375), .ZN(n6353) );
  OAI21_X1 U7336 ( .B1(n6487), .B2(n6369), .A(n6353), .ZN(U3200) );
  AOI22_X1 U7337 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6375), .ZN(n6354) );
  OAI21_X1 U7338 ( .B1(n6487), .B2(n6373), .A(n6354), .ZN(U3201) );
  AOI22_X1 U7339 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6364), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6375), .ZN(n6355) );
  OAI21_X1 U7340 ( .B1(n6357), .B2(n6369), .A(n6355), .ZN(U3202) );
  AOI22_X1 U7341 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6375), .ZN(n6356) );
  OAI21_X1 U7342 ( .B1(n6357), .B2(n6373), .A(n6356), .ZN(U3203) );
  AOI22_X1 U7343 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6375), .ZN(n6358) );
  OAI21_X1 U7344 ( .B1(n6359), .B2(n6373), .A(n6358), .ZN(U3204) );
  AOI22_X1 U7345 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6364), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6375), .ZN(n6360) );
  OAI21_X1 U7346 ( .B1(n6361), .B2(n6369), .A(n6360), .ZN(U3205) );
  AOI22_X1 U7347 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6364), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6375), .ZN(n6362) );
  OAI21_X1 U7348 ( .B1(n6583), .B2(n6369), .A(n6362), .ZN(U3206) );
  AOI22_X1 U7349 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6364), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6375), .ZN(n6363) );
  OAI21_X1 U7350 ( .B1(n6504), .B2(n6369), .A(n6363), .ZN(U3207) );
  AOI22_X1 U7351 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6364), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6375), .ZN(n6365) );
  OAI21_X1 U7352 ( .B1(n6639), .B2(n6369), .A(n6365), .ZN(U3208) );
  INV_X1 U7353 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6495) );
  OAI222_X1 U7354 ( .A1(n6373), .A2(n6639), .B1(n6495), .B2(n6429), .C1(n6367), 
        .C2(n6369), .ZN(U3209) );
  AOI22_X1 U7355 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6375), .ZN(n6366) );
  OAI21_X1 U7356 ( .B1(n6367), .B2(n6373), .A(n6366), .ZN(U3210) );
  AOI22_X1 U7357 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6375), .ZN(n6368) );
  OAI21_X1 U7358 ( .B1(n5016), .B2(n6373), .A(n6368), .ZN(U3211) );
  INV_X1 U7359 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6695) );
  OAI222_X1 U7360 ( .A1(n6373), .A2(n6370), .B1(n6695), .B2(n6429), .C1(n6374), 
        .C2(n6369), .ZN(U3212) );
  AOI22_X1 U7361 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6371), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6375), .ZN(n6372) );
  OAI21_X1 U7362 ( .B1(n6374), .B2(n6373), .A(n6372), .ZN(U3213) );
  MUX2_X1 U7363 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6429), .Z(U3445) );
  MUX2_X1 U7364 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6429), .Z(U3446) );
  MUX2_X1 U7365 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6429), .Z(U3447) );
  INV_X1 U7366 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6413) );
  INV_X1 U7367 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6668) );
  AOI22_X1 U7368 ( .A1(n6429), .A2(n6413), .B1(n6668), .B2(n6375), .ZN(U3448)
         );
  INV_X1 U7369 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6377) );
  INV_X1 U7370 ( .A(n6378), .ZN(n6376) );
  AOI21_X1 U7371 ( .B1(n6750), .B2(n6377), .A(n6376), .ZN(U3451) );
  OAI21_X1 U7372 ( .B1(n6380), .B2(n6379), .A(n6378), .ZN(U3452) );
  OAI211_X1 U7373 ( .C1(n6384), .C2(n6383), .A(n6382), .B(n6381), .ZN(U3453)
         );
  INV_X1 U7374 ( .A(n6385), .ZN(n6388) );
  OAI22_X1 U7375 ( .A1(n6388), .A2(n6396), .B1(n6387), .B2(n6386), .ZN(n6390)
         );
  MUX2_X1 U7376 ( .A(n6390), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6389), 
        .Z(U3456) );
  OAI22_X1 U7377 ( .A1(n6391), .A2(n6396), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6431), .ZN(n6393) );
  OAI22_X1 U7378 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6394), .B1(n6393), .B2(n6392), .ZN(n6395) );
  OAI21_X1 U7379 ( .B1(n6397), .B2(n6396), .A(n6395), .ZN(U3461) );
  INV_X1 U7380 ( .A(n6403), .ZN(n6406) );
  XNOR2_X1 U7381 ( .A(n4263), .B(n6398), .ZN(n6402) );
  INV_X1 U7382 ( .A(n6399), .ZN(n6400) );
  AOI22_X1 U7383 ( .A1(n6402), .A2(n6432), .B1(n6401), .B2(n6400), .ZN(n6404)
         );
  AOI22_X1 U7384 ( .A1(n6406), .A2(n6405), .B1(n6404), .B2(n6403), .ZN(U3463)
         );
  AOI21_X1 U7385 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6408) );
  AOI22_X1 U7386 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6408), .B2(n6407), .ZN(n6411) );
  INV_X1 U7387 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6410) );
  AOI22_X1 U7388 ( .A1(n6414), .A2(n6411), .B1(n6410), .B2(n6409), .ZN(U3468)
         );
  OAI21_X1 U7389 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6414), .ZN(n6412) );
  OAI21_X1 U7390 ( .B1(n6414), .B2(n6413), .A(n6412), .ZN(U3469) );
  INV_X1 U7391 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6502) );
  MUX2_X1 U7392 ( .A(W_R_N_REG_SCAN_IN), .B(n6502), .S(n6429), .Z(U3470) );
  INV_X1 U7393 ( .A(MORE_REG_SCAN_IN), .ZN(n6416) );
  INV_X1 U7394 ( .A(n6418), .ZN(n6415) );
  AOI22_X1 U7395 ( .A1(n6418), .A2(n6417), .B1(n6416), .B2(n6415), .ZN(U3471)
         );
  AOI211_X1 U7396 ( .C1(n6421), .C2(n6420), .A(n6419), .B(n6434), .ZN(n6428)
         );
  OAI211_X1 U7397 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6423), .A(n6422), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6425) );
  AOI21_X1 U7398 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6425), .A(n6424), .ZN(
        n6427) );
  NAND2_X1 U7399 ( .A1(n6428), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6426) );
  OAI21_X1 U7400 ( .B1(n6428), .B2(n6427), .A(n6426), .ZN(U3472) );
  MUX2_X1 U7401 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6429), .Z(U3473) );
  AOI211_X1 U7402 ( .C1(n6432), .C2(n6431), .A(READREQUEST_REG_SCAN_IN), .B(
        n6430), .ZN(n6436) );
  AOI22_X1 U7403 ( .A1(n6436), .A2(n6435), .B1(n6434), .B2(n6433), .ZN(U3474)
         );
  NOR2_X1 U7404 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n6447) );
  NOR4_X1 U7405 ( .A1(EAX_REG_13__SCAN_IN), .A2(ADDRESS_REG_28__SCAN_IN), .A3(
        ADDRESS_REG_0__SCAN_IN), .A4(ADDRESS_REG_5__SCAN_IN), .ZN(n6445) );
  NOR4_X1 U7406 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6437) );
  NAND3_X1 U7407 ( .A1(n6437), .A2(n6734), .A3(n6679), .ZN(n6443) );
  NOR4_X1 U7408 ( .A1(UWORD_REG_5__SCAN_IN), .A2(UWORD_REG_0__SCAN_IN), .A3(
        LWORD_REG_14__SCAN_IN), .A4(DATAO_REG_13__SCAN_IN), .ZN(n6441) );
  NOR4_X1 U7409 ( .A1(DATAI_15_), .A2(DATAO_REG_10__SCAN_IN), .A3(
        LWORD_REG_3__SCAN_IN), .A4(DATAO_REG_1__SCAN_IN), .ZN(n6440) );
  NOR4_X1 U7410 ( .A1(EBX_REG_13__SCAN_IN), .A2(EAX_REG_18__SCAN_IN), .A3(
        DATAI_2_), .A4(DATAI_16_), .ZN(n6439) );
  NOR4_X1 U7411 ( .A1(EAX_REG_15__SCAN_IN), .A2(EAX_REG_16__SCAN_IN), .A3(
        DATAO_REG_29__SCAN_IN), .A4(DATAO_REG_24__SCAN_IN), .ZN(n6438) );
  NAND4_X1 U7412 ( .A1(n6441), .A2(n6440), .A3(n6439), .A4(n6438), .ZN(n6442)
         );
  NOR4_X1 U7413 ( .A1(STATE2_REG_2__SCAN_IN), .A2(EAX_REG_11__SCAN_IN), .A3(
        n6443), .A4(n6442), .ZN(n6444) );
  NAND4_X1 U7414 ( .A1(n6447), .A2(n6446), .A3(n6445), .A4(n6444), .ZN(n6479)
         );
  NOR4_X1 U7415 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(DATAI_11_), .A3(
        DATAI_6_), .A4(DATAI_21_), .ZN(n6451) );
  NOR4_X1 U7416 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(
        INSTQUEUE_REG_9__6__SCAN_IN), .A3(INSTQUEUE_REG_2__6__SCAN_IN), .A4(
        INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6450) );
  NOR4_X1 U7417 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .A3(REIP_REG_15__SCAN_IN), .A4(n6482), 
        .ZN(n6449) );
  NOR4_X1 U7418 ( .A1(EBX_REG_20__SCAN_IN), .A2(REIP_REG_31__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(DATAI_30_), .ZN(n6448) );
  NAND4_X1 U7419 ( .A1(n6451), .A2(n6450), .A3(n6449), .A4(n6448), .ZN(n6478)
         );
  NOR4_X1 U7420 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(INSTADDRPOINTER_REG_19__SCAN_IN), 
        .A4(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6455) );
  NOR4_X1 U7421 ( .A1(EBX_REG_23__SCAN_IN), .A2(EBX_REG_18__SCAN_IN), .A3(
        EBX_REG_16__SCAN_IN), .A4(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6454)
         );
  NOR4_X1 U7422 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(
        INSTQUEUE_REG_9__5__SCAN_IN), .A3(INSTQUEUE_REG_8__5__SCAN_IN), .A4(
        INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6453) );
  NOR4_X1 U7423 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(
        INSTQUEUE_REG_8__0__SCAN_IN), .A3(INSTQUEUE_REG_3__2__SCAN_IN), .A4(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6452) );
  NAND4_X1 U7424 ( .A1(n6455), .A2(n6454), .A3(n6453), .A4(n6452), .ZN(n6477)
         );
  NAND4_X1 U7425 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(DATAO_REG_27__SCAN_IN), .A3(UWORD_REG_7__SCAN_IN), .A4(DATAO_REG_18__SCAN_IN), .ZN(n6459) );
  NAND4_X1 U7426 ( .A1(EBX_REG_9__SCAN_IN), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), 
        .A3(DATAO_REG_23__SCAN_IN), .A4(DATAO_REG_11__SCAN_IN), .ZN(n6458) );
  NAND4_X1 U7427 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(
        INSTQUEUE_REG_7__2__SCAN_IN), .A3(PHYADDRPOINTER_REG_21__SCAN_IN), 
        .A4(REIP_REG_17__SCAN_IN), .ZN(n6457) );
  NAND4_X1 U7428 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(
        INSTQUEUE_REG_3__0__SCAN_IN), .A3(REIP_REG_12__SCAN_IN), .A4(
        REIP_REG_4__SCAN_IN), .ZN(n6456) );
  NOR4_X1 U7429 ( .A1(n6459), .A2(n6458), .A3(n6457), .A4(n6456), .ZN(n6475)
         );
  NAND4_X1 U7430 ( .A1(READREQUEST_REG_SCAN_IN), .A2(DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6463)
         );
  NAND4_X1 U7431 ( .A1(ADDRESS_REG_25__SCAN_IN), .A2(ADDRESS_REG_6__SCAN_IN), 
        .A3(BE_N_REG_0__SCAN_IN), .A4(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6462)
         );
  NAND4_X1 U7432 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .A4(EAX_REG_9__SCAN_IN), .ZN(n6461) );
  NAND4_X1 U7433 ( .A1(STATE_REG_2__SCAN_IN), .A2(EBX_REG_3__SCAN_IN), .A3(
        DATAWIDTH_REG_23__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6460)
         );
  NOR4_X1 U7434 ( .A1(n6463), .A2(n6462), .A3(n6461), .A4(n6460), .ZN(n6474)
         );
  NAND4_X1 U7435 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(
        INSTQUEUE_REG_2__7__SCAN_IN), .A3(EAX_REG_27__SCAN_IN), .A4(DATAI_4_), 
        .ZN(n6467) );
  NAND4_X1 U7436 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(
        INSTQUEUE_REG_15__6__SCAN_IN), .A3(INSTQUEUE_REG_11__6__SCAN_IN), .A4(
        INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6466) );
  NAND4_X1 U7437 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_27__SCAN_IN), .A3(REIP_REG_24__SCAN_IN), .A4(
        DATAO_REG_31__SCAN_IN), .ZN(n6465) );
  NAND4_X1 U7438 ( .A1(EBX_REG_28__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .A3(EAX_REG_28__SCAN_IN), .A4(
        DATAI_24_), .ZN(n6464) );
  NOR4_X1 U7439 ( .A1(n6467), .A2(n6466), .A3(n6465), .A4(n6464), .ZN(n6473)
         );
  NAND4_X1 U7440 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(
        INSTQUEUE_REG_8__2__SCAN_IN), .A3(INSTQUEUE_REG_9__2__SCAN_IN), .A4(
        INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6471) );
  NAND4_X1 U7441 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(
        INSTQUEUE_REG_15__2__SCAN_IN), .A3(INSTQUEUE_REG_4__2__SCAN_IN), .A4(
        INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6470) );
  NAND4_X1 U7442 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        INSTQUEUE_REG_9__4__SCAN_IN), .A3(INSTQUEUE_REG_13__6__SCAN_IN), .A4(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6469) );
  NAND4_X1 U7443 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(
        INSTQUEUE_REG_12__1__SCAN_IN), .A3(INSTQUEUE_REG_13__3__SCAN_IN), .A4(
        INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6468) );
  NOR4_X1 U7444 ( .A1(n6471), .A2(n6470), .A3(n6469), .A4(n6468), .ZN(n6472)
         );
  NAND4_X1 U7445 ( .A1(n6475), .A2(n6474), .A3(n6473), .A4(n6472), .ZN(n6476)
         );
  NOR4_X1 U7446 ( .A1(n6479), .A2(n6478), .A3(n6477), .A4(n6476), .ZN(n6749)
         );
  AOI22_X1 U7447 ( .A1(n6482), .A2(keyinput101), .B1(n6481), .B2(keyinput99), 
        .ZN(n6480) );
  OAI221_X1 U7448 ( .B1(n6482), .B2(keyinput101), .C1(n6481), .C2(keyinput99), 
        .A(n6480), .ZN(n6493) );
  INV_X1 U7449 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6484) );
  AOI22_X1 U7450 ( .A1(n3934), .A2(keyinput64), .B1(keyinput39), .B2(n6484), 
        .ZN(n6483) );
  OAI221_X1 U7451 ( .B1(n3934), .B2(keyinput64), .C1(n6484), .C2(keyinput39), 
        .A(n6483), .ZN(n6492) );
  AOI22_X1 U7452 ( .A1(n6487), .A2(keyinput47), .B1(keyinput127), .B2(n6486), 
        .ZN(n6485) );
  OAI221_X1 U7453 ( .B1(n6487), .B2(keyinput47), .C1(n6486), .C2(keyinput127), 
        .A(n6485), .ZN(n6491) );
  INV_X1 U7454 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n6489) );
  AOI22_X1 U7455 ( .A1(n6489), .A2(keyinput57), .B1(n4487), .B2(keyinput120), 
        .ZN(n6488) );
  OAI221_X1 U7456 ( .B1(n6489), .B2(keyinput57), .C1(n4487), .C2(keyinput120), 
        .A(n6488), .ZN(n6490) );
  NOR4_X1 U7457 ( .A1(n6493), .A2(n6492), .A3(n6491), .A4(n6490), .ZN(n6545)
         );
  AOI22_X1 U7458 ( .A1(n6496), .A2(keyinput13), .B1(n6495), .B2(keyinput5), 
        .ZN(n6494) );
  OAI221_X1 U7459 ( .B1(n6496), .B2(keyinput13), .C1(n6495), .C2(keyinput5), 
        .A(n6494), .ZN(n6509) );
  INV_X1 U7460 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n6498) );
  AOI22_X1 U7461 ( .A1(n6499), .A2(keyinput44), .B1(keyinput119), .B2(n6498), 
        .ZN(n6497) );
  OAI221_X1 U7462 ( .B1(n6499), .B2(keyinput44), .C1(n6498), .C2(keyinput119), 
        .A(n6497), .ZN(n6508) );
  AOI22_X1 U7463 ( .A1(n6502), .A2(keyinput125), .B1(n6501), .B2(keyinput74), 
        .ZN(n6500) );
  OAI221_X1 U7464 ( .B1(n6502), .B2(keyinput125), .C1(n6501), .C2(keyinput74), 
        .A(n6500), .ZN(n6507) );
  AOI22_X1 U7465 ( .A1(n6505), .A2(keyinput92), .B1(keyinput88), .B2(n6504), 
        .ZN(n6503) );
  OAI221_X1 U7466 ( .B1(n6505), .B2(keyinput92), .C1(n6504), .C2(keyinput88), 
        .A(n6503), .ZN(n6506) );
  NOR4_X1 U7467 ( .A1(n6509), .A2(n6508), .A3(n6507), .A4(n6506), .ZN(n6544)
         );
  INV_X1 U7468 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6511) );
  AOI22_X1 U7469 ( .A1(n6512), .A2(keyinput53), .B1(n6511), .B2(keyinput87), 
        .ZN(n6510) );
  OAI221_X1 U7470 ( .B1(n6512), .B2(keyinput53), .C1(n6511), .C2(keyinput87), 
        .A(n6510), .ZN(n6525) );
  INV_X1 U7471 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6514) );
  AOI22_X1 U7472 ( .A1(n6515), .A2(keyinput108), .B1(n6514), .B2(keyinput60), 
        .ZN(n6513) );
  OAI221_X1 U7473 ( .B1(n6515), .B2(keyinput108), .C1(n6514), .C2(keyinput60), 
        .A(n6513), .ZN(n6524) );
  AOI22_X1 U7474 ( .A1(n6518), .A2(keyinput27), .B1(n6517), .B2(keyinput112), 
        .ZN(n6516) );
  OAI221_X1 U7475 ( .B1(n6518), .B2(keyinput27), .C1(n6517), .C2(keyinput112), 
        .A(n6516), .ZN(n6523) );
  INV_X1 U7476 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6521) );
  INV_X1 U7477 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6520) );
  AOI22_X1 U7478 ( .A1(n6521), .A2(keyinput100), .B1(keyinput114), .B2(n6520), 
        .ZN(n6519) );
  OAI221_X1 U7479 ( .B1(n6521), .B2(keyinput100), .C1(n6520), .C2(keyinput114), 
        .A(n6519), .ZN(n6522) );
  NOR4_X1 U7480 ( .A1(n6525), .A2(n6524), .A3(n6523), .A4(n6522), .ZN(n6543)
         );
  AOI22_X1 U7481 ( .A1(n6528), .A2(keyinput109), .B1(keyinput122), .B2(n6527), 
        .ZN(n6526) );
  OAI221_X1 U7482 ( .B1(n6528), .B2(keyinput109), .C1(n6527), .C2(keyinput122), 
        .A(n6526), .ZN(n6541) );
  INV_X1 U7483 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6531) );
  AOI22_X1 U7484 ( .A1(n6531), .A2(keyinput4), .B1(keyinput83), .B2(n6530), 
        .ZN(n6529) );
  OAI221_X1 U7485 ( .B1(n6531), .B2(keyinput4), .C1(n6530), .C2(keyinput83), 
        .A(n6529), .ZN(n6540) );
  INV_X1 U7486 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6534) );
  INV_X1 U7487 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6533) );
  AOI22_X1 U7488 ( .A1(n6534), .A2(keyinput50), .B1(n6533), .B2(keyinput116), 
        .ZN(n6532) );
  OAI221_X1 U7489 ( .B1(n6534), .B2(keyinput50), .C1(n6533), .C2(keyinput116), 
        .A(n6532), .ZN(n6539) );
  INV_X1 U7490 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6537) );
  AOI22_X1 U7491 ( .A1(n6537), .A2(keyinput80), .B1(keyinput56), .B2(n6536), 
        .ZN(n6535) );
  OAI221_X1 U7492 ( .B1(n6537), .B2(keyinput80), .C1(n6536), .C2(keyinput56), 
        .A(n6535), .ZN(n6538) );
  NOR4_X1 U7493 ( .A1(n6541), .A2(n6540), .A3(n6539), .A4(n6538), .ZN(n6542)
         );
  NAND4_X1 U7494 ( .A1(n6545), .A2(n6544), .A3(n6543), .A4(n6542), .ZN(n6747)
         );
  INV_X1 U7495 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6548) );
  INV_X1 U7496 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6547) );
  AOI22_X1 U7497 ( .A1(n6548), .A2(keyinput98), .B1(n6547), .B2(keyinput14), 
        .ZN(n6546) );
  OAI221_X1 U7498 ( .B1(n6548), .B2(keyinput98), .C1(n6547), .C2(keyinput14), 
        .A(n6546), .ZN(n6560) );
  AOI22_X1 U7499 ( .A1(n3944), .A2(keyinput107), .B1(n6550), .B2(keyinput115), 
        .ZN(n6549) );
  OAI221_X1 U7500 ( .B1(n3944), .B2(keyinput107), .C1(n6550), .C2(keyinput115), 
        .A(n6549), .ZN(n6559) );
  AOI22_X1 U7501 ( .A1(n6553), .A2(keyinput121), .B1(n6552), .B2(keyinput124), 
        .ZN(n6551) );
  OAI221_X1 U7502 ( .B1(n6553), .B2(keyinput121), .C1(n6552), .C2(keyinput124), 
        .A(n6551), .ZN(n6558) );
  INV_X1 U7503 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6556) );
  INV_X1 U7504 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6555) );
  AOI22_X1 U7505 ( .A1(n6556), .A2(keyinput52), .B1(keyinput23), .B2(n6555), 
        .ZN(n6554) );
  OAI221_X1 U7506 ( .B1(n6556), .B2(keyinput52), .C1(n6555), .C2(keyinput23), 
        .A(n6554), .ZN(n6557) );
  NOR4_X1 U7507 ( .A1(n6560), .A2(n6559), .A3(n6558), .A4(n6557), .ZN(n6611)
         );
  INV_X1 U7508 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6563) );
  AOI22_X1 U7509 ( .A1(n6563), .A2(keyinput66), .B1(keyinput63), .B2(n6562), 
        .ZN(n6561) );
  OAI221_X1 U7510 ( .B1(n6563), .B2(keyinput66), .C1(n6562), .C2(keyinput63), 
        .A(n6561), .ZN(n6576) );
  INV_X1 U7511 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6566) );
  INV_X1 U7512 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6565) );
  AOI22_X1 U7513 ( .A1(n6566), .A2(keyinput48), .B1(keyinput62), .B2(n6565), 
        .ZN(n6564) );
  OAI221_X1 U7514 ( .B1(n6566), .B2(keyinput48), .C1(n6565), .C2(keyinput62), 
        .A(n6564), .ZN(n6575) );
  INV_X1 U7515 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n6569) );
  AOI22_X1 U7516 ( .A1(n6569), .A2(keyinput31), .B1(keyinput91), .B2(n6568), 
        .ZN(n6567) );
  OAI221_X1 U7517 ( .B1(n6569), .B2(keyinput31), .C1(n6568), .C2(keyinput91), 
        .A(n6567), .ZN(n6574) );
  OAI221_X1 U7518 ( .B1(n6572), .B2(keyinput118), .C1(n6571), .C2(keyinput46), 
        .A(n6570), .ZN(n6573) );
  NOR4_X1 U7519 ( .A1(n6576), .A2(n6575), .A3(n6574), .A4(n6573), .ZN(n6610)
         );
  INV_X1 U7520 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6578) );
  AOI22_X1 U7521 ( .A1(n6579), .A2(keyinput84), .B1(n6578), .B2(keyinput20), 
        .ZN(n6577) );
  OAI221_X1 U7522 ( .B1(n6579), .B2(keyinput84), .C1(n6578), .C2(keyinput20), 
        .A(n6577), .ZN(n6591) );
  INV_X1 U7523 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6581) );
  AOI22_X1 U7524 ( .A1(n6581), .A2(keyinput61), .B1(keyinput28), .B2(n4850), 
        .ZN(n6580) );
  OAI221_X1 U7525 ( .B1(n6581), .B2(keyinput61), .C1(n4850), .C2(keyinput28), 
        .A(n6580), .ZN(n6590) );
  INV_X1 U7526 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n6584) );
  AOI22_X1 U7527 ( .A1(n6584), .A2(keyinput2), .B1(n6583), .B2(keyinput0), 
        .ZN(n6582) );
  OAI221_X1 U7528 ( .B1(n6584), .B2(keyinput2), .C1(n6583), .C2(keyinput0), 
        .A(n6582), .ZN(n6589) );
  INV_X1 U7529 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U7530 ( .A1(n6587), .A2(keyinput69), .B1(n6586), .B2(keyinput68), 
        .ZN(n6585) );
  OAI221_X1 U7531 ( .B1(n6587), .B2(keyinput69), .C1(n6586), .C2(keyinput68), 
        .A(n6585), .ZN(n6588) );
  NOR4_X1 U7532 ( .A1(n6591), .A2(n6590), .A3(n6589), .A4(n6588), .ZN(n6609)
         );
  INV_X1 U7533 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6594) );
  AOI22_X1 U7534 ( .A1(n6594), .A2(keyinput49), .B1(keyinput10), .B2(n6593), 
        .ZN(n6592) );
  OAI221_X1 U7535 ( .B1(n6594), .B2(keyinput49), .C1(n6593), .C2(keyinput10), 
        .A(n6592), .ZN(n6607) );
  AOI22_X1 U7536 ( .A1(n6597), .A2(keyinput3), .B1(n6596), .B2(keyinput104), 
        .ZN(n6595) );
  OAI221_X1 U7537 ( .B1(n6597), .B2(keyinput3), .C1(n6596), .C2(keyinput104), 
        .A(n6595), .ZN(n6606) );
  INV_X1 U7538 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6599) );
  AOI22_X1 U7539 ( .A1(n6600), .A2(keyinput73), .B1(n6599), .B2(keyinput54), 
        .ZN(n6598) );
  OAI221_X1 U7540 ( .B1(n6600), .B2(keyinput73), .C1(n6599), .C2(keyinput54), 
        .A(n6598), .ZN(n6605) );
  INV_X1 U7541 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6603) );
  INV_X1 U7542 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6602) );
  AOI22_X1 U7543 ( .A1(n6603), .A2(keyinput106), .B1(n6602), .B2(keyinput90), 
        .ZN(n6601) );
  OAI221_X1 U7544 ( .B1(n6603), .B2(keyinput106), .C1(n6602), .C2(keyinput90), 
        .A(n6601), .ZN(n6604) );
  NOR4_X1 U7545 ( .A1(n6607), .A2(n6606), .A3(n6605), .A4(n6604), .ZN(n6608)
         );
  NAND4_X1 U7546 ( .A1(n6611), .A2(n6610), .A3(n6609), .A4(n6608), .ZN(n6746)
         );
  INV_X1 U7547 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6614) );
  AOI22_X1 U7548 ( .A1(n6614), .A2(keyinput59), .B1(keyinput71), .B2(n6613), 
        .ZN(n6612) );
  OAI221_X1 U7549 ( .B1(n6614), .B2(keyinput59), .C1(n6613), .C2(keyinput71), 
        .A(n6612), .ZN(n6627) );
  AOI22_X1 U7550 ( .A1(n6617), .A2(keyinput41), .B1(keyinput33), .B2(n6616), 
        .ZN(n6615) );
  OAI221_X1 U7551 ( .B1(n6617), .B2(keyinput41), .C1(n6616), .C2(keyinput33), 
        .A(n6615), .ZN(n6626) );
  INV_X1 U7552 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n6620) );
  INV_X1 U7553 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6619) );
  AOI22_X1 U7554 ( .A1(n6620), .A2(keyinput95), .B1(n6619), .B2(keyinput45), 
        .ZN(n6618) );
  OAI221_X1 U7555 ( .B1(n6620), .B2(keyinput95), .C1(n6619), .C2(keyinput45), 
        .A(n6618), .ZN(n6625) );
  INV_X1 U7556 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6623) );
  AOI22_X1 U7557 ( .A1(n6623), .A2(keyinput123), .B1(keyinput113), .B2(n6622), 
        .ZN(n6621) );
  OAI221_X1 U7558 ( .B1(n6623), .B2(keyinput123), .C1(n6622), .C2(keyinput113), 
        .A(n6621), .ZN(n6624) );
  NOR4_X1 U7559 ( .A1(n6627), .A2(n6626), .A3(n6625), .A4(n6624), .ZN(n6676)
         );
  AOI22_X1 U7560 ( .A1(n6630), .A2(keyinput89), .B1(keyinput103), .B2(n6629), 
        .ZN(n6628) );
  OAI221_X1 U7561 ( .B1(n6630), .B2(keyinput89), .C1(n6629), .C2(keyinput103), 
        .A(n6628), .ZN(n6643) );
  INV_X1 U7562 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6636) );
  INV_X1 U7563 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n6635) );
  AOI22_X1 U7564 ( .A1(n6636), .A2(keyinput94), .B1(n6635), .B2(keyinput43), 
        .ZN(n6634) );
  OAI221_X1 U7565 ( .B1(n6636), .B2(keyinput94), .C1(n6635), .C2(keyinput43), 
        .A(n6634), .ZN(n6641) );
  AOI22_X1 U7566 ( .A1(n6639), .A2(keyinput51), .B1(n6638), .B2(keyinput85), 
        .ZN(n6637) );
  OAI221_X1 U7567 ( .B1(n6639), .B2(keyinput51), .C1(n6638), .C2(keyinput85), 
        .A(n6637), .ZN(n6640) );
  NOR4_X1 U7568 ( .A1(n6643), .A2(n6642), .A3(n6641), .A4(n6640), .ZN(n6675)
         );
  INV_X1 U7569 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6646) );
  AOI22_X1 U7570 ( .A1(n6646), .A2(keyinput111), .B1(keyinput11), .B2(n6645), 
        .ZN(n6644) );
  OAI221_X1 U7571 ( .B1(n6646), .B2(keyinput111), .C1(n6645), .C2(keyinput11), 
        .A(n6644), .ZN(n6659) );
  INV_X1 U7572 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n6649) );
  AOI22_X1 U7573 ( .A1(n6649), .A2(keyinput40), .B1(n6648), .B2(keyinput42), 
        .ZN(n6647) );
  OAI221_X1 U7574 ( .B1(n6649), .B2(keyinput40), .C1(n6648), .C2(keyinput42), 
        .A(n6647), .ZN(n6658) );
  INV_X1 U7575 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n6652) );
  AOI22_X1 U7576 ( .A1(n6652), .A2(keyinput30), .B1(n6651), .B2(keyinput9), 
        .ZN(n6650) );
  OAI221_X1 U7577 ( .B1(n6652), .B2(keyinput30), .C1(n6651), .C2(keyinput9), 
        .A(n6650), .ZN(n6657) );
  INV_X1 U7578 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6654) );
  AOI22_X1 U7579 ( .A1(n6655), .A2(keyinput29), .B1(n6654), .B2(keyinput105), 
        .ZN(n6653) );
  OAI221_X1 U7580 ( .B1(n6655), .B2(keyinput29), .C1(n6654), .C2(keyinput105), 
        .A(n6653), .ZN(n6656) );
  NOR4_X1 U7581 ( .A1(n6659), .A2(n6658), .A3(n6657), .A4(n6656), .ZN(n6674)
         );
  INV_X1 U7582 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6661) );
  AOI22_X1 U7583 ( .A1(n4722), .A2(keyinput77), .B1(n6661), .B2(keyinput36), 
        .ZN(n6660) );
  OAI221_X1 U7584 ( .B1(n4722), .B2(keyinput77), .C1(n6661), .C2(keyinput36), 
        .A(n6660), .ZN(n6672) );
  AOI22_X1 U7585 ( .A1(n6663), .A2(keyinput81), .B1(n4897), .B2(keyinput79), 
        .ZN(n6662) );
  OAI221_X1 U7586 ( .B1(n6663), .B2(keyinput81), .C1(n4897), .C2(keyinput79), 
        .A(n6662), .ZN(n6671) );
  INV_X1 U7587 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n6665) );
  AOI22_X1 U7588 ( .A1(n6665), .A2(keyinput117), .B1(n4994), .B2(keyinput22), 
        .ZN(n6664) );
  OAI221_X1 U7589 ( .B1(n6665), .B2(keyinput117), .C1(n4994), .C2(keyinput22), 
        .A(n6664), .ZN(n6670) );
  AOI22_X1 U7590 ( .A1(n6668), .A2(keyinput12), .B1(n6667), .B2(keyinput25), 
        .ZN(n6666) );
  OAI221_X1 U7591 ( .B1(n6668), .B2(keyinput12), .C1(n6667), .C2(keyinput25), 
        .A(n6666), .ZN(n6669) );
  NOR4_X1 U7592 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n6673)
         );
  NAND4_X1 U7593 ( .A1(n6676), .A2(n6675), .A3(n6674), .A4(n6673), .ZN(n6745)
         );
  AOI22_X1 U7594 ( .A1(n6679), .A2(keyinput96), .B1(keyinput38), .B2(n6678), 
        .ZN(n6677) );
  OAI221_X1 U7595 ( .B1(n6679), .B2(keyinput96), .C1(n6678), .C2(keyinput38), 
        .A(n6677), .ZN(n6692) );
  INV_X1 U7596 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6681) );
  AOI22_X1 U7597 ( .A1(n6682), .A2(keyinput6), .B1(n6681), .B2(keyinput97), 
        .ZN(n6680) );
  OAI221_X1 U7598 ( .B1(n6682), .B2(keyinput6), .C1(n6681), .C2(keyinput97), 
        .A(n6680), .ZN(n6691) );
  INV_X1 U7599 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6685) );
  AOI22_X1 U7600 ( .A1(n6685), .A2(keyinput35), .B1(n6684), .B2(keyinput82), 
        .ZN(n6683) );
  OAI221_X1 U7601 ( .B1(n6685), .B2(keyinput35), .C1(n6684), .C2(keyinput82), 
        .A(n6683), .ZN(n6690) );
  INV_X1 U7602 ( .A(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n6688) );
  INV_X1 U7603 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6687) );
  AOI22_X1 U7604 ( .A1(n6688), .A2(keyinput58), .B1(n6687), .B2(keyinput78), 
        .ZN(n6686) );
  OAI221_X1 U7605 ( .B1(n6688), .B2(keyinput58), .C1(n6687), .C2(keyinput78), 
        .A(n6686), .ZN(n6689) );
  NOR4_X1 U7606 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n6743)
         );
  INV_X1 U7607 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6694) );
  AOI22_X1 U7608 ( .A1(n6695), .A2(keyinput93), .B1(n6694), .B2(keyinput15), 
        .ZN(n6693) );
  OAI221_X1 U7609 ( .B1(n6695), .B2(keyinput93), .C1(n6694), .C2(keyinput15), 
        .A(n6693), .ZN(n6708) );
  INV_X1 U7610 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6698) );
  AOI22_X1 U7611 ( .A1(n6698), .A2(keyinput76), .B1(keyinput16), .B2(n6697), 
        .ZN(n6696) );
  OAI221_X1 U7612 ( .B1(n6698), .B2(keyinput76), .C1(n6697), .C2(keyinput16), 
        .A(n6696), .ZN(n6707) );
  AOI22_X1 U7613 ( .A1(n6701), .A2(keyinput102), .B1(keyinput86), .B2(n6700), 
        .ZN(n6699) );
  OAI221_X1 U7614 ( .B1(n6701), .B2(keyinput102), .C1(n6700), .C2(keyinput86), 
        .A(n6699), .ZN(n6706) );
  INV_X1 U7615 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6704) );
  AOI22_X1 U7616 ( .A1(n6704), .A2(keyinput18), .B1(keyinput32), .B2(n6703), 
        .ZN(n6702) );
  OAI221_X1 U7617 ( .B1(n6704), .B2(keyinput18), .C1(n6703), .C2(keyinput32), 
        .A(n6702), .ZN(n6705) );
  NOR4_X1 U7618 ( .A1(n6708), .A2(n6707), .A3(n6706), .A4(n6705), .ZN(n6742)
         );
  INV_X1 U7619 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6710) );
  AOI22_X1 U7620 ( .A1(n6711), .A2(keyinput55), .B1(n6710), .B2(keyinput110), 
        .ZN(n6709) );
  OAI221_X1 U7621 ( .B1(n6711), .B2(keyinput55), .C1(n6710), .C2(keyinput110), 
        .A(n6709), .ZN(n6724) );
  INV_X1 U7622 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n6714) );
  INV_X1 U7623 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6713) );
  AOI22_X1 U7624 ( .A1(n6714), .A2(keyinput75), .B1(n6713), .B2(keyinput26), 
        .ZN(n6712) );
  OAI221_X1 U7625 ( .B1(n6714), .B2(keyinput75), .C1(n6713), .C2(keyinput26), 
        .A(n6712), .ZN(n6723) );
  INV_X1 U7626 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6717) );
  INV_X1 U7627 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6716) );
  AOI22_X1 U7628 ( .A1(n6717), .A2(keyinput67), .B1(keyinput65), .B2(n6716), 
        .ZN(n6715) );
  OAI221_X1 U7629 ( .B1(n6717), .B2(keyinput67), .C1(n6716), .C2(keyinput65), 
        .A(n6715), .ZN(n6722) );
  AOI22_X1 U7630 ( .A1(n6720), .A2(keyinput24), .B1(keyinput1), .B2(n6719), 
        .ZN(n6718) );
  OAI221_X1 U7631 ( .B1(n6720), .B2(keyinput24), .C1(n6719), .C2(keyinput1), 
        .A(n6718), .ZN(n6721) );
  NOR4_X1 U7632 ( .A1(n6724), .A2(n6723), .A3(n6722), .A4(n6721), .ZN(n6741)
         );
  INV_X1 U7633 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n6726) );
  AOI22_X1 U7634 ( .A1(n6726), .A2(keyinput70), .B1(n4450), .B2(keyinput8), 
        .ZN(n6725) );
  OAI221_X1 U7635 ( .B1(n6726), .B2(keyinput70), .C1(n4450), .C2(keyinput8), 
        .A(n6725), .ZN(n6739) );
  INV_X1 U7636 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n6728) );
  AOI22_X1 U7637 ( .A1(n6729), .A2(keyinput126), .B1(keyinput37), .B2(n6728), 
        .ZN(n6727) );
  OAI221_X1 U7638 ( .B1(n6729), .B2(keyinput126), .C1(n6728), .C2(keyinput37), 
        .A(n6727), .ZN(n6738) );
  AOI22_X1 U7639 ( .A1(n6732), .A2(keyinput21), .B1(n6731), .B2(keyinput7), 
        .ZN(n6730) );
  OAI221_X1 U7640 ( .B1(n6732), .B2(keyinput21), .C1(n6731), .C2(keyinput7), 
        .A(n6730), .ZN(n6737) );
  INV_X1 U7641 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6735) );
  AOI22_X1 U7642 ( .A1(n6735), .A2(keyinput17), .B1(n6734), .B2(keyinput19), 
        .ZN(n6733) );
  OAI221_X1 U7643 ( .B1(n6735), .B2(keyinput17), .C1(n6734), .C2(keyinput19), 
        .A(n6733), .ZN(n6736) );
  NOR4_X1 U7644 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6740)
         );
  NAND4_X1 U7645 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6744)
         );
  NOR4_X1 U7646 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6748)
         );
  XOR2_X1 U7647 ( .A(n6749), .B(n6748), .Z(n6752) );
  NAND2_X1 U7648 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6750), .ZN(n6751) );
  XNOR2_X1 U7649 ( .A(n6752), .B(n6751), .ZN(U3153) );
  AND2_X2 U4621 ( .A1(n5158), .A2(n4992), .ZN(n5136) );
  OAI21_X1 U3602 ( .B1(n4239), .B2(STATE2_REG_0__SCAN_IN), .A(n3281), .ZN(
        n3337) );
  CLKBUF_X1 U3776 ( .A(n4598), .Z(n4609) );
  CLKBUF_X2 U3827 ( .A(n3993), .Z(n3096) );
  CLKBUF_X1 U3970 ( .A(n4822), .Z(n4947) );
  CLKBUF_X1 U4220 ( .A(n5658), .Z(n5648) );
endmodule

