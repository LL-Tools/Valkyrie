

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689;

  INV_X4 U4915 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AND4_X1 U4916 ( .A1(n6118), .A2(n6117), .A3(n6116), .A4(n6115), .ZN(n9375)
         );
  NAND2_X1 U4917 ( .A1(n6107), .A2(n6106), .ZN(n7566) );
  AND4_X1 U4918 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n7691)
         );
  NAND2_X2 U4919 ( .A1(n7074), .A2(n8295), .ZN(n6366) );
  AND2_X2 U4920 ( .A1(n6038), .A2(n6035), .ZN(n6856) );
  NAND2_X1 U4921 ( .A1(n6009), .A2(n6008), .ZN(n9601) );
  INV_X1 U4922 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6226) );
  INV_X4 U4923 ( .A(n10163), .ZN(n4856) );
  INV_X1 U4924 ( .A(n6079), .ZN(n6478) );
  AND2_X2 U4925 ( .A1(n4862), .A2(n6707), .ZN(n9046) );
  INV_X1 U4926 ( .A(n8544), .ZN(n5711) );
  MUX2_X1 U4927 ( .A(n8639), .B(n8636), .S(n8760), .Z(n8637) );
  AND3_X1 U4928 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5443) );
  INV_X1 U4929 ( .A(n7546), .ZN(n4854) );
  NAND2_X1 U4930 ( .A1(n7371), .A2(n6186), .ZN(n7374) );
  AND2_X1 U4932 ( .A1(n6091), .A2(n6090), .ZN(n10507) );
  OR2_X1 U4933 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  NAND4_X1 U4934 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n10536)
         );
  NAND2_X2 U4935 ( .A1(n5899), .A2(n6785), .ZN(n6646) );
  CLKBUF_X3 U4936 ( .A(n5403), .Z(n4851) );
  NOR2_X2 U4937 ( .A1(n5812), .A2(n5811), .ZN(n5832) );
  OAI21_X4 U4938 ( .B1(n5721), .B2(n5720), .A(n5719), .ZN(n5736) );
  OAI21_X2 U4939 ( .B1(n5683), .B2(n5164), .A(n5161), .ZN(n5721) );
  XNOR2_X2 U4940 ( .A(n5890), .B(n5889), .ZN(n9041) );
  OAI22_X2 U4941 ( .A1(n9550), .A2(n9431), .B1(n9571), .B2(n9682), .ZN(n9539)
         );
  CLKBUF_X1 U4942 ( .A(n5403), .Z(n4850) );
  NAND2_X1 U4943 ( .A1(n5336), .A2(n5337), .ZN(n5403) );
  AND2_X1 U4944 ( .A1(n4862), .A2(n6707), .ZN(n4852) );
  XNOR2_X1 U4945 ( .A(n9375), .B(n7566), .ZN(n8497) );
  NAND2_X1 U4946 ( .A1(n6020), .A2(n8340), .ZN(n4853) );
  NAND2_X2 U4947 ( .A1(n6020), .A2(n8340), .ZN(n6079) );
  XNOR2_X1 U4948 ( .A(n10527), .B(n10536), .ZN(n8499) );
  XNOR2_X2 U4950 ( .A(n6034), .B(n6033), .ZN(n6035) );
  AOI211_X2 U4951 ( .C1(n8611), .C2(n8675), .A(n10076), .B(n8610), .ZN(n8617)
         );
  NAND2_X2 U4952 ( .A1(n5496), .A2(n5495), .ZN(n8277) );
  NAND2_X1 U4953 ( .A1(n7374), .A2(n5190), .ZN(n10613) );
  NAND2_X1 U4954 ( .A1(n6722), .A2(n10160), .ZN(n9863) );
  NOR2_X1 U4955 ( .A1(n6948), .A2(n6483), .ZN(n6068) );
  OR2_X1 U4956 ( .A1(n6914), .A2(n7326), .ZN(n8778) );
  INV_X1 U4957 ( .A(n7633), .ZN(n10478) );
  INV_X1 U4958 ( .A(n6911), .ZN(n7326) );
  NAND4_X1 U4959 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(n9377)
         );
  INV_X1 U4960 ( .A(n9041), .ZN(n8825) );
  CLKBUF_X2 U4961 ( .A(P1_U4006), .Z(n4857) );
  CLKBUF_X2 U4962 ( .A(n5441), .Z(n5883) );
  OR3_X1 U4963 ( .A1(n8096), .A2(n7866), .A3(n8058), .ZN(n6885) );
  INV_X4 U4965 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  OR2_X1 U4966 ( .A1(n6441), .A2(n5201), .ZN(n5198) );
  NAND2_X1 U4967 ( .A1(n5267), .A2(n5266), .ZN(n9460) );
  XNOR2_X1 U4968 ( .A(n6426), .B(n6424), .ZN(n9077) );
  NAND2_X1 U4969 ( .A1(n9115), .A2(n6413), .ZN(n6426) );
  OAI21_X1 U4970 ( .B1(n8226), .B2(n5213), .A(n5210), .ZN(n4939) );
  NOR2_X1 U4971 ( .A1(n4871), .A2(n8324), .ZN(n5107) );
  INV_X1 U4972 ( .A(n9986), .ZN(n8678) );
  OAI21_X1 U4973 ( .B1(n5942), .B2(n5060), .A(n5058), .ZN(n10133) );
  AOI21_X1 U4974 ( .B1(n5212), .B2(n5214), .A(n5211), .ZN(n5210) );
  NAND2_X1 U4975 ( .A1(n5935), .A2(n5934), .ZN(n7887) );
  INV_X1 U4976 ( .A(n6382), .ZN(n5211) );
  NAND2_X1 U4977 ( .A1(n5740), .A2(n5739), .ZN(n10217) );
  NAND2_X1 U4978 ( .A1(n6172), .A2(n10562), .ZN(n7371) );
  NAND2_X1 U4979 ( .A1(n6352), .A2(n6351), .ZN(n9700) );
  NAND2_X1 U4980 ( .A1(n6323), .A2(n6322), .ZN(n9710) );
  NAND2_X1 U4981 ( .A1(n6231), .A2(n6230), .ZN(n8975) );
  NAND3_X1 U4982 ( .A1(n4955), .A2(n7181), .A3(n7182), .ZN(n7335) );
  NAND2_X1 U4983 ( .A1(n7100), .A2(n5029), .ZN(n7412) );
  NAND2_X1 U4984 ( .A1(n7101), .A2(n5916), .ZN(n7100) );
  NAND2_X1 U4985 ( .A1(n5537), .A2(n5536), .ZN(n10596) );
  NAND2_X2 U4986 ( .A1(n6126), .A2(n6125), .ZN(n10527) );
  OAI21_X1 U4987 ( .B1(n5487), .B2(n5151), .A(n5149), .ZN(n5526) );
  NAND2_X1 U4988 ( .A1(n5472), .A2(n5471), .ZN(n5487) );
  INV_X2 U4989 ( .A(n10657), .ZN(n4855) );
  AOI21_X1 U4990 ( .B1(n6946), .B2(n6945), .A(n6944), .ZN(n7619) );
  INV_X4 U4991 ( .A(n7385), .ZN(n6912) );
  NAND4_X2 U4992 ( .A1(n5389), .A2(n5388), .A3(n5387), .A4(n5386), .ZN(n9900)
         );
  NAND2_X1 U4993 ( .A1(n5400), .A2(n5399), .ZN(n5420) );
  NAND2_X1 U4994 ( .A1(n6708), .A2(n6885), .ZN(n7385) );
  NAND4_X1 U4995 ( .A1(n5440), .A2(n5439), .A3(n5438), .A4(n5437), .ZN(n9898)
         );
  NAND2_X2 U4996 ( .A1(n5188), .A2(n10467), .ZN(n8527) );
  INV_X1 U4997 ( .A(n6895), .ZN(n6708) );
  NAND2_X1 U4998 ( .A1(n5068), .A2(n4880), .ZN(n7633) );
  NAND2_X1 U4999 ( .A1(n5003), .A2(n4891), .ZN(n7546) );
  NAND2_X1 U5000 ( .A1(n7527), .A2(n9601), .ZN(n6539) );
  INV_X1 U5001 ( .A(n8532), .ZN(n8537) );
  NAND2_X1 U5002 ( .A1(n5895), .A2(n5709), .ZN(n9944) );
  NAND2_X1 U5003 ( .A1(n5338), .A2(n5337), .ZN(n5441) );
  OR2_X1 U5004 ( .A1(n4850), .A2(n6671), .ZN(n5343) );
  AND2_X2 U5005 ( .A1(n5338), .A2(n5339), .ZN(n6624) );
  NAND2_X1 U5006 ( .A1(n6008), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5189) );
  MUX2_X1 U5008 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5708), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5709) );
  NAND2_X2 U5009 ( .A1(n6646), .A2(n5356), .ZN(n8544) );
  AND2_X1 U5010 ( .A1(n5463), .A2(n5466), .ZN(n5465) );
  NAND2_X1 U5011 ( .A1(n6503), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6509) );
  XNOR2_X1 U5012 ( .A(n5968), .B(n5967), .ZN(n8096) );
  NAND2_X1 U5013 ( .A1(n10285), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5330) );
  INV_X2 U5014 ( .A(n9740), .ZN(n8538) );
  OR2_X1 U5015 ( .A1(n6032), .A2(n6515), .ZN(n6034) );
  XNOR2_X1 U5016 ( .A(n6025), .B(n6024), .ZN(n6547) );
  OR2_X1 U5017 ( .A1(n5332), .A2(n5331), .ZN(n5334) );
  INV_X2 U5018 ( .A(n6639), .ZN(n4858) );
  AND2_X1 U5019 ( .A1(n5345), .A2(n5346), .ZN(n5332) );
  NAND2_X1 U5020 ( .A1(n5073), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6025) );
  AND4_X1 U5021 ( .A1(n5171), .A2(n5170), .A3(n5175), .A4(n5033), .ZN(n5345)
         );
  AND3_X1 U5022 ( .A1(n5325), .A2(n5326), .A3(n5169), .ZN(n5171) );
  AND2_X1 U5023 ( .A1(n4877), .A2(n6086), .ZN(n5071) );
  AND2_X1 U5024 ( .A1(n5327), .A2(n5551), .ZN(n5170) );
  NAND2_X1 U5025 ( .A1(n5443), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5479) );
  AND2_X1 U5026 ( .A1(n5969), .A2(n5987), .ZN(n5169) );
  AND3_X1 U5027 ( .A1(n5318), .A2(n5317), .A3(n5316), .ZN(n5551) );
  INV_X1 U5028 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5969) );
  NOR2_X1 U5029 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6001) );
  INV_X1 U5030 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5594) );
  INV_X1 U5031 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5987) );
  NOR2_X1 U5032 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5323) );
  NOR2_X1 U5033 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5319) );
  NOR2_X1 U5034 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5320) );
  NOR2_X1 U5035 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5316) );
  NOR2_X1 U5036 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5317) );
  NOR2_X1 U5037 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5318) );
  NOR2_X1 U5038 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5304) );
  INV_X1 U5039 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5374) );
  INV_X1 U5040 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6227) );
  INV_X1 U5041 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6010) );
  INV_X1 U5042 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6270) );
  NAND2_X2 U5043 ( .A1(n7343), .A2(n7344), .ZN(n7513) );
  NAND2_X2 U5044 ( .A1(n7348), .A2(n7346), .ZN(n7343) );
  NAND2_X1 U5045 ( .A1(n7486), .A2(n5958), .ZN(n6895) );
  CLKBUF_X1 U5046 ( .A(n5361), .Z(n4859) );
  BUF_X4 U5047 ( .A(n5361), .Z(n4860) );
  INV_X8 U5048 ( .A(n7385), .ZN(n9042) );
  NAND2_X2 U5049 ( .A1(n5959), .A2(n6701), .ZN(n6896) );
  NAND2_X1 U5050 ( .A1(n6896), .A2(n6895), .ZN(n7173) );
  INV_X1 U5051 ( .A(n7514), .ZN(n4862) );
  XNOR2_X2 U5052 ( .A(n5330), .B(n5329), .ZN(n5336) );
  NAND2_X1 U5053 ( .A1(n5573), .A2(n5572), .ZN(n5590) );
  NAND2_X1 U5054 ( .A1(n6895), .A2(n6885), .ZN(n7514) );
  NOR2_X1 U5055 ( .A1(n5943), .A2(n5064), .ZN(n5063) );
  INV_X1 U5056 ( .A(n5941), .ZN(n5064) );
  INV_X1 U5057 ( .A(n5259), .ZN(n5258) );
  NAND2_X1 U5058 ( .A1(n5631), .A2(n9285), .ZN(n5645) );
  NOR2_X1 U5059 ( .A1(n5504), .A2(n5153), .ZN(n5152) );
  INV_X1 U5060 ( .A(n5489), .ZN(n5153) );
  NAND2_X1 U5061 ( .A1(n5490), .A2(n9300), .ZN(n5506) );
  INV_X1 U5062 ( .A(n6319), .ZN(n5226) );
  AND2_X1 U5063 ( .A1(n8335), .A2(n8482), .ZN(n8491) );
  AND2_X1 U5064 ( .A1(n9661), .A2(n9479), .ZN(n8492) );
  OR2_X1 U5065 ( .A1(n9703), .A2(n9596), .ZN(n8358) );
  OR2_X1 U5066 ( .A1(n8989), .A2(n8970), .ZN(n8436) );
  INV_X1 U5067 ( .A(n7554), .ZN(n5100) );
  NOR2_X1 U5068 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6063) );
  AND2_X1 U5069 ( .A1(n5242), .A2(n9842), .ZN(n5241) );
  OR2_X1 U5070 ( .A1(n5244), .A2(n9778), .ZN(n5240) );
  NAND2_X1 U5071 ( .A1(n9843), .A2(n5243), .ZN(n5242) );
  NAND2_X1 U5072 ( .A1(n5253), .A2(n5252), .ZN(n5251) );
  INV_X1 U5073 ( .A(n7511), .ZN(n5252) );
  INV_X1 U5074 ( .A(n7512), .ZN(n5253) );
  NAND2_X1 U5075 ( .A1(n4888), .A2(n7789), .ZN(n5248) );
  INV_X1 U5076 ( .A(n5250), .ZN(n5249) );
  AOI22_X1 U5077 ( .A1(n6912), .A2(n6902), .B1(n8234), .B2(n8776), .ZN(n6903)
         );
  NAND2_X1 U5078 ( .A1(n8845), .A2(n8844), .ZN(n8847) );
  OR2_X1 U5079 ( .A1(n10179), .A2(n9987), .ZN(n8628) );
  OR2_X1 U5080 ( .A1(n10196), .A2(n9997), .ZN(n8750) );
  NOR2_X1 U5081 ( .A1(n10143), .A2(n5002), .ZN(n5001) );
  INV_X1 U5082 ( .A(n8687), .ZN(n5002) );
  AND2_X1 U5083 ( .A1(n10143), .A2(n5065), .ZN(n5061) );
  OR2_X1 U5084 ( .A1(n10239), .A2(n9887), .ZN(n5065) );
  NOR2_X1 U5085 ( .A1(n8655), .A2(n5030), .ZN(n5029) );
  INV_X1 U5086 ( .A(n5917), .ZN(n5030) );
  NAND2_X1 U5087 ( .A1(n5787), .A2(n5131), .ZN(n5133) );
  NOR2_X1 U5088 ( .A1(n5802), .A2(n5132), .ZN(n5131) );
  INV_X1 U5089 ( .A(n5786), .ZN(n5132) );
  AOI21_X1 U5090 ( .B1(n5128), .B2(n5749), .A(n4914), .ZN(n5127) );
  NOR2_X1 U5091 ( .A1(n5735), .A2(n5129), .ZN(n5128) );
  INV_X1 U5092 ( .A(n5737), .ZN(n5129) );
  AND2_X1 U5093 ( .A1(n5228), .A2(n5613), .ZN(n4958) );
  NAND2_X1 U5094 ( .A1(n5590), .A2(n5575), .ZN(n5588) );
  XNOR2_X1 U5095 ( .A(n5566), .B(SI_11_), .ZN(n5565) );
  NAND2_X1 U5096 ( .A1(n5545), .A2(n5305), .ZN(n5547) );
  INV_X1 U5097 ( .A(n8085), .ZN(n5227) );
  INV_X2 U5098 ( .A(n8527), .ZN(n6483) );
  XNOR2_X1 U5099 ( .A(n8525), .B(n4972), .ZN(n4971) );
  INV_X1 U5100 ( .A(n8490), .ZN(n4972) );
  INV_X1 U5101 ( .A(n6109), .ZN(n6855) );
  NOR2_X1 U5102 ( .A1(n9450), .A2(n9423), .ZN(n9422) );
  AOI21_X1 U5103 ( .B1(n5269), .B2(n5272), .A(n4916), .ZN(n5266) );
  OR2_X1 U5104 ( .A1(n9682), .A2(n9092), .ZN(n8351) );
  INV_X1 U5105 ( .A(n5281), .ZN(n5280) );
  OAI21_X1 U5106 ( .B1(n8512), .B2(n5286), .A(n5285), .ZN(n5281) );
  OR2_X1 U5107 ( .A1(n9718), .A2(n9369), .ZN(n5285) );
  INV_X1 U5108 ( .A(n6366), .ZN(n6350) );
  INV_X1 U5109 ( .A(n7074), .ZN(n7022) );
  NAND2_X1 U5110 ( .A1(n7690), .A2(n5101), .ZN(n7606) );
  OR2_X1 U5111 ( .A1(n7058), .A2(n6547), .ZN(n9597) );
  NAND2_X1 U5112 ( .A1(n7074), .A2(n5356), .ZN(n6104) );
  NAND2_X1 U5113 ( .A1(n9742), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6031) );
  AND2_X1 U5114 ( .A1(n5215), .A2(n4895), .ZN(n5072) );
  INV_X1 U5115 ( .A(n6646), .ZN(n5710) );
  NAND2_X1 U5116 ( .A1(n6646), .A2(n8295), .ZN(n5428) );
  NAND2_X1 U5117 ( .A1(n7251), .A2(n7252), .ZN(n7250) );
  NAND2_X1 U5118 ( .A1(n5860), .A2(n5859), .ZN(n5875) );
  OR2_X1 U5119 ( .A1(n5345), .A2(n5331), .ZN(n5347) );
  INV_X1 U5120 ( .A(n8430), .ZN(n4960) );
  NAND2_X1 U5121 ( .A1(n4963), .A2(n4962), .ZN(n4961) );
  NOR2_X1 U5122 ( .A1(n8431), .A2(n7911), .ZN(n4962) );
  NAND2_X1 U5123 ( .A1(n4964), .A2(n8414), .ZN(n4963) );
  AND2_X1 U5124 ( .A1(n5080), .A2(n8446), .ZN(n4975) );
  NOR2_X1 U5125 ( .A1(n4873), .A2(n9477), .ZN(n5097) );
  INV_X1 U5126 ( .A(n8499), .ZN(n7569) );
  NAND2_X1 U5127 ( .A1(n4934), .A2(n6427), .ZN(n6440) );
  NAND2_X1 U5128 ( .A1(n9077), .A2(n9076), .ZN(n4934) );
  NAND2_X1 U5129 ( .A1(n8343), .A2(n8537), .ZN(n8485) );
  NAND2_X1 U5130 ( .A1(n8520), .A2(n8485), .ZN(n5142) );
  NAND2_X1 U5131 ( .A1(n8331), .A2(n8479), .ZN(n8332) );
  INV_X1 U5132 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5066) );
  OR2_X1 U5133 ( .A1(n9645), .A2(n8330), .ZN(n8479) );
  NOR2_X1 U5134 ( .A1(n9667), .A2(n9661), .ZN(n5012) );
  NOR2_X1 U5135 ( .A1(n9661), .A2(n9479), .ZN(n8493) );
  OR2_X1 U5136 ( .A1(n9676), .A2(n9558), .ZN(n8352) );
  AOI21_X1 U5137 ( .B1(n8146), .B2(n8441), .A(n5088), .ZN(n5087) );
  INV_X1 U5138 ( .A(n8445), .ZN(n5088) );
  OR2_X1 U5139 ( .A1(n9710), .A2(n8182), .ZN(n8363) );
  AND2_X1 U5140 ( .A1(n9714), .A2(n9368), .ZN(n5284) );
  INV_X1 U5141 ( .A(n8512), .ZN(n5282) );
  OAI21_X1 U5142 ( .B1(n5101), .B2(n5100), .A(n7555), .ZN(n5099) );
  NOR2_X1 U5143 ( .A1(n8497), .A2(n5102), .ZN(n5101) );
  INV_X1 U5144 ( .A(n7553), .ZN(n5102) );
  NOR2_X1 U5145 ( .A1(n8522), .A2(n9601), .ZN(n8343) );
  NAND2_X1 U5146 ( .A1(n6948), .A2(n7633), .ZN(n8377) );
  NOR2_X1 U5147 ( .A1(n9541), .A2(n9670), .ZN(n9507) );
  NAND2_X1 U5148 ( .A1(n8504), .A2(n7587), .ZN(n5265) );
  OR2_X1 U5149 ( .A1(n8497), .A2(n7568), .ZN(n7650) );
  OR2_X1 U5150 ( .A1(n9001), .A2(n9000), .ZN(n9007) );
  XNOR2_X1 U5151 ( .A(n6897), .B(n8946), .ZN(n7178) );
  INV_X1 U5152 ( .A(n8207), .ZN(n8210) );
  INV_X1 U5153 ( .A(n5956), .ZN(n5037) );
  OR2_X1 U5154 ( .A1(n5963), .A2(n9961), .ZN(n8629) );
  OR2_X1 U5155 ( .A1(n10007), .A2(n10026), .ZN(n8751) );
  INV_X1 U5156 ( .A(n10014), .ZN(n5057) );
  OR2_X1 U5157 ( .A1(n10201), .A2(n10025), .ZN(n8745) );
  OR2_X1 U5158 ( .A1(n10211), .A2(n10091), .ZN(n8695) );
  NAND2_X1 U5159 ( .A1(n5942), .A2(n5063), .ZN(n5062) );
  OR2_X1 U5160 ( .A1(n10246), .A2(n5179), .ZN(n5178) );
  AND2_X1 U5161 ( .A1(n8739), .A2(n8702), .ZN(n8669) );
  OR2_X1 U5162 ( .A1(n10249), .A2(n10257), .ZN(n5179) );
  NOR2_X1 U5163 ( .A1(n5932), .A2(n4980), .ZN(n4979) );
  INV_X1 U5164 ( .A(n8706), .ZN(n4982) );
  OR2_X1 U5165 ( .A1(n6892), .A2(n10485), .ZN(n8785) );
  NAND2_X1 U5166 ( .A1(n5879), .A2(n5878), .ZN(n8287) );
  INV_X1 U5167 ( .A(n5768), .ZN(n5122) );
  NAND2_X1 U5168 ( .A1(n5254), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5892) );
  NOR2_X1 U5169 ( .A1(n5256), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U5170 ( .A1(n5258), .A2(n5257), .ZN(n5256) );
  AND2_X1 U5171 ( .A1(n5737), .A2(n5724), .ZN(n5735) );
  AOI21_X1 U5172 ( .B1(n5163), .B2(n5162), .A(n4915), .ZN(n5161) );
  INV_X1 U5173 ( .A(n5685), .ZN(n5162) );
  OAI21_X1 U5174 ( .B1(n5610), .B2(n4875), .A(n5134), .ZN(n5665) );
  INV_X1 U5175 ( .A(n5135), .ZN(n5134) );
  OAI21_X1 U5176 ( .B1(n5138), .B2(n4875), .A(n5645), .ZN(n5135) );
  AND2_X1 U5177 ( .A1(n5666), .A2(n5650), .ZN(n5664) );
  NOR2_X1 U5178 ( .A1(n5629), .A2(n5139), .ZN(n5138) );
  INV_X1 U5179 ( .A(n5609), .ZN(n5139) );
  INV_X1 U5180 ( .A(n5626), .ZN(n5629) );
  XNOR2_X1 U5181 ( .A(n5627), .B(n9163), .ZN(n5626) );
  INV_X1 U5182 ( .A(n5156), .ZN(n5155) );
  OAI21_X1 U5183 ( .B1(n5159), .B2(n4876), .A(n5590), .ZN(n5156) );
  NOR2_X1 U5184 ( .A1(n5569), .A2(n5160), .ZN(n5159) );
  INV_X1 U5185 ( .A(n5546), .ZN(n5160) );
  INV_X1 U5186 ( .A(n5565), .ZN(n5569) );
  NAND2_X1 U5187 ( .A1(n5567), .A2(SI_11_), .ZN(n5568) );
  NAND2_X1 U5188 ( .A1(n5528), .A2(n5527), .ZN(n5545) );
  NAND2_X1 U5189 ( .A1(n5526), .A2(n5313), .ZN(n5528) );
  AND2_X1 U5190 ( .A1(n5546), .A2(n5532), .ZN(n5305) );
  NAND2_X1 U5191 ( .A1(n5506), .A2(n5492), .ZN(n5504) );
  XNOR2_X1 U5192 ( .A(n5425), .B(SI_5_), .ZN(n5451) );
  AND2_X1 U5193 ( .A1(n4929), .A2(n6099), .ZN(n10494) );
  OR2_X1 U5194 ( .A1(n6084), .A2(n6085), .ZN(n4929) );
  OR2_X1 U5195 ( .A1(n6354), .A2(n6353), .ZN(n6370) );
  OR2_X1 U5196 ( .A1(n6247), .A2(n6235), .ZN(n6276) );
  NAND2_X1 U5197 ( .A1(n10613), .A2(n6209), .ZN(n7502) );
  NAND2_X1 U5198 ( .A1(n4853), .A2(n4854), .ZN(n5192) );
  NOR2_X1 U5199 ( .A1(n4854), .A2(n5195), .ZN(n5194) );
  NOR2_X1 U5200 ( .A1(n5225), .A2(n4941), .ZN(n4940) );
  INV_X1 U5201 ( .A(n6297), .ZN(n4941) );
  NAND2_X1 U5202 ( .A1(n4933), .A2(n4932), .ZN(n6441) );
  INV_X1 U5203 ( .A(n6439), .ZN(n4932) );
  INV_X1 U5204 ( .A(n6440), .ZN(n4933) );
  NAND2_X1 U5205 ( .A1(n6275), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6307) );
  INV_X1 U5206 ( .A(n6276), .ZN(n6275) );
  AOI21_X1 U5207 ( .B1(n8990), .B2(n5206), .A(n4879), .ZN(n5205) );
  INV_X1 U5208 ( .A(n6266), .ZN(n5206) );
  AND2_X1 U5209 ( .A1(n8532), .A2(n5187), .ZN(n7024) );
  NAND2_X1 U5210 ( .A1(n8303), .A2(n8302), .ZN(n9423) );
  OR2_X1 U5211 ( .A1(n9645), .A2(n9449), .ZN(n9450) );
  AND2_X1 U5212 ( .A1(n8479), .A2(n8480), .ZN(n9440) );
  XNOR2_X1 U5213 ( .A(n9650), .B(n9480), .ZN(n9438) );
  OR2_X1 U5214 ( .A1(n9655), .A2(n9142), .ZN(n8472) );
  INV_X1 U5215 ( .A(n9438), .ZN(n9465) );
  OAI21_X1 U5216 ( .B1(n9560), .B2(n5107), .A(n5104), .ZN(n8327) );
  INV_X1 U5217 ( .A(n5105), .ZN(n5104) );
  NOR2_X1 U5218 ( .A1(n9490), .A2(n9504), .ZN(n5273) );
  OR2_X1 U5219 ( .A1(n9667), .A2(n9528), .ZN(n9488) );
  NOR2_X1 U5220 ( .A1(n8493), .A2(n8492), .ZN(n9490) );
  OR2_X1 U5221 ( .A1(n9670), .A2(n9107), .ZN(n9501) );
  INV_X1 U5222 ( .A(n5103), .ZN(n9502) );
  AOI21_X1 U5223 ( .B1(n9560), .B2(n5108), .A(n5107), .ZN(n5103) );
  OR2_X1 U5224 ( .A1(n9670), .A2(n9536), .ZN(n9433) );
  NAND2_X1 U5225 ( .A1(n9560), .A2(n5106), .ZN(n9535) );
  INV_X1 U5226 ( .A(n5109), .ZN(n5106) );
  NAND2_X1 U5227 ( .A1(n5076), .A2(n5074), .ZN(n8321) );
  NOR2_X1 U5228 ( .A1(n4874), .A2(n5075), .ZN(n5074) );
  OR2_X1 U5229 ( .A1(n9692), .A2(n9598), .ZN(n8454) );
  OR2_X1 U5230 ( .A1(n9581), .A2(n9598), .ZN(n5307) );
  NOR2_X1 U5231 ( .A1(n9568), .A2(n5292), .ZN(n5291) );
  INV_X1 U5232 ( .A(n5307), .ZN(n5292) );
  NAND2_X1 U5233 ( .A1(n8454), .A2(n8450), .ZN(n9582) );
  NAND2_X1 U5234 ( .A1(n9577), .A2(n9582), .ZN(n9576) );
  INV_X1 U5235 ( .A(n5087), .ZN(n5085) );
  AOI21_X1 U5236 ( .B1(n5087), .B2(n5084), .A(n5083), .ZN(n5082) );
  INV_X1 U5237 ( .A(n8444), .ZN(n5083) );
  INV_X1 U5238 ( .A(n8441), .ZN(n5084) );
  AND2_X1 U5239 ( .A1(n5280), .A2(n5278), .ZN(n5277) );
  INV_X1 U5240 ( .A(n8513), .ZN(n5278) );
  NAND2_X1 U5241 ( .A1(n8133), .A2(n5282), .ZN(n5279) );
  AND2_X1 U5242 ( .A1(n8445), .A2(n8444), .ZN(n8513) );
  AND2_X1 U5243 ( .A1(n8440), .A2(n8441), .ZN(n8512) );
  OR2_X1 U5244 ( .A1(n10668), .A2(n8991), .ZN(n5314) );
  AND2_X1 U5245 ( .A1(n8436), .A2(n8437), .ZN(n8510) );
  AND4_X1 U5246 ( .A1(n6282), .A2(n6281), .A3(n6280), .A4(n6279), .ZN(n8970)
         );
  NAND2_X1 U5247 ( .A1(n7910), .A2(n5297), .ZN(n7919) );
  AND2_X1 U5248 ( .A1(n7911), .A2(n7909), .ZN(n5297) );
  INV_X1 U5249 ( .A(n6215), .ZN(n6214) );
  AOI21_X1 U5250 ( .B1(n4863), .B2(n5091), .A(n4899), .ZN(n5090) );
  INV_X1 U5251 ( .A(n8401), .ZN(n5091) );
  NAND2_X1 U5252 ( .A1(n5093), .A2(n8401), .ZN(n5092) );
  INV_X1 U5253 ( .A(n7674), .ZN(n5093) );
  INV_X1 U5254 ( .A(n8501), .ZN(n7573) );
  AND4_X1 U5255 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .ZN(n7656)
         );
  NAND2_X1 U5256 ( .A1(n7552), .A2(n7551), .ZN(n7690) );
  XNOR2_X1 U5257 ( .A(n9377), .B(n10507), .ZN(n8495) );
  NOR2_X1 U5258 ( .A1(n7628), .A2(n7633), .ZN(n7627) );
  INV_X1 U5259 ( .A(n9597), .ZN(n9624) );
  AND2_X1 U5260 ( .A1(n7024), .A2(n6547), .ZN(n9626) );
  INV_X1 U5261 ( .A(n8989), .ZN(n10677) );
  NAND2_X1 U5262 ( .A1(n7617), .A2(n10477), .ZN(n10682) );
  AND2_X1 U5263 ( .A1(n10467), .A2(n7527), .ZN(n10528) );
  AND2_X1 U5264 ( .A1(n6590), .A2(n10423), .ZN(n10299) );
  NAND2_X1 U5265 ( .A1(n6027), .A2(n6024), .ZN(n5296) );
  INV_X1 U5266 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6024) );
  NOR2_X1 U5267 ( .A1(n6503), .A2(n6504), .ZN(n6513) );
  XNOR2_X1 U5268 ( .A(n6509), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8532) );
  AND2_X1 U5269 ( .A1(n8868), .A2(n8858), .ZN(n5237) );
  NOR2_X1 U5270 ( .A1(n8209), .A2(n4946), .ZN(n4945) );
  INV_X1 U5271 ( .A(n8215), .ZN(n4946) );
  XNOR2_X1 U5272 ( .A(n8237), .B(n9017), .ZN(n8844) );
  XNOR2_X1 U5273 ( .A(n8946), .B(n7388), .ZN(n7512) );
  OR2_X1 U5274 ( .A1(n5436), .A2(n7104), .ZN(n5448) );
  INV_X1 U5275 ( .A(n5441), .ZN(n5442) );
  OR2_X1 U5276 ( .A1(n4851), .A2(n6676), .ZN(n5405) );
  NOR2_X1 U5277 ( .A1(n8680), .A2(n5956), .ZN(n5038) );
  NAND2_X1 U5278 ( .A1(n8680), .A2(n5037), .ZN(n5036) );
  NOR2_X1 U5279 ( .A1(n10016), .A2(n5183), .ZN(n9969) );
  INV_X1 U5280 ( .A(n5185), .ZN(n5183) );
  OAI22_X1 U5281 ( .A1(n9977), .A2(n8678), .B1(n5955), .B2(n9884), .ZN(n9966)
         );
  NAND2_X1 U5282 ( .A1(n4996), .A2(n8758), .ZN(n4995) );
  INV_X1 U5283 ( .A(n4997), .ZN(n4996) );
  OAI21_X1 U5284 ( .B1(n5057), .B2(n5056), .A(n5054), .ZN(n9977) );
  INV_X1 U5285 ( .A(n5055), .ZN(n5054) );
  OAI22_X1 U5286 ( .A1(n10024), .A2(n5056), .B1(n10026), .B2(n10189), .ZN(
        n5055) );
  NAND2_X1 U5287 ( .A1(n4913), .A2(n5954), .ZN(n5056) );
  NAND2_X1 U5288 ( .A1(n8750), .A2(n8748), .ZN(n10024) );
  NAND2_X1 U5289 ( .A1(n5057), .A2(n10024), .ZN(n10012) );
  AOI21_X1 U5290 ( .B1(n4864), .B2(n5053), .A(n5048), .ZN(n5047) );
  INV_X1 U5291 ( .A(n8612), .ZN(n5048) );
  AOI21_X1 U5292 ( .B1(n5951), .B2(n5052), .A(n4890), .ZN(n5051) );
  INV_X1 U5293 ( .A(n5949), .ZN(n5052) );
  NOR2_X1 U5294 ( .A1(n10205), .A2(n10069), .ZN(n10058) );
  OR2_X1 U5295 ( .A1(n10222), .A2(n9782), .ZN(n10086) );
  AOI21_X1 U5296 ( .B1(n5061), .B2(n5059), .A(n4878), .ZN(n5058) );
  INV_X1 U5297 ( .A(n5061), .ZN(n5060) );
  NOR2_X1 U5298 ( .A1(n10159), .A2(n10226), .ZN(n10125) );
  INV_X1 U5299 ( .A(n4999), .ZN(n4998) );
  AOI21_X1 U5300 ( .B1(n5001), .B2(n8672), .A(n5000), .ZN(n4999) );
  INV_X1 U5301 ( .A(n8705), .ZN(n5000) );
  OR2_X1 U5302 ( .A1(n10231), .A2(n10157), .ZN(n10159) );
  OR2_X1 U5303 ( .A1(n8253), .A2(n8672), .ZN(n8251) );
  NAND2_X1 U5304 ( .A1(n7961), .A2(n4889), .ZN(n8159) );
  NAND2_X1 U5305 ( .A1(n7887), .A2(n5031), .ZN(n8153) );
  NOR2_X1 U5306 ( .A1(n4883), .A2(n5032), .ZN(n5031) );
  INV_X1 U5307 ( .A(n5936), .ZN(n5032) );
  NAND2_X1 U5308 ( .A1(n5580), .A2(n5579), .ZN(n8203) );
  AOI21_X1 U5309 ( .B1(n5929), .B2(n5043), .A(n4897), .ZN(n5042) );
  AND2_X1 U5310 ( .A1(n7084), .A2(n5915), .ZN(n7101) );
  AND2_X1 U5311 ( .A1(n8785), .A2(n5912), .ZN(n7265) );
  AND2_X1 U5312 ( .A1(n7257), .A2(n5360), .ZN(n5166) );
  AND2_X1 U5313 ( .A1(n6712), .A2(n7040), .ZN(n7248) );
  NAND2_X1 U5314 ( .A1(n5898), .A2(n5897), .ZN(n10152) );
  INV_X1 U5315 ( .A(n10111), .ZN(n10146) );
  NAND2_X1 U5316 ( .A1(n8546), .A2(n8545), .ZN(n10176) );
  INV_X1 U5317 ( .A(n7275), .ZN(n10485) );
  INV_X1 U5318 ( .A(n10651), .ZN(n10597) );
  NAND2_X1 U5319 ( .A1(n8287), .A2(n5146), .ZN(n5144) );
  AOI21_X1 U5320 ( .B1(n5146), .B2(n5148), .A(n4924), .ZN(n5143) );
  XNOR2_X1 U5321 ( .A(n5827), .B(n5826), .ZN(n8081) );
  NAND2_X1 U5322 ( .A1(n5787), .A2(n5786), .ZN(n5803) );
  NOR2_X1 U5323 ( .A1(n5259), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n4957) );
  INV_X1 U5324 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5409) );
  XNOR2_X1 U5325 ( .A(n5378), .B(n5358), .ZN(n5377) );
  AND2_X1 U5326 ( .A1(n6407), .A2(n6406), .ZN(n9092) );
  NAND2_X1 U5327 ( .A1(n6244), .A2(n6243), .ZN(n7932) );
  NAND2_X1 U5328 ( .A1(n6315), .A2(n7835), .ZN(n7840) );
  NAND2_X1 U5329 ( .A1(n7737), .A2(n6297), .ZN(n6315) );
  INV_X1 U5330 ( .A(n8140), .ZN(n9714) );
  NAND2_X1 U5331 ( .A1(n6119), .A2(n7478), .ZN(n8964) );
  NAND2_X1 U5332 ( .A1(n6288), .A2(n6287), .ZN(n9718) );
  NAND2_X1 U5333 ( .A1(n4971), .A2(n4970), .ZN(n4969) );
  NAND2_X1 U5334 ( .A1(n4968), .A2(n6483), .ZN(n4967) );
  AND2_X1 U5335 ( .A1(n6344), .A2(n6343), .ZN(n9596) );
  AND2_X1 U5336 ( .A1(n6067), .A2(n6080), .ZN(n10454) );
  INV_X1 U5337 ( .A(n9601), .ZN(n8339) );
  NAND2_X1 U5338 ( .A1(n8301), .A2(n8300), .ZN(n9636) );
  XNOR2_X1 U5339 ( .A(n9422), .B(n5007), .ZN(n9638) );
  INV_X1 U5340 ( .A(n9636), .ZN(n5007) );
  NAND2_X1 U5341 ( .A1(n9448), .A2(n9447), .ZN(n9647) );
  NAND2_X1 U5342 ( .A1(n9443), .A2(n9629), .ZN(n9448) );
  NAND2_X1 U5343 ( .A1(n6026), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U5344 ( .A1(n5862), .A2(n5861), .ZN(n10179) );
  OR2_X1 U5345 ( .A1(n9032), .A2(n9029), .ZN(n9030) );
  NAND2_X1 U5346 ( .A1(n8999), .A2(n9028), .ZN(n9031) );
  AND2_X1 U5347 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  AOI21_X1 U5348 ( .B1(n4954), .B2(n4951), .A(n4949), .ZN(n4948) );
  NAND2_X1 U5349 ( .A1(n5809), .A2(n5808), .ZN(n10196) );
  INV_X1 U5350 ( .A(n7337), .ZN(n10514) );
  NAND2_X1 U5351 ( .A1(n5556), .A2(n5555), .ZN(n8078) );
  OR2_X1 U5352 ( .A1(n8544), .A2(n6604), .ZN(n5383) );
  AND2_X1 U5353 ( .A1(n6891), .A2(n6890), .ZN(n9876) );
  OR2_X1 U5354 ( .A1(n5441), .A2(n5335), .ZN(n5344) );
  OR2_X1 U5355 ( .A1(n5445), .A2(n5340), .ZN(n5341) );
  NAND2_X1 U5356 ( .A1(n6624), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5342) );
  XNOR2_X1 U5357 ( .A(n5350), .B(n5349), .ZN(n6785) );
  AOI21_X1 U5358 ( .B1(n10290), .B2(n8541), .A(n8540), .ZN(n9952) );
  NAND2_X1 U5359 ( .A1(n10160), .A2(n7106), .ZN(n10163) );
  NAND2_X1 U5360 ( .A1(n5067), .A2(n4881), .ZN(n8374) );
  NAND2_X1 U5361 ( .A1(n8408), .A2(n4965), .ZN(n4964) );
  NOR2_X1 U5362 ( .A1(n4966), .A2(n8410), .ZN(n4965) );
  INV_X1 U5363 ( .A(n8406), .ZN(n4966) );
  NAND2_X1 U5364 ( .A1(n4961), .A2(n4959), .ZN(n8435) );
  NOR2_X1 U5365 ( .A1(n7913), .A2(n4960), .ZN(n4959) );
  AOI21_X1 U5366 ( .B1(n4976), .B2(n4975), .A(n4973), .ZN(n8448) );
  INV_X1 U5367 ( .A(n8485), .ZN(n8478) );
  INV_X1 U5368 ( .A(n9843), .ZN(n5244) );
  INV_X1 U5369 ( .A(n5628), .ZN(n5136) );
  INV_X1 U5370 ( .A(n5568), .ZN(n5157) );
  NAND2_X1 U5371 ( .A1(n5508), .A2(n9296), .ZN(n5527) );
  OR2_X1 U5372 ( .A1(n5462), .A2(n5461), .ZN(n5466) );
  INV_X1 U5373 ( .A(n5460), .ZN(n5461) );
  AND2_X1 U5374 ( .A1(n5468), .A2(n5467), .ZN(n5469) );
  INV_X1 U5375 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5114) );
  INV_X1 U5376 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5115) );
  INV_X1 U5377 ( .A(n6400), .ZN(n6399) );
  OR2_X1 U5378 ( .A1(n6448), .A2(n7631), .ZN(n6059) );
  NAND2_X1 U5379 ( .A1(n5094), .A2(n5095), .ZN(n9442) );
  NAND2_X1 U5380 ( .A1(n4904), .A2(n5096), .ZN(n5095) );
  INV_X1 U5381 ( .A(n4873), .ZN(n5096) );
  NOR2_X1 U5382 ( .A1(n5009), .A2(n9650), .ZN(n5008) );
  INV_X1 U5383 ( .A(n5010), .ZN(n5009) );
  AOI21_X1 U5384 ( .B1(n5271), .B2(n5270), .A(n8328), .ZN(n5269) );
  INV_X1 U5385 ( .A(n5273), .ZN(n5270) );
  OAI21_X1 U5386 ( .B1(n5107), .B2(n5108), .A(n8346), .ZN(n5105) );
  NOR2_X1 U5387 ( .A1(n9655), .A2(n5011), .ZN(n5010) );
  INV_X1 U5388 ( .A(n5012), .ZN(n5011) );
  NOR2_X1 U5389 ( .A1(n4871), .A2(n5109), .ZN(n5108) );
  NAND2_X1 U5390 ( .A1(n9538), .A2(n8351), .ZN(n5109) );
  INV_X1 U5391 ( .A(n8454), .ZN(n5075) );
  INV_X1 U5392 ( .A(n9430), .ZN(n5293) );
  AND2_X1 U5393 ( .A1(n5293), .A2(n9582), .ZN(n5290) );
  NOR2_X1 U5394 ( .A1(n10555), .A2(n10544), .ZN(n5019) );
  NAND2_X1 U5395 ( .A1(n5188), .A2(n5187), .ZN(n6019) );
  INV_X1 U5396 ( .A(n6539), .ZN(n5188) );
  NAND2_X1 U5397 ( .A1(n9507), .A2(n9515), .ZN(n9508) );
  AND2_X1 U5398 ( .A1(n7680), .A2(n5015), .ZN(n7711) );
  NOR2_X1 U5399 ( .A1(n10620), .A2(n5017), .ZN(n5015) );
  AND2_X1 U5400 ( .A1(n7604), .A2(n7567), .ZN(n7649) );
  INV_X1 U5401 ( .A(n7650), .ZN(n7570) );
  NOR2_X1 U5402 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n6002) );
  NAND2_X1 U5403 ( .A1(n5999), .A2(n5218), .ZN(n5216) );
  INV_X1 U5404 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5218) );
  OR2_X1 U5405 ( .A1(n6139), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6156) );
  NOR2_X1 U5406 ( .A1(n9767), .A2(n9768), .ZN(n5233) );
  NOR2_X1 U5407 ( .A1(n5233), .A2(n5232), .ZN(n5231) );
  INV_X1 U5408 ( .A(n9856), .ZN(n5232) );
  NOR2_X1 U5409 ( .A1(n5186), .A2(n10179), .ZN(n5185) );
  NAND2_X1 U5410 ( .A1(n9984), .A2(n10189), .ZN(n5186) );
  AOI21_X1 U5411 ( .B1(n5766), .B2(n8614), .A(n8698), .ZN(n4991) );
  NAND2_X1 U5412 ( .A1(n5741), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5759) );
  INV_X1 U5413 ( .A(n5063), .ZN(n5059) );
  NOR2_X1 U5414 ( .A1(n8664), .A2(n5928), .ZN(n5041) );
  INV_X1 U5415 ( .A(n5927), .ZN(n5043) );
  INV_X1 U5416 ( .A(n7265), .ZN(n8651) );
  INV_X1 U5417 ( .A(n8290), .ZN(n5148) );
  INV_X1 U5418 ( .A(n5147), .ZN(n5146) );
  OAI21_X1 U5419 ( .B1(n8286), .B2(n5148), .A(n8291), .ZN(n5147) );
  AND2_X1 U5420 ( .A1(n4882), .A2(n5349), .ZN(n5033) );
  NAND2_X1 U5421 ( .A1(n5594), .A2(n5322), .ZN(n5611) );
  NAND2_X1 U5422 ( .A1(n5260), .A2(n5707), .ZN(n5259) );
  INV_X1 U5423 ( .A(n5309), .ZN(n5260) );
  NOR2_X1 U5424 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(n5611), .ZN(n5228) );
  NAND2_X1 U5425 ( .A1(n5577), .A2(n5553), .ZN(n5578) );
  AOI21_X1 U5426 ( .B1(n5485), .B2(n5152), .A(n5150), .ZN(n5149) );
  INV_X1 U5427 ( .A(n5152), .ZN(n5151) );
  INV_X1 U5428 ( .A(n5506), .ZN(n5150) );
  XNOR2_X1 U5429 ( .A(n5459), .B(SI_6_), .ZN(n5460) );
  NAND2_X1 U5430 ( .A1(n5357), .A2(n6051), .ZN(n5378) );
  NAND2_X1 U5431 ( .A1(n8967), .A2(n5208), .ZN(n10539) );
  NOR2_X1 U5432 ( .A1(n10541), .A2(n5209), .ZN(n5208) );
  INV_X1 U5433 ( .A(n6138), .ZN(n5209) );
  INV_X1 U5434 ( .A(n6370), .ZN(n6369) );
  NAND2_X1 U5435 ( .A1(n7005), .A2(n6073), .ZN(n4930) );
  INV_X1 U5436 ( .A(n8226), .ZN(n6364) );
  INV_X1 U5437 ( .A(n6365), .ZN(n5214) );
  AND2_X1 U5438 ( .A1(n6208), .A2(n6190), .ZN(n5190) );
  AOI21_X1 U5439 ( .B1(n5224), .B2(n5223), .A(n5222), .ZN(n5221) );
  INV_X1 U5440 ( .A(n7951), .ZN(n5222) );
  XNOR2_X1 U5441 ( .A(n5193), .B(n10507), .ZN(n7476) );
  NAND2_X1 U5442 ( .A1(n9098), .A2(n5200), .ZN(n5199) );
  INV_X1 U5443 ( .A(n6438), .ZN(n5200) );
  INV_X1 U5444 ( .A(n10500), .ZN(n10609) );
  OR2_X1 U5445 ( .A1(n7451), .A2(n7449), .ZN(n6557) );
  INV_X1 U5446 ( .A(n8528), .ZN(n4968) );
  NOR2_X1 U5447 ( .A1(n10467), .A2(n8524), .ZN(n4970) );
  AND2_X1 U5448 ( .A1(n5141), .A2(n5140), .ZN(n8525) );
  NAND2_X1 U5449 ( .A1(n8487), .A2(n8488), .ZN(n5140) );
  OAI211_X1 U5450 ( .C1(n8491), .C2(n8485), .A(n8489), .B(n5142), .ZN(n5141)
         );
  NOR4_X1 U5451 ( .A1(n8520), .A2(n8519), .A3(n8518), .A4(n9438), .ZN(n8521)
         );
  AND4_X1 U5452 ( .A1(n6203), .A2(n6202), .A3(n6201), .A4(n6200), .ZN(n7590)
         );
  NOR2_X1 U5453 ( .A1(n6004), .A2(n6005), .ZN(n5219) );
  NAND2_X1 U5454 ( .A1(n8308), .A2(n8307), .ZN(n9645) );
  AND2_X1 U5455 ( .A1(n6499), .A2(n6498), .ZN(n9480) );
  NAND2_X1 U5456 ( .A1(n9501), .A2(n8347), .ZN(n9526) );
  NAND2_X1 U5457 ( .A1(n5025), .A2(n5020), .ZN(n9541) );
  NOR2_X1 U5458 ( .A1(n9589), .A2(n5021), .ZN(n5020) );
  NAND2_X1 U5459 ( .A1(n9554), .A2(n9546), .ZN(n5021) );
  NAND2_X1 U5460 ( .A1(n8322), .A2(n9431), .ZN(n9560) );
  NOR2_X1 U5461 ( .A1(n5022), .A2(n9589), .ZN(n9551) );
  OR2_X1 U5462 ( .A1(n5024), .A2(n9682), .ZN(n5022) );
  NAND2_X1 U5463 ( .A1(n5289), .A2(n5287), .ZN(n9550) );
  NAND2_X1 U5464 ( .A1(n5288), .A2(n5293), .ZN(n5287) );
  NAND2_X1 U5465 ( .A1(n9577), .A2(n5290), .ZN(n5289) );
  INV_X1 U5466 ( .A(n5291), .ZN(n5288) );
  OR2_X1 U5467 ( .A1(n9613), .A2(n9700), .ZN(n9589) );
  NAND2_X1 U5468 ( .A1(n5079), .A2(n5077), .ZN(n9623) );
  AOI21_X1 U5469 ( .B1(n4867), .B2(n5085), .A(n5078), .ZN(n5077) );
  INV_X1 U5470 ( .A(n8363), .ZN(n5078) );
  AND2_X1 U5471 ( .A1(n8310), .A2(n8309), .ZN(n9612) );
  NAND2_X1 U5472 ( .A1(n9612), .A2(n9621), .ZN(n9613) );
  NAND2_X1 U5473 ( .A1(n6324), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6354) );
  OAI21_X1 U5474 ( .B1(n5277), .B2(n5284), .A(n5275), .ZN(n8183) );
  INV_X1 U5475 ( .A(n5284), .ZN(n5276) );
  NOR2_X1 U5476 ( .A1(n8165), .A2(n9714), .ZN(n8309) );
  NAND2_X1 U5477 ( .A1(n8137), .A2(n10677), .ZN(n8167) );
  OR2_X1 U5478 ( .A1(n8167), .A2(n9718), .ZN(n8165) );
  AND2_X1 U5479 ( .A1(n7926), .A2(n10668), .ZN(n8137) );
  NOR2_X1 U5480 ( .A1(n7925), .A2(n7932), .ZN(n7926) );
  OR2_X1 U5481 ( .A1(n6197), .A2(n7234), .ZN(n6215) );
  NAND2_X1 U5482 ( .A1(n5262), .A2(n5261), .ZN(n7578) );
  NAND2_X1 U5483 ( .A1(n7680), .A2(n5019), .ZN(n7664) );
  NAND2_X1 U5484 ( .A1(n5092), .A2(n4863), .ZN(n7662) );
  NAND2_X1 U5485 ( .A1(n7680), .A2(n10547), .ZN(n7682) );
  AND2_X1 U5486 ( .A1(n7648), .A2(n8395), .ZN(n7680) );
  NAND2_X1 U5487 ( .A1(n7557), .A2(n7556), .ZN(n7674) );
  OAI21_X1 U5488 ( .B1(n7690), .B2(n5100), .A(n5098), .ZN(n7557) );
  INV_X1 U5489 ( .A(n5099), .ZN(n5098) );
  NOR2_X1 U5490 ( .A1(n7697), .A2(n7566), .ZN(n7648) );
  OR2_X1 U5491 ( .A1(n7696), .A2(n8382), .ZN(n7697) );
  NAND2_X1 U5492 ( .A1(n7529), .A2(n4854), .ZN(n7628) );
  NAND2_X1 U5493 ( .A1(n6429), .A2(n6428), .ZN(n9670) );
  NAND2_X1 U5494 ( .A1(n6415), .A2(n6414), .ZN(n9676) );
  INV_X1 U5495 ( .A(n8975), .ZN(n10668) );
  AND2_X1 U5496 ( .A1(n7919), .A2(n7912), .ZN(n7914) );
  NAND2_X1 U5497 ( .A1(n5264), .A2(n7586), .ZN(n7588) );
  INV_X1 U5498 ( .A(n5265), .ZN(n5264) );
  AND2_X1 U5499 ( .A1(n7572), .A2(n7571), .ZN(n10531) );
  OR2_X1 U5500 ( .A1(n6866), .A2(P2_U3152), .ZN(n7008) );
  INV_X1 U5501 ( .A(n6005), .ZN(n5217) );
  NOR2_X1 U5502 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5998) );
  NAND2_X1 U5503 ( .A1(n5304), .A2(n6012), .ZN(n6013) );
  INV_X1 U5504 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6021) );
  INV_X1 U5505 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U5506 ( .A1(n7512), .A2(n7511), .ZN(n5250) );
  INV_X1 U5507 ( .A(n5779), .ZN(n5780) );
  NAND2_X1 U5508 ( .A1(n5780), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5792) );
  INV_X1 U5509 ( .A(n9046), .ZN(n9019) );
  OR2_X1 U5510 ( .A1(n9013), .A2(n9012), .ZN(n9029) );
  OR2_X1 U5511 ( .A1(n9011), .A2(n9010), .ZN(n9012) );
  INV_X1 U5512 ( .A(n9832), .ZN(n4949) );
  NAND2_X1 U5513 ( .A1(n9865), .A2(n8855), .ZN(n5238) );
  NAND2_X1 U5514 ( .A1(n5793), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5812) );
  INV_X1 U5515 ( .A(n8925), .ZN(n8922) );
  NAND2_X1 U5516 ( .A1(n7177), .A2(n7176), .ZN(n4955) );
  NAND2_X1 U5517 ( .A1(n4903), .A2(n5248), .ZN(n5247) );
  AOI21_X1 U5518 ( .B1(n5231), .B2(n4953), .A(n4952), .ZN(n4951) );
  NOR2_X1 U5519 ( .A1(n5233), .A2(n5234), .ZN(n4952) );
  NAND2_X1 U5520 ( .A1(n9767), .A2(n9768), .ZN(n5234) );
  NOR2_X1 U5521 ( .A1(n5231), .A2(n5230), .ZN(n4954) );
  NOR2_X1 U5522 ( .A1(n5233), .A2(n8885), .ZN(n5230) );
  OR2_X1 U5523 ( .A1(n5601), .A2(n5600), .ZN(n5618) );
  INV_X1 U5524 ( .A(n5759), .ZN(n5760) );
  NAND2_X1 U5525 ( .A1(n5760), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5779) );
  NOR2_X1 U5526 ( .A1(n5559), .A2(n5558), .ZN(n5581) );
  NAND2_X1 U5527 ( .A1(n8884), .A2(n8885), .ZN(n9857) );
  NAND2_X1 U5528 ( .A1(n9857), .A2(n9856), .ZN(n9855) );
  NOR2_X1 U5529 ( .A1(n5691), .A2(n9850), .ZN(n5714) );
  NOR2_X1 U5530 ( .A1(n5618), .A2(n7437), .ZN(n5637) );
  AND2_X1 U5531 ( .A1(n5637), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5655) );
  INV_X1 U5532 ( .A(n4851), .ZN(n5848) );
  NOR2_X1 U5533 ( .A1(n10016), .A2(n5184), .ZN(n9953) );
  NAND2_X1 U5534 ( .A1(n6580), .A2(n5185), .ZN(n5184) );
  NOR2_X1 U5535 ( .A1(n9986), .A2(n8754), .ZN(n4997) );
  NAND2_X1 U5536 ( .A1(n9993), .A2(n8753), .ZN(n9985) );
  OR2_X1 U5537 ( .A1(n10016), .A2(n5186), .ZN(n9978) );
  NAND2_X1 U5538 ( .A1(n8758), .A2(n8756), .ZN(n9986) );
  NOR2_X1 U5539 ( .A1(n10022), .A2(n5820), .ZN(n9994) );
  INV_X1 U5540 ( .A(n9884), .ZN(n9998) );
  INV_X1 U5541 ( .A(n9885), .ZN(n10026) );
  AOI21_X1 U5542 ( .B1(n4991), .B2(n8744), .A(n4989), .ZN(n4988) );
  INV_X1 U5543 ( .A(n8747), .ZN(n4989) );
  OR2_X1 U5544 ( .A1(n10074), .A2(n4990), .ZN(n4987) );
  INV_X1 U5545 ( .A(n4991), .ZN(n4990) );
  AND2_X1 U5546 ( .A1(n4987), .A2(n4985), .ZN(n10022) );
  NOR2_X1 U5547 ( .A1(n10024), .A2(n4986), .ZN(n4985) );
  INV_X1 U5548 ( .A(n4988), .ZN(n4986) );
  OR2_X1 U5549 ( .A1(n10042), .A2(n10196), .ZN(n10016) );
  AND2_X1 U5550 ( .A1(n8745), .A2(n8747), .ZN(n10035) );
  NOR2_X1 U5551 ( .A1(n10053), .A2(n8744), .ZN(n10034) );
  NOR2_X1 U5552 ( .A1(n10074), .A2(n5766), .ZN(n10053) );
  NAND2_X1 U5553 ( .A1(n5168), .A2(n5167), .ZN(n10069) );
  NAND2_X1 U5554 ( .A1(n10125), .A2(n10106), .ZN(n10100) );
  NAND2_X1 U5555 ( .A1(n10086), .A2(n8604), .ZN(n10109) );
  NAND2_X1 U5556 ( .A1(n8251), .A2(n8687), .ZN(n10144) );
  NAND2_X1 U5557 ( .A1(n5062), .A2(n5061), .ZN(n10142) );
  NAND2_X1 U5558 ( .A1(n5062), .A2(n5065), .ZN(n10140) );
  OR2_X1 U5559 ( .A1(n5674), .A2(n5673), .ZN(n5691) );
  NAND2_X1 U5560 ( .A1(n5655), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U5561 ( .A1(n5177), .A2(n5176), .ZN(n10157) );
  NOR2_X1 U5562 ( .A1(n5178), .A2(n10239), .ZN(n5176) );
  NAND2_X1 U5563 ( .A1(n8103), .A2(n8669), .ZN(n5663) );
  NOR2_X1 U5564 ( .A1(n7967), .A2(n5178), .ZN(n8256) );
  INV_X1 U5565 ( .A(n8669), .ZN(n8104) );
  NOR2_X1 U5566 ( .A1(n7967), .A2(n5179), .ZN(n8155) );
  AND2_X1 U5567 ( .A1(n8730), .A2(n8707), .ZN(n8649) );
  AOI21_X1 U5568 ( .B1(n8665), .B2(n4983), .A(n4982), .ZN(n4981) );
  INV_X1 U5569 ( .A(n8725), .ZN(n4983) );
  AND2_X1 U5570 ( .A1(n7823), .A2(n10652), .ZN(n7890) );
  AND2_X1 U5571 ( .A1(n7640), .A2(n10632), .ZN(n7823) );
  OR2_X1 U5572 ( .A1(n5539), .A2(n5538), .ZN(n5559) );
  OR2_X1 U5573 ( .A1(n5519), .A2(n5518), .ZN(n5539) );
  AOI21_X1 U5574 ( .B1(n7399), .B2(n4992), .A(n5300), .ZN(n7490) );
  NOR2_X1 U5575 ( .A1(n4894), .A2(n4993), .ZN(n4992) );
  INV_X1 U5576 ( .A(n8709), .ZN(n4993) );
  NOR2_X1 U5577 ( .A1(n8044), .A2(n10596), .ZN(n7640) );
  AND4_X1 U5578 ( .A1(n5503), .A2(n5502), .A3(n5501), .A4(n5500), .ZN(n8040)
         );
  NAND2_X1 U5579 ( .A1(n7421), .A2(n4866), .ZN(n8043) );
  AND2_X1 U5580 ( .A1(n7399), .A2(n8709), .ZN(n8037) );
  NAND2_X1 U5581 ( .A1(n7421), .A2(n4865), .ZN(n7756) );
  NAND2_X1 U5582 ( .A1(n7401), .A2(n7400), .ZN(n7399) );
  AND2_X1 U5583 ( .A1(n7421), .A2(n7443), .ZN(n7422) );
  NAND2_X1 U5584 ( .A1(n7100), .A2(n5917), .ZN(n7410) );
  NOR2_X1 U5585 ( .A1(n7105), .A2(n10514), .ZN(n7421) );
  NAND2_X1 U5586 ( .A1(n7269), .A2(n10485), .ZN(n7271) );
  AND2_X1 U5587 ( .A1(n5909), .A2(n5908), .ZN(n6972) );
  OR2_X1 U5588 ( .A1(n6902), .A2(n8776), .ZN(n5907) );
  NAND2_X1 U5589 ( .A1(n6972), .A2(n5910), .ZN(n6971) );
  NOR2_X1 U5590 ( .A1(n6911), .A2(n7256), .ZN(n7269) );
  INV_X1 U5591 ( .A(n5353), .ZN(n4977) );
  NAND2_X1 U5592 ( .A1(n5044), .A2(n5927), .ZN(n7496) );
  NAND2_X1 U5593 ( .A1(n5926), .A2(n4918), .ZN(n5044) );
  XNOR2_X1 U5594 ( .A(n8292), .B(n8291), .ZN(n8542) );
  NAND2_X1 U5595 ( .A1(n5145), .A2(n8290), .ZN(n8292) );
  XNOR2_X1 U5596 ( .A(n8287), .B(n8286), .ZN(n8305) );
  AOI21_X1 U5597 ( .B1(n5842), .B2(n5841), .A(n5840), .ZN(n5858) );
  INV_X1 U5598 ( .A(n5839), .ZN(n5840) );
  NAND2_X1 U5599 ( .A1(n5133), .A2(n5801), .ZN(n5821) );
  AND2_X1 U5600 ( .A1(n5327), .A2(n5551), .ZN(n5174) );
  AOI21_X1 U5601 ( .B1(n4870), .B2(n5130), .A(n5121), .ZN(n5120) );
  INV_X1 U5602 ( .A(n5767), .ZN(n5121) );
  NAND2_X1 U5603 ( .A1(n5123), .A2(n5127), .ZN(n5769) );
  NAND2_X1 U5604 ( .A1(n5125), .A2(n5124), .ZN(n5123) );
  NAND2_X1 U5605 ( .A1(n5126), .A2(n5737), .ZN(n5751) );
  NAND2_X1 U5606 ( .A1(n5137), .A2(n5628), .ZN(n5647) );
  NAND2_X1 U5607 ( .A1(n5610), .A2(n5138), .ZN(n5137) );
  NAND2_X1 U5608 ( .A1(n5158), .A2(n5568), .ZN(n5589) );
  NAND2_X1 U5609 ( .A1(n5547), .A2(n5159), .ZN(n5158) );
  NAND2_X1 U5610 ( .A1(n5547), .A2(n5546), .ZN(n5570) );
  NAND2_X1 U5611 ( .A1(n5154), .A2(n5489), .ZN(n5505) );
  OR2_X1 U5612 ( .A1(n5432), .A2(n5431), .ZN(n5473) );
  NAND2_X1 U5613 ( .A1(n5359), .A2(SI_0_), .ZN(n5366) );
  AND4_X1 U5614 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n10538)
         );
  NAND2_X1 U5615 ( .A1(n8967), .A2(n6138), .ZN(n10540) );
  AND2_X1 U5616 ( .A1(n6470), .A2(n6469), .ZN(n9479) );
  NAND2_X1 U5617 ( .A1(n7374), .A2(n6190), .ZN(n10616) );
  NAND2_X1 U5618 ( .A1(n6364), .A2(n6363), .ZN(n8266) );
  AND4_X1 U5619 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n10557)
         );
  AND4_X1 U5620 ( .A1(n6220), .A2(n6219), .A3(n6218), .A4(n6217), .ZN(n10612)
         );
  NAND2_X1 U5621 ( .A1(n9108), .A2(n6441), .ZN(n9097) );
  NAND2_X1 U5622 ( .A1(n7840), .A2(n6319), .ZN(n7954) );
  AND2_X1 U5623 ( .A1(n6423), .A2(n6422), .ZN(n9558) );
  OR2_X1 U5624 ( .A1(n9106), .A2(n6438), .ZN(n9108) );
  INV_X1 U5625 ( .A(n6870), .ZN(n7032) );
  INV_X1 U5626 ( .A(n10615), .ZN(n10561) );
  NAND2_X1 U5627 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  NAND2_X1 U5628 ( .A1(n5220), .A2(n5221), .ZN(n8088) );
  NAND2_X1 U5629 ( .A1(n6338), .A2(n6337), .ZN(n9703) );
  INV_X1 U5630 ( .A(n9102), .ZN(n9137) );
  NAND2_X1 U5631 ( .A1(n5205), .A2(n5207), .ZN(n5202) );
  NAND2_X1 U5632 ( .A1(n8968), .A2(n6266), .ZN(n5204) );
  AND4_X1 U5633 ( .A1(n6240), .A2(n6239), .A3(n6238), .A4(n6237), .ZN(n8991)
         );
  OR2_X1 U5634 ( .A1(n6109), .A2(n6092), .ZN(n6097) );
  CLKBUF_X1 U5635 ( .A(n6943), .Z(n9379) );
  INV_X1 U5636 ( .A(n10449), .ZN(n10425) );
  AND2_X1 U5637 ( .A1(n7067), .A2(n6547), .ZN(n10455) );
  AOI21_X1 U5638 ( .B1(n9468), .B2(n9629), .A(n9467), .ZN(n9653) );
  AND2_X1 U5639 ( .A1(n9482), .A2(n8472), .ZN(n9466) );
  NAND2_X1 U5640 ( .A1(n5268), .A2(n5271), .ZN(n9472) );
  NAND2_X1 U5641 ( .A1(n9499), .A2(n5273), .ZN(n5268) );
  NAND2_X1 U5642 ( .A1(n6461), .A2(n6460), .ZN(n9661) );
  NAND2_X1 U5643 ( .A1(n8081), .A2(n8304), .ZN(n6461) );
  AOI21_X1 U5644 ( .B1(n9499), .B2(n9435), .A(n9434), .ZN(n9487) );
  NAND2_X1 U5645 ( .A1(n5076), .A2(n8454), .ZN(n9569) );
  NAND2_X1 U5646 ( .A1(n9576), .A2(n5307), .ZN(n9565) );
  NAND2_X1 U5647 ( .A1(n5081), .A2(n5082), .ZN(n8316) );
  OR2_X1 U5648 ( .A1(n8172), .A2(n5085), .ZN(n5081) );
  NAND2_X1 U5649 ( .A1(n5086), .A2(n8441), .ZN(n8190) );
  OR2_X1 U5650 ( .A1(n8172), .A2(n8146), .ZN(n5086) );
  AND2_X1 U5651 ( .A1(n6303), .A2(n6302), .ZN(n8140) );
  NAND2_X1 U5652 ( .A1(n5279), .A2(n5280), .ZN(n8135) );
  AND2_X1 U5653 ( .A1(n5277), .A2(n5279), .ZN(n8181) );
  NOR2_X1 U5654 ( .A1(n8133), .A2(n5283), .ZN(n8164) );
  NAND2_X1 U5655 ( .A1(n6274), .A2(n6273), .ZN(n8989) );
  AND2_X1 U5656 ( .A1(n7913), .A2(n7912), .ZN(n5298) );
  AND2_X1 U5657 ( .A1(n7910), .A2(n7909), .ZN(n7920) );
  NAND2_X1 U5658 ( .A1(n7606), .A2(n7554), .ZN(n7655) );
  OAI22_X1 U5659 ( .A1(n6366), .A2(n6594), .B1(n7074), .B2(n6593), .ZN(n5069)
         );
  INV_X1 U5660 ( .A(n5004), .ZN(n5003) );
  OAI22_X1 U5661 ( .A1(n6104), .A2(n6596), .B1(n7074), .B2(n7071), .ZN(n5004)
         );
  NAND2_X1 U5662 ( .A1(n10299), .A2(n7455), .ZN(n9592) );
  INV_X1 U5663 ( .A(n9620), .ZN(n9606) );
  CLKBUF_X1 U5664 ( .A(n9517), .Z(n9457) );
  OAI21_X1 U5665 ( .B1(n9638), .B2(n10678), .A(n9637), .ZN(n9723) );
  NOR2_X1 U5666 ( .A1(n9647), .A2(n5110), .ZN(n9648) );
  NAND2_X1 U5667 ( .A1(n5301), .A2(n4911), .ZN(n5110) );
  INV_X1 U5668 ( .A(n5296), .ZN(n5295) );
  NAND2_X1 U5669 ( .A1(n6507), .A2(n6026), .ZN(n8083) );
  NAND2_X1 U5670 ( .A1(n5777), .A2(n5776), .ZN(n10205) );
  NAND2_X1 U5671 ( .A1(n9855), .A2(n9859), .ZN(n9770) );
  NAND2_X1 U5672 ( .A1(n5713), .A2(n5712), .ZN(n10226) );
  CLKBUF_X1 U5673 ( .A(n7811), .Z(n7945) );
  NAND2_X1 U5674 ( .A1(n5238), .A2(n8858), .ZN(n9800) );
  NAND2_X1 U5675 ( .A1(n7335), .A2(n5235), .ZN(n7348) );
  NOR2_X1 U5676 ( .A1(n5236), .A2(n7341), .ZN(n5235) );
  INV_X1 U5677 ( .A(n7334), .ZN(n5236) );
  NAND2_X1 U5678 ( .A1(n5790), .A2(n5789), .ZN(n10201) );
  NAND2_X1 U5679 ( .A1(n4955), .A2(n7181), .ZN(n7184) );
  NAND2_X1 U5680 ( .A1(n5727), .A2(n5726), .ZN(n10222) );
  NAND2_X1 U5681 ( .A1(n4943), .A2(n8833), .ZN(n4942) );
  INV_X1 U5682 ( .A(n4945), .ZN(n4943) );
  NAND2_X1 U5683 ( .A1(n5599), .A2(n5598), .ZN(n10261) );
  NAND2_X1 U5684 ( .A1(n5245), .A2(n9777), .ZN(n9841) );
  NAND2_X1 U5685 ( .A1(n5239), .A2(n5246), .ZN(n5245) );
  INV_X1 U5686 ( .A(n9776), .ZN(n5239) );
  AND2_X1 U5687 ( .A1(n8822), .A2(n6923), .ZN(n9873) );
  NAND2_X1 U5688 ( .A1(n8886), .A2(n4953), .ZN(n9859) );
  INV_X1 U5689 ( .A(n8884), .ZN(n8886) );
  OR2_X1 U5690 ( .A1(n8763), .A2(n8641), .ZN(n8642) );
  NAND4_X1 U5691 ( .A1(n5484), .A2(n5483), .A3(n5482), .A4(n5481), .ZN(n9897)
         );
  NAND4_X1 U5692 ( .A1(n5450), .A2(n5449), .A3(n5448), .A4(n5447), .ZN(n9899)
         );
  OR2_X1 U5693 ( .A1(n5883), .A2(n7168), .ZN(n5387) );
  OR2_X1 U5694 ( .A1(n5436), .A2(n6660), .ZN(n5407) );
  NOR2_X1 U5695 ( .A1(n5306), .A2(n5406), .ZN(n5408) );
  OR2_X1 U5696 ( .A1(n5441), .A2(n5368), .ZN(n5371) );
  NAND2_X1 U5697 ( .A1(n6624), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5370) );
  OR2_X1 U5698 ( .A1(n4850), .A2(n6673), .ZN(n5369) );
  OR2_X1 U5699 ( .A1(n5403), .A2(n6713), .ZN(n5365) );
  AND2_X1 U5700 ( .A1(n5452), .A2(n5392), .ZN(n6784) );
  INV_X1 U5701 ( .A(n10176), .ZN(n9954) );
  NAND2_X1 U5702 ( .A1(n8680), .A2(n9959), .ZN(n5039) );
  OAI21_X1 U5703 ( .B1(n8680), .B2(n4900), .A(n5036), .ZN(n5035) );
  NAND2_X1 U5704 ( .A1(n10012), .A2(n5954), .ZN(n9996) );
  NAND2_X1 U5705 ( .A1(n5049), .A2(n5051), .ZN(n10064) );
  NAND2_X1 U5706 ( .A1(n5050), .A2(n5951), .ZN(n5049) );
  NAND2_X1 U5707 ( .A1(n5950), .A2(n5949), .ZN(n10068) );
  NAND2_X1 U5708 ( .A1(n5690), .A2(n5689), .ZN(n10231) );
  NAND2_X1 U5709 ( .A1(n5942), .A2(n5941), .ZN(n8250) );
  AND2_X1 U5710 ( .A1(n7961), .A2(n8731), .ZN(n5299) );
  NAND2_X1 U5711 ( .A1(n5931), .A2(n4893), .ZN(n10648) );
  NAND2_X1 U5712 ( .A1(n7637), .A2(n8663), .ZN(n4984) );
  AND2_X1 U5713 ( .A1(n5455), .A2(n5454), .ZN(n7337) );
  OR2_X1 U5714 ( .A1(n8544), .A2(n6608), .ZN(n5413) );
  OR2_X1 U5715 ( .A1(n10600), .A2(n6570), .ZN(n10160) );
  AND2_X1 U5716 ( .A1(n10163), .A2(n6576), .ZN(n10137) );
  NAND2_X1 U5717 ( .A1(n10181), .A2(n5960), .ZN(n10182) );
  XNOR2_X1 U5718 ( .A(n8299), .B(n8298), .ZN(n10290) );
  NAND2_X1 U5719 ( .A1(n5144), .A2(n5143), .ZN(n8299) );
  XNOR2_X1 U5720 ( .A(n5875), .B(n5874), .ZN(n8195) );
  XNOR2_X1 U5721 ( .A(n5858), .B(n5857), .ZN(n8111) );
  XNOR2_X1 U5722 ( .A(n5896), .B(n5257), .ZN(n7486) );
  INV_X1 U5723 ( .A(n6784), .ZN(n6677) );
  NOR2_X1 U5724 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5373) );
  CLKBUF_X1 U5725 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n10292) );
  NAND2_X1 U5726 ( .A1(n5118), .A2(n7023), .ZN(n5116) );
  INV_X1 U5727 ( .A(n5005), .ZN(P2_U3519) );
  AOI21_X1 U5728 ( .B1(n9723), .B2(n10689), .A(n5006), .ZN(n5005) );
  NOR2_X1 U5729 ( .A1(n10689), .A2(n6691), .ZN(n5006) );
  AOI21_X1 U5730 ( .B1(n9033), .B2(n9032), .A(n9050), .ZN(n9038) );
  AND2_X1 U5731 ( .A1(n8502), .A2(n8400), .ZN(n4863) );
  INV_X1 U5732 ( .A(n8522), .ZN(n5187) );
  AND2_X1 U5733 ( .A1(n5051), .A2(n4896), .ZN(n4864) );
  AND2_X1 U5734 ( .A1(n7406), .A2(n7443), .ZN(n4865) );
  AND2_X1 U5735 ( .A1(n4865), .A2(n5182), .ZN(n4866) );
  AND2_X1 U5736 ( .A1(n5082), .A2(n5080), .ZN(n4867) );
  INV_X1 U5737 ( .A(n5272), .ZN(n5271) );
  OAI22_X1 U5738 ( .A1(n9490), .A2(n5274), .B1(n9436), .B2(n9661), .ZN(n5272)
         );
  INV_X1 U5739 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6515) );
  AND2_X1 U5740 ( .A1(n8723), .A2(n8720), .ZN(n8664) );
  AND2_X1 U5741 ( .A1(n8728), .A2(n8725), .ZN(n8663) );
  INV_X1 U5742 ( .A(n8663), .ZN(n4980) );
  NAND2_X1 U5743 ( .A1(n6384), .A2(n6383), .ZN(n9687) );
  AND2_X1 U5744 ( .A1(n7789), .A2(n5251), .ZN(n4868) );
  AND2_X1 U5745 ( .A1(n4866), .A2(n5181), .ZN(n4869) );
  AND2_X1 U5746 ( .A1(n5127), .A2(n5122), .ZN(n4870) );
  NOR2_X1 U5747 ( .A1(n9667), .A2(n9133), .ZN(n9434) );
  NOR2_X1 U5748 ( .A1(n9589), .A2(n5024), .ZN(n5023) );
  INV_X1 U5749 ( .A(n8990), .ZN(n5207) );
  NOR2_X1 U5750 ( .A1(n9435), .A2(n9501), .ZN(n4871) );
  AND2_X1 U5751 ( .A1(n6086), .A2(n5999), .ZN(n6088) );
  NAND2_X1 U5752 ( .A1(n5408), .A2(n5407), .ZN(n6892) );
  NAND2_X1 U5753 ( .A1(n4947), .A2(n4945), .ZN(n8233) );
  INV_X2 U5754 ( .A(n5445), .ZN(n5361) );
  AND2_X1 U5755 ( .A1(n5046), .A2(n5047), .ZN(n4872) );
  AND2_X1 U5756 ( .A1(n9650), .A2(n9480), .ZN(n4873) );
  INV_X1 U5757 ( .A(n5225), .ZN(n5224) );
  OR2_X1 U5758 ( .A1(n7950), .A2(n5226), .ZN(n5225) );
  NOR2_X1 U5759 ( .A1(n9687), .A2(n9557), .ZN(n4874) );
  OR2_X1 U5760 ( .A1(n5646), .A2(n5136), .ZN(n4875) );
  OR2_X1 U5761 ( .A1(n5588), .A2(n5157), .ZN(n4876) );
  OR2_X1 U5762 ( .A1(n5955), .A2(n9998), .ZN(n8758) );
  AND3_X1 U5763 ( .A1(n5374), .A2(n5229), .A3(n5352), .ZN(n5390) );
  XNOR2_X1 U5764 ( .A(n9700), .B(n9428), .ZN(n9602) );
  INV_X1 U5765 ( .A(n9602), .ZN(n4974) );
  NAND2_X1 U5766 ( .A1(n6398), .A2(n6397), .ZN(n9682) );
  NAND2_X1 U5767 ( .A1(n5424), .A2(n5423), .ZN(n5464) );
  NAND2_X1 U5768 ( .A1(n5636), .A2(n5635), .ZN(n10249) );
  INV_X1 U5769 ( .A(n8364), .ZN(n5080) );
  AND4_X1 U5770 ( .A1(n6012), .A2(n6023), .A3(n6535), .A4(n6505), .ZN(n4877)
         );
  INV_X1 U5771 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U5772 ( .A1(n8997), .A2(n6035), .ZN(n6093) );
  AND2_X1 U5773 ( .A1(n10231), .A2(n10121), .ZN(n4878) );
  AND2_X1 U5774 ( .A1(n7743), .A2(n6284), .ZN(n4879) );
  AND2_X1 U5775 ( .A1(n6063), .A2(n5998), .ZN(n6086) );
  OR2_X1 U5776 ( .A1(n6104), .A2(n6605), .ZN(n4880) );
  OR2_X1 U5777 ( .A1(n8478), .A2(n8368), .ZN(n4881) );
  NAND2_X1 U5778 ( .A1(n9031), .A2(n9030), .ZN(n9050) );
  NOR2_X1 U5779 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4882) );
  NAND2_X1 U5780 ( .A1(n6443), .A2(n6442), .ZN(n9667) );
  NAND2_X1 U5781 ( .A1(n9488), .A2(n8463), .ZN(n9435) );
  NOR2_X1 U5782 ( .A1(n10257), .A2(n9890), .ZN(n4883) );
  AND2_X1 U5783 ( .A1(n9560), .A2(n8351), .ZN(n4884) );
  AND2_X1 U5784 ( .A1(n9993), .A2(n4997), .ZN(n4885) );
  AND2_X1 U5785 ( .A1(n5202), .A2(n7742), .ZN(n4886) );
  AND2_X1 U5786 ( .A1(n5925), .A2(n5041), .ZN(n4887) );
  OR2_X1 U5787 ( .A1(n7803), .A2(n5249), .ZN(n4888) );
  NAND2_X1 U5788 ( .A1(n6543), .A2(n6542), .ZN(n9650) );
  NAND2_X1 U5789 ( .A1(n5672), .A2(n5671), .ZN(n10239) );
  AND2_X1 U5790 ( .A1(n5644), .A2(n8731), .ZN(n4889) );
  AND2_X1 U5791 ( .A1(n10211), .A2(n10055), .ZN(n4890) );
  NAND2_X1 U5792 ( .A1(n9507), .A2(n5010), .ZN(n5013) );
  NAND2_X1 U5793 ( .A1(n9507), .A2(n5012), .ZN(n5014) );
  INV_X1 U5794 ( .A(n5023), .ZN(n5027) );
  OR2_X1 U5795 ( .A1(n6366), .A2(n6591), .ZN(n4891) );
  AND2_X1 U5796 ( .A1(n7569), .A2(n7649), .ZN(n4892) );
  INV_X1 U5797 ( .A(n9431), .ZN(n9555) );
  AND2_X1 U5798 ( .A1(n8351), .A2(n8350), .ZN(n9431) );
  AND2_X1 U5799 ( .A1(n5932), .A2(n5930), .ZN(n4893) );
  INV_X1 U5800 ( .A(n5951), .ZN(n5053) );
  NAND2_X1 U5801 ( .A1(n8708), .A2(n8721), .ZN(n4894) );
  AND4_X1 U5802 ( .A1(n5304), .A2(n6022), .A3(n6508), .A4(n6021), .ZN(n4895)
         );
  NAND2_X1 U5803 ( .A1(n10205), .A2(n10037), .ZN(n4896) );
  NOR2_X1 U5804 ( .A1(n10596), .A2(n9894), .ZN(n4897) );
  NAND2_X1 U5805 ( .A1(n8472), .A2(n8471), .ZN(n9477) );
  INV_X1 U5806 ( .A(n9477), .ZN(n8328) );
  OR2_X1 U5807 ( .A1(n5706), .A2(n5309), .ZN(n4898) );
  OR2_X1 U5808 ( .A1(n8504), .A2(n7591), .ZN(n4899) );
  INV_X1 U5809 ( .A(n5213), .ZN(n5212) );
  OAI21_X1 U5810 ( .B1(n6363), .B2(n5214), .A(n8264), .ZN(n5213) );
  AND2_X1 U5811 ( .A1(n9965), .A2(n5037), .ZN(n4900) );
  XNOR2_X1 U5812 ( .A(n5488), .B(SI_7_), .ZN(n5485) );
  INV_X1 U5813 ( .A(n8208), .ZN(n8209) );
  AND2_X1 U5814 ( .A1(n8729), .A2(n8706), .ZN(n8665) );
  INV_X1 U5815 ( .A(n8665), .ZN(n5932) );
  INV_X1 U5816 ( .A(n9434), .ZN(n5274) );
  NAND3_X1 U5817 ( .A1(n5174), .A2(n5172), .A3(n5552), .ZN(n4901) );
  AND4_X1 U5818 ( .A1(n5217), .A2(n4877), .A3(n6027), .A4(n6086), .ZN(n4902)
         );
  INV_X1 U5819 ( .A(n5017), .ZN(n5016) );
  NAND2_X1 U5820 ( .A1(n5019), .A2(n5018), .ZN(n5017) );
  INV_X1 U5821 ( .A(n5286), .ZN(n5283) );
  NAND2_X1 U5822 ( .A1(n10677), .A2(n8970), .ZN(n5286) );
  INV_X1 U5823 ( .A(n5025), .ZN(n5024) );
  NOR2_X1 U5824 ( .A1(n9687), .A2(n9692), .ZN(n5025) );
  NAND2_X1 U5825 ( .A1(n5197), .A2(n5196), .ZN(n9096) );
  INV_X1 U5826 ( .A(n9098), .ZN(n5201) );
  AND2_X1 U5827 ( .A1(n8352), .A2(n9525), .ZN(n9538) );
  OR2_X1 U5828 ( .A1(n7791), .A2(n7941), .ZN(n4903) );
  NAND2_X1 U5829 ( .A1(n9465), .A2(n8472), .ZN(n4904) );
  NAND2_X1 U5830 ( .A1(n5654), .A2(n5653), .ZN(n10246) );
  AND2_X1 U5831 ( .A1(n8758), .A2(n9995), .ZN(n4905) );
  AND2_X1 U5832 ( .A1(n8210), .A2(n8833), .ZN(n4906) );
  AND2_X1 U5833 ( .A1(n5227), .A2(n5221), .ZN(n4907) );
  AND2_X1 U5834 ( .A1(n5295), .A2(n6033), .ZN(n4908) );
  AND2_X1 U5835 ( .A1(n7804), .A2(n5250), .ZN(n4909) );
  AND2_X1 U5836 ( .A1(n5282), .A2(n5276), .ZN(n4910) );
  INV_X1 U5837 ( .A(n8655), .ZN(n5918) );
  AND2_X1 U5838 ( .A1(n8551), .A2(n8789), .ZN(n8655) );
  INV_X1 U5839 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5257) );
  INV_X1 U5840 ( .A(n8885), .ZN(n4953) );
  NAND2_X1 U5841 ( .A1(n5847), .A2(n5846), .ZN(n5955) );
  OAI21_X1 U5842 ( .B1(n6364), .B2(n5214), .A(n5212), .ZN(n8268) );
  NAND2_X1 U5843 ( .A1(n4939), .A2(n9085), .ZN(n9088) );
  NAND2_X1 U5844 ( .A1(n6017), .A2(n6021), .ZN(n6503) );
  AND2_X1 U5845 ( .A1(n5577), .A2(n4958), .ZN(n5652) );
  AND3_X1 U5846 ( .A1(n5217), .A2(n5215), .A3(n6086), .ZN(n6300) );
  NAND2_X1 U5847 ( .A1(n4944), .A2(n4942), .ZN(n8845) );
  NAND2_X1 U5848 ( .A1(n7887), .A2(n5936), .ZN(n7960) );
  OR2_X1 U5849 ( .A1(n9454), .A2(n10676), .ZN(n4911) );
  AND2_X1 U5850 ( .A1(n5577), .A2(n5228), .ZN(n5614) );
  INV_X1 U5851 ( .A(n9777), .ZN(n5243) );
  NAND2_X1 U5852 ( .A1(n5830), .A2(n5829), .ZN(n10007) );
  NAND2_X1 U5853 ( .A1(n5219), .A2(n6088), .ZN(n6298) );
  NAND2_X1 U5854 ( .A1(n10007), .A2(n10026), .ZN(n8753) );
  OR2_X1 U5855 ( .A1(n10588), .A2(n10557), .ZN(n8407) );
  INV_X1 U5856 ( .A(n5168), .ZN(n10084) );
  NOR2_X1 U5857 ( .A1(n10217), .A2(n10100), .ZN(n5168) );
  INV_X1 U5858 ( .A(n9959), .ZN(n9965) );
  NAND2_X1 U5859 ( .A1(n8628), .A2(n8757), .ZN(n9959) );
  INV_X1 U5860 ( .A(n5130), .ZN(n5124) );
  NAND2_X1 U5861 ( .A1(n5749), .A2(n5737), .ZN(n5130) );
  NAND2_X1 U5862 ( .A1(n6477), .A2(n6476), .ZN(n9655) );
  AND2_X1 U5863 ( .A1(n9576), .A2(n5291), .ZN(n4912) );
  OR2_X1 U5864 ( .A1(n10007), .A2(n9885), .ZN(n4913) );
  AND2_X1 U5865 ( .A1(n5750), .A2(SI_21_), .ZN(n4914) );
  AND2_X1 U5866 ( .A1(n5698), .A2(SI_18_), .ZN(n4915) );
  INV_X1 U5867 ( .A(n5164), .ZN(n5163) );
  NAND2_X1 U5868 ( .A1(n5165), .A2(n5696), .ZN(n5164) );
  AND2_X1 U5869 ( .A1(n9476), .A2(n9142), .ZN(n4916) );
  NAND2_X1 U5870 ( .A1(n5881), .A2(n5880), .ZN(n5963) );
  AND2_X1 U5871 ( .A1(n8251), .A2(n5001), .ZN(n4917) );
  INV_X1 U5872 ( .A(n9778), .ZN(n5246) );
  AND2_X1 U5873 ( .A1(n8906), .A2(n8907), .ZN(n9778) );
  AND2_X1 U5874 ( .A1(n5894), .A2(n5893), .ZN(n5958) );
  INV_X1 U5875 ( .A(n9687), .ZN(n5026) );
  INV_X1 U5876 ( .A(n7835), .ZN(n5223) );
  NAND2_X1 U5877 ( .A1(n7919), .A2(n5298), .ZN(n7973) );
  NAND2_X1 U5878 ( .A1(n5204), .A2(n8990), .ZN(n7741) );
  NAND2_X1 U5879 ( .A1(n4984), .A2(n8725), .ZN(n7821) );
  NAND2_X1 U5880 ( .A1(n4956), .A2(n5250), .ZN(n7802) );
  NAND2_X1 U5881 ( .A1(n5757), .A2(n5756), .ZN(n10211) );
  INV_X1 U5882 ( .A(n10211), .ZN(n5167) );
  NAND2_X1 U5883 ( .A1(n5931), .A2(n5930), .ZN(n7828) );
  AND2_X1 U5884 ( .A1(n5925), .A2(n5045), .ZN(n4918) );
  NOR2_X1 U5885 ( .A1(n7967), .A2(n10257), .ZN(n5180) );
  AND2_X1 U5886 ( .A1(n8425), .A2(n8426), .ZN(n8508) );
  NAND2_X1 U5887 ( .A1(n8037), .A2(n8708), .ZN(n4919) );
  AND2_X1 U5888 ( .A1(n7680), .A2(n5016), .ZN(n4920) );
  AND2_X1 U5889 ( .A1(n7690), .A2(n7553), .ZN(n4921) );
  AND2_X1 U5890 ( .A1(n5823), .A2(n5801), .ZN(n4922) );
  AND2_X1 U5891 ( .A1(n5092), .A2(n8400), .ZN(n4923) );
  INV_X1 U5892 ( .A(n10581), .ZN(n5181) );
  INV_X1 U5893 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5112) );
  OAI21_X1 U5894 ( .B1(n6937), .B2(n6936), .A(n6917), .ZN(n7177) );
  INV_X1 U5895 ( .A(n8277), .ZN(n5182) );
  NAND2_X1 U5896 ( .A1(n6176), .A2(n6175), .ZN(n10588) );
  INV_X1 U5897 ( .A(n10588), .ZN(n5018) );
  XNOR2_X1 U5898 ( .A(n6054), .B(n6055), .ZN(n7013) );
  AND2_X1 U5899 ( .A1(n8294), .A2(n9258), .ZN(n4924) );
  OR2_X1 U5900 ( .A1(n8534), .A2(n8533), .ZN(n4925) );
  INV_X1 U5901 ( .A(n8340), .ZN(n5195) );
  AND2_X1 U5902 ( .A1(n5195), .A2(n7023), .ZN(n4926) );
  INV_X1 U5903 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8127) );
  INV_X2 U5904 ( .A(n10289), .ZN(n9064) );
  NAND2_X1 U5905 ( .A1(n4927), .A2(n9650), .ZN(n6565) );
  NAND2_X1 U5906 ( .A1(n4928), .A2(n6546), .ZN(n4927) );
  NAND2_X1 U5907 ( .A1(n6544), .A2(n10561), .ZN(n4928) );
  XNOR2_X1 U5908 ( .A(n6502), .B(n6501), .ZN(n6544) );
  INV_X1 U5909 ( .A(n6084), .ZN(n7045) );
  NAND2_X1 U5910 ( .A1(n4930), .A2(n10494), .ZN(n7044) );
  NAND2_X1 U5911 ( .A1(n6072), .A2(n4931), .ZN(n7005) );
  INV_X1 U5912 ( .A(n7006), .ZN(n4931) );
  NAND2_X1 U5913 ( .A1(n4935), .A2(n9066), .ZN(n9069) );
  NAND2_X1 U5914 ( .A1(n9065), .A2(n6475), .ZN(n4935) );
  NAND2_X1 U5915 ( .A1(n4936), .A2(n9127), .ZN(n9065) );
  NAND2_X1 U5916 ( .A1(n5198), .A2(n4937), .ZN(n4936) );
  INV_X1 U5917 ( .A(n4938), .ZN(n4937) );
  OAI21_X1 U5918 ( .B1(n9106), .B2(n5199), .A(n6459), .ZN(n4938) );
  NAND2_X1 U5919 ( .A1(n7737), .A2(n4940), .ZN(n5220) );
  NAND2_X1 U5920 ( .A1(n5220), .A2(n4907), .ZN(n6349) );
  NAND2_X1 U5921 ( .A1(n8211), .A2(n4906), .ZN(n4944) );
  NAND2_X1 U5922 ( .A1(n8211), .A2(n8210), .ZN(n4947) );
  AND2_X1 U5923 ( .A1(n4947), .A2(n8208), .ZN(n8214) );
  OAI21_X1 U5924 ( .B1(n8884), .B2(n4954), .A(n4951), .ZN(n9834) );
  NAND2_X1 U5925 ( .A1(n4950), .A2(n4948), .ZN(n8900) );
  NAND2_X1 U5926 ( .A1(n8884), .A2(n4951), .ZN(n4950) );
  NAND2_X1 U5927 ( .A1(n7513), .A2(n5251), .ZN(n4956) );
  NAND2_X1 U5928 ( .A1(n4956), .A2(n4909), .ZN(n7806) );
  NAND3_X1 U5929 ( .A1(n5577), .A2(n4958), .A3(n5651), .ZN(n5706) );
  NAND3_X1 U5930 ( .A1(n5577), .A2(n4958), .A3(n4957), .ZN(n5895) );
  INV_X1 U5931 ( .A(n6015), .ZN(n6017) );
  NAND2_X1 U5932 ( .A1(n6300), .A2(n6023), .ZN(n6014) );
  NAND3_X1 U5933 ( .A1(n8526), .A2(n4969), .A3(n4967), .ZN(n5118) );
  NAND3_X1 U5934 ( .A1(n9610), .A2(n8447), .A3(n4974), .ZN(n4973) );
  NAND3_X1 U5935 ( .A1(n8443), .A2(n8513), .A3(n8442), .ZN(n4976) );
  NAND2_X2 U5936 ( .A1(n4977), .A2(n5360), .ZN(n8776) );
  NAND2_X1 U5937 ( .A1(n5166), .A2(n4977), .ZN(n7256) );
  NAND2_X1 U5938 ( .A1(n7637), .A2(n4979), .ZN(n4978) );
  NAND2_X1 U5939 ( .A1(n4978), .A2(n4981), .ZN(n7885) );
  NAND2_X1 U5940 ( .A1(n4987), .A2(n4988), .ZN(n10023) );
  NAND2_X1 U5941 ( .A1(n8159), .A2(n8736), .ZN(n8103) );
  INV_X1 U5942 ( .A(n8658), .ZN(n7400) );
  INV_X1 U5943 ( .A(n5458), .ZN(n7401) );
  NAND2_X1 U5944 ( .A1(n4994), .A2(n4995), .ZN(n9960) );
  NAND2_X1 U5945 ( .A1(n9994), .A2(n4905), .ZN(n4994) );
  NAND2_X1 U5946 ( .A1(n9994), .A2(n9995), .ZN(n9993) );
  AOI21_X1 U5947 ( .B1(n8253), .B2(n5001), .A(n4998), .ZN(n10119) );
  NAND2_X1 U5948 ( .A1(n9507), .A2(n5008), .ZN(n9449) );
  INV_X1 U5949 ( .A(n5014), .ZN(n9493) );
  INV_X1 U5950 ( .A(n5013), .ZN(n9473) );
  NOR2_X1 U5951 ( .A1(n9589), .A2(n9692), .ZN(n5028) );
  INV_X1 U5952 ( .A(n5028), .ZN(n9578) );
  NAND2_X1 U5953 ( .A1(n10648), .A2(n5933), .ZN(n7889) );
  NAND4_X1 U5954 ( .A1(n5171), .A2(n5170), .A3(n5175), .A4(n4882), .ZN(n5348)
         );
  NAND3_X1 U5955 ( .A1(n5171), .A2(n5170), .A3(n5175), .ZN(n5966) );
  NOR2_X1 U5956 ( .A1(n9966), .A2(n9965), .ZN(n9964) );
  INV_X1 U5957 ( .A(n6584), .ZN(n5961) );
  OAI211_X1 U5958 ( .C1(n9966), .C2(n5039), .A(n5034), .B(n5035), .ZN(n6584)
         );
  NAND2_X1 U5959 ( .A1(n9966), .A2(n5038), .ZN(n5034) );
  NAND2_X1 U5960 ( .A1(n5926), .A2(n4887), .ZN(n5040) );
  NAND2_X1 U5961 ( .A1(n5040), .A2(n5042), .ZN(n7639) );
  NAND2_X1 U5962 ( .A1(n5926), .A2(n5925), .ZN(n8042) );
  INV_X1 U5963 ( .A(n5928), .ZN(n5045) );
  INV_X1 U5964 ( .A(n5950), .ZN(n5050) );
  NAND2_X1 U5965 ( .A1(n5950), .A2(n4864), .ZN(n5046) );
  XNOR2_X2 U5966 ( .A(n6902), .B(n8776), .ZN(n7251) );
  INV_X1 U5967 ( .A(n5550), .ZN(n5175) );
  OR2_X1 U5968 ( .A1(n5919), .A2(n7749), .ZN(n5921) );
  NAND4_X1 U5969 ( .A1(n6226), .A2(n6227), .A3(n6270), .A4(n5066), .ZN(n6004)
         );
  INV_X1 U5970 ( .A(n6952), .ZN(n6953) );
  OAI21_X1 U5971 ( .B1(n6952), .B2(n7619), .A(n7618), .ZN(n10483) );
  NAND2_X1 U5972 ( .A1(n7621), .A2(n6952), .ZN(n7622) );
  OR2_X1 U5973 ( .A1(n8369), .A2(n6952), .ZN(n5067) );
  INV_X1 U5974 ( .A(n5069), .ZN(n5068) );
  NAND2_X1 U5975 ( .A1(n5072), .A2(n4902), .ZN(n5073) );
  NAND2_X1 U5976 ( .A1(n5070), .A2(n5072), .ZN(n6026) );
  AND2_X1 U5977 ( .A1(n5071), .A2(n5217), .ZN(n5070) );
  NAND2_X1 U5978 ( .A1(n9583), .A2(n8319), .ZN(n5076) );
  NAND2_X1 U5979 ( .A1(n8172), .A2(n4867), .ZN(n5079) );
  NAND2_X1 U5980 ( .A1(n7674), .A2(n4863), .ZN(n5089) );
  NAND2_X1 U5981 ( .A1(n5089), .A2(n5090), .ZN(n7560) );
  XNOR2_X1 U5982 ( .A(n9442), .B(n9441), .ZN(n9443) );
  NAND2_X1 U5983 ( .A1(n8329), .A2(n5097), .ZN(n5094) );
  NAND2_X1 U5984 ( .A1(n8329), .A2(n8328), .ZN(n9482) );
  NAND2_X2 U5985 ( .A1(n5113), .A2(n5111), .ZN(n5359) );
  NAND3_X1 U5986 ( .A1(n5112), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5111) );
  NAND3_X1 U5987 ( .A1(n8127), .A2(n5115), .A3(n5114), .ZN(n5113) );
  NAND2_X1 U5988 ( .A1(n8529), .A2(n4926), .ZN(n5117) );
  NAND3_X1 U5989 ( .A1(n5117), .A2(n5116), .A3(n4925), .ZN(P2_U3244) );
  NAND2_X1 U5990 ( .A1(n5119), .A2(n5120), .ZN(n5774) );
  NAND2_X1 U5991 ( .A1(n5736), .A2(n4870), .ZN(n5119) );
  NAND2_X1 U5992 ( .A1(n5736), .A2(n5735), .ZN(n5126) );
  INV_X1 U5993 ( .A(n5736), .ZN(n5125) );
  NAND2_X1 U5994 ( .A1(n5133), .A2(n4922), .ZN(n5842) );
  NAND2_X1 U5995 ( .A1(n5610), .A2(n5609), .ZN(n5630) );
  NAND2_X1 U5996 ( .A1(n5665), .A2(n5664), .ZN(n5667) );
  NAND2_X1 U5997 ( .A1(n8287), .A2(n8286), .ZN(n5145) );
  NAND2_X1 U5998 ( .A1(n5487), .A2(n5486), .ZN(n5154) );
  OAI21_X2 U5999 ( .B1(n5547), .B2(n4876), .A(n5155), .ZN(n5608) );
  OAI21_X1 U6000 ( .B1(n5683), .B2(n5682), .A(n5685), .ZN(n5697) );
  NAND2_X1 U6001 ( .A1(n5682), .A2(n5685), .ZN(n5165) );
  AND3_X1 U6002 ( .A1(n5325), .A2(n5326), .A3(n5987), .ZN(n5172) );
  NAND4_X1 U6003 ( .A1(n5174), .A2(n5552), .A3(n5326), .A4(n5325), .ZN(n5173)
         );
  INV_X1 U6004 ( .A(n7967), .ZN(n5177) );
  INV_X1 U6005 ( .A(n5180), .ZN(n8156) );
  NAND2_X1 U6006 ( .A1(n4869), .A2(n7421), .ZN(n8044) );
  NOR2_X1 U6007 ( .A1(n10016), .A2(n10007), .ZN(n10003) );
  NAND2_X1 U6008 ( .A1(n7044), .A2(n6100), .ZN(n7050) );
  NAND2_X1 U6009 ( .A1(n9088), .A2(n6409), .ZN(n9115) );
  XNOR2_X2 U6010 ( .A(n5189), .B(n6010), .ZN(n7527) );
  NAND2_X1 U6011 ( .A1(n5192), .A2(n5191), .ZN(n6054) );
  NAND2_X1 U6012 ( .A1(n5194), .A2(n6020), .ZN(n5191) );
  NAND2_X1 U6013 ( .A1(n6020), .A2(n8340), .ZN(n5193) );
  NAND2_X1 U6014 ( .A1(n7013), .A2(n7015), .ZN(n7014) );
  NAND2_X1 U6015 ( .A1(n9106), .A2(n6441), .ZN(n5196) );
  AOI21_X1 U6016 ( .B1(n6441), .B2(n6438), .A(n5201), .ZN(n5197) );
  NAND2_X1 U6017 ( .A1(n8968), .A2(n5205), .ZN(n5203) );
  NAND2_X2 U6018 ( .A1(n5203), .A2(n4886), .ZN(n7737) );
  NAND2_X1 U6019 ( .A1(n6134), .A2(n8960), .ZN(n8967) );
  NOR2_X1 U6020 ( .A1(n6004), .A2(n5216), .ZN(n5215) );
  INV_X2 U6021 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6022 ( .A1(n7335), .A2(n7334), .ZN(n7342) );
  NAND2_X1 U6023 ( .A1(n5238), .A2(n5237), .ZN(n9797) );
  OAI21_X1 U6024 ( .B1(n9776), .B2(n5240), .A(n5241), .ZN(n8926) );
  AOI21_X1 U6025 ( .B1(n7513), .B2(n4868), .A(n5247), .ZN(n7810) );
  NAND2_X1 U6026 ( .A1(n5652), .A2(n5255), .ZN(n5254) );
  NAND2_X1 U6027 ( .A1(n7578), .A2(n8505), .ZN(n7716) );
  NAND2_X1 U6028 ( .A1(n5265), .A2(n7577), .ZN(n5261) );
  NAND2_X1 U6029 ( .A1(n5263), .A2(n7669), .ZN(n5262) );
  AND2_X1 U6030 ( .A1(n7576), .A2(n7577), .ZN(n5263) );
  NAND2_X1 U6031 ( .A1(n7669), .A2(n7576), .ZN(n7586) );
  NAND3_X1 U6032 ( .A1(n7572), .A2(n7571), .A3(n8393), .ZN(n7678) );
  NAND2_X1 U6033 ( .A1(n9499), .A2(n5269), .ZN(n5267) );
  NAND2_X1 U6034 ( .A1(n8133), .A2(n4910), .ZN(n5275) );
  INV_X1 U6035 ( .A(n6026), .ZN(n5294) );
  NAND2_X1 U6036 ( .A1(n5294), .A2(n4908), .ZN(n9742) );
  NOR2_X1 U6037 ( .A1(n6026), .A2(n5296), .ZN(n6032) );
  NAND2_X2 U6038 ( .A1(n5336), .A2(n5339), .ZN(n5445) );
  NAND2_X1 U6039 ( .A1(n8332), .A2(n9643), .ZN(n8333) );
  NAND2_X1 U6040 ( .A1(n8321), .A2(n8320), .ZN(n9556) );
  NOR2_X1 U6041 ( .A1(n10194), .A2(n6896), .ZN(n10000) );
  NAND2_X1 U6042 ( .A1(n5842), .A2(n5838), .ZN(n5827) );
  NAND2_X1 U6043 ( .A1(n5875), .A2(n5874), .ZN(n5879) );
  NAND2_X1 U6044 ( .A1(n5961), .A2(n5960), .ZN(n5965) );
  NAND2_X1 U6045 ( .A1(n4859), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6046 ( .A1(n7560), .A2(n7559), .ZN(n7705) );
  NAND2_X1 U6047 ( .A1(n8338), .A2(n8342), .ZN(n8528) );
  AND2_X1 U6048 ( .A1(n7810), .A2(n7812), .ZN(n7809) );
  NAND2_X1 U6049 ( .A1(n6263), .A2(n6262), .ZN(n8968) );
  OR2_X1 U6050 ( .A1(n6868), .A2(n5187), .ZN(n6020) );
  CLKBUF_X1 U6051 ( .A(n6539), .Z(n8530) );
  NAND2_X1 U6052 ( .A1(n5774), .A2(n5773), .ZN(n5787) );
  NAND2_X1 U6053 ( .A1(n8926), .A2(n8925), .ZN(n9759) );
  NAND2_X1 U6054 ( .A1(n8927), .A2(n9759), .ZN(n8999) );
  NAND2_X1 U6055 ( .A1(n5390), .A2(n5328), .ZN(n5550) );
  OAI21_X1 U6056 ( .B1(n8845), .B2(n8844), .A(n8843), .ZN(n8848) );
  OAI22_X1 U6057 ( .A1(n8544), .A2(n6597), .B1(n6646), .B2(n6672), .ZN(n5353)
         );
  INV_X1 U6058 ( .A(n5451), .ZN(n5463) );
  XNOR2_X1 U6059 ( .A(n5821), .B(n5822), .ZN(n8054) );
  AOI22_X1 U6060 ( .A1(n9611), .A2(n9622), .B1(n9621), .B2(n9596), .ZN(n9603)
         );
  OAI21_X1 U6061 ( .B1(n10119), .B2(n10132), .A(n8699), .ZN(n10108) );
  INV_X1 U6062 ( .A(n5339), .ZN(n5337) );
  AOI22_X1 U6063 ( .A1(n9460), .A2(n9438), .B1(n9464), .B2(n9480), .ZN(n9439)
         );
  INV_X1 U6064 ( .A(n5336), .ZN(n5338) );
  INV_X1 U6065 ( .A(n6038), .ZN(n8997) );
  NOR2_X2 U6066 ( .A1(n7974), .A2(n8510), .ZN(n8133) );
  NOR2_X1 U6067 ( .A1(n5525), .A2(n8719), .ZN(n5300) );
  OR2_X1 U6068 ( .A1(n9646), .A2(n10678), .ZN(n5301) );
  OR2_X1 U6069 ( .A1(n6574), .A2(n4856), .ZN(n5302) );
  OR2_X1 U6070 ( .A1(n6584), .A2(n10134), .ZN(n5303) );
  INV_X1 U6071 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5329) );
  AND2_X1 U6072 ( .A1(n8788), .A2(n8714), .ZN(n8653) );
  INV_X1 U6073 ( .A(n8653), .ZN(n5916) );
  INV_X1 U6074 ( .A(n8668), .ZN(n5644) );
  AND2_X1 U6075 ( .A1(n4860), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5306) );
  AND2_X1 U6076 ( .A1(n8530), .A2(n10467), .ZN(n10554) );
  INV_X1 U6077 ( .A(n9594), .ZN(n9629) );
  OR2_X1 U6078 ( .A1(n9429), .A2(n9428), .ZN(n5308) );
  NAND3_X1 U6079 ( .A1(n5705), .A2(n5704), .A3(n5703), .ZN(n5309) );
  OR2_X1 U6080 ( .A1(n10656), .A2(n5996), .ZN(n5310) );
  OR2_X1 U6081 ( .A1(n4855), .A2(n5882), .ZN(n5311) );
  AND2_X1 U6082 ( .A1(n6896), .A2(n10600), .ZN(n10580) );
  INV_X1 U6083 ( .A(n9370), .ZN(n9143) );
  NAND4_X2 U6084 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n6914)
         );
  AND2_X1 U6085 ( .A1(n5609), .A2(n5593), .ZN(n5312) );
  AND2_X1 U6086 ( .A1(n5527), .A2(n5510), .ZN(n5313) );
  AND2_X1 U6087 ( .A1(n6454), .A2(n6453), .ZN(n9528) );
  INV_X1 U6088 ( .A(n10024), .ZN(n10015) );
  INV_X1 U6089 ( .A(n8649), .ZN(n5934) );
  INV_X1 U6090 ( .A(n8495), .ZN(n7551) );
  NOR2_X1 U6091 ( .A1(n8206), .A2(n8207), .ZN(n5315) );
  AND2_X1 U6092 ( .A1(n5324), .A2(n5323), .ZN(n5325) );
  INV_X1 U6093 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5322) );
  INV_X1 U6094 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6012) );
  INV_X1 U6095 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5999) );
  INV_X1 U6096 ( .A(n6245), .ZN(n6234) );
  INV_X1 U6097 ( .A(n6325), .ZN(n6324) );
  INV_X1 U6098 ( .A(n7185), .ZN(n7182) );
  INV_X1 U6099 ( .A(n7941), .ZN(n7807) );
  NAND2_X1 U6100 ( .A1(n8629), .A2(n8810), .ZN(n8680) );
  AND2_X1 U6101 ( .A1(n10179), .A2(n9883), .ZN(n5956) );
  INV_X1 U6102 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U6103 ( .A1(n6973), .A2(n8778), .ZN(n7264) );
  INV_X1 U6104 ( .A(n5822), .ZN(n5823) );
  INV_X1 U6105 ( .A(n5485), .ZN(n5486) );
  OR2_X1 U6106 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  AND2_X1 U6107 ( .A1(n6489), .A2(n6488), .ZN(n9066) );
  NAND2_X1 U6108 ( .A1(n6234), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6247) );
  OR2_X1 U6109 ( .A1(n6416), .A2(n9247), .ZN(n6430) );
  INV_X1 U6110 ( .A(n10617), .ZN(n6208) );
  AND2_X1 U6111 ( .A1(n6475), .A2(n6474), .ZN(n9127) );
  OR2_X1 U6112 ( .A1(n6307), .A2(n6306), .ZN(n6325) );
  INV_X1 U6113 ( .A(n6856), .ZN(n6160) );
  OR2_X1 U6114 ( .A1(n6093), .A2(n6058), .ZN(n6060) );
  AND2_X1 U6115 ( .A1(n7208), .A2(n7159), .ZN(n7160) );
  AND2_X1 U6116 ( .A1(n6493), .A2(n6548), .ZN(n9462) );
  NAND2_X1 U6117 ( .A1(n6214), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6245) );
  AND3_X1 U6118 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n6128) );
  INV_X1 U6119 ( .A(n8508), .ZN(n7911) );
  INV_X1 U6120 ( .A(n9799), .ZN(n8868) );
  AOI22_X1 U6121 ( .A1(n6914), .A2(n6912), .B1(n8234), .B2(n6911), .ZN(n6913)
         );
  INV_X1 U6122 ( .A(n5792), .ZN(n5793) );
  INV_X1 U6123 ( .A(n8680), .ZN(n5957) );
  NAND2_X1 U6124 ( .A1(n8780), .A2(n8778), .ZN(n5910) );
  INV_X1 U6125 ( .A(n9883), .ZN(n9987) );
  INV_X1 U6126 ( .A(n10035), .ZN(n5952) );
  NAND2_X1 U6127 ( .A1(n5858), .A2(n5857), .ZN(n5860) );
  NAND2_X1 U6128 ( .A1(n5608), .A2(n5312), .ZN(n5610) );
  NAND2_X1 U6129 ( .A1(n5530), .A2(n5529), .ZN(n5546) );
  INV_X1 U6130 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6144) );
  OR2_X1 U6131 ( .A1(n6179), .A2(n6178), .ZN(n6197) );
  INV_X1 U6132 ( .A(n10621), .ZN(n6546) );
  OR2_X1 U6133 ( .A1(n6385), .A2(n9334), .ZN(n6400) );
  OR2_X1 U6134 ( .A1(n6430), .A2(n9110), .ZN(n6446) );
  OR2_X1 U6135 ( .A1(n6557), .A2(n6556), .ZN(n9102) );
  INV_X1 U6136 ( .A(n6692), .ZN(n6857) );
  OR2_X1 U6137 ( .A1(n6109), .A2(n6127), .ZN(n6133) );
  OR2_X1 U6138 ( .A1(n7206), .A2(n7205), .ZN(n7208) );
  AND2_X1 U6139 ( .A1(n7214), .A2(n7138), .ZN(n7140) );
  AND2_X1 U6140 ( .A1(n6437), .A2(n6436), .ZN(n9107) );
  AND2_X1 U6141 ( .A1(n8340), .A2(n8490), .ZN(n9594) );
  NOR2_X1 U6142 ( .A1(n8083), .A2(n6520), .ZN(n10297) );
  INV_X1 U6143 ( .A(n6300), .ZN(n6320) );
  NAND2_X1 U6144 ( .A1(n8195), .A2(n8541), .ZN(n5862) );
  NAND2_X1 U6145 ( .A1(n8999), .A2(n9826), .ZN(n9787) );
  NAND2_X1 U6146 ( .A1(n8081), .A2(n8541), .ZN(n5830) );
  AND2_X1 U6147 ( .A1(n5728), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5741) );
  AND2_X1 U6148 ( .A1(n5714), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5728) );
  AND2_X1 U6149 ( .A1(n9966), .A2(n9965), .ZN(n9967) );
  INV_X1 U6150 ( .A(n10038), .ZN(n9997) );
  INV_X1 U6151 ( .A(n5910), .ZN(n6974) );
  INV_X1 U6152 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5996) );
  AND2_X1 U6153 ( .A1(n8751), .A2(n8753), .ZN(n9995) );
  OR2_X1 U6154 ( .A1(n8645), .A2(n6920), .ZN(n10111) );
  NOR2_X1 U6155 ( .A1(n6145), .A2(n6144), .ZN(n6161) );
  AND2_X1 U6156 ( .A1(n10570), .A2(n10554), .ZN(n10621) );
  INV_X1 U6157 ( .A(n6448), .ZN(n6553) );
  AND4_X1 U6158 ( .A1(n6294), .A2(n6293), .A3(n6292), .A4(n6291), .ZN(n8134)
         );
  AND4_X1 U6159 ( .A1(n6252), .A2(n6251), .A3(n6250), .A4(n6249), .ZN(n8976)
         );
  OR2_X1 U6160 ( .A1(n7212), .A2(n7211), .ZN(n7214) );
  INV_X1 U6161 ( .A(n10554), .ZN(n10676) );
  NOR2_X1 U6162 ( .A1(n9539), .A2(n9538), .ZN(n9681) );
  INV_X1 U6163 ( .A(n10682), .ZN(n10666) );
  AND2_X1 U6164 ( .A1(n8537), .A2(n8522), .ZN(n10467) );
  AND2_X1 U6165 ( .A1(n6850), .A2(n6724), .ZN(n9853) );
  AOI21_X1 U6166 ( .B1(n8644), .B2(n8643), .A(n8642), .ZN(n8772) );
  INV_X2 U6167 ( .A(n5428), .ZN(n8541) );
  NOR2_X1 U6168 ( .A1(n9964), .A2(n9967), .ZN(n10181) );
  INV_X1 U6169 ( .A(n10149), .ZN(n10120) );
  OR2_X1 U6170 ( .A1(n6852), .A2(n8816), .ZN(n10633) );
  OR2_X1 U6171 ( .A1(n8631), .A2(n8816), .ZN(n10600) );
  AND2_X1 U6172 ( .A1(n5993), .A2(n5992), .ZN(n6567) );
  XNOR2_X1 U6173 ( .A(n5421), .B(SI_4_), .ZN(n5419) );
  INV_X1 U6174 ( .A(n9143), .ZN(P2_U3966) );
  INV_X1 U6175 ( .A(n10455), .ZN(n10426) );
  INV_X1 U6176 ( .A(n10685), .ZN(n10684) );
  INV_X1 U6177 ( .A(n10689), .ZN(n10686) );
  OR2_X1 U6178 ( .A1(n6518), .A2(n6517), .ZN(n8055) );
  AOI21_X1 U6179 ( .B1(n6582), .B2(n10137), .A(n6581), .ZN(n6585) );
  AND2_X1 U6180 ( .A1(n10155), .A2(n10154), .ZN(n10237) );
  AND2_X1 U6181 ( .A1(n6885), .A2(n6586), .ZN(n10295) );
  NOR2_X1 U6182 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5321) );
  AND3_X1 U6183 ( .A1(n5321), .A2(n5320), .A3(n5319), .ZN(n5327) );
  INV_X1 U6184 ( .A(n5611), .ZN(n5326) );
  NOR2_X1 U6185 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5324) );
  NOR2_X1 U6186 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5328) );
  INV_X1 U6187 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5346) );
  INV_X1 U6188 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6189 ( .A1(n5332), .A2(n5333), .ZN(n10285) );
  INV_X1 U6190 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5331) );
  XNOR2_X2 U6191 ( .A(n5334), .B(n5333), .ZN(n5339) );
  INV_X1 U6192 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5335) );
  INV_X1 U6193 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6671) );
  INV_X1 U6194 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5340) );
  NAND4_X4 U6195 ( .A1(n5344), .A2(n5343), .A3(n5342), .A4(n5341), .ZN(n6902)
         );
  XNOR2_X2 U6196 ( .A(n5347), .B(n5346), .ZN(n5899) );
  NAND2_X1 U6197 ( .A1(n5348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5350) );
  INV_X1 U6198 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5349) );
  INV_X2 U6199 ( .A(n5359), .ZN(n5356) );
  INV_X4 U6200 ( .A(n5356), .ZN(n8295) );
  INV_X1 U6201 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6597) );
  INV_X1 U6202 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6203 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n10292), .ZN(n5351) );
  XNOR2_X1 U6204 ( .A(n5352), .B(n5351), .ZN(n6672) );
  INV_X1 U6205 ( .A(n5366), .ZN(n5354) );
  NAND2_X1 U6206 ( .A1(n5354), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5357) );
  AND2_X1 U6207 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6208 ( .A1(n5356), .A2(n5355), .ZN(n6051) );
  INV_X1 U6209 ( .A(SI_1_), .ZN(n5358) );
  MUX2_X1 U6210 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5359), .Z(n5376) );
  XNOR2_X1 U6211 ( .A(n5377), .B(n5376), .ZN(n6596) );
  OR2_X1 U6212 ( .A1(n5428), .A2(n6596), .ZN(n5360) );
  INV_X1 U6213 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6713) );
  INV_X1 U6214 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6727) );
  OR2_X1 U6215 ( .A1(n5441), .A2(n6727), .ZN(n5364) );
  NAND2_X1 U6216 ( .A1(n6624), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5363) );
  NAND4_X2 U6217 ( .A1(n5365), .A2(n5364), .A3(n5363), .A4(n5362), .ZN(n6712)
         );
  XNOR2_X1 U6218 ( .A(n5366), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10293) );
  MUX2_X1 U6219 ( .A(n10292), .B(n10293), .S(n6646), .Z(n7040) );
  INV_X1 U6220 ( .A(n7040), .ZN(n7257) );
  NOR2_X1 U6221 ( .A1(n6712), .A2(n7257), .ZN(n7252) );
  INV_X1 U6222 ( .A(n8776), .ZN(n10472) );
  OR2_X1 U6223 ( .A1(n6902), .A2(n10472), .ZN(n5367) );
  NAND2_X1 U6224 ( .A1(n7250), .A2(n5367), .ZN(n8782) );
  NAND2_X1 U6225 ( .A1(n4860), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5372) );
  INV_X1 U6226 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5368) );
  INV_X1 U6227 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6673) );
  OR2_X1 U6228 ( .A1(n5373), .A2(n5331), .ZN(n5375) );
  XNOR2_X1 U6229 ( .A(n5375), .B(n5374), .ZN(n6791) );
  INV_X1 U6230 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U6231 ( .A1(n5377), .A2(n5376), .ZN(n5380) );
  NAND2_X1 U6232 ( .A1(n5378), .A2(SI_1_), .ZN(n5379) );
  NAND2_X1 U6233 ( .A1(n5380), .A2(n5379), .ZN(n5394) );
  MUX2_X1 U6234 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5359), .Z(n5395) );
  INV_X1 U6235 ( .A(SI_2_), .ZN(n5381) );
  XNOR2_X1 U6236 ( .A(n5395), .B(n5381), .ZN(n5393) );
  XNOR2_X1 U6237 ( .A(n5394), .B(n5393), .ZN(n6605) );
  OR2_X1 U6238 ( .A1(n5428), .A2(n6605), .ZN(n5382) );
  OAI211_X2 U6239 ( .C1(n6646), .C2(n6791), .A(n5383), .B(n5382), .ZN(n6911)
         );
  NAND2_X1 U6240 ( .A1(n6914), .A2(n7326), .ZN(n8780) );
  NAND2_X1 U6241 ( .A1(n8782), .A2(n6974), .ZN(n6973) );
  NAND2_X1 U6242 ( .A1(n4860), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5389) );
  INV_X1 U6243 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5384) );
  OR2_X1 U6244 ( .A1(n4851), .A2(n5384), .ZN(n5388) );
  XNOR2_X1 U6245 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7168) );
  INV_X2 U6246 ( .A(n6624), .ZN(n5436) );
  INV_X1 U6247 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5385) );
  OR2_X1 U6248 ( .A1(n5436), .A2(n5385), .ZN(n5386) );
  NAND2_X1 U6249 ( .A1(n5390), .A2(n5409), .ZN(n5432) );
  NAND2_X1 U6250 ( .A1(n5432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5391) );
  INV_X1 U6251 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6252 ( .A1(n5391), .A2(n5430), .ZN(n5452) );
  OR2_X1 U6253 ( .A1(n5391), .A2(n5430), .ZN(n5392) );
  NAND2_X1 U6254 ( .A1(n5394), .A2(n5393), .ZN(n5397) );
  NAND2_X1 U6255 ( .A1(n5395), .A2(SI_2_), .ZN(n5396) );
  NAND2_X1 U6256 ( .A1(n5397), .A2(n5396), .ZN(n5412) );
  MUX2_X1 U6257 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5359), .Z(n5398) );
  INV_X1 U6258 ( .A(SI_3_), .ZN(n9308) );
  XNOR2_X1 U6259 ( .A(n5398), .B(n9308), .ZN(n5411) );
  NAND2_X1 U6260 ( .A1(n5412), .A2(n5411), .ZN(n5400) );
  NAND2_X1 U6261 ( .A1(n5398), .A2(SI_3_), .ZN(n5399) );
  INV_X1 U6262 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6595) );
  INV_X1 U6263 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6606) );
  MUX2_X1 U6264 ( .A(n6595), .B(n6606), .S(n8295), .Z(n5421) );
  XNOR2_X1 U6265 ( .A(n5420), .B(n5419), .ZN(n6607) );
  OR2_X1 U6266 ( .A1(n6607), .A2(n5428), .ZN(n5402) );
  OR2_X1 U6267 ( .A1(n8544), .A2(n6606), .ZN(n5401) );
  OAI211_X1 U6268 ( .C1(n6646), .C2(n6677), .A(n5402), .B(n5401), .ZN(n7175)
         );
  INV_X1 U6269 ( .A(n7175), .ZN(n7318) );
  NAND2_X1 U6270 ( .A1(n9900), .A2(n7318), .ZN(n5914) );
  INV_X1 U6271 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6676) );
  OR2_X1 U6272 ( .A1(n5441), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6273 ( .A1(n5405), .A2(n5404), .ZN(n5406) );
  INV_X1 U6274 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6660) );
  OR2_X1 U6275 ( .A1(n5390), .A2(n5331), .ZN(n5410) );
  XNOR2_X1 U6276 ( .A(n5410), .B(n5409), .ZN(n6748) );
  XNOR2_X1 U6277 ( .A(n5412), .B(n5411), .ZN(n6609) );
  OR2_X1 U6278 ( .A1(n5428), .A2(n6609), .ZN(n5414) );
  INV_X1 U6279 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6608) );
  OAI211_X1 U6280 ( .C1(n6646), .C2(n6748), .A(n5414), .B(n5413), .ZN(n7275)
         );
  NAND2_X1 U6281 ( .A1(n6892), .A2(n10485), .ZN(n5912) );
  AND2_X1 U6282 ( .A1(n5914), .A2(n5912), .ZN(n8783) );
  NAND2_X1 U6283 ( .A1(n7264), .A2(n8783), .ZN(n5418) );
  INV_X1 U6284 ( .A(n8785), .ZN(n5415) );
  NAND2_X1 U6285 ( .A1(n5415), .A2(n5914), .ZN(n5416) );
  OR2_X1 U6286 ( .A1(n9900), .A2(n7318), .ZN(n8787) );
  AND2_X1 U6287 ( .A1(n5416), .A2(n8787), .ZN(n5417) );
  NAND2_X1 U6288 ( .A1(n5418), .A2(n5417), .ZN(n7102) );
  NAND2_X1 U6289 ( .A1(n5420), .A2(n5419), .ZN(n5424) );
  INV_X1 U6290 ( .A(n5421), .ZN(n5422) );
  NAND2_X1 U6291 ( .A1(n5422), .A2(SI_4_), .ZN(n5423) );
  MUX2_X1 U6292 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8295), .Z(n5425) );
  NAND2_X1 U6293 ( .A1(n5464), .A2(n5463), .ZN(n5426) );
  NAND2_X1 U6294 ( .A1(n5425), .A2(SI_5_), .ZN(n5468) );
  NAND2_X1 U6295 ( .A1(n5426), .A2(n5468), .ZN(n5427) );
  MUX2_X1 U6296 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5359), .Z(n5459) );
  XNOR2_X1 U6297 ( .A(n5427), .B(n5460), .ZN(n6610) );
  NAND2_X1 U6298 ( .A1(n6610), .A2(n8541), .ZN(n5435) );
  INV_X1 U6299 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6300 ( .A1(n5430), .A2(n5429), .ZN(n5431) );
  NAND2_X1 U6301 ( .A1(n5473), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5433) );
  XNOR2_X1 U6302 ( .A(n5433), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U6303 ( .A1(n5711), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5710), .B2(
        n10379), .ZN(n5434) );
  NAND2_X1 U6304 ( .A1(n5435), .A2(n5434), .ZN(n7424) );
  NAND2_X1 U6305 ( .A1(n4860), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5440) );
  INV_X1 U6306 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6669) );
  OR2_X1 U6307 ( .A1(n4851), .A2(n6669), .ZN(n5439) );
  OAI21_X1 U6308 ( .B1(n5443), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5479), .ZN(
        n7442) );
  OR2_X1 U6309 ( .A1(n5883), .A2(n7442), .ZN(n5438) );
  OR2_X1 U6310 ( .A1(n5436), .A2(n6656), .ZN(n5437) );
  INV_X1 U6311 ( .A(n9898), .ZN(n5456) );
  NAND2_X1 U6312 ( .A1(n7424), .A2(n5456), .ZN(n8789) );
  AOI21_X1 U6313 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5444) );
  NOR2_X1 U6314 ( .A1(n5444), .A2(n5443), .ZN(n7107) );
  NAND2_X1 U6315 ( .A1(n5442), .A2(n7107), .ZN(n5450) );
  INV_X1 U6316 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6670) );
  OR2_X1 U6317 ( .A1(n4851), .A2(n6670), .ZN(n5449) );
  INV_X1 U6318 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7104) );
  INV_X1 U6319 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5446) );
  OR2_X1 U6320 ( .A1(n5445), .A2(n5446), .ZN(n5447) );
  XNOR2_X1 U6321 ( .A(n5464), .B(n5451), .ZN(n6600) );
  NAND2_X1 U6322 ( .A1(n6600), .A2(n8541), .ZN(n5455) );
  NAND2_X1 U6323 ( .A1(n5452), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5453) );
  XNOR2_X1 U6324 ( .A(n5453), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10405) );
  AOI22_X1 U6325 ( .A1(n5711), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5710), .B2(
        n10405), .ZN(n5454) );
  OR2_X1 U6326 ( .A1(n9899), .A2(n7337), .ZN(n8788) );
  NAND2_X1 U6327 ( .A1(n8789), .A2(n8788), .ZN(n8715) );
  OR2_X1 U6328 ( .A1(n5456), .A2(n7424), .ZN(n8551) );
  NAND2_X1 U6329 ( .A1(n9899), .A2(n7337), .ZN(n8714) );
  NAND2_X1 U6330 ( .A1(n8551), .A2(n8714), .ZN(n5457) );
  NAND2_X1 U6331 ( .A1(n5457), .A2(n8789), .ZN(n8790) );
  OAI21_X1 U6332 ( .B1(n7102), .B2(n8715), .A(n8790), .ZN(n5458) );
  NAND2_X1 U6333 ( .A1(n5459), .A2(SI_6_), .ZN(n5467) );
  INV_X1 U6334 ( .A(n5467), .ZN(n5462) );
  NAND2_X1 U6335 ( .A1(n5465), .A2(n5464), .ZN(n5472) );
  INV_X1 U6336 ( .A(n5466), .ZN(n5470) );
  MUX2_X1 U6337 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8295), .Z(n5488) );
  XNOR2_X1 U6338 ( .A(n5487), .B(n5485), .ZN(n6614) );
  NAND2_X1 U6339 ( .A1(n6614), .A2(n8541), .ZN(n5476) );
  NOR2_X1 U6340 ( .A1(n5473), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5494) );
  OR2_X1 U6341 ( .A1(n5494), .A2(n5331), .ZN(n5474) );
  XNOR2_X1 U6342 ( .A(n5474), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6762) );
  AOI22_X1 U6343 ( .A1(n5711), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5710), .B2(
        n6762), .ZN(n5475) );
  NAND2_X1 U6344 ( .A1(n5476), .A2(n5475), .ZN(n7523) );
  NAND2_X1 U6345 ( .A1(n4860), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5484) );
  INV_X1 U6346 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5477) );
  OR2_X1 U6347 ( .A1(n4851), .A2(n5477), .ZN(n5483) );
  AND2_X1 U6348 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  NOR2_X2 U6349 ( .A1(n5479), .A2(n5478), .ZN(n5497) );
  OR2_X1 U6350 ( .A1(n5480), .A2(n5497), .ZN(n7521) );
  OR2_X1 U6351 ( .A1(n5883), .A2(n7521), .ZN(n5482) );
  INV_X1 U6352 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7403) );
  OR2_X1 U6353 ( .A1(n5436), .A2(n7403), .ZN(n5481) );
  INV_X1 U6354 ( .A(n9897), .ZN(n7413) );
  OR2_X1 U6355 ( .A1(n7523), .A2(n7413), .ZN(n8791) );
  NAND2_X1 U6356 ( .A1(n7523), .A2(n7413), .ZN(n8709) );
  NAND2_X1 U6357 ( .A1(n8791), .A2(n8709), .ZN(n8658) );
  NAND2_X1 U6358 ( .A1(n5488), .A2(SI_7_), .ZN(n5489) );
  INV_X1 U6359 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6618) );
  INV_X1 U6360 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6619) );
  MUX2_X1 U6361 ( .A(n6618), .B(n6619), .S(n8295), .Z(n5490) );
  INV_X1 U6362 ( .A(SI_8_), .ZN(n9300) );
  INV_X1 U6363 ( .A(n5490), .ZN(n5491) );
  NAND2_X1 U6364 ( .A1(n5491), .A2(SI_8_), .ZN(n5492) );
  XNOR2_X1 U6365 ( .A(n5505), .B(n5504), .ZN(n6617) );
  NAND2_X1 U6366 ( .A1(n6617), .A2(n8541), .ZN(n5496) );
  INV_X1 U6367 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U6368 ( .A1(n5494), .A2(n5493), .ZN(n5533) );
  NAND2_X1 U6369 ( .A1(n5533), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5512) );
  XNOR2_X1 U6370 ( .A(n5512), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6816) );
  AOI22_X1 U6371 ( .A1(n5711), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5710), .B2(
        n6816), .ZN(n5495) );
  NAND2_X1 U6372 ( .A1(n4860), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5503) );
  OR2_X1 U6373 ( .A1(n4851), .A2(n7764), .ZN(n5502) );
  NAND2_X1 U6374 ( .A1(n5497), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5519) );
  OR2_X1 U6375 ( .A1(n5497), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6376 ( .A1(n5519), .A2(n5498), .ZN(n8278) );
  OR2_X1 U6377 ( .A1(n5883), .A2(n8278), .ZN(n5501) );
  INV_X1 U6378 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5499) );
  OR2_X1 U6379 ( .A1(n5436), .A2(n5499), .ZN(n5500) );
  NAND2_X1 U6380 ( .A1(n8277), .A2(n8040), .ZN(n8708) );
  INV_X1 U6381 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6622) );
  INV_X1 U6382 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5507) );
  MUX2_X1 U6383 ( .A(n6622), .B(n5507), .S(n8295), .Z(n5508) );
  INV_X1 U6384 ( .A(SI_9_), .ZN(n9296) );
  INV_X1 U6385 ( .A(n5508), .ZN(n5509) );
  NAND2_X1 U6386 ( .A1(n5509), .A2(SI_9_), .ZN(n5510) );
  XNOR2_X1 U6387 ( .A(n5526), .B(n5313), .ZN(n6621) );
  NAND2_X1 U6388 ( .A1(n6621), .A2(n8541), .ZN(n5516) );
  INV_X1 U6389 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U6390 ( .A1(n5512), .A2(n5511), .ZN(n5513) );
  NAND2_X1 U6391 ( .A1(n5513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5514) );
  XNOR2_X1 U6392 ( .A(n5514), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6841) );
  AOI22_X1 U6393 ( .A1(n5711), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5710), .B2(
        n6841), .ZN(n5515) );
  NAND2_X1 U6394 ( .A1(n5516), .A2(n5515), .ZN(n10581) );
  NAND2_X1 U6395 ( .A1(n4860), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5524) );
  INV_X1 U6396 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5517) );
  OR2_X1 U6397 ( .A1(n4851), .A2(n5517), .ZN(n5523) );
  INV_X1 U6398 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U6399 ( .A1(n5519), .A2(n5518), .ZN(n5520) );
  NAND2_X1 U6400 ( .A1(n5539), .A2(n5520), .ZN(n8046) );
  OR2_X1 U6401 ( .A1(n5883), .A2(n8046), .ZN(n5522) );
  INV_X1 U6402 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6815) );
  OR2_X1 U6403 ( .A1(n5436), .A2(n6815), .ZN(n5521) );
  NAND4_X1 U6404 ( .A1(n5524), .A2(n5523), .A3(n5522), .A4(n5521), .ZN(n9895)
         );
  INV_X1 U6405 ( .A(n9895), .ZN(n7795) );
  NAND2_X1 U6406 ( .A1(n10581), .A2(n7795), .ZN(n8721) );
  INV_X1 U6407 ( .A(n8721), .ZN(n5525) );
  OR2_X1 U6408 ( .A1(n10581), .A2(n7795), .ZN(n8561) );
  OR2_X1 U6409 ( .A1(n8277), .A2(n8040), .ZN(n8557) );
  AND2_X1 U6410 ( .A1(n8561), .A2(n8557), .ZN(n8719) );
  INV_X1 U6411 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6632) );
  INV_X1 U6412 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6635) );
  MUX2_X1 U6413 ( .A(n6632), .B(n6635), .S(n8295), .Z(n5530) );
  INV_X1 U6414 ( .A(SI_10_), .ZN(n5529) );
  INV_X1 U6415 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U6416 ( .A1(n5531), .A2(SI_10_), .ZN(n5532) );
  XNOR2_X1 U6417 ( .A(n5545), .B(n5305), .ZN(n6631) );
  NAND2_X1 U6418 ( .A1(n6631), .A2(n8541), .ZN(n5537) );
  OR3_X1 U6419 ( .A1(n5533), .A2(P1_IR_REG_8__SCAN_IN), .A3(
        P1_IR_REG_9__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U6420 ( .A1(n5534), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5535) );
  XNOR2_X1 U6421 ( .A(n5535), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U6422 ( .A1(n5711), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5710), .B2(
        n10391), .ZN(n5536) );
  NAND2_X1 U6423 ( .A1(n4860), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5544) );
  INV_X1 U6424 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6811) );
  OR2_X1 U6425 ( .A1(n4851), .A2(n6811), .ZN(n5543) );
  INV_X1 U6426 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7493) );
  OR2_X1 U6427 ( .A1(n5436), .A2(n7493), .ZN(n5542) );
  INV_X1 U6428 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6429 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  NAND2_X1 U6430 ( .A1(n5559), .A2(n5540), .ZN(n8033) );
  OR2_X1 U6431 ( .A1(n5883), .A2(n8033), .ZN(n5541) );
  NAND4_X1 U6432 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .ZN(n9894)
         );
  INV_X1 U6433 ( .A(n9894), .ZN(n8041) );
  OR2_X1 U6434 ( .A1(n10596), .A2(n8041), .ZN(n8723) );
  NAND2_X1 U6435 ( .A1(n10596), .A2(n8041), .ZN(n8720) );
  NAND2_X1 U6436 ( .A1(n7490), .A2(n8664), .ZN(n7489) );
  NAND2_X1 U6437 ( .A1(n7489), .A2(n8720), .ZN(n7637) );
  INV_X1 U6438 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5549) );
  INV_X1 U6439 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5548) );
  MUX2_X1 U6440 ( .A(n5549), .B(n5548), .S(n8295), .Z(n5566) );
  XNOR2_X1 U6441 ( .A(n5570), .B(n5565), .ZN(n6633) );
  NAND2_X1 U6442 ( .A1(n6633), .A2(n8541), .ZN(n5556) );
  INV_X1 U6443 ( .A(n5550), .ZN(n5552) );
  NAND2_X1 U6444 ( .A1(n5552), .A2(n5551), .ZN(n5576) );
  NAND2_X1 U6445 ( .A1(n5576), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5554) );
  INV_X1 U6446 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5553) );
  XNOR2_X1 U6447 ( .A(n5554), .B(n5553), .ZN(n6823) );
  INV_X1 U6448 ( .A(n6823), .ZN(n6986) );
  AOI22_X1 U6449 ( .A1(n5711), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5710), .B2(
        n6986), .ZN(n5555) );
  NAND2_X1 U6450 ( .A1(n4860), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5564) );
  INV_X1 U6451 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5557) );
  OR2_X1 U6452 ( .A1(n4851), .A2(n5557), .ZN(n5563) );
  INV_X1 U6453 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5558) );
  AND2_X1 U6454 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  OR2_X1 U6455 ( .A1(n5560), .A2(n5581), .ZN(n8076) );
  OR2_X1 U6456 ( .A1(n5883), .A2(n8076), .ZN(n5562) );
  INV_X1 U6457 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6822) );
  OR2_X1 U6458 ( .A1(n5436), .A2(n6822), .ZN(n5561) );
  NAND4_X1 U6459 ( .A1(n5564), .A2(n5563), .A3(n5562), .A4(n5561), .ZN(n9893)
         );
  INV_X1 U6460 ( .A(n9893), .ZN(n8062) );
  OR2_X1 U6461 ( .A1(n8078), .A2(n8062), .ZN(n8728) );
  NAND2_X1 U6462 ( .A1(n8078), .A2(n8062), .ZN(n8725) );
  INV_X1 U6463 ( .A(n5566), .ZN(n5567) );
  INV_X1 U6464 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5571) );
  INV_X1 U6465 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6642) );
  MUX2_X1 U6466 ( .A(n5571), .B(n6642), .S(n8295), .Z(n5573) );
  INV_X1 U6467 ( .A(SI_12_), .ZN(n5572) );
  INV_X1 U6468 ( .A(n5573), .ZN(n5574) );
  NAND2_X1 U6469 ( .A1(n5574), .A2(SI_12_), .ZN(n5575) );
  XNOR2_X1 U6470 ( .A(n5589), .B(n5588), .ZN(n6638) );
  NAND2_X1 U6471 ( .A1(n6638), .A2(n8541), .ZN(n5580) );
  INV_X1 U6472 ( .A(n5576), .ZN(n5577) );
  NAND2_X1 U6473 ( .A1(n5578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5595) );
  XNOR2_X1 U6474 ( .A(n5595), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7120) );
  AOI22_X1 U6475 ( .A1(n5711), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5710), .B2(
        n7120), .ZN(n5579) );
  NAND2_X1 U6476 ( .A1(n4860), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5587) );
  INV_X1 U6477 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6989) );
  OR2_X1 U6478 ( .A1(n4851), .A2(n6989), .ZN(n5586) );
  NAND2_X1 U6479 ( .A1(n5581), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5601) );
  OR2_X1 U6480 ( .A1(n5581), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U6481 ( .A1(n5601), .A2(n5582), .ZN(n8220) );
  OR2_X1 U6482 ( .A1(n5883), .A2(n8220), .ZN(n5585) );
  INV_X1 U6483 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5583) );
  OR2_X1 U6484 ( .A1(n5436), .A2(n5583), .ZN(n5584) );
  NAND4_X1 U6485 ( .A1(n5587), .A2(n5586), .A3(n5585), .A4(n5584), .ZN(n9892)
         );
  INV_X1 U6486 ( .A(n9892), .ZN(n8201) );
  OR2_X1 U6487 ( .A1(n8203), .A2(n8201), .ZN(n8729) );
  NAND2_X1 U6488 ( .A1(n8203), .A2(n8201), .ZN(n8706) );
  INV_X1 U6489 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6655) );
  MUX2_X1 U6490 ( .A(n6655), .B(n6970), .S(n8295), .Z(n5591) );
  INV_X1 U6491 ( .A(SI_13_), .ZN(n9283) );
  NAND2_X1 U6492 ( .A1(n5591), .A2(n9283), .ZN(n5609) );
  INV_X1 U6493 ( .A(n5591), .ZN(n5592) );
  NAND2_X1 U6494 ( .A1(n5592), .A2(SI_13_), .ZN(n5593) );
  XNOR2_X1 U6495 ( .A(n5608), .B(n5312), .ZN(n6654) );
  NAND2_X1 U6496 ( .A1(n6654), .A2(n8541), .ZN(n5599) );
  NAND2_X1 U6497 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  NAND2_X1 U6498 ( .A1(n5596), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5597) );
  XNOR2_X1 U6499 ( .A(n5597), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7436) );
  AOI22_X1 U6500 ( .A1(n5711), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5710), .B2(
        n7436), .ZN(n5598) );
  NAND2_X1 U6501 ( .A1(n4860), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5607) );
  INV_X1 U6502 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7118) );
  OR2_X1 U6503 ( .A1(n4851), .A2(n7118), .ZN(n5606) );
  INV_X1 U6504 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U6505 ( .A1(n5601), .A2(n5600), .ZN(n5602) );
  NAND2_X1 U6506 ( .A1(n5618), .A2(n5602), .ZN(n8245) );
  OR2_X1 U6507 ( .A1(n5883), .A2(n8245), .ZN(n5605) );
  INV_X1 U6508 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5603) );
  OR2_X1 U6509 ( .A1(n5436), .A2(n5603), .ZN(n5604) );
  NAND4_X1 U6510 ( .A1(n5607), .A2(n5606), .A3(n5605), .A4(n5604), .ZN(n9891)
         );
  INV_X1 U6511 ( .A(n9891), .ZN(n9754) );
  OR2_X1 U6512 ( .A1(n10261), .A2(n9754), .ZN(n8730) );
  NAND2_X1 U6513 ( .A1(n10261), .A2(n9754), .ZN(n8707) );
  NAND2_X1 U6514 ( .A1(n7885), .A2(n8649), .ZN(n7963) );
  MUX2_X1 U6515 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n8295), .Z(n5627) );
  INV_X1 U6516 ( .A(SI_14_), .ZN(n9163) );
  XNOR2_X1 U6517 ( .A(n5630), .B(n5626), .ZN(n6729) );
  NAND2_X1 U6518 ( .A1(n6729), .A2(n8541), .ZN(n5617) );
  NOR2_X1 U6519 ( .A1(n5614), .A2(n5331), .ZN(n5612) );
  MUX2_X1 U6520 ( .A(n5331), .B(n5612), .S(P1_IR_REG_14__SCAN_IN), .Z(n5615)
         );
  INV_X1 U6521 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5613) );
  NOR2_X1 U6522 ( .A1(n5615), .A2(n5652), .ZN(n7731) );
  AOI22_X1 U6523 ( .A1(n5711), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5710), .B2(
        n7731), .ZN(n5616) );
  NAND2_X2 U6524 ( .A1(n5617), .A2(n5616), .ZN(n10257) );
  INV_X1 U6525 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7437) );
  AND2_X1 U6526 ( .A1(n5618), .A2(n7437), .ZN(n5619) );
  NOR2_X1 U6527 ( .A1(n5637), .A2(n5619), .ZN(n9750) );
  NAND2_X1 U6528 ( .A1(n5442), .A2(n9750), .ZN(n5624) );
  INV_X1 U6529 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7722) );
  OR2_X1 U6530 ( .A1(n4851), .A2(n7722), .ZN(n5623) );
  INV_X1 U6531 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7430) );
  OR2_X1 U6532 ( .A1(n5436), .A2(n7430), .ZN(n5622) );
  INV_X1 U6533 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5620) );
  OR2_X1 U6534 ( .A1(n5445), .A2(n5620), .ZN(n5621) );
  NAND4_X1 U6535 ( .A1(n5624), .A2(n5623), .A3(n5622), .A4(n5621), .ZN(n9890)
         );
  INV_X1 U6536 ( .A(n9890), .ZN(n8242) );
  OR2_X1 U6537 ( .A1(n10257), .A2(n8242), .ZN(n8731) );
  NAND2_X1 U6538 ( .A1(n10257), .A2(n8242), .ZN(n8735) );
  NAND2_X1 U6539 ( .A1(n8731), .A2(n8735), .ZN(n8667) );
  INV_X1 U6540 ( .A(n8707), .ZN(n8568) );
  NOR2_X1 U6541 ( .A1(n8667), .A2(n8568), .ZN(n5625) );
  NAND2_X1 U6542 ( .A1(n7963), .A2(n5625), .ZN(n7961) );
  NAND2_X1 U6543 ( .A1(n5627), .A2(SI_14_), .ZN(n5628) );
  INV_X1 U6544 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6883) );
  INV_X1 U6545 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6881) );
  MUX2_X1 U6546 ( .A(n6883), .B(n6881), .S(n8295), .Z(n5631) );
  INV_X1 U6547 ( .A(SI_15_), .ZN(n9285) );
  INV_X1 U6548 ( .A(n5631), .ZN(n5632) );
  NAND2_X1 U6549 ( .A1(n5632), .A2(SI_15_), .ZN(n5633) );
  NAND2_X1 U6550 ( .A1(n5645), .A2(n5633), .ZN(n5646) );
  XNOR2_X1 U6551 ( .A(n5647), .B(n5646), .ZN(n6880) );
  NAND2_X1 U6552 ( .A1(n6880), .A2(n8541), .ZN(n5636) );
  OR2_X1 U6553 ( .A1(n5652), .A2(n5331), .ZN(n5634) );
  INV_X1 U6554 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5651) );
  XNOR2_X1 U6555 ( .A(n5634), .B(n5651), .ZN(n7875) );
  INV_X1 U6556 ( .A(n7875), .ZN(n7729) );
  AOI22_X1 U6557 ( .A1(n5711), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5710), .B2(
        n7729), .ZN(n5635) );
  NOR2_X1 U6558 ( .A1(n5637), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5638) );
  OR2_X1 U6559 ( .A1(n5655), .A2(n5638), .ZN(n9875) );
  INV_X1 U6560 ( .A(n9875), .ZN(n8157) );
  NAND2_X1 U6561 ( .A1(n5442), .A2(n8157), .ZN(n5643) );
  INV_X1 U6562 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7726) );
  OR2_X1 U6563 ( .A1(n4851), .A2(n7726), .ZN(n5642) );
  INV_X1 U6564 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5639) );
  OR2_X1 U6565 ( .A1(n5445), .A2(n5639), .ZN(n5641) );
  INV_X1 U6566 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7733) );
  OR2_X1 U6567 ( .A1(n5436), .A2(n7733), .ZN(n5640) );
  NAND4_X1 U6568 ( .A1(n5643), .A2(n5642), .A3(n5641), .A4(n5640), .ZN(n9889)
         );
  INV_X1 U6569 ( .A(n9889), .ZN(n8853) );
  OR2_X1 U6570 ( .A1(n10249), .A2(n8853), .ZN(n8738) );
  NAND2_X1 U6571 ( .A1(n10249), .A2(n8853), .ZN(n8736) );
  NAND2_X1 U6572 ( .A1(n8738), .A2(n8736), .ZN(n8668) );
  INV_X1 U6573 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6967) );
  INV_X1 U6574 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6982) );
  MUX2_X1 U6575 ( .A(n6967), .B(n6982), .S(n8295), .Z(n5648) );
  INV_X1 U6576 ( .A(SI_16_), .ZN(n9282) );
  NAND2_X1 U6577 ( .A1(n5648), .A2(n9282), .ZN(n5666) );
  INV_X1 U6578 ( .A(n5648), .ZN(n5649) );
  NAND2_X1 U6579 ( .A1(n5649), .A2(SI_16_), .ZN(n5650) );
  XNOR2_X1 U6580 ( .A(n5665), .B(n5664), .ZN(n6966) );
  NAND2_X1 U6581 ( .A1(n6966), .A2(n8541), .ZN(n5654) );
  NAND2_X1 U6582 ( .A1(n5706), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5669) );
  XNOR2_X1 U6583 ( .A(n5669), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9908) );
  AOI22_X1 U6584 ( .A1(n5711), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5710), .B2(
        n9908), .ZN(n5653) );
  OR2_X1 U6585 ( .A1(n5655), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5656) );
  AND2_X1 U6586 ( .A1(n5674), .A2(n5656), .ZN(n9807) );
  NAND2_X1 U6587 ( .A1(n5442), .A2(n9807), .ZN(n5662) );
  NAND2_X1 U6588 ( .A1(n5848), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5661) );
  INV_X1 U6589 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5657) );
  OR2_X1 U6590 ( .A1(n5445), .A2(n5657), .ZN(n5660) );
  INV_X1 U6591 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5658) );
  OR2_X1 U6592 ( .A1(n5436), .A2(n5658), .ZN(n5659) );
  NAND4_X1 U6593 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .ZN(n9888)
         );
  INV_X1 U6594 ( .A(n9888), .ZN(n9870) );
  OR2_X1 U6595 ( .A1(n10246), .A2(n9870), .ZN(n8739) );
  NAND2_X1 U6596 ( .A1(n10246), .A2(n9870), .ZN(n8702) );
  NAND2_X1 U6597 ( .A1(n5663), .A2(n8702), .ZN(n8253) );
  NAND2_X2 U6598 ( .A1(n5667), .A2(n5666), .ZN(n5683) );
  MUX2_X1 U6599 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n8295), .Z(n5684) );
  INV_X1 U6600 ( .A(SI_17_), .ZN(n5668) );
  XNOR2_X1 U6601 ( .A(n5684), .B(n5668), .ZN(n5681) );
  XNOR2_X1 U6602 ( .A(n5683), .B(n5681), .ZN(n7001) );
  NAND2_X1 U6603 ( .A1(n7001), .A2(n8541), .ZN(n5672) );
  INV_X1 U6604 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U6605 ( .A1(n5669), .A2(n5704), .ZN(n5670) );
  NAND2_X1 U6606 ( .A1(n5670), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5686) );
  XNOR2_X1 U6607 ( .A(n5686), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U6608 ( .A1(n5711), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9919), .B2(
        n5710), .ZN(n5671) );
  INV_X1 U6609 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U6610 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  NAND2_X1 U6611 ( .A1(n5691), .A2(n5675), .ZN(n9819) );
  NAND2_X1 U6612 ( .A1(n4860), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5676) );
  OAI21_X1 U6613 ( .B1(n9819), .B2(n5883), .A(n5676), .ZN(n5680) );
  INV_X1 U6614 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U6615 ( .A1(n6624), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5677) );
  OAI21_X1 U6616 ( .B1(n5678), .B2(n5403), .A(n5677), .ZN(n5679) );
  OR2_X1 U6617 ( .A1(n5680), .A2(n5679), .ZN(n9887) );
  INV_X1 U6618 ( .A(n9887), .ZN(n10150) );
  OR2_X1 U6619 ( .A1(n10239), .A2(n10150), .ZN(n8687) );
  NAND2_X1 U6620 ( .A1(n10239), .A2(n10150), .ZN(n8703) );
  NAND2_X1 U6621 ( .A1(n8687), .A2(n8703), .ZN(n8672) );
  INV_X1 U6622 ( .A(n5681), .ZN(n5682) );
  NAND2_X1 U6623 ( .A1(n5684), .A2(SI_17_), .ZN(n5685) );
  MUX2_X1 U6624 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n8295), .Z(n5698) );
  XNOR2_X1 U6625 ( .A(n5698), .B(SI_18_), .ZN(n5695) );
  XNOR2_X1 U6626 ( .A(n5697), .B(n5695), .ZN(n7037) );
  NAND2_X1 U6627 ( .A1(n7037), .A2(n8541), .ZN(n5690) );
  INV_X1 U6628 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U6629 ( .A1(n5686), .A2(n5705), .ZN(n5687) );
  NAND2_X1 U6630 ( .A1(n5687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5688) );
  XNOR2_X1 U6631 ( .A(n5688), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U6632 ( .A1(n9935), .A2(n5710), .B1(n5711), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5689) );
  INV_X1 U6633 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9850) );
  AND2_X1 U6634 ( .A1(n5691), .A2(n9850), .ZN(n5692) );
  OR2_X1 U6635 ( .A1(n5692), .A2(n5714), .ZN(n10161) );
  AOI22_X1 U6636 ( .A1(n4860), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n5848), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U6637 ( .A1(n6624), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5693) );
  OAI211_X1 U6638 ( .C1(n10161), .C2(n5883), .A(n5694), .B(n5693), .ZN(n10121)
         );
  INV_X1 U6639 ( .A(n10121), .ZN(n9818) );
  OR2_X1 U6640 ( .A1(n10231), .A2(n9818), .ZN(n8688) );
  NAND2_X1 U6641 ( .A1(n10231), .A2(n9818), .ZN(n8705) );
  NAND2_X1 U6642 ( .A1(n8688), .A2(n8705), .ZN(n10143) );
  INV_X1 U6643 ( .A(n5695), .ZN(n5696) );
  INV_X1 U6644 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8315) );
  INV_X1 U6645 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n5699) );
  MUX2_X1 U6646 ( .A(n8315), .B(n5699), .S(n8295), .Z(n5700) );
  INV_X1 U6647 ( .A(SI_19_), .ZN(n9280) );
  NAND2_X1 U6648 ( .A1(n5700), .A2(n9280), .ZN(n5719) );
  INV_X1 U6649 ( .A(n5700), .ZN(n5701) );
  NAND2_X1 U6650 ( .A1(n5701), .A2(SI_19_), .ZN(n5702) );
  NAND2_X1 U6651 ( .A1(n5719), .A2(n5702), .ZN(n5720) );
  XNOR2_X1 U6652 ( .A(n5721), .B(n5720), .ZN(n7331) );
  NAND2_X1 U6653 ( .A1(n7331), .A2(n8541), .ZN(n5713) );
  INV_X1 U6654 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5703) );
  INV_X1 U6655 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6656 ( .A1(n4898), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5708) );
  INV_X2 U6657 ( .A(n9944), .ZN(n10095) );
  AOI22_X1 U6658 ( .A1(n5711), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10095), 
        .B2(n5710), .ZN(n5712) );
  NOR2_X1 U6659 ( .A1(n5714), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5715) );
  OR2_X1 U6660 ( .A1(n5728), .A2(n5715), .ZN(n10126) );
  AOI22_X1 U6661 ( .A1(n4860), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n5848), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n5718) );
  INV_X1 U6662 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5716) );
  OR2_X1 U6663 ( .A1(n5436), .A2(n5716), .ZN(n5717) );
  OAI211_X1 U6664 ( .C1(n10126), .C2(n5883), .A(n5718), .B(n5717), .ZN(n10147)
         );
  INV_X1 U6665 ( .A(n10147), .ZN(n10110) );
  OR2_X1 U6666 ( .A1(n10226), .A2(n10110), .ZN(n8691) );
  NAND2_X1 U6667 ( .A1(n10226), .A2(n10110), .ZN(n8699) );
  NAND2_X1 U6668 ( .A1(n8691), .A2(n8699), .ZN(n10132) );
  INV_X1 U6669 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7526) );
  INV_X1 U6670 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n5725) );
  MUX2_X1 U6671 ( .A(n7526), .B(n5725), .S(n8295), .Z(n5722) );
  INV_X1 U6672 ( .A(SI_20_), .ZN(n9277) );
  NAND2_X1 U6673 ( .A1(n5722), .A2(n9277), .ZN(n5737) );
  INV_X1 U6674 ( .A(n5722), .ZN(n5723) );
  NAND2_X1 U6675 ( .A1(n5723), .A2(SI_20_), .ZN(n5724) );
  XNOR2_X1 U6676 ( .A(n5736), .B(n5735), .ZN(n7485) );
  NAND2_X1 U6677 ( .A1(n7485), .A2(n8541), .ZN(n5727) );
  OR2_X1 U6678 ( .A1(n8544), .A2(n5725), .ZN(n5726) );
  NOR2_X1 U6679 ( .A1(n5728), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5729) );
  OR2_X1 U6680 ( .A1(n5741), .A2(n5729), .ZN(n10103) );
  INV_X1 U6681 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U6682 ( .A1(n6624), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U6683 ( .A1(n5848), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5730) );
  OAI211_X1 U6684 ( .C1(n5445), .C2(n5732), .A(n5731), .B(n5730), .ZN(n5733)
         );
  INV_X1 U6685 ( .A(n5733), .ZN(n5734) );
  OAI21_X1 U6686 ( .B1(n10103), .B2(n5883), .A(n5734), .ZN(n10122) );
  INV_X1 U6687 ( .A(n10122), .ZN(n9782) );
  NAND2_X1 U6688 ( .A1(n10222), .A2(n9782), .ZN(n8604) );
  NOR2_X1 U6689 ( .A1(n10108), .A2(n10109), .ZN(n10085) );
  MUX2_X1 U6690 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n8295), .Z(n5750) );
  INV_X1 U6691 ( .A(SI_21_), .ZN(n5738) );
  XNOR2_X1 U6692 ( .A(n5750), .B(n5738), .ZN(n5749) );
  XNOR2_X1 U6693 ( .A(n5751), .B(n5749), .ZN(n7487) );
  NAND2_X1 U6694 ( .A1(n7487), .A2(n8541), .ZN(n5740) );
  INV_X1 U6695 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7509) );
  OR2_X1 U6696 ( .A1(n8544), .A2(n7509), .ZN(n5739) );
  OR2_X1 U6697 ( .A1(n5741), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5742) );
  AND2_X1 U6698 ( .A1(n5742), .A2(n5759), .ZN(n10092) );
  NAND2_X1 U6699 ( .A1(n10092), .A2(n5442), .ZN(n5748) );
  INV_X1 U6700 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U6701 ( .A1(n5848), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U6702 ( .A1(n6624), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5743) );
  OAI211_X1 U6703 ( .C1(n5745), .C2(n5445), .A(n5744), .B(n5743), .ZN(n5746)
         );
  INV_X1 U6704 ( .A(n5746), .ZN(n5747) );
  NAND2_X1 U6705 ( .A1(n5748), .A2(n5747), .ZN(n9886) );
  INV_X1 U6706 ( .A(n9886), .ZN(n10112) );
  OR2_X1 U6707 ( .A1(n10217), .A2(n10112), .ZN(n8606) );
  NAND2_X1 U6708 ( .A1(n8606), .A2(n10086), .ZN(n8694) );
  NAND2_X1 U6709 ( .A1(n10217), .A2(n10112), .ZN(n8607) );
  OAI21_X1 U6710 ( .B1(n10085), .B2(n8694), .A(n8607), .ZN(n10075) );
  INV_X1 U6711 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8539) );
  INV_X1 U6712 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9039) );
  MUX2_X1 U6713 ( .A(n8539), .B(n9039), .S(n8295), .Z(n5753) );
  INV_X1 U6714 ( .A(SI_22_), .ZN(n5752) );
  NAND2_X1 U6715 ( .A1(n5753), .A2(n5752), .ZN(n5767) );
  INV_X1 U6716 ( .A(n5753), .ZN(n5754) );
  NAND2_X1 U6717 ( .A1(n5754), .A2(SI_22_), .ZN(n5755) );
  NAND2_X1 U6718 ( .A1(n5767), .A2(n5755), .ZN(n5768) );
  XNOR2_X1 U6719 ( .A(n5769), .B(n5768), .ZN(n8536) );
  NAND2_X1 U6720 ( .A1(n8536), .A2(n8541), .ZN(n5757) );
  OR2_X1 U6721 ( .A1(n8544), .A2(n9039), .ZN(n5756) );
  NAND2_X1 U6722 ( .A1(n5848), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5765) );
  INV_X1 U6723 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n5758) );
  OR2_X1 U6724 ( .A1(n5445), .A2(n5758), .ZN(n5764) );
  OAI21_X1 U6725 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n5760), .A(n5779), .ZN(
        n10071) );
  OR2_X1 U6726 ( .A1(n5883), .A2(n10071), .ZN(n5763) );
  INV_X1 U6727 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5761) );
  OR2_X1 U6728 ( .A1(n5436), .A2(n5761), .ZN(n5762) );
  NAND4_X1 U6729 ( .A1(n5765), .A2(n5764), .A3(n5763), .A4(n5762), .ZN(n10055)
         );
  INV_X1 U6730 ( .A(n10055), .ZN(n10091) );
  NAND2_X1 U6731 ( .A1(n10211), .A2(n10091), .ZN(n8685) );
  NAND2_X1 U6732 ( .A1(n8695), .A2(n8685), .ZN(n10076) );
  NOR2_X1 U6733 ( .A1(n10075), .A2(n10076), .ZN(n10074) );
  INV_X1 U6734 ( .A(n8695), .ZN(n5766) );
  INV_X1 U6735 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7779) );
  INV_X1 U6736 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7783) );
  MUX2_X1 U6737 ( .A(n7779), .B(n7783), .S(n8295), .Z(n5770) );
  INV_X1 U6738 ( .A(SI_23_), .ZN(n9254) );
  NAND2_X1 U6739 ( .A1(n5770), .A2(n9254), .ZN(n5786) );
  INV_X1 U6740 ( .A(n5770), .ZN(n5771) );
  NAND2_X1 U6741 ( .A1(n5771), .A2(SI_23_), .ZN(n5772) );
  AND2_X1 U6742 ( .A1(n5786), .A2(n5772), .ZN(n5773) );
  OR2_X1 U6743 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  NAND2_X1 U6744 ( .A1(n5787), .A2(n5775), .ZN(n7780) );
  NAND2_X1 U6745 ( .A1(n7780), .A2(n8541), .ZN(n5777) );
  OR2_X1 U6746 ( .A1(n8544), .A2(n7783), .ZN(n5776) );
  NAND2_X1 U6747 ( .A1(n5848), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5785) );
  INV_X1 U6748 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n5778) );
  OR2_X1 U6749 ( .A1(n5445), .A2(n5778), .ZN(n5784) );
  OAI21_X1 U6750 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n5780), .A(n5792), .ZN(
        n10059) );
  OR2_X1 U6751 ( .A1(n5883), .A2(n10059), .ZN(n5783) );
  INV_X1 U6752 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5781) );
  OR2_X1 U6753 ( .A1(n5436), .A2(n5781), .ZN(n5782) );
  NAND4_X1 U6754 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n10037)
         );
  INV_X1 U6755 ( .A(n10037), .ZN(n10077) );
  AND2_X1 U6756 ( .A1(n10205), .A2(n10077), .ZN(n8744) );
  MUX2_X1 U6757 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n8295), .Z(n5800) );
  INV_X1 U6758 ( .A(SI_24_), .ZN(n9271) );
  XNOR2_X1 U6759 ( .A(n5800), .B(n9271), .ZN(n5799) );
  XNOR2_X1 U6760 ( .A(n5803), .B(n5799), .ZN(n7841) );
  NAND2_X1 U6761 ( .A1(n7841), .A2(n8541), .ZN(n5790) );
  INV_X1 U6762 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5788) );
  OR2_X1 U6763 ( .A1(n8544), .A2(n5788), .ZN(n5789) );
  NAND2_X1 U6764 ( .A1(n5848), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5798) );
  INV_X1 U6765 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5791) );
  OR2_X1 U6766 ( .A1(n5445), .A2(n5791), .ZN(n5797) );
  OAI21_X1 U6767 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n5793), .A(n5812), .ZN(
        n10044) );
  OR2_X1 U6768 ( .A1(n5883), .A2(n10044), .ZN(n5796) );
  INV_X1 U6769 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5794) );
  OR2_X1 U6770 ( .A1(n5436), .A2(n5794), .ZN(n5795) );
  NAND4_X1 U6771 ( .A1(n5798), .A2(n5797), .A3(n5796), .A4(n5795), .ZN(n10054)
         );
  INV_X1 U6772 ( .A(n10054), .ZN(n10025) );
  OR2_X1 U6773 ( .A1(n10205), .A2(n10077), .ZN(n10032) );
  NAND2_X1 U6774 ( .A1(n8745), .A2(n10032), .ZN(n8698) );
  NAND2_X1 U6775 ( .A1(n10201), .A2(n10025), .ZN(n8747) );
  INV_X1 U6776 ( .A(n5799), .ZN(n5802) );
  NAND2_X1 U6777 ( .A1(n5800), .A2(SI_24_), .ZN(n5801) );
  INV_X1 U6778 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8056) );
  INV_X1 U6779 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5807) );
  MUX2_X1 U6780 ( .A(n8056), .B(n5807), .S(n8295), .Z(n5804) );
  INV_X1 U6781 ( .A(SI_25_), .ZN(n9184) );
  NAND2_X1 U6782 ( .A1(n5804), .A2(n9184), .ZN(n5838) );
  INV_X1 U6783 ( .A(n5804), .ZN(n5805) );
  NAND2_X1 U6784 ( .A1(n5805), .A2(SI_25_), .ZN(n5806) );
  NAND2_X1 U6785 ( .A1(n5838), .A2(n5806), .ZN(n5822) );
  NAND2_X1 U6786 ( .A1(n8054), .A2(n8541), .ZN(n5809) );
  OR2_X1 U6787 ( .A1(n8544), .A2(n5807), .ZN(n5808) );
  NAND2_X1 U6788 ( .A1(n4860), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5819) );
  INV_X1 U6789 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5810) );
  OR2_X1 U6790 ( .A1(n4851), .A2(n5810), .ZN(n5818) );
  INV_X1 U6791 ( .A(n5812), .ZN(n5814) );
  INV_X1 U6792 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5811) );
  INV_X1 U6793 ( .A(n5832), .ZN(n5813) );
  OAI21_X1 U6794 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n5814), .A(n5813), .ZN(
        n10018) );
  OR2_X1 U6795 ( .A1(n5883), .A2(n10018), .ZN(n5817) );
  INV_X1 U6796 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5815) );
  OR2_X1 U6797 ( .A1(n5436), .A2(n5815), .ZN(n5816) );
  NAND4_X1 U6798 ( .A1(n5819), .A2(n5818), .A3(n5817), .A4(n5816), .ZN(n10038)
         );
  NAND2_X1 U6799 ( .A1(n10196), .A2(n9997), .ZN(n8748) );
  INV_X1 U6800 ( .A(n8750), .ZN(n5820) );
  INV_X1 U6801 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8082) );
  INV_X1 U6802 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5828) );
  MUX2_X1 U6803 ( .A(n8082), .B(n5828), .S(n8295), .Z(n5824) );
  INV_X1 U6804 ( .A(SI_26_), .ZN(n9172) );
  NAND2_X1 U6805 ( .A1(n5824), .A2(n9172), .ZN(n5837) );
  INV_X1 U6806 ( .A(n5824), .ZN(n5825) );
  NAND2_X1 U6807 ( .A1(n5825), .A2(SI_26_), .ZN(n5839) );
  AND2_X1 U6808 ( .A1(n5837), .A2(n5839), .ZN(n5826) );
  OR2_X1 U6809 ( .A1(n8544), .A2(n5828), .ZN(n5829) );
  NAND2_X1 U6810 ( .A1(n5848), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5836) );
  INV_X1 U6811 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n5831) );
  OR2_X1 U6812 ( .A1(n5445), .A2(n5831), .ZN(n5835) );
  NAND2_X1 U6813 ( .A1(n5832), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5850) );
  OAI21_X1 U6814 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n5832), .A(n5850), .ZN(
        n10004) );
  OR2_X1 U6815 ( .A1(n5883), .A2(n10004), .ZN(n5834) );
  INV_X1 U6816 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10005) );
  OR2_X1 U6817 ( .A1(n5436), .A2(n10005), .ZN(n5833) );
  NAND4_X1 U6818 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n5833), .ZN(n9885)
         );
  AND2_X1 U6819 ( .A1(n5838), .A2(n5837), .ZN(n5841) );
  INV_X1 U6820 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8112) );
  INV_X1 U6821 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8110) );
  MUX2_X1 U6822 ( .A(n8112), .B(n8110), .S(n8295), .Z(n5843) );
  INV_X1 U6823 ( .A(SI_27_), .ZN(n9173) );
  NAND2_X1 U6824 ( .A1(n5843), .A2(n9173), .ZN(n5859) );
  INV_X1 U6825 ( .A(n5843), .ZN(n5844) );
  NAND2_X1 U6826 ( .A1(n5844), .A2(SI_27_), .ZN(n5845) );
  AND2_X1 U6827 ( .A1(n5859), .A2(n5845), .ZN(n5857) );
  NAND2_X1 U6828 ( .A1(n8111), .A2(n8541), .ZN(n5847) );
  OR2_X1 U6829 ( .A1(n8544), .A2(n8110), .ZN(n5846) );
  NAND2_X1 U6830 ( .A1(n5848), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5856) );
  INV_X1 U6831 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5849) );
  OR2_X1 U6832 ( .A1(n5445), .A2(n5849), .ZN(n5855) );
  INV_X1 U6833 ( .A(n5850), .ZN(n5851) );
  NAND2_X1 U6834 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n5851), .ZN(n5866) );
  OAI21_X1 U6835 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n5851), .A(n5866), .ZN(
        n9981) );
  OR2_X1 U6836 ( .A1(n5883), .A2(n9981), .ZN(n5854) );
  INV_X1 U6837 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5852) );
  OR2_X1 U6838 ( .A1(n5436), .A2(n5852), .ZN(n5853) );
  NAND4_X1 U6839 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n9884)
         );
  NAND2_X1 U6840 ( .A1(n5955), .A2(n9998), .ZN(n8756) );
  MUX2_X1 U6841 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n8295), .Z(n5876) );
  INV_X1 U6842 ( .A(SI_28_), .ZN(n9263) );
  XNOR2_X1 U6843 ( .A(n5876), .B(n9263), .ZN(n5874) );
  INV_X1 U6844 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8180) );
  OR2_X1 U6845 ( .A1(n8544), .A2(n8180), .ZN(n5861) );
  NAND2_X1 U6846 ( .A1(n4860), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5872) );
  INV_X1 U6847 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5863) );
  OR2_X1 U6848 ( .A1(n5403), .A2(n5863), .ZN(n5871) );
  INV_X1 U6849 ( .A(n5866), .ZN(n5864) );
  NAND2_X1 U6850 ( .A1(n5864), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6577) );
  INV_X1 U6851 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U6852 ( .A1(n5866), .A2(n5865), .ZN(n5867) );
  NAND2_X1 U6853 ( .A1(n6577), .A2(n5867), .ZN(n9970) );
  OR2_X1 U6854 ( .A1(n5883), .A2(n9970), .ZN(n5870) );
  INV_X1 U6855 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5868) );
  OR2_X1 U6856 ( .A1(n5436), .A2(n5868), .ZN(n5869) );
  NAND4_X1 U6857 ( .A1(n5872), .A2(n5871), .A3(n5870), .A4(n5869), .ZN(n9883)
         );
  NAND2_X1 U6858 ( .A1(n10179), .A2(n9987), .ZN(n8757) );
  NOR2_X1 U6859 ( .A1(n9960), .A2(n9959), .ZN(n9958) );
  INV_X1 U6860 ( .A(n8628), .ZN(n5873) );
  NOR2_X1 U6861 ( .A1(n9958), .A2(n5873), .ZN(n5888) );
  INV_X1 U6862 ( .A(n5876), .ZN(n5877) );
  NAND2_X1 U6863 ( .A1(n5877), .A2(n9263), .ZN(n5878) );
  MUX2_X1 U6864 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n8295), .Z(n8288) );
  INV_X1 U6865 ( .A(SI_29_), .ZN(n9260) );
  XNOR2_X1 U6866 ( .A(n8288), .B(n9260), .ZN(n8286) );
  NAND2_X1 U6867 ( .A1(n8305), .A2(n8541), .ZN(n5881) );
  INV_X1 U6868 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9061) );
  OR2_X1 U6869 ( .A1(n8544), .A2(n9061), .ZN(n5880) );
  NAND2_X1 U6870 ( .A1(n6624), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5887) );
  INV_X1 U6871 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5882) );
  OR2_X1 U6872 ( .A1(n5445), .A2(n5882), .ZN(n5886) );
  OR2_X1 U6873 ( .A1(n4851), .A2(n5996), .ZN(n5885) );
  OR2_X1 U6874 ( .A1(n5883), .A2(n6577), .ZN(n5884) );
  NAND4_X1 U6875 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n9882)
         );
  INV_X1 U6876 ( .A(n9882), .ZN(n9961) );
  NAND2_X1 U6877 ( .A1(n5963), .A2(n9961), .ZN(n8810) );
  XNOR2_X1 U6878 ( .A(n5888), .B(n5957), .ZN(n5906) );
  INV_X1 U6879 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U6880 ( .A1(n5892), .A2(n5891), .ZN(n5893) );
  NAND2_X1 U6881 ( .A1(n5893), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5890) );
  INV_X1 U6882 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5889) );
  OR2_X1 U6883 ( .A1(n9041), .A2(n9944), .ZN(n5898) );
  OR2_X1 U6884 ( .A1(n5892), .A2(n5891), .ZN(n5894) );
  NAND2_X1 U6885 ( .A1(n5895), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5896) );
  INV_X1 U6886 ( .A(n7486), .ZN(n8816) );
  NAND2_X1 U6887 ( .A1(n5958), .A2(n8816), .ZN(n5897) );
  NAND2_X1 U6888 ( .A1(n8825), .A2(n5958), .ZN(n8645) );
  OR2_X1 U6889 ( .A1(n8645), .A2(n5899), .ZN(n10149) );
  INV_X1 U6890 ( .A(n5899), .ZN(n6920) );
  INV_X1 U6891 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U6892 ( .A1(n6624), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5902) );
  INV_X1 U6893 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5900) );
  OR2_X1 U6894 ( .A1(n5403), .A2(n5900), .ZN(n5901) );
  OAI211_X1 U6895 ( .C1(n5445), .C2(n5903), .A(n5902), .B(n5901), .ZN(n9881)
         );
  INV_X1 U6896 ( .A(n6785), .ZN(n8821) );
  NAND2_X1 U6897 ( .A1(n8821), .A2(P1_B_REG_SCAN_IN), .ZN(n9946) );
  NAND2_X1 U6898 ( .A1(n9881), .A2(n9946), .ZN(n5904) );
  OAI22_X1 U6899 ( .A1(n9987), .A2(n10149), .B1(n10111), .B2(n5904), .ZN(n5905) );
  AOI21_X1 U6900 ( .B1(n5906), .B2(n10152), .A(n5905), .ZN(n6574) );
  NAND2_X1 U6901 ( .A1(n7248), .A2(n5907), .ZN(n5909) );
  NAND2_X1 U6902 ( .A1(n6902), .A2(n8776), .ZN(n5908) );
  OR2_X1 U6903 ( .A1(n6914), .A2(n6911), .ZN(n5911) );
  NAND2_X1 U6904 ( .A1(n6971), .A2(n5911), .ZN(n7262) );
  NAND2_X1 U6905 ( .A1(n7262), .A2(n8651), .ZN(n7261) );
  OR2_X1 U6906 ( .A1(n6892), .A2(n7275), .ZN(n5913) );
  NAND2_X1 U6907 ( .A1(n7261), .A2(n5913), .ZN(n7085) );
  AND2_X1 U6908 ( .A1(n8787), .A2(n5914), .ZN(n8656) );
  INV_X1 U6909 ( .A(n8656), .ZN(n7088) );
  NAND2_X1 U6910 ( .A1(n7085), .A2(n7088), .ZN(n7084) );
  OR2_X1 U6911 ( .A1(n9900), .A2(n7175), .ZN(n5915) );
  NAND2_X1 U6912 ( .A1(n10514), .A2(n9899), .ZN(n5917) );
  OR2_X1 U6913 ( .A1(n7424), .A2(n9898), .ZN(n7396) );
  INV_X1 U6914 ( .A(n8040), .ZN(n9896) );
  NAND2_X1 U6915 ( .A1(n8277), .A2(n9896), .ZN(n5922) );
  INV_X1 U6916 ( .A(n5922), .ZN(n5919) );
  NAND2_X1 U6917 ( .A1(n8557), .A2(n8708), .ZN(n8659) );
  OR2_X1 U6918 ( .A1(n7523), .A2(n9897), .ZN(n7748) );
  AND2_X1 U6919 ( .A1(n8659), .A2(n7748), .ZN(n7749) );
  AND2_X1 U6920 ( .A1(n7396), .A2(n5921), .ZN(n5920) );
  NAND2_X1 U6921 ( .A1(n7412), .A2(n5920), .ZN(n5926) );
  INV_X1 U6922 ( .A(n5921), .ZN(n5924) );
  AND2_X1 U6923 ( .A1(n8658), .A2(n5922), .ZN(n5923) );
  OR2_X1 U6924 ( .A1(n5924), .A2(n5923), .ZN(n5925) );
  AND2_X1 U6925 ( .A1(n10581), .A2(n9895), .ZN(n5928) );
  OR2_X1 U6926 ( .A1(n10581), .A2(n9895), .ZN(n5927) );
  INV_X1 U6927 ( .A(n8664), .ZN(n5929) );
  NAND2_X1 U6928 ( .A1(n7639), .A2(n4980), .ZN(n5931) );
  OR2_X1 U6929 ( .A1(n8078), .A2(n9893), .ZN(n5930) );
  NAND2_X1 U6930 ( .A1(n8203), .A2(n9892), .ZN(n5933) );
  INV_X1 U6931 ( .A(n7889), .ZN(n5935) );
  OR2_X1 U6932 ( .A1(n10261), .A2(n9891), .ZN(n5936) );
  NAND2_X1 U6933 ( .A1(n10257), .A2(n9890), .ZN(n8152) );
  NAND2_X1 U6934 ( .A1(n10249), .A2(n9889), .ZN(n5938) );
  AND2_X1 U6935 ( .A1(n8152), .A2(n5938), .ZN(n5937) );
  NAND2_X1 U6936 ( .A1(n8153), .A2(n5937), .ZN(n8098) );
  INV_X1 U6937 ( .A(n5938), .ZN(n5939) );
  OR2_X1 U6938 ( .A1(n5939), .A2(n8668), .ZN(n8097) );
  AND2_X1 U6939 ( .A1(n8104), .A2(n8097), .ZN(n5940) );
  NAND2_X1 U6940 ( .A1(n8098), .A2(n5940), .ZN(n5942) );
  NAND2_X1 U6941 ( .A1(n10246), .A2(n9888), .ZN(n5941) );
  AND2_X1 U6942 ( .A1(n10239), .A2(n9887), .ZN(n5943) );
  INV_X1 U6943 ( .A(n10143), .ZN(n10139) );
  OR2_X1 U6944 ( .A1(n10226), .A2(n10147), .ZN(n5944) );
  NAND2_X1 U6945 ( .A1(n10133), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U6946 ( .A1(n10226), .A2(n10147), .ZN(n5945) );
  NAND2_X1 U6947 ( .A1(n5946), .A2(n5945), .ZN(n10099) );
  NAND2_X1 U6948 ( .A1(n10099), .A2(n10109), .ZN(n5948) );
  NAND2_X1 U6949 ( .A1(n10222), .A2(n10122), .ZN(n5947) );
  NAND2_X1 U6950 ( .A1(n5948), .A2(n5947), .ZN(n10083) );
  NAND2_X1 U6951 ( .A1(n8606), .A2(n8607), .ZN(n10088) );
  NAND2_X1 U6952 ( .A1(n10083), .A2(n10088), .ZN(n5950) );
  NAND2_X1 U6953 ( .A1(n10217), .A2(n9886), .ZN(n5949) );
  OR2_X1 U6954 ( .A1(n10211), .A2(n10055), .ZN(n5951) );
  OR2_X1 U6955 ( .A1(n10205), .A2(n10037), .ZN(n8612) );
  NAND2_X1 U6956 ( .A1(n4872), .A2(n5952), .ZN(n10040) );
  NAND2_X1 U6957 ( .A1(n10201), .A2(n10054), .ZN(n5953) );
  NAND2_X1 U6958 ( .A1(n10040), .A2(n5953), .ZN(n10014) );
  OR2_X1 U6959 ( .A1(n10196), .A2(n10038), .ZN(n5954) );
  INV_X1 U6960 ( .A(n10007), .ZN(n10189) );
  AOI21_X1 U6961 ( .B1(n9041), .B2(n6895), .A(n10095), .ZN(n5959) );
  NAND2_X1 U6962 ( .A1(n8825), .A2(n6708), .ZN(n6701) );
  NAND2_X2 U6963 ( .A1(n9041), .A2(n10095), .ZN(n8631) );
  INV_X1 U6964 ( .A(n10580), .ZN(n5960) );
  INV_X1 U6965 ( .A(n5955), .ZN(n9984) );
  INV_X1 U6966 ( .A(n10201), .ZN(n10048) );
  INV_X1 U6967 ( .A(n10222), .ZN(n10106) );
  INV_X1 U6968 ( .A(n10239), .ZN(n9825) );
  INV_X1 U6969 ( .A(n10246), .ZN(n9803) );
  OR2_X1 U6970 ( .A1(n7271), .A2(n7175), .ZN(n7105) );
  INV_X1 U6971 ( .A(n7424), .ZN(n7443) );
  INV_X1 U6972 ( .A(n7523), .ZN(n7406) );
  INV_X1 U6973 ( .A(n8078), .ZN(n10632) );
  INV_X1 U6974 ( .A(n8203), .ZN(n10652) );
  INV_X1 U6975 ( .A(n10261), .ZN(n7895) );
  NAND2_X1 U6976 ( .A1(n7890), .A2(n7895), .ZN(n7967) );
  NAND2_X1 U6977 ( .A1(n10048), .A2(n10058), .ZN(n10042) );
  INV_X1 U6978 ( .A(n9969), .ZN(n5962) );
  INV_X1 U6979 ( .A(n5963), .ZN(n6580) );
  AOI21_X1 U6980 ( .B1(n5963), .B2(n5962), .A(n9953), .ZN(n6582) );
  INV_X1 U6981 ( .A(n5958), .ZN(n8762) );
  NAND2_X1 U6982 ( .A1(n9041), .A2(n8762), .ZN(n6852) );
  INV_X1 U6983 ( .A(n10633), .ZN(n10250) );
  AND2_X1 U6984 ( .A1(n7486), .A2(n9944), .ZN(n8819) );
  OR2_X1 U6985 ( .A1(n6852), .A2(n8819), .ZN(n10651) );
  AOI22_X1 U6986 ( .A1(n6582), .A2(n10250), .B1(n10597), .B2(n5963), .ZN(n5964) );
  NAND3_X1 U6987 ( .A1(n6574), .A2(n5965), .A3(n5964), .ZN(n6568) );
  OR2_X1 U6988 ( .A1(n8645), .A2(n8819), .ZN(n6886) );
  NAND2_X1 U6989 ( .A1(n5966), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5972) );
  INV_X1 U6990 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U6991 ( .A1(n5972), .A2(n5971), .ZN(n5974) );
  NAND2_X1 U6992 ( .A1(n5974), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  INV_X1 U6993 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U6994 ( .A1(n4901), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5970) );
  XNOR2_X1 U6995 ( .A(n5970), .B(n5969), .ZN(n7866) );
  OR2_X1 U6996 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  NAND2_X1 U6997 ( .A1(n5974), .A2(n5973), .ZN(n8058) );
  NAND3_X1 U6998 ( .A1(n8058), .A2(P1_B_REG_SCAN_IN), .A3(n7866), .ZN(n5975)
         );
  OAI21_X1 U6999 ( .B1(P1_B_REG_SCAN_IN), .B2(n7866), .A(n5975), .ZN(n5976) );
  OR2_X1 U7000 ( .A1(n8096), .A2(n5976), .ZN(n10294) );
  NOR4_X1 U7001 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5985) );
  NOR4_X1 U7002 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5984) );
  OR4_X1 U7003 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n5982) );
  NOR4_X1 U7004 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5980) );
  NOR4_X1 U7005 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5979) );
  NOR4_X1 U7006 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5978) );
  NOR4_X1 U7007 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5977) );
  NAND4_X1 U7008 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(n5981)
         );
  NOR4_X1 U7009 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n5982), .A4(n5981), .ZN(n5983) );
  AND3_X1 U7010 ( .A1(n5985), .A2(n5984), .A3(n5983), .ZN(n5986) );
  NOR2_X1 U7011 ( .A1(n10294), .A2(n5986), .ZN(n6571) );
  INV_X1 U7012 ( .A(n6571), .ZN(n5990) );
  NAND2_X1 U7013 ( .A1(n5173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U7014 ( .A(n5988), .B(n5987), .ZN(n7781) );
  AND2_X1 U7015 ( .A1(n7781), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6586) );
  NAND2_X1 U7016 ( .A1(n8096), .A2(n8058), .ZN(n5989) );
  OAI21_X1 U7017 ( .B1(n10294), .B2(P1_D_REG_1__SCAN_IN), .A(n5989), .ZN(n6599) );
  AND3_X1 U7018 ( .A1(n5990), .A2(n10295), .A3(n6599), .ZN(n5991) );
  AND2_X1 U7019 ( .A1(n6886), .A2(n5991), .ZN(n5993) );
  OR2_X1 U7020 ( .A1(n10600), .A2(n5958), .ZN(n5992) );
  INV_X1 U7021 ( .A(n8096), .ZN(n5995) );
  INV_X1 U7022 ( .A(n7866), .ZN(n5994) );
  OAI22_X1 U7023 ( .A1(n10294), .A2(P1_D_REG_0__SCAN_IN), .B1(n5995), .B2(
        n5994), .ZN(n6698) );
  INV_X1 U7024 ( .A(n6698), .ZN(n10284) );
  NAND2_X1 U7025 ( .A1(n6567), .A2(n10284), .ZN(n10655) );
  INV_X2 U7026 ( .A(n10655), .ZN(n10656) );
  NAND2_X1 U7027 ( .A1(n6568), .A2(n10656), .ZN(n5997) );
  NAND2_X1 U7028 ( .A1(n5997), .A2(n5310), .ZN(P1_U3552) );
  NOR2_X1 U7029 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6003) );
  INV_X1 U7030 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6000) );
  NAND4_X1 U7031 ( .A1(n6003), .A2(n6002), .A3(n6001), .A4(n6000), .ZN(n6005)
         );
  INV_X1 U7032 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7033 ( .A1(n6014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7034 ( .A1(n6336), .A2(n6012), .ZN(n6006) );
  NAND2_X1 U7035 ( .A1(n6006), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7036 ( .A1(n6007), .A2(n6011), .ZN(n6008) );
  OR2_X1 U7037 ( .A1(n6007), .A2(n6011), .ZN(n6009) );
  NAND2_X1 U7038 ( .A1(n6015), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6016) );
  XNOR2_X1 U7039 ( .A(n6016), .B(n6021), .ZN(n8522) );
  NAND2_X1 U7040 ( .A1(n8532), .A2(n9601), .ZN(n6018) );
  NAND2_X1 U7041 ( .A1(n6019), .A2(n6018), .ZN(n6868) );
  INV_X1 U7042 ( .A(n7527), .ZN(n8524) );
  NAND2_X1 U7043 ( .A1(n8524), .A2(n5187), .ZN(n8340) );
  NOR2_X1 U7044 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n6022) );
  INV_X1 U7045 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6535) );
  INV_X1 U7046 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6505) );
  INV_X1 U7047 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6027) );
  XNOR2_X2 U7048 ( .A(n6028), .B(n6027), .ZN(n7063) );
  INV_X1 U7049 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7050 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6029) );
  XNOR2_X1 U7051 ( .A(n6030), .B(n6029), .ZN(n7071) );
  INV_X1 U7052 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6591) );
  INV_X1 U7053 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6033) );
  INV_X1 U7054 ( .A(n6035), .ZN(n6037) );
  NAND2_X2 U7055 ( .A1(n8997), .A2(n6037), .ZN(n6109) );
  INV_X1 U7056 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7070) );
  OR2_X1 U7057 ( .A1(n6109), .A2(n7070), .ZN(n6042) );
  NAND2_X1 U7058 ( .A1(n6856), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6041) );
  INV_X1 U7059 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6036) );
  OR2_X1 U7060 ( .A1(n6093), .A2(n6036), .ZN(n6040) );
  INV_X1 U7061 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9332) );
  OR2_X1 U7062 ( .A1(n6448), .A2(n9332), .ZN(n6039) );
  NAND4_X1 U7063 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n6943)
         );
  NAND2_X1 U7064 ( .A1(n9379), .A2(n8527), .ZN(n6055) );
  NAND2_X1 U7065 ( .A1(n6856), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6048) );
  INV_X1 U7066 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7533) );
  OR2_X1 U7067 ( .A1(n6448), .A2(n7533), .ZN(n6047) );
  INV_X1 U7068 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6043) );
  OR2_X1 U7069 ( .A1(n6093), .A2(n6043), .ZN(n6046) );
  INV_X1 U7070 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6044) );
  OR2_X1 U7071 ( .A1(n6109), .A2(n6044), .ZN(n6045) );
  NAND4_X1 U7072 ( .A1(n6048), .A2(n6047), .A3(n6046), .A4(n6045), .ZN(n6870)
         );
  INV_X1 U7073 ( .A(SI_0_), .ZN(n6050) );
  INV_X1 U7074 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6049) );
  OAI21_X1 U7075 ( .B1(n8295), .B2(n6050), .A(n6049), .ZN(n6052) );
  AND2_X1 U7076 ( .A1(n6052), .A2(n6051), .ZN(n9745) );
  MUX2_X1 U7077 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9745), .S(n7074), .Z(n10468)
         );
  AND2_X1 U7078 ( .A1(n6870), .A2(n10468), .ZN(n6945) );
  NAND2_X1 U7079 ( .A1(n6945), .A2(n8527), .ZN(n7033) );
  INV_X1 U7080 ( .A(n10468), .ZN(n7529) );
  NAND2_X1 U7081 ( .A1(n5193), .A2(n7529), .ZN(n6053) );
  AND2_X1 U7082 ( .A1(n7033), .A2(n6053), .ZN(n7015) );
  INV_X1 U7083 ( .A(n6054), .ZN(n6056) );
  NAND2_X1 U7084 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  NAND2_X1 U7085 ( .A1(n7014), .A2(n6057), .ZN(n7007) );
  INV_X1 U7086 ( .A(n7007), .ZN(n6072) );
  INV_X1 U7087 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7069) );
  OR2_X1 U7088 ( .A1(n6109), .A2(n7069), .ZN(n6062) );
  NAND2_X1 U7089 ( .A1(n6856), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6061) );
  INV_X1 U7090 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6058) );
  INV_X1 U7091 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7631) );
  AND4_X2 U7092 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n6948)
         );
  OR2_X1 U7093 ( .A1(n6063), .A2(n6515), .ZN(n6066) );
  INV_X1 U7094 ( .A(n6066), .ZN(n6064) );
  NAND2_X1 U7095 ( .A1(n6064), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n6067) );
  INV_X1 U7096 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7097 ( .A1(n6066), .A2(n6065), .ZN(n6080) );
  INV_X1 U7098 ( .A(n10454), .ZN(n6593) );
  INV_X1 U7099 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6594) );
  XNOR2_X1 U7100 ( .A(n5193), .B(n10478), .ZN(n10493) );
  NAND2_X1 U7101 ( .A1(n6068), .A2(n10493), .ZN(n6073) );
  INV_X1 U7102 ( .A(n10493), .ZN(n6070) );
  INV_X1 U7103 ( .A(n6068), .ZN(n6069) );
  NAND2_X1 U7104 ( .A1(n6073), .A2(n6071), .ZN(n7006) );
  NAND2_X1 U7105 ( .A1(n6856), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6078) );
  OR2_X1 U7106 ( .A1(n6448), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6077) );
  INV_X1 U7107 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6074) );
  OR2_X1 U7108 ( .A1(n6093), .A2(n6074), .ZN(n6076) );
  INV_X1 U7109 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7073) );
  OR2_X1 U7110 ( .A1(n6109), .A2(n7073), .ZN(n6075) );
  NOR2_X1 U7111 ( .A1(n7691), .A2(n6483), .ZN(n6085) );
  NAND2_X1 U7112 ( .A1(n6080), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6081) );
  XNOR2_X1 U7113 ( .A(n6081), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7143) );
  INV_X1 U7114 ( .A(n7143), .ZN(n7081) );
  OR2_X1 U7115 ( .A1(n6609), .A2(n6104), .ZN(n6083) );
  INV_X1 U7116 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6592) );
  OR2_X1 U7117 ( .A1(n6366), .A2(n6592), .ZN(n6082) );
  OAI211_X1 U7118 ( .C1(n7074), .C2(n7081), .A(n6083), .B(n6082), .ZN(n6960)
         );
  INV_X1 U7119 ( .A(n6960), .ZN(n10502) );
  XNOR2_X1 U7120 ( .A(n5193), .B(n10502), .ZN(n6084) );
  NAND2_X1 U7121 ( .A1(n6085), .A2(n6084), .ZN(n6099) );
  OR2_X1 U7122 ( .A1(n6607), .A2(n6104), .ZN(n6091) );
  NOR2_X1 U7123 ( .A1(n6086), .A2(n6515), .ZN(n6087) );
  MUX2_X1 U7124 ( .A(n6515), .B(n6087), .S(P2_IR_REG_4__SCAN_IN), .Z(n6089) );
  NOR2_X1 U7125 ( .A1(n6089), .A2(n6088), .ZN(n7146) );
  AOI22_X1 U7126 ( .A1(n6350), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7022), .B2(
        n7146), .ZN(n6090) );
  NAND2_X1 U7127 ( .A1(n6856), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6098) );
  INV_X1 U7128 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6092) );
  INV_X1 U7129 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6094) );
  OR2_X1 U7130 ( .A1(n6093), .A2(n6094), .ZN(n6096) );
  XNOR2_X1 U7131 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7699) );
  OR2_X1 U7132 ( .A1(n6448), .A2(n7699), .ZN(n6095) );
  NAND2_X1 U7133 ( .A1(n9377), .A2(n8527), .ZN(n6101) );
  XNOR2_X1 U7134 ( .A(n7476), .B(n6101), .ZN(n7054) );
  AND2_X1 U7135 ( .A1(n7054), .A2(n6099), .ZN(n6100) );
  INV_X1 U7136 ( .A(n7476), .ZN(n6102) );
  NAND2_X1 U7137 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  NAND2_X1 U7138 ( .A1(n7050), .A2(n6103), .ZN(n6119) );
  INV_X2 U7139 ( .A(n6104), .ZN(n8304) );
  NAND2_X1 U7140 ( .A1(n6600), .A2(n8304), .ZN(n6107) );
  OR2_X1 U7141 ( .A1(n6088), .A2(n6515), .ZN(n6105) );
  XNOR2_X1 U7142 ( .A(n6105), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7147) );
  AOI22_X1 U7143 ( .A1(n6350), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7022), .B2(
        n7147), .ZN(n6106) );
  XNOR2_X1 U7144 ( .A(n7566), .B(n6079), .ZN(n8961) );
  NAND2_X1 U7145 ( .A1(n6856), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6118) );
  INV_X1 U7146 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6108) );
  OR2_X1 U7147 ( .A1(n6109), .A2(n6108), .ZN(n6117) );
  INV_X1 U7148 ( .A(n6128), .ZN(n6113) );
  INV_X1 U7149 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7150 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6110) );
  NAND2_X1 U7151 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  NAND2_X1 U7152 ( .A1(n6113), .A2(n6112), .ZN(n7612) );
  OR2_X1 U7153 ( .A1(n6448), .A2(n7612), .ZN(n6116) );
  INV_X1 U7154 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6114) );
  OR2_X1 U7155 ( .A1(n6093), .A2(n6114), .ZN(n6115) );
  NOR2_X1 U7156 ( .A1(n9375), .A2(n6483), .ZN(n6120) );
  XNOR2_X1 U7157 ( .A(n8961), .B(n6120), .ZN(n7478) );
  INV_X1 U7158 ( .A(n6120), .ZN(n6121) );
  NAND2_X1 U7159 ( .A1(n8961), .A2(n6121), .ZN(n6122) );
  NAND2_X1 U7160 ( .A1(n8964), .A2(n6122), .ZN(n6134) );
  NAND2_X1 U7161 ( .A1(n6610), .A2(n8304), .ZN(n6126) );
  INV_X1 U7162 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7163 ( .A1(n6088), .A2(n6123), .ZN(n6139) );
  NAND2_X1 U7164 ( .A1(n6139), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6124) );
  XNOR2_X1 U7165 ( .A(n6124), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7150) );
  AOI22_X1 U7166 ( .A1(n6350), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7022), .B2(
        n7150), .ZN(n6125) );
  XNOR2_X1 U7167 ( .A(n10527), .B(n6478), .ZN(n6135) );
  INV_X1 U7168 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6127) );
  INV_X1 U7169 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7659) );
  OR2_X1 U7170 ( .A1(n6160), .A2(n7659), .ZN(n6132) );
  NAND2_X1 U7171 ( .A1(n6128), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6145) );
  OAI21_X1 U7172 ( .B1(n6128), .B2(P2_REG3_REG_6__SCAN_IN), .A(n6145), .ZN(
        n8955) );
  OR2_X1 U7173 ( .A1(n6448), .A2(n8955), .ZN(n6131) );
  INV_X1 U7174 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6129) );
  OR2_X1 U7175 ( .A1(n6093), .A2(n6129), .ZN(n6130) );
  NAND2_X1 U7176 ( .A1(n10536), .A2(n8527), .ZN(n6136) );
  XNOR2_X1 U7177 ( .A(n6135), .B(n6136), .ZN(n8960) );
  INV_X1 U7178 ( .A(n6135), .ZN(n6137) );
  NAND2_X1 U7179 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  NAND2_X1 U7180 ( .A1(n6614), .A2(n8304), .ZN(n6142) );
  NAND2_X1 U7181 ( .A1(n6156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6140) );
  XNOR2_X1 U7182 ( .A(n6140), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7152) );
  AOI22_X1 U7183 ( .A1(n6350), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7022), .B2(
        n7152), .ZN(n6141) );
  NAND2_X1 U7184 ( .A1(n6142), .A2(n6141), .ZN(n10544) );
  XNOR2_X1 U7185 ( .A(n10544), .B(n6478), .ZN(n10559) );
  NAND2_X1 U7186 ( .A1(n6856), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6150) );
  INV_X1 U7187 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7151) );
  OR2_X1 U7188 ( .A1(n6109), .A2(n7151), .ZN(n6149) );
  INV_X1 U7189 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6143) );
  OR2_X1 U7190 ( .A1(n6692), .A2(n6143), .ZN(n6148) );
  AND2_X1 U7191 ( .A1(n6145), .A2(n6144), .ZN(n6146) );
  OR2_X1 U7192 ( .A1(n6146), .A2(n6161), .ZN(n10546) );
  OR2_X1 U7193 ( .A1(n6448), .A2(n10546), .ZN(n6147) );
  NOR2_X1 U7194 ( .A1(n7656), .A2(n6483), .ZN(n6151) );
  NAND2_X1 U7195 ( .A1(n10559), .A2(n6151), .ZN(n6155) );
  INV_X1 U7196 ( .A(n10559), .ZN(n6153) );
  INV_X1 U7197 ( .A(n6151), .ZN(n6152) );
  NAND2_X1 U7198 ( .A1(n6153), .A2(n6152), .ZN(n6154) );
  NAND2_X1 U7199 ( .A1(n6155), .A2(n6154), .ZN(n10541) );
  NAND2_X1 U7200 ( .A1(n10539), .A2(n6155), .ZN(n6172) );
  NAND2_X1 U7201 ( .A1(n6617), .A2(n8304), .ZN(n6159) );
  NOR2_X1 U7202 ( .A1(n6156), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6174) );
  OR2_X1 U7203 ( .A1(n6174), .A2(n6515), .ZN(n6157) );
  XNOR2_X1 U7204 ( .A(n6157), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7153) );
  AOI22_X1 U7205 ( .A1(n6350), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7022), .B2(
        n7153), .ZN(n6158) );
  NAND2_X1 U7206 ( .A1(n6159), .A2(n6158), .ZN(n10555) );
  XNOR2_X1 U7207 ( .A(n10555), .B(n6478), .ZN(n6168) );
  NAND2_X1 U7208 ( .A1(n6855), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6167) );
  INV_X1 U7209 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7132) );
  OR2_X1 U7210 ( .A1(n6160), .A2(n7132), .ZN(n6166) );
  NAND2_X1 U7211 ( .A1(n6161), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6179) );
  OR2_X1 U7212 ( .A1(n6161), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7213 ( .A1(n6179), .A2(n6162), .ZN(n10572) );
  OR2_X1 U7214 ( .A1(n6448), .A2(n10572), .ZN(n6165) );
  INV_X1 U7215 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6163) );
  OR2_X1 U7216 ( .A1(n6692), .A2(n6163), .ZN(n6164) );
  NOR2_X1 U7217 ( .A1(n10538), .A2(n6483), .ZN(n6169) );
  NAND2_X1 U7218 ( .A1(n6168), .A2(n6169), .ZN(n6185) );
  INV_X1 U7219 ( .A(n6168), .ZN(n7372) );
  INV_X1 U7220 ( .A(n6169), .ZN(n6170) );
  NAND2_X1 U7221 ( .A1(n7372), .A2(n6170), .ZN(n6171) );
  AND2_X1 U7222 ( .A1(n6185), .A2(n6171), .ZN(n10562) );
  NAND2_X1 U7223 ( .A1(n6621), .A2(n8304), .ZN(n6176) );
  INV_X1 U7224 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7225 ( .A1(n6174), .A2(n6173), .ZN(n6229) );
  NAND2_X1 U7226 ( .A1(n6229), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6191) );
  XNOR2_X1 U7227 ( .A(n6191), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7154) );
  AOI22_X1 U7228 ( .A1(n6350), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7022), .B2(
        n7154), .ZN(n6175) );
  XNOR2_X1 U7229 ( .A(n10588), .B(n6079), .ZN(n6189) );
  NAND2_X1 U7230 ( .A1(n6856), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6184) );
  INV_X1 U7231 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6177) );
  OR2_X1 U7232 ( .A1(n6692), .A2(n6177), .ZN(n6183) );
  INV_X1 U7233 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7234 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  NAND2_X1 U7235 ( .A1(n6197), .A2(n6180), .ZN(n7596) );
  OR2_X1 U7236 ( .A1(n6448), .A2(n7596), .ZN(n6182) );
  INV_X1 U7237 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7155) );
  OR2_X1 U7238 ( .A1(n6109), .A2(n7155), .ZN(n6181) );
  NOR2_X1 U7239 ( .A1(n10557), .A2(n6483), .ZN(n6187) );
  XNOR2_X1 U7240 ( .A(n6189), .B(n6187), .ZN(n7382) );
  AND2_X1 U7241 ( .A1(n7382), .A2(n6185), .ZN(n6186) );
  INV_X1 U7242 ( .A(n6187), .ZN(n6188) );
  NAND2_X1 U7243 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  NAND2_X1 U7244 ( .A1(n6631), .A2(n8304), .ZN(n6196) );
  NAND2_X1 U7245 ( .A1(n6191), .A2(n6227), .ZN(n6192) );
  NAND2_X1 U7246 ( .A1(n6192), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7247 ( .A1(n6193), .A2(n6226), .ZN(n6210) );
  OR2_X1 U7248 ( .A1(n6193), .A2(n6226), .ZN(n6194) );
  AND2_X1 U7249 ( .A1(n6210), .A2(n6194), .ZN(n7242) );
  AOI22_X1 U7250 ( .A1(n6350), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7242), .B2(
        n7022), .ZN(n6195) );
  NAND2_X1 U7251 ( .A1(n6196), .A2(n6195), .ZN(n10620) );
  XNOR2_X1 U7252 ( .A(n10620), .B(n6478), .ZN(n6204) );
  NAND2_X1 U7253 ( .A1(n6856), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6203) );
  INV_X1 U7254 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7142) );
  OR2_X1 U7255 ( .A1(n6109), .A2(n7142), .ZN(n6202) );
  INV_X1 U7256 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U7257 ( .A1(n6197), .A2(n7234), .ZN(n6198) );
  NAND2_X1 U7258 ( .A1(n6215), .A2(n6198), .ZN(n10624) );
  OR2_X1 U7259 ( .A1(n6448), .A2(n10624), .ZN(n6201) );
  INV_X1 U7260 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6199) );
  OR2_X1 U7261 ( .A1(n6692), .A2(n6199), .ZN(n6200) );
  NOR2_X1 U7262 ( .A1(n7590), .A2(n6483), .ZN(n6205) );
  NAND2_X1 U7263 ( .A1(n6204), .A2(n6205), .ZN(n6209) );
  INV_X1 U7264 ( .A(n6204), .ZN(n7500) );
  INV_X1 U7265 ( .A(n6205), .ZN(n6206) );
  NAND2_X1 U7266 ( .A1(n7500), .A2(n6206), .ZN(n6207) );
  NAND2_X1 U7267 ( .A1(n6209), .A2(n6207), .ZN(n10617) );
  NAND2_X1 U7268 ( .A1(n6633), .A2(n8304), .ZN(n6213) );
  NAND2_X1 U7269 ( .A1(n6210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6211) );
  XNOR2_X1 U7270 ( .A(n6211), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9402) );
  AOI22_X1 U7271 ( .A1(n9402), .A2(n7022), .B1(n6350), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7272 ( .A1(n6213), .A2(n6212), .ZN(n7908) );
  XNOR2_X1 U7273 ( .A(n7908), .B(n6478), .ZN(n6221) );
  NAND2_X1 U7274 ( .A1(n6857), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6220) );
  INV_X1 U7275 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7141) );
  OR2_X1 U7276 ( .A1(n6109), .A2(n7141), .ZN(n6219) );
  INV_X1 U7277 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7136) );
  OR2_X1 U7278 ( .A1(n6160), .A2(n7136), .ZN(n6218) );
  NAND2_X1 U7279 ( .A1(n6215), .A2(n9400), .ZN(n6216) );
  NAND2_X1 U7280 ( .A1(n6245), .A2(n6216), .ZN(n7710) );
  OR2_X1 U7281 ( .A1(n6448), .A2(n7710), .ZN(n6217) );
  NOR2_X1 U7282 ( .A1(n10612), .A2(n6483), .ZN(n6222) );
  NAND2_X1 U7283 ( .A1(n6221), .A2(n6222), .ZN(n6258) );
  INV_X1 U7284 ( .A(n6221), .ZN(n7765) );
  INV_X1 U7285 ( .A(n6222), .ZN(n6223) );
  NAND2_X1 U7286 ( .A1(n7765), .A2(n6223), .ZN(n6224) );
  AND2_X1 U7287 ( .A1(n6258), .A2(n6224), .ZN(n7501) );
  NAND2_X1 U7288 ( .A1(n6654), .A2(n8304), .ZN(n6231) );
  INV_X1 U7289 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6225) );
  NAND3_X1 U7290 ( .A1(n6227), .A2(n6226), .A3(n6225), .ZN(n6228) );
  OR2_X1 U7291 ( .A1(n6229), .A2(n6228), .ZN(n6241) );
  OAI21_X1 U7292 ( .B1(n6241), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6268) );
  XNOR2_X1 U7293 ( .A(n6268), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7362) );
  AOI22_X1 U7294 ( .A1(n7362), .A2(n7022), .B1(n6350), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6230) );
  XNOR2_X1 U7295 ( .A(n8975), .B(n6079), .ZN(n8992) );
  NAND2_X1 U7296 ( .A1(n6857), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6240) );
  INV_X1 U7297 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6232) );
  OR2_X1 U7298 ( .A1(n6160), .A2(n6232), .ZN(n6239) );
  INV_X1 U7299 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6233) );
  OR2_X1 U7300 ( .A1(n6109), .A2(n6233), .ZN(n6238) );
  INV_X1 U7301 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U7302 ( .A1(n6247), .A2(n6235), .ZN(n6236) );
  NAND2_X1 U7303 ( .A1(n6276), .A2(n6236), .ZN(n8973) );
  OR2_X1 U7304 ( .A1(n6448), .A2(n8973), .ZN(n6237) );
  NOR2_X1 U7305 ( .A1(n8991), .A2(n6483), .ZN(n6264) );
  XNOR2_X1 U7306 ( .A(n8992), .B(n6264), .ZN(n6259) );
  INV_X1 U7307 ( .A(n6259), .ZN(n8979) );
  NAND2_X1 U7308 ( .A1(n6638), .A2(n8304), .ZN(n6244) );
  NAND2_X1 U7309 ( .A1(n6241), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6242) );
  XNOR2_X1 U7310 ( .A(n6242), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7204) );
  AOI22_X1 U7311 ( .A1(n6350), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7022), .B2(
        n7204), .ZN(n6243) );
  XNOR2_X1 U7312 ( .A(n7932), .B(n6079), .ZN(n8977) );
  NAND2_X1 U7313 ( .A1(n6855), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6252) );
  INV_X1 U7314 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7930) );
  OR2_X1 U7315 ( .A1(n6160), .A2(n7930), .ZN(n6251) );
  INV_X1 U7316 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U7317 ( .A1(n6245), .A2(n9337), .ZN(n6246) );
  NAND2_X1 U7318 ( .A1(n6247), .A2(n6246), .ZN(n7929) );
  OR2_X1 U7319 ( .A1(n6448), .A2(n7929), .ZN(n6250) );
  INV_X1 U7320 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6248) );
  OR2_X1 U7321 ( .A1(n6692), .A2(n6248), .ZN(n6249) );
  NOR2_X1 U7322 ( .A1(n8976), .A2(n6483), .ZN(n6257) );
  INV_X1 U7323 ( .A(n6257), .ZN(n6253) );
  NAND2_X1 U7324 ( .A1(n8977), .A2(n6253), .ZN(n6254) );
  OR2_X1 U7325 ( .A1(n8979), .A2(n6254), .ZN(n6256) );
  AND2_X1 U7326 ( .A1(n7501), .A2(n6256), .ZN(n6255) );
  NAND2_X1 U7327 ( .A1(n7502), .A2(n6255), .ZN(n6263) );
  INV_X1 U7328 ( .A(n6256), .ZN(n6261) );
  XNOR2_X1 U7329 ( .A(n8977), .B(n6257), .ZN(n7777) );
  AND2_X1 U7330 ( .A1(n7777), .A2(n6258), .ZN(n7771) );
  AND2_X1 U7331 ( .A1(n7771), .A2(n6259), .ZN(n6260) );
  OR2_X1 U7332 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  INV_X1 U7333 ( .A(n6264), .ZN(n6265) );
  NAND2_X1 U7334 ( .A1(n8992), .A2(n6265), .ZN(n6266) );
  NAND2_X1 U7335 ( .A1(n6729), .A2(n8304), .ZN(n6274) );
  INV_X1 U7336 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U7337 ( .A1(n6268), .A2(n6267), .ZN(n6269) );
  NAND2_X1 U7338 ( .A1(n6269), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7339 ( .A1(n6271), .A2(n6270), .ZN(n6285) );
  OR2_X1 U7340 ( .A1(n6271), .A2(n6270), .ZN(n6272) );
  AND2_X1 U7341 ( .A1(n6285), .A2(n6272), .ZN(n7855) );
  AOI22_X1 U7342 ( .A1(n7855), .A2(n7022), .B1(n6350), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6273) );
  XNOR2_X1 U7343 ( .A(n8989), .B(n6079), .ZN(n7743) );
  NAND2_X1 U7344 ( .A1(n6857), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6282) );
  INV_X1 U7345 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7977) );
  OR2_X1 U7346 ( .A1(n6160), .A2(n7977), .ZN(n6281) );
  INV_X1 U7347 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U7348 ( .A1(n6276), .A2(n9325), .ZN(n6277) );
  NAND2_X1 U7349 ( .A1(n6307), .A2(n6277), .ZN(n8983) );
  OR2_X1 U7350 ( .A1(n6448), .A2(n8983), .ZN(n6280) );
  INV_X1 U7351 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6278) );
  OR2_X1 U7352 ( .A1(n6109), .A2(n6278), .ZN(n6279) );
  NOR2_X1 U7353 ( .A1(n8970), .A2(n6483), .ZN(n6283) );
  XNOR2_X1 U7354 ( .A(n7743), .B(n6283), .ZN(n8990) );
  INV_X1 U7355 ( .A(n6283), .ZN(n6284) );
  NAND2_X1 U7356 ( .A1(n6880), .A2(n8304), .ZN(n6288) );
  NAND2_X1 U7357 ( .A1(n6285), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6286) );
  XNOR2_X1 U7358 ( .A(n6286), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9417) );
  AOI22_X1 U7359 ( .A1(n9417), .A2(n7022), .B1(n6350), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6287) );
  XNOR2_X1 U7360 ( .A(n9718), .B(n6079), .ZN(n7836) );
  NAND2_X1 U7361 ( .A1(n6857), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6294) );
  INV_X1 U7362 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6289) );
  OR2_X1 U7363 ( .A1(n6160), .A2(n6289), .ZN(n6293) );
  INV_X1 U7364 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6305) );
  XNOR2_X1 U7365 ( .A(n6307), .B(n6305), .ZN(n8168) );
  OR2_X1 U7366 ( .A1(n6448), .A2(n8168), .ZN(n6292) );
  INV_X1 U7367 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6290) );
  OR2_X1 U7368 ( .A1(n6109), .A2(n6290), .ZN(n6291) );
  NOR2_X1 U7369 ( .A1(n8134), .A2(n6483), .ZN(n6295) );
  XNOR2_X1 U7370 ( .A(n7836), .B(n6295), .ZN(n7742) );
  INV_X1 U7371 ( .A(n6295), .ZN(n6296) );
  NAND2_X1 U7372 ( .A1(n7836), .A2(n6296), .ZN(n6297) );
  NAND2_X1 U7373 ( .A1(n6966), .A2(n8304), .ZN(n6303) );
  NAND2_X1 U7374 ( .A1(n6298), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6299) );
  MUX2_X1 U7375 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6299), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6301) );
  AND2_X1 U7376 ( .A1(n6301), .A2(n6320), .ZN(n7983) );
  AOI22_X1 U7377 ( .A1(n6350), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7022), .B2(
        n7983), .ZN(n6302) );
  XNOR2_X1 U7378 ( .A(n8140), .B(n6079), .ZN(n6316) );
  INV_X1 U7379 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6304) );
  OAI21_X1 U7380 ( .B1(n6307), .B2(n6305), .A(n6304), .ZN(n6308) );
  NAND2_X1 U7381 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n6306) );
  AND2_X1 U7382 ( .A1(n6308), .A2(n6325), .ZN(n8138) );
  NAND2_X1 U7383 ( .A1(n8138), .A2(n6553), .ZN(n6314) );
  NAND2_X1 U7384 ( .A1(n6855), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6313) );
  INV_X1 U7385 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6309) );
  OR2_X1 U7386 ( .A1(n6160), .A2(n6309), .ZN(n6312) );
  INV_X1 U7387 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6310) );
  OR2_X1 U7388 ( .A1(n6692), .A2(n6310), .ZN(n6311) );
  NAND4_X1 U7389 ( .A1(n6314), .A2(n6313), .A3(n6312), .A4(n6311), .ZN(n9368)
         );
  NAND2_X1 U7390 ( .A1(n9368), .A2(n8527), .ZN(n6317) );
  XNOR2_X1 U7391 ( .A(n6316), .B(n6317), .ZN(n7835) );
  INV_X1 U7392 ( .A(n6316), .ZN(n6318) );
  NAND2_X1 U7393 ( .A1(n6318), .A2(n6317), .ZN(n6319) );
  NAND2_X1 U7394 ( .A1(n7001), .A2(n8304), .ZN(n6323) );
  NAND2_X1 U7395 ( .A1(n6320), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6321) );
  XNOR2_X1 U7396 ( .A(n6321), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8016) );
  AOI22_X1 U7397 ( .A1(n6350), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7022), .B2(
        n8016), .ZN(n6322) );
  XNOR2_X1 U7398 ( .A(n9710), .B(n6079), .ZN(n6332) );
  INV_X1 U7399 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U7400 ( .A1(n6325), .A2(n9340), .ZN(n6326) );
  NAND2_X1 U7401 ( .A1(n6354), .A2(n6326), .ZN(n8186) );
  OR2_X1 U7402 ( .A1(n8186), .A2(n6448), .ZN(n6331) );
  INV_X1 U7403 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7993) );
  OR2_X1 U7404 ( .A1(n6109), .A2(n7993), .ZN(n6328) );
  INV_X1 U7405 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8187) );
  OR2_X1 U7406 ( .A1(n6160), .A2(n8187), .ZN(n6327) );
  AND2_X1 U7407 ( .A1(n6328), .A2(n6327), .ZN(n6330) );
  NAND2_X1 U7408 ( .A1(n6857), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6329) );
  AND3_X1 U7409 ( .A1(n6331), .A2(n6330), .A3(n6329), .ZN(n8182) );
  INV_X1 U7410 ( .A(n8182), .ZN(n9625) );
  NAND2_X1 U7411 ( .A1(n9625), .A2(n8527), .ZN(n6333) );
  AND2_X1 U7412 ( .A1(n6332), .A2(n6333), .ZN(n7950) );
  INV_X1 U7413 ( .A(n6332), .ZN(n6335) );
  INV_X1 U7414 ( .A(n6333), .ZN(n6334) );
  NAND2_X1 U7415 ( .A1(n6335), .A2(n6334), .ZN(n7951) );
  NAND2_X1 U7416 ( .A1(n7037), .A2(n8304), .ZN(n6338) );
  XNOR2_X1 U7417 ( .A(n6336), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8119) );
  AOI22_X1 U7418 ( .A1(n6350), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7022), .B2(
        n8119), .ZN(n6337) );
  XNOR2_X1 U7419 ( .A(n9703), .B(n6478), .ZN(n6345) );
  XNOR2_X1 U7420 ( .A(n6354), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n9617) );
  NAND2_X1 U7421 ( .A1(n9617), .A2(n6553), .ZN(n6344) );
  INV_X1 U7422 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6341) );
  NAND2_X1 U7423 ( .A1(n6855), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7424 ( .A1(n6856), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6339) );
  OAI211_X1 U7425 ( .C1(n6341), .C2(n6692), .A(n6340), .B(n6339), .ZN(n6342)
         );
  INV_X1 U7426 ( .A(n6342), .ZN(n6343) );
  NOR2_X1 U7427 ( .A1(n9596), .A2(n6483), .ZN(n6346) );
  AND2_X1 U7428 ( .A1(n6345), .A2(n6346), .ZN(n8085) );
  INV_X1 U7429 ( .A(n6345), .ZN(n6348) );
  INV_X1 U7430 ( .A(n6346), .ZN(n6347) );
  NAND2_X1 U7431 ( .A1(n6348), .A2(n6347), .ZN(n8084) );
  NAND2_X1 U7432 ( .A1(n6349), .A2(n8084), .ZN(n8226) );
  NAND2_X1 U7433 ( .A1(n7331), .A2(n8304), .ZN(n6352) );
  AOI22_X1 U7434 ( .A1(n6350), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8339), .B2(
        n7022), .ZN(n6351) );
  XNOR2_X1 U7435 ( .A(n9700), .B(n6478), .ZN(n6359) );
  INV_X1 U7436 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7998) );
  INV_X1 U7437 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9248) );
  OAI21_X1 U7438 ( .B1(n6354), .B2(n7998), .A(n9248), .ZN(n6355) );
  NAND2_X1 U7439 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n6353) );
  NAND2_X1 U7440 ( .A1(n6355), .A2(n6370), .ZN(n9591) );
  OR2_X1 U7441 ( .A1(n9591), .A2(n6448), .ZN(n6358) );
  AOI22_X1 U7442 ( .A1(n6857), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n6856), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U7443 ( .A1(n6855), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6356) );
  AND3_X1 U7444 ( .A1(n6358), .A2(n6357), .A3(n6356), .ZN(n9428) );
  NOR2_X1 U7445 ( .A1(n9428), .A2(n6483), .ZN(n6360) );
  NAND2_X1 U7446 ( .A1(n6359), .A2(n6360), .ZN(n6365) );
  INV_X1 U7447 ( .A(n6359), .ZN(n8267) );
  INV_X1 U7448 ( .A(n6360), .ZN(n6361) );
  NAND2_X1 U7449 ( .A1(n8267), .A2(n6361), .ZN(n6362) );
  NAND2_X1 U7450 ( .A1(n6365), .A2(n6362), .ZN(n8225) );
  INV_X1 U7451 ( .A(n8225), .ZN(n6363) );
  NAND2_X1 U7452 ( .A1(n7485), .A2(n8304), .ZN(n6368) );
  OR2_X1 U7453 ( .A1(n6366), .A2(n7526), .ZN(n6367) );
  NAND2_X2 U7454 ( .A1(n6368), .A2(n6367), .ZN(n9692) );
  XNOR2_X1 U7455 ( .A(n9692), .B(n6478), .ZN(n6378) );
  NAND2_X1 U7456 ( .A1(n6369), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6385) );
  INV_X1 U7457 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9237) );
  NAND2_X1 U7458 ( .A1(n6370), .A2(n9237), .ZN(n6371) );
  NAND2_X1 U7459 ( .A1(n6385), .A2(n6371), .ZN(n8271) );
  OR2_X1 U7460 ( .A1(n8271), .A2(n6448), .ZN(n6377) );
  INV_X1 U7461 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U7462 ( .A1(n6855), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7463 ( .A1(n6856), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6372) );
  OAI211_X1 U7464 ( .C1(n6374), .C2(n6692), .A(n6373), .B(n6372), .ZN(n6375)
         );
  INV_X1 U7465 ( .A(n6375), .ZN(n6376) );
  AND2_X1 U7466 ( .A1(n6377), .A2(n6376), .ZN(n9598) );
  NOR2_X1 U7467 ( .A1(n9598), .A2(n6483), .ZN(n6379) );
  NAND2_X1 U7468 ( .A1(n6378), .A2(n6379), .ZN(n6382) );
  INV_X1 U7469 ( .A(n6378), .ZN(n9087) );
  INV_X1 U7470 ( .A(n6379), .ZN(n6380) );
  NAND2_X1 U7471 ( .A1(n9087), .A2(n6380), .ZN(n6381) );
  AND2_X1 U7472 ( .A1(n6382), .A2(n6381), .ZN(n8264) );
  NAND2_X1 U7473 ( .A1(n7487), .A2(n8304), .ZN(n6384) );
  INV_X1 U7474 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7488) );
  OR2_X1 U7475 ( .A1(n6366), .A2(n7488), .ZN(n6383) );
  XNOR2_X1 U7476 ( .A(n9687), .B(n6478), .ZN(n6393) );
  INV_X1 U7477 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U7478 ( .A1(n6385), .A2(n9334), .ZN(n6386) );
  AND2_X1 U7479 ( .A1(n6400), .A2(n6386), .ZN(n9566) );
  NAND2_X1 U7480 ( .A1(n9566), .A2(n6553), .ZN(n6392) );
  INV_X1 U7481 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U7482 ( .A1(n6855), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U7483 ( .A1(n6856), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6387) );
  OAI211_X1 U7484 ( .C1(n6389), .C2(n6692), .A(n6388), .B(n6387), .ZN(n6390)
         );
  INV_X1 U7485 ( .A(n6390), .ZN(n6391) );
  NAND2_X1 U7486 ( .A1(n6392), .A2(n6391), .ZN(n9584) );
  AND2_X1 U7487 ( .A1(n9584), .A2(n8527), .ZN(n6394) );
  NAND2_X1 U7488 ( .A1(n6393), .A2(n6394), .ZN(n6408) );
  INV_X1 U7489 ( .A(n6393), .ZN(n9116) );
  INV_X1 U7490 ( .A(n6394), .ZN(n6395) );
  NAND2_X1 U7491 ( .A1(n9116), .A2(n6395), .ZN(n6396) );
  AND2_X1 U7492 ( .A1(n6408), .A2(n6396), .ZN(n9085) );
  NAND2_X1 U7493 ( .A1(n8536), .A2(n8304), .ZN(n6398) );
  OR2_X1 U7494 ( .A1(n6366), .A2(n8539), .ZN(n6397) );
  XNOR2_X1 U7495 ( .A(n9682), .B(n6478), .ZN(n6410) );
  NAND2_X1 U7496 ( .A1(n6399), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6416) );
  INV_X1 U7497 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9352) );
  NAND2_X1 U7498 ( .A1(n6400), .A2(n9352), .ZN(n6401) );
  NAND2_X1 U7499 ( .A1(n6416), .A2(n6401), .ZN(n9119) );
  OR2_X1 U7500 ( .A1(n9119), .A2(n6448), .ZN(n6407) );
  INV_X1 U7501 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U7502 ( .A1(n6856), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6403) );
  NAND2_X1 U7503 ( .A1(n6855), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6402) );
  OAI211_X1 U7504 ( .C1(n6404), .C2(n6692), .A(n6403), .B(n6402), .ZN(n6405)
         );
  INV_X1 U7505 ( .A(n6405), .ZN(n6406) );
  INV_X1 U7506 ( .A(n9092), .ZN(n9571) );
  NAND2_X1 U7507 ( .A1(n9571), .A2(n8527), .ZN(n6411) );
  XNOR2_X1 U7508 ( .A(n6410), .B(n6411), .ZN(n9117) );
  AND2_X1 U7509 ( .A1(n9117), .A2(n6408), .ZN(n6409) );
  INV_X1 U7510 ( .A(n6410), .ZN(n6412) );
  NAND2_X1 U7511 ( .A1(n6412), .A2(n6411), .ZN(n6413) );
  NAND2_X1 U7512 ( .A1(n7780), .A2(n8304), .ZN(n6415) );
  OR2_X1 U7513 ( .A1(n6366), .A2(n7779), .ZN(n6414) );
  XNOR2_X1 U7514 ( .A(n9676), .B(n6478), .ZN(n6424) );
  INV_X1 U7515 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U7516 ( .A1(n6416), .A2(n9247), .ZN(n6417) );
  NAND2_X1 U7517 ( .A1(n6430), .A2(n6417), .ZN(n9080) );
  OR2_X1 U7518 ( .A1(n9080), .A2(n6448), .ZN(n6423) );
  INV_X1 U7519 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U7520 ( .A1(n6856), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U7521 ( .A1(n6855), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6418) );
  OAI211_X1 U7522 ( .C1(n6692), .C2(n6420), .A(n6419), .B(n6418), .ZN(n6421)
         );
  INV_X1 U7523 ( .A(n6421), .ZN(n6422) );
  INV_X1 U7524 ( .A(n9558), .ZN(n9432) );
  NAND2_X1 U7525 ( .A1(n9432), .A2(n8527), .ZN(n9076) );
  INV_X1 U7526 ( .A(n6424), .ZN(n6425) );
  NAND2_X1 U7527 ( .A1(n6426), .A2(n6425), .ZN(n6427) );
  NAND2_X1 U7528 ( .A1(n7841), .A2(n8304), .ZN(n6429) );
  INV_X1 U7529 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7842) );
  OR2_X1 U7530 ( .A1(n6366), .A2(n7842), .ZN(n6428) );
  XNOR2_X1 U7531 ( .A(n9670), .B(n6079), .ZN(n6439) );
  XNOR2_X1 U7532 ( .A(n6440), .B(n6439), .ZN(n9106) );
  INV_X1 U7533 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U7534 ( .A1(n6430), .A2(n9110), .ZN(n6431) );
  AND2_X1 U7535 ( .A1(n6446), .A2(n6431), .ZN(n9522) );
  NAND2_X1 U7536 ( .A1(n9522), .A2(n6553), .ZN(n6437) );
  INV_X1 U7537 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U7538 ( .A1(n6856), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U7539 ( .A1(n6855), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6432) );
  OAI211_X1 U7540 ( .C1(n6692), .C2(n6434), .A(n6433), .B(n6432), .ZN(n6435)
         );
  INV_X1 U7541 ( .A(n6435), .ZN(n6436) );
  OR2_X1 U7542 ( .A1(n9107), .A2(n6483), .ZN(n6438) );
  NAND2_X1 U7543 ( .A1(n8054), .A2(n8304), .ZN(n6443) );
  OR2_X1 U7544 ( .A1(n6366), .A2(n8056), .ZN(n6442) );
  XNOR2_X1 U7545 ( .A(n9667), .B(n6478), .ZN(n6455) );
  INV_X1 U7546 ( .A(n6446), .ZN(n6444) );
  NAND2_X1 U7547 ( .A1(n6444), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6463) );
  INV_X1 U7548 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U7549 ( .A1(n6446), .A2(n6445), .ZN(n6447) );
  NAND2_X1 U7550 ( .A1(n6463), .A2(n6447), .ZN(n9100) );
  OR2_X1 U7551 ( .A1(n9100), .A2(n6448), .ZN(n6454) );
  INV_X1 U7552 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U7553 ( .A1(n6855), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U7554 ( .A1(n6856), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6449) );
  OAI211_X1 U7555 ( .C1(n6451), .C2(n6692), .A(n6450), .B(n6449), .ZN(n6452)
         );
  INV_X1 U7556 ( .A(n6452), .ZN(n6453) );
  NOR2_X1 U7557 ( .A1(n9528), .A2(n6483), .ZN(n6456) );
  NAND2_X1 U7558 ( .A1(n6455), .A2(n6456), .ZN(n6459) );
  INV_X1 U7559 ( .A(n6455), .ZN(n9130) );
  INV_X1 U7560 ( .A(n6456), .ZN(n6457) );
  NAND2_X1 U7561 ( .A1(n9130), .A2(n6457), .ZN(n6458) );
  AND2_X1 U7562 ( .A1(n6459), .A2(n6458), .ZN(n9098) );
  OR2_X1 U7563 ( .A1(n6366), .A2(n8082), .ZN(n6460) );
  XNOR2_X1 U7564 ( .A(n9661), .B(n6478), .ZN(n6471) );
  INV_X1 U7565 ( .A(n6463), .ZN(n6462) );
  NAND2_X1 U7566 ( .A1(n6462), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6492) );
  INV_X1 U7567 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U7568 ( .A1(n6463), .A2(n9361), .ZN(n6464) );
  NAND2_X1 U7569 ( .A1(n6492), .A2(n6464), .ZN(n9495) );
  OR2_X1 U7570 ( .A1(n9495), .A2(n6448), .ZN(n6470) );
  INV_X1 U7571 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7572 ( .A1(n6855), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U7573 ( .A1(n6856), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6465) );
  OAI211_X1 U7574 ( .C1(n6467), .C2(n6692), .A(n6466), .B(n6465), .ZN(n6468)
         );
  INV_X1 U7575 ( .A(n6468), .ZN(n6469) );
  NOR2_X1 U7576 ( .A1(n9479), .A2(n6483), .ZN(n6472) );
  NAND2_X1 U7577 ( .A1(n6471), .A2(n6472), .ZN(n6475) );
  INV_X1 U7578 ( .A(n6471), .ZN(n9068) );
  INV_X1 U7579 ( .A(n6472), .ZN(n6473) );
  NAND2_X1 U7580 ( .A1(n9068), .A2(n6473), .ZN(n6474) );
  NAND2_X1 U7581 ( .A1(n8111), .A2(n8304), .ZN(n6477) );
  OR2_X1 U7582 ( .A1(n6366), .A2(n8112), .ZN(n6476) );
  XNOR2_X1 U7583 ( .A(n9655), .B(n6478), .ZN(n6484) );
  XNOR2_X1 U7584 ( .A(n6492), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9474) );
  INV_X1 U7585 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U7586 ( .A1(n6856), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U7587 ( .A1(n6855), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6479) );
  OAI211_X1 U7588 ( .C1(n6692), .C2(n6481), .A(n6480), .B(n6479), .ZN(n6482)
         );
  AOI21_X1 U7589 ( .B1(n9474), .B2(n6553), .A(n6482), .ZN(n9142) );
  NOR2_X1 U7590 ( .A1(n9142), .A2(n6483), .ZN(n6485) );
  NAND2_X1 U7591 ( .A1(n6484), .A2(n6485), .ZN(n6489) );
  INV_X1 U7592 ( .A(n6484), .ZN(n6487) );
  INV_X1 U7593 ( .A(n6485), .ZN(n6486) );
  NAND2_X1 U7594 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  NAND2_X1 U7595 ( .A1(n9069), .A2(n6489), .ZN(n6502) );
  INV_X1 U7596 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6490) );
  OAI21_X1 U7597 ( .B1(n6492), .B2(n9322), .A(n6490), .ZN(n6493) );
  NAND2_X1 U7598 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6491) );
  OR2_X1 U7599 ( .A1(n6492), .A2(n6491), .ZN(n6548) );
  NAND2_X1 U7600 ( .A1(n9462), .A2(n6553), .ZN(n6499) );
  INV_X1 U7601 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U7602 ( .A1(n6855), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U7603 ( .A1(n6856), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6494) );
  OAI211_X1 U7604 ( .C1(n6496), .C2(n6692), .A(n6495), .B(n6494), .ZN(n6497)
         );
  INV_X1 U7605 ( .A(n6497), .ZN(n6498) );
  INV_X1 U7606 ( .A(n9480), .ZN(n9141) );
  NAND2_X1 U7607 ( .A1(n9141), .A2(n8527), .ZN(n6500) );
  MUX2_X1 U7608 ( .A(n9141), .B(n6500), .S(n6079), .Z(n6501) );
  INV_X1 U7609 ( .A(n6544), .ZN(n6541) );
  INV_X1 U7610 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6511) );
  NAND3_X1 U7611 ( .A1(n6508), .A2(n6535), .A3(n6511), .ZN(n6504) );
  NAND2_X1 U7612 ( .A1(n6513), .A2(n6505), .ZN(n6516) );
  NAND2_X1 U7613 ( .A1(n6516), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6506) );
  MUX2_X1 U7614 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6506), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6507) );
  NAND2_X1 U7615 ( .A1(n6509), .A2(n6508), .ZN(n6510) );
  NAND2_X1 U7616 ( .A1(n6510), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U7617 ( .A1(n6536), .A2(n6535), .ZN(n6538) );
  NAND2_X1 U7618 ( .A1(n6538), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6512) );
  XNOR2_X1 U7619 ( .A(n6512), .B(n6511), .ZN(n7843) );
  INV_X1 U7620 ( .A(n7843), .ZN(n6534) );
  INV_X1 U7621 ( .A(P2_B_REG_SCAN_IN), .ZN(n8311) );
  NOR2_X1 U7622 ( .A1(n6513), .A2(n6515), .ZN(n6514) );
  MUX2_X1 U7623 ( .A(n6515), .B(n6514), .S(P2_IR_REG_25__SCAN_IN), .Z(n6518)
         );
  INV_X1 U7624 ( .A(n6516), .ZN(n6517) );
  OAI221_X1 U7625 ( .B1(n6534), .B2(P2_B_REG_SCAN_IN), .C1(n7843), .C2(n8311), 
        .A(n8055), .ZN(n6519) );
  INV_X1 U7626 ( .A(n6519), .ZN(n6520) );
  INV_X1 U7627 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10422) );
  NAND2_X1 U7628 ( .A1(n10297), .A2(n10422), .ZN(n6522) );
  AND2_X1 U7629 ( .A1(n7843), .A2(n8083), .ZN(n10424) );
  INV_X1 U7630 ( .A(n10424), .ZN(n6521) );
  NAND2_X1 U7631 ( .A1(n6522), .A2(n6521), .ZN(n7451) );
  INV_X1 U7632 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10300) );
  AND2_X1 U7633 ( .A1(n8083), .A2(n8055), .ZN(n10301) );
  AOI21_X1 U7634 ( .B1(n10300), .B2(n10297), .A(n10301), .ZN(n6864) );
  NOR4_X1 U7635 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6526) );
  NOR4_X1 U7636 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6525) );
  NOR4_X1 U7637 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6524) );
  NOR4_X1 U7638 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6523) );
  NAND4_X1 U7639 ( .A1(n6526), .A2(n6525), .A3(n6524), .A4(n6523), .ZN(n6532)
         );
  NOR2_X1 U7640 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6530) );
  NOR4_X1 U7641 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6529) );
  NOR4_X1 U7642 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6528) );
  NOR4_X1 U7643 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6527) );
  NAND4_X1 U7644 ( .A1(n6530), .A2(n6529), .A3(n6528), .A4(n6527), .ZN(n6531)
         );
  OAI21_X1 U7645 ( .B1(n6532), .B2(n6531), .A(n10297), .ZN(n6863) );
  NAND2_X1 U7646 ( .A1(n6864), .A2(n6863), .ZN(n7449) );
  NOR2_X1 U7647 ( .A1(n8083), .A2(n8055), .ZN(n6533) );
  NAND2_X1 U7648 ( .A1(n6534), .A2(n6533), .ZN(n6590) );
  OR2_X1 U7649 ( .A1(n6536), .A2(n6535), .ZN(n6537) );
  AND2_X1 U7650 ( .A1(n6538), .A2(n6537), .ZN(n7021) );
  NOR2_X1 U7651 ( .A1(n7021), .A2(P2_U3152), .ZN(n10423) );
  INV_X1 U7652 ( .A(n7024), .ZN(n7058) );
  NAND3_X1 U7653 ( .A1(n10299), .A2(n10676), .A3(n7058), .ZN(n6540) );
  OR2_X2 U7654 ( .A1(n6557), .A2(n6540), .ZN(n10615) );
  NAND2_X1 U7655 ( .A1(n6541), .A2(n10561), .ZN(n6566) );
  NAND2_X1 U7656 ( .A1(n8195), .A2(n8304), .ZN(n6543) );
  INV_X1 U7657 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8196) );
  OR2_X1 U7658 ( .A1(n6366), .A2(n8196), .ZN(n6542) );
  NAND2_X1 U7659 ( .A1(n6557), .A2(n8524), .ZN(n6545) );
  AND2_X1 U7660 ( .A1(n6545), .A2(n10299), .ZN(n10570) );
  OR2_X1 U7661 ( .A1(n9142), .A2(n9597), .ZN(n6555) );
  INV_X1 U7662 ( .A(n6548), .ZN(n9452) );
  INV_X1 U7663 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U7664 ( .A1(n6856), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U7665 ( .A1(n6855), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6549) );
  OAI211_X1 U7666 ( .C1(n6692), .C2(n6551), .A(n6550), .B(n6549), .ZN(n6552)
         );
  AOI21_X1 U7667 ( .B1(n9452), .B2(n6553), .A(n6552), .ZN(n8330) );
  INV_X1 U7668 ( .A(n9626), .ZN(n9599) );
  OR2_X1 U7669 ( .A1(n8330), .A2(n9599), .ZN(n6554) );
  NAND2_X1 U7670 ( .A1(n6555), .A2(n6554), .ZN(n9467) );
  INV_X1 U7671 ( .A(n9467), .ZN(n6562) );
  NAND2_X1 U7672 ( .A1(n10299), .A2(n5188), .ZN(n6556) );
  NAND2_X1 U7673 ( .A1(n10528), .A2(n8339), .ZN(n7454) );
  NAND2_X1 U7674 ( .A1(n6557), .A2(n7454), .ZN(n7009) );
  AOI21_X1 U7675 ( .B1(n7024), .B2(n8530), .A(n7021), .ZN(n6558) );
  NAND2_X1 U7676 ( .A1(n6590), .A2(n6558), .ZN(n6866) );
  INV_X1 U7677 ( .A(n6866), .ZN(n6559) );
  NAND2_X1 U7678 ( .A1(n7009), .A2(n6559), .ZN(n6560) );
  NAND2_X1 U7679 ( .A1(n6560), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10623) );
  INV_X1 U7680 ( .A(n10623), .ZN(n9121) );
  AOI22_X1 U7681 ( .A1(n9462), .A2(n9121), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6561) );
  OAI21_X1 U7682 ( .B1(n6562), .B2(n9102), .A(n6561), .ZN(n6563) );
  INV_X1 U7683 ( .A(n6563), .ZN(n6564) );
  OAI211_X1 U7684 ( .C1(n6566), .C2(n9650), .A(n6565), .B(n6564), .ZN(P2_U3222) );
  NAND2_X1 U7685 ( .A1(n6567), .A2(n6698), .ZN(n10657) );
  NAND2_X1 U7686 ( .A1(n6568), .A2(n4855), .ZN(n6569) );
  NAND2_X1 U7687 ( .A1(n6569), .A2(n5311), .ZN(P1_U3520) );
  NAND2_X1 U7688 ( .A1(n8762), .A2(n10295), .ZN(n6570) );
  OR2_X1 U7689 ( .A1(n6599), .A2(n6571), .ZN(n6699) );
  NAND2_X1 U7690 ( .A1(n6698), .A2(n10295), .ZN(n6572) );
  NOR2_X1 U7691 ( .A1(n6699), .A2(n6572), .ZN(n6573) );
  NAND2_X1 U7692 ( .A1(n6886), .A2(n6573), .ZN(n7106) );
  INV_X1 U7693 ( .A(n8819), .ZN(n6575) );
  NOR2_X1 U7694 ( .A1(n6852), .A2(n6575), .ZN(n6576) );
  OR2_X1 U7695 ( .A1(n6852), .A2(n7486), .ZN(n6703) );
  INV_X1 U7696 ( .A(n6703), .ZN(n6721) );
  NAND2_X1 U7697 ( .A1(n10163), .A2(n6721), .ZN(n10130) );
  INV_X1 U7698 ( .A(n10160), .ZN(n10128) );
  INV_X1 U7699 ( .A(n6577), .ZN(n6578) );
  AOI22_X1 U7700 ( .A1(n4856), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n10128), .B2(
        n6578), .ZN(n6579) );
  OAI21_X1 U7701 ( .B1(n6580), .B2(n10130), .A(n6579), .ZN(n6581) );
  NAND2_X1 U7702 ( .A1(n6708), .A2(n10095), .ZN(n7249) );
  NAND2_X1 U7703 ( .A1(n6896), .A2(n7249), .ZN(n6583) );
  NAND2_X1 U7704 ( .A1(n10163), .A2(n6583), .ZN(n10134) );
  NAND3_X1 U7705 ( .A1(n5302), .A2(n6585), .A3(n5303), .ZN(P1_U3355) );
  INV_X1 U7706 ( .A(n6586), .ZN(n6587) );
  NOR2_X1 U7707 ( .A1(n6885), .A2(n6587), .ZN(P1_U4006) );
  NAND2_X1 U7708 ( .A1(n8645), .A2(n6885), .ZN(n6588) );
  NAND2_X1 U7709 ( .A1(n6588), .A2(n7781), .ZN(n6667) );
  NAND2_X1 U7710 ( .A1(n6667), .A2(n6646), .ZN(n6589) );
  NAND2_X1 U7711 ( .A1(n6589), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  OR2_X1 U7712 ( .A1(n6590), .A2(P2_U3152), .ZN(n7059) );
  NOR2_X2 U7713 ( .A1(n7059), .A2(n7021), .ZN(n9370) );
  AND2_X1 U7714 ( .A1(n8295), .A2(P2_U3152), .ZN(n6639) );
  NOR2_X1 U7715 ( .A1(n8295), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9740) );
  OAI222_X1 U7716 ( .A1(n4858), .A2(n6591), .B1(n8538), .B2(n6596), .C1(
        P2_U3152), .C2(n7071), .ZN(P2_U3357) );
  OAI222_X1 U7717 ( .A1(n4858), .A2(n6592), .B1(n8538), .B2(n6609), .C1(
        P2_U3152), .C2(n7081), .ZN(P2_U3355) );
  OAI222_X1 U7718 ( .A1(n4858), .A2(n6594), .B1(n8538), .B2(n6605), .C1(
        P2_U3152), .C2(n6593), .ZN(P2_U3356) );
  INV_X1 U7719 ( .A(n7146), .ZN(n7203) );
  OAI222_X1 U7720 ( .A1(n4858), .A2(n6595), .B1(n8538), .B2(n6607), .C1(
        P2_U3152), .C2(n7203), .ZN(P2_U3354) );
  NAND2_X1 U7721 ( .A1(n5356), .A2(P1_U3084), .ZN(n9060) );
  AND2_X1 U7722 ( .A1(n8295), .A2(P1_U3084), .ZN(n10289) );
  OAI222_X1 U7723 ( .A1(n9060), .A2(n6597), .B1(n9064), .B2(n6596), .C1(n6672), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  INV_X1 U7724 ( .A(n10295), .ZN(n6718) );
  NAND2_X1 U7725 ( .A1(n6718), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6598) );
  OAI21_X1 U7726 ( .B1(n6718), .B2(n6599), .A(n6598), .ZN(P1_U3441) );
  INV_X1 U7727 ( .A(n6600), .ZN(n6602) );
  INV_X1 U7728 ( .A(n9060), .ZN(n7038) );
  AOI22_X1 U7729 ( .A1(n10405), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n7038), .ZN(n6601) );
  OAI21_X1 U7730 ( .B1(n6602), .B2(n9064), .A(n6601), .ZN(P1_U3348) );
  INV_X1 U7731 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6603) );
  INV_X1 U7732 ( .A(n7147), .ZN(n7229) );
  OAI222_X1 U7733 ( .A1(n4858), .A2(n6603), .B1(n8538), .B2(n6602), .C1(
        P2_U3152), .C2(n7229), .ZN(P2_U3353) );
  INV_X1 U7734 ( .A(n7038), .ZN(n10286) );
  OAI222_X1 U7735 ( .A1(n6791), .A2(P1_U3084), .B1(n9064), .B2(n6605), .C1(
        n6604), .C2(n10286), .ZN(P1_U3351) );
  OAI222_X1 U7736 ( .A1(n6677), .A2(P1_U3084), .B1(n9064), .B2(n6607), .C1(
        n6606), .C2(n10286), .ZN(P1_U3349) );
  OAI222_X1 U7737 ( .A1(n6748), .A2(P1_U3084), .B1(n9064), .B2(n6609), .C1(
        n6608), .C2(n10286), .ZN(P1_U3350) );
  INV_X1 U7738 ( .A(n10379), .ZN(n6611) );
  INV_X1 U7739 ( .A(n6610), .ZN(n6612) );
  INV_X1 U7740 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7190) );
  OAI222_X1 U7741 ( .A1(n6611), .A2(P1_U3084), .B1(n9064), .B2(n6612), .C1(
        n9060), .C2(n7190), .ZN(P1_U3347) );
  INV_X1 U7742 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6613) );
  INV_X1 U7743 ( .A(n7150), .ZN(n7288) );
  OAI222_X1 U7744 ( .A1(n4858), .A2(n6613), .B1(n8538), .B2(n6612), .C1(
        P2_U3152), .C2(n7288), .ZN(P2_U3352) );
  INV_X1 U7745 ( .A(n6762), .ZN(n6680) );
  INV_X1 U7746 ( .A(n6614), .ZN(n6615) );
  INV_X1 U7747 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6696) );
  OAI222_X1 U7748 ( .A1(n6680), .A2(P1_U3084), .B1(n9064), .B2(n6615), .C1(
        n9060), .C2(n6696), .ZN(P1_U3346) );
  INV_X1 U7749 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6616) );
  INV_X1 U7750 ( .A(n7152), .ZN(n7301) );
  OAI222_X1 U7751 ( .A1(n4858), .A2(n6616), .B1(n8538), .B2(n6615), .C1(
        P2_U3152), .C2(n7301), .ZN(P2_U3351) );
  INV_X1 U7752 ( .A(n6617), .ZN(n6620) );
  INV_X1 U7753 ( .A(n7153), .ZN(n7313) );
  OAI222_X1 U7754 ( .A1(n4858), .A2(n6618), .B1(n8538), .B2(n6620), .C1(
        P2_U3152), .C2(n7313), .ZN(P2_U3350) );
  INV_X1 U7755 ( .A(n6816), .ZN(n6809) );
  OAI222_X1 U7756 ( .A1(n6809), .A2(P1_U3084), .B1(n9064), .B2(n6620), .C1(
        n6619), .C2(n10286), .ZN(P1_U3345) );
  INV_X1 U7757 ( .A(n6621), .ZN(n6623) );
  INV_X1 U7758 ( .A(n7154), .ZN(n9381) );
  OAI222_X1 U7759 ( .A1(n8538), .A2(n6623), .B1(n9381), .B2(P2_U3152), .C1(
        n6622), .C2(n4858), .ZN(P2_U3349) );
  INV_X1 U7760 ( .A(n6841), .ZN(n6819) );
  OAI222_X1 U7761 ( .A1(n6819), .A2(P1_U3084), .B1(n10286), .B2(n5507), .C1(
        n6623), .C2(n9064), .ZN(P1_U3344) );
  INV_X1 U7762 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6630) );
  INV_X1 U7763 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U7764 ( .A1(n6624), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6627) );
  INV_X1 U7765 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6625) );
  OR2_X1 U7766 ( .A1(n4851), .A2(n6625), .ZN(n6626) );
  OAI211_X1 U7767 ( .C1(n5445), .C2(n6628), .A(n6627), .B(n6626), .ZN(n9947)
         );
  NAND2_X1 U7768 ( .A1(n9947), .A2(n4857), .ZN(n6629) );
  OAI21_X1 U7769 ( .B1(n4857), .B2(n6630), .A(n6629), .ZN(P1_U3586) );
  INV_X1 U7770 ( .A(n6631), .ZN(n6636) );
  INV_X1 U7771 ( .A(n7242), .ZN(n7156) );
  OAI222_X1 U7772 ( .A1(n8538), .A2(n6636), .B1(n7156), .B2(P2_U3152), .C1(
        n6632), .C2(n4858), .ZN(P2_U3348) );
  INV_X1 U7773 ( .A(n6633), .ZN(n6637) );
  AOI22_X1 U7774 ( .A1(n9402), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n6639), .ZN(n6634) );
  OAI21_X1 U7775 ( .B1(n6637), .B2(n8538), .A(n6634), .ZN(P2_U3347) );
  INV_X1 U7776 ( .A(n10391), .ZN(n6812) );
  OAI222_X1 U7777 ( .A1(P1_U3084), .A2(n6812), .B1(n9064), .B2(n6636), .C1(
        n6635), .C2(n10286), .ZN(P1_U3343) );
  OAI222_X1 U7778 ( .A1(n6823), .A2(P1_U3084), .B1(n10286), .B2(n5548), .C1(
        n6637), .C2(n9064), .ZN(P1_U3342) );
  INV_X1 U7779 ( .A(n6638), .ZN(n6641) );
  AOI22_X1 U7780 ( .A1(n7204), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n6639), .ZN(n6640) );
  OAI21_X1 U7781 ( .B1(n6641), .B2(n8538), .A(n6640), .ZN(P2_U3346) );
  INV_X1 U7782 ( .A(n7120), .ZN(n6994) );
  OAI222_X1 U7783 ( .A1(n9060), .A2(n6642), .B1(n9064), .B2(n6641), .C1(n6994), 
        .C2(P1_U3084), .ZN(P1_U3341) );
  INV_X1 U7784 ( .A(n7781), .ZN(n6643) );
  NOR2_X1 U7785 ( .A1(n6885), .A2(n6643), .ZN(n6644) );
  OR2_X1 U7786 ( .A1(P1_U3083), .A2(n6644), .ZN(n9929) );
  INV_X1 U7787 ( .A(n9929), .ZN(n10407) );
  NAND2_X1 U7788 ( .A1(n10407), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n6653) );
  OR2_X1 U7789 ( .A1(n5899), .A2(P1_U3084), .ZN(n8178) );
  NOR2_X1 U7790 ( .A1(n8178), .A2(n8821), .ZN(n6645) );
  NAND2_X1 U7791 ( .A1(n6667), .A2(n6645), .ZN(n10395) );
  INV_X1 U7792 ( .A(n6667), .ZN(n6648) );
  OAI21_X1 U7793 ( .B1(n6785), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6920), .ZN(
        n6649) );
  OAI211_X1 U7794 ( .C1(n6649), .C2(n5229), .A(P1_STATE_REG_SCAN_IN), .B(n6646), .ZN(n6647) );
  OAI22_X1 U7795 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(n10395), .B1(n6648), .B2(
        n6647), .ZN(n6651) );
  NAND2_X1 U7796 ( .A1(n6649), .A2(n5229), .ZN(n6788) );
  NAND3_X1 U7797 ( .A1(n6785), .A2(n5229), .A3(n6713), .ZN(n6650) );
  NAND3_X1 U7798 ( .A1(n6651), .A2(n6788), .A3(n6650), .ZN(n6652) );
  OAI211_X1 U7799 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6727), .A(n6653), .B(n6652), .ZN(P1_U3241) );
  INV_X1 U7800 ( .A(n6654), .ZN(n6697) );
  INV_X1 U7801 ( .A(n7362), .ZN(n7358) );
  OAI222_X1 U7802 ( .A1(n8538), .A2(n6697), .B1(n7358), .B2(P2_U3152), .C1(
        n6655), .C2(n4858), .ZN(P2_U3345) );
  NAND2_X1 U7803 ( .A1(n10379), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6663) );
  INV_X1 U7804 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6656) );
  MUX2_X1 U7805 ( .A(n6656), .B(P1_REG2_REG_6__SCAN_IN), .S(n10379), .Z(n6657)
         );
  INV_X1 U7806 ( .A(n6657), .ZN(n10382) );
  NOR2_X1 U7807 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n10405), .ZN(n6662) );
  XNOR2_X1 U7808 ( .A(n6672), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6738) );
  AND2_X1 U7809 ( .A1(n10292), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U7810 ( .A1(n6738), .A2(n6658), .ZN(n6737) );
  INV_X1 U7811 ( .A(n6672), .ZN(n6736) );
  NAND2_X1 U7812 ( .A1(n6736), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U7813 ( .A1(n6737), .A2(n6659), .ZN(n6799) );
  XNOR2_X1 U7814 ( .A(n6791), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6800) );
  INV_X1 U7815 ( .A(n6791), .ZN(n6805) );
  AOI22_X1 U7816 ( .A1(n6799), .A2(n6800), .B1(n6805), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n6752) );
  MUX2_X1 U7817 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6660), .S(n6748), .Z(n6751)
         );
  OR2_X1 U7818 ( .A1(n6752), .A2(n6751), .ZN(n6749) );
  OAI21_X1 U7819 ( .B1(n6748), .B2(n6660), .A(n6749), .ZN(n6779) );
  AOI22_X1 U7820 ( .A1(n6784), .A2(n5385), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n6677), .ZN(n6778) );
  NOR2_X1 U7821 ( .A1(n6779), .A2(n6778), .ZN(n6777) );
  AOI21_X1 U7822 ( .B1(n6677), .B2(n5385), .A(n6777), .ZN(n10409) );
  MUX2_X1 U7823 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7104), .S(n10405), .Z(n6661)
         );
  INV_X1 U7824 ( .A(n6661), .ZN(n10410) );
  NOR2_X1 U7825 ( .A1(n10409), .A2(n10410), .ZN(n10408) );
  NOR2_X1 U7826 ( .A1(n6662), .A2(n10408), .ZN(n10383) );
  NAND2_X1 U7827 ( .A1(n10382), .A2(n10383), .ZN(n10381) );
  NAND2_X1 U7828 ( .A1(n6663), .A2(n10381), .ZN(n6665) );
  MUX2_X1 U7829 ( .A(n7403), .B(P1_REG2_REG_7__SCAN_IN), .S(n6762), .Z(n6664)
         );
  NOR2_X1 U7830 ( .A1(n6665), .A2(n6664), .ZN(n6763) );
  AOI21_X1 U7831 ( .B1(n6665), .B2(n6664), .A(n6763), .ZN(n6686) );
  NAND2_X1 U7832 ( .A1(n8821), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8108) );
  INV_X1 U7833 ( .A(n8108), .ZN(n6666) );
  NAND2_X1 U7834 ( .A1(n6667), .A2(n6666), .ZN(n6827) );
  OR2_X1 U7835 ( .A1(n6827), .A2(n5899), .ZN(n10412) );
  AND2_X1 U7836 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7518) );
  OR2_X1 U7837 ( .A1(n6827), .A2(n6920), .ZN(n9943) );
  NOR2_X1 U7838 ( .A1(n9943), .A2(n6680), .ZN(n6668) );
  AOI211_X1 U7839 ( .C1(n10407), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7518), .B(
        n6668), .ZN(n6685) );
  NAND2_X1 U7840 ( .A1(n10379), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6679) );
  MUX2_X1 U7841 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6669), .S(n10379), .Z(n10385) );
  NAND2_X1 U7842 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n10405), .ZN(n6678) );
  MUX2_X1 U7843 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6670), .S(n10405), .Z(n10415) );
  MUX2_X1 U7844 ( .A(n6671), .B(P1_REG1_REG_1__SCAN_IN), .S(n6672), .Z(n6732)
         );
  AND2_X1 U7845 ( .A1(n10292), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6733) );
  AND2_X1 U7846 ( .A1(n6732), .A2(n6733), .ZN(n6731) );
  NOR2_X1 U7847 ( .A1(n6672), .A2(n6671), .ZN(n6792) );
  MUX2_X1 U7848 ( .A(n6673), .B(P1_REG1_REG_2__SCAN_IN), .S(n6791), .Z(n6674)
         );
  OAI21_X1 U7849 ( .B1(n6731), .B2(n6792), .A(n6674), .ZN(n6797) );
  NAND2_X1 U7850 ( .A1(n6805), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6743) );
  MUX2_X1 U7851 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6676), .S(n6748), .Z(n6744)
         );
  AOI21_X1 U7852 ( .B1(n6797), .B2(n6743), .A(n6744), .ZN(n6675) );
  INV_X1 U7853 ( .A(n6675), .ZN(n6746) );
  OAI21_X1 U7854 ( .B1(n6748), .B2(n6676), .A(n6746), .ZN(n6775) );
  AOI22_X1 U7855 ( .A1(n6784), .A2(n5384), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n6677), .ZN(n6774) );
  NOR2_X1 U7856 ( .A1(n6775), .A2(n6774), .ZN(n6773) );
  AOI21_X1 U7857 ( .B1(n6677), .B2(n5384), .A(n6773), .ZN(n10416) );
  NAND2_X1 U7858 ( .A1(n10415), .A2(n10416), .ZN(n10413) );
  NAND2_X1 U7859 ( .A1(n6678), .A2(n10413), .ZN(n10386) );
  NAND2_X1 U7860 ( .A1(n10385), .A2(n10386), .ZN(n10384) );
  NAND2_X1 U7861 ( .A1(n6679), .A2(n10384), .ZN(n6682) );
  AOI22_X1 U7862 ( .A1(n6762), .A2(n5477), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n6680), .ZN(n6681) );
  NOR2_X1 U7863 ( .A1(n6682), .A2(n6681), .ZN(n6756) );
  AOI21_X1 U7864 ( .B1(n6682), .B2(n6681), .A(n6756), .ZN(n6683) );
  OR2_X1 U7865 ( .A1(n6683), .A2(n10395), .ZN(n6684) );
  OAI211_X1 U7866 ( .C1(n6686), .C2(n10412), .A(n6685), .B(n6684), .ZN(
        P1_U3248) );
  INV_X1 U7867 ( .A(n10557), .ZN(n10608) );
  NAND2_X1 U7868 ( .A1(n9370), .A2(n10608), .ZN(n6687) );
  OAI21_X1 U7869 ( .B1(n9370), .B2(n5507), .A(n6687), .ZN(P2_U3561) );
  INV_X1 U7870 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6694) );
  INV_X1 U7871 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U7872 ( .A1(n6856), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6690) );
  INV_X1 U7873 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6688) );
  OR2_X1 U7874 ( .A1(n6109), .A2(n6688), .ZN(n6689) );
  OAI211_X1 U7875 ( .C1(n6692), .C2(n6691), .A(n6690), .B(n6689), .ZN(n8486)
         );
  NAND2_X1 U7876 ( .A1(n9370), .A2(n8486), .ZN(n6693) );
  OAI21_X1 U7877 ( .B1(n9370), .B2(n6694), .A(n6693), .ZN(P2_U3583) );
  INV_X1 U7878 ( .A(n7656), .ZN(n10558) );
  NAND2_X1 U7879 ( .A1(n9370), .A2(n10558), .ZN(n6695) );
  OAI21_X1 U7880 ( .B1(n9370), .B2(n6696), .A(n6695), .ZN(P2_U3559) );
  INV_X1 U7881 ( .A(n7436), .ZN(n7127) );
  INV_X1 U7882 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6970) );
  OAI222_X1 U7883 ( .A1(n7127), .A2(P1_U3084), .B1(n10286), .B2(n6970), .C1(
        n6697), .C2(n9064), .ZN(P1_U3340) );
  NOR2_X1 U7884 ( .A1(n6699), .A2(n6698), .ZN(n6923) );
  INV_X1 U7885 ( .A(n6923), .ZN(n6719) );
  NAND2_X1 U7886 ( .A1(n10651), .A2(n6719), .ZN(n6700) );
  AND3_X1 U7887 ( .A1(n6700), .A2(n10295), .A3(n6886), .ZN(n6706) );
  INV_X1 U7888 ( .A(n6701), .ZN(n6702) );
  NAND2_X1 U7889 ( .A1(n6702), .A2(n9944), .ZN(n6922) );
  NAND2_X1 U7890 ( .A1(n6922), .A2(n6703), .ZN(n6705) );
  AND2_X1 U7891 ( .A1(n6719), .A2(n10295), .ZN(n6704) );
  NAND2_X1 U7892 ( .A1(n6705), .A2(n6704), .ZN(n6890) );
  NAND2_X1 U7893 ( .A1(n6706), .A2(n6890), .ZN(n6938) );
  INV_X1 U7894 ( .A(n6938), .ZN(n6728) );
  INV_X2 U7895 ( .A(n7514), .ZN(n8234) );
  NAND2_X1 U7896 ( .A1(n9041), .A2(n8819), .ZN(n6707) );
  NAND2_X1 U7897 ( .A1(n4852), .A2(n6712), .ZN(n6711) );
  NOR2_X1 U7898 ( .A1(n6885), .A2(n5229), .ZN(n6709) );
  AOI21_X1 U7899 ( .B1(n6912), .B2(n7040), .A(n6709), .ZN(n6710) );
  AND2_X1 U7900 ( .A1(n6711), .A2(n6710), .ZN(n6717) );
  NAND2_X1 U7901 ( .A1(n6912), .A2(n6712), .ZN(n6716) );
  NOR2_X1 U7902 ( .A1(n6885), .A2(n6713), .ZN(n6714) );
  AOI21_X1 U7903 ( .B1(n4862), .B2(n7040), .A(n6714), .ZN(n6715) );
  NAND2_X1 U7904 ( .A1(n6716), .A2(n6715), .ZN(n6898) );
  NAND2_X1 U7905 ( .A1(n6717), .A2(n6898), .ZN(n6900) );
  OAI21_X1 U7906 ( .B1(n6717), .B2(n6898), .A(n6900), .ZN(n6786) );
  NAND2_X1 U7907 ( .A1(n10651), .A2(n8645), .ZN(n6888) );
  OR2_X1 U7908 ( .A1(n6719), .A2(n6718), .ZN(n6723) );
  OR2_X2 U7909 ( .A1(n6888), .A2(n6723), .ZN(n9879) );
  INV_X1 U7910 ( .A(n9879), .ZN(n9815) );
  NAND2_X1 U7911 ( .A1(n6786), .A2(n9815), .ZN(n6726) );
  INV_X1 U7912 ( .A(n6723), .ZN(n6720) );
  NAND2_X1 U7913 ( .A1(n6721), .A2(n6720), .ZN(n6722) );
  INV_X1 U7914 ( .A(n6922), .ZN(n6850) );
  NOR2_X1 U7915 ( .A1(n6723), .A2(n6920), .ZN(n6724) );
  AOI22_X1 U7916 ( .A1(n7040), .A2(n9863), .B1(n9853), .B2(n6902), .ZN(n6725)
         );
  OAI211_X1 U7917 ( .C1(n6728), .C2(n6727), .A(n6726), .B(n6725), .ZN(P1_U3230) );
  INV_X1 U7918 ( .A(n6729), .ZN(n6742) );
  INV_X1 U7919 ( .A(n7855), .ZN(n7845) );
  INV_X1 U7920 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6730) );
  OAI222_X1 U7921 ( .A1(n8538), .A2(n6742), .B1(n7845), .B2(P2_U3152), .C1(
        n6730), .C2(n4858), .ZN(P2_U3344) );
  INV_X1 U7922 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6741) );
  INV_X1 U7923 ( .A(n9943), .ZN(n10406) );
  INV_X1 U7924 ( .A(n6731), .ZN(n6794) );
  OAI21_X1 U7925 ( .B1(n6733), .B2(n6732), .A(n6794), .ZN(n6734) );
  OAI22_X1 U7926 ( .A1(n10395), .A2(n6734), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5335), .ZN(n6735) );
  AOI21_X1 U7927 ( .B1(n6736), .B2(n10406), .A(n6735), .ZN(n6740) );
  NAND2_X1 U7928 ( .A1(n10292), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6787) );
  INV_X1 U7929 ( .A(n10412), .ZN(n10398) );
  OAI211_X1 U7930 ( .C1(n6738), .C2(n6658), .A(n10398), .B(n6737), .ZN(n6739)
         );
  OAI211_X1 U7931 ( .C1(n9929), .C2(n6741), .A(n6740), .B(n6739), .ZN(P1_U3242) );
  INV_X1 U7932 ( .A(n7731), .ZN(n7721) );
  INV_X1 U7933 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7028) );
  OAI222_X1 U7934 ( .A1(n7721), .A2(P1_U3084), .B1(n10286), .B2(n7028), .C1(
        n6742), .C2(n9064), .ZN(P1_U3339) );
  INV_X1 U7935 ( .A(n10395), .ZN(n10414) );
  NAND3_X1 U7936 ( .A1(n6744), .A2(n6797), .A3(n6743), .ZN(n6745) );
  NAND3_X1 U7937 ( .A1(n10414), .A2(n6746), .A3(n6745), .ZN(n6747) );
  NAND2_X1 U7938 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6919) );
  OAI211_X1 U7939 ( .C1(n9943), .C2(n6748), .A(n6747), .B(n6919), .ZN(n6754)
         );
  INV_X1 U7940 ( .A(n6749), .ZN(n6750) );
  AOI211_X1 U7941 ( .C1(n6752), .C2(n6751), .A(n6750), .B(n10412), .ZN(n6753)
         );
  AOI211_X1 U7942 ( .C1(n10407), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n6754), .B(
        n6753), .ZN(n6755) );
  INV_X1 U7943 ( .A(n6755), .ZN(P1_U3244) );
  NOR2_X1 U7944 ( .A1(n6762), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6757) );
  NOR2_X1 U7945 ( .A1(n6757), .A2(n6756), .ZN(n6759) );
  INV_X1 U7946 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7764) );
  AOI22_X1 U7947 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6809), .B1(n6816), .B2(
        n7764), .ZN(n6758) );
  NOR2_X1 U7948 ( .A1(n6759), .A2(n6758), .ZN(n6808) );
  AOI21_X1 U7949 ( .B1(n6759), .B2(n6758), .A(n6808), .ZN(n6772) );
  INV_X1 U7950 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6760) );
  NOR2_X1 U7951 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6760), .ZN(n7937) );
  INV_X1 U7952 ( .A(n7937), .ZN(n6761) );
  OAI21_X1 U7953 ( .B1(n9943), .B2(n6809), .A(n6761), .ZN(n6770) );
  NOR2_X1 U7954 ( .A1(n6762), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6764) );
  NOR2_X1 U7955 ( .A1(n6764), .A2(n6763), .ZN(n6767) );
  MUX2_X1 U7956 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n5499), .S(n6816), .Z(n6765)
         );
  INV_X1 U7957 ( .A(n6765), .ZN(n6766) );
  NOR2_X1 U7958 ( .A1(n6767), .A2(n6766), .ZN(n6817) );
  AOI21_X1 U7959 ( .B1(n6767), .B2(n6766), .A(n6817), .ZN(n6768) );
  NOR2_X1 U7960 ( .A1(n6768), .A2(n10412), .ZN(n6769) );
  AOI211_X1 U7961 ( .C1(n10407), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n6770), .B(
        n6769), .ZN(n6771) );
  OAI21_X1 U7962 ( .B1(n6772), .B2(n10395), .A(n6771), .ZN(P1_U3249) );
  AOI21_X1 U7963 ( .B1(n6775), .B2(n6774), .A(n6773), .ZN(n6776) );
  NAND2_X1 U7964 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7169) );
  OAI21_X1 U7965 ( .B1(n10395), .B2(n6776), .A(n7169), .ZN(n6783) );
  INV_X1 U7966 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6781) );
  AOI21_X1 U7967 ( .B1(n6779), .B2(n6778), .A(n6777), .ZN(n6780) );
  OAI22_X1 U7968 ( .A1(n9929), .A2(n6781), .B1(n10412), .B2(n6780), .ZN(n6782)
         );
  AOI211_X1 U7969 ( .C1(n6784), .C2(n10406), .A(n6783), .B(n6782), .ZN(n6790)
         );
  MUX2_X1 U7970 ( .A(n6787), .B(n6786), .S(n6785), .Z(n6789) );
  OAI211_X1 U7971 ( .C1(n6789), .C2(n5899), .A(n4857), .B(n6788), .ZN(n6806)
         );
  NAND2_X1 U7972 ( .A1(n6790), .A2(n6806), .ZN(P1_U3245) );
  MUX2_X1 U7973 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6673), .S(n6791), .Z(n6795)
         );
  INV_X1 U7974 ( .A(n6792), .ZN(n6793) );
  NAND3_X1 U7975 ( .A1(n6795), .A2(n6794), .A3(n6793), .ZN(n6796) );
  NAND3_X1 U7976 ( .A1(n10414), .A2(n6797), .A3(n6796), .ZN(n6798) );
  OAI21_X1 U7977 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n5368), .A(n6798), .ZN(n6804) );
  INV_X1 U7978 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6802) );
  XNOR2_X1 U7979 ( .A(n6800), .B(n6799), .ZN(n6801) );
  OAI22_X1 U7980 ( .A1(n9929), .A2(n6802), .B1(n10412), .B2(n6801), .ZN(n6803)
         );
  AOI211_X1 U7981 ( .C1(n6805), .C2(n10406), .A(n6804), .B(n6803), .ZN(n6807)
         );
  NAND2_X1 U7982 ( .A1(n6807), .A2(n6806), .ZN(P1_U3243) );
  AOI21_X1 U7983 ( .B1(n7764), .B2(n6809), .A(n6808), .ZN(n6837) );
  AOI22_X1 U7984 ( .A1(n6841), .A2(n5517), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6819), .ZN(n6836) );
  NOR2_X1 U7985 ( .A1(n6837), .A2(n6836), .ZN(n6835) );
  NOR2_X1 U7986 ( .A1(n6841), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6810) );
  NOR2_X1 U7987 ( .A1(n6835), .A2(n6810), .ZN(n10394) );
  MUX2_X1 U7988 ( .A(n6811), .B(P1_REG1_REG_10__SCAN_IN), .S(n10391), .Z(
        n10393) );
  NOR2_X1 U7989 ( .A1(n10394), .A2(n10393), .ZN(n10392) );
  AOI21_X1 U7990 ( .B1(n6811), .B2(n6812), .A(n10392), .ZN(n6987) );
  NOR2_X1 U7991 ( .A1(n6823), .A2(n5557), .ZN(n6988) );
  AOI21_X1 U7992 ( .B1(n6823), .B2(n5557), .A(n6988), .ZN(n6813) );
  XNOR2_X1 U7993 ( .A(n6987), .B(n6813), .ZN(n6834) );
  NAND2_X1 U7994 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n10391), .ZN(n6820) );
  MUX2_X1 U7995 ( .A(n7493), .B(P1_REG2_REG_10__SCAN_IN), .S(n10391), .Z(n6814) );
  INV_X1 U7996 ( .A(n6814), .ZN(n10399) );
  MUX2_X1 U7997 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n6815), .S(n6841), .Z(n6839)
         );
  NOR2_X1 U7998 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6816), .ZN(n6818) );
  NOR2_X1 U7999 ( .A1(n6818), .A2(n6817), .ZN(n6840) );
  NAND2_X1 U8000 ( .A1(n6839), .A2(n6840), .ZN(n6838) );
  OAI21_X1 U8001 ( .B1(n6819), .B2(n6815), .A(n6838), .ZN(n10400) );
  NAND2_X1 U8002 ( .A1(n10399), .A2(n10400), .ZN(n10397) );
  NAND2_X1 U8003 ( .A1(n6820), .A2(n10397), .ZN(n6826) );
  INV_X1 U8004 ( .A(n6826), .ZN(n6824) );
  OAI21_X1 U8005 ( .B1(n6824), .B2(n6822), .A(n6823), .ZN(n6821) );
  OAI21_X1 U8006 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6826), .A(n6821), .ZN(
        n6997) );
  NAND3_X1 U8007 ( .A1(n6824), .A2(n6823), .A3(n6822), .ZN(n6825) );
  NAND3_X1 U8008 ( .A1(n6997), .A2(n10398), .A3(n6825), .ZN(n6833) );
  NAND2_X1 U8009 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6826), .ZN(n6828) );
  OAI21_X1 U8010 ( .B1(n6828), .B2(n6827), .A(n9943), .ZN(n6831) );
  AND2_X1 U8011 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8074) );
  INV_X1 U8012 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6829) );
  NOR2_X1 U8013 ( .A1(n9929), .A2(n6829), .ZN(n6830) );
  AOI211_X1 U8014 ( .C1(n6986), .C2(n6831), .A(n8074), .B(n6830), .ZN(n6832)
         );
  OAI211_X1 U8015 ( .C1(n6834), .C2(n10395), .A(n6833), .B(n6832), .ZN(
        P1_U3252) );
  AOI21_X1 U8016 ( .B1(n6837), .B2(n6836), .A(n6835), .ZN(n6847) );
  INV_X1 U8017 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6844) );
  OAI211_X1 U8018 ( .C1(n6840), .C2(n6839), .A(n10398), .B(n6838), .ZN(n6843)
         );
  AND2_X1 U8019 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7815) );
  AOI21_X1 U8020 ( .B1(n10406), .B2(n6841), .A(n7815), .ZN(n6842) );
  OAI211_X1 U8021 ( .C1(n9929), .C2(n6844), .A(n6843), .B(n6842), .ZN(n6845)
         );
  INV_X1 U8022 ( .A(n6845), .ZN(n6846) );
  OAI21_X1 U8023 ( .B1(n6847), .B2(n10395), .A(n6846), .ZN(P1_U3250) );
  INV_X1 U8024 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6854) );
  INV_X1 U8025 ( .A(n7252), .ZN(n6848) );
  NAND2_X1 U8026 ( .A1(n6712), .A2(n7257), .ZN(n8775) );
  NAND2_X1 U8027 ( .A1(n6848), .A2(n8775), .ZN(n8652) );
  INV_X1 U8028 ( .A(n6852), .ZN(n6849) );
  NOR2_X1 U8029 ( .A1(n6850), .A2(n6849), .ZN(n6851) );
  AOI22_X1 U8030 ( .A1(n8652), .A2(n6851), .B1(n10146), .B2(n6902), .ZN(n7043)
         );
  OAI21_X1 U8031 ( .B1(n6852), .B2(n7257), .A(n7043), .ZN(n10265) );
  NAND2_X1 U8032 ( .A1(n10265), .A2(n4855), .ZN(n6853) );
  OAI21_X1 U8033 ( .B1(n4855), .B2(n6854), .A(n6853), .ZN(P1_U3454) );
  NAND2_X1 U8034 ( .A1(n6855), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U8035 ( .A1(n6856), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8036 ( .A1(n6857), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6858) );
  AND3_X1 U8037 ( .A1(n6860), .A2(n6859), .A3(n6858), .ZN(n9444) );
  NAND2_X1 U8038 ( .A1(n9143), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6861) );
  OAI21_X1 U8039 ( .B1(n9143), .B2(n9444), .A(n6861), .ZN(P2_U3582) );
  NAND2_X1 U8040 ( .A1(n9143), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n6862) );
  OAI21_X1 U8041 ( .B1(n9143), .B2(n9596), .A(n6862), .ZN(P2_U3570) );
  NAND2_X1 U8042 ( .A1(n6863), .A2(n7454), .ZN(n6865) );
  NOR2_X1 U8043 ( .A1(n6865), .A2(n6864), .ZN(n6877) );
  NOR2_X1 U8044 ( .A1(n7008), .A2(n7451), .ZN(n6867) );
  AND2_X2 U8045 ( .A1(n6877), .A2(n6867), .ZN(n10685) );
  OR2_X1 U8046 ( .A1(n7058), .A2(n8524), .ZN(n6869) );
  NAND2_X1 U8047 ( .A1(n6868), .A2(n6869), .ZN(n7617) );
  NAND3_X1 U8048 ( .A1(n7527), .A2(n8339), .A3(n8537), .ZN(n10477) );
  INV_X1 U8049 ( .A(n6943), .ZN(n7620) );
  NAND2_X1 U8050 ( .A1(n7620), .A2(n7546), .ZN(n8371) );
  NAND2_X1 U8051 ( .A1(n9379), .A2(n4854), .ZN(n8366) );
  AND2_X1 U8052 ( .A1(n8371), .A2(n8366), .ZN(n8494) );
  XOR2_X1 U8053 ( .A(n6945), .B(n8494), .Z(n7542) );
  NAND2_X1 U8054 ( .A1(n8532), .A2(n8339), .ZN(n8490) );
  NAND2_X1 U8055 ( .A1(n7032), .A2(n10468), .ZN(n7530) );
  XOR2_X1 U8056 ( .A(n8494), .B(n7530), .Z(n6871) );
  INV_X1 U8057 ( .A(n6948), .ZN(n6947) );
  AOI222_X1 U8058 ( .A1(n9629), .A2(n6871), .B1(n6947), .B2(n9626), .C1(n6870), 
        .C2(n9624), .ZN(n7549) );
  INV_X1 U8059 ( .A(n7628), .ZN(n6872) );
  AOI21_X1 U8060 ( .B1(n10468), .B2(n7546), .A(n6872), .ZN(n7545) );
  AOI22_X1 U8061 ( .A1(n7545), .A2(n10528), .B1(n10554), .B2(n7546), .ZN(n6873) );
  OAI211_X1 U8062 ( .C1(n10666), .C2(n7542), .A(n7549), .B(n6873), .ZN(n6878)
         );
  NAND2_X1 U8063 ( .A1(n6878), .A2(n10685), .ZN(n6874) );
  OAI21_X1 U8064 ( .B1(n10685), .B2(n7070), .A(n6874), .ZN(P2_U3521) );
  INV_X1 U8065 ( .A(n7451), .ZN(n6875) );
  NOR2_X1 U8066 ( .A1(n6875), .A2(n7008), .ZN(n6876) );
  AND2_X2 U8067 ( .A1(n6877), .A2(n6876), .ZN(n10689) );
  NAND2_X1 U8068 ( .A1(n6878), .A2(n10689), .ZN(n6879) );
  OAI21_X1 U8069 ( .B1(n10689), .B2(n6036), .A(n6879), .ZN(P2_U3454) );
  INV_X1 U8070 ( .A(n6880), .ZN(n6882) );
  OAI222_X1 U8071 ( .A1(n7875), .A2(P1_U3084), .B1(n9064), .B2(n6882), .C1(
        n6881), .C2(n10286), .ZN(P1_U3338) );
  INV_X1 U8072 ( .A(n9417), .ZN(n7856) );
  OAI222_X1 U8073 ( .A1(n4858), .A2(n6883), .B1(n8538), .B2(n6882), .C1(
        P2_U3152), .C2(n7856), .ZN(P2_U3343) );
  NAND2_X1 U8074 ( .A1(n10037), .A2(n4857), .ZN(n6884) );
  OAI21_X1 U8075 ( .B1(n4857), .B2(n7779), .A(n6884), .ZN(P1_U3578) );
  AND3_X1 U8076 ( .A1(n6886), .A2(n6885), .A3(n7781), .ZN(n6887) );
  OAI21_X1 U8077 ( .B1(n6888), .B2(n6923), .A(n6887), .ZN(n6889) );
  NAND2_X1 U8078 ( .A1(n6889), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6891) );
  NAND2_X1 U8079 ( .A1(n6912), .A2(n6892), .ZN(n6894) );
  NAND2_X1 U8080 ( .A1(n4862), .A2(n7275), .ZN(n6893) );
  NAND2_X1 U8081 ( .A1(n6894), .A2(n6893), .ZN(n6897) );
  AOI22_X1 U8082 ( .A1(n9046), .A2(n6892), .B1(n9042), .B2(n7275), .ZN(n7179)
         );
  XNOR2_X1 U8083 ( .A(n7178), .B(n7179), .ZN(n7176) );
  INV_X1 U8084 ( .A(n6898), .ZN(n6899) );
  NAND2_X1 U8085 ( .A1(n6899), .A2(n7173), .ZN(n6901) );
  NAND2_X1 U8086 ( .A1(n6901), .A2(n6900), .ZN(n6907) );
  XNOR2_X1 U8087 ( .A(n6903), .B(n7173), .ZN(n6906) );
  NAND2_X1 U8088 ( .A1(n6907), .A2(n6906), .ZN(n6929) );
  NAND2_X1 U8089 ( .A1(n9046), .A2(n6902), .ZN(n6905) );
  NAND2_X1 U8090 ( .A1(n9042), .A2(n8776), .ZN(n6904) );
  NAND2_X1 U8091 ( .A1(n6905), .A2(n6904), .ZN(n6932) );
  NAND2_X1 U8092 ( .A1(n6929), .A2(n6932), .ZN(n6910) );
  INV_X1 U8093 ( .A(n6906), .ZN(n6909) );
  INV_X1 U8094 ( .A(n6907), .ZN(n6908) );
  NAND2_X1 U8095 ( .A1(n6909), .A2(n6908), .ZN(n6930) );
  NAND2_X1 U8096 ( .A1(n6910), .A2(n6930), .ZN(n6937) );
  XNOR2_X1 U8097 ( .A(n6913), .B(n7173), .ZN(n6916) );
  AOI22_X1 U8098 ( .A1(n9046), .A2(n6914), .B1(n9042), .B2(n6911), .ZN(n6915)
         );
  XNOR2_X1 U8099 ( .A(n6916), .B(n6915), .ZN(n6936) );
  NAND2_X1 U8100 ( .A1(n6916), .A2(n6915), .ZN(n6917) );
  XNOR2_X1 U8101 ( .A(n7176), .B(n7177), .ZN(n6918) );
  NAND2_X1 U8102 ( .A1(n6918), .A2(n9815), .ZN(n6928) );
  INV_X1 U8103 ( .A(n6919), .ZN(n6926) );
  NAND2_X1 U8104 ( .A1(n10295), .A2(n6920), .ZN(n6921) );
  NOR2_X1 U8105 ( .A1(n6922), .A2(n6921), .ZN(n8822) );
  INV_X1 U8106 ( .A(n9873), .ZN(n9851) );
  INV_X1 U8107 ( .A(n6914), .ZN(n6924) );
  INV_X1 U8108 ( .A(n9863), .ZN(n9824) );
  OAI22_X1 U8109 ( .A1(n9851), .A2(n6924), .B1(n10485), .B2(n9824), .ZN(n6925)
         );
  AOI211_X1 U8110 ( .C1(n9853), .C2(n9900), .A(n6926), .B(n6925), .ZN(n6927)
         );
  OAI211_X1 U8111 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9876), .A(n6928), .B(
        n6927), .ZN(P1_U3216) );
  NAND2_X1 U8112 ( .A1(n6930), .A2(n6929), .ZN(n6931) );
  XOR2_X1 U8113 ( .A(n6932), .B(n6931), .Z(n6935) );
  AOI22_X1 U8114 ( .A1(n9873), .A2(n6712), .B1(n9853), .B2(n6914), .ZN(n6934)
         );
  AOI22_X1 U8115 ( .A1(n6938), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9863), .B2(
        n8776), .ZN(n6933) );
  OAI211_X1 U8116 ( .C1(n6935), .C2(n9879), .A(n6934), .B(n6933), .ZN(P1_U3220) );
  XOR2_X1 U8117 ( .A(n6937), .B(n6936), .Z(n6941) );
  AOI22_X1 U8118 ( .A1(n9873), .A2(n6902), .B1(n9853), .B2(n6892), .ZN(n6940)
         );
  AOI22_X1 U8119 ( .A1(n6938), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n9863), .B2(
        n6911), .ZN(n6939) );
  OAI211_X1 U8120 ( .C1(n6941), .C2(n9879), .A(n6940), .B(n6939), .ZN(P1_U3235) );
  NAND2_X1 U8121 ( .A1(n9143), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6942) );
  OAI21_X1 U8122 ( .B1(n8330), .B2(n9143), .A(n6942), .ZN(P2_U3581) );
  NAND2_X1 U8123 ( .A1(n7620), .A2(n4854), .ZN(n6946) );
  AND2_X1 U8124 ( .A1(n6943), .A2(n7546), .ZN(n6944) );
  NAND2_X1 U8125 ( .A1(n6947), .A2(n10478), .ZN(n8368) );
  NAND2_X1 U8126 ( .A1(n8368), .A2(n8377), .ZN(n6952) );
  NAND2_X1 U8127 ( .A1(n7619), .A2(n6952), .ZN(n7618) );
  NAND2_X1 U8128 ( .A1(n6948), .A2(n10478), .ZN(n6949) );
  NAND2_X1 U8129 ( .A1(n7618), .A2(n6949), .ZN(n6950) );
  NAND2_X1 U8130 ( .A1(n7691), .A2(n6960), .ZN(n8378) );
  INV_X1 U8131 ( .A(n7691), .ZN(n9378) );
  NAND2_X1 U8132 ( .A1(n9378), .A2(n10502), .ZN(n8379) );
  NAND2_X1 U8133 ( .A1(n8378), .A2(n8379), .ZN(n8496) );
  NAND2_X1 U8134 ( .A1(n6950), .A2(n8496), .ZN(n7565) );
  OAI21_X1 U8135 ( .B1(n6950), .B2(n8496), .A(n7565), .ZN(n7464) );
  INV_X1 U8136 ( .A(n7464), .ZN(n6962) );
  INV_X1 U8137 ( .A(n8496), .ZN(n8375) );
  NAND2_X1 U8138 ( .A1(n7530), .A2(n8371), .ZN(n6951) );
  NAND2_X1 U8139 ( .A1(n6951), .A2(n8366), .ZN(n7621) );
  INV_X1 U8140 ( .A(n7621), .ZN(n6954) );
  NAND2_X1 U8141 ( .A1(n6954), .A2(n6953), .ZN(n7623) );
  NAND2_X1 U8142 ( .A1(n7623), .A2(n8377), .ZN(n6955) );
  NAND2_X1 U8143 ( .A1(n6955), .A2(n8375), .ZN(n7550) );
  OAI21_X1 U8144 ( .B1(n8375), .B2(n6955), .A(n7550), .ZN(n6958) );
  INV_X1 U8145 ( .A(n9377), .ZN(n10501) );
  OAI22_X1 U8146 ( .A1(n10501), .A2(n9599), .B1(n6948), .B2(n9597), .ZN(n6957)
         );
  NOR2_X1 U8147 ( .A1(n6962), .A2(n7617), .ZN(n6956) );
  AOI211_X1 U8148 ( .C1(n9629), .C2(n6958), .A(n6957), .B(n6956), .ZN(n7466)
         );
  OR2_X1 U8149 ( .A1(n7627), .A2(n10502), .ZN(n6959) );
  NAND2_X1 U8150 ( .A1(n7627), .A2(n10502), .ZN(n7696) );
  AND2_X1 U8151 ( .A1(n6959), .A2(n7696), .ZN(n7460) );
  AOI22_X1 U8152 ( .A1(n7460), .A2(n10528), .B1(n10554), .B2(n6960), .ZN(n6961) );
  OAI211_X1 U8153 ( .C1(n6962), .C2(n10477), .A(n7466), .B(n6961), .ZN(n6964)
         );
  NAND2_X1 U8154 ( .A1(n6964), .A2(n10685), .ZN(n6963) );
  OAI21_X1 U8155 ( .B1(n10685), .B2(n7073), .A(n6963), .ZN(P2_U3523) );
  NAND2_X1 U8156 ( .A1(n6964), .A2(n10689), .ZN(n6965) );
  OAI21_X1 U8157 ( .B1(n10689), .B2(n6074), .A(n6965), .ZN(P2_U3460) );
  INV_X1 U8158 ( .A(n6966), .ZN(n6983) );
  INV_X1 U8159 ( .A(n7983), .ZN(n7849) );
  OAI222_X1 U8160 ( .A1(n8538), .A2(n6983), .B1(n7849), .B2(P2_U3152), .C1(
        n6967), .C2(n4858), .ZN(P2_U3342) );
  INV_X1 U8161 ( .A(n8991), .ZN(n6968) );
  NAND2_X1 U8162 ( .A1(n9370), .A2(n6968), .ZN(n6969) );
  OAI21_X1 U8163 ( .B1(n9370), .B2(n6970), .A(n6969), .ZN(P2_U3565) );
  INV_X1 U8164 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6981) );
  OAI21_X1 U8165 ( .B1(n6972), .B2(n5910), .A(n6971), .ZN(n7328) );
  INV_X1 U8166 ( .A(n7328), .ZN(n6979) );
  OAI21_X1 U8167 ( .B1(n6974), .B2(n8782), .A(n6973), .ZN(n6977) );
  AOI22_X1 U8168 ( .A1(n10146), .A2(n6892), .B1(n10120), .B2(n6902), .ZN(n6975) );
  OAI21_X1 U8169 ( .B1(n6979), .B2(n6896), .A(n6975), .ZN(n6976) );
  AOI21_X1 U8170 ( .B1(n10152), .B2(n6977), .A(n6976), .ZN(n7330) );
  AOI21_X1 U8171 ( .B1(n6911), .B2(n7256), .A(n7269), .ZN(n7323) );
  AOI22_X1 U8172 ( .A1(n7323), .A2(n10250), .B1(n10597), .B2(n6911), .ZN(n6978) );
  OAI211_X1 U8173 ( .C1(n6979), .C2(n10600), .A(n7330), .B(n6978), .ZN(n6984)
         );
  NAND2_X1 U8174 ( .A1(n6984), .A2(n4855), .ZN(n6980) );
  OAI21_X1 U8175 ( .B1(n4855), .B2(n6981), .A(n6980), .ZN(P1_U3460) );
  INV_X1 U8176 ( .A(n9908), .ZN(n7881) );
  OAI222_X1 U8177 ( .A1(P1_U3084), .A2(n7881), .B1(n9064), .B2(n6983), .C1(
        n6982), .C2(n10286), .ZN(P1_U3337) );
  NAND2_X1 U8178 ( .A1(n6984), .A2(n10656), .ZN(n6985) );
  OAI21_X1 U8179 ( .B1(n10656), .B2(n6673), .A(n6985), .ZN(P1_U3525) );
  NAND2_X1 U8180 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8219) );
  OAI22_X1 U8181 ( .A1(n6988), .A2(n6987), .B1(n6986), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n6991) );
  MUX2_X1 U8182 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6989), .S(n7120), .Z(n6990)
         );
  NAND2_X1 U8183 ( .A1(n6990), .A2(n6991), .ZN(n7119) );
  OAI21_X1 U8184 ( .B1(n6991), .B2(n6990), .A(n7119), .ZN(n6992) );
  NAND2_X1 U8185 ( .A1(n10414), .A2(n6992), .ZN(n6993) );
  OAI211_X1 U8186 ( .C1(n9943), .C2(n6994), .A(n8219), .B(n6993), .ZN(n6999)
         );
  NAND2_X1 U8187 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7120), .ZN(n6995) );
  OAI21_X1 U8188 ( .B1(n7120), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6995), .ZN(
        n6996) );
  NOR2_X1 U8189 ( .A1(n6996), .A2(n6997), .ZN(n7113) );
  AOI211_X1 U8190 ( .C1(n6997), .C2(n6996), .A(n7113), .B(n10412), .ZN(n6998)
         );
  AOI211_X1 U8191 ( .C1(n10407), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6999), .B(
        n6998), .ZN(n7000) );
  INV_X1 U8192 ( .A(n7000), .ZN(P1_U3253) );
  INV_X1 U8193 ( .A(n7001), .ZN(n7004) );
  AOI22_X1 U8194 ( .A1(n9919), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7038), .ZN(n7002) );
  OAI21_X1 U8195 ( .B1(n7004), .B2(n9064), .A(n7002), .ZN(P1_U3336) );
  INV_X1 U8196 ( .A(n8016), .ZN(n7992) );
  INV_X1 U8197 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7003) );
  OAI222_X1 U8198 ( .A1(n8538), .A2(n7004), .B1(n7992), .B2(P2_U3152), .C1(
        n7003), .C2(n4858), .ZN(P2_U3341) );
  INV_X1 U8199 ( .A(n7005), .ZN(n10495) );
  AOI211_X1 U8200 ( .C1(n7007), .C2(n7006), .A(n10615), .B(n10495), .ZN(n7012)
         );
  NAND2_X1 U8201 ( .A1(n9137), .A2(n9624), .ZN(n10500) );
  INV_X1 U8202 ( .A(n7008), .ZN(n7453) );
  NAND2_X1 U8203 ( .A1(n7009), .A2(n7453), .ZN(n7031) );
  INV_X1 U8204 ( .A(n7031), .ZN(n7016) );
  OAI22_X1 U8205 ( .A1(n7620), .A2(n10500), .B1(n7016), .B2(n7631), .ZN(n7011)
         );
  NAND2_X1 U8206 ( .A1(n9137), .A2(n9626), .ZN(n10611) );
  OAI22_X1 U8207 ( .A1(n6546), .A2(n10478), .B1(n7691), .B2(n10611), .ZN(n7010) );
  OR3_X1 U8208 ( .A1(n7012), .A2(n7011), .A3(n7010), .ZN(P2_U3239) );
  OAI21_X1 U8209 ( .B1(n7013), .B2(n7015), .A(n7014), .ZN(n7019) );
  OAI22_X1 U8210 ( .A1(n7032), .A2(n10500), .B1(n7016), .B2(n9332), .ZN(n7018)
         );
  OAI22_X1 U8211 ( .A1(n6546), .A2(n4854), .B1(n6948), .B2(n10611), .ZN(n7017)
         );
  AOI211_X1 U8212 ( .C1(n10561), .C2(n7019), .A(n7018), .B(n7017), .ZN(n7020)
         );
  INV_X1 U8213 ( .A(n7020), .ZN(P2_U3224) );
  NAND2_X1 U8214 ( .A1(n7021), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8535) );
  INV_X1 U8215 ( .A(n8535), .ZN(n7023) );
  OAI21_X1 U8216 ( .B1(n10299), .B2(n7023), .A(n7022), .ZN(n7026) );
  NAND2_X1 U8217 ( .A1(n10299), .A2(n7024), .ZN(n7025) );
  NAND2_X1 U8218 ( .A1(n7026), .A2(n7025), .ZN(n10448) );
  NOR2_X1 U8219 ( .A1(n10448), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8220 ( .A(n8970), .ZN(n8173) );
  NAND2_X1 U8221 ( .A1(n9370), .A2(n8173), .ZN(n7027) );
  OAI21_X1 U8222 ( .B1(P2_U3966), .B2(n7028), .A(n7027), .ZN(P2_U3566) );
  INV_X1 U8223 ( .A(n10612), .ZN(n7907) );
  NAND2_X1 U8224 ( .A1(n9370), .A2(n7907), .ZN(n7029) );
  OAI21_X1 U8225 ( .B1(P2_U3966), .B2(n5548), .A(n7029), .ZN(P2_U3563) );
  INV_X1 U8226 ( .A(n9428), .ZN(n9627) );
  NAND2_X1 U8227 ( .A1(n9370), .A2(n9627), .ZN(n7030) );
  OAI21_X1 U8228 ( .B1(P2_U3966), .B2(n5699), .A(n7030), .ZN(P2_U3571) );
  INV_X1 U8229 ( .A(n10611), .ZN(n8984) );
  AOI22_X1 U8230 ( .A1(n8984), .A2(n9379), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n7031), .ZN(n7036) );
  NAND2_X1 U8231 ( .A1(n10561), .A2(n8527), .ZN(n9129) );
  OAI22_X1 U8232 ( .A1(n9129), .A2(n7032), .B1(n7529), .B2(n10615), .ZN(n7034)
         );
  NAND2_X1 U8233 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  OAI211_X1 U8234 ( .C1(n7529), .C2(n6546), .A(n7036), .B(n7035), .ZN(P2_U3234) );
  INV_X1 U8235 ( .A(n7037), .ZN(n7111) );
  AOI22_X1 U8236 ( .A1(n9935), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7038), .ZN(n7039) );
  OAI21_X1 U8237 ( .B1(n7111), .B2(n9064), .A(n7039), .ZN(P1_U3335) );
  AOI22_X1 U8238 ( .A1(n4856), .A2(P1_REG2_REG_0__SCAN_IN), .B1(n10128), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n7042) );
  INV_X1 U8239 ( .A(n10130), .ZN(n10165) );
  OAI21_X1 U8240 ( .B1(n10165), .B2(n10137), .A(n7040), .ZN(n7041) );
  OAI211_X1 U8241 ( .C1(n7043), .C2(n4856), .A(n7042), .B(n7041), .ZN(P1_U3291) );
  INV_X1 U8242 ( .A(n7044), .ZN(n10496) );
  NOR3_X1 U8243 ( .A1(n9129), .A2(n7691), .A3(n7045), .ZN(n7046) );
  AOI21_X1 U8244 ( .B1(n10496), .B2(n10561), .A(n7046), .ZN(n7053) );
  INV_X1 U8245 ( .A(n7699), .ZN(n7049) );
  NAND2_X1 U8246 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7191) );
  OAI21_X1 U8247 ( .B1(n10611), .B2(n9375), .A(n7191), .ZN(n7048) );
  OAI22_X1 U8248 ( .A1(n6546), .A2(n10507), .B1(n7691), .B2(n10500), .ZN(n7047) );
  AOI211_X1 U8249 ( .C1(n7049), .C2(n9121), .A(n7048), .B(n7047), .ZN(n7052)
         );
  INV_X1 U8250 ( .A(n7050), .ZN(n7479) );
  NAND2_X1 U8251 ( .A1(n7479), .A2(n10561), .ZN(n7051) );
  OAI211_X1 U8252 ( .C1(n7054), .C2(n7053), .A(n7052), .B(n7051), .ZN(P2_U3232) );
  INV_X1 U8253 ( .A(n7071), .ZN(n10438) );
  INV_X1 U8254 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7055) );
  MUX2_X1 U8255 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7055), .S(n7071), .Z(n10434)
         );
  NAND2_X1 U8256 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10433) );
  NOR2_X1 U8257 ( .A1(n10434), .A2(n10433), .ZN(n10435) );
  AOI21_X1 U8258 ( .B1(n10438), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10435), .ZN(
        n10452) );
  NAND2_X1 U8259 ( .A1(n10454), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7056) );
  OAI21_X1 U8260 ( .B1(n10454), .B2(P2_REG2_REG_2__SCAN_IN), .A(n7056), .ZN(
        n10451) );
  NOR2_X1 U8261 ( .A1(n10452), .A2(n10451), .ZN(n10450) );
  AOI21_X1 U8262 ( .B1(n10454), .B2(P2_REG2_REG_2__SCAN_IN), .A(n10450), .ZN(
        n7066) );
  NAND2_X1 U8263 ( .A1(n7143), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7057) );
  OAI21_X1 U8264 ( .B1(n7143), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7057), .ZN(
        n7065) );
  NOR2_X1 U8265 ( .A1(n7066), .A2(n7065), .ZN(n7129) );
  NAND2_X1 U8266 ( .A1(n10299), .A2(n7058), .ZN(n7061) );
  AND2_X1 U8267 ( .A1(n7059), .A2(n8535), .ZN(n7060) );
  NAND2_X1 U8268 ( .A1(n7061), .A2(n7060), .ZN(n7076) );
  NAND2_X1 U8269 ( .A1(n7076), .A2(n7074), .ZN(n7062) );
  NAND2_X1 U8270 ( .A1(n9143), .A2(n7062), .ZN(n7067) );
  NOR2_X1 U8271 ( .A1(n6547), .A2(n7063), .ZN(n7064) );
  NAND2_X1 U8272 ( .A1(n7067), .A2(n7064), .ZN(n10449) );
  AOI211_X1 U8273 ( .C1(n7066), .C2(n7065), .A(n7129), .B(n10449), .ZN(n7083)
         );
  INV_X1 U8274 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10499) );
  NOR2_X1 U8275 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10499), .ZN(n7068) );
  AOI21_X1 U8276 ( .B1(n10448), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7068), .ZN(
        n7080) );
  NAND2_X1 U8277 ( .A1(n10454), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7072) );
  MUX2_X1 U8278 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7069), .S(n10454), .Z(n10459) );
  MUX2_X1 U8279 ( .A(n7070), .B(P2_REG1_REG_1__SCAN_IN), .S(n7071), .Z(n10444)
         );
  NAND3_X1 U8280 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n10444), .ZN(n10443) );
  OAI21_X1 U8281 ( .B1(n7071), .B2(n7070), .A(n10443), .ZN(n10458) );
  NAND2_X1 U8282 ( .A1(n10459), .A2(n10458), .ZN(n10456) );
  NAND2_X1 U8283 ( .A1(n7072), .A2(n10456), .ZN(n7078) );
  MUX2_X1 U8284 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7073), .S(n7143), .Z(n7077)
         );
  AND2_X1 U8285 ( .A1(n7063), .A2(n7074), .ZN(n7075) );
  NAND2_X1 U8286 ( .A1(n7076), .A2(n7075), .ZN(n10427) );
  INV_X1 U8287 ( .A(n10427), .ZN(n10457) );
  NAND2_X1 U8288 ( .A1(n7077), .A2(n7078), .ZN(n7144) );
  OAI211_X1 U8289 ( .C1(n7078), .C2(n7077), .A(n10457), .B(n7144), .ZN(n7079)
         );
  OAI211_X1 U8290 ( .C1(n10426), .C2(n7081), .A(n7080), .B(n7079), .ZN(n7082)
         );
  OR2_X1 U8291 ( .A1(n7083), .A2(n7082), .ZN(P2_U3248) );
  INV_X1 U8292 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7097) );
  OAI21_X1 U8293 ( .B1(n7085), .B2(n7088), .A(n7084), .ZN(n7320) );
  INV_X1 U8294 ( .A(n7320), .ZN(n7095) );
  INV_X1 U8295 ( .A(n6896), .ZN(n10604) );
  INV_X1 U8296 ( .A(n9899), .ZN(n7414) );
  INV_X1 U8297 ( .A(n6892), .ZN(n7086) );
  OAI22_X1 U8298 ( .A1(n7414), .A2(n10111), .B1(n10149), .B2(n7086), .ZN(n7092) );
  NAND2_X1 U8299 ( .A1(n7264), .A2(n7265), .ZN(n7263) );
  NAND2_X1 U8300 ( .A1(n7263), .A2(n8785), .ZN(n7087) );
  NAND2_X1 U8301 ( .A1(n7087), .A2(n8656), .ZN(n7090) );
  NAND3_X1 U8302 ( .A1(n7263), .A2(n8785), .A3(n7088), .ZN(n7089) );
  INV_X1 U8303 ( .A(n10152), .ZN(n10107) );
  AOI21_X1 U8304 ( .B1(n7090), .B2(n7089), .A(n10107), .ZN(n7091) );
  AOI211_X1 U8305 ( .C1(n10604), .C2(n7320), .A(n7092), .B(n7091), .ZN(n7322)
         );
  INV_X1 U8306 ( .A(n7105), .ZN(n7093) );
  AOI21_X1 U8307 ( .B1(n7175), .B2(n7271), .A(n7093), .ZN(n7314) );
  AOI22_X1 U8308 ( .A1(n7314), .A2(n10250), .B1(n10597), .B2(n7175), .ZN(n7094) );
  OAI211_X1 U8309 ( .C1(n7095), .C2(n10600), .A(n7322), .B(n7094), .ZN(n7098)
         );
  NAND2_X1 U8310 ( .A1(n7098), .A2(n4855), .ZN(n7096) );
  OAI21_X1 U8311 ( .B1(n4855), .B2(n7097), .A(n7096), .ZN(P1_U3466) );
  NAND2_X1 U8312 ( .A1(n7098), .A2(n10656), .ZN(n7099) );
  OAI21_X1 U8313 ( .B1(n10656), .B2(n5384), .A(n7099), .ZN(P1_U3527) );
  OAI21_X1 U8314 ( .B1(n7101), .B2(n5916), .A(n7100), .ZN(n10517) );
  XNOR2_X1 U8315 ( .A(n7102), .B(n8653), .ZN(n7103) );
  AOI222_X1 U8316 ( .A1(n10152), .A2(n7103), .B1(n9898), .B2(n10146), .C1(
        n9900), .C2(n10120), .ZN(n10516) );
  MUX2_X1 U8317 ( .A(n7104), .B(n10516), .S(n10163), .Z(n7110) );
  AOI211_X1 U8318 ( .C1(n10514), .C2(n7105), .A(n10633), .B(n7421), .ZN(n10513) );
  NOR2_X1 U8319 ( .A1(n7106), .A2(n10095), .ZN(n10117) );
  INV_X1 U8320 ( .A(n7107), .ZN(n7353) );
  OAI22_X1 U8321 ( .A1(n10130), .A2(n7337), .B1(n10160), .B2(n7353), .ZN(n7108) );
  AOI21_X1 U8322 ( .B1(n10513), .B2(n10117), .A(n7108), .ZN(n7109) );
  OAI211_X1 U8323 ( .C1(n10134), .C2(n10517), .A(n7110), .B(n7109), .ZN(
        P1_U3286) );
  INV_X1 U8324 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7112) );
  INV_X1 U8325 ( .A(n8119), .ZN(n8116) );
  OAI222_X1 U8326 ( .A1(n4858), .A2(n7112), .B1(n8538), .B2(n7111), .C1(
        P2_U3152), .C2(n8116), .ZN(P2_U3340) );
  AOI21_X1 U8327 ( .B1(n7120), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7113), .ZN(
        n7116) );
  NAND2_X1 U8328 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7436), .ZN(n7114) );
  OAI21_X1 U8329 ( .B1(n7436), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7114), .ZN(
        n7115) );
  NOR2_X1 U8330 ( .A1(n7116), .A2(n7115), .ZN(n7431) );
  AOI211_X1 U8331 ( .C1(n7116), .C2(n7115), .A(n7431), .B(n10412), .ZN(n7117)
         );
  AOI21_X1 U8332 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n10407), .A(n7117), .ZN(
        n7126) );
  XNOR2_X1 U8333 ( .A(n7436), .B(n7118), .ZN(n7122) );
  OAI21_X1 U8334 ( .B1(n7120), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7119), .ZN(
        n7121) );
  NAND2_X1 U8335 ( .A1(n7122), .A2(n7121), .ZN(n7435) );
  OAI21_X1 U8336 ( .B1(n7122), .B2(n7121), .A(n7435), .ZN(n7124) );
  NAND2_X1 U8337 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8241) );
  INV_X1 U8338 ( .A(n8241), .ZN(n7123) );
  AOI21_X1 U8339 ( .B1(n10414), .B2(n7124), .A(n7123), .ZN(n7125) );
  OAI211_X1 U8340 ( .C1(n7127), .C2(n9943), .A(n7126), .B(n7125), .ZN(P1_U3254) );
  OR2_X1 U8341 ( .A1(n9402), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7137) );
  INV_X1 U8342 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7683) );
  INV_X1 U8343 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7131) );
  INV_X1 U8344 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7128) );
  MUX2_X1 U8345 ( .A(n7128), .B(P2_REG2_REG_4__SCAN_IN), .S(n7146), .Z(n7198)
         );
  AOI21_X1 U8346 ( .B1(n7143), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7129), .ZN(
        n7199) );
  NOR2_X1 U8347 ( .A1(n7198), .A2(n7199), .ZN(n7197) );
  AOI21_X1 U8348 ( .B1(n7146), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7197), .ZN(
        n7224) );
  NAND2_X1 U8349 ( .A1(n7147), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7130) );
  OAI21_X1 U8350 ( .B1(n7147), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7130), .ZN(
        n7223) );
  OR2_X1 U8351 ( .A1(n7224), .A2(n7223), .ZN(n7226) );
  OAI21_X1 U8352 ( .B1(n7229), .B2(n7131), .A(n7226), .ZN(n7284) );
  MUX2_X1 U8353 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7659), .S(n7150), .Z(n7285)
         );
  NAND2_X1 U8354 ( .A1(n7284), .A2(n7285), .ZN(n7283) );
  OAI21_X1 U8355 ( .B1(n7288), .B2(n7659), .A(n7283), .ZN(n7297) );
  MUX2_X1 U8356 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7683), .S(n7152), .Z(n7298)
         );
  NAND2_X1 U8357 ( .A1(n7297), .A2(n7298), .ZN(n7296) );
  OAI21_X1 U8358 ( .B1(n7683), .B2(n7301), .A(n7296), .ZN(n7309) );
  MUX2_X1 U8359 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7132), .S(n7153), .Z(n7310)
         );
  NAND2_X1 U8360 ( .A1(n7309), .A2(n7310), .ZN(n7308) );
  OAI21_X1 U8361 ( .B1(n7132), .B2(n7313), .A(n7308), .ZN(n9386) );
  INV_X1 U8362 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7133) );
  MUX2_X1 U8363 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7133), .S(n7154), .Z(n9387)
         );
  AND2_X1 U8364 ( .A1(n9386), .A2(n9387), .ZN(n9384) );
  AOI21_X1 U8365 ( .B1(n7154), .B2(P2_REG2_REG_9__SCAN_IN), .A(n9384), .ZN(
        n7239) );
  INV_X1 U8366 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7134) );
  MUX2_X1 U8367 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7134), .S(n7242), .Z(n7135)
         );
  INV_X1 U8368 ( .A(n7135), .ZN(n7238) );
  NOR2_X1 U8369 ( .A1(n7239), .A2(n7238), .ZN(n7237) );
  AOI21_X1 U8370 ( .B1(n7242), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7237), .ZN(
        n9397) );
  MUX2_X1 U8371 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7136), .S(n9402), .Z(n9398)
         );
  NAND2_X1 U8372 ( .A1(n9397), .A2(n9398), .ZN(n9396) );
  NAND2_X1 U8373 ( .A1(n7137), .A2(n9396), .ZN(n7212) );
  MUX2_X1 U8374 ( .A(n7930), .B(P2_REG2_REG_12__SCAN_IN), .S(n7204), .Z(n7211)
         );
  NAND2_X1 U8375 ( .A1(n7204), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7138) );
  AOI22_X1 U8376 ( .A1(n7362), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n6232), .B2(
        n7358), .ZN(n7139) );
  NAND2_X1 U8377 ( .A1(n7140), .A2(n7139), .ZN(n7361) );
  OAI21_X1 U8378 ( .B1(n7140), .B2(n7139), .A(n7361), .ZN(n7166) );
  AOI22_X1 U8379 ( .A1(n7362), .A2(n6233), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7358), .ZN(n7161) );
  NAND2_X1 U8380 ( .A1(n9402), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7157) );
  MUX2_X1 U8381 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7141), .S(n9402), .Z(n9404)
         );
  MUX2_X1 U8382 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7142), .S(n7242), .Z(n7244)
         );
  NAND2_X1 U8383 ( .A1(n7147), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7149) );
  NAND2_X1 U8384 ( .A1(n7143), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7145) );
  AND2_X1 U8385 ( .A1(n7145), .A2(n7144), .ZN(n7194) );
  MUX2_X1 U8386 ( .A(n6092), .B(P2_REG1_REG_4__SCAN_IN), .S(n7146), .Z(n7193)
         );
  NOR2_X1 U8387 ( .A1(n7194), .A2(n7193), .ZN(n7192) );
  AOI21_X1 U8388 ( .B1(n7146), .B2(P2_REG1_REG_4__SCAN_IN), .A(n7192), .ZN(
        n7219) );
  MUX2_X1 U8389 ( .A(n6108), .B(P2_REG1_REG_5__SCAN_IN), .S(n7147), .Z(n7218)
         );
  OR2_X1 U8390 ( .A1(n7219), .A2(n7218), .ZN(n7148) );
  AND2_X1 U8391 ( .A1(n7149), .A2(n7148), .ZN(n7280) );
  MUX2_X1 U8392 ( .A(n6127), .B(P2_REG1_REG_6__SCAN_IN), .S(n7150), .Z(n7279)
         );
  NOR2_X1 U8393 ( .A1(n7280), .A2(n7279), .ZN(n7291) );
  NOR2_X1 U8394 ( .A1(n7288), .A2(n6127), .ZN(n7290) );
  MUX2_X1 U8395 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7151), .S(n7152), .Z(n7289)
         );
  OAI21_X1 U8396 ( .B1(n7291), .B2(n7290), .A(n7289), .ZN(n7304) );
  NAND2_X1 U8397 ( .A1(n7152), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7303) );
  INV_X1 U8398 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10578) );
  MUX2_X1 U8399 ( .A(n10578), .B(P2_REG1_REG_8__SCAN_IN), .S(n7153), .Z(n7302)
         );
  AOI21_X1 U8400 ( .B1(n7304), .B2(n7303), .A(n7302), .ZN(n9390) );
  NOR2_X1 U8401 ( .A1(n7313), .A2(n10578), .ZN(n9389) );
  MUX2_X1 U8402 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7155), .S(n7154), .Z(n9388)
         );
  OAI21_X1 U8403 ( .B1(n9390), .B2(n9389), .A(n9388), .ZN(n9392) );
  OAI21_X1 U8404 ( .B1(n7155), .B2(n9381), .A(n9392), .ZN(n7245) );
  NAND2_X1 U8405 ( .A1(n7244), .A2(n7245), .ZN(n7243) );
  OAI21_X1 U8406 ( .B1(n7156), .B2(n7142), .A(n7243), .ZN(n9405) );
  NAND2_X1 U8407 ( .A1(n9404), .A2(n9405), .ZN(n9403) );
  NAND2_X1 U8408 ( .A1(n7157), .A2(n9403), .ZN(n7206) );
  INV_X1 U8409 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7158) );
  MUX2_X1 U8410 ( .A(n7158), .B(P2_REG1_REG_12__SCAN_IN), .S(n7204), .Z(n7205)
         );
  OR2_X1 U8411 ( .A1(n7204), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7159) );
  NOR2_X1 U8412 ( .A1(n7160), .A2(n7161), .ZN(n7357) );
  AOI21_X1 U8413 ( .B1(n7161), .B2(n7160), .A(n7357), .ZN(n7163) );
  NAND2_X1 U8414 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8969) );
  NAND2_X1 U8415 ( .A1(n10448), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7162) );
  OAI211_X1 U8416 ( .C1(n10427), .C2(n7163), .A(n8969), .B(n7162), .ZN(n7165)
         );
  NOR2_X1 U8417 ( .A1(n10426), .A2(n7358), .ZN(n7164) );
  AOI211_X1 U8418 ( .C1(n10425), .C2(n7166), .A(n7165), .B(n7164), .ZN(n7167)
         );
  INV_X1 U8419 ( .A(n7167), .ZN(P2_U3258) );
  INV_X1 U8420 ( .A(n7168), .ZN(n7315) );
  INV_X1 U8421 ( .A(n9876), .ZN(n9806) );
  NAND2_X1 U8422 ( .A1(n9873), .A2(n6892), .ZN(n7172) );
  INV_X1 U8423 ( .A(n7169), .ZN(n7170) );
  AOI21_X1 U8424 ( .B1(n9853), .B2(n9899), .A(n7170), .ZN(n7171) );
  OAI211_X1 U8425 ( .C1(n7318), .C2(n9824), .A(n7172), .B(n7171), .ZN(n7187)
         );
  AOI22_X1 U8426 ( .A1(n9042), .A2(n9900), .B1(n8234), .B2(n7175), .ZN(n7174)
         );
  BUF_X4 U8427 ( .A(n7173), .Z(n8946) );
  XNOR2_X1 U8428 ( .A(n7174), .B(n8946), .ZN(n7333) );
  AOI22_X1 U8429 ( .A1(n9046), .A2(n9900), .B1(n9042), .B2(n7175), .ZN(n7332)
         );
  XNOR2_X1 U8430 ( .A(n7333), .B(n7332), .ZN(n7185) );
  INV_X1 U8431 ( .A(n7178), .ZN(n7180) );
  NAND2_X1 U8432 ( .A1(n7180), .A2(n7179), .ZN(n7181) );
  INV_X1 U8433 ( .A(n7335), .ZN(n7183) );
  AOI211_X1 U8434 ( .C1(n7185), .C2(n7184), .A(n9879), .B(n7183), .ZN(n7186)
         );
  AOI211_X1 U8435 ( .C1(n7315), .C2(n9806), .A(n7187), .B(n7186), .ZN(n7188)
         );
  INV_X1 U8436 ( .A(n7188), .ZN(P1_U3228) );
  NAND2_X1 U8437 ( .A1(P2_U3966), .A2(n10536), .ZN(n7189) );
  OAI21_X1 U8438 ( .B1(n9370), .B2(n7190), .A(n7189), .ZN(P2_U3558) );
  INV_X1 U8439 ( .A(n7191), .ZN(n7196) );
  AOI211_X1 U8440 ( .C1(n7194), .C2(n7193), .A(n7192), .B(n10427), .ZN(n7195)
         );
  AOI211_X1 U8441 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10448), .A(n7196), .B(
        n7195), .ZN(n7202) );
  AOI211_X1 U8442 ( .C1(n7199), .C2(n7198), .A(n7197), .B(n10449), .ZN(n7200)
         );
  INV_X1 U8443 ( .A(n7200), .ZN(n7201) );
  OAI211_X1 U8444 ( .C1(n10426), .C2(n7203), .A(n7202), .B(n7201), .ZN(
        P2_U3249) );
  INV_X1 U8445 ( .A(n7204), .ZN(n7217) );
  NAND2_X1 U8446 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7768) );
  INV_X1 U8447 ( .A(n7768), .ZN(n7210) );
  NAND2_X1 U8448 ( .A1(n7206), .A2(n7205), .ZN(n7207) );
  AOI21_X1 U8449 ( .B1(n7208), .B2(n7207), .A(n10427), .ZN(n7209) );
  AOI211_X1 U8450 ( .C1(P2_ADDR_REG_12__SCAN_IN), .C2(n10448), .A(n7210), .B(
        n7209), .ZN(n7216) );
  NAND2_X1 U8451 ( .A1(n7212), .A2(n7211), .ZN(n7213) );
  NAND3_X1 U8452 ( .A1(n10425), .A2(n7214), .A3(n7213), .ZN(n7215) );
  OAI211_X1 U8453 ( .C1(n10426), .C2(n7217), .A(n7216), .B(n7215), .ZN(
        P2_U3257) );
  NAND2_X1 U8454 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7473) );
  INV_X1 U8455 ( .A(n7473), .ZN(n7222) );
  XNOR2_X1 U8456 ( .A(n7219), .B(n7218), .ZN(n7220) );
  NOR2_X1 U8457 ( .A1(n10427), .A2(n7220), .ZN(n7221) );
  AOI211_X1 U8458 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n10448), .A(n7222), .B(
        n7221), .ZN(n7228) );
  NAND2_X1 U8459 ( .A1(n7224), .A2(n7223), .ZN(n7225) );
  NAND3_X1 U8460 ( .A1(n10425), .A2(n7226), .A3(n7225), .ZN(n7227) );
  OAI211_X1 U8461 ( .C1(n10426), .C2(n7229), .A(n7228), .B(n7227), .ZN(
        P2_U3250) );
  INV_X1 U8462 ( .A(n9107), .ZN(n9536) );
  NAND2_X1 U8463 ( .A1(n9536), .A2(P2_U3966), .ZN(n7230) );
  OAI21_X1 U8464 ( .B1(n5788), .B2(P2_U3966), .A(n7230), .ZN(P2_U3576) );
  INV_X1 U8465 ( .A(n9479), .ZN(n9436) );
  NAND2_X1 U8466 ( .A1(n9436), .A2(P2_U3966), .ZN(n7231) );
  OAI21_X1 U8467 ( .B1(n5828), .B2(P2_U3966), .A(n7231), .ZN(P2_U3578) );
  INV_X1 U8468 ( .A(n9528), .ZN(n9133) );
  NAND2_X1 U8469 ( .A1(n9133), .A2(P2_U3966), .ZN(n7232) );
  OAI21_X1 U8470 ( .B1(n5807), .B2(P2_U3966), .A(n7232), .ZN(P2_U3577) );
  INV_X1 U8471 ( .A(n9598), .ZN(n9570) );
  NAND2_X1 U8472 ( .A1(n9570), .A2(P2_U3966), .ZN(n7233) );
  OAI21_X1 U8473 ( .B1(n9370), .B2(n5725), .A(n7233), .ZN(P2_U3572) );
  NOR2_X1 U8474 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7234), .ZN(n7235) );
  AOI21_X1 U8475 ( .B1(n10448), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7235), .ZN(
        n7236) );
  INV_X1 U8476 ( .A(n7236), .ZN(n7241) );
  AOI211_X1 U8477 ( .C1(n7239), .C2(n7238), .A(n7237), .B(n10449), .ZN(n7240)
         );
  AOI211_X1 U8478 ( .C1(n10455), .C2(n7242), .A(n7241), .B(n7240), .ZN(n7247)
         );
  OAI211_X1 U8479 ( .C1(n7245), .C2(n7244), .A(n10457), .B(n7243), .ZN(n7246)
         );
  NAND2_X1 U8480 ( .A1(n7247), .A2(n7246), .ZN(P2_U3255) );
  INV_X1 U8481 ( .A(n7251), .ZN(n8650) );
  XNOR2_X1 U8482 ( .A(n8650), .B(n7248), .ZN(n10470) );
  NOR2_X1 U8483 ( .A1(n4856), .A2(n7249), .ZN(n10169) );
  INV_X1 U8484 ( .A(n10169), .ZN(n8282) );
  AOI22_X1 U8485 ( .A1(n10120), .A2(n6712), .B1(n10146), .B2(n6914), .ZN(n7255) );
  OAI21_X1 U8486 ( .B1(n7252), .B2(n7251), .A(n7250), .ZN(n7253) );
  NAND2_X1 U8487 ( .A1(n7253), .A2(n10152), .ZN(n7254) );
  OAI211_X1 U8488 ( .C1(n10470), .C2(n6896), .A(n7255), .B(n7254), .ZN(n10473)
         );
  OAI211_X1 U8489 ( .C1(n10472), .C2(n7257), .A(n10250), .B(n7256), .ZN(n10471) );
  OAI22_X1 U8490 ( .A1(n10471), .A2(n10095), .B1(n5335), .B2(n10160), .ZN(
        n7258) );
  OAI21_X1 U8491 ( .B1(n10473), .B2(n7258), .A(n10163), .ZN(n7260) );
  AOI22_X1 U8492 ( .A1(n10165), .A2(n8776), .B1(n4856), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7259) );
  OAI211_X1 U8493 ( .C1(n10470), .C2(n8282), .A(n7260), .B(n7259), .ZN(
        P1_U3290) );
  OAI21_X1 U8494 ( .B1(n7262), .B2(n8651), .A(n7261), .ZN(n10489) );
  INV_X1 U8495 ( .A(n10489), .ZN(n7278) );
  AOI22_X1 U8496 ( .A1(n10120), .A2(n6914), .B1(n10146), .B2(n9900), .ZN(n7268) );
  OAI21_X1 U8497 ( .B1(n7265), .B2(n7264), .A(n7263), .ZN(n7266) );
  NAND2_X1 U8498 ( .A1(n7266), .A2(n10152), .ZN(n7267) );
  OAI211_X1 U8499 ( .C1(n7278), .C2(n6896), .A(n7268), .B(n7267), .ZN(n10487)
         );
  NAND2_X1 U8500 ( .A1(n10487), .A2(n10163), .ZN(n7277) );
  INV_X1 U8501 ( .A(n10137), .ZN(n10167) );
  OR2_X1 U8502 ( .A1(n7269), .A2(n10485), .ZN(n7270) );
  NAND2_X1 U8503 ( .A1(n7271), .A2(n7270), .ZN(n10486) );
  INV_X1 U8504 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7272) );
  AOI22_X1 U8505 ( .A1(n4856), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10128), .B2(
        n7272), .ZN(n7273) );
  OAI21_X1 U8506 ( .B1(n10167), .B2(n10486), .A(n7273), .ZN(n7274) );
  AOI21_X1 U8507 ( .B1(n10165), .B2(n7275), .A(n7274), .ZN(n7276) );
  OAI211_X1 U8508 ( .C1(n7278), .C2(n8282), .A(n7277), .B(n7276), .ZN(P1_U3288) );
  NAND2_X1 U8509 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8956) );
  INV_X1 U8510 ( .A(n8956), .ZN(n7282) );
  AOI211_X1 U8511 ( .C1(n7280), .C2(n7279), .A(n7291), .B(n10427), .ZN(n7281)
         );
  AOI211_X1 U8512 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n10448), .A(n7282), .B(
        n7281), .ZN(n7287) );
  OAI211_X1 U8513 ( .C1(n7285), .C2(n7284), .A(n10425), .B(n7283), .ZN(n7286)
         );
  OAI211_X1 U8514 ( .C1(n10426), .C2(n7288), .A(n7287), .B(n7286), .ZN(
        P2_U3251) );
  NOR2_X1 U8515 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6144), .ZN(n7295) );
  INV_X1 U8516 ( .A(n7304), .ZN(n7293) );
  NOR3_X1 U8517 ( .A1(n7291), .A2(n7290), .A3(n7289), .ZN(n7292) );
  NOR3_X1 U8518 ( .A1(n7293), .A2(n7292), .A3(n10427), .ZN(n7294) );
  AOI211_X1 U8519 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n10448), .A(n7295), .B(
        n7294), .ZN(n7300) );
  OAI211_X1 U8520 ( .C1(n7298), .C2(n7297), .A(n10425), .B(n7296), .ZN(n7299)
         );
  OAI211_X1 U8521 ( .C1(n10426), .C2(n7301), .A(n7300), .B(n7299), .ZN(
        P2_U3252) );
  INV_X1 U8522 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9157) );
  NOR2_X1 U8523 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9157), .ZN(n7307) );
  AND3_X1 U8524 ( .A1(n7304), .A2(n7303), .A3(n7302), .ZN(n7305) );
  NOR3_X1 U8525 ( .A1(n9390), .A2(n7305), .A3(n10427), .ZN(n7306) );
  AOI211_X1 U8526 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10448), .A(n7307), .B(
        n7306), .ZN(n7312) );
  OAI211_X1 U8527 ( .C1(n7310), .C2(n7309), .A(n10425), .B(n7308), .ZN(n7311)
         );
  OAI211_X1 U8528 ( .C1(n10426), .C2(n7313), .A(n7312), .B(n7311), .ZN(
        P2_U3253) );
  NAND2_X1 U8529 ( .A1(n7314), .A2(n10137), .ZN(n7317) );
  AOI22_X1 U8530 ( .A1(n4856), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n10128), .B2(
        n7315), .ZN(n7316) );
  OAI211_X1 U8531 ( .C1(n7318), .C2(n10130), .A(n7317), .B(n7316), .ZN(n7319)
         );
  AOI21_X1 U8532 ( .B1(n7320), .B2(n10169), .A(n7319), .ZN(n7321) );
  OAI21_X1 U8533 ( .B1(n7322), .B2(n4856), .A(n7321), .ZN(P1_U3287) );
  AOI22_X1 U8534 ( .A1(n4856), .A2(P1_REG2_REG_2__SCAN_IN), .B1(n10128), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7325) );
  NAND2_X1 U8535 ( .A1(n10137), .A2(n7323), .ZN(n7324) );
  OAI211_X1 U8536 ( .C1(n7326), .C2(n10130), .A(n7325), .B(n7324), .ZN(n7327)
         );
  AOI21_X1 U8537 ( .B1(n10169), .B2(n7328), .A(n7327), .ZN(n7329) );
  OAI21_X1 U8538 ( .B1(n7330), .B2(n4856), .A(n7329), .ZN(P1_U3289) );
  INV_X1 U8539 ( .A(n7331), .ZN(n8314) );
  OAI222_X1 U8540 ( .A1(n9944), .A2(P1_U3084), .B1(n9064), .B2(n8314), .C1(
        n9060), .C2(n5699), .ZN(P1_U3334) );
  OR2_X1 U8541 ( .A1(n7333), .A2(n7332), .ZN(n7334) );
  NAND2_X1 U8542 ( .A1(n9042), .A2(n9899), .ZN(n7336) );
  OAI21_X1 U8543 ( .B1(n7337), .B2(n7514), .A(n7336), .ZN(n7338) );
  XNOR2_X1 U8544 ( .A(n8946), .B(n7338), .ZN(n7341) );
  NAND2_X1 U8545 ( .A1(n9046), .A2(n9899), .ZN(n7340) );
  NAND2_X1 U8546 ( .A1(n9042), .A2(n10514), .ZN(n7339) );
  NAND2_X1 U8547 ( .A1(n7340), .A2(n7339), .ZN(n7346) );
  NAND2_X1 U8548 ( .A1(n7342), .A2(n7341), .ZN(n7344) );
  INV_X1 U8549 ( .A(n7513), .ZN(n7349) );
  INV_X1 U8550 ( .A(n7343), .ZN(n7345) );
  NAND2_X1 U8551 ( .A1(n7345), .A2(n7344), .ZN(n7347) );
  AOI22_X1 U8552 ( .A1(n7349), .A2(n7348), .B1(n7347), .B2(n7346), .ZN(n7356)
         );
  NAND2_X1 U8553 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10419) );
  INV_X1 U8554 ( .A(n10419), .ZN(n7350) );
  AOI21_X1 U8555 ( .B1(n9853), .B2(n9898), .A(n7350), .ZN(n7352) );
  NAND2_X1 U8556 ( .A1(n9873), .A2(n9900), .ZN(n7351) );
  OAI211_X1 U8557 ( .C1(n9876), .C2(n7353), .A(n7352), .B(n7351), .ZN(n7354)
         );
  AOI21_X1 U8558 ( .B1(n10514), .B2(n9863), .A(n7354), .ZN(n7355) );
  OAI21_X1 U8559 ( .B1(n7356), .B2(n9879), .A(n7355), .ZN(P1_U3225) );
  AOI21_X1 U8560 ( .B1(n7358), .B2(n6233), .A(n7357), .ZN(n7360) );
  AOI22_X1 U8561 ( .A1(n7855), .A2(n6278), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7845), .ZN(n7359) );
  NOR2_X1 U8562 ( .A1(n7360), .A2(n7359), .ZN(n7844) );
  AOI21_X1 U8563 ( .B1(n7360), .B2(n7359), .A(n7844), .ZN(n7370) );
  AOI22_X1 U8564 ( .A1(n7855), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7977), .B2(
        n7845), .ZN(n7364) );
  OAI21_X1 U8565 ( .B1(n7362), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7361), .ZN(
        n7363) );
  NAND2_X1 U8566 ( .A1(n7364), .A2(n7363), .ZN(n7854) );
  OAI21_X1 U8567 ( .B1(n7364), .B2(n7363), .A(n7854), .ZN(n7368) );
  INV_X1 U8568 ( .A(n10448), .ZN(n8001) );
  INV_X1 U8569 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7366) );
  NAND2_X1 U8570 ( .A1(n10455), .A2(n7855), .ZN(n7365) );
  NAND2_X1 U8571 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8985) );
  OAI211_X1 U8572 ( .C1(n8001), .C2(n7366), .A(n7365), .B(n8985), .ZN(n7367)
         );
  AOI21_X1 U8573 ( .B1(n7368), .B2(n10425), .A(n7367), .ZN(n7369) );
  OAI21_X1 U8574 ( .B1(n7370), .B2(n10427), .A(n7369), .ZN(P2_U3259) );
  INV_X1 U8575 ( .A(n7371), .ZN(n10564) );
  NOR3_X1 U8576 ( .A1(n7372), .A2(n10538), .A3(n9129), .ZN(n7373) );
  AOI21_X1 U8577 ( .B1(n10564), .B2(n10561), .A(n7373), .ZN(n7381) );
  NOR2_X1 U8578 ( .A1(n7374), .A2(n10615), .ZN(n7379) );
  AND2_X1 U8579 ( .A1(n10588), .A2(n10621), .ZN(n7378) );
  NOR2_X1 U8580 ( .A1(n10623), .A2(n7596), .ZN(n7377) );
  INV_X1 U8581 ( .A(n10538), .ZN(n9374) );
  NAND2_X1 U8582 ( .A1(n10609), .A2(n9374), .ZN(n7375) );
  NAND2_X1 U8583 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n9380) );
  OAI211_X1 U8584 ( .C1(n7590), .C2(n10611), .A(n7375), .B(n9380), .ZN(n7376)
         );
  NOR4_X1 U8585 ( .A1(n7379), .A2(n7378), .A3(n7377), .A4(n7376), .ZN(n7380)
         );
  OAI21_X1 U8586 ( .B1(n7382), .B2(n7381), .A(n7380), .ZN(P2_U3233) );
  NAND2_X1 U8587 ( .A1(n9046), .A2(n9898), .ZN(n7384) );
  NAND2_X1 U8588 ( .A1(n7424), .A2(n9042), .ZN(n7383) );
  NAND2_X1 U8589 ( .A1(n7384), .A2(n7383), .ZN(n7511) );
  NAND2_X1 U8590 ( .A1(n7424), .A2(n4862), .ZN(n7387) );
  NAND2_X1 U8591 ( .A1(n9042), .A2(n9898), .ZN(n7386) );
  NAND2_X1 U8592 ( .A1(n7387), .A2(n7386), .ZN(n7388) );
  XOR2_X1 U8593 ( .A(n7511), .B(n7512), .Z(n7389) );
  XNOR2_X1 U8594 ( .A(n7513), .B(n7389), .ZN(n7395) );
  INV_X1 U8595 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7390) );
  NOR2_X1 U8596 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7390), .ZN(n10380) );
  AOI21_X1 U8597 ( .B1(n9853), .B2(n9897), .A(n10380), .ZN(n7392) );
  NAND2_X1 U8598 ( .A1(n9873), .A2(n9899), .ZN(n7391) );
  OAI211_X1 U8599 ( .C1(n9876), .C2(n7442), .A(n7392), .B(n7391), .ZN(n7393)
         );
  AOI21_X1 U8600 ( .B1(n7424), .B2(n9863), .A(n7393), .ZN(n7394) );
  OAI21_X1 U8601 ( .B1(n7395), .B2(n9879), .A(n7394), .ZN(P1_U3237) );
  NAND2_X1 U8602 ( .A1(n7412), .A2(n7396), .ZN(n7397) );
  NAND2_X1 U8603 ( .A1(n7397), .A2(n8658), .ZN(n7750) );
  OAI21_X1 U8604 ( .B1(n7397), .B2(n8658), .A(n7750), .ZN(n7398) );
  INV_X1 U8605 ( .A(n7398), .ZN(n7470) );
  OAI21_X1 U8606 ( .B1(n7401), .B2(n7400), .A(n7399), .ZN(n7402) );
  AOI222_X1 U8607 ( .A1(n10152), .A2(n7402), .B1(n9898), .B2(n10120), .C1(
        n9896), .C2(n10146), .ZN(n7469) );
  MUX2_X1 U8608 ( .A(n7403), .B(n7469), .S(n10163), .Z(n7409) );
  INV_X1 U8609 ( .A(n7422), .ZN(n7405) );
  INV_X1 U8610 ( .A(n7756), .ZN(n7404) );
  AOI211_X1 U8611 ( .C1(n7523), .C2(n7405), .A(n10633), .B(n7404), .ZN(n7467)
         );
  OAI22_X1 U8612 ( .A1(n10130), .A2(n7406), .B1(n7521), .B2(n10160), .ZN(n7407) );
  AOI21_X1 U8613 ( .B1(n7467), .B2(n10117), .A(n7407), .ZN(n7408) );
  OAI211_X1 U8614 ( .C1(n10134), .C2(n7470), .A(n7409), .B(n7408), .ZN(
        P1_U3284) );
  INV_X1 U8615 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7427) );
  NAND2_X1 U8616 ( .A1(n7410), .A2(n8655), .ZN(n7411) );
  NAND2_X1 U8617 ( .A1(n7412), .A2(n7411), .ZN(n7416) );
  INV_X1 U8618 ( .A(n7416), .ZN(n7448) );
  OAI22_X1 U8619 ( .A1(n7414), .A2(n10149), .B1(n10111), .B2(n7413), .ZN(n7415) );
  AOI21_X1 U8620 ( .B1(n7416), .B2(n10604), .A(n7415), .ZN(n7420) );
  INV_X1 U8621 ( .A(n8788), .ZN(n7417) );
  AOI21_X1 U8622 ( .B1(n7102), .B2(n8714), .A(n7417), .ZN(n8550) );
  XNOR2_X1 U8623 ( .A(n8550), .B(n5918), .ZN(n7418) );
  NAND2_X1 U8624 ( .A1(n7418), .A2(n10152), .ZN(n7419) );
  AND2_X1 U8625 ( .A1(n7420), .A2(n7419), .ZN(n7441) );
  INV_X1 U8626 ( .A(n7421), .ZN(n7423) );
  AOI21_X1 U8627 ( .B1(n7424), .B2(n7423), .A(n7422), .ZN(n7445) );
  AOI22_X1 U8628 ( .A1(n7445), .A2(n10250), .B1(n10597), .B2(n7424), .ZN(n7425) );
  OAI211_X1 U8629 ( .C1(n7448), .C2(n10600), .A(n7441), .B(n7425), .ZN(n7428)
         );
  NAND2_X1 U8630 ( .A1(n7428), .A2(n4855), .ZN(n7426) );
  OAI21_X1 U8631 ( .B1(n4855), .B2(n7427), .A(n7426), .ZN(P1_U3472) );
  NAND2_X1 U8632 ( .A1(n7428), .A2(n10656), .ZN(n7429) );
  OAI21_X1 U8633 ( .B1(n10656), .B2(n6669), .A(n7429), .ZN(P1_U3529) );
  XNOR2_X1 U8634 ( .A(n7731), .B(n7430), .ZN(n7433) );
  AOI21_X1 U8635 ( .B1(n7436), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7431), .ZN(
        n7432) );
  NAND2_X1 U8636 ( .A1(n7433), .A2(n7432), .ZN(n7730) );
  OAI21_X1 U8637 ( .B1(n7433), .B2(n7432), .A(n7730), .ZN(n7434) );
  AOI22_X1 U8638 ( .A1(n10407), .A2(P1_ADDR_REG_14__SCAN_IN), .B1(n10398), 
        .B2(n7434), .ZN(n7440) );
  XNOR2_X1 U8639 ( .A(n7731), .B(n7722), .ZN(n7724) );
  OAI21_X1 U8640 ( .B1(n7436), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7435), .ZN(
        n7723) );
  XNOR2_X1 U8641 ( .A(n7724), .B(n7723), .ZN(n7438) );
  NOR2_X1 U8642 ( .A1(n7437), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9751) );
  AOI21_X1 U8643 ( .B1(n10414), .B2(n7438), .A(n9751), .ZN(n7439) );
  OAI211_X1 U8644 ( .C1(n7721), .C2(n9943), .A(n7440), .B(n7439), .ZN(P1_U3255) );
  MUX2_X1 U8645 ( .A(n7441), .B(n6656), .S(n4856), .Z(n7447) );
  OAI22_X1 U8646 ( .A1(n10130), .A2(n7443), .B1(n7442), .B2(n10160), .ZN(n7444) );
  AOI21_X1 U8647 ( .B1(n7445), .B2(n10137), .A(n7444), .ZN(n7446) );
  OAI211_X1 U8648 ( .C1(n7448), .C2(n8282), .A(n7447), .B(n7446), .ZN(P1_U3285) );
  INV_X1 U8649 ( .A(n7449), .ZN(n7450) );
  AND2_X1 U8650 ( .A1(n7451), .A2(n7450), .ZN(n7452) );
  NAND2_X1 U8651 ( .A1(n7453), .A2(n7452), .ZN(n7459) );
  INV_X1 U8652 ( .A(n7454), .ZN(n7455) );
  NAND2_X1 U8653 ( .A1(n7459), .A2(n9592), .ZN(n9517) );
  INV_X2 U8654 ( .A(n9517), .ZN(n9618) );
  NAND2_X1 U8655 ( .A1(n7527), .A2(n8343), .ZN(n7535) );
  OR2_X1 U8656 ( .A1(n9618), .A2(n7535), .ZN(n7601) );
  INV_X1 U8657 ( .A(n7601), .ZN(n7634) );
  AND2_X1 U8658 ( .A1(n8524), .A2(n10467), .ZN(n7456) );
  NAND2_X1 U8659 ( .A1(n9457), .A2(n7456), .ZN(n9620) );
  INV_X1 U8660 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7457) );
  OAI22_X1 U8661 ( .A1(n9457), .A2(n7457), .B1(n9592), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n7458) );
  INV_X1 U8662 ( .A(n7458), .ZN(n7462) );
  OR2_X1 U8663 ( .A1(n7459), .A2(n8527), .ZN(n9451) );
  INV_X1 U8664 ( .A(n9451), .ZN(n9632) );
  NAND2_X1 U8665 ( .A1(n9632), .A2(n7460), .ZN(n7461) );
  OAI211_X1 U8666 ( .C1(n10502), .C2(n9620), .A(n7462), .B(n7461), .ZN(n7463)
         );
  AOI21_X1 U8667 ( .B1(n7634), .B2(n7464), .A(n7463), .ZN(n7465) );
  OAI21_X1 U8668 ( .B1(n7466), .B2(n9618), .A(n7465), .ZN(P2_U3293) );
  INV_X1 U8669 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7472) );
  AOI21_X1 U8670 ( .B1(n10597), .B2(n7523), .A(n7467), .ZN(n7468) );
  OAI211_X1 U8671 ( .C1(n10580), .C2(n7470), .A(n7469), .B(n7468), .ZN(n7483)
         );
  NAND2_X1 U8672 ( .A1(n7483), .A2(n4855), .ZN(n7471) );
  OAI21_X1 U8673 ( .B1(n4855), .B2(n7472), .A(n7471), .ZN(P1_U3475) );
  INV_X1 U8674 ( .A(n10536), .ZN(n8394) );
  OAI21_X1 U8675 ( .B1(n10611), .B2(n8394), .A(n7473), .ZN(n7474) );
  AOI21_X1 U8676 ( .B1(n10609), .B2(n9377), .A(n7474), .ZN(n7475) );
  OAI21_X1 U8677 ( .B1(n7612), .B2(n10623), .A(n7475), .ZN(n7481) );
  INV_X1 U8678 ( .A(n9129), .ZN(n10560) );
  AOI22_X1 U8679 ( .A1(n10560), .A2(n9377), .B1(n10561), .B2(n7476), .ZN(n7477) );
  NOR3_X1 U8680 ( .A1(n7479), .A2(n7478), .A3(n7477), .ZN(n7480) );
  AOI211_X1 U8681 ( .C1(n10621), .C2(n7566), .A(n7481), .B(n7480), .ZN(n7482)
         );
  OAI21_X1 U8682 ( .B1(n8964), .B2(n10615), .A(n7482), .ZN(P2_U3229) );
  NAND2_X1 U8683 ( .A1(n7483), .A2(n10656), .ZN(n7484) );
  OAI21_X1 U8684 ( .B1(n10656), .B2(n5477), .A(n7484), .ZN(P1_U3530) );
  INV_X1 U8685 ( .A(n7485), .ZN(n7528) );
  OAI222_X1 U8686 ( .A1(n7486), .A2(P1_U3084), .B1(n10286), .B2(n5725), .C1(
        n7528), .C2(n9064), .ZN(P1_U3333) );
  INV_X1 U8687 ( .A(n7487), .ZN(n7510) );
  OAI222_X1 U8688 ( .A1(n8538), .A2(n7510), .B1(P2_U3152), .B2(n8522), .C1(
        n7488), .C2(n4858), .ZN(P2_U3337) );
  OAI21_X1 U8689 ( .B1(n8664), .B2(n7490), .A(n7489), .ZN(n7491) );
  AOI222_X1 U8690 ( .A1(n10152), .A2(n7491), .B1(n9893), .B2(n10146), .C1(
        n9895), .C2(n10120), .ZN(n10599) );
  AOI211_X1 U8691 ( .C1(n10596), .C2(n8044), .A(n10633), .B(n7640), .ZN(n10595) );
  INV_X1 U8692 ( .A(n10596), .ZN(n7492) );
  NOR2_X1 U8693 ( .A1(n7492), .A2(n10130), .ZN(n7495) );
  OAI22_X1 U8694 ( .A1(n10163), .A2(n7493), .B1(n8033), .B2(n10160), .ZN(n7494) );
  AOI211_X1 U8695 ( .C1(n10595), .C2(n10117), .A(n7495), .B(n7494), .ZN(n7498)
         );
  XNOR2_X1 U8696 ( .A(n7496), .B(n8664), .ZN(n10601) );
  INV_X1 U8697 ( .A(n10601), .ZN(n10603) );
  INV_X1 U8698 ( .A(n10134), .ZN(n10050) );
  NAND2_X1 U8699 ( .A1(n10603), .A2(n10050), .ZN(n7497) );
  OAI211_X1 U8700 ( .C1(n10599), .C2(n4856), .A(n7498), .B(n7497), .ZN(
        P1_U3281) );
  INV_X1 U8701 ( .A(n7908), .ZN(n10642) );
  INV_X1 U8702 ( .A(n7501), .ZN(n7499) );
  AOI21_X1 U8703 ( .B1(n10613), .B2(n7499), .A(n10615), .ZN(n7504) );
  NOR3_X1 U8704 ( .A1(n7500), .A2(n7590), .A3(n9129), .ZN(n7503) );
  NAND2_X1 U8705 ( .A1(n7502), .A2(n7501), .ZN(n7772) );
  OAI21_X1 U8706 ( .B1(n7504), .B2(n7503), .A(n7772), .ZN(n7508) );
  INV_X1 U8707 ( .A(n8976), .ZN(n9371) );
  NOR2_X1 U8708 ( .A1(n10623), .A2(n7710), .ZN(n7506) );
  INV_X1 U8709 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9400) );
  OAI22_X1 U8710 ( .A1(n10500), .A2(n7590), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9400), .ZN(n7505) );
  AOI211_X1 U8711 ( .C1(n8984), .C2(n9371), .A(n7506), .B(n7505), .ZN(n7507)
         );
  OAI211_X1 U8712 ( .C1(n10642), .C2(n6546), .A(n7508), .B(n7507), .ZN(
        P2_U3238) );
  OAI222_X1 U8713 ( .A1(P1_U3084), .A2(n8762), .B1(n9064), .B2(n7510), .C1(
        n7509), .C2(n10286), .ZN(P1_U3332) );
  NAND2_X1 U8714 ( .A1(n7523), .A2(n8234), .ZN(n7516) );
  NAND2_X1 U8715 ( .A1(n9042), .A2(n9897), .ZN(n7515) );
  NAND2_X1 U8716 ( .A1(n7516), .A2(n7515), .ZN(n7517) );
  INV_X4 U8717 ( .A(n8946), .ZN(n9017) );
  XNOR2_X1 U8718 ( .A(n7517), .B(n9017), .ZN(n7785) );
  AOI22_X1 U8719 ( .A1(n7523), .A2(n9042), .B1(n9046), .B2(n9897), .ZN(n7784)
         );
  XNOR2_X1 U8720 ( .A(n7785), .B(n7784), .ZN(n7803) );
  XOR2_X1 U8721 ( .A(n7802), .B(n7803), .Z(n7525) );
  AOI21_X1 U8722 ( .B1(n9853), .B2(n9896), .A(n7518), .ZN(n7520) );
  NAND2_X1 U8723 ( .A1(n9873), .A2(n9898), .ZN(n7519) );
  OAI211_X1 U8724 ( .C1(n9876), .C2(n7521), .A(n7520), .B(n7519), .ZN(n7522)
         );
  AOI21_X1 U8725 ( .B1(n7523), .B2(n9863), .A(n7522), .ZN(n7524) );
  OAI21_X1 U8726 ( .B1(n7525), .B2(n9879), .A(n7524), .ZN(P1_U3211) );
  OAI222_X1 U8727 ( .A1(n8538), .A2(n7528), .B1(P2_U3152), .B2(n7527), .C1(
        n7526), .C2(n4858), .ZN(P2_U3338) );
  NAND2_X1 U8728 ( .A1(n6870), .A2(n7529), .ZN(n8365) );
  AND2_X1 U8729 ( .A1(n7530), .A2(n8365), .ZN(n10463) );
  OR2_X1 U8730 ( .A1(n10463), .A2(n9594), .ZN(n7532) );
  NAND2_X1 U8731 ( .A1(n9379), .A2(n9626), .ZN(n7531) );
  AND2_X1 U8732 ( .A1(n7532), .A2(n7531), .ZN(n10464) );
  OAI21_X1 U8733 ( .B1(n7533), .B2(n9592), .A(n10464), .ZN(n7539) );
  INV_X1 U8734 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7534) );
  NOR2_X1 U8735 ( .A1(n9457), .A2(n7534), .ZN(n7538) );
  NAND2_X1 U8736 ( .A1(n7617), .A2(n7535), .ZN(n7536) );
  NAND2_X1 U8737 ( .A1(n9457), .A2(n7536), .ZN(n9634) );
  NOR2_X1 U8738 ( .A1(n9634), .A2(n10463), .ZN(n7537) );
  AOI211_X1 U8739 ( .C1(n9457), .C2(n7539), .A(n7538), .B(n7537), .ZN(n7541)
         );
  OAI21_X1 U8740 ( .B1(n9606), .B2(n9632), .A(n10468), .ZN(n7540) );
  NAND2_X1 U8741 ( .A1(n7541), .A2(n7540), .ZN(P2_U3296) );
  OAI22_X1 U8742 ( .A1(n7542), .A2(n9634), .B1(n7055), .B2(n9457), .ZN(n7544)
         );
  NOR2_X1 U8743 ( .A1(n9592), .A2(n9332), .ZN(n7543) );
  AOI211_X1 U8744 ( .C1(n9632), .C2(n7545), .A(n7544), .B(n7543), .ZN(n7548)
         );
  NAND2_X1 U8745 ( .A1(n9606), .A2(n7546), .ZN(n7547) );
  OAI211_X1 U8746 ( .C1(n7549), .C2(n9618), .A(n7548), .B(n7547), .ZN(P2_U3295) );
  NAND2_X1 U8747 ( .A1(n7550), .A2(n8378), .ZN(n7688) );
  INV_X1 U8748 ( .A(n7688), .ZN(n7552) );
  NAND2_X1 U8749 ( .A1(n9377), .A2(n10507), .ZN(n7553) );
  INV_X1 U8750 ( .A(n8497), .ZN(n8386) );
  NAND2_X1 U8751 ( .A1(n9375), .A2(n7566), .ZN(n7554) );
  OR2_X1 U8752 ( .A1(n10527), .A2(n8394), .ZN(n7555) );
  NAND2_X1 U8753 ( .A1(n10527), .A2(n8394), .ZN(n7556) );
  NAND2_X1 U8754 ( .A1(n10544), .A2(n7656), .ZN(n8401) );
  OR2_X1 U8755 ( .A1(n10544), .A2(n7656), .ZN(n8400) );
  OR2_X1 U8756 ( .A1(n10555), .A2(n10538), .ZN(n8404) );
  NAND2_X1 U8757 ( .A1(n10555), .A2(n10538), .ZN(n8405) );
  AND2_X2 U8758 ( .A1(n8404), .A2(n8405), .ZN(n8502) );
  NAND2_X1 U8759 ( .A1(n10588), .A2(n10557), .ZN(n8417) );
  NAND2_X1 U8760 ( .A1(n8407), .A2(n8417), .ZN(n8504) );
  INV_X1 U8761 ( .A(n8405), .ZN(n7591) );
  NAND2_X1 U8762 ( .A1(n7560), .A2(n8407), .ZN(n7558) );
  OR2_X1 U8763 ( .A1(n10620), .A2(n7590), .ZN(n8413) );
  NAND2_X1 U8764 ( .A1(n10620), .A2(n7590), .ZN(n8415) );
  NAND2_X1 U8765 ( .A1(n8413), .A2(n8415), .ZN(n8505) );
  NAND2_X1 U8766 ( .A1(n7558), .A2(n8505), .ZN(n7561) );
  INV_X1 U8767 ( .A(n8407), .ZN(n8410) );
  NOR2_X1 U8768 ( .A1(n8505), .A2(n8410), .ZN(n7559) );
  AOI21_X1 U8769 ( .B1(n7561), .B2(n7705), .A(n9594), .ZN(n7563) );
  OAI22_X1 U8770 ( .A1(n10612), .A2(n9599), .B1(n10557), .B2(n9597), .ZN(n7562) );
  OR2_X1 U8771 ( .A1(n7563), .A2(n7562), .ZN(n10628) );
  INV_X1 U8772 ( .A(n10628), .ZN(n7585) );
  NAND2_X1 U8773 ( .A1(n7691), .A2(n10502), .ZN(n7564) );
  NAND2_X1 U8774 ( .A1(n7565), .A2(n7564), .ZN(n7695) );
  NAND2_X1 U8775 ( .A1(n7695), .A2(n8495), .ZN(n7603) );
  NAND2_X1 U8776 ( .A1(n10501), .A2(n10507), .ZN(n7604) );
  INV_X1 U8777 ( .A(n7566), .ZN(n10522) );
  NAND2_X1 U8778 ( .A1(n10522), .A2(n9375), .ZN(n7567) );
  NAND2_X1 U8779 ( .A1(n7603), .A2(n4892), .ZN(n7572) );
  INV_X1 U8780 ( .A(n7567), .ZN(n7568) );
  NAND2_X1 U8781 ( .A1(n7570), .A2(n7569), .ZN(n7571) );
  NAND2_X1 U8782 ( .A1(n10527), .A2(n10536), .ZN(n8393) );
  INV_X1 U8783 ( .A(n7678), .ZN(n7574) );
  AND2_X1 U8784 ( .A1(n8400), .A2(n8401), .ZN(n8501) );
  NAND2_X1 U8785 ( .A1(n7574), .A2(n7573), .ZN(n7669) );
  INV_X1 U8786 ( .A(n8502), .ZN(n7575) );
  OR2_X1 U8787 ( .A1(n10544), .A2(n10558), .ZN(n7670) );
  AND2_X1 U8788 ( .A1(n7575), .A2(n7670), .ZN(n7576) );
  NAND2_X1 U8789 ( .A1(n10555), .A2(n9374), .ZN(n7587) );
  OR2_X1 U8790 ( .A1(n10588), .A2(n10608), .ZN(n7577) );
  NOR2_X1 U8791 ( .A1(n7578), .A2(n8505), .ZN(n10625) );
  INV_X1 U8792 ( .A(n10625), .ZN(n7579) );
  INV_X1 U8793 ( .A(n9634), .ZN(n9605) );
  NAND3_X1 U8794 ( .A1(n7579), .A2(n9605), .A3(n7716), .ZN(n7584) );
  OAI22_X1 U8795 ( .A1(n9457), .A2(n7134), .B1(n10624), .B2(n9592), .ZN(n7582)
         );
  INV_X1 U8796 ( .A(n10620), .ZN(n10626) );
  INV_X1 U8797 ( .A(n10507), .ZN(n8382) );
  INV_X1 U8798 ( .A(n10527), .ZN(n8395) );
  INV_X1 U8799 ( .A(n10544), .ZN(n10547) );
  INV_X1 U8800 ( .A(n7711), .ZN(n7580) );
  OAI21_X1 U8801 ( .B1(n10626), .B2(n4920), .A(n7580), .ZN(n10627) );
  NOR2_X1 U8802 ( .A1(n10627), .A2(n9451), .ZN(n7581) );
  AOI211_X1 U8803 ( .C1(n9606), .C2(n10620), .A(n7582), .B(n7581), .ZN(n7583)
         );
  OAI211_X1 U8804 ( .C1(n9618), .C2(n7585), .A(n7584), .B(n7583), .ZN(P2_U3286) );
  AND2_X1 U8805 ( .A1(n7586), .A2(n7587), .ZN(n7589) );
  OAI21_X1 U8806 ( .B1(n7589), .B2(n8504), .A(n7588), .ZN(n10592) );
  INV_X1 U8807 ( .A(n10592), .ZN(n7602) );
  INV_X1 U8808 ( .A(n7590), .ZN(n9372) );
  AOI22_X1 U8809 ( .A1(n9624), .A2(n9374), .B1(n9372), .B2(n9626), .ZN(n7595)
         );
  INV_X1 U8810 ( .A(n7662), .ZN(n7592) );
  OAI21_X1 U8811 ( .B1(n7592), .B2(n7591), .A(n8504), .ZN(n7593) );
  NAND3_X1 U8812 ( .A1(n7593), .A2(n9629), .A3(n7560), .ZN(n7594) );
  OAI211_X1 U8813 ( .C1(n7602), .C2(n7617), .A(n7595), .B(n7594), .ZN(n10590)
         );
  NAND2_X1 U8814 ( .A1(n10590), .A2(n9517), .ZN(n7600) );
  OAI22_X1 U8815 ( .A1(n9457), .A2(n7133), .B1(n7596), .B2(n9592), .ZN(n7598)
         );
  XNOR2_X1 U8816 ( .A(n7664), .B(n10588), .ZN(n10589) );
  NOR2_X1 U8817 ( .A1(n10589), .A2(n9451), .ZN(n7597) );
  AOI211_X1 U8818 ( .C1(n9606), .C2(n10588), .A(n7598), .B(n7597), .ZN(n7599)
         );
  OAI211_X1 U8819 ( .C1(n7602), .C2(n7601), .A(n7600), .B(n7599), .ZN(P2_U3287) );
  NAND2_X1 U8820 ( .A1(n7603), .A2(n7604), .ZN(n7605) );
  XNOR2_X1 U8821 ( .A(n7605), .B(n8497), .ZN(n10520) );
  INV_X1 U8822 ( .A(n10520), .ZN(n7616) );
  OAI21_X1 U8823 ( .B1(n4921), .B2(n8386), .A(n7606), .ZN(n7607) );
  NAND2_X1 U8824 ( .A1(n7607), .A2(n9629), .ZN(n7609) );
  AOI22_X1 U8825 ( .A1(n9624), .A2(n9377), .B1(n10536), .B2(n9626), .ZN(n7608)
         );
  NAND2_X1 U8826 ( .A1(n7609), .A2(n7608), .ZN(n10525) );
  NAND2_X1 U8827 ( .A1(n7697), .A2(n7566), .ZN(n7610) );
  NAND2_X1 U8828 ( .A1(n7610), .A2(n10528), .ZN(n7611) );
  OR2_X1 U8829 ( .A1(n7611), .A2(n7648), .ZN(n10521) );
  OAI22_X1 U8830 ( .A1(n10521), .A2(n8339), .B1(n9592), .B2(n7612), .ZN(n7613)
         );
  OAI21_X1 U8831 ( .B1(n10525), .B2(n7613), .A(n9457), .ZN(n7615) );
  AOI22_X1 U8832 ( .A1(n9606), .A2(n7566), .B1(P2_REG2_REG_5__SCAN_IN), .B2(
        n9618), .ZN(n7614) );
  OAI211_X1 U8833 ( .C1(n9634), .C2(n7616), .A(n7615), .B(n7614), .ZN(P2_U3291) );
  INV_X1 U8834 ( .A(n7617), .ZN(n7626) );
  OAI22_X1 U8835 ( .A1(n7620), .A2(n9597), .B1(n7691), .B2(n9599), .ZN(n7625)
         );
  AOI21_X1 U8836 ( .B1(n7623), .B2(n7622), .A(n9594), .ZN(n7624) );
  AOI211_X1 U8837 ( .C1(n7626), .C2(n10483), .A(n7625), .B(n7624), .ZN(n10480)
         );
  INV_X1 U8838 ( .A(n7627), .ZN(n7630) );
  NAND2_X1 U8839 ( .A1(n7628), .A2(n7633), .ZN(n7629) );
  NAND2_X1 U8840 ( .A1(n7630), .A2(n7629), .ZN(n10479) );
  OAI22_X1 U8841 ( .A1(n9451), .A2(n10479), .B1(n7631), .B2(n9592), .ZN(n7632)
         );
  AOI21_X1 U8842 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n9618), .A(n7632), .ZN(
        n7636) );
  AOI22_X1 U8843 ( .A1(n7634), .A2(n10483), .B1(n9606), .B2(n7633), .ZN(n7635)
         );
  OAI211_X1 U8844 ( .C1(n10480), .C2(n9618), .A(n7636), .B(n7635), .ZN(
        P2_U3294) );
  XNOR2_X1 U8845 ( .A(n7637), .B(n4980), .ZN(n7638) );
  OAI222_X1 U8846 ( .A1(n10111), .A2(n8201), .B1(n10149), .B2(n8041), .C1(
        n7638), .C2(n10107), .ZN(n10635) );
  INV_X1 U8847 ( .A(n10635), .ZN(n7647) );
  XNOR2_X1 U8848 ( .A(n7639), .B(n4980), .ZN(n10637) );
  NOR2_X1 U8849 ( .A1(n7640), .A2(n10632), .ZN(n7641) );
  OR2_X1 U8850 ( .A1(n7823), .A2(n7641), .ZN(n10634) );
  INV_X1 U8851 ( .A(n8076), .ZN(n7642) );
  AOI22_X1 U8852 ( .A1(n4856), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n10128), .B2(
        n7642), .ZN(n7644) );
  NAND2_X1 U8853 ( .A1(n8078), .A2(n10165), .ZN(n7643) );
  OAI211_X1 U8854 ( .C1(n10634), .C2(n10167), .A(n7644), .B(n7643), .ZN(n7645)
         );
  AOI21_X1 U8855 ( .B1(n10637), .B2(n10050), .A(n7645), .ZN(n7646) );
  OAI21_X1 U8856 ( .B1(n7647), .B2(n4856), .A(n7646), .ZN(P1_U3280) );
  XNOR2_X1 U8857 ( .A(n7648), .B(n10527), .ZN(n10529) );
  OAI22_X1 U8858 ( .A1(n9620), .A2(n8395), .B1(n8955), .B2(n9592), .ZN(n7654)
         );
  NAND2_X1 U8859 ( .A1(n7603), .A2(n7649), .ZN(n7651) );
  AND2_X1 U8860 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  NAND2_X1 U8861 ( .A1(n7652), .A2(n8499), .ZN(n10530) );
  AND3_X1 U8862 ( .A1(n10531), .A2(n9605), .A3(n10530), .ZN(n7653) );
  AOI211_X1 U8863 ( .C1(n9632), .C2(n10529), .A(n7654), .B(n7653), .ZN(n7661)
         );
  XNOR2_X1 U8864 ( .A(n8499), .B(n7655), .ZN(n7658) );
  OAI22_X1 U8865 ( .A1(n9375), .A2(n9597), .B1(n7656), .B2(n9599), .ZN(n7657)
         );
  AOI21_X1 U8866 ( .B1(n7658), .B2(n9629), .A(n7657), .ZN(n10534) );
  MUX2_X1 U8867 ( .A(n7659), .B(n10534), .S(n9457), .Z(n7660) );
  NAND2_X1 U8868 ( .A1(n7661), .A2(n7660), .ZN(P2_U3290) );
  OAI21_X1 U8869 ( .B1(n8502), .B2(n4923), .A(n7662), .ZN(n7663) );
  AOI222_X1 U8870 ( .A1(n9629), .A2(n7663), .B1(n10608), .B2(n9626), .C1(
        n10558), .C2(n9624), .ZN(n10577) );
  INV_X1 U8871 ( .A(n10528), .ZN(n10678) );
  AOI21_X1 U8872 ( .B1(n7682), .B2(n10555), .A(n10678), .ZN(n7665) );
  NAND2_X1 U8873 ( .A1(n7665), .A2(n7664), .ZN(n10575) );
  AND2_X1 U8874 ( .A1(n9457), .A2(n9601), .ZN(n9511) );
  INV_X1 U8875 ( .A(n9511), .ZN(n7712) );
  OAI22_X1 U8876 ( .A1(n9457), .A2(n7132), .B1(n10572), .B2(n9592), .ZN(n7666)
         );
  AOI21_X1 U8877 ( .B1(n9606), .B2(n10555), .A(n7666), .ZN(n7667) );
  OAI21_X1 U8878 ( .B1(n10575), .B2(n7712), .A(n7667), .ZN(n7668) );
  INV_X1 U8879 ( .A(n7668), .ZN(n7673) );
  NAND2_X1 U8880 ( .A1(n7669), .A2(n7670), .ZN(n7671) );
  NAND2_X1 U8881 ( .A1(n7671), .A2(n8502), .ZN(n10573) );
  NAND3_X1 U8882 ( .A1(n7586), .A2(n9605), .A3(n10573), .ZN(n7672) );
  OAI211_X1 U8883 ( .C1(n10577), .C2(n9618), .A(n7673), .B(n7672), .ZN(
        P2_U3288) );
  XNOR2_X1 U8884 ( .A(n7674), .B(n8501), .ZN(n7677) );
  NAND2_X1 U8885 ( .A1(n10536), .A2(n9624), .ZN(n7675) );
  OAI21_X1 U8886 ( .B1(n10538), .B2(n9599), .A(n7675), .ZN(n7676) );
  AOI21_X1 U8887 ( .B1(n7677), .B2(n9629), .A(n7676), .ZN(n10552) );
  NAND2_X1 U8888 ( .A1(n7678), .A2(n8501), .ZN(n7679) );
  NAND2_X1 U8889 ( .A1(n7669), .A2(n7679), .ZN(n10550) );
  OR2_X1 U8890 ( .A1(n7680), .A2(n10547), .ZN(n7681) );
  NAND2_X1 U8891 ( .A1(n7682), .A2(n7681), .ZN(n10548) );
  OAI22_X1 U8892 ( .A1(n9457), .A2(n7683), .B1(n10546), .B2(n9592), .ZN(n7684)
         );
  AOI21_X1 U8893 ( .B1(n9606), .B2(n10544), .A(n7684), .ZN(n7685) );
  OAI21_X1 U8894 ( .B1(n9451), .B2(n10548), .A(n7685), .ZN(n7686) );
  AOI21_X1 U8895 ( .B1(n10550), .B2(n9605), .A(n7686), .ZN(n7687) );
  OAI21_X1 U8896 ( .B1(n10552), .B2(n9618), .A(n7687), .ZN(P2_U3289) );
  NAND2_X1 U8897 ( .A1(n7688), .A2(n8495), .ZN(n7689) );
  NAND3_X1 U8898 ( .A1(n7690), .A2(n9629), .A3(n7689), .ZN(n7694) );
  OAI22_X1 U8899 ( .A1(n9375), .A2(n9599), .B1(n7691), .B2(n9597), .ZN(n7692)
         );
  INV_X1 U8900 ( .A(n7692), .ZN(n7693) );
  NAND2_X1 U8901 ( .A1(n7694), .A2(n7693), .ZN(n10509) );
  INV_X1 U8902 ( .A(n10509), .ZN(n7704) );
  OAI21_X1 U8903 ( .B1(n7695), .B2(n8495), .A(n7603), .ZN(n10511) );
  INV_X1 U8904 ( .A(n7696), .ZN(n7698) );
  OAI21_X1 U8905 ( .B1(n7698), .B2(n10507), .A(n7697), .ZN(n10508) );
  OAI22_X1 U8906 ( .A1(n7128), .A2(n9457), .B1(n7699), .B2(n9592), .ZN(n7700)
         );
  AOI21_X1 U8907 ( .B1(n9606), .B2(n8382), .A(n7700), .ZN(n7701) );
  OAI21_X1 U8908 ( .B1(n9451), .B2(n10508), .A(n7701), .ZN(n7702) );
  AOI21_X1 U8909 ( .B1(n9605), .B2(n10511), .A(n7702), .ZN(n7703) );
  OAI21_X1 U8910 ( .B1(n9618), .B2(n7704), .A(n7703), .ZN(P2_U3292) );
  NAND2_X1 U8911 ( .A1(n7705), .A2(n8415), .ZN(n7707) );
  OR2_X1 U8912 ( .A1(n7908), .A2(n10612), .ZN(n8421) );
  NAND2_X1 U8913 ( .A1(n7908), .A2(n10612), .ZN(n8416) );
  NAND2_X1 U8914 ( .A1(n8421), .A2(n8416), .ZN(n8506) );
  INV_X1 U8915 ( .A(n8506), .ZN(n7706) );
  NAND2_X1 U8916 ( .A1(n7707), .A2(n7706), .ZN(n7899) );
  NAND3_X1 U8917 ( .A1(n7705), .A2(n8506), .A3(n8415), .ZN(n7708) );
  NAND2_X1 U8918 ( .A1(n7899), .A2(n7708), .ZN(n7709) );
  AOI222_X1 U8919 ( .A1(n9629), .A2(n7709), .B1(n9372), .B2(n9624), .C1(n9371), 
        .C2(n9626), .ZN(n10641) );
  OAI22_X1 U8920 ( .A1(n9457), .A2(n7136), .B1(n7710), .B2(n9592), .ZN(n7714)
         );
  NAND2_X1 U8921 ( .A1(n7711), .A2(n10642), .ZN(n7925) );
  OAI211_X1 U8922 ( .C1(n7711), .C2(n10642), .A(n10528), .B(n7925), .ZN(n10640) );
  NOR2_X1 U8923 ( .A1(n10640), .A2(n7712), .ZN(n7713) );
  AOI211_X1 U8924 ( .C1(n9606), .C2(n7908), .A(n7714), .B(n7713), .ZN(n7720)
         );
  NAND2_X1 U8925 ( .A1(n10620), .A2(n9372), .ZN(n7715) );
  NAND2_X1 U8926 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  NAND2_X1 U8927 ( .A1(n7717), .A2(n8506), .ZN(n7910) );
  OAI21_X1 U8928 ( .B1(n7717), .B2(n8506), .A(n7910), .ZN(n7718) );
  INV_X1 U8929 ( .A(n7718), .ZN(n10644) );
  NAND2_X1 U8930 ( .A1(n10644), .A2(n9605), .ZN(n7719) );
  OAI211_X1 U8931 ( .C1(n10641), .C2(n9618), .A(n7720), .B(n7719), .ZN(
        P2_U3285) );
  NAND2_X1 U8932 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9869) );
  INV_X1 U8933 ( .A(n9869), .ZN(n7728) );
  AOI22_X1 U8934 ( .A1(n7724), .A2(n7723), .B1(n7722), .B2(n7721), .ZN(n7873)
         );
  XNOR2_X1 U8935 ( .A(n7873), .B(n7729), .ZN(n7725) );
  NOR2_X1 U8936 ( .A1(n7726), .A2(n7725), .ZN(n7876) );
  AOI211_X1 U8937 ( .C1(n7726), .C2(n7725), .A(n7876), .B(n10395), .ZN(n7727)
         );
  AOI211_X1 U8938 ( .C1(n7729), .C2(n10406), .A(n7728), .B(n7727), .ZN(n7736)
         );
  OAI21_X1 U8939 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7731), .A(n7730), .ZN(
        n7867) );
  XNOR2_X1 U8940 ( .A(n7867), .B(n7875), .ZN(n7732) );
  NOR2_X1 U8941 ( .A1(n7733), .A2(n7732), .ZN(n7868) );
  AOI211_X1 U8942 ( .C1(n7733), .C2(n7732), .A(n7868), .B(n10412), .ZN(n7734)
         );
  AOI21_X1 U8943 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n10407), .A(n7734), .ZN(
        n7735) );
  NAND2_X1 U8944 ( .A1(n7736), .A2(n7735), .ZN(P1_U3256) );
  INV_X1 U8945 ( .A(n9368), .ZN(n8192) );
  NAND2_X1 U8946 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n9412) );
  OAI21_X1 U8947 ( .B1(n10611), .B2(n8192), .A(n9412), .ZN(n7738) );
  AOI21_X1 U8948 ( .B1(n10609), .B2(n8173), .A(n7738), .ZN(n7739) );
  OAI21_X1 U8949 ( .B1(n8168), .B2(n10623), .A(n7739), .ZN(n7740) );
  AOI21_X1 U8950 ( .B1(n9718), .B2(n10621), .A(n7740), .ZN(n7747) );
  INV_X1 U8951 ( .A(n7742), .ZN(n7745) );
  OAI22_X1 U8952 ( .A1(n7743), .A2(n10615), .B1(n8970), .B2(n9129), .ZN(n7744)
         );
  NAND3_X1 U8953 ( .A1(n7741), .A2(n7745), .A3(n7744), .ZN(n7746) );
  OAI211_X1 U8954 ( .C1(n7737), .C2(n10615), .A(n7747), .B(n7746), .ZN(
        P2_U3243) );
  INV_X1 U8955 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7761) );
  AND2_X1 U8956 ( .A1(n7750), .A2(n7748), .ZN(n7752) );
  NAND2_X1 U8957 ( .A1(n7750), .A2(n7749), .ZN(n7751) );
  OAI21_X1 U8958 ( .B1(n7752), .B2(n8659), .A(n7751), .ZN(n8283) );
  INV_X1 U8959 ( .A(n8659), .ZN(n8556) );
  XNOR2_X1 U8960 ( .A(n8037), .B(n8556), .ZN(n7755) );
  OR2_X1 U8961 ( .A1(n8283), .A2(n6896), .ZN(n7754) );
  AOI22_X1 U8962 ( .A1(n10120), .A2(n9897), .B1(n10146), .B2(n9895), .ZN(n7753) );
  OAI211_X1 U8963 ( .C1(n10107), .C2(n7755), .A(n7754), .B(n7753), .ZN(n8276)
         );
  INV_X1 U8964 ( .A(n8276), .ZN(n7759) );
  NAND2_X1 U8965 ( .A1(n7756), .A2(n8277), .ZN(n7757) );
  AND2_X1 U8966 ( .A1(n8043), .A2(n7757), .ZN(n8280) );
  AOI22_X1 U8967 ( .A1(n8280), .A2(n10250), .B1(n10597), .B2(n8277), .ZN(n7758) );
  OAI211_X1 U8968 ( .C1(n10600), .C2(n8283), .A(n7759), .B(n7758), .ZN(n7762)
         );
  NAND2_X1 U8969 ( .A1(n7762), .A2(n4855), .ZN(n7760) );
  OAI21_X1 U8970 ( .B1(n4855), .B2(n7761), .A(n7760), .ZN(P1_U3478) );
  NAND2_X1 U8971 ( .A1(n7762), .A2(n10656), .ZN(n7763) );
  OAI21_X1 U8972 ( .B1(n10656), .B2(n7764), .A(n7763), .ZN(P1_U3531) );
  INV_X1 U8973 ( .A(n7772), .ZN(n7767) );
  NOR3_X1 U8974 ( .A1(n7765), .A2(n10612), .A3(n9129), .ZN(n7766) );
  AOI21_X1 U8975 ( .B1(n7767), .B2(n10561), .A(n7766), .ZN(n7776) );
  OAI21_X1 U8976 ( .B1(n10611), .B2(n8991), .A(n7768), .ZN(n7769) );
  AOI21_X1 U8977 ( .B1(n10609), .B2(n7907), .A(n7769), .ZN(n7770) );
  OAI21_X1 U8978 ( .B1(n7929), .B2(n10623), .A(n7770), .ZN(n7774) );
  NAND2_X1 U8979 ( .A1(n7772), .A2(n7771), .ZN(n8980) );
  NOR2_X1 U8980 ( .A1(n8980), .A2(n10615), .ZN(n7773) );
  AOI211_X1 U8981 ( .C1(n10621), .C2(n7932), .A(n7774), .B(n7773), .ZN(n7775)
         );
  OAI21_X1 U8982 ( .B1(n7777), .B2(n7776), .A(n7775), .ZN(P2_U3226) );
  NAND2_X1 U8983 ( .A1(n7780), .A2(n9740), .ZN(n7778) );
  OAI211_X1 U8984 ( .C1(n7779), .C2(n4858), .A(n7778), .B(n8535), .ZN(P2_U3335) );
  NAND2_X1 U8985 ( .A1(n7780), .A2(n10289), .ZN(n7782) );
  OR2_X1 U8986 ( .A1(n7781), .A2(P1_U3084), .ZN(n8824) );
  OAI211_X1 U8987 ( .C1(n7783), .C2(n10286), .A(n7782), .B(n8824), .ZN(
        P1_U3330) );
  NAND2_X1 U8988 ( .A1(n7785), .A2(n7784), .ZN(n7805) );
  NAND2_X1 U8989 ( .A1(n8277), .A2(n8234), .ZN(n7787) );
  NAND2_X1 U8990 ( .A1(n9042), .A2(n9896), .ZN(n7786) );
  NAND2_X1 U8991 ( .A1(n7787), .A2(n7786), .ZN(n7788) );
  XNOR2_X1 U8992 ( .A(n7788), .B(n8946), .ZN(n7942) );
  AND2_X1 U8993 ( .A1(n7805), .A2(n7942), .ZN(n7789) );
  INV_X1 U8994 ( .A(n7942), .ZN(n7791) );
  NOR2_X1 U8995 ( .A1(n8040), .A2(n9019), .ZN(n7790) );
  AOI21_X1 U8996 ( .B1(n8277), .B2(n9042), .A(n7790), .ZN(n7941) );
  NAND2_X1 U8997 ( .A1(n10581), .A2(n8234), .ZN(n7793) );
  NAND2_X1 U8998 ( .A1(n9042), .A2(n9895), .ZN(n7792) );
  NAND2_X1 U8999 ( .A1(n7793), .A2(n7792), .ZN(n7794) );
  XNOR2_X1 U9000 ( .A(n7794), .B(n9017), .ZN(n7797) );
  NOR2_X1 U9001 ( .A1(n7795), .A2(n9019), .ZN(n7796) );
  AOI21_X1 U9002 ( .B1(n10581), .B2(n9042), .A(n7796), .ZN(n7798) );
  NAND2_X1 U9003 ( .A1(n7797), .A2(n7798), .ZN(n8021) );
  INV_X1 U9004 ( .A(n7797), .ZN(n7800) );
  INV_X1 U9005 ( .A(n7798), .ZN(n7799) );
  NAND2_X1 U9006 ( .A1(n7800), .A2(n7799), .ZN(n7801) );
  AND2_X1 U9007 ( .A1(n8021), .A2(n7801), .ZN(n7812) );
  INV_X1 U9008 ( .A(n7803), .ZN(n7804) );
  NAND2_X1 U9009 ( .A1(n7806), .A2(n7805), .ZN(n7940) );
  INV_X1 U9010 ( .A(n7940), .ZN(n7808) );
  NAND2_X1 U9011 ( .A1(n7808), .A2(n7807), .ZN(n7811) );
  NAND2_X1 U9012 ( .A1(n7809), .A2(n7811), .ZN(n8022) );
  INV_X1 U9013 ( .A(n8022), .ZN(n7814) );
  AOI21_X1 U9014 ( .B1(n7810), .B2(n7945), .A(n7812), .ZN(n7813) );
  OAI21_X1 U9015 ( .B1(n7814), .B2(n7813), .A(n9815), .ZN(n7820) );
  AOI21_X1 U9016 ( .B1(n9853), .B2(n9894), .A(n7815), .ZN(n7817) );
  NAND2_X1 U9017 ( .A1(n9873), .A2(n9896), .ZN(n7816) );
  OAI211_X1 U9018 ( .C1(n9876), .C2(n8046), .A(n7817), .B(n7816), .ZN(n7818)
         );
  AOI21_X1 U9019 ( .B1(n10581), .B2(n9863), .A(n7818), .ZN(n7819) );
  NAND2_X1 U9020 ( .A1(n7820), .A2(n7819), .ZN(P1_U3229) );
  XOR2_X1 U9021 ( .A(n7821), .B(n8665), .Z(n7822) );
  OAI222_X1 U9022 ( .A1(n10111), .A2(n9754), .B1(n10149), .B2(n8062), .C1(
        n7822), .C2(n10107), .ZN(n10654) );
  OAI21_X1 U9023 ( .B1(n7823), .B2(n10652), .A(n10250), .ZN(n7824) );
  OR2_X1 U9024 ( .A1(n7890), .A2(n7824), .ZN(n10649) );
  INV_X1 U9025 ( .A(n8220), .ZN(n7825) );
  AOI22_X1 U9026 ( .A1(n4856), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n10128), .B2(
        n7825), .ZN(n7827) );
  NAND2_X1 U9027 ( .A1(n8203), .A2(n10165), .ZN(n7826) );
  OAI211_X1 U9028 ( .C1(n10649), .C2(n8050), .A(n7827), .B(n7826), .ZN(n7830)
         );
  NAND2_X1 U9029 ( .A1(n7828), .A2(n8665), .ZN(n10647) );
  AND3_X1 U9030 ( .A1(n10648), .A2(n10050), .A3(n10647), .ZN(n7829) );
  AOI211_X1 U9031 ( .C1(n10163), .C2(n10654), .A(n7830), .B(n7829), .ZN(n7831)
         );
  INV_X1 U9032 ( .A(n7831), .ZN(P1_U3279) );
  INV_X1 U9033 ( .A(n8138), .ZN(n7833) );
  OAI22_X1 U9034 ( .A1(n8182), .A2(n9599), .B1(n8134), .B2(n9597), .ZN(n8147)
         );
  AOI22_X1 U9035 ( .A1(n9137), .A2(n8147), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n7832) );
  OAI21_X1 U9036 ( .B1(n7833), .B2(n10623), .A(n7832), .ZN(n7834) );
  AOI21_X1 U9037 ( .B1(n9714), .B2(n10621), .A(n7834), .ZN(n7839) );
  OAI22_X1 U9038 ( .A1(n7836), .A2(n10615), .B1(n8134), .B2(n9129), .ZN(n7837)
         );
  NAND3_X1 U9039 ( .A1(n7737), .A2(n5223), .A3(n7837), .ZN(n7838) );
  OAI211_X1 U9040 ( .C1(n7840), .C2(n10615), .A(n7839), .B(n7838), .ZN(
        P2_U3228) );
  INV_X1 U9041 ( .A(n7841), .ZN(n7865) );
  OAI222_X1 U9042 ( .A1(n8538), .A2(n7865), .B1(P2_U3152), .B2(n7843), .C1(
        n7842), .C2(n4858), .ZN(P2_U3334) );
  AOI21_X1 U9043 ( .B1(n7845), .B2(n6278), .A(n7844), .ZN(n7846) );
  NAND2_X1 U9044 ( .A1(n9417), .A2(n7846), .ZN(n7847) );
  XNOR2_X1 U9045 ( .A(n7846), .B(n7856), .ZN(n9411) );
  NAND2_X1 U9046 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9411), .ZN(n9410) );
  NAND2_X1 U9047 ( .A1(n7847), .A2(n9410), .ZN(n7851) );
  INV_X1 U9048 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U9049 ( .A1(n7849), .A2(n7848), .ZN(n7987) );
  OAI21_X1 U9050 ( .B1(n7849), .B2(n7848), .A(n7987), .ZN(n7850) );
  NOR2_X1 U9051 ( .A1(n7851), .A2(n7850), .ZN(n7989) );
  AOI21_X1 U9052 ( .B1(n7851), .B2(n7850), .A(n7989), .ZN(n7864) );
  NOR2_X1 U9053 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6304), .ZN(n7852) );
  AOI21_X1 U9054 ( .B1(n10448), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7852), .ZN(
        n7853) );
  INV_X1 U9055 ( .A(n7853), .ZN(n7862) );
  OAI21_X1 U9056 ( .B1(n7855), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7854), .ZN(
        n7857) );
  NAND2_X1 U9057 ( .A1(n7856), .A2(n7857), .ZN(n7858) );
  XNOR2_X1 U9058 ( .A(n7857), .B(n9417), .ZN(n9415) );
  NAND2_X1 U9059 ( .A1(n9415), .A2(n6289), .ZN(n9414) );
  NAND2_X1 U9060 ( .A1(n7858), .A2(n9414), .ZN(n7860) );
  XNOR2_X1 U9061 ( .A(n7983), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n7859) );
  NOR2_X1 U9062 ( .A1(n7860), .A2(n7859), .ZN(n7982) );
  AOI211_X1 U9063 ( .C1(n7860), .C2(n7859), .A(n10449), .B(n7982), .ZN(n7861)
         );
  AOI211_X1 U9064 ( .C1(n10455), .C2(n7983), .A(n7862), .B(n7861), .ZN(n7863)
         );
  OAI21_X1 U9065 ( .B1(n7864), .B2(n10427), .A(n7863), .ZN(P2_U3261) );
  OAI222_X1 U9066 ( .A1(P1_U3084), .A2(n7866), .B1(n10286), .B2(n5788), .C1(
        n7865), .C2(n9064), .ZN(P1_U3329) );
  NOR2_X1 U9067 ( .A1(n7875), .A2(n7867), .ZN(n7869) );
  NOR2_X1 U9068 ( .A1(n7869), .A2(n7868), .ZN(n7872) );
  NAND2_X1 U9069 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9908), .ZN(n7870) );
  OAI21_X1 U9070 ( .B1(n9908), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7870), .ZN(
        n7871) );
  NOR2_X1 U9071 ( .A1(n7872), .A2(n7871), .ZN(n9907) );
  AOI211_X1 U9072 ( .C1(n7872), .C2(n7871), .A(n9907), .B(n10412), .ZN(n7884)
         );
  INV_X1 U9073 ( .A(n7873), .ZN(n7874) );
  NOR2_X1 U9074 ( .A1(n7875), .A2(n7874), .ZN(n7877) );
  NOR2_X1 U9075 ( .A1(n7877), .A2(n7876), .ZN(n7879) );
  XNOR2_X1 U9076 ( .A(n9908), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7878) );
  NOR2_X1 U9077 ( .A1(n7879), .A2(n7878), .ZN(n9902) );
  AOI211_X1 U9078 ( .C1(n7879), .C2(n7878), .A(n9902), .B(n10395), .ZN(n7883)
         );
  NAND2_X1 U9079 ( .A1(n10407), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7880) );
  NAND2_X1 U9080 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9801) );
  OAI211_X1 U9081 ( .C1(n7881), .C2(n9943), .A(n7880), .B(n9801), .ZN(n7882)
         );
  OR3_X1 U9082 ( .A1(n7884), .A2(n7883), .A3(n7882), .ZN(P1_U3257) );
  OAI21_X1 U9083 ( .B1(n8649), .B2(n7885), .A(n7963), .ZN(n7886) );
  AOI222_X1 U9084 ( .A1(n10152), .A2(n7886), .B1(n9890), .B2(n10146), .C1(
        n9892), .C2(n10120), .ZN(n10263) );
  INV_X1 U9085 ( .A(n7887), .ZN(n7888) );
  AOI21_X1 U9086 ( .B1(n8649), .B2(n7889), .A(n7888), .ZN(n10264) );
  INV_X1 U9087 ( .A(n10264), .ZN(n7897) );
  OR2_X1 U9088 ( .A1(n7890), .A2(n7895), .ZN(n7891) );
  AND3_X1 U9089 ( .A1(n7891), .A2(n7967), .A3(n10250), .ZN(n10260) );
  NAND2_X1 U9090 ( .A1(n10260), .A2(n10117), .ZN(n7894) );
  INV_X1 U9091 ( .A(n8245), .ZN(n7892) );
  AOI22_X1 U9092 ( .A1(n4856), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n10128), .B2(
        n7892), .ZN(n7893) );
  OAI211_X1 U9093 ( .C1(n7895), .C2(n10130), .A(n7894), .B(n7893), .ZN(n7896)
         );
  AOI21_X1 U9094 ( .B1(n7897), .B2(n10050), .A(n7896), .ZN(n7898) );
  OAI21_X1 U9095 ( .B1(n4856), .B2(n10263), .A(n7898), .ZN(P1_U3278) );
  NAND2_X1 U9096 ( .A1(n7899), .A2(n8416), .ZN(n7900) );
  OR2_X1 U9097 ( .A1(n7932), .A2(n8976), .ZN(n8425) );
  NAND2_X1 U9098 ( .A1(n7932), .A2(n8976), .ZN(n8426) );
  NAND2_X1 U9099 ( .A1(n7900), .A2(n8508), .ZN(n7921) );
  NAND2_X1 U9100 ( .A1(n7921), .A2(n8426), .ZN(n7901) );
  OR2_X1 U9101 ( .A1(n8975), .A2(n8991), .ZN(n8433) );
  NAND2_X1 U9102 ( .A1(n8975), .A2(n8991), .ZN(n8432) );
  NAND2_X1 U9103 ( .A1(n8433), .A2(n8432), .ZN(n7913) );
  INV_X1 U9104 ( .A(n7913), .ZN(n8509) );
  NAND2_X1 U9105 ( .A1(n7901), .A2(n8509), .ZN(n8144) );
  NAND3_X1 U9106 ( .A1(n7921), .A2(n7913), .A3(n8426), .ZN(n7902) );
  AND2_X1 U9107 ( .A1(n8144), .A2(n7902), .ZN(n7903) );
  OAI222_X1 U9108 ( .A1(n9597), .A2(n8976), .B1(n9599), .B2(n8970), .C1(n9594), 
        .C2(n7903), .ZN(n10670) );
  INV_X1 U9109 ( .A(n10670), .ZN(n7918) );
  OAI22_X1 U9110 ( .A1(n9457), .A2(n6232), .B1(n8973), .B2(n9592), .ZN(n7906)
         );
  INV_X1 U9111 ( .A(n8137), .ZN(n7904) );
  OAI21_X1 U9112 ( .B1(n10668), .B2(n7926), .A(n7904), .ZN(n10669) );
  NOR2_X1 U9113 ( .A1(n10669), .A2(n9451), .ZN(n7905) );
  AOI211_X1 U9114 ( .C1(n9606), .C2(n8975), .A(n7906), .B(n7905), .ZN(n7917)
         );
  NAND2_X1 U9115 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  OR2_X1 U9116 ( .A1(n7932), .A2(n9371), .ZN(n7912) );
  NOR2_X1 U9117 ( .A1(n7914), .A2(n7913), .ZN(n10667) );
  INV_X1 U9118 ( .A(n10667), .ZN(n7915) );
  NAND3_X1 U9119 ( .A1(n7915), .A2(n9605), .A3(n7973), .ZN(n7916) );
  OAI211_X1 U9120 ( .C1(n7918), .C2(n9618), .A(n7917), .B(n7916), .ZN(P2_U3283) );
  OAI21_X1 U9121 ( .B1(n7920), .B2(n7911), .A(n7919), .ZN(n10664) );
  INV_X1 U9122 ( .A(n10664), .ZN(n7936) );
  INV_X1 U9123 ( .A(n8416), .ZN(n8424) );
  NOR2_X1 U9124 ( .A1(n8508), .A2(n8424), .ZN(n7923) );
  INV_X1 U9125 ( .A(n7921), .ZN(n7922) );
  AOI21_X1 U9126 ( .B1(n7923), .B2(n7899), .A(n7922), .ZN(n7924) );
  OAI222_X1 U9127 ( .A1(n9597), .A2(n10612), .B1(n9599), .B2(n8991), .C1(n9594), .C2(n7924), .ZN(n10662) );
  INV_X1 U9128 ( .A(n7932), .ZN(n10660) );
  INV_X1 U9129 ( .A(n7925), .ZN(n7928) );
  INV_X1 U9130 ( .A(n7926), .ZN(n7927) );
  OAI21_X1 U9131 ( .B1(n10660), .B2(n7928), .A(n7927), .ZN(n10661) );
  OAI22_X1 U9132 ( .A1(n9457), .A2(n7930), .B1(n7929), .B2(n9592), .ZN(n7931)
         );
  AOI21_X1 U9133 ( .B1(n7932), .B2(n9606), .A(n7931), .ZN(n7933) );
  OAI21_X1 U9134 ( .B1(n10661), .B2(n9451), .A(n7933), .ZN(n7934) );
  AOI21_X1 U9135 ( .B1(n10662), .B2(n9457), .A(n7934), .ZN(n7935) );
  OAI21_X1 U9136 ( .B1(n7936), .B2(n9634), .A(n7935), .ZN(P2_U3284) );
  AOI21_X1 U9137 ( .B1(n9853), .B2(n9895), .A(n7937), .ZN(n7939) );
  NAND2_X1 U9138 ( .A1(n9873), .A2(n9897), .ZN(n7938) );
  OAI211_X1 U9139 ( .C1(n9876), .C2(n8278), .A(n7939), .B(n7938), .ZN(n7948)
         );
  INV_X1 U9140 ( .A(n7810), .ZN(n7946) );
  NAND2_X1 U9141 ( .A1(n7940), .A2(n7941), .ZN(n7943) );
  AOI21_X1 U9142 ( .B1(n7945), .B2(n7943), .A(n7942), .ZN(n7944) );
  AOI211_X1 U9143 ( .C1(n7946), .C2(n7945), .A(n9879), .B(n7944), .ZN(n7947)
         );
  AOI211_X1 U9144 ( .C1(n8277), .C2(n9863), .A(n7948), .B(n7947), .ZN(n7949)
         );
  INV_X1 U9145 ( .A(n7949), .ZN(P1_U3219) );
  INV_X1 U9146 ( .A(n7950), .ZN(n7952) );
  NAND2_X1 U9147 ( .A1(n7952), .A2(n7951), .ZN(n7953) );
  XNOR2_X1 U9148 ( .A(n7954), .B(n7953), .ZN(n7959) );
  NOR2_X1 U9149 ( .A1(n10623), .A2(n8186), .ZN(n7957) );
  NAND2_X1 U9150 ( .A1(n10609), .A2(n9368), .ZN(n7955) );
  NAND2_X1 U9151 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n8008) );
  OAI211_X1 U9152 ( .C1(n9596), .C2(n10611), .A(n7955), .B(n8008), .ZN(n7956)
         );
  AOI211_X1 U9153 ( .C1(n9710), .C2(n10621), .A(n7957), .B(n7956), .ZN(n7958)
         );
  OAI21_X1 U9154 ( .B1(n7959), .B2(n10615), .A(n7958), .ZN(P2_U3230) );
  XOR2_X1 U9155 ( .A(n7960), .B(n8667), .Z(n10259) );
  NAND2_X1 U9156 ( .A1(n7961), .A2(n10152), .ZN(n7966) );
  INV_X1 U9157 ( .A(n8667), .ZN(n7962) );
  AOI21_X1 U9158 ( .B1(n7963), .B2(n8707), .A(n7962), .ZN(n7965) );
  AOI22_X1 U9159 ( .A1(n10146), .A2(n9889), .B1(n10120), .B2(n9891), .ZN(n7964) );
  OAI21_X1 U9160 ( .B1(n7966), .B2(n7965), .A(n7964), .ZN(n10255) );
  INV_X1 U9161 ( .A(n10257), .ZN(n7970) );
  AOI211_X1 U9162 ( .C1(n10257), .C2(n7967), .A(n10633), .B(n5180), .ZN(n10256) );
  NAND2_X1 U9163 ( .A1(n10256), .A2(n10117), .ZN(n7969) );
  AOI22_X1 U9164 ( .A1(n4856), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n10128), .B2(
        n9750), .ZN(n7968) );
  OAI211_X1 U9165 ( .C1(n7970), .C2(n10130), .A(n7969), .B(n7968), .ZN(n7971)
         );
  AOI21_X1 U9166 ( .B1(n10255), .B2(n10163), .A(n7971), .ZN(n7972) );
  OAI21_X1 U9167 ( .B1(n10259), .B2(n10134), .A(n7972), .ZN(P1_U3277) );
  NAND2_X1 U9168 ( .A1(n8989), .A2(n8970), .ZN(n8437) );
  NAND2_X1 U9169 ( .A1(n7973), .A2(n5314), .ZN(n7974) );
  AOI21_X1 U9170 ( .B1(n8510), .B2(n7974), .A(n8133), .ZN(n10675) );
  NAND2_X1 U9171 ( .A1(n8144), .A2(n8432), .ZN(n7975) );
  INV_X1 U9172 ( .A(n8510), .ZN(n8142) );
  XNOR2_X1 U9173 ( .A(n7975), .B(n8142), .ZN(n7976) );
  OAI222_X1 U9174 ( .A1(n9597), .A2(n8991), .B1(n9599), .B2(n8134), .C1(n7976), 
        .C2(n9594), .ZN(n10681) );
  XNOR2_X1 U9175 ( .A(n10677), .B(n8137), .ZN(n10679) );
  OAI22_X1 U9176 ( .A1(n9457), .A2(n7977), .B1(n8983), .B2(n9592), .ZN(n7978)
         );
  AOI21_X1 U9177 ( .B1(n8989), .B2(n9606), .A(n7978), .ZN(n7979) );
  OAI21_X1 U9178 ( .B1(n10679), .B2(n9451), .A(n7979), .ZN(n7980) );
  AOI21_X1 U9179 ( .B1(n10681), .B2(n9517), .A(n7980), .ZN(n7981) );
  OAI21_X1 U9180 ( .B1(n10675), .B2(n9634), .A(n7981), .ZN(P2_U3282) );
  AOI21_X1 U9181 ( .B1(n7983), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7982), .ZN(
        n8013) );
  OR2_X1 U9182 ( .A1(n8016), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U9183 ( .A1(n8016), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U9184 ( .A1(n7985), .A2(n7984), .ZN(n8012) );
  NOR2_X1 U9185 ( .A1(n8013), .A2(n8012), .ZN(n8011) );
  AOI21_X1 U9186 ( .B1(n8016), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8011), .ZN(
        n8115) );
  XNOR2_X1 U9187 ( .A(n8119), .B(P2_REG2_REG_18__SCAN_IN), .ZN(n7986) );
  XNOR2_X1 U9188 ( .A(n8115), .B(n7986), .ZN(n8005) );
  INV_X1 U9189 ( .A(n7987), .ZN(n7988) );
  NOR2_X1 U9190 ( .A1(n7989), .A2(n7988), .ZN(n8006) );
  XNOR2_X1 U9191 ( .A(n8016), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8007) );
  INV_X1 U9192 ( .A(n8007), .ZN(n7990) );
  NAND2_X1 U9193 ( .A1(n8006), .A2(n7990), .ZN(n7991) );
  OAI21_X1 U9194 ( .B1(n7993), .B2(n7992), .A(n7991), .ZN(n7996) );
  INV_X1 U9195 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U9196 ( .A1(n8116), .A2(n7994), .ZN(n8122) );
  OAI21_X1 U9197 ( .B1(n8116), .B2(n7994), .A(n8122), .ZN(n7995) );
  NOR2_X1 U9198 ( .A1(n7995), .A2(n7996), .ZN(n8124) );
  AOI21_X1 U9199 ( .B1(n7996), .B2(n7995), .A(n8124), .ZN(n7997) );
  NOR2_X1 U9200 ( .A1(n10427), .A2(n7997), .ZN(n8003) );
  INV_X1 U9201 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8000) );
  NOR2_X1 U9202 ( .A1(n7998), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8089) );
  INV_X1 U9203 ( .A(n8089), .ZN(n7999) );
  OAI21_X1 U9204 ( .B1(n8001), .B2(n8000), .A(n7999), .ZN(n8002) );
  AOI211_X1 U9205 ( .C1(n10455), .C2(n8119), .A(n8003), .B(n8002), .ZN(n8004)
         );
  OAI21_X1 U9206 ( .B1(n8005), .B2(n10449), .A(n8004), .ZN(P2_U3263) );
  XOR2_X1 U9207 ( .A(n8007), .B(n8006), .Z(n8018) );
  INV_X1 U9208 ( .A(n8008), .ZN(n8009) );
  AOI21_X1 U9209 ( .B1(n10448), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8009), .ZN(
        n8010) );
  INV_X1 U9210 ( .A(n8010), .ZN(n8015) );
  AOI211_X1 U9211 ( .C1(n8013), .C2(n8012), .A(n10449), .B(n8011), .ZN(n8014)
         );
  AOI211_X1 U9212 ( .C1(n10455), .C2(n8016), .A(n8015), .B(n8014), .ZN(n8017)
         );
  OAI21_X1 U9213 ( .B1(n10427), .B2(n8018), .A(n8017), .ZN(P2_U3262) );
  NAND2_X1 U9214 ( .A1(n10596), .A2(n9042), .ZN(n8020) );
  NAND2_X1 U9215 ( .A1(n9046), .A2(n9894), .ZN(n8019) );
  NAND2_X1 U9216 ( .A1(n8020), .A2(n8019), .ZN(n8069) );
  NAND2_X1 U9217 ( .A1(n8022), .A2(n8021), .ZN(n8029) );
  INV_X1 U9218 ( .A(n8029), .ZN(n8027) );
  NAND2_X1 U9219 ( .A1(n10596), .A2(n8234), .ZN(n8024) );
  NAND2_X1 U9220 ( .A1(n9042), .A2(n9894), .ZN(n8023) );
  NAND2_X1 U9221 ( .A1(n8024), .A2(n8023), .ZN(n8025) );
  XNOR2_X1 U9222 ( .A(n8025), .B(n9017), .ZN(n8028) );
  INV_X1 U9223 ( .A(n8028), .ZN(n8026) );
  NAND2_X1 U9224 ( .A1(n8027), .A2(n8026), .ZN(n8071) );
  NAND2_X1 U9225 ( .A1(n8029), .A2(n8028), .ZN(n8070) );
  NAND2_X1 U9226 ( .A1(n8071), .A2(n8070), .ZN(n8030) );
  XOR2_X1 U9227 ( .A(n8069), .B(n8030), .Z(n8036) );
  INV_X1 U9228 ( .A(n9853), .ZN(n9871) );
  NAND2_X1 U9229 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10403) );
  OAI21_X1 U9230 ( .B1(n9871), .B2(n8062), .A(n10403), .ZN(n8031) );
  AOI21_X1 U9231 ( .B1(n9873), .B2(n9895), .A(n8031), .ZN(n8032) );
  OAI21_X1 U9232 ( .B1(n9876), .B2(n8033), .A(n8032), .ZN(n8034) );
  AOI21_X1 U9233 ( .B1(n10596), .B2(n9863), .A(n8034), .ZN(n8035) );
  OAI21_X1 U9234 ( .B1(n8036), .B2(n9879), .A(n8035), .ZN(P1_U3215) );
  NAND2_X1 U9235 ( .A1(n4919), .A2(n8557), .ZN(n8038) );
  AND2_X1 U9236 ( .A1(n8561), .A2(n8721), .ZN(n8657) );
  XNOR2_X1 U9237 ( .A(n8038), .B(n8657), .ZN(n8039) );
  OAI222_X1 U9238 ( .A1(n10111), .A2(n8041), .B1(n10149), .B2(n8040), .C1(
        n10107), .C2(n8039), .ZN(n10583) );
  INV_X1 U9239 ( .A(n10583), .ZN(n8053) );
  XNOR2_X1 U9240 ( .A(n8042), .B(n8657), .ZN(n10585) );
  AOI21_X1 U9241 ( .B1(n8043), .B2(n10581), .A(n10633), .ZN(n8045) );
  NAND2_X1 U9242 ( .A1(n8045), .A2(n8044), .ZN(n10582) );
  INV_X1 U9243 ( .A(n10117), .ZN(n8050) );
  INV_X1 U9244 ( .A(n8046), .ZN(n8047) );
  AOI22_X1 U9245 ( .A1(n4856), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n10128), .B2(
        n8047), .ZN(n8049) );
  NAND2_X1 U9246 ( .A1(n10581), .A2(n10165), .ZN(n8048) );
  OAI211_X1 U9247 ( .C1(n10582), .C2(n8050), .A(n8049), .B(n8048), .ZN(n8051)
         );
  AOI21_X1 U9248 ( .B1(n10585), .B2(n10050), .A(n8051), .ZN(n8052) );
  OAI21_X1 U9249 ( .B1(n8053), .B2(n4856), .A(n8052), .ZN(P1_U3282) );
  INV_X1 U9250 ( .A(n8054), .ZN(n8057) );
  OAI222_X1 U9251 ( .A1(n4858), .A2(n8056), .B1(n8538), .B2(n8057), .C1(n8055), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9252 ( .A1(P1_U3084), .A2(n8058), .B1(n9064), .B2(n8057), .C1(
        n9060), .C2(n5807), .ZN(P1_U3328) );
  NAND2_X1 U9253 ( .A1(n8078), .A2(n8234), .ZN(n8060) );
  NAND2_X1 U9254 ( .A1(n9042), .A2(n9893), .ZN(n8059) );
  NAND2_X1 U9255 ( .A1(n8060), .A2(n8059), .ZN(n8061) );
  XNOR2_X1 U9256 ( .A(n8061), .B(n9017), .ZN(n8064) );
  NOR2_X1 U9257 ( .A1(n8062), .A2(n9019), .ZN(n8063) );
  AOI21_X1 U9258 ( .B1(n8078), .B2(n9042), .A(n8063), .ZN(n8065) );
  NAND2_X1 U9259 ( .A1(n8064), .A2(n8065), .ZN(n8208) );
  INV_X1 U9260 ( .A(n8064), .ZN(n8067) );
  INV_X1 U9261 ( .A(n8065), .ZN(n8066) );
  NAND2_X1 U9262 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U9263 ( .A1(n8208), .A2(n8068), .ZN(n8207) );
  NAND2_X1 U9264 ( .A1(n8070), .A2(n8069), .ZN(n8072) );
  NAND2_X1 U9265 ( .A1(n8072), .A2(n8071), .ZN(n8206) );
  AOI21_X1 U9266 ( .B1(n8207), .B2(n8206), .A(n5315), .ZN(n8080) );
  NOR2_X1 U9267 ( .A1(n9871), .A2(n8201), .ZN(n8073) );
  AOI211_X1 U9268 ( .C1(n9873), .C2(n9894), .A(n8074), .B(n8073), .ZN(n8075)
         );
  OAI21_X1 U9269 ( .B1(n9876), .B2(n8076), .A(n8075), .ZN(n8077) );
  AOI21_X1 U9270 ( .B1(n8078), .B2(n9863), .A(n8077), .ZN(n8079) );
  OAI21_X1 U9271 ( .B1(n8080), .B2(n9879), .A(n8079), .ZN(P1_U3234) );
  INV_X1 U9272 ( .A(n8081), .ZN(n8095) );
  OAI222_X1 U9273 ( .A1(n8538), .A2(n8095), .B1(P2_U3152), .B2(n8083), .C1(
        n8082), .C2(n4858), .ZN(P2_U3332) );
  INV_X1 U9274 ( .A(n8084), .ZN(n8086) );
  NOR2_X1 U9275 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  XNOR2_X1 U9276 ( .A(n8088), .B(n8087), .ZN(n8094) );
  AOI21_X1 U9277 ( .B1(n10609), .B2(n9625), .A(n8089), .ZN(n8091) );
  NAND2_X1 U9278 ( .A1(n9121), .A2(n9617), .ZN(n8090) );
  OAI211_X1 U9279 ( .C1(n9428), .C2(n10611), .A(n8091), .B(n8090), .ZN(n8092)
         );
  AOI21_X1 U9280 ( .B1(n9703), .B2(n10621), .A(n8092), .ZN(n8093) );
  OAI21_X1 U9281 ( .B1(n8094), .B2(n10615), .A(n8093), .ZN(P2_U3240) );
  OAI222_X1 U9282 ( .A1(P1_U3084), .A2(n8096), .B1(n10286), .B2(n5828), .C1(
        n8095), .C2(n9064), .ZN(P1_U3327) );
  AND2_X1 U9283 ( .A1(n8098), .A2(n8097), .ZN(n8099) );
  XNOR2_X1 U9284 ( .A(n8099), .B(n8104), .ZN(n10248) );
  OAI21_X1 U9285 ( .B1(n8155), .B2(n9803), .A(n10250), .ZN(n8100) );
  NOR2_X1 U9286 ( .A1(n8100), .A2(n8256), .ZN(n10245) );
  AOI22_X1 U9287 ( .A1(n4856), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10128), .B2(
        n9807), .ZN(n8101) );
  OAI21_X1 U9288 ( .B1(n9803), .B2(n10130), .A(n8101), .ZN(n8102) );
  AOI21_X1 U9289 ( .B1(n10245), .B2(n10117), .A(n8102), .ZN(n8107) );
  XNOR2_X1 U9290 ( .A(n8103), .B(n8104), .ZN(n8105) );
  OAI222_X1 U9291 ( .A1(n10111), .A2(n10150), .B1(n10149), .B2(n8853), .C1(
        n8105), .C2(n10107), .ZN(n10244) );
  NAND2_X1 U9292 ( .A1(n10244), .A2(n10163), .ZN(n8106) );
  OAI211_X1 U9293 ( .C1(n10248), .C2(n10134), .A(n8107), .B(n8106), .ZN(
        P1_U3275) );
  NAND2_X1 U9294 ( .A1(n8111), .A2(n10289), .ZN(n8109) );
  OAI211_X1 U9295 ( .C1(n9060), .C2(n8110), .A(n8109), .B(n8108), .ZN(P1_U3326) );
  INV_X1 U9296 ( .A(n8111), .ZN(n8113) );
  OAI222_X1 U9297 ( .A1(n8538), .A2(n8113), .B1(n7063), .B2(P2_U3152), .C1(
        n8112), .C2(n4858), .ZN(P2_U3331) );
  INV_X1 U9298 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8114) );
  MUX2_X1 U9299 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8114), .S(n8339), .Z(n8121)
         );
  INV_X1 U9300 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8117) );
  AOI21_X1 U9301 ( .B1(n8117), .B2(n8116), .A(n8115), .ZN(n8118) );
  AOI21_X1 U9302 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8119), .A(n8118), .ZN(
        n8120) );
  XOR2_X1 U9303 ( .A(n8121), .B(n8120), .Z(n8132) );
  INV_X1 U9304 ( .A(n8122), .ZN(n8123) );
  NOR2_X1 U9305 ( .A1(n8124), .A2(n8123), .ZN(n8126) );
  XNOR2_X1 U9306 ( .A(n9601), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8125) );
  XNOR2_X1 U9307 ( .A(n8126), .B(n8125), .ZN(n8129) );
  NAND2_X1 U9308 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U9309 ( .A1(n10448), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8128) );
  OAI211_X1 U9310 ( .C1(n10427), .C2(n8129), .A(n8228), .B(n8128), .ZN(n8130)
         );
  AOI21_X1 U9311 ( .B1(n10455), .B2(n8339), .A(n8130), .ZN(n8131) );
  OAI21_X1 U9312 ( .B1(n8132), .B2(n10449), .A(n8131), .ZN(P2_U3264) );
  NAND2_X1 U9313 ( .A1(n8140), .A2(n9368), .ZN(n8445) );
  NAND2_X1 U9314 ( .A1(n9714), .A2(n8192), .ZN(n8444) );
  OR2_X1 U9315 ( .A1(n9718), .A2(n8134), .ZN(n8440) );
  NAND2_X1 U9316 ( .A1(n9718), .A2(n8134), .ZN(n8441) );
  INV_X1 U9317 ( .A(n8134), .ZN(n9369) );
  AOI21_X1 U9318 ( .B1(n8513), .B2(n8135), .A(n8181), .ZN(n8136) );
  INV_X1 U9319 ( .A(n8136), .ZN(n9717) );
  AOI211_X1 U9320 ( .C1(n9714), .C2(n8165), .A(n10678), .B(n8309), .ZN(n9713)
         );
  INV_X1 U9321 ( .A(n9592), .ZN(n9616) );
  AOI22_X1 U9322 ( .A1(n9618), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8138), .B2(
        n9616), .ZN(n8139) );
  OAI21_X1 U9323 ( .B1(n8140), .B2(n9620), .A(n8139), .ZN(n8150) );
  INV_X1 U9324 ( .A(n8432), .ZN(n8141) );
  NOR2_X1 U9325 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  NAND2_X1 U9326 ( .A1(n8144), .A2(n8143), .ZN(n8145) );
  NAND2_X1 U9327 ( .A1(n8145), .A2(n8436), .ZN(n8172) );
  INV_X1 U9328 ( .A(n8440), .ZN(n8146) );
  XNOR2_X1 U9329 ( .A(n8190), .B(n8513), .ZN(n8148) );
  AOI21_X1 U9330 ( .B1(n8148), .B2(n9629), .A(n8147), .ZN(n9716) );
  NOR2_X1 U9331 ( .A1(n9716), .A2(n9618), .ZN(n8149) );
  AOI211_X1 U9332 ( .C1(n9713), .C2(n9511), .A(n8150), .B(n8149), .ZN(n8151)
         );
  OAI21_X1 U9333 ( .B1(n9717), .B2(n9634), .A(n8151), .ZN(P2_U3280) );
  NAND2_X1 U9334 ( .A1(n8153), .A2(n8152), .ZN(n8154) );
  XNOR2_X1 U9335 ( .A(n8154), .B(n8668), .ZN(n10254) );
  AOI21_X1 U9336 ( .B1(n10249), .B2(n8156), .A(n8155), .ZN(n10251) );
  INV_X1 U9337 ( .A(n10249), .ZN(n8576) );
  AOI22_X1 U9338 ( .A1(n4856), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10128), .B2(
        n8157), .ZN(n8158) );
  OAI21_X1 U9339 ( .B1(n8576), .B2(n10130), .A(n8158), .ZN(n8162) );
  OAI21_X1 U9340 ( .B1(n5299), .B2(n5644), .A(n8159), .ZN(n8160) );
  AOI222_X1 U9341 ( .A1(n10152), .A2(n8160), .B1(n9888), .B2(n10146), .C1(
        n9890), .C2(n10120), .ZN(n10253) );
  NOR2_X1 U9342 ( .A1(n10253), .A2(n4856), .ZN(n8161) );
  AOI211_X1 U9343 ( .C1(n10251), .C2(n10137), .A(n8162), .B(n8161), .ZN(n8163)
         );
  OAI21_X1 U9344 ( .B1(n10134), .B2(n10254), .A(n8163), .ZN(P1_U3276) );
  XOR2_X1 U9345 ( .A(n8512), .B(n8164), .Z(n9722) );
  INV_X1 U9346 ( .A(n8165), .ZN(n8166) );
  AOI21_X1 U9347 ( .B1(n9718), .B2(n8167), .A(n8166), .ZN(n9719) );
  INV_X1 U9348 ( .A(n9718), .ZN(n8171) );
  INV_X1 U9349 ( .A(n8168), .ZN(n8169) );
  AOI22_X1 U9350 ( .A1(n9618), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8169), .B2(
        n9616), .ZN(n8170) );
  OAI21_X1 U9351 ( .B1(n8171), .B2(n9620), .A(n8170), .ZN(n8176) );
  XOR2_X1 U9352 ( .A(n8512), .B(n8172), .Z(n8174) );
  AOI222_X1 U9353 ( .A1(n9629), .A2(n8174), .B1(n9368), .B2(n9626), .C1(n8173), 
        .C2(n9624), .ZN(n9721) );
  NOR2_X1 U9354 ( .A1(n9721), .A2(n9618), .ZN(n8175) );
  AOI211_X1 U9355 ( .C1(n9719), .C2(n9632), .A(n8176), .B(n8175), .ZN(n8177)
         );
  OAI21_X1 U9356 ( .B1(n9722), .B2(n9634), .A(n8177), .ZN(P2_U3281) );
  NAND2_X1 U9357 ( .A1(n8195), .A2(n10289), .ZN(n8179) );
  OAI211_X1 U9358 ( .C1(n9060), .C2(n8180), .A(n8179), .B(n8178), .ZN(P1_U3325) );
  NAND2_X1 U9359 ( .A1(n9710), .A2(n8182), .ZN(n8362) );
  NAND2_X1 U9360 ( .A1(n8363), .A2(n8362), .ZN(n8364) );
  NAND2_X1 U9361 ( .A1(n8183), .A2(n8364), .ZN(n9427) );
  OAI21_X1 U9362 ( .B1(n8183), .B2(n8364), .A(n9427), .ZN(n8184) );
  INV_X1 U9363 ( .A(n8184), .ZN(n9712) );
  INV_X1 U9364 ( .A(n9710), .ZN(n8310) );
  XNOR2_X1 U9365 ( .A(n8310), .B(n8309), .ZN(n8185) );
  NOR2_X1 U9366 ( .A1(n8185), .A2(n10678), .ZN(n9709) );
  NOR2_X1 U9367 ( .A1(n8310), .A2(n9620), .ZN(n8189) );
  OAI22_X1 U9368 ( .A1(n9457), .A2(n8187), .B1(n8186), .B2(n9592), .ZN(n8188)
         );
  AOI211_X1 U9369 ( .C1(n9709), .C2(n9511), .A(n8189), .B(n8188), .ZN(n8194)
         );
  XNOR2_X1 U9370 ( .A(n8316), .B(n8364), .ZN(n8191) );
  OAI222_X1 U9371 ( .A1(n9599), .A2(n9596), .B1(n9597), .B2(n8192), .C1(n8191), 
        .C2(n9594), .ZN(n9708) );
  NAND2_X1 U9372 ( .A1(n9708), .A2(n9457), .ZN(n8193) );
  OAI211_X1 U9373 ( .C1(n9712), .C2(n9634), .A(n8194), .B(n8193), .ZN(P2_U3279) );
  INV_X1 U9374 ( .A(n8195), .ZN(n8197) );
  OAI222_X1 U9375 ( .A1(n8538), .A2(n8197), .B1(n6547), .B2(P2_U3152), .C1(
        n8196), .C2(n4858), .ZN(P2_U3330) );
  NAND2_X1 U9376 ( .A1(n8203), .A2(n8234), .ZN(n8199) );
  NAND2_X1 U9377 ( .A1(n9042), .A2(n9892), .ZN(n8198) );
  NAND2_X1 U9378 ( .A1(n8199), .A2(n8198), .ZN(n8200) );
  XNOR2_X1 U9379 ( .A(n8200), .B(n9017), .ZN(n8213) );
  INV_X1 U9380 ( .A(n8213), .ZN(n8205) );
  NOR2_X1 U9381 ( .A1(n8201), .A2(n9019), .ZN(n8202) );
  AOI21_X1 U9382 ( .B1(n8203), .B2(n9042), .A(n8202), .ZN(n8212) );
  INV_X1 U9383 ( .A(n8212), .ZN(n8204) );
  NAND2_X1 U9384 ( .A1(n8205), .A2(n8204), .ZN(n8833) );
  INV_X1 U9385 ( .A(n8833), .ZN(n8218) );
  INV_X1 U9386 ( .A(n8206), .ZN(n8211) );
  NAND2_X1 U9387 ( .A1(n8213), .A2(n8212), .ZN(n8215) );
  AOI21_X1 U9388 ( .B1(n8833), .B2(n8215), .A(n8214), .ZN(n8216) );
  NOR2_X1 U9389 ( .A1(n8216), .A2(n9879), .ZN(n8217) );
  OAI21_X1 U9390 ( .B1(n8218), .B2(n8233), .A(n8217), .ZN(n8224) );
  OAI21_X1 U9391 ( .B1(n9871), .B2(n9754), .A(n8219), .ZN(n8222) );
  NOR2_X1 U9392 ( .A1(n9876), .A2(n8220), .ZN(n8221) );
  AOI211_X1 U9393 ( .C1(n9873), .C2(n9893), .A(n8222), .B(n8221), .ZN(n8223)
         );
  OAI211_X1 U9394 ( .C1(n10652), .C2(n9824), .A(n8224), .B(n8223), .ZN(
        P1_U3222) );
  INV_X1 U9395 ( .A(n9700), .ZN(n9429) );
  AOI21_X1 U9396 ( .B1(n8226), .B2(n8225), .A(n10615), .ZN(n8227) );
  NAND2_X1 U9397 ( .A1(n8227), .A2(n8266), .ZN(n8232) );
  NOR2_X1 U9398 ( .A1(n10623), .A2(n9591), .ZN(n8230) );
  OAI21_X1 U9399 ( .B1(n10500), .B2(n9596), .A(n8228), .ZN(n8229) );
  AOI211_X1 U9400 ( .C1(n8984), .C2(n9570), .A(n8230), .B(n8229), .ZN(n8231)
         );
  OAI211_X1 U9401 ( .C1(n9429), .C2(n6546), .A(n8232), .B(n8231), .ZN(P2_U3221) );
  NAND2_X1 U9402 ( .A1(n10261), .A2(n8234), .ZN(n8236) );
  NAND2_X1 U9403 ( .A1(n9042), .A2(n9891), .ZN(n8235) );
  NAND2_X1 U9404 ( .A1(n8236), .A2(n8235), .ZN(n8237) );
  NAND2_X1 U9405 ( .A1(n10261), .A2(n9042), .ZN(n8239) );
  NAND2_X1 U9406 ( .A1(n9046), .A2(n9891), .ZN(n8238) );
  NAND2_X1 U9407 ( .A1(n8239), .A2(n8238), .ZN(n8829) );
  INV_X1 U9408 ( .A(n8829), .ZN(n8843) );
  XNOR2_X1 U9409 ( .A(n8844), .B(n8843), .ZN(n8240) );
  XNOR2_X1 U9410 ( .A(n8845), .B(n8240), .ZN(n8248) );
  OAI21_X1 U9411 ( .B1(n9871), .B2(n8242), .A(n8241), .ZN(n8243) );
  AOI21_X1 U9412 ( .B1(n9873), .B2(n9892), .A(n8243), .ZN(n8244) );
  OAI21_X1 U9413 ( .B1(n9876), .B2(n8245), .A(n8244), .ZN(n8246) );
  AOI21_X1 U9414 ( .B1(n10261), .B2(n9863), .A(n8246), .ZN(n8247) );
  OAI21_X1 U9415 ( .B1(n8248), .B2(n9879), .A(n8247), .ZN(P1_U3232) );
  INV_X1 U9416 ( .A(n8672), .ZN(n8249) );
  XNOR2_X1 U9417 ( .A(n8250), .B(n8249), .ZN(n10238) );
  OAI22_X1 U9418 ( .A1(n9818), .A2(n10111), .B1(n9870), .B2(n10149), .ZN(n8255) );
  INV_X1 U9419 ( .A(n8251), .ZN(n8252) );
  AOI211_X1 U9420 ( .C1(n8672), .C2(n8253), .A(n10107), .B(n8252), .ZN(n8254)
         );
  AOI211_X1 U9421 ( .C1(n10238), .C2(n10604), .A(n8255), .B(n8254), .ZN(n10242) );
  INV_X1 U9422 ( .A(n8256), .ZN(n8258) );
  INV_X1 U9423 ( .A(n10157), .ZN(n8257) );
  AOI21_X1 U9424 ( .B1(n10239), .B2(n8258), .A(n8257), .ZN(n10240) );
  NOR2_X1 U9425 ( .A1(n9825), .A2(n10130), .ZN(n8261) );
  INV_X1 U9426 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8259) );
  OAI22_X1 U9427 ( .A1(n10163), .A2(n8259), .B1(n9819), .B2(n10160), .ZN(n8260) );
  AOI211_X1 U9428 ( .C1(n10240), .C2(n10137), .A(n8261), .B(n8260), .ZN(n8263)
         );
  NAND2_X1 U9429 ( .A1(n10238), .A2(n10169), .ZN(n8262) );
  OAI211_X1 U9430 ( .C1(n10242), .C2(n4856), .A(n8263), .B(n8262), .ZN(
        P1_U3274) );
  INV_X1 U9431 ( .A(n8305), .ZN(n9063) );
  INV_X1 U9432 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8306) );
  OAI222_X1 U9433 ( .A1(n8538), .A2(n9063), .B1(n6035), .B2(P2_U3152), .C1(
        n8306), .C2(n4858), .ZN(P2_U3329) );
  INV_X1 U9434 ( .A(n9692), .ZN(n9581) );
  INV_X1 U9435 ( .A(n8264), .ZN(n8265) );
  AOI21_X1 U9436 ( .B1(n8266), .B2(n8265), .A(n10615), .ZN(n8270) );
  NOR3_X1 U9437 ( .A1(n8267), .A2(n9428), .A3(n9129), .ZN(n8269) );
  OAI21_X1 U9438 ( .B1(n8270), .B2(n8269), .A(n8268), .ZN(n8275) );
  INV_X1 U9439 ( .A(n8271), .ZN(n9579) );
  INV_X1 U9440 ( .A(n9584), .ZN(n9557) );
  AOI22_X1 U9441 ( .A1(n10609), .A2(n9627), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8272) );
  OAI21_X1 U9442 ( .B1(n9557), .B2(n10611), .A(n8272), .ZN(n8273) );
  AOI21_X1 U9443 ( .B1(n9579), .B2(n9121), .A(n8273), .ZN(n8274) );
  OAI211_X1 U9444 ( .C1(n9581), .C2(n6546), .A(n8275), .B(n8274), .ZN(P2_U3235) );
  MUX2_X1 U9445 ( .A(n8276), .B(P1_REG2_REG_8__SCAN_IN), .S(n4856), .Z(n8285)
         );
  OAI22_X1 U9446 ( .A1(n5182), .A2(n10130), .B1(n10160), .B2(n8278), .ZN(n8279) );
  AOI21_X1 U9447 ( .B1(n8280), .B2(n10137), .A(n8279), .ZN(n8281) );
  OAI21_X1 U9448 ( .B1(n8283), .B2(n8282), .A(n8281), .ZN(n8284) );
  OR2_X1 U9449 ( .A1(n8285), .A2(n8284), .ZN(P1_U3283) );
  INV_X1 U9450 ( .A(n8288), .ZN(n8289) );
  NAND2_X1 U9451 ( .A1(n8289), .A2(n9260), .ZN(n8290) );
  MUX2_X1 U9452 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n8295), .Z(n8293) );
  INV_X1 U9453 ( .A(SI_30_), .ZN(n9258) );
  XNOR2_X1 U9454 ( .A(n8293), .B(n9258), .ZN(n8291) );
  INV_X1 U9455 ( .A(n8542), .ZN(n8998) );
  INV_X1 U9456 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8543) );
  OAI222_X1 U9457 ( .A1(n9064), .A2(n8998), .B1(n5336), .B2(P1_U3084), .C1(
        n8543), .C2(n9060), .ZN(P1_U3323) );
  INV_X1 U9458 ( .A(n8293), .ZN(n8294) );
  MUX2_X1 U9459 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n8295), .Z(n8297) );
  INV_X1 U9460 ( .A(SI_31_), .ZN(n8296) );
  XNOR2_X1 U9461 ( .A(n8297), .B(n8296), .ZN(n8298) );
  NAND2_X1 U9462 ( .A1(n10290), .A2(n8304), .ZN(n8301) );
  OR2_X1 U9463 ( .A1(n6366), .A2(n6630), .ZN(n8300) );
  NAND2_X1 U9464 ( .A1(n8542), .A2(n8304), .ZN(n8303) );
  INV_X1 U9465 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8996) );
  OR2_X1 U9466 ( .A1(n6366), .A2(n8996), .ZN(n8302) );
  NAND2_X1 U9467 ( .A1(n8305), .A2(n8304), .ZN(n8308) );
  OR2_X1 U9468 ( .A1(n6366), .A2(n8306), .ZN(n8307) );
  INV_X1 U9469 ( .A(n9650), .ZN(n9464) );
  INV_X1 U9470 ( .A(n9655), .ZN(n9476) );
  INV_X1 U9471 ( .A(n9676), .ZN(n9546) );
  INV_X1 U9472 ( .A(n9682), .ZN(n9554) );
  INV_X1 U9473 ( .A(n9703), .ZN(n9621) );
  INV_X1 U9474 ( .A(n8486), .ZN(n8337) );
  OAI21_X1 U9475 ( .B1(n7063), .B2(n8311), .A(n9626), .ZN(n9445) );
  NOR2_X1 U9476 ( .A1(n8337), .A2(n9445), .ZN(n9635) );
  INV_X1 U9477 ( .A(n9635), .ZN(n9641) );
  NOR2_X1 U9478 ( .A1(n9618), .A2(n9641), .ZN(n9424) );
  AOI21_X1 U9479 ( .B1(n9618), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9424), .ZN(
        n8313) );
  NAND2_X1 U9480 ( .A1(n9636), .A2(n9606), .ZN(n8312) );
  OAI211_X1 U9481 ( .C1(n9638), .C2(n9451), .A(n8313), .B(n8312), .ZN(P2_U3265) );
  OAI222_X1 U9482 ( .A1(n4858), .A2(n8315), .B1(n8538), .B2(n8314), .C1(n9601), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U9483 ( .A1(n9703), .A2(n9596), .ZN(n8359) );
  NAND2_X1 U9484 ( .A1(n8358), .A2(n8359), .ZN(n9622) );
  INV_X1 U9485 ( .A(n9622), .ZN(n9610) );
  NAND2_X1 U9486 ( .A1(n9623), .A2(n9610), .ZN(n8317) );
  NAND2_X1 U9487 ( .A1(n8317), .A2(n8358), .ZN(n9593) );
  NAND2_X1 U9488 ( .A1(n9593), .A2(n4974), .ZN(n8318) );
  OR2_X1 U9489 ( .A1(n9700), .A2(n9428), .ZN(n8357) );
  NAND2_X1 U9490 ( .A1(n8318), .A2(n8357), .ZN(n9583) );
  NAND2_X1 U9491 ( .A1(n9692), .A2(n9598), .ZN(n8450) );
  INV_X1 U9492 ( .A(n9582), .ZN(n8319) );
  NAND2_X1 U9493 ( .A1(n9687), .A2(n9557), .ZN(n8320) );
  INV_X1 U9494 ( .A(n9556), .ZN(n8322) );
  NAND2_X1 U9495 ( .A1(n9682), .A2(n9092), .ZN(n8350) );
  NAND2_X1 U9496 ( .A1(n9676), .A2(n9558), .ZN(n9525) );
  NAND2_X1 U9497 ( .A1(n9670), .A2(n9107), .ZN(n8347) );
  INV_X1 U9498 ( .A(n9526), .ZN(n8323) );
  AND2_X1 U9499 ( .A1(n8323), .A2(n9525), .ZN(n9500) );
  NAND2_X1 U9500 ( .A1(n9667), .A2(n9528), .ZN(n8463) );
  INV_X1 U9501 ( .A(n9435), .ZN(n9504) );
  AND2_X1 U9502 ( .A1(n9500), .A2(n9504), .ZN(n8324) );
  INV_X1 U9503 ( .A(n8493), .ZN(n8325) );
  AND2_X1 U9504 ( .A1(n8325), .A2(n9488), .ZN(n8346) );
  INV_X1 U9505 ( .A(n8492), .ZN(n8326) );
  NAND2_X1 U9506 ( .A1(n8327), .A2(n8326), .ZN(n9478) );
  INV_X1 U9507 ( .A(n9478), .ZN(n8329) );
  NAND2_X1 U9508 ( .A1(n9655), .A2(n9142), .ZN(n8471) );
  NAND2_X1 U9509 ( .A1(n9645), .A2(n8330), .ZN(n8480) );
  NAND2_X1 U9510 ( .A1(n9442), .A2(n8480), .ZN(n8331) );
  NOR2_X1 U9511 ( .A1(n9423), .A2(n9444), .ZN(n8341) );
  OAI22_X1 U9512 ( .A1(n8332), .A2(n8341), .B1(n8522), .B2(n8486), .ZN(n8334)
         );
  NAND2_X1 U9513 ( .A1(n8334), .A2(n8333), .ZN(n8336) );
  OR2_X1 U9514 ( .A1(n9636), .A2(n8337), .ZN(n8335) );
  NAND2_X1 U9515 ( .A1(n9423), .A2(n9444), .ZN(n8482) );
  NAND2_X1 U9516 ( .A1(n8336), .A2(n8491), .ZN(n8338) );
  NAND2_X1 U9517 ( .A1(n9636), .A2(n8337), .ZN(n8342) );
  XNOR2_X1 U9518 ( .A(n8528), .B(n8339), .ZN(n8529) );
  INV_X1 U9519 ( .A(n8341), .ZN(n8483) );
  NAND2_X1 U9520 ( .A1(n8342), .A2(n8483), .ZN(n8520) );
  INV_X1 U9521 ( .A(n8463), .ZN(n8344) );
  NOR2_X1 U9522 ( .A1(n8492), .A2(n8344), .ZN(n8345) );
  MUX2_X1 U9523 ( .A(n8346), .B(n8345), .S(n8478), .Z(n8470) );
  AND2_X1 U9524 ( .A1(n8347), .A2(n9525), .ZN(n8349) );
  AND2_X1 U9525 ( .A1(n9501), .A2(n8352), .ZN(n8348) );
  MUX2_X1 U9526 ( .A(n8349), .B(n8348), .S(n8478), .Z(n8462) );
  INV_X1 U9527 ( .A(n8350), .ZN(n8354) );
  NAND2_X1 U9528 ( .A1(n8352), .A2(n8351), .ZN(n8353) );
  MUX2_X1 U9529 ( .A(n8354), .B(n8353), .S(n8485), .Z(n8356) );
  INV_X1 U9530 ( .A(n9525), .ZN(n8355) );
  NOR2_X1 U9531 ( .A1(n8356), .A2(n8355), .ZN(n8460) );
  OAI211_X1 U9532 ( .C1(n9602), .C2(n8358), .A(n8454), .B(n8357), .ZN(n8361)
         );
  OAI22_X1 U9533 ( .A1(n9602), .A2(n8359), .B1(n9429), .B2(n9627), .ZN(n8360)
         );
  MUX2_X1 U9534 ( .A(n8361), .B(n8360), .S(n8485), .Z(n8449) );
  MUX2_X1 U9535 ( .A(n8363), .B(n8362), .S(n8478), .Z(n8447) );
  AND2_X1 U9536 ( .A1(n8366), .A2(n8365), .ZN(n8370) );
  NAND2_X1 U9537 ( .A1(n8370), .A2(n5187), .ZN(n8367) );
  AOI21_X1 U9538 ( .B1(n7621), .B2(n8367), .A(n8478), .ZN(n8369) );
  INV_X1 U9539 ( .A(n8370), .ZN(n8372) );
  NAND3_X1 U9540 ( .A1(n8372), .A2(n8371), .A3(n8478), .ZN(n8373) );
  NAND2_X1 U9541 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  OAI211_X1 U9542 ( .C1(n8377), .C2(n8485), .A(n8376), .B(n8375), .ZN(n8381)
         );
  MUX2_X1 U9543 ( .A(n8379), .B(n8378), .S(n8485), .Z(n8380) );
  NAND3_X1 U9544 ( .A1(n8381), .A2(n7551), .A3(n8380), .ZN(n8387) );
  NAND2_X1 U9545 ( .A1(n8382), .A2(n8478), .ZN(n8384) );
  NAND2_X1 U9546 ( .A1(n10507), .A2(n8485), .ZN(n8383) );
  MUX2_X1 U9547 ( .A(n8384), .B(n8383), .S(n9377), .Z(n8385) );
  NAND3_X1 U9548 ( .A1(n8387), .A2(n8386), .A3(n8385), .ZN(n8391) );
  OR2_X1 U9549 ( .A1(n7566), .A2(n8485), .ZN(n8389) );
  NAND2_X1 U9550 ( .A1(n7566), .A2(n8485), .ZN(n8388) );
  MUX2_X1 U9551 ( .A(n8389), .B(n8388), .S(n9375), .Z(n8390) );
  NAND2_X1 U9552 ( .A1(n8391), .A2(n8390), .ZN(n8396) );
  MUX2_X1 U9553 ( .A(n10536), .B(n10527), .S(n8485), .Z(n8392) );
  OAI21_X1 U9554 ( .B1(n8396), .B2(n8393), .A(n8392), .ZN(n8398) );
  NAND3_X1 U9555 ( .A1(n8396), .A2(n8395), .A3(n8394), .ZN(n8397) );
  NAND2_X1 U9556 ( .A1(n8398), .A2(n8397), .ZN(n8399) );
  NAND2_X1 U9557 ( .A1(n8399), .A2(n8501), .ZN(n8403) );
  MUX2_X1 U9558 ( .A(n8401), .B(n8400), .S(n8478), .Z(n8402) );
  NAND3_X1 U9559 ( .A1(n8403), .A2(n8502), .A3(n8402), .ZN(n8408) );
  MUX2_X1 U9560 ( .A(n8405), .B(n8404), .S(n8485), .Z(n8406) );
  NAND2_X1 U9561 ( .A1(n8415), .A2(n8417), .ZN(n8409) );
  MUX2_X1 U9562 ( .A(n8410), .B(n8409), .S(n8485), .Z(n8412) );
  INV_X1 U9563 ( .A(n8413), .ZN(n8411) );
  NOR2_X1 U9564 ( .A1(n8412), .A2(n8411), .ZN(n8414) );
  NAND2_X1 U9565 ( .A1(n8421), .A2(n8413), .ZN(n8420) );
  INV_X1 U9566 ( .A(n8414), .ZN(n8418) );
  OAI211_X1 U9567 ( .C1(n8418), .C2(n8417), .A(n8416), .B(n8415), .ZN(n8419)
         );
  MUX2_X1 U9568 ( .A(n8420), .B(n8419), .S(n8478), .Z(n8431) );
  INV_X1 U9569 ( .A(n8421), .ZN(n8422) );
  NAND2_X1 U9570 ( .A1(n8426), .A2(n8422), .ZN(n8423) );
  AND2_X1 U9571 ( .A1(n8423), .A2(n8425), .ZN(n8429) );
  NAND2_X1 U9572 ( .A1(n8425), .A2(n8424), .ZN(n8427) );
  AND2_X1 U9573 ( .A1(n8427), .A2(n8426), .ZN(n8428) );
  MUX2_X1 U9574 ( .A(n8429), .B(n8428), .S(n8485), .Z(n8430) );
  MUX2_X1 U9575 ( .A(n8433), .B(n8432), .S(n8478), .Z(n8434) );
  NAND3_X1 U9576 ( .A1(n8435), .A2(n8510), .A3(n8434), .ZN(n8439) );
  MUX2_X1 U9577 ( .A(n8437), .B(n8436), .S(n8478), .Z(n8438) );
  NAND3_X1 U9578 ( .A1(n8512), .A2(n8439), .A3(n8438), .ZN(n8443) );
  MUX2_X1 U9579 ( .A(n8441), .B(n8440), .S(n8485), .Z(n8442) );
  MUX2_X1 U9580 ( .A(n8445), .B(n8444), .S(n8485), .Z(n8446) );
  NOR2_X1 U9581 ( .A1(n8449), .A2(n8448), .ZN(n8451) );
  MUX2_X1 U9582 ( .A(n8478), .B(n8451), .S(n8450), .Z(n8458) );
  MUX2_X1 U9583 ( .A(n9584), .B(n9687), .S(n8478), .Z(n8455) );
  NAND2_X1 U9584 ( .A1(n9687), .A2(n9584), .ZN(n8452) );
  NAND2_X1 U9585 ( .A1(n8455), .A2(n8452), .ZN(n8453) );
  OAI21_X1 U9586 ( .B1(n8478), .B2(n8454), .A(n8453), .ZN(n8457) );
  NOR2_X1 U9587 ( .A1(n9687), .A2(n9584), .ZN(n9430) );
  OR2_X1 U9588 ( .A1(n8455), .A2(n9430), .ZN(n8456) );
  OAI211_X1 U9589 ( .C1(n8458), .C2(n8457), .A(n9431), .B(n8456), .ZN(n8459)
         );
  NAND2_X1 U9590 ( .A1(n8460), .A2(n8459), .ZN(n8461) );
  NAND2_X1 U9591 ( .A1(n8462), .A2(n8461), .ZN(n8464) );
  INV_X1 U9592 ( .A(n9670), .ZN(n9524) );
  AOI21_X1 U9593 ( .B1(n8464), .B2(n9524), .A(n9435), .ZN(n8467) );
  AND2_X1 U9594 ( .A1(n8463), .A2(n8485), .ZN(n8466) );
  OAI211_X1 U9595 ( .C1(n9536), .C2(n8485), .A(n8464), .B(n9501), .ZN(n8465)
         );
  OAI21_X1 U9596 ( .B1(n8467), .B2(n8466), .A(n8465), .ZN(n8469) );
  MUX2_X1 U9597 ( .A(n8492), .B(n8493), .S(n8478), .Z(n8468) );
  AOI21_X1 U9598 ( .B1(n8470), .B2(n8469), .A(n8468), .ZN(n8474) );
  MUX2_X1 U9599 ( .A(n8472), .B(n8471), .S(n8485), .Z(n8473) );
  OAI211_X1 U9600 ( .C1(n8474), .C2(n9477), .A(n9465), .B(n8473), .ZN(n8477)
         );
  OR3_X1 U9601 ( .A1(n9650), .A2(n9480), .A3(n8478), .ZN(n8476) );
  NAND3_X1 U9602 ( .A1(n9650), .A2(n9480), .A3(n8478), .ZN(n8475) );
  NAND4_X1 U9603 ( .A1(n8477), .A2(n9440), .A3(n8476), .A4(n8475), .ZN(n8484)
         );
  MUX2_X1 U9604 ( .A(n8480), .B(n8479), .S(n8478), .Z(n8481) );
  NAND4_X1 U9605 ( .A1(n8484), .A2(n8483), .A3(n8482), .A4(n8481), .ZN(n8489)
         );
  NAND2_X1 U9606 ( .A1(n9636), .A2(n8486), .ZN(n8488) );
  MUX2_X1 U9607 ( .A(n9636), .B(n8486), .S(n8485), .Z(n8487) );
  INV_X1 U9608 ( .A(n8491), .ZN(n8519) );
  NAND4_X1 U9609 ( .A1(n6953), .A2(n8524), .A3(n10463), .A4(n8494), .ZN(n8498)
         );
  NOR4_X1 U9610 ( .A1(n8498), .A2(n8497), .A3(n8496), .A4(n8495), .ZN(n8500)
         );
  NAND4_X1 U9611 ( .A1(n8502), .A2(n8501), .A3(n8500), .A4(n8499), .ZN(n8503)
         );
  NOR4_X1 U9612 ( .A1(n8506), .A2(n8505), .A3(n8504), .A4(n8503), .ZN(n8507)
         );
  AND4_X1 U9613 ( .A1(n8510), .A2(n8509), .A3(n8508), .A4(n8507), .ZN(n8511)
         );
  NAND4_X1 U9614 ( .A1(n5080), .A2(n8513), .A3(n8512), .A4(n8511), .ZN(n8514)
         );
  NOR4_X1 U9615 ( .A1(n9582), .A2(n9602), .A3(n9622), .A4(n8514), .ZN(n8515)
         );
  XNOR2_X1 U9616 ( .A(n9687), .B(n9584), .ZN(n9568) );
  NAND4_X1 U9617 ( .A1(n9538), .A2(n9431), .A3(n8515), .A4(n9568), .ZN(n8516)
         );
  NOR3_X1 U9618 ( .A1(n9435), .A2(n9526), .A3(n8516), .ZN(n8517) );
  NAND4_X1 U9619 ( .A1(n9440), .A2(n8328), .A3(n9490), .A4(n8517), .ZN(n8518)
         );
  XNOR2_X1 U9620 ( .A(n8521), .B(n9601), .ZN(n8523) );
  OAI211_X1 U9621 ( .C1(n8525), .C2(n8524), .A(n8523), .B(n8522), .ZN(n8526)
         );
  INV_X1 U9622 ( .A(n10299), .ZN(n8531) );
  NOR4_X1 U9623 ( .A1(n8531), .A2(n8530), .A3(n7063), .A4(n9597), .ZN(n8534)
         );
  OAI21_X1 U9624 ( .B1(n8535), .B2(n8532), .A(P2_B_REG_SCAN_IN), .ZN(n8533) );
  INV_X1 U9625 ( .A(n8536), .ZN(n9040) );
  OAI222_X1 U9626 ( .A1(n4858), .A2(n8539), .B1(n8538), .B2(n9040), .C1(n8537), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9627 ( .A(n8631), .ZN(n8639) );
  NOR2_X1 U9628 ( .A1(n8544), .A2(n6694), .ZN(n8540) );
  NAND2_X1 U9629 ( .A1(n8542), .A2(n8541), .ZN(n8546) );
  OR2_X1 U9630 ( .A1(n8544), .A2(n8543), .ZN(n8545) );
  INV_X1 U9631 ( .A(n9881), .ZN(n8647) );
  OR2_X1 U9632 ( .A1(n10176), .A2(n8647), .ZN(n8648) );
  MUX2_X1 U9633 ( .A(n8758), .B(n8756), .S(n8631), .Z(n8625) );
  MUX2_X1 U9634 ( .A(n8753), .B(n8751), .S(n8631), .Z(n8623) );
  MUX2_X1 U9635 ( .A(n8750), .B(n8748), .S(n8631), .Z(n8621) );
  INV_X1 U9636 ( .A(n7102), .ZN(n8548) );
  INV_X1 U9637 ( .A(n8714), .ZN(n8547) );
  AOI21_X1 U9638 ( .B1(n8548), .B2(n8788), .A(n8547), .ZN(n8549) );
  MUX2_X1 U9639 ( .A(n8550), .B(n8549), .S(n8631), .Z(n8554) );
  NAND2_X1 U9640 ( .A1(n8791), .A2(n8551), .ZN(n8716) );
  NAND2_X1 U9641 ( .A1(n8709), .A2(n8789), .ZN(n8552) );
  MUX2_X1 U9642 ( .A(n8716), .B(n8552), .S(n8631), .Z(n8553) );
  AOI21_X1 U9643 ( .B1(n8554), .B2(n8655), .A(n8553), .ZN(n8560) );
  MUX2_X1 U9644 ( .A(n8709), .B(n8791), .S(n8631), .Z(n8555) );
  NAND2_X1 U9645 ( .A1(n8556), .A2(n8555), .ZN(n8559) );
  MUX2_X1 U9646 ( .A(n8557), .B(n8708), .S(n8631), .Z(n8558) );
  OAI211_X1 U9647 ( .C1(n8560), .C2(n8559), .A(n8657), .B(n8558), .ZN(n8563)
         );
  MUX2_X1 U9648 ( .A(n8721), .B(n8561), .S(n8631), .Z(n8562) );
  NAND3_X1 U9649 ( .A1(n8563), .A2(n8664), .A3(n8562), .ZN(n8565) );
  MUX2_X1 U9650 ( .A(n8723), .B(n8720), .S(n8631), .Z(n8564) );
  NAND3_X1 U9651 ( .A1(n8565), .A2(n8663), .A3(n8564), .ZN(n8567) );
  MUX2_X1 U9652 ( .A(n8725), .B(n8728), .S(n8631), .Z(n8566) );
  NAND3_X1 U9653 ( .A1(n8567), .A2(n8665), .A3(n8566), .ZN(n8569) );
  AOI21_X1 U9654 ( .B1(n8569), .B2(n8729), .A(n8568), .ZN(n8571) );
  INV_X1 U9655 ( .A(n8730), .ZN(n8581) );
  AOI21_X1 U9656 ( .B1(n8569), .B2(n8706), .A(n8581), .ZN(n8570) );
  MUX2_X1 U9657 ( .A(n8571), .B(n8570), .S(n8631), .Z(n8572) );
  NOR2_X1 U9658 ( .A1(n8572), .A2(n8667), .ZN(n8594) );
  NAND4_X1 U9659 ( .A1(n8702), .A2(n8639), .A3(n8735), .A4(n8736), .ZN(n8592)
         );
  NOR2_X1 U9660 ( .A1(n8639), .A2(n9889), .ZN(n8573) );
  NAND2_X1 U9661 ( .A1(n10249), .A2(n8573), .ZN(n8580) );
  OAI21_X1 U9662 ( .B1(n8639), .B2(n9888), .A(n8580), .ZN(n8590) );
  AND2_X1 U9663 ( .A1(n8639), .A2(n9888), .ZN(n8585) );
  INV_X1 U9664 ( .A(n8585), .ZN(n8574) );
  AOI21_X1 U9665 ( .B1(n8730), .B2(n8853), .A(n8574), .ZN(n8575) );
  OAI211_X1 U9666 ( .C1(n9889), .C2(n8735), .A(n8576), .B(n8575), .ZN(n8579)
         );
  NAND2_X1 U9667 ( .A1(n8639), .A2(n9889), .ZN(n8583) );
  INV_X1 U9668 ( .A(n8583), .ZN(n8577) );
  NAND4_X1 U9669 ( .A1(n8735), .A2(n8581), .A3(n8577), .A4(n9888), .ZN(n8578)
         );
  OAI211_X1 U9670 ( .C1(n8580), .C2(n9888), .A(n8579), .B(n8578), .ZN(n8589)
         );
  NOR2_X1 U9671 ( .A1(n8730), .A2(n8583), .ZN(n8586) );
  NAND3_X1 U9672 ( .A1(n8735), .A2(n8639), .A3(n8581), .ZN(n8582) );
  AOI21_X1 U9673 ( .B1(n8583), .B2(n8582), .A(n10249), .ZN(n8584) );
  AOI211_X1 U9674 ( .C1(n8586), .C2(n8735), .A(n8585), .B(n8584), .ZN(n8587)
         );
  NOR2_X1 U9675 ( .A1(n8587), .A2(n10246), .ZN(n8588) );
  AOI211_X1 U9676 ( .C1(n10246), .C2(n8590), .A(n8589), .B(n8588), .ZN(n8591)
         );
  OAI21_X1 U9677 ( .B1(n8594), .B2(n8592), .A(n8591), .ZN(n8596) );
  NAND4_X1 U9678 ( .A1(n8739), .A2(n8631), .A3(n8731), .A4(n8738), .ZN(n8593)
         );
  AOI21_X1 U9679 ( .B1(n8594), .B2(n8707), .A(n8593), .ZN(n8595) );
  NOR2_X1 U9680 ( .A1(n8596), .A2(n8595), .ZN(n8598) );
  MUX2_X1 U9681 ( .A(n8687), .B(n8703), .S(n8631), .Z(n8597) );
  OAI211_X1 U9682 ( .C1(n8598), .C2(n8672), .A(n10139), .B(n8597), .ZN(n8601)
         );
  INV_X1 U9683 ( .A(n10132), .ZN(n8600) );
  MUX2_X1 U9684 ( .A(n8705), .B(n8688), .S(n8631), .Z(n8599) );
  NAND3_X1 U9685 ( .A1(n8601), .A2(n8600), .A3(n8599), .ZN(n8603) );
  MUX2_X1 U9686 ( .A(n8691), .B(n8699), .S(n8631), .Z(n8602) );
  NAND2_X1 U9687 ( .A1(n8603), .A2(n8602), .ZN(n8611) );
  NOR2_X1 U9688 ( .A1(n10088), .A2(n10109), .ZN(n8675) );
  AND2_X1 U9689 ( .A1(n8694), .A2(n8607), .ZN(n8609) );
  INV_X1 U9690 ( .A(n8604), .ZN(n8605) );
  NAND2_X1 U9691 ( .A1(n8606), .A2(n8605), .ZN(n8608) );
  NAND2_X1 U9692 ( .A1(n8608), .A2(n8607), .ZN(n8684) );
  MUX2_X1 U9693 ( .A(n8609), .B(n8684), .S(n8631), .Z(n8610) );
  NAND2_X1 U9694 ( .A1(n4896), .A2(n8612), .ZN(n10063) );
  MUX2_X1 U9695 ( .A(n8685), .B(n8695), .S(n8631), .Z(n8613) );
  NAND2_X1 U9696 ( .A1(n10063), .A2(n8613), .ZN(n8616) );
  INV_X1 U9697 ( .A(n8744), .ZN(n8614) );
  MUX2_X1 U9698 ( .A(n10032), .B(n8614), .S(n8631), .Z(n8615) );
  OAI211_X1 U9699 ( .C1(n8617), .C2(n8616), .A(n10035), .B(n8615), .ZN(n8619)
         );
  MUX2_X1 U9700 ( .A(n8747), .B(n8745), .S(n8631), .Z(n8618) );
  NAND3_X1 U9701 ( .A1(n10015), .A2(n8619), .A3(n8618), .ZN(n8620) );
  NAND3_X1 U9702 ( .A1(n9995), .A2(n8621), .A3(n8620), .ZN(n8622) );
  NAND3_X1 U9703 ( .A1(n8678), .A2(n8623), .A3(n8622), .ZN(n8624) );
  AND3_X1 U9704 ( .A1(n9965), .A2(n8625), .A3(n8624), .ZN(n8630) );
  INV_X1 U9705 ( .A(n8630), .ZN(n8626) );
  NAND3_X1 U9706 ( .A1(n8626), .A2(n8810), .A3(n8757), .ZN(n8627) );
  NAND2_X1 U9707 ( .A1(n8627), .A2(n8629), .ZN(n8633) );
  NAND2_X1 U9708 ( .A1(n8629), .A2(n8628), .ZN(n8805) );
  OAI21_X1 U9709 ( .B1(n8630), .B2(n8805), .A(n8810), .ZN(n8632) );
  MUX2_X1 U9710 ( .A(n8633), .B(n8632), .S(n8631), .Z(n8634) );
  OAI21_X1 U9711 ( .B1(n9952), .B2(n8648), .A(n8634), .ZN(n8636) );
  NAND2_X1 U9712 ( .A1(n9947), .A2(n9881), .ZN(n8635) );
  NAND2_X1 U9713 ( .A1(n10176), .A2(n8635), .ZN(n8760) );
  INV_X1 U9714 ( .A(n9952), .ZN(n10172) );
  INV_X1 U9715 ( .A(n9947), .ZN(n8638) );
  OR2_X1 U9716 ( .A1(n10172), .A2(n8638), .ZN(n8640) );
  AND2_X1 U9717 ( .A1(n10172), .A2(n8638), .ZN(n8681) );
  AOI21_X1 U9718 ( .B1(n8637), .B2(n8640), .A(n8681), .ZN(n8646) );
  INV_X1 U9719 ( .A(n8646), .ZN(n8644) );
  INV_X1 U9720 ( .A(n8681), .ZN(n8813) );
  OAI21_X1 U9721 ( .B1(n8648), .B2(n8638), .A(n8813), .ZN(n8683) );
  NAND2_X1 U9722 ( .A1(n8683), .A2(n8639), .ZN(n8643) );
  INV_X1 U9723 ( .A(n8640), .ZN(n8763) );
  NAND2_X1 U9724 ( .A1(n5958), .A2(n9041), .ZN(n8641) );
  NOR3_X1 U9725 ( .A1(n8646), .A2(n9944), .A3(n8645), .ZN(n8771) );
  AOI21_X1 U9726 ( .B1(n8647), .B2(n10176), .A(n8763), .ZN(n8812) );
  INV_X1 U9727 ( .A(n8648), .ZN(n8809) );
  INV_X1 U9728 ( .A(n10076), .ZN(n8674) );
  NOR4_X1 U9729 ( .A1(n5910), .A2(n8652), .A3(n8651), .A4(n8650), .ZN(n8654)
         );
  NAND4_X1 U9730 ( .A1(n8656), .A2(n8655), .A3(n8654), .A4(n8653), .ZN(n8661)
         );
  INV_X1 U9731 ( .A(n8657), .ZN(n8660) );
  NOR4_X1 U9732 ( .A1(n8661), .A2(n8660), .A3(n8659), .A4(n8658), .ZN(n8662)
         );
  NAND4_X1 U9733 ( .A1(n8665), .A2(n8664), .A3(n8663), .A4(n8662), .ZN(n8666)
         );
  NOR4_X1 U9734 ( .A1(n8668), .A2(n8667), .A3(n5934), .A4(n8666), .ZN(n8670)
         );
  NAND2_X1 U9735 ( .A1(n8670), .A2(n8669), .ZN(n8671) );
  NOR4_X1 U9736 ( .A1(n10132), .A2(n10143), .A3(n8672), .A4(n8671), .ZN(n8673)
         );
  NAND4_X1 U9737 ( .A1(n10063), .A2(n8675), .A3(n8674), .A4(n8673), .ZN(n8676)
         );
  NOR3_X1 U9738 ( .A1(n10024), .A2(n5952), .A3(n8676), .ZN(n8677) );
  NAND4_X1 U9739 ( .A1(n9965), .A2(n8678), .A3(n9995), .A4(n8677), .ZN(n8679)
         );
  NOR4_X1 U9740 ( .A1(n8681), .A2(n8809), .A3(n8680), .A4(n8679), .ZN(n8682)
         );
  AOI21_X1 U9741 ( .B1(n8812), .B2(n8682), .A(n5958), .ZN(n8767) );
  INV_X1 U9742 ( .A(n8683), .ZN(n8765) );
  INV_X1 U9743 ( .A(n8684), .ZN(n8686) );
  NAND2_X1 U9744 ( .A1(n8686), .A2(n8685), .ZN(n8701) );
  NAND2_X1 U9745 ( .A1(n8688), .A2(n8687), .ZN(n8689) );
  NAND2_X1 U9746 ( .A1(n8689), .A2(n8705), .ZN(n8690) );
  NAND2_X1 U9747 ( .A1(n8691), .A2(n8690), .ZN(n8692) );
  AND2_X1 U9748 ( .A1(n8692), .A2(n8699), .ZN(n8693) );
  NOR2_X1 U9749 ( .A1(n8694), .A2(n8693), .ZN(n8696) );
  OAI21_X1 U9750 ( .B1(n8701), .B2(n8696), .A(n8695), .ZN(n8697) );
  NOR2_X1 U9751 ( .A1(n8698), .A2(n8697), .ZN(n8799) );
  INV_X1 U9752 ( .A(n8699), .ZN(n8700) );
  NOR2_X1 U9753 ( .A1(n8701), .A2(n8700), .ZN(n8798) );
  AND2_X1 U9754 ( .A1(n8703), .A2(n8702), .ZN(n8704) );
  NAND2_X1 U9755 ( .A1(n8705), .A2(n8704), .ZN(n8741) );
  INV_X1 U9756 ( .A(n8736), .ZN(n8713) );
  NAND2_X1 U9757 ( .A1(n8707), .A2(n8706), .ZN(n8733) );
  INV_X1 U9758 ( .A(n8733), .ZN(n8711) );
  AND4_X1 U9759 ( .A1(n8720), .A2(n8709), .A3(n8708), .A4(n8721), .ZN(n8710)
         );
  NAND4_X1 U9760 ( .A1(n8735), .A2(n8711), .A3(n8710), .A4(n8725), .ZN(n8712)
         );
  OR3_X1 U9761 ( .A1(n8741), .A2(n8713), .A3(n8712), .ZN(n8774) );
  NAND2_X1 U9762 ( .A1(n7102), .A2(n8714), .ZN(n8718) );
  INV_X1 U9763 ( .A(n8715), .ZN(n8717) );
  AOI21_X1 U9764 ( .B1(n8718), .B2(n8717), .A(n8716), .ZN(n8742) );
  INV_X1 U9765 ( .A(n8719), .ZN(n8722) );
  NAND3_X1 U9766 ( .A1(n8722), .A2(n8721), .A3(n8720), .ZN(n8724) );
  NAND2_X1 U9767 ( .A1(n8724), .A2(n8723), .ZN(n8726) );
  NAND2_X1 U9768 ( .A1(n8726), .A2(n8725), .ZN(n8727) );
  AND3_X1 U9769 ( .A1(n8729), .A2(n8728), .A3(n8727), .ZN(n8732) );
  OAI211_X1 U9770 ( .C1(n8733), .C2(n8732), .A(n8731), .B(n8730), .ZN(n8734)
         );
  NAND3_X1 U9771 ( .A1(n8736), .A2(n8735), .A3(n8734), .ZN(n8737) );
  AND3_X1 U9772 ( .A1(n8739), .A2(n8738), .A3(n8737), .ZN(n8740) );
  OR2_X1 U9773 ( .A1(n8741), .A2(n8740), .ZN(n8794) );
  OAI21_X1 U9774 ( .B1(n8774), .B2(n8742), .A(n8794), .ZN(n8743) );
  NAND2_X1 U9775 ( .A1(n8798), .A2(n8743), .ZN(n8749) );
  NAND2_X1 U9776 ( .A1(n8745), .A2(n8744), .ZN(n8746) );
  NAND3_X1 U9777 ( .A1(n8748), .A2(n8747), .A3(n8746), .ZN(n8773) );
  AOI21_X1 U9778 ( .B1(n8799), .B2(n8749), .A(n8773), .ZN(n8752) );
  NAND2_X1 U9779 ( .A1(n8751), .A2(n8750), .ZN(n8802) );
  NOR2_X1 U9780 ( .A1(n8752), .A2(n8802), .ZN(n8759) );
  INV_X1 U9781 ( .A(n8753), .ZN(n8754) );
  NAND2_X1 U9782 ( .A1(n8758), .A2(n8754), .ZN(n8755) );
  NAND3_X1 U9783 ( .A1(n8757), .A2(n8756), .A3(n8755), .ZN(n8807) );
  AOI21_X1 U9784 ( .B1(n8759), .B2(n8758), .A(n8807), .ZN(n8761) );
  OAI211_X1 U9785 ( .C1(n8761), .C2(n8805), .A(n8810), .B(n8760), .ZN(n8764)
         );
  AOI211_X1 U9786 ( .C1(n8765), .C2(n8764), .A(n8763), .B(n8762), .ZN(n8766)
         );
  NOR3_X1 U9787 ( .A1(n8767), .A2(n8766), .A3(n10095), .ZN(n8770) );
  INV_X1 U9788 ( .A(n8767), .ZN(n8768) );
  OAI21_X1 U9789 ( .B1(n8768), .B2(n9944), .A(n8816), .ZN(n8769) );
  NOR4_X1 U9790 ( .A1(n8772), .A2(n8771), .A3(n8770), .A4(n8769), .ZN(n8828)
         );
  INV_X1 U9791 ( .A(n8773), .ZN(n8804) );
  INV_X1 U9792 ( .A(n8774), .ZN(n8797) );
  INV_X1 U9793 ( .A(n6902), .ZN(n8777) );
  OAI211_X1 U9794 ( .C1(n8777), .C2(n8776), .A(n5958), .B(n8775), .ZN(n8779)
         );
  NAND2_X1 U9795 ( .A1(n8779), .A2(n8778), .ZN(n8781) );
  OAI21_X1 U9796 ( .B1(n8782), .B2(n8781), .A(n8780), .ZN(n8786) );
  INV_X1 U9797 ( .A(n8783), .ZN(n8784) );
  AOI21_X1 U9798 ( .B1(n8786), .B2(n8785), .A(n8784), .ZN(n8793) );
  NAND3_X1 U9799 ( .A1(n8789), .A2(n8788), .A3(n8787), .ZN(n8792) );
  OAI211_X1 U9800 ( .C1(n8793), .C2(n8792), .A(n8791), .B(n8790), .ZN(n8796)
         );
  INV_X1 U9801 ( .A(n8794), .ZN(n8795) );
  AOI21_X1 U9802 ( .B1(n8797), .B2(n8796), .A(n8795), .ZN(n8801) );
  INV_X1 U9803 ( .A(n8798), .ZN(n8800) );
  OAI21_X1 U9804 ( .B1(n8801), .B2(n8800), .A(n8799), .ZN(n8803) );
  AOI211_X1 U9805 ( .C1(n8804), .C2(n8803), .A(n8802), .B(n9986), .ZN(n8808)
         );
  INV_X1 U9806 ( .A(n8805), .ZN(n8806) );
  OAI21_X1 U9807 ( .B1(n8808), .B2(n8807), .A(n8806), .ZN(n8811) );
  AOI21_X1 U9808 ( .B1(n8811), .B2(n8810), .A(n8809), .ZN(n8815) );
  INV_X1 U9809 ( .A(n8812), .ZN(n8814) );
  OAI21_X1 U9810 ( .B1(n8815), .B2(n8814), .A(n8813), .ZN(n8818) );
  NOR3_X1 U9811 ( .A1(n8818), .A2(n8816), .A3(n9944), .ZN(n8817) );
  AOI211_X1 U9812 ( .C1(n8819), .C2(n8818), .A(n8824), .B(n8817), .ZN(n8820)
         );
  INV_X1 U9813 ( .A(n8820), .ZN(n8827) );
  NAND2_X1 U9814 ( .A1(n8822), .A2(n8821), .ZN(n8823) );
  OAI211_X1 U9815 ( .C1(n8825), .C2(n8824), .A(n8823), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8826) );
  OAI21_X1 U9816 ( .B1(n8828), .B2(n8827), .A(n8826), .ZN(P1_U3240) );
  NAND2_X1 U9817 ( .A1(n8847), .A2(n8829), .ZN(n8840) );
  NAND2_X1 U9818 ( .A1(n10257), .A2(n8234), .ZN(n8831) );
  NAND2_X1 U9819 ( .A1(n9042), .A2(n9890), .ZN(n8830) );
  NAND2_X1 U9820 ( .A1(n8831), .A2(n8830), .ZN(n8832) );
  XNOR2_X1 U9821 ( .A(n8832), .B(n9017), .ZN(n8835) );
  AND2_X1 U9822 ( .A1(n8833), .A2(n8835), .ZN(n8834) );
  NAND2_X1 U9823 ( .A1(n8233), .A2(n8834), .ZN(n8838) );
  INV_X1 U9824 ( .A(n8835), .ZN(n8846) );
  INV_X1 U9825 ( .A(n8844), .ZN(n8836) );
  OR2_X1 U9826 ( .A1(n8846), .A2(n8836), .ZN(n8837) );
  NAND2_X1 U9827 ( .A1(n8838), .A2(n8837), .ZN(n8839) );
  NAND2_X1 U9828 ( .A1(n8840), .A2(n8839), .ZN(n9746) );
  NAND2_X1 U9829 ( .A1(n10257), .A2(n9042), .ZN(n8842) );
  NAND2_X1 U9830 ( .A1(n9046), .A2(n9890), .ZN(n8841) );
  NAND2_X1 U9831 ( .A1(n8842), .A2(n8841), .ZN(n9749) );
  NAND2_X1 U9832 ( .A1(n9746), .A2(n9749), .ZN(n8849) );
  NAND3_X1 U9833 ( .A1(n8848), .A2(n8847), .A3(n8846), .ZN(n9747) );
  NAND2_X1 U9834 ( .A1(n8849), .A2(n9747), .ZN(n9865) );
  NAND2_X1 U9835 ( .A1(n10249), .A2(n8234), .ZN(n8851) );
  NAND2_X1 U9836 ( .A1(n9042), .A2(n9889), .ZN(n8850) );
  NAND2_X1 U9837 ( .A1(n8851), .A2(n8850), .ZN(n8852) );
  XNOR2_X1 U9838 ( .A(n8852), .B(n9017), .ZN(n9867) );
  NOR2_X1 U9839 ( .A1(n8853), .A2(n9019), .ZN(n8854) );
  AOI21_X1 U9840 ( .B1(n10249), .B2(n9042), .A(n8854), .ZN(n8856) );
  NAND2_X1 U9841 ( .A1(n9867), .A2(n8856), .ZN(n8855) );
  INV_X1 U9842 ( .A(n9867), .ZN(n8857) );
  INV_X1 U9843 ( .A(n8856), .ZN(n9866) );
  NAND2_X1 U9844 ( .A1(n8857), .A2(n9866), .ZN(n8858) );
  NAND2_X1 U9845 ( .A1(n10246), .A2(n8234), .ZN(n8860) );
  NAND2_X1 U9846 ( .A1(n9042), .A2(n9888), .ZN(n8859) );
  NAND2_X1 U9847 ( .A1(n8860), .A2(n8859), .ZN(n8861) );
  XNOR2_X1 U9848 ( .A(n8861), .B(n9017), .ZN(n8863) );
  NOR2_X1 U9849 ( .A1(n9870), .A2(n9019), .ZN(n8862) );
  AOI21_X1 U9850 ( .B1(n10246), .B2(n9042), .A(n8862), .ZN(n8864) );
  NAND2_X1 U9851 ( .A1(n8863), .A2(n8864), .ZN(n8869) );
  INV_X1 U9852 ( .A(n8863), .ZN(n8866) );
  INV_X1 U9853 ( .A(n8864), .ZN(n8865) );
  NAND2_X1 U9854 ( .A1(n8866), .A2(n8865), .ZN(n8867) );
  NAND2_X1 U9855 ( .A1(n8869), .A2(n8867), .ZN(n9799) );
  NAND2_X1 U9856 ( .A1(n9797), .A2(n8869), .ZN(n9812) );
  NAND2_X1 U9857 ( .A1(n10239), .A2(n8234), .ZN(n8871) );
  NAND2_X1 U9858 ( .A1(n9887), .A2(n9042), .ZN(n8870) );
  NAND2_X1 U9859 ( .A1(n8871), .A2(n8870), .ZN(n8872) );
  XNOR2_X1 U9860 ( .A(n8872), .B(n8946), .ZN(n8875) );
  NAND2_X1 U9861 ( .A1(n10239), .A2(n9042), .ZN(n8874) );
  NAND2_X1 U9862 ( .A1(n9046), .A2(n9887), .ZN(n8873) );
  NAND2_X1 U9863 ( .A1(n8874), .A2(n8873), .ZN(n8876) );
  NAND2_X1 U9864 ( .A1(n8875), .A2(n8876), .ZN(n9813) );
  NAND2_X1 U9865 ( .A1(n9812), .A2(n9813), .ZN(n9810) );
  INV_X1 U9866 ( .A(n8875), .ZN(n8878) );
  INV_X1 U9867 ( .A(n8876), .ZN(n8877) );
  NAND2_X1 U9868 ( .A1(n8878), .A2(n8877), .ZN(n9814) );
  NAND2_X1 U9869 ( .A1(n9810), .A2(n9814), .ZN(n8884) );
  NAND2_X1 U9870 ( .A1(n10231), .A2(n8234), .ZN(n8880) );
  NAND2_X1 U9871 ( .A1(n10121), .A2(n9042), .ZN(n8879) );
  NAND2_X1 U9872 ( .A1(n8880), .A2(n8879), .ZN(n8881) );
  XNOR2_X1 U9873 ( .A(n8881), .B(n9017), .ZN(n8885) );
  NAND2_X1 U9874 ( .A1(n10231), .A2(n9042), .ZN(n8883) );
  NAND2_X1 U9875 ( .A1(n10121), .A2(n9046), .ZN(n8882) );
  NAND2_X1 U9876 ( .A1(n8883), .A2(n8882), .ZN(n9856) );
  NAND2_X1 U9877 ( .A1(n10226), .A2(n8234), .ZN(n8888) );
  NAND2_X1 U9878 ( .A1(n10147), .A2(n9042), .ZN(n8887) );
  NAND2_X1 U9879 ( .A1(n8888), .A2(n8887), .ZN(n8889) );
  XNOR2_X1 U9880 ( .A(n8889), .B(n8946), .ZN(n9767) );
  NAND2_X1 U9881 ( .A1(n10226), .A2(n9042), .ZN(n8891) );
  NAND2_X1 U9882 ( .A1(n10147), .A2(n9046), .ZN(n8890) );
  NAND2_X1 U9883 ( .A1(n8891), .A2(n8890), .ZN(n9768) );
  NAND2_X1 U9884 ( .A1(n10222), .A2(n8234), .ZN(n8893) );
  NAND2_X1 U9885 ( .A1(n10122), .A2(n9042), .ZN(n8892) );
  NAND2_X1 U9886 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  XNOR2_X1 U9887 ( .A(n8894), .B(n9017), .ZN(n8896) );
  AND2_X1 U9888 ( .A1(n10122), .A2(n9046), .ZN(n8895) );
  AOI21_X1 U9889 ( .B1(n10222), .B2(n9042), .A(n8895), .ZN(n8897) );
  NAND2_X1 U9890 ( .A1(n8896), .A2(n8897), .ZN(n9832) );
  INV_X1 U9891 ( .A(n8896), .ZN(n8899) );
  INV_X1 U9892 ( .A(n8897), .ZN(n8898) );
  NAND2_X1 U9893 ( .A1(n8899), .A2(n8898), .ZN(n9833) );
  NAND2_X1 U9894 ( .A1(n8900), .A2(n9833), .ZN(n9776) );
  NAND2_X1 U9895 ( .A1(n10217), .A2(n8234), .ZN(n8902) );
  NAND2_X1 U9896 ( .A1(n9886), .A2(n9042), .ZN(n8901) );
  NAND2_X1 U9897 ( .A1(n8902), .A2(n8901), .ZN(n8903) );
  XNOR2_X1 U9898 ( .A(n8903), .B(n8946), .ZN(n8906) );
  NAND2_X1 U9899 ( .A1(n10217), .A2(n9042), .ZN(n8905) );
  NAND2_X1 U9900 ( .A1(n9886), .A2(n9046), .ZN(n8904) );
  NAND2_X1 U9901 ( .A1(n8905), .A2(n8904), .ZN(n8907) );
  INV_X1 U9902 ( .A(n8906), .ZN(n8909) );
  INV_X1 U9903 ( .A(n8907), .ZN(n8908) );
  NAND2_X1 U9904 ( .A1(n8909), .A2(n8908), .ZN(n9777) );
  NAND2_X1 U9905 ( .A1(n10211), .A2(n8234), .ZN(n8911) );
  NAND2_X1 U9906 ( .A1(n9042), .A2(n10055), .ZN(n8910) );
  NAND2_X1 U9907 ( .A1(n8911), .A2(n8910), .ZN(n8912) );
  XNOR2_X1 U9908 ( .A(n8912), .B(n8946), .ZN(n8915) );
  NAND2_X1 U9909 ( .A1(n10211), .A2(n9042), .ZN(n8914) );
  NAND2_X1 U9910 ( .A1(n9046), .A2(n10055), .ZN(n8913) );
  NAND2_X1 U9911 ( .A1(n8914), .A2(n8913), .ZN(n8916) );
  NAND2_X1 U9912 ( .A1(n8915), .A2(n8916), .ZN(n9843) );
  INV_X1 U9913 ( .A(n8915), .ZN(n8918) );
  INV_X1 U9914 ( .A(n8916), .ZN(n8917) );
  NAND2_X1 U9915 ( .A1(n8918), .A2(n8917), .ZN(n9842) );
  INV_X1 U9916 ( .A(n8926), .ZN(n8923) );
  NAND2_X1 U9917 ( .A1(n10205), .A2(n8234), .ZN(n8920) );
  NAND2_X1 U9918 ( .A1(n9042), .A2(n10037), .ZN(n8919) );
  NAND2_X1 U9919 ( .A1(n8920), .A2(n8919), .ZN(n8921) );
  XNOR2_X1 U9920 ( .A(n8921), .B(n9017), .ZN(n8925) );
  NAND2_X1 U9921 ( .A1(n8923), .A2(n8922), .ZN(n9758) );
  NOR2_X1 U9922 ( .A1(n10077), .A2(n9019), .ZN(n8924) );
  AOI21_X1 U9923 ( .B1(n10205), .B2(n9042), .A(n8924), .ZN(n9760) );
  NAND2_X1 U9924 ( .A1(n9758), .A2(n9760), .ZN(n8927) );
  NAND2_X1 U9925 ( .A1(n10201), .A2(n8234), .ZN(n8929) );
  NAND2_X1 U9926 ( .A1(n9042), .A2(n10054), .ZN(n8928) );
  NAND2_X1 U9927 ( .A1(n8929), .A2(n8928), .ZN(n8930) );
  XNOR2_X1 U9928 ( .A(n8930), .B(n8946), .ZN(n8932) );
  NOR2_X1 U9929 ( .A1(n10025), .A2(n9019), .ZN(n8931) );
  AOI21_X1 U9930 ( .B1(n10201), .B2(n9042), .A(n8931), .ZN(n8933) );
  XNOR2_X1 U9931 ( .A(n8932), .B(n8933), .ZN(n9826) );
  INV_X1 U9932 ( .A(n8932), .ZN(n8934) );
  NAND2_X1 U9933 ( .A1(n8934), .A2(n8933), .ZN(n9786) );
  INV_X1 U9934 ( .A(n9786), .ZN(n8940) );
  NAND2_X1 U9935 ( .A1(n10196), .A2(n8234), .ZN(n8936) );
  NAND2_X1 U9936 ( .A1(n9042), .A2(n10038), .ZN(n8935) );
  NAND2_X1 U9937 ( .A1(n8936), .A2(n8935), .ZN(n8937) );
  XNOR2_X1 U9938 ( .A(n8937), .B(n9017), .ZN(n9789) );
  NOR2_X1 U9939 ( .A1(n9997), .A2(n9019), .ZN(n8938) );
  AOI21_X1 U9940 ( .B1(n10196), .B2(n9042), .A(n8938), .ZN(n9788) );
  AND2_X1 U9941 ( .A1(n9789), .A2(n9788), .ZN(n8939) );
  NOR2_X1 U9942 ( .A1(n8940), .A2(n8939), .ZN(n9009) );
  NAND2_X1 U9943 ( .A1(n9787), .A2(n9009), .ZN(n8943) );
  INV_X1 U9944 ( .A(n9789), .ZN(n8942) );
  INV_X1 U9945 ( .A(n9788), .ZN(n8941) );
  NAND2_X1 U9946 ( .A1(n8942), .A2(n8941), .ZN(n9000) );
  NAND2_X1 U9947 ( .A1(n8943), .A2(n9000), .ZN(n8949) );
  NAND2_X1 U9948 ( .A1(n10007), .A2(n4862), .ZN(n8945) );
  NAND2_X1 U9949 ( .A1(n9042), .A2(n9885), .ZN(n8944) );
  NAND2_X1 U9950 ( .A1(n8945), .A2(n8944), .ZN(n8947) );
  XNOR2_X1 U9951 ( .A(n8947), .B(n8946), .ZN(n9004) );
  NOR2_X1 U9952 ( .A1(n10026), .A2(n9019), .ZN(n8948) );
  AOI21_X1 U9953 ( .B1(n10007), .B2(n9042), .A(n8948), .ZN(n9002) );
  XNOR2_X1 U9954 ( .A(n9004), .B(n9002), .ZN(n9008) );
  XNOR2_X1 U9955 ( .A(n8949), .B(n9008), .ZN(n8954) );
  AOI22_X1 U9956 ( .A1(n9853), .A2(n9884), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8951) );
  NAND2_X1 U9957 ( .A1(n9873), .A2(n10038), .ZN(n8950) );
  OAI211_X1 U9958 ( .C1(n9876), .C2(n10004), .A(n8951), .B(n8950), .ZN(n8952)
         );
  AOI21_X1 U9959 ( .B1(n10007), .B2(n9863), .A(n8952), .ZN(n8953) );
  OAI21_X1 U9960 ( .B1(n8954), .B2(n9879), .A(n8953), .ZN(P1_U3238) );
  NOR2_X1 U9961 ( .A1(n10623), .A2(n8955), .ZN(n8959) );
  NAND2_X1 U9962 ( .A1(n8984), .A2(n10558), .ZN(n8957) );
  OAI211_X1 U9963 ( .C1(n9375), .C2(n10500), .A(n8957), .B(n8956), .ZN(n8958)
         );
  AOI211_X1 U9964 ( .C1(n10621), .C2(n10527), .A(n8959), .B(n8958), .ZN(n8966)
         );
  INV_X1 U9965 ( .A(n8960), .ZN(n8963) );
  OAI22_X1 U9966 ( .A1(n9129), .A2(n9375), .B1(n10615), .B2(n8961), .ZN(n8962)
         );
  NAND3_X1 U9967 ( .A1(n8964), .A2(n8963), .A3(n8962), .ZN(n8965) );
  OAI211_X1 U9968 ( .C1(n8967), .C2(n10615), .A(n8966), .B(n8965), .ZN(
        P2_U3241) );
  OAI21_X1 U9969 ( .B1(n10611), .B2(n8970), .A(n8969), .ZN(n8971) );
  AOI21_X1 U9970 ( .B1(n10609), .B2(n9371), .A(n8971), .ZN(n8972) );
  OAI21_X1 U9971 ( .B1(n8973), .B2(n10623), .A(n8972), .ZN(n8974) );
  AOI21_X1 U9972 ( .B1(n8975), .B2(n10621), .A(n8974), .ZN(n8982) );
  OAI22_X1 U9973 ( .A1(n8977), .A2(n10615), .B1(n8976), .B2(n9129), .ZN(n8978)
         );
  NAND3_X1 U9974 ( .A1(n8980), .A2(n8979), .A3(n8978), .ZN(n8981) );
  OAI211_X1 U9975 ( .C1(n8968), .C2(n10615), .A(n8982), .B(n8981), .ZN(
        P2_U3236) );
  NOR2_X1 U9976 ( .A1(n10623), .A2(n8983), .ZN(n8988) );
  NAND2_X1 U9977 ( .A1(n8984), .A2(n9369), .ZN(n8986) );
  OAI211_X1 U9978 ( .C1(n8991), .C2(n10500), .A(n8986), .B(n8985), .ZN(n8987)
         );
  AOI211_X1 U9979 ( .C1(n8989), .C2(n10621), .A(n8988), .B(n8987), .ZN(n8995)
         );
  OAI22_X1 U9980 ( .A1(n8992), .A2(n10615), .B1(n8991), .B2(n9129), .ZN(n8993)
         );
  NAND3_X1 U9981 ( .A1(n8968), .A2(n5207), .A3(n8993), .ZN(n8994) );
  OAI211_X1 U9982 ( .C1(n7741), .C2(n10615), .A(n8995), .B(n8994), .ZN(
        P2_U3217) );
  OAI222_X1 U9983 ( .A1(n8538), .A2(n8998), .B1(n8997), .B2(P2_U3152), .C1(
        n8996), .C2(n4858), .ZN(P2_U3328) );
  INV_X1 U9984 ( .A(n9008), .ZN(n9001) );
  AND2_X1 U9985 ( .A1(n9826), .A2(n9007), .ZN(n9005) );
  INV_X1 U9986 ( .A(n9002), .ZN(n9003) );
  NAND2_X1 U9987 ( .A1(n9004), .A2(n9003), .ZN(n9006) );
  AND2_X1 U9988 ( .A1(n9005), .A2(n9006), .ZN(n9027) );
  INV_X1 U9989 ( .A(n9006), .ZN(n9013) );
  INV_X1 U9990 ( .A(n9007), .ZN(n9011) );
  AND2_X1 U9991 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  INV_X1 U9992 ( .A(n9029), .ZN(n9014) );
  AOI21_X1 U9993 ( .B1(n8999), .B2(n9027), .A(n9014), .ZN(n9033) );
  NAND2_X1 U9994 ( .A1(n5955), .A2(n8234), .ZN(n9016) );
  NAND2_X1 U9995 ( .A1(n9042), .A2(n9884), .ZN(n9015) );
  NAND2_X1 U9996 ( .A1(n9016), .A2(n9015), .ZN(n9018) );
  XNOR2_X1 U9997 ( .A(n9018), .B(n9017), .ZN(n9021) );
  NOR2_X1 U9998 ( .A1(n9998), .A2(n9019), .ZN(n9020) );
  AOI21_X1 U9999 ( .B1(n5955), .B2(n9042), .A(n9020), .ZN(n9022) );
  NAND2_X1 U10000 ( .A1(n9021), .A2(n9022), .ZN(n9053) );
  INV_X1 U10001 ( .A(n9021), .ZN(n9024) );
  INV_X1 U10002 ( .A(n9022), .ZN(n9023) );
  NAND2_X1 U10003 ( .A1(n9024), .A2(n9023), .ZN(n9025) );
  NAND2_X1 U10004 ( .A1(n9053), .A2(n9025), .ZN(n9032) );
  INV_X1 U10005 ( .A(n9032), .ZN(n9026) );
  AOI22_X1 U10006 ( .A1(n9853), .A2(n9883), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9035) );
  NAND2_X1 U10007 ( .A1(n9873), .A2(n9885), .ZN(n9034) );
  OAI211_X1 U10008 ( .C1(n9876), .C2(n9981), .A(n9035), .B(n9034), .ZN(n9036)
         );
  AOI21_X1 U10009 ( .B1(n5955), .B2(n9863), .A(n9036), .ZN(n9037) );
  OAI21_X1 U10010 ( .B1(n9038), .B2(n9879), .A(n9037), .ZN(P1_U3212) );
  OAI222_X1 U10011 ( .A1(n9041), .A2(P1_U3084), .B1(n9064), .B2(n9040), .C1(
        n9039), .C2(n9060), .ZN(P1_U3331) );
  NAND2_X1 U10012 ( .A1(n10179), .A2(n4862), .ZN(n9044) );
  NAND2_X1 U10013 ( .A1(n9042), .A2(n9883), .ZN(n9043) );
  NAND2_X1 U10014 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  XNOR2_X1 U10015 ( .A(n9045), .B(n8946), .ZN(n9048) );
  AOI22_X1 U10016 ( .A1(n10179), .A2(n9042), .B1(n9046), .B2(n9883), .ZN(n9047) );
  XNOR2_X1 U10017 ( .A(n9048), .B(n9047), .ZN(n9049) );
  INV_X1 U10018 ( .A(n9049), .ZN(n9054) );
  NAND3_X1 U10019 ( .A1(n9054), .A2(n9815), .A3(n9053), .ZN(n9059) );
  NAND3_X1 U10020 ( .A1(n9050), .A2(n9815), .A3(n9049), .ZN(n9058) );
  AOI22_X1 U10021 ( .A1(n9853), .A2(n9882), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n9052) );
  NAND2_X1 U10022 ( .A1(n9873), .A2(n9884), .ZN(n9051) );
  OAI211_X1 U10023 ( .C1(n9876), .C2(n9970), .A(n9052), .B(n9051), .ZN(n9056)
         );
  NOR3_X1 U10024 ( .A1(n9054), .A2(n9879), .A3(n9053), .ZN(n9055) );
  AOI211_X1 U10025 ( .C1(n9863), .C2(n10179), .A(n9056), .B(n9055), .ZN(n9057)
         );
  OAI211_X1 U10026 ( .C1(n9050), .C2(n9059), .A(n9058), .B(n9057), .ZN(
        P1_U3218) );
  OAI222_X1 U10027 ( .A1(n9064), .A2(n9063), .B1(n5339), .B2(P1_U3084), .C1(
        n9061), .C2(n9060), .ZN(P1_U3324) );
  INV_X1 U10028 ( .A(n9066), .ZN(n9067) );
  AOI21_X1 U10029 ( .B1(n9065), .B2(n9067), .A(n10615), .ZN(n9071) );
  NOR3_X1 U10030 ( .A1(n9068), .A2(n9479), .A3(n9129), .ZN(n9070) );
  OAI21_X1 U10031 ( .B1(n9071), .B2(n9070), .A(n9069), .ZN(n9075) );
  OAI22_X1 U10032 ( .A1(n9479), .A2(n10500), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9322), .ZN(n9073) );
  NOR2_X1 U10033 ( .A1(n9480), .A2(n10611), .ZN(n9072) );
  AOI211_X1 U10034 ( .C1(n9121), .C2(n9474), .A(n9073), .B(n9072), .ZN(n9074)
         );
  OAI211_X1 U10035 ( .C1(n9476), .C2(n6546), .A(n9075), .B(n9074), .ZN(
        P2_U3216) );
  NAND2_X1 U10036 ( .A1(n9432), .A2(n10560), .ZN(n9079) );
  NAND2_X1 U10037 ( .A1(n9076), .A2(n10561), .ZN(n9078) );
  MUX2_X1 U10038 ( .A(n9079), .B(n9078), .S(n9077), .Z(n9084) );
  INV_X1 U10039 ( .A(n9080), .ZN(n9544) );
  NOR2_X1 U10040 ( .A1(n10500), .A2(n9092), .ZN(n9082) );
  OAI22_X1 U10041 ( .A1(n9107), .A2(n10611), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9247), .ZN(n9081) );
  AOI211_X1 U10042 ( .C1(n9121), .C2(n9544), .A(n9082), .B(n9081), .ZN(n9083)
         );
  OAI211_X1 U10043 ( .C1(n9546), .C2(n6546), .A(n9084), .B(n9083), .ZN(
        P2_U3218) );
  INV_X1 U10044 ( .A(n9085), .ZN(n9086) );
  AOI21_X1 U10045 ( .B1(n8268), .B2(n9086), .A(n10615), .ZN(n9090) );
  NOR3_X1 U10046 ( .A1(n9087), .A2(n9598), .A3(n9129), .ZN(n9089) );
  OAI21_X1 U10047 ( .B1(n9090), .B2(n9089), .A(n9088), .ZN(n9095) );
  AOI22_X1 U10048 ( .A1(n10609), .A2(n9570), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3152), .ZN(n9091) );
  OAI21_X1 U10049 ( .B1(n9092), .B2(n10611), .A(n9091), .ZN(n9093) );
  AOI21_X1 U10050 ( .B1(n9566), .B2(n9121), .A(n9093), .ZN(n9094) );
  OAI211_X1 U10051 ( .C1(n5026), .C2(n6546), .A(n9095), .B(n9094), .ZN(
        P2_U3225) );
  OAI211_X1 U10052 ( .C1(n9098), .C2(n9097), .A(n9096), .B(n10561), .ZN(n9105)
         );
  NOR2_X1 U10053 ( .A1(n9107), .A2(n9597), .ZN(n9099) );
  AOI21_X1 U10054 ( .B1(n9436), .B2(n9626), .A(n9099), .ZN(n9505) );
  INV_X1 U10055 ( .A(n9100), .ZN(n9512) );
  AOI22_X1 U10056 ( .A1(n9512), .A2(n9121), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n9101) );
  OAI21_X1 U10057 ( .B1(n9505), .B2(n9102), .A(n9101), .ZN(n9103) );
  AOI21_X1 U10058 ( .B1(n9667), .B2(n10621), .A(n9103), .ZN(n9104) );
  NAND2_X1 U10059 ( .A1(n9105), .A2(n9104), .ZN(P2_U3227) );
  OAI22_X1 U10060 ( .A1(n9106), .A2(n10615), .B1(n9107), .B2(n9129), .ZN(n9109) );
  NAND2_X1 U10061 ( .A1(n9109), .A2(n9108), .ZN(n9114) );
  OAI22_X1 U10062 ( .A1(n9558), .A2(n10500), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9110), .ZN(n9112) );
  NOR2_X1 U10063 ( .A1(n9528), .A2(n10611), .ZN(n9111) );
  AOI211_X1 U10064 ( .C1(n9121), .C2(n9522), .A(n9112), .B(n9111), .ZN(n9113)
         );
  OAI211_X1 U10065 ( .C1(n9524), .C2(n6546), .A(n9114), .B(n9113), .ZN(
        P2_U3231) );
  OAI21_X1 U10066 ( .B1(n9117), .B2(n9088), .A(n9115), .ZN(n9125) );
  NOR3_X1 U10067 ( .A1(n9117), .A2(n9116), .A3(n9129), .ZN(n9118) );
  OAI21_X1 U10068 ( .B1(n9118), .B2(n10609), .A(n9584), .ZN(n9123) );
  INV_X1 U10069 ( .A(n9119), .ZN(n9552) );
  OAI22_X1 U10070 ( .A1(n9558), .A2(n10611), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9352), .ZN(n9120) );
  AOI21_X1 U10071 ( .B1(n9552), .B2(n9121), .A(n9120), .ZN(n9122) );
  OAI211_X1 U10072 ( .C1(n9554), .C2(n6546), .A(n9123), .B(n9122), .ZN(n9124)
         );
  AOI21_X1 U10073 ( .B1(n9125), .B2(n10561), .A(n9124), .ZN(n9126) );
  INV_X1 U10074 ( .A(n9126), .ZN(P2_U3237) );
  INV_X1 U10075 ( .A(n9661), .ZN(n9140) );
  INV_X1 U10076 ( .A(n9127), .ZN(n9128) );
  AOI21_X1 U10077 ( .B1(n9096), .B2(n9128), .A(n10615), .ZN(n9132) );
  NOR3_X1 U10078 ( .A1(n9130), .A2(n9528), .A3(n9129), .ZN(n9131) );
  OAI21_X1 U10079 ( .B1(n9132), .B2(n9131), .A(n9065), .ZN(n9139) );
  OR2_X1 U10080 ( .A1(n9142), .A2(n9599), .ZN(n9135) );
  NAND2_X1 U10081 ( .A1(n9133), .A2(n9624), .ZN(n9134) );
  NAND2_X1 U10082 ( .A1(n9135), .A2(n9134), .ZN(n9491) );
  OAI22_X1 U10083 ( .A1(n9495), .A2(n10623), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9361), .ZN(n9136) );
  AOI21_X1 U10084 ( .B1(n9491), .B2(n9137), .A(n9136), .ZN(n9138) );
  OAI211_X1 U10085 ( .C1(n9140), .C2(n6546), .A(n9139), .B(n9138), .ZN(
        P2_U3242) );
  MUX2_X1 U10086 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9141), .S(P2_U3966), .Z(
        P2_U3580) );
  INV_X1 U10087 ( .A(n9142), .ZN(n9437) );
  MUX2_X1 U10088 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9437), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10089 ( .A(n9432), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9143), .Z(
        P2_U3575) );
  MUX2_X1 U10090 ( .A(n9571), .B(P2_DATAO_REG_22__SCAN_IN), .S(n9143), .Z(
        P2_U3574) );
  MUX2_X1 U10091 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9584), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10092 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9625), .S(n9370), .Z(
        n9367) );
  INV_X1 U10093 ( .A(keyinput_127), .ZN(n9145) );
  XOR2_X1 U10094 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_126), .Z(n9144) );
  AOI221_X1 U10095 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(n9145), .C1(n6305), 
        .C2(keyinput_127), .A(n9144), .ZN(n9365) );
  AOI22_X1 U10096 ( .A1(n6178), .A2(keyinput_117), .B1(keyinput_114), .B2(
        n9340), .ZN(n9146) );
  OAI221_X1 U10097 ( .B1(n6178), .B2(keyinput_117), .C1(n9340), .C2(
        keyinput_114), .A(n9146), .ZN(n9153) );
  AOI22_X1 U10098 ( .A1(n6445), .A2(keyinput_111), .B1(n6304), .B2(
        keyinput_112), .ZN(n9147) );
  OAI221_X1 U10099 ( .B1(n6445), .B2(keyinput_111), .C1(n6304), .C2(
        keyinput_112), .A(n9147), .ZN(n9152) );
  AOI22_X1 U10100 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_118), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_116), .ZN(n9148) );
  OAI221_X1 U10101 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_116), .A(n9148), .ZN(n9151) );
  AOI22_X1 U10102 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_115), .B1(
        P2_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .ZN(n9149) );
  OAI221_X1 U10103 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_113), .A(n9149), .ZN(n9150) );
  NOR4_X1 U10104 ( .A1(n9153), .A2(n9152), .A3(n9151), .A4(n9150), .ZN(n9234)
         );
  INV_X1 U10105 ( .A(keyinput_110), .ZN(n9232) );
  INV_X1 U10106 ( .A(keyinput_109), .ZN(n9230) );
  INV_X1 U10107 ( .A(keyinput_108), .ZN(n9228) );
  OAI22_X1 U10108 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_102), .B1(
        keyinput_106), .B2(P2_REG3_REG_28__SCAN_IN), .ZN(n9154) );
  AOI221_X1 U10109 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_102), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_106), .A(n9154), .ZN(n9226) );
  OAI22_X1 U10110 ( .A1(n10499), .A2(keyinput_104), .B1(keyinput_103), .B2(
        P2_REG3_REG_10__SCAN_IN), .ZN(n9155) );
  AOI221_X1 U10111 ( .B1(n10499), .B2(keyinput_104), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_103), .A(n9155), .ZN(n9225) );
  OAI22_X1 U10112 ( .A1(n9157), .A2(keyinput_107), .B1(n9248), .B2(
        keyinput_105), .ZN(n9156) );
  AOI221_X1 U10113 ( .B1(n9157), .B2(keyinput_107), .C1(keyinput_105), .C2(
        n9248), .A(n9156), .ZN(n9224) );
  INV_X1 U10114 ( .A(keyinput_101), .ZN(n9222) );
  INV_X1 U10115 ( .A(keyinput_96), .ZN(n9158) );
  MUX2_X1 U10116 ( .A(keyinput_96), .B(n9158), .S(SI_0_), .Z(n9159) );
  INV_X1 U10117 ( .A(n9159), .ZN(n9216) );
  INV_X1 U10118 ( .A(keyinput_93), .ZN(n9207) );
  INV_X1 U10119 ( .A(SI_6_), .ZN(n9161) );
  OAI22_X1 U10120 ( .A1(n9161), .A2(keyinput_90), .B1(keyinput_89), .B2(SI_7_), 
        .ZN(n9160) );
  AOI221_X1 U10121 ( .B1(n9161), .B2(keyinput_90), .C1(SI_7_), .C2(keyinput_89), .A(n9160), .ZN(n9205) );
  INV_X1 U10122 ( .A(SI_11_), .ZN(n9292) );
  OAI22_X1 U10123 ( .A1(n9285), .A2(keyinput_81), .B1(n9163), .B2(keyinput_82), 
        .ZN(n9162) );
  AOI221_X1 U10124 ( .B1(n9285), .B2(keyinput_81), .C1(keyinput_82), .C2(n9163), .A(n9162), .ZN(n9169) );
  OAI22_X1 U10125 ( .A1(SI_18_), .A2(keyinput_78), .B1(keyinput_79), .B2(
        SI_17_), .ZN(n9164) );
  AOI221_X1 U10126 ( .B1(SI_18_), .B2(keyinput_78), .C1(SI_17_), .C2(
        keyinput_79), .A(n9164), .ZN(n9168) );
  OAI22_X1 U10127 ( .A1(SI_16_), .A2(keyinput_80), .B1(SI_12_), .B2(
        keyinput_84), .ZN(n9165) );
  AOI221_X1 U10128 ( .B1(SI_16_), .B2(keyinput_80), .C1(keyinput_84), .C2(
        SI_12_), .A(n9165), .ZN(n9167) );
  XNOR2_X1 U10129 ( .A(SI_13_), .B(keyinput_83), .ZN(n9166) );
  NAND4_X1 U10130 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .ZN(n9195)
         );
  INV_X1 U10131 ( .A(keyinput_77), .ZN(n9193) );
  INV_X1 U10132 ( .A(keyinput_76), .ZN(n9191) );
  AOI22_X1 U10133 ( .A1(SI_22_), .A2(keyinput_74), .B1(SI_23_), .B2(
        keyinput_73), .ZN(n9170) );
  OAI221_X1 U10134 ( .B1(SI_22_), .B2(keyinput_74), .C1(SI_23_), .C2(
        keyinput_73), .A(n9170), .ZN(n9188) );
  INV_X1 U10135 ( .A(keyinput_72), .ZN(n9186) );
  OAI22_X1 U10136 ( .A1(n9173), .A2(keyinput_69), .B1(n9172), .B2(keyinput_70), 
        .ZN(n9171) );
  AOI221_X1 U10137 ( .B1(n9173), .B2(keyinput_69), .C1(keyinput_70), .C2(n9172), .A(n9171), .ZN(n9182) );
  INV_X1 U10138 ( .A(keyinput_68), .ZN(n9180) );
  INV_X1 U10139 ( .A(keyinput_67), .ZN(n9178) );
  INV_X1 U10140 ( .A(keyinput_66), .ZN(n9176) );
  OAI22_X1 U10141 ( .A1(SI_31_), .A2(keyinput_65), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_64), .ZN(n9174) );
  AOI221_X1 U10142 ( .B1(SI_31_), .B2(keyinput_65), .C1(keyinput_64), .C2(
        P2_WR_REG_SCAN_IN), .A(n9174), .ZN(n9175) );
  OAI221_X1 U10143 ( .B1(SI_30_), .B2(keyinput_66), .C1(n9258), .C2(n9176), 
        .A(n9175), .ZN(n9177) );
  OAI221_X1 U10144 ( .B1(SI_29_), .B2(n9178), .C1(n9260), .C2(keyinput_67), 
        .A(n9177), .ZN(n9179) );
  OAI221_X1 U10145 ( .B1(SI_28_), .B2(n9180), .C1(n9263), .C2(keyinput_68), 
        .A(n9179), .ZN(n9181) );
  OAI211_X1 U10146 ( .C1(n9184), .C2(keyinput_71), .A(n9182), .B(n9181), .ZN(
        n9183) );
  AOI21_X1 U10147 ( .B1(n9184), .B2(keyinput_71), .A(n9183), .ZN(n9185) );
  AOI221_X1 U10148 ( .B1(SI_24_), .B2(n9186), .C1(n9271), .C2(keyinput_72), 
        .A(n9185), .ZN(n9187) );
  OAI22_X1 U10149 ( .A1(n9188), .A2(n9187), .B1(keyinput_75), .B2(SI_21_), 
        .ZN(n9189) );
  AOI21_X1 U10150 ( .B1(keyinput_75), .B2(SI_21_), .A(n9189), .ZN(n9190) );
  AOI221_X1 U10151 ( .B1(SI_20_), .B2(keyinput_76), .C1(n9277), .C2(n9191), 
        .A(n9190), .ZN(n9192) );
  AOI221_X1 U10152 ( .B1(SI_19_), .B2(keyinput_77), .C1(n9280), .C2(n9193), 
        .A(n9192), .ZN(n9194) );
  OAI22_X1 U10153 ( .A1(keyinput_85), .A2(n9292), .B1(n9195), .B2(n9194), .ZN(
        n9196) );
  AOI21_X1 U10154 ( .B1(keyinput_85), .B2(n9292), .A(n9196), .ZN(n9199) );
  AOI22_X1 U10155 ( .A1(SI_8_), .A2(keyinput_88), .B1(n9296), .B2(keyinput_87), 
        .ZN(n9197) );
  OAI221_X1 U10156 ( .B1(SI_8_), .B2(keyinput_88), .C1(n9296), .C2(keyinput_87), .A(n9197), .ZN(n9198) );
  AOI211_X1 U10157 ( .C1(SI_10_), .C2(keyinput_86), .A(n9199), .B(n9198), .ZN(
        n9200) );
  OAI21_X1 U10158 ( .B1(SI_10_), .B2(keyinput_86), .A(n9200), .ZN(n9204) );
  INV_X1 U10159 ( .A(SI_5_), .ZN(n9202) );
  INV_X1 U10160 ( .A(SI_4_), .ZN(n9302) );
  AOI22_X1 U10161 ( .A1(n9202), .A2(keyinput_91), .B1(keyinput_92), .B2(n9302), 
        .ZN(n9201) );
  OAI221_X1 U10162 ( .B1(n9202), .B2(keyinput_91), .C1(n9302), .C2(keyinput_92), .A(n9201), .ZN(n9203) );
  AOI21_X1 U10163 ( .B1(n9205), .B2(n9204), .A(n9203), .ZN(n9206) );
  AOI221_X1 U10164 ( .B1(SI_3_), .B2(keyinput_93), .C1(n9308), .C2(n9207), .A(
        n9206), .ZN(n9213) );
  INV_X1 U10165 ( .A(keyinput_94), .ZN(n9208) );
  MUX2_X1 U10166 ( .A(keyinput_94), .B(n9208), .S(SI_2_), .Z(n9212) );
  INV_X1 U10167 ( .A(keyinput_95), .ZN(n9209) );
  MUX2_X1 U10168 ( .A(n9209), .B(keyinput_95), .S(SI_1_), .Z(n9210) );
  INV_X1 U10169 ( .A(n9210), .ZN(n9211) );
  OAI21_X1 U10170 ( .B1(n9213), .B2(n9212), .A(n9211), .ZN(n9215) );
  INV_X1 U10171 ( .A(keyinput_97), .ZN(n9214) );
  AOI222_X1 U10172 ( .A1(n9216), .A2(n9215), .B1(P2_RD_REG_SCAN_IN), .B2(n9214), .C1(n5112), .C2(keyinput_97), .ZN(n9219) );
  AOI22_X1 U10173 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_100), .B1(n6144), .B2(keyinput_99), .ZN(n9217) );
  OAI221_X1 U10174 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .C1(
        n6144), .C2(keyinput_99), .A(n9217), .ZN(n9218) );
  AOI211_X1 U10175 ( .C1(P2_STATE_REG_SCAN_IN), .C2(keyinput_98), .A(n9219), 
        .B(n9218), .ZN(n9220) );
  OAI21_X1 U10176 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_98), .A(n9220), 
        .ZN(n9221) );
  OAI221_X1 U10177 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .C1(
        n9325), .C2(n9222), .A(n9221), .ZN(n9223) );
  NAND4_X1 U10178 ( .A1(n9226), .A2(n9225), .A3(n9224), .A4(n9223), .ZN(n9227)
         );
  OAI221_X1 U10179 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_108), .C1(n9332), .C2(n9228), .A(n9227), .ZN(n9229) );
  OAI221_X1 U10180 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(n9230), .C1(n9334), 
        .C2(keyinput_109), .A(n9229), .ZN(n9231) );
  OAI221_X1 U10181 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .C1(
        n9337), .C2(n9232), .A(n9231), .ZN(n9233) );
  AOI22_X1 U10182 ( .A1(n9234), .A2(n9233), .B1(keyinput_120), .B2(n6235), 
        .ZN(n9235) );
  OAI21_X1 U10183 ( .B1(keyinput_120), .B2(n6235), .A(n9235), .ZN(n9243) );
  AOI22_X1 U10184 ( .A1(n9352), .A2(keyinput_121), .B1(n9237), .B2(
        keyinput_119), .ZN(n9236) );
  OAI221_X1 U10185 ( .B1(n9352), .B2(keyinput_121), .C1(n9237), .C2(
        keyinput_119), .A(n9236), .ZN(n9242) );
  OAI22_X1 U10186 ( .A1(n7631), .A2(keyinput_123), .B1(keyinput_122), .B2(
        P2_REG3_REG_11__SCAN_IN), .ZN(n9238) );
  AOI221_X1 U10187 ( .B1(n7631), .B2(keyinput_123), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_122), .A(n9238), .ZN(n9241) );
  OAI22_X1 U10188 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_125), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .ZN(n9239) );
  AOI221_X1 U10189 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .C1(
        keyinput_124), .C2(P2_REG3_REG_18__SCAN_IN), .A(n9239), .ZN(n9240) );
  OAI211_X1 U10190 ( .C1(n9243), .C2(n9242), .A(n9241), .B(n9240), .ZN(n9364)
         );
  INV_X1 U10191 ( .A(keyinput_46), .ZN(n9338) );
  INV_X1 U10192 ( .A(keyinput_45), .ZN(n9335) );
  INV_X1 U10193 ( .A(keyinput_44), .ZN(n9331) );
  OAI22_X1 U10194 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_39), .B1(
        keyinput_42), .B2(P2_REG3_REG_28__SCAN_IN), .ZN(n9244) );
  AOI221_X1 U10195 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_42), .A(n9244), .ZN(n9329) );
  OAI22_X1 U10196 ( .A1(n10499), .A2(keyinput_40), .B1(keyinput_43), .B2(
        P2_REG3_REG_8__SCAN_IN), .ZN(n9245) );
  AOI221_X1 U10197 ( .B1(n10499), .B2(keyinput_40), .C1(P2_REG3_REG_8__SCAN_IN), .C2(keyinput_43), .A(n9245), .ZN(n9328) );
  OAI22_X1 U10198 ( .A1(n9248), .A2(keyinput_41), .B1(n9247), .B2(keyinput_38), 
        .ZN(n9246) );
  AOI221_X1 U10199 ( .B1(n9248), .B2(keyinput_41), .C1(keyinput_38), .C2(n9247), .A(n9246), .ZN(n9327) );
  INV_X1 U10200 ( .A(keyinput_37), .ZN(n9324) );
  INV_X1 U10201 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9322) );
  INV_X1 U10202 ( .A(keyinput_32), .ZN(n9249) );
  MUX2_X1 U10203 ( .A(keyinput_32), .B(n9249), .S(SI_0_), .Z(n9250) );
  INV_X1 U10204 ( .A(n9250), .ZN(n9317) );
  INV_X1 U10205 ( .A(keyinput_29), .ZN(n9307) );
  INV_X1 U10206 ( .A(SI_7_), .ZN(n9252) );
  OAI22_X1 U10207 ( .A1(n9252), .A2(keyinput_25), .B1(keyinput_26), .B2(SI_6_), 
        .ZN(n9251) );
  AOI221_X1 U10208 ( .B1(n9252), .B2(keyinput_25), .C1(SI_6_), .C2(keyinput_26), .A(n9251), .ZN(n9305) );
  INV_X1 U10209 ( .A(keyinput_13), .ZN(n9279) );
  INV_X1 U10210 ( .A(keyinput_12), .ZN(n9276) );
  OAI22_X1 U10211 ( .A1(n9254), .A2(keyinput_9), .B1(SI_22_), .B2(keyinput_10), 
        .ZN(n9253) );
  AOI221_X1 U10212 ( .B1(n9254), .B2(keyinput_9), .C1(keyinput_10), .C2(SI_22_), .A(n9253), .ZN(n9273) );
  INV_X1 U10213 ( .A(keyinput_8), .ZN(n9270) );
  INV_X1 U10214 ( .A(keyinput_4), .ZN(n9264) );
  INV_X1 U10215 ( .A(keyinput_3), .ZN(n9261) );
  INV_X1 U10216 ( .A(keyinput_2), .ZN(n9257) );
  AOI22_X1 U10217 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n9255) );
  OAI221_X1 U10218 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n9255), .ZN(n9256) );
  AOI221_X1 U10219 ( .B1(SI_30_), .B2(keyinput_2), .C1(n9258), .C2(n9257), .A(
        n9256), .ZN(n9259) );
  AOI221_X1 U10220 ( .B1(SI_29_), .B2(n9261), .C1(n9260), .C2(keyinput_3), .A(
        n9259), .ZN(n9262) );
  AOI221_X1 U10221 ( .B1(SI_28_), .B2(n9264), .C1(n9263), .C2(keyinput_4), .A(
        n9262), .ZN(n9267) );
  AOI22_X1 U10222 ( .A1(SI_25_), .A2(keyinput_7), .B1(SI_26_), .B2(keyinput_6), 
        .ZN(n9265) );
  OAI221_X1 U10223 ( .B1(SI_25_), .B2(keyinput_7), .C1(SI_26_), .C2(keyinput_6), .A(n9265), .ZN(n9266) );
  AOI211_X1 U10224 ( .C1(SI_27_), .C2(keyinput_5), .A(n9267), .B(n9266), .ZN(
        n9268) );
  OAI21_X1 U10225 ( .B1(SI_27_), .B2(keyinput_5), .A(n9268), .ZN(n9269) );
  OAI221_X1 U10226 ( .B1(SI_24_), .B2(keyinput_8), .C1(n9271), .C2(n9270), .A(
        n9269), .ZN(n9272) );
  AOI22_X1 U10227 ( .A1(n9273), .A2(n9272), .B1(keyinput_11), .B2(SI_21_), 
        .ZN(n9274) );
  OAI21_X1 U10228 ( .B1(keyinput_11), .B2(SI_21_), .A(n9274), .ZN(n9275) );
  OAI221_X1 U10229 ( .B1(SI_20_), .B2(keyinput_12), .C1(n9277), .C2(n9276), 
        .A(n9275), .ZN(n9278) );
  OAI221_X1 U10230 ( .B1(SI_19_), .B2(keyinput_13), .C1(n9280), .C2(n9279), 
        .A(n9278), .ZN(n9294) );
  XOR2_X1 U10231 ( .A(SI_14_), .B(keyinput_18), .Z(n9290) );
  AOI22_X1 U10232 ( .A1(n9283), .A2(keyinput_19), .B1(n9282), .B2(keyinput_16), 
        .ZN(n9281) );
  OAI221_X1 U10233 ( .B1(n9283), .B2(keyinput_19), .C1(n9282), .C2(keyinput_16), .A(n9281), .ZN(n9289) );
  AOI22_X1 U10234 ( .A1(SI_12_), .A2(keyinput_20), .B1(n9285), .B2(keyinput_17), .ZN(n9284) );
  OAI221_X1 U10235 ( .B1(SI_12_), .B2(keyinput_20), .C1(n9285), .C2(
        keyinput_17), .A(n9284), .ZN(n9288) );
  AOI22_X1 U10236 ( .A1(SI_17_), .A2(keyinput_15), .B1(SI_18_), .B2(
        keyinput_14), .ZN(n9286) );
  OAI221_X1 U10237 ( .B1(SI_17_), .B2(keyinput_15), .C1(SI_18_), .C2(
        keyinput_14), .A(n9286), .ZN(n9287) );
  NOR4_X1 U10238 ( .A1(n9290), .A2(n9289), .A3(n9288), .A4(n9287), .ZN(n9293)
         );
  NOR2_X1 U10239 ( .A1(n9292), .A2(keyinput_21), .ZN(n9291) );
  AOI221_X1 U10240 ( .B1(n9294), .B2(n9293), .C1(keyinput_21), .C2(n9292), .A(
        n9291), .ZN(n9298) );
  AOI22_X1 U10241 ( .A1(SI_10_), .A2(keyinput_22), .B1(n9296), .B2(keyinput_23), .ZN(n9295) );
  OAI221_X1 U10242 ( .B1(SI_10_), .B2(keyinput_22), .C1(n9296), .C2(
        keyinput_23), .A(n9295), .ZN(n9297) );
  AOI211_X1 U10243 ( .C1(n9300), .C2(keyinput_24), .A(n9298), .B(n9297), .ZN(
        n9299) );
  OAI21_X1 U10244 ( .B1(n9300), .B2(keyinput_24), .A(n9299), .ZN(n9304) );
  AOI22_X1 U10245 ( .A1(SI_5_), .A2(keyinput_27), .B1(n9302), .B2(keyinput_28), 
        .ZN(n9301) );
  OAI221_X1 U10246 ( .B1(SI_5_), .B2(keyinput_27), .C1(n9302), .C2(keyinput_28), .A(n9301), .ZN(n9303) );
  AOI21_X1 U10247 ( .B1(n9305), .B2(n9304), .A(n9303), .ZN(n9306) );
  AOI221_X1 U10248 ( .B1(SI_3_), .B2(keyinput_29), .C1(n9308), .C2(n9307), .A(
        n9306), .ZN(n9314) );
  INV_X1 U10249 ( .A(keyinput_30), .ZN(n9309) );
  MUX2_X1 U10250 ( .A(n9309), .B(keyinput_30), .S(SI_2_), .Z(n9313) );
  INV_X1 U10251 ( .A(keyinput_31), .ZN(n9310) );
  MUX2_X1 U10252 ( .A(n9310), .B(keyinput_31), .S(SI_1_), .Z(n9311) );
  INV_X1 U10253 ( .A(n9311), .ZN(n9312) );
  OAI21_X1 U10254 ( .B1(n9314), .B2(n9313), .A(n9312), .ZN(n9316) );
  INV_X1 U10255 ( .A(keyinput_33), .ZN(n9315) );
  AOI222_X1 U10256 ( .A1(n9317), .A2(n9316), .B1(n5112), .B2(n9315), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_33), .ZN(n9320) );
  AOI22_X1 U10257 ( .A1(n6144), .A2(keyinput_35), .B1(keyinput_34), .B2(
        P2_U3152), .ZN(n9318) );
  OAI221_X1 U10258 ( .B1(n6144), .B2(keyinput_35), .C1(P2_U3152), .C2(
        keyinput_34), .A(n9318), .ZN(n9319) );
  AOI211_X1 U10259 ( .C1(n9322), .C2(keyinput_36), .A(n9320), .B(n9319), .ZN(
        n9321) );
  OAI21_X1 U10260 ( .B1(n9322), .B2(keyinput_36), .A(n9321), .ZN(n9323) );
  OAI221_X1 U10261 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(n9325), .C2(n9324), .A(n9323), .ZN(n9326) );
  NAND4_X1 U10262 ( .A1(n9329), .A2(n9328), .A3(n9327), .A4(n9326), .ZN(n9330)
         );
  OAI221_X1 U10263 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .C1(n9332), 
        .C2(n9331), .A(n9330), .ZN(n9333) );
  OAI221_X1 U10264 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(n9335), .C1(n9334), 
        .C2(keyinput_45), .A(n9333), .ZN(n9336) );
  OAI221_X1 U10265 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(n9338), .C1(n9337), 
        .C2(keyinput_46), .A(n9336), .ZN(n9350) );
  AOI22_X1 U10266 ( .A1(n6445), .A2(keyinput_47), .B1(n9340), .B2(keyinput_50), 
        .ZN(n9339) );
  OAI221_X1 U10267 ( .B1(n6445), .B2(keyinput_47), .C1(n9340), .C2(keyinput_50), .A(n9339), .ZN(n9347) );
  AOI22_X1 U10268 ( .A1(n6111), .A2(keyinput_49), .B1(keyinput_48), .B2(n6304), 
        .ZN(n9341) );
  OAI221_X1 U10269 ( .B1(n6111), .B2(keyinput_49), .C1(n6304), .C2(keyinput_48), .A(n9341), .ZN(n9346) );
  AOI22_X1 U10270 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_53), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .ZN(n9342) );
  OAI221_X1 U10271 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_52), .A(n9342), .ZN(n9345) );
  AOI22_X1 U10272 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_54), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .ZN(n9343) );
  OAI221_X1 U10273 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_51), .A(n9343), .ZN(n9344) );
  NOR4_X1 U10274 ( .A1(n9347), .A2(n9346), .A3(n9345), .A4(n9344), .ZN(n9349)
         );
  NOR2_X1 U10275 ( .A1(keyinput_55), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n9348)
         );
  AOI221_X1 U10276 ( .B1(n9350), .B2(n9349), .C1(P2_REG3_REG_20__SCAN_IN), 
        .C2(keyinput_55), .A(n9348), .ZN(n9359) );
  OAI22_X1 U10277 ( .A1(n6235), .A2(keyinput_56), .B1(n9352), .B2(keyinput_57), 
        .ZN(n9351) );
  AOI221_X1 U10278 ( .B1(n6235), .B2(keyinput_56), .C1(keyinput_57), .C2(n9352), .A(n9351), .ZN(n9358) );
  INV_X1 U10279 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9354) );
  AOI22_X1 U10280 ( .A1(n7998), .A2(keyinput_60), .B1(n9354), .B2(keyinput_61), 
        .ZN(n9353) );
  OAI221_X1 U10281 ( .B1(n7998), .B2(keyinput_60), .C1(n9354), .C2(keyinput_61), .A(n9353), .ZN(n9357) );
  AOI22_X1 U10282 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(n9400), 
        .B2(keyinput_58), .ZN(n9355) );
  OAI221_X1 U10283 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(n9400), 
        .C2(keyinput_58), .A(n9355), .ZN(n9356) );
  AOI211_X1 U10284 ( .C1(n9359), .C2(n9358), .A(n9357), .B(n9356), .ZN(n9363)
         );
  AOI22_X1 U10285 ( .A1(n6305), .A2(keyinput_63), .B1(keyinput_62), .B2(n9361), 
        .ZN(n9360) );
  OAI221_X1 U10286 ( .B1(n6305), .B2(keyinput_63), .C1(n9361), .C2(keyinput_62), .A(n9360), .ZN(n9362) );
  AOI211_X1 U10287 ( .C1(n9365), .C2(n9364), .A(n9363), .B(n9362), .ZN(n9366)
         );
  XOR2_X1 U10288 ( .A(n9367), .B(n9366), .Z(P2_U3569) );
  MUX2_X1 U10289 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9368), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10290 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9369), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10291 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9371), .S(n9370), .Z(
        P2_U3564) );
  MUX2_X1 U10292 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9372), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10293 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n9374), .S(P2_U3966), .Z(
        P2_U3560) );
  INV_X1 U10294 ( .A(n9375), .ZN(n9376) );
  MUX2_X1 U10295 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n9376), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10296 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n9377), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10297 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9378), .S(n9370), .Z(
        P2_U3555) );
  MUX2_X1 U10298 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6947), .S(n9370), .Z(
        P2_U3554) );
  MUX2_X1 U10299 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9379), .S(n9370), .Z(
        P2_U3553) );
  MUX2_X1 U10300 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6870), .S(n9370), .Z(
        P2_U3552) );
  INV_X1 U10301 ( .A(n9380), .ZN(n9383) );
  NOR2_X1 U10302 ( .A1(n10426), .A2(n9381), .ZN(n9382) );
  AOI211_X1 U10303 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n10448), .A(n9383), .B(
        n9382), .ZN(n9395) );
  INV_X1 U10304 ( .A(n9384), .ZN(n9385) );
  OAI211_X1 U10305 ( .C1(n9387), .C2(n9386), .A(n10425), .B(n9385), .ZN(n9394)
         );
  OR3_X1 U10306 ( .A1(n9390), .A2(n9389), .A3(n9388), .ZN(n9391) );
  NAND3_X1 U10307 ( .A1(n9392), .A2(n10457), .A3(n9391), .ZN(n9393) );
  NAND3_X1 U10308 ( .A1(n9395), .A2(n9394), .A3(n9393), .ZN(P2_U3254) );
  OAI21_X1 U10309 ( .B1(n9398), .B2(n9397), .A(n9396), .ZN(n9399) );
  NAND2_X1 U10310 ( .A1(n10425), .A2(n9399), .ZN(n9409) );
  NOR2_X1 U10311 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9400), .ZN(n9401) );
  AOI21_X1 U10312 ( .B1(n10448), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9401), .ZN(
        n9408) );
  NAND2_X1 U10313 ( .A1(n10455), .A2(n9402), .ZN(n9407) );
  OAI211_X1 U10314 ( .C1(n9405), .C2(n9404), .A(n10457), .B(n9403), .ZN(n9406)
         );
  NAND4_X1 U10315 ( .A1(n9409), .A2(n9408), .A3(n9407), .A4(n9406), .ZN(
        P2_U3256) );
  OAI211_X1 U10316 ( .C1(n9411), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10457), .B(
        n9410), .ZN(n9421) );
  INV_X1 U10317 ( .A(n9412), .ZN(n9413) );
  AOI21_X1 U10318 ( .B1(n10448), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n9413), .ZN(
        n9420) );
  OAI21_X1 U10319 ( .B1(n9415), .B2(n6289), .A(n9414), .ZN(n9416) );
  NAND2_X1 U10320 ( .A1(n9416), .A2(n10425), .ZN(n9419) );
  NAND2_X1 U10321 ( .A1(n10455), .A2(n9417), .ZN(n9418) );
  NAND4_X1 U10322 ( .A1(n9421), .A2(n9420), .A3(n9419), .A4(n9418), .ZN(
        P2_U3260) );
  INV_X1 U10323 ( .A(n9423), .ZN(n9643) );
  INV_X1 U10324 ( .A(n9422), .ZN(n9640) );
  NAND2_X1 U10325 ( .A1(n9423), .A2(n9450), .ZN(n9639) );
  NAND3_X1 U10326 ( .A1(n9640), .A2(n9632), .A3(n9639), .ZN(n9426) );
  AOI21_X1 U10327 ( .B1(n9618), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9424), .ZN(
        n9425) );
  OAI211_X1 U10328 ( .C1(n9643), .C2(n9620), .A(n9426), .B(n9425), .ZN(
        P2_U3266) );
  OAI21_X1 U10329 ( .B1(n9710), .B2(n9625), .A(n9427), .ZN(n9611) );
  NAND2_X1 U10330 ( .A1(n9603), .A2(n9602), .ZN(n9604) );
  NAND2_X1 U10331 ( .A1(n9604), .A2(n5308), .ZN(n9577) );
  AOI21_X1 U10332 ( .B1(n9432), .B2(n9676), .A(n9681), .ZN(n9520) );
  NAND2_X1 U10333 ( .A1(n9520), .A2(n9526), .ZN(n9519) );
  NAND2_X1 U10334 ( .A1(n9519), .A2(n9433), .ZN(n9499) );
  INV_X1 U10335 ( .A(n9667), .ZN(n9515) );
  XNOR2_X1 U10336 ( .A(n9439), .B(n9440), .ZN(n9644) );
  INV_X1 U10337 ( .A(n9644), .ZN(n9459) );
  INV_X1 U10338 ( .A(n9440), .ZN(n9441) );
  OAI22_X1 U10339 ( .A1(n9480), .A2(n9597), .B1(n9445), .B2(n9444), .ZN(n9446)
         );
  INV_X1 U10340 ( .A(n9446), .ZN(n9447) );
  INV_X1 U10341 ( .A(n9645), .ZN(n9454) );
  INV_X1 U10342 ( .A(n9449), .ZN(n9461) );
  OAI21_X1 U10343 ( .B1(n9454), .B2(n9461), .A(n9450), .ZN(n9646) );
  NOR2_X1 U10344 ( .A1(n9646), .A2(n9451), .ZN(n9456) );
  AOI22_X1 U10345 ( .A1(n9452), .A2(n9616), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9618), .ZN(n9453) );
  OAI21_X1 U10346 ( .B1(n9454), .B2(n9620), .A(n9453), .ZN(n9455) );
  AOI211_X1 U10347 ( .C1(n9647), .C2(n9457), .A(n9456), .B(n9455), .ZN(n9458)
         );
  OAI21_X1 U10348 ( .B1(n9459), .B2(n9634), .A(n9458), .ZN(P2_U3267) );
  XNOR2_X1 U10349 ( .A(n9460), .B(n9465), .ZN(n9654) );
  AOI21_X1 U10350 ( .B1(n9650), .B2(n5013), .A(n9461), .ZN(n9651) );
  AOI22_X1 U10351 ( .A1(n9462), .A2(n9616), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9618), .ZN(n9463) );
  OAI21_X1 U10352 ( .B1(n9464), .B2(n9620), .A(n9463), .ZN(n9470) );
  XNOR2_X1 U10353 ( .A(n9466), .B(n9465), .ZN(n9468) );
  NOR2_X1 U10354 ( .A1(n9653), .A2(n9618), .ZN(n9469) );
  AOI211_X1 U10355 ( .C1(n9632), .C2(n9651), .A(n9470), .B(n9469), .ZN(n9471)
         );
  OAI21_X1 U10356 ( .B1(n9654), .B2(n9634), .A(n9471), .ZN(P2_U3268) );
  XNOR2_X1 U10357 ( .A(n9472), .B(n8328), .ZN(n9659) );
  AOI21_X1 U10358 ( .B1(n9655), .B2(n5014), .A(n9473), .ZN(n9656) );
  AOI22_X1 U10359 ( .A1(n9474), .A2(n9616), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9618), .ZN(n9475) );
  OAI21_X1 U10360 ( .B1(n9476), .B2(n9620), .A(n9475), .ZN(n9485) );
  AOI21_X1 U10361 ( .B1(n9478), .B2(n9477), .A(n9594), .ZN(n9483) );
  OAI22_X1 U10362 ( .A1(n9480), .A2(n9599), .B1(n9479), .B2(n9597), .ZN(n9481)
         );
  AOI21_X1 U10363 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9658) );
  NOR2_X1 U10364 ( .A1(n9658), .A2(n9618), .ZN(n9484) );
  AOI211_X1 U10365 ( .C1(n9632), .C2(n9656), .A(n9485), .B(n9484), .ZN(n9486)
         );
  OAI21_X1 U10366 ( .B1(n9659), .B2(n9634), .A(n9486), .ZN(P2_U3269) );
  XOR2_X1 U10367 ( .A(n9490), .B(n9487), .Z(n9664) );
  AOI22_X1 U10368 ( .A1(n9661), .A2(n9606), .B1(n9618), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U10369 ( .A1(n9502), .A2(n9488), .ZN(n9489) );
  XOR2_X1 U10370 ( .A(n9490), .B(n9489), .Z(n9492) );
  AOI21_X1 U10371 ( .B1(n9492), .B2(n9629), .A(n9491), .ZN(n9663) );
  AOI211_X1 U10372 ( .C1(n9661), .C2(n9508), .A(n10678), .B(n9493), .ZN(n9660)
         );
  NAND2_X1 U10373 ( .A1(n9660), .A2(n9601), .ZN(n9494) );
  OAI211_X1 U10374 ( .C1(n9592), .C2(n9495), .A(n9663), .B(n9494), .ZN(n9496)
         );
  NAND2_X1 U10375 ( .A1(n9496), .A2(n9517), .ZN(n9497) );
  OAI211_X1 U10376 ( .C1(n9664), .C2(n9634), .A(n9498), .B(n9497), .ZN(
        P2_U3270) );
  XNOR2_X1 U10377 ( .A(n9499), .B(n9504), .ZN(n9669) );
  NAND2_X1 U10378 ( .A1(n9535), .A2(n9500), .ZN(n9530) );
  NAND2_X1 U10379 ( .A1(n9530), .A2(n9501), .ZN(n9503) );
  OAI211_X1 U10380 ( .C1(n9504), .C2(n9503), .A(n9502), .B(n9629), .ZN(n9506)
         );
  NAND2_X1 U10381 ( .A1(n9506), .A2(n9505), .ZN(n9665) );
  INV_X1 U10382 ( .A(n9507), .ZN(n9510) );
  INV_X1 U10383 ( .A(n9508), .ZN(n9509) );
  AOI211_X1 U10384 ( .C1(n9667), .C2(n9510), .A(n10678), .B(n9509), .ZN(n9666)
         );
  NAND2_X1 U10385 ( .A1(n9666), .A2(n9511), .ZN(n9514) );
  AOI22_X1 U10386 ( .A1(n9512), .A2(n9616), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9618), .ZN(n9513) );
  OAI211_X1 U10387 ( .C1(n9515), .C2(n9620), .A(n9514), .B(n9513), .ZN(n9516)
         );
  AOI21_X1 U10388 ( .B1(n9665), .B2(n9517), .A(n9516), .ZN(n9518) );
  OAI21_X1 U10389 ( .B1(n9669), .B2(n9634), .A(n9518), .ZN(P2_U3271) );
  OAI21_X1 U10390 ( .B1(n9520), .B2(n9526), .A(n9519), .ZN(n9521) );
  INV_X1 U10391 ( .A(n9521), .ZN(n9674) );
  XNOR2_X1 U10392 ( .A(n9524), .B(n9541), .ZN(n9671) );
  AOI22_X1 U10393 ( .A1(n9522), .A2(n9616), .B1(n9618), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n9523) );
  OAI21_X1 U10394 ( .B1(n9524), .B2(n9620), .A(n9523), .ZN(n9533) );
  NAND2_X1 U10395 ( .A1(n9535), .A2(n9525), .ZN(n9527) );
  AOI21_X1 U10396 ( .B1(n9527), .B2(n9526), .A(n9594), .ZN(n9531) );
  OAI22_X1 U10397 ( .A1(n9528), .A2(n9599), .B1(n9558), .B2(n9597), .ZN(n9529)
         );
  AOI21_X1 U10398 ( .B1(n9531), .B2(n9530), .A(n9529), .ZN(n9673) );
  NOR2_X1 U10399 ( .A1(n9673), .A2(n9618), .ZN(n9532) );
  AOI211_X1 U10400 ( .C1(n9671), .C2(n9632), .A(n9533), .B(n9532), .ZN(n9534)
         );
  OAI21_X1 U10401 ( .B1(n9674), .B2(n9634), .A(n9534), .ZN(P2_U3272) );
  OAI21_X1 U10402 ( .B1(n4884), .B2(n9538), .A(n9535), .ZN(n9537) );
  AOI222_X1 U10403 ( .A1(n9629), .A2(n9537), .B1(n9571), .B2(n9624), .C1(n9536), .C2(n9626), .ZN(n9679) );
  INV_X1 U10404 ( .A(n9681), .ZN(n9540) );
  NAND2_X1 U10405 ( .A1(n9539), .A2(n9538), .ZN(n9675) );
  NAND3_X1 U10406 ( .A1(n9540), .A2(n9605), .A3(n9675), .ZN(n9549) );
  INV_X1 U10407 ( .A(n9551), .ZN(n9543) );
  INV_X1 U10408 ( .A(n9541), .ZN(n9542) );
  AOI21_X1 U10409 ( .B1(n9676), .B2(n9543), .A(n9542), .ZN(n9677) );
  AOI22_X1 U10410 ( .A1(n9618), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9544), .B2(
        n9616), .ZN(n9545) );
  OAI21_X1 U10411 ( .B1(n9546), .B2(n9620), .A(n9545), .ZN(n9547) );
  AOI21_X1 U10412 ( .B1(n9677), .B2(n9632), .A(n9547), .ZN(n9548) );
  OAI211_X1 U10413 ( .C1(n9618), .C2(n9679), .A(n9549), .B(n9548), .ZN(
        P2_U3273) );
  XNOR2_X1 U10414 ( .A(n9550), .B(n9555), .ZN(n9686) );
  AOI21_X1 U10415 ( .B1(n9682), .B2(n5027), .A(n9551), .ZN(n9683) );
  AOI22_X1 U10416 ( .A1(n9618), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9552), .B2(
        n9616), .ZN(n9553) );
  OAI21_X1 U10417 ( .B1(n9554), .B2(n9620), .A(n9553), .ZN(n9563) );
  AOI21_X1 U10418 ( .B1(n9556), .B2(n9555), .A(n9594), .ZN(n9561) );
  OAI22_X1 U10419 ( .A1(n9558), .A2(n9599), .B1(n9557), .B2(n9597), .ZN(n9559)
         );
  AOI21_X1 U10420 ( .B1(n9561), .B2(n9560), .A(n9559), .ZN(n9685) );
  NOR2_X1 U10421 ( .A1(n9685), .A2(n9618), .ZN(n9562) );
  AOI211_X1 U10422 ( .C1(n9683), .C2(n9632), .A(n9563), .B(n9562), .ZN(n9564)
         );
  OAI21_X1 U10423 ( .B1(n9686), .B2(n9634), .A(n9564), .ZN(P2_U3274) );
  AOI21_X1 U10424 ( .B1(n9568), .B2(n9565), .A(n4912), .ZN(n9691) );
  AOI21_X1 U10425 ( .B1(n9687), .B2(n9578), .A(n5023), .ZN(n9688) );
  AOI22_X1 U10426 ( .A1(n9618), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9566), .B2(
        n9616), .ZN(n9567) );
  OAI21_X1 U10427 ( .B1(n5026), .B2(n9620), .A(n9567), .ZN(n9574) );
  XOR2_X1 U10428 ( .A(n9569), .B(n9568), .Z(n9572) );
  AOI222_X1 U10429 ( .A1(n9629), .A2(n9572), .B1(n9571), .B2(n9626), .C1(n9570), .C2(n9624), .ZN(n9690) );
  NOR2_X1 U10430 ( .A1(n9690), .A2(n9618), .ZN(n9573) );
  AOI211_X1 U10431 ( .C1(n9688), .C2(n9632), .A(n9574), .B(n9573), .ZN(n9575)
         );
  OAI21_X1 U10432 ( .B1(n9691), .B2(n9634), .A(n9575), .ZN(P2_U3275) );
  OAI21_X1 U10433 ( .B1(n9577), .B2(n9582), .A(n9576), .ZN(n9696) );
  AOI21_X1 U10434 ( .B1(n9692), .B2(n9589), .A(n5028), .ZN(n9693) );
  AOI22_X1 U10435 ( .A1(n9618), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9579), .B2(
        n9616), .ZN(n9580) );
  OAI21_X1 U10436 ( .B1(n9581), .B2(n9620), .A(n9580), .ZN(n9587) );
  XNOR2_X1 U10437 ( .A(n9583), .B(n9582), .ZN(n9585) );
  AOI222_X1 U10438 ( .A1(n9629), .A2(n9585), .B1(n9627), .B2(n9624), .C1(n9584), .C2(n9626), .ZN(n9695) );
  NOR2_X1 U10439 ( .A1(n9695), .A2(n9618), .ZN(n9586) );
  AOI211_X1 U10440 ( .C1(n9693), .C2(n9632), .A(n9587), .B(n9586), .ZN(n9588)
         );
  OAI21_X1 U10441 ( .B1(n9696), .B2(n9634), .A(n9588), .ZN(P2_U3276) );
  INV_X1 U10442 ( .A(n9589), .ZN(n9590) );
  AOI211_X1 U10443 ( .C1(n9700), .C2(n9613), .A(n10678), .B(n9590), .ZN(n9699)
         );
  NOR2_X1 U10444 ( .A1(n9592), .A2(n9591), .ZN(n9600) );
  XNOR2_X1 U10445 ( .A(n9593), .B(n4974), .ZN(n9595) );
  OAI222_X1 U10446 ( .A1(n9599), .A2(n9598), .B1(n9597), .B2(n9596), .C1(n9595), .C2(n9594), .ZN(n9698) );
  AOI211_X1 U10447 ( .C1(n9699), .C2(n9601), .A(n9600), .B(n9698), .ZN(n9609)
         );
  OR2_X1 U10448 ( .A1(n9603), .A2(n9602), .ZN(n9697) );
  NAND3_X1 U10449 ( .A1(n9697), .A2(n9604), .A3(n9605), .ZN(n9608) );
  AOI22_X1 U10450 ( .A1(n9700), .A2(n9606), .B1(n9618), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n9607) );
  OAI211_X1 U10451 ( .C1(n9618), .C2(n9609), .A(n9608), .B(n9607), .ZN(
        P2_U3277) );
  XNOR2_X1 U10452 ( .A(n9611), .B(n9610), .ZN(n9707) );
  INV_X1 U10453 ( .A(n9612), .ZN(n9615) );
  INV_X1 U10454 ( .A(n9613), .ZN(n9614) );
  AOI21_X1 U10455 ( .B1(n9703), .B2(n9615), .A(n9614), .ZN(n9704) );
  AOI22_X1 U10456 ( .A1(n9618), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9617), .B2(
        n9616), .ZN(n9619) );
  OAI21_X1 U10457 ( .B1(n9621), .B2(n9620), .A(n9619), .ZN(n9631) );
  XNOR2_X1 U10458 ( .A(n9623), .B(n9622), .ZN(n9628) );
  AOI222_X1 U10459 ( .A1(n9629), .A2(n9628), .B1(n9627), .B2(n9626), .C1(n9625), .C2(n9624), .ZN(n9706) );
  NOR2_X1 U10460 ( .A1(n9706), .A2(n9618), .ZN(n9630) );
  AOI211_X1 U10461 ( .C1(n9704), .C2(n9632), .A(n9631), .B(n9630), .ZN(n9633)
         );
  OAI21_X1 U10462 ( .B1(n9707), .B2(n9634), .A(n9633), .ZN(P2_U3278) );
  AOI21_X1 U10463 ( .B1(n9636), .B2(n10554), .A(n9635), .ZN(n9637) );
  MUX2_X1 U10464 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9723), .S(n10685), .Z(
        P2_U3551) );
  NAND3_X1 U10465 ( .A1(n9640), .A2(n10528), .A3(n9639), .ZN(n9642) );
  OAI211_X1 U10466 ( .C1(n9643), .C2(n10676), .A(n9642), .B(n9641), .ZN(n9724)
         );
  MUX2_X1 U10467 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9724), .S(n10685), .Z(
        P2_U3550) );
  NAND2_X1 U10468 ( .A1(n9644), .A2(n10682), .ZN(n9649) );
  NAND2_X1 U10469 ( .A1(n9649), .A2(n9648), .ZN(n9725) );
  MUX2_X1 U10470 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9725), .S(n10685), .Z(
        P2_U3549) );
  AOI22_X1 U10471 ( .A1(n9651), .A2(n10528), .B1(n10554), .B2(n9650), .ZN(
        n9652) );
  OAI211_X1 U10472 ( .C1(n9654), .C2(n10666), .A(n9653), .B(n9652), .ZN(n9726)
         );
  MUX2_X1 U10473 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9726), .S(n10685), .Z(
        P2_U3548) );
  AOI22_X1 U10474 ( .A1(n9656), .A2(n10528), .B1(n10554), .B2(n9655), .ZN(
        n9657) );
  OAI211_X1 U10475 ( .C1(n9659), .C2(n10666), .A(n9658), .B(n9657), .ZN(n9727)
         );
  MUX2_X1 U10476 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9727), .S(n10685), .Z(
        P2_U3547) );
  AOI21_X1 U10477 ( .B1(n10554), .B2(n9661), .A(n9660), .ZN(n9662) );
  OAI211_X1 U10478 ( .C1(n9664), .C2(n10666), .A(n9663), .B(n9662), .ZN(n9728)
         );
  MUX2_X1 U10479 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9728), .S(n10685), .Z(
        P2_U3546) );
  AOI211_X1 U10480 ( .C1(n10554), .C2(n9667), .A(n9666), .B(n9665), .ZN(n9668)
         );
  OAI21_X1 U10481 ( .B1(n9669), .B2(n10666), .A(n9668), .ZN(n9729) );
  MUX2_X1 U10482 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9729), .S(n10685), .Z(
        P2_U3545) );
  AOI22_X1 U10483 ( .A1(n9671), .A2(n10528), .B1(n10554), .B2(n9670), .ZN(
        n9672) );
  OAI211_X1 U10484 ( .C1(n9674), .C2(n10666), .A(n9673), .B(n9672), .ZN(n9730)
         );
  MUX2_X1 U10485 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9730), .S(n10685), .Z(
        P2_U3544) );
  NAND2_X1 U10486 ( .A1(n9675), .A2(n10682), .ZN(n9680) );
  AOI22_X1 U10487 ( .A1(n9677), .A2(n10528), .B1(n10554), .B2(n9676), .ZN(
        n9678) );
  OAI211_X1 U10488 ( .C1(n9681), .C2(n9680), .A(n9679), .B(n9678), .ZN(n9731)
         );
  MUX2_X1 U10489 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9731), .S(n10685), .Z(
        P2_U3543) );
  AOI22_X1 U10490 ( .A1(n9683), .A2(n10528), .B1(n10554), .B2(n9682), .ZN(
        n9684) );
  OAI211_X1 U10491 ( .C1(n9686), .C2(n10666), .A(n9685), .B(n9684), .ZN(n9732)
         );
  MUX2_X1 U10492 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9732), .S(n10685), .Z(
        P2_U3542) );
  AOI22_X1 U10493 ( .A1(n9688), .A2(n10528), .B1(n10554), .B2(n9687), .ZN(
        n9689) );
  OAI211_X1 U10494 ( .C1(n9691), .C2(n10666), .A(n9690), .B(n9689), .ZN(n9733)
         );
  MUX2_X1 U10495 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9733), .S(n10685), .Z(
        P2_U3541) );
  AOI22_X1 U10496 ( .A1(n9693), .A2(n10528), .B1(n10554), .B2(n9692), .ZN(
        n9694) );
  OAI211_X1 U10497 ( .C1(n9696), .C2(n10666), .A(n9695), .B(n9694), .ZN(n9734)
         );
  MUX2_X1 U10498 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9734), .S(n10685), .Z(
        P2_U3540) );
  NAND3_X1 U10499 ( .A1(n9697), .A2(n9604), .A3(n10682), .ZN(n9702) );
  AOI211_X1 U10500 ( .C1(n10554), .C2(n9700), .A(n9699), .B(n9698), .ZN(n9701)
         );
  NAND2_X1 U10501 ( .A1(n9702), .A2(n9701), .ZN(n9735) );
  MUX2_X1 U10502 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9735), .S(n10685), .Z(
        P2_U3539) );
  AOI22_X1 U10503 ( .A1(n9704), .A2(n10528), .B1(n10554), .B2(n9703), .ZN(
        n9705) );
  OAI211_X1 U10504 ( .C1(n9707), .C2(n10666), .A(n9706), .B(n9705), .ZN(n9736)
         );
  MUX2_X1 U10505 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9736), .S(n10685), .Z(
        P2_U3538) );
  AOI211_X1 U10506 ( .C1(n10554), .C2(n9710), .A(n9709), .B(n9708), .ZN(n9711)
         );
  OAI21_X1 U10507 ( .B1(n9712), .B2(n10666), .A(n9711), .ZN(n9737) );
  MUX2_X1 U10508 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9737), .S(n10685), .Z(
        P2_U3537) );
  AOI21_X1 U10509 ( .B1(n10554), .B2(n9714), .A(n9713), .ZN(n9715) );
  OAI211_X1 U10510 ( .C1(n9717), .C2(n10666), .A(n9716), .B(n9715), .ZN(n9738)
         );
  MUX2_X1 U10511 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9738), .S(n10685), .Z(
        P2_U3536) );
  AOI22_X1 U10512 ( .A1(n9719), .A2(n10528), .B1(n10554), .B2(n9718), .ZN(
        n9720) );
  OAI211_X1 U10513 ( .C1(n9722), .C2(n10666), .A(n9721), .B(n9720), .ZN(n9739)
         );
  MUX2_X1 U10514 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9739), .S(n10685), .Z(
        P2_U3535) );
  MUX2_X1 U10515 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9724), .S(n10689), .Z(
        P2_U3518) );
  MUX2_X1 U10516 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9725), .S(n10689), .Z(
        P2_U3517) );
  MUX2_X1 U10517 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9726), .S(n10689), .Z(
        P2_U3516) );
  MUX2_X1 U10518 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9727), .S(n10689), .Z(
        P2_U3515) );
  MUX2_X1 U10519 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9728), .S(n10689), .Z(
        P2_U3514) );
  MUX2_X1 U10520 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9729), .S(n10689), .Z(
        P2_U3513) );
  MUX2_X1 U10521 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9730), .S(n10689), .Z(
        P2_U3512) );
  MUX2_X1 U10522 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9731), .S(n10689), .Z(
        P2_U3511) );
  MUX2_X1 U10523 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9732), .S(n10689), .Z(
        P2_U3510) );
  MUX2_X1 U10524 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9733), .S(n10689), .Z(
        P2_U3509) );
  MUX2_X1 U10525 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9734), .S(n10689), .Z(
        P2_U3508) );
  MUX2_X1 U10526 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9735), .S(n10689), .Z(
        P2_U3507) );
  MUX2_X1 U10527 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9736), .S(n10689), .Z(
        P2_U3505) );
  MUX2_X1 U10528 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9737), .S(n10689), .Z(
        P2_U3502) );
  MUX2_X1 U10529 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9738), .S(n10689), .Z(
        P2_U3499) );
  MUX2_X1 U10530 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9739), .S(n10689), .Z(
        P2_U3496) );
  NAND2_X1 U10531 ( .A1(n10290), .A2(n9740), .ZN(n9744) );
  NAND2_X1 U10532 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_STATE_REG_SCAN_IN), 
        .ZN(n9741) );
  OR3_X1 U10533 ( .A1(n9742), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9741), .ZN(
        n9743) );
  OAI211_X1 U10534 ( .C1(n6630), .C2(n4858), .A(n9744), .B(n9743), .ZN(
        P2_U3327) );
  MUX2_X1 U10535 ( .A(n9745), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10536 ( .A1(n9746), .A2(n9747), .ZN(n9748) );
  XOR2_X1 U10537 ( .A(n9749), .B(n9748), .Z(n9757) );
  NAND2_X1 U10538 ( .A1(n9806), .A2(n9750), .ZN(n9753) );
  AOI21_X1 U10539 ( .B1(n9853), .B2(n9889), .A(n9751), .ZN(n9752) );
  OAI211_X1 U10540 ( .C1(n9754), .C2(n9851), .A(n9753), .B(n9752), .ZN(n9755)
         );
  AOI21_X1 U10541 ( .B1(n10257), .B2(n9863), .A(n9755), .ZN(n9756) );
  OAI21_X1 U10542 ( .B1(n9757), .B2(n9879), .A(n9756), .ZN(P1_U3213) );
  NAND2_X1 U10543 ( .A1(n9758), .A2(n9759), .ZN(n9761) );
  XNOR2_X1 U10544 ( .A(n9761), .B(n9760), .ZN(n9766) );
  AOI22_X1 U10545 ( .A1(n9853), .A2(n10054), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9763) );
  NAND2_X1 U10546 ( .A1(n9873), .A2(n10055), .ZN(n9762) );
  OAI211_X1 U10547 ( .C1(n9876), .C2(n10059), .A(n9763), .B(n9762), .ZN(n9764)
         );
  AOI21_X1 U10548 ( .B1(n10205), .B2(n9863), .A(n9764), .ZN(n9765) );
  OAI21_X1 U10549 ( .B1(n9766), .B2(n9879), .A(n9765), .ZN(P1_U3214) );
  XOR2_X1 U10550 ( .A(n9768), .B(n9767), .Z(n9769) );
  XNOR2_X1 U10551 ( .A(n9770), .B(n9769), .ZN(n9775) );
  NOR2_X1 U10552 ( .A1(n9876), .A2(n10126), .ZN(n9773) );
  NAND2_X1 U10553 ( .A1(n10122), .A2(n9853), .ZN(n9771) );
  NAND2_X1 U10554 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9938) );
  OAI211_X1 U10555 ( .C1(n9851), .C2(n9818), .A(n9771), .B(n9938), .ZN(n9772)
         );
  AOI211_X1 U10556 ( .C1(n10226), .C2(n9863), .A(n9773), .B(n9772), .ZN(n9774)
         );
  OAI21_X1 U10557 ( .B1(n9775), .B2(n9879), .A(n9774), .ZN(P1_U3217) );
  NOR2_X1 U10558 ( .A1(n5243), .A2(n9778), .ZN(n9779) );
  XNOR2_X1 U10559 ( .A(n9776), .B(n9779), .ZN(n9785) );
  NAND2_X1 U10560 ( .A1(n9806), .A2(n10092), .ZN(n9781) );
  AOI22_X1 U10561 ( .A1(n9853), .A2(n10055), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9780) );
  OAI211_X1 U10562 ( .C1(n9782), .C2(n9851), .A(n9781), .B(n9780), .ZN(n9783)
         );
  AOI21_X1 U10563 ( .B1(n10217), .B2(n9863), .A(n9783), .ZN(n9784) );
  OAI21_X1 U10564 ( .B1(n9785), .B2(n9879), .A(n9784), .ZN(P1_U3221) );
  NAND2_X1 U10565 ( .A1(n9787), .A2(n9786), .ZN(n9791) );
  XNOR2_X1 U10566 ( .A(n9789), .B(n9788), .ZN(n9790) );
  XNOR2_X1 U10567 ( .A(n9791), .B(n9790), .ZN(n9796) );
  AOI22_X1 U10568 ( .A1(n9853), .A2(n9885), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9793) );
  NAND2_X1 U10569 ( .A1(n9873), .A2(n10054), .ZN(n9792) );
  OAI211_X1 U10570 ( .C1(n9876), .C2(n10018), .A(n9793), .B(n9792), .ZN(n9794)
         );
  AOI21_X1 U10571 ( .B1(n10196), .B2(n9863), .A(n9794), .ZN(n9795) );
  OAI21_X1 U10572 ( .B1(n9796), .B2(n9879), .A(n9795), .ZN(P1_U3223) );
  INV_X1 U10573 ( .A(n9797), .ZN(n9798) );
  AOI21_X1 U10574 ( .B1(n9800), .B2(n9799), .A(n9798), .ZN(n9809) );
  NAND2_X1 U10575 ( .A1(n9873), .A2(n9889), .ZN(n9802) );
  OAI211_X1 U10576 ( .C1(n10150), .C2(n9871), .A(n9802), .B(n9801), .ZN(n9805)
         );
  NOR2_X1 U10577 ( .A1(n9803), .A2(n9824), .ZN(n9804) );
  AOI211_X1 U10578 ( .C1(n9807), .C2(n9806), .A(n9805), .B(n9804), .ZN(n9808)
         );
  OAI21_X1 U10579 ( .B1(n9809), .B2(n9879), .A(n9808), .ZN(P1_U3224) );
  INV_X1 U10580 ( .A(n9814), .ZN(n9811) );
  NOR2_X1 U10581 ( .A1(n9810), .A2(n9811), .ZN(n9817) );
  AOI21_X1 U10582 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9816) );
  OAI21_X1 U10583 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9823) );
  NAND2_X1 U10584 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9901) );
  OAI21_X1 U10585 ( .B1(n9871), .B2(n9818), .A(n9901), .ZN(n9821) );
  NOR2_X1 U10586 ( .A1(n9876), .A2(n9819), .ZN(n9820) );
  AOI211_X1 U10587 ( .C1(n9873), .C2(n9888), .A(n9821), .B(n9820), .ZN(n9822)
         );
  OAI211_X1 U10588 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9822), .ZN(
        P1_U3226) );
  XOR2_X1 U10589 ( .A(n9826), .B(n8999), .Z(n9831) );
  AOI22_X1 U10590 ( .A1(n9853), .A2(n10038), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9828) );
  NAND2_X1 U10591 ( .A1(n9873), .A2(n10037), .ZN(n9827) );
  OAI211_X1 U10592 ( .C1(n9876), .C2(n10044), .A(n9828), .B(n9827), .ZN(n9829)
         );
  AOI21_X1 U10593 ( .B1(n10201), .B2(n9863), .A(n9829), .ZN(n9830) );
  OAI21_X1 U10594 ( .B1(n9831), .B2(n9879), .A(n9830), .ZN(P1_U3227) );
  NAND2_X1 U10595 ( .A1(n9833), .A2(n9832), .ZN(n9835) );
  XOR2_X1 U10596 ( .A(n9835), .B(n9834), .Z(n9840) );
  AOI22_X1 U10597 ( .A1(n9886), .A2(n9853), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9837) );
  NAND2_X1 U10598 ( .A1(n9873), .A2(n10147), .ZN(n9836) );
  OAI211_X1 U10599 ( .C1(n9876), .C2(n10103), .A(n9837), .B(n9836), .ZN(n9838)
         );
  AOI21_X1 U10600 ( .B1(n10222), .B2(n9863), .A(n9838), .ZN(n9839) );
  OAI21_X1 U10601 ( .B1(n9840), .B2(n9879), .A(n9839), .ZN(P1_U3231) );
  NAND2_X1 U10602 ( .A1(n9843), .A2(n9842), .ZN(n9844) );
  XNOR2_X1 U10603 ( .A(n9841), .B(n9844), .ZN(n9849) );
  NAND2_X1 U10604 ( .A1(n9886), .A2(n9873), .ZN(n9846) );
  AOI22_X1 U10605 ( .A1(n9853), .A2(n10037), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9845) );
  OAI211_X1 U10606 ( .C1(n9876), .C2(n10071), .A(n9846), .B(n9845), .ZN(n9847)
         );
  AOI21_X1 U10607 ( .B1(n10211), .B2(n9863), .A(n9847), .ZN(n9848) );
  OAI21_X1 U10608 ( .B1(n9849), .B2(n9879), .A(n9848), .ZN(P1_U3233) );
  NOR2_X1 U10609 ( .A1(n9850), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9925) );
  NOR2_X1 U10610 ( .A1(n9851), .A2(n10150), .ZN(n9852) );
  AOI211_X1 U10611 ( .C1(n9853), .C2(n10147), .A(n9925), .B(n9852), .ZN(n9854)
         );
  OAI21_X1 U10612 ( .B1(n9876), .B2(n10161), .A(n9854), .ZN(n9862) );
  INV_X1 U10613 ( .A(n9855), .ZN(n9860) );
  AOI21_X1 U10614 ( .B1(n9859), .B2(n9857), .A(n9856), .ZN(n9858) );
  AOI211_X1 U10615 ( .C1(n9860), .C2(n9859), .A(n9879), .B(n9858), .ZN(n9861)
         );
  AOI211_X1 U10616 ( .C1(n10231), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9864)
         );
  INV_X1 U10617 ( .A(n9864), .ZN(P1_U3236) );
  XNOR2_X1 U10618 ( .A(n9867), .B(n9866), .ZN(n9868) );
  XNOR2_X1 U10619 ( .A(n9865), .B(n9868), .ZN(n9880) );
  OAI21_X1 U10620 ( .B1(n9871), .B2(n9870), .A(n9869), .ZN(n9872) );
  AOI21_X1 U10621 ( .B1(n9873), .B2(n9890), .A(n9872), .ZN(n9874) );
  OAI21_X1 U10622 ( .B1(n9876), .B2(n9875), .A(n9874), .ZN(n9877) );
  AOI21_X1 U10623 ( .B1(n10249), .B2(n9863), .A(n9877), .ZN(n9878) );
  OAI21_X1 U10624 ( .B1(n9880), .B2(n9879), .A(n9878), .ZN(P1_U3239) );
  MUX2_X1 U10625 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9881), .S(n4857), .Z(
        P1_U3585) );
  MUX2_X1 U10626 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9882), .S(n4857), .Z(
        P1_U3584) );
  MUX2_X1 U10627 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9883), .S(n4857), .Z(
        P1_U3583) );
  MUX2_X1 U10628 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9884), .S(n4857), .Z(
        P1_U3582) );
  MUX2_X1 U10629 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9885), .S(n4857), .Z(
        P1_U3581) );
  MUX2_X1 U10630 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10038), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10631 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10054), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10632 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10055), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10633 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9886), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10634 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10122), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10635 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10147), .S(n4857), .Z(
        P1_U3574) );
  MUX2_X1 U10636 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10121), .S(n4857), .Z(
        P1_U3573) );
  MUX2_X1 U10637 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9887), .S(n4857), .Z(
        P1_U3572) );
  MUX2_X1 U10638 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9888), .S(n4857), .Z(
        P1_U3571) );
  MUX2_X1 U10639 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9889), .S(n4857), .Z(
        P1_U3570) );
  MUX2_X1 U10640 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9890), .S(n4857), .Z(
        P1_U3569) );
  MUX2_X1 U10641 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9891), .S(n4857), .Z(
        P1_U3568) );
  MUX2_X1 U10642 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9892), .S(n4857), .Z(
        P1_U3567) );
  MUX2_X1 U10643 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9893), .S(n4857), .Z(
        P1_U3566) );
  MUX2_X1 U10644 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9894), .S(n4857), .Z(
        P1_U3565) );
  MUX2_X1 U10645 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9895), .S(n4857), .Z(
        P1_U3564) );
  MUX2_X1 U10646 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9896), .S(n4857), .Z(
        P1_U3563) );
  MUX2_X1 U10647 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9897), .S(n4857), .Z(
        P1_U3562) );
  MUX2_X1 U10648 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9898), .S(n4857), .Z(
        P1_U3561) );
  MUX2_X1 U10649 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9899), .S(n4857), .Z(
        P1_U3560) );
  MUX2_X1 U10650 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9900), .S(n4857), .Z(
        P1_U3559) );
  MUX2_X1 U10651 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n6892), .S(n4857), .Z(
        P1_U3558) );
  MUX2_X1 U10652 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6914), .S(n4857), .Z(
        P1_U3557) );
  MUX2_X1 U10653 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6902), .S(n4857), .Z(
        P1_U3556) );
  MUX2_X1 U10654 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6712), .S(n4857), .Z(
        P1_U3555) );
  INV_X1 U10655 ( .A(n9901), .ZN(n9906) );
  AOI21_X1 U10656 ( .B1(n9908), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9902), .ZN(
        n9904) );
  XNOR2_X1 U10657 ( .A(n9919), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9903) );
  NOR2_X1 U10658 ( .A1(n9904), .A2(n9903), .ZN(n9915) );
  AOI211_X1 U10659 ( .C1(n9904), .C2(n9903), .A(n9915), .B(n10395), .ZN(n9905)
         );
  AOI211_X1 U10660 ( .C1(n9919), .C2(n10406), .A(n9906), .B(n9905), .ZN(n9914)
         );
  AOI21_X1 U10661 ( .B1(n9908), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9907), .ZN(
        n9911) );
  NAND2_X1 U10662 ( .A1(n9919), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9909) );
  OAI21_X1 U10663 ( .B1(n9919), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9909), .ZN(
        n9910) );
  NOR2_X1 U10664 ( .A1(n9911), .A2(n9910), .ZN(n9918) );
  AOI211_X1 U10665 ( .C1(n9911), .C2(n9910), .A(n9918), .B(n10412), .ZN(n9912)
         );
  AOI21_X1 U10666 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n10407), .A(n9912), .ZN(
        n9913) );
  NAND2_X1 U10667 ( .A1(n9914), .A2(n9913), .ZN(P1_U3258) );
  INV_X1 U10668 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9928) );
  XOR2_X1 U10669 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9935), .Z(n9917) );
  AOI21_X1 U10670 ( .B1(n9919), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9915), .ZN(
        n9916) );
  NAND2_X1 U10671 ( .A1(n9916), .A2(n9917), .ZN(n9934) );
  OAI21_X1 U10672 ( .B1(n9917), .B2(n9916), .A(n9934), .ZN(n9924) );
  AOI21_X1 U10673 ( .B1(n9919), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9918), .ZN(
        n9922) );
  NAND2_X1 U10674 ( .A1(n9935), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9920) );
  OAI21_X1 U10675 ( .B1(n9935), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9920), .ZN(
        n9921) );
  NOR2_X1 U10676 ( .A1(n9922), .A2(n9921), .ZN(n9930) );
  AOI211_X1 U10677 ( .C1(n9922), .C2(n9921), .A(n9930), .B(n10412), .ZN(n9923)
         );
  AOI21_X1 U10678 ( .B1(n10414), .B2(n9924), .A(n9923), .ZN(n9927) );
  AOI21_X1 U10679 ( .B1(n10406), .B2(n9935), .A(n9925), .ZN(n9926) );
  OAI211_X1 U10680 ( .C1(n9929), .C2(n9928), .A(n9927), .B(n9926), .ZN(
        P1_U3259) );
  MUX2_X1 U10681 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n5716), .S(n9944), .Z(n9932) );
  AOI21_X1 U10682 ( .B1(n9935), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9930), .ZN(
        n9931) );
  XOR2_X1 U10683 ( .A(n9932), .B(n9931), .Z(n9933) );
  AOI22_X1 U10684 ( .A1(n10407), .A2(P1_ADDR_REG_19__SCAN_IN), .B1(n10398), 
        .B2(n9933), .ZN(n9942) );
  OAI21_X1 U10685 ( .B1(n9935), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9934), .ZN(
        n9937) );
  XNOR2_X1 U10686 ( .A(n9944), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9936) );
  XNOR2_X1 U10687 ( .A(n9937), .B(n9936), .ZN(n9940) );
  INV_X1 U10688 ( .A(n9938), .ZN(n9939) );
  AOI21_X1 U10689 ( .B1(n10414), .B2(n9940), .A(n9939), .ZN(n9941) );
  OAI211_X1 U10690 ( .C1(n9944), .C2(n9943), .A(n9942), .B(n9941), .ZN(
        P1_U3260) );
  NAND2_X1 U10691 ( .A1(n9954), .A2(n9953), .ZN(n9945) );
  XNOR2_X1 U10692 ( .A(n9952), .B(n9945), .ZN(n10171) );
  NAND2_X1 U10693 ( .A1(n10171), .A2(n10137), .ZN(n9951) );
  NAND2_X1 U10694 ( .A1(n9947), .A2(n9946), .ZN(n9948) );
  NOR2_X1 U10695 ( .A1(n10111), .A2(n9948), .ZN(n10175) );
  INV_X1 U10696 ( .A(n10175), .ZN(n9949) );
  NOR2_X1 U10697 ( .A1(n9949), .A2(n4856), .ZN(n9956) );
  AOI21_X1 U10698 ( .B1(n4856), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9956), .ZN(
        n9950) );
  OAI211_X1 U10699 ( .C1(n9952), .C2(n10130), .A(n9951), .B(n9950), .ZN(
        P1_U3261) );
  XNOR2_X1 U10700 ( .A(n9954), .B(n9953), .ZN(n10178) );
  NOR2_X1 U10701 ( .A1(n9954), .A2(n10130), .ZN(n9955) );
  AOI211_X1 U10702 ( .C1(n4856), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9956), .B(
        n9955), .ZN(n9957) );
  OAI21_X1 U10703 ( .B1(n10167), .B2(n10178), .A(n9957), .ZN(P1_U3262) );
  AOI211_X1 U10704 ( .C1(n9960), .C2(n9959), .A(n10107), .B(n9958), .ZN(n9963)
         );
  OAI22_X1 U10705 ( .A1(n9961), .A2(n10111), .B1(n10149), .B2(n9998), .ZN(
        n9962) );
  NOR2_X1 U10706 ( .A1(n9963), .A2(n9962), .ZN(n10184) );
  INV_X1 U10707 ( .A(n10179), .ZN(n9974) );
  AND2_X1 U10708 ( .A1(n9978), .A2(n10179), .ZN(n9968) );
  NOR2_X1 U10709 ( .A1(n9969), .A2(n9968), .ZN(n10180) );
  NAND2_X1 U10710 ( .A1(n10180), .A2(n10137), .ZN(n9973) );
  INV_X1 U10711 ( .A(n9970), .ZN(n9971) );
  AOI22_X1 U10712 ( .A1(n4856), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n10128), 
        .B2(n9971), .ZN(n9972) );
  OAI211_X1 U10713 ( .C1(n9974), .C2(n10130), .A(n9973), .B(n9972), .ZN(n9975)
         );
  AOI21_X1 U10714 ( .B1(n10181), .B2(n10050), .A(n9975), .ZN(n9976) );
  OAI21_X1 U10715 ( .B1(n10184), .B2(n4856), .A(n9976), .ZN(P1_U3263) );
  XNOR2_X1 U10716 ( .A(n9977), .B(n9986), .ZN(n10188) );
  INV_X1 U10717 ( .A(n10003), .ZN(n9980) );
  INV_X1 U10718 ( .A(n9978), .ZN(n9979) );
  AOI211_X1 U10719 ( .C1(n5955), .C2(n9980), .A(n10633), .B(n9979), .ZN(n10185) );
  INV_X1 U10720 ( .A(n9981), .ZN(n9982) );
  AOI22_X1 U10721 ( .A1(n4856), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10128), 
        .B2(n9982), .ZN(n9983) );
  OAI21_X1 U10722 ( .B1(n9984), .B2(n10130), .A(n9983), .ZN(n9991) );
  AOI211_X1 U10723 ( .C1(n9986), .C2(n9985), .A(n10107), .B(n4885), .ZN(n9989)
         );
  OAI22_X1 U10724 ( .A1(n9987), .A2(n10111), .B1(n10149), .B2(n10026), .ZN(
        n9988) );
  NOR2_X1 U10725 ( .A1(n9989), .A2(n9988), .ZN(n10187) );
  NOR2_X1 U10726 ( .A1(n10187), .A2(n4856), .ZN(n9990) );
  AOI211_X1 U10727 ( .C1(n10185), .C2(n10117), .A(n9991), .B(n9990), .ZN(n9992) );
  OAI21_X1 U10728 ( .B1(n10134), .B2(n10188), .A(n9992), .ZN(P1_U3264) );
  OAI21_X1 U10729 ( .B1(n9995), .B2(n9994), .A(n9993), .ZN(n10001) );
  XNOR2_X2 U10730 ( .A(n9996), .B(n9995), .ZN(n10194) );
  OAI22_X1 U10731 ( .A1(n9998), .A2(n10111), .B1(n10149), .B2(n9997), .ZN(
        n9999) );
  AOI211_X2 U10732 ( .C1(n10001), .C2(n10152), .A(n10000), .B(n9999), .ZN(
        n10193) );
  INV_X1 U10733 ( .A(n10194), .ZN(n10010) );
  AND2_X1 U10734 ( .A1(n10007), .A2(n10016), .ZN(n10002) );
  OR2_X1 U10735 ( .A1(n10003), .A2(n10002), .ZN(n10190) );
  OAI22_X1 U10736 ( .A1(n10163), .A2(n10005), .B1(n10004), .B2(n10160), .ZN(
        n10006) );
  AOI21_X1 U10737 ( .B1(n10007), .B2(n10165), .A(n10006), .ZN(n10008) );
  OAI21_X1 U10738 ( .B1(n10190), .B2(n10167), .A(n10008), .ZN(n10009) );
  AOI21_X1 U10739 ( .B1(n10010), .B2(n10169), .A(n10009), .ZN(n10011) );
  OAI21_X1 U10740 ( .B1(n10193), .B2(n4856), .A(n10011), .ZN(P1_U3265) );
  INV_X1 U10741 ( .A(n10012), .ZN(n10013) );
  AOI21_X1 U10742 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(n10199) );
  INV_X1 U10743 ( .A(n10016), .ZN(n10017) );
  AOI211_X1 U10744 ( .C1(n10196), .C2(n10042), .A(n10633), .B(n10017), .ZN(
        n10195) );
  INV_X1 U10745 ( .A(n10196), .ZN(n10021) );
  INV_X1 U10746 ( .A(n10018), .ZN(n10019) );
  AOI22_X1 U10747 ( .A1(n4856), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10128), 
        .B2(n10019), .ZN(n10020) );
  OAI21_X1 U10748 ( .B1(n10021), .B2(n10130), .A(n10020), .ZN(n10030) );
  AOI211_X1 U10749 ( .C1(n10024), .C2(n10023), .A(n10107), .B(n10022), .ZN(
        n10028) );
  OAI22_X1 U10750 ( .A1(n10026), .A2(n10111), .B1(n10149), .B2(n10025), .ZN(
        n10027) );
  NOR2_X1 U10751 ( .A1(n10028), .A2(n10027), .ZN(n10198) );
  NOR2_X1 U10752 ( .A1(n10198), .A2(n4856), .ZN(n10029) );
  AOI211_X1 U10753 ( .C1(n10195), .C2(n10117), .A(n10030), .B(n10029), .ZN(
        n10031) );
  OAI21_X1 U10754 ( .B1(n10199), .B2(n10134), .A(n10031), .ZN(P1_U3266) );
  INV_X1 U10755 ( .A(n10032), .ZN(n10033) );
  NOR2_X1 U10756 ( .A1(n10034), .A2(n10033), .ZN(n10036) );
  XNOR2_X1 U10757 ( .A(n10036), .B(n10035), .ZN(n10039) );
  AOI222_X1 U10758 ( .A1(n10152), .A2(n10039), .B1(n10038), .B2(n10146), .C1(
        n10037), .C2(n10120), .ZN(n10203) );
  OAI21_X1 U10759 ( .B1(n4872), .B2(n5952), .A(n10040), .ZN(n10204) );
  INV_X1 U10760 ( .A(n10204), .ZN(n10051) );
  INV_X1 U10761 ( .A(n10058), .ZN(n10041) );
  AOI21_X1 U10762 ( .B1(n10041), .B2(n10201), .A(n10633), .ZN(n10043) );
  AND2_X1 U10763 ( .A1(n10043), .A2(n10042), .ZN(n10200) );
  NAND2_X1 U10764 ( .A1(n10200), .A2(n10117), .ZN(n10047) );
  INV_X1 U10765 ( .A(n10044), .ZN(n10045) );
  AOI22_X1 U10766 ( .A1(n4856), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n10128), 
        .B2(n10045), .ZN(n10046) );
  OAI211_X1 U10767 ( .C1(n10048), .C2(n10130), .A(n10047), .B(n10046), .ZN(
        n10049) );
  AOI21_X1 U10768 ( .B1(n10051), .B2(n10050), .A(n10049), .ZN(n10052) );
  OAI21_X1 U10769 ( .B1(n10203), .B2(n4856), .A(n10052), .ZN(P1_U3267) );
  XNOR2_X1 U10770 ( .A(n10053), .B(n10063), .ZN(n10056) );
  AOI222_X1 U10771 ( .A1(n10152), .A2(n10056), .B1(n10055), .B2(n10120), .C1(
        n10054), .C2(n10146), .ZN(n10208) );
  AND2_X1 U10772 ( .A1(n10205), .A2(n10069), .ZN(n10057) );
  NOR2_X1 U10773 ( .A1(n10058), .A2(n10057), .ZN(n10206) );
  INV_X1 U10774 ( .A(n10205), .ZN(n10062) );
  INV_X1 U10775 ( .A(n10059), .ZN(n10060) );
  AOI22_X1 U10776 ( .A1(n4856), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10128), 
        .B2(n10060), .ZN(n10061) );
  OAI21_X1 U10777 ( .B1(n10062), .B2(n10130), .A(n10061), .ZN(n10066) );
  XOR2_X1 U10778 ( .A(n10064), .B(n10063), .Z(n10209) );
  NOR2_X1 U10779 ( .A1(n10209), .A2(n10134), .ZN(n10065) );
  AOI211_X1 U10780 ( .C1(n10206), .C2(n10137), .A(n10066), .B(n10065), .ZN(
        n10067) );
  OAI21_X1 U10781 ( .B1(n10208), .B2(n4856), .A(n10067), .ZN(P1_U3268) );
  XNOR2_X1 U10782 ( .A(n10068), .B(n10076), .ZN(n10214) );
  INV_X1 U10783 ( .A(n10069), .ZN(n10070) );
  AOI211_X1 U10784 ( .C1(n10211), .C2(n10084), .A(n10633), .B(n10070), .ZN(
        n10210) );
  INV_X1 U10785 ( .A(n10071), .ZN(n10072) );
  AOI22_X1 U10786 ( .A1(n4856), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10128), 
        .B2(n10072), .ZN(n10073) );
  OAI21_X1 U10787 ( .B1(n5167), .B2(n10130), .A(n10073), .ZN(n10081) );
  AOI211_X1 U10788 ( .C1(n10076), .C2(n10075), .A(n10107), .B(n10074), .ZN(
        n10079) );
  OAI22_X1 U10789 ( .A1(n10112), .A2(n10149), .B1(n10077), .B2(n10111), .ZN(
        n10078) );
  NOR2_X1 U10790 ( .A1(n10079), .A2(n10078), .ZN(n10213) );
  NOR2_X1 U10791 ( .A1(n10213), .A2(n4856), .ZN(n10080) );
  AOI211_X1 U10792 ( .C1(n10210), .C2(n10117), .A(n10081), .B(n10080), .ZN(
        n10082) );
  OAI21_X1 U10793 ( .B1(n10134), .B2(n10214), .A(n10082), .ZN(P1_U3269) );
  XNOR2_X1 U10794 ( .A(n10083), .B(n10088), .ZN(n10220) );
  AOI211_X1 U10795 ( .C1(n10217), .C2(n10100), .A(n10633), .B(n5168), .ZN(
        n10215) );
  INV_X1 U10796 ( .A(n10215), .ZN(n10094) );
  INV_X1 U10797 ( .A(n10085), .ZN(n10087) );
  NAND2_X1 U10798 ( .A1(n10087), .A2(n10086), .ZN(n10089) );
  XNOR2_X1 U10799 ( .A(n10089), .B(n10088), .ZN(n10090) );
  AOI22_X1 U10800 ( .A1(n10090), .A2(n10152), .B1(n10120), .B2(n10122), .ZN(
        n10219) );
  NOR2_X1 U10801 ( .A1(n10111), .A2(n10091), .ZN(n10216) );
  AOI21_X1 U10802 ( .B1(n10092), .B2(n10128), .A(n10216), .ZN(n10093) );
  OAI211_X1 U10803 ( .C1(n10095), .C2(n10094), .A(n10219), .B(n10093), .ZN(
        n10096) );
  NAND2_X1 U10804 ( .A1(n10096), .A2(n10163), .ZN(n10098) );
  AOI22_X1 U10805 ( .A1(n10217), .A2(n10165), .B1(n4856), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n10097) );
  OAI211_X1 U10806 ( .C1(n10220), .C2(n10134), .A(n10098), .B(n10097), .ZN(
        P1_U3270) );
  XNOR2_X1 U10807 ( .A(n10099), .B(n10109), .ZN(n10225) );
  INV_X1 U10808 ( .A(n10125), .ZN(n10102) );
  INV_X1 U10809 ( .A(n10100), .ZN(n10101) );
  AOI211_X1 U10810 ( .C1(n10222), .C2(n10102), .A(n10633), .B(n10101), .ZN(
        n10221) );
  INV_X1 U10811 ( .A(n10103), .ZN(n10104) );
  AOI22_X1 U10812 ( .A1(n10104), .A2(n10128), .B1(n4856), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n10105) );
  OAI21_X1 U10813 ( .B1(n10106), .B2(n10130), .A(n10105), .ZN(n10116) );
  AOI211_X1 U10814 ( .C1(n10109), .C2(n10108), .A(n10107), .B(n10085), .ZN(
        n10114) );
  OAI22_X1 U10815 ( .A1(n10112), .A2(n10111), .B1(n10110), .B2(n10149), .ZN(
        n10113) );
  NOR2_X1 U10816 ( .A1(n10114), .A2(n10113), .ZN(n10224) );
  NOR2_X1 U10817 ( .A1(n10224), .A2(n4856), .ZN(n10115) );
  AOI211_X1 U10818 ( .C1(n10221), .C2(n10117), .A(n10116), .B(n10115), .ZN(
        n10118) );
  OAI21_X1 U10819 ( .B1(n10134), .B2(n10225), .A(n10118), .ZN(P1_U3271) );
  XNOR2_X1 U10820 ( .A(n10119), .B(n10132), .ZN(n10123) );
  AOI222_X1 U10821 ( .A1(n10152), .A2(n10123), .B1(n10122), .B2(n10146), .C1(
        n10121), .C2(n10120), .ZN(n10229) );
  AND2_X1 U10822 ( .A1(n10226), .A2(n10159), .ZN(n10124) );
  NOR2_X1 U10823 ( .A1(n10125), .A2(n10124), .ZN(n10227) );
  INV_X1 U10824 ( .A(n10226), .ZN(n10131) );
  INV_X1 U10825 ( .A(n10126), .ZN(n10127) );
  AOI22_X1 U10826 ( .A1(n4856), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10128), 
        .B2(n10127), .ZN(n10129) );
  OAI21_X1 U10827 ( .B1(n10131), .B2(n10130), .A(n10129), .ZN(n10136) );
  XNOR2_X1 U10828 ( .A(n10133), .B(n10132), .ZN(n10230) );
  NOR2_X1 U10829 ( .A1(n10230), .A2(n10134), .ZN(n10135) );
  AOI211_X1 U10830 ( .C1(n10227), .C2(n10137), .A(n10136), .B(n10135), .ZN(
        n10138) );
  OAI21_X1 U10831 ( .B1(n4856), .B2(n10229), .A(n10138), .ZN(P1_U3272) );
  NAND2_X1 U10832 ( .A1(n10140), .A2(n10139), .ZN(n10141) );
  NAND2_X1 U10833 ( .A1(n10142), .A2(n10141), .ZN(n10156) );
  OR2_X1 U10834 ( .A1(n10156), .A2(n6896), .ZN(n10155) );
  AND2_X1 U10835 ( .A1(n10144), .A2(n10143), .ZN(n10145) );
  OR2_X1 U10836 ( .A1(n4917), .A2(n10145), .ZN(n10153) );
  NAND2_X1 U10837 ( .A1(n10147), .A2(n10146), .ZN(n10148) );
  OAI21_X1 U10838 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(n10151) );
  AOI21_X1 U10839 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(n10154) );
  INV_X1 U10840 ( .A(n10156), .ZN(n10235) );
  NAND2_X1 U10841 ( .A1(n10231), .A2(n10157), .ZN(n10158) );
  NAND2_X1 U10842 ( .A1(n10159), .A2(n10158), .ZN(n10233) );
  INV_X1 U10843 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10162) );
  OAI22_X1 U10844 ( .A1(n10163), .A2(n10162), .B1(n10161), .B2(n10160), .ZN(
        n10164) );
  AOI21_X1 U10845 ( .B1(n10231), .B2(n10165), .A(n10164), .ZN(n10166) );
  OAI21_X1 U10846 ( .B1(n10233), .B2(n10167), .A(n10166), .ZN(n10168) );
  AOI21_X1 U10847 ( .B1(n10235), .B2(n10169), .A(n10168), .ZN(n10170) );
  OAI21_X1 U10848 ( .B1(n10237), .B2(n4856), .A(n10170), .ZN(P1_U3273) );
  NAND2_X1 U10849 ( .A1(n10171), .A2(n10250), .ZN(n10174) );
  AOI21_X1 U10850 ( .B1(n10172), .B2(n10597), .A(n10175), .ZN(n10173) );
  NAND2_X1 U10851 ( .A1(n10174), .A2(n10173), .ZN(n10266) );
  MUX2_X1 U10852 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10266), .S(n10656), .Z(
        P1_U3554) );
  AOI21_X1 U10853 ( .B1(n10176), .B2(n10597), .A(n10175), .ZN(n10177) );
  OAI21_X1 U10854 ( .B1(n10178), .B2(n10633), .A(n10177), .ZN(n10267) );
  MUX2_X1 U10855 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10267), .S(n10656), .Z(
        P1_U3553) );
  AOI22_X1 U10856 ( .A1(n10180), .A2(n10250), .B1(n10597), .B2(n10179), .ZN(
        n10183) );
  NAND3_X1 U10857 ( .A1(n10184), .A2(n10183), .A3(n10182), .ZN(n10268) );
  MUX2_X1 U10858 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10268), .S(n10656), .Z(
        P1_U3551) );
  AOI21_X1 U10859 ( .B1(n10597), .B2(n5955), .A(n10185), .ZN(n10186) );
  OAI211_X1 U10860 ( .C1(n10580), .C2(n10188), .A(n10187), .B(n10186), .ZN(
        n10269) );
  MUX2_X1 U10861 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10269), .S(n10656), .Z(
        P1_U3550) );
  OAI22_X1 U10862 ( .A1(n10190), .A2(n10633), .B1(n10189), .B2(n10651), .ZN(
        n10191) );
  INV_X1 U10863 ( .A(n10191), .ZN(n10192) );
  OAI211_X1 U10864 ( .C1(n10194), .C2(n10600), .A(n10193), .B(n10192), .ZN(
        n10270) );
  MUX2_X1 U10865 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10270), .S(n10656), .Z(
        P1_U3549) );
  AOI21_X1 U10866 ( .B1(n10597), .B2(n10196), .A(n10195), .ZN(n10197) );
  OAI211_X1 U10867 ( .C1(n10580), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        n10271) );
  MUX2_X1 U10868 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10271), .S(n10656), .Z(
        P1_U3548) );
  AOI21_X1 U10869 ( .B1(n10597), .B2(n10201), .A(n10200), .ZN(n10202) );
  OAI211_X1 U10870 ( .C1(n10580), .C2(n10204), .A(n10203), .B(n10202), .ZN(
        n10272) );
  MUX2_X1 U10871 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10272), .S(n10656), .Z(
        P1_U3547) );
  AOI22_X1 U10872 ( .A1(n10206), .A2(n10250), .B1(n10597), .B2(n10205), .ZN(
        n10207) );
  OAI211_X1 U10873 ( .C1(n10580), .C2(n10209), .A(n10208), .B(n10207), .ZN(
        n10273) );
  MUX2_X1 U10874 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10273), .S(n10656), .Z(
        P1_U3546) );
  AOI21_X1 U10875 ( .B1(n10597), .B2(n10211), .A(n10210), .ZN(n10212) );
  OAI211_X1 U10876 ( .C1(n10580), .C2(n10214), .A(n10213), .B(n10212), .ZN(
        n10274) );
  MUX2_X1 U10877 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10274), .S(n10656), .Z(
        P1_U3545) );
  AOI211_X1 U10878 ( .C1(n10597), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        n10218) );
  OAI211_X1 U10879 ( .C1(n10580), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        n10275) );
  MUX2_X1 U10880 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10275), .S(n10656), .Z(
        P1_U3544) );
  AOI21_X1 U10881 ( .B1(n10597), .B2(n10222), .A(n10221), .ZN(n10223) );
  OAI211_X1 U10882 ( .C1(n10580), .C2(n10225), .A(n10224), .B(n10223), .ZN(
        n10276) );
  MUX2_X1 U10883 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10276), .S(n10656), .Z(
        P1_U3543) );
  AOI22_X1 U10884 ( .A1(n10227), .A2(n10250), .B1(n10597), .B2(n10226), .ZN(
        n10228) );
  OAI211_X1 U10885 ( .C1(n10580), .C2(n10230), .A(n10229), .B(n10228), .ZN(
        n10277) );
  MUX2_X1 U10886 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10277), .S(n10656), .Z(
        P1_U3542) );
  INV_X1 U10887 ( .A(n10600), .ZN(n10490) );
  INV_X1 U10888 ( .A(n10231), .ZN(n10232) );
  OAI22_X1 U10889 ( .A1(n10233), .A2(n10633), .B1(n10232), .B2(n10651), .ZN(
        n10234) );
  AOI21_X1 U10890 ( .B1(n10235), .B2(n10490), .A(n10234), .ZN(n10236) );
  NAND2_X1 U10891 ( .A1(n10237), .A2(n10236), .ZN(n10278) );
  MUX2_X1 U10892 ( .A(n10278), .B(P1_REG1_REG_18__SCAN_IN), .S(n10655), .Z(
        P1_U3541) );
  INV_X1 U10893 ( .A(n10238), .ZN(n10243) );
  AOI22_X1 U10894 ( .A1(n10240), .A2(n10250), .B1(n10597), .B2(n10239), .ZN(
        n10241) );
  OAI211_X1 U10895 ( .C1(n10600), .C2(n10243), .A(n10242), .B(n10241), .ZN(
        n10279) );
  MUX2_X1 U10896 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10279), .S(n10656), .Z(
        P1_U3540) );
  AOI211_X1 U10897 ( .C1(n10597), .C2(n10246), .A(n10245), .B(n10244), .ZN(
        n10247) );
  OAI21_X1 U10898 ( .B1(n10580), .B2(n10248), .A(n10247), .ZN(n10280) );
  MUX2_X1 U10899 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10280), .S(n10656), .Z(
        P1_U3539) );
  AOI22_X1 U10900 ( .A1(n10251), .A2(n10250), .B1(n10597), .B2(n10249), .ZN(
        n10252) );
  OAI211_X1 U10901 ( .C1(n10254), .C2(n10580), .A(n10253), .B(n10252), .ZN(
        n10281) );
  MUX2_X1 U10902 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10281), .S(n10656), .Z(
        P1_U3538) );
  AOI211_X1 U10903 ( .C1(n10597), .C2(n10257), .A(n10256), .B(n10255), .ZN(
        n10258) );
  OAI21_X1 U10904 ( .B1(n10259), .B2(n10580), .A(n10258), .ZN(n10282) );
  MUX2_X1 U10905 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10282), .S(n10656), .Z(
        P1_U3537) );
  AOI21_X1 U10906 ( .B1(n10597), .B2(n10261), .A(n10260), .ZN(n10262) );
  OAI211_X1 U10907 ( .C1(n10264), .C2(n10580), .A(n10263), .B(n10262), .ZN(
        n10283) );
  MUX2_X1 U10908 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10283), .S(n10656), .Z(
        P1_U3536) );
  MUX2_X1 U10909 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10265), .S(n10656), .Z(
        P1_U3523) );
  MUX2_X1 U10910 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10266), .S(n4855), .Z(
        P1_U3522) );
  MUX2_X1 U10911 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10267), .S(n4855), .Z(
        P1_U3521) );
  MUX2_X1 U10912 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10268), .S(n4855), .Z(
        P1_U3519) );
  MUX2_X1 U10913 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10269), .S(n4855), .Z(
        P1_U3518) );
  MUX2_X1 U10914 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10270), .S(n4855), .Z(
        P1_U3517) );
  MUX2_X1 U10915 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10271), .S(n4855), .Z(
        P1_U3516) );
  MUX2_X1 U10916 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10272), .S(n4855), .Z(
        P1_U3515) );
  MUX2_X1 U10917 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10273), .S(n4855), .Z(
        P1_U3514) );
  MUX2_X1 U10918 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10274), .S(n4855), .Z(
        P1_U3513) );
  MUX2_X1 U10919 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10275), .S(n4855), .Z(
        P1_U3512) );
  MUX2_X1 U10920 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10276), .S(n4855), .Z(
        P1_U3511) );
  MUX2_X1 U10921 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10277), .S(n4855), .Z(
        P1_U3510) );
  MUX2_X1 U10922 ( .A(n10278), .B(P1_REG0_REG_18__SCAN_IN), .S(n10657), .Z(
        P1_U3508) );
  MUX2_X1 U10923 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10279), .S(n4855), .Z(
        P1_U3505) );
  MUX2_X1 U10924 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10280), .S(n4855), .Z(
        P1_U3502) );
  MUX2_X1 U10925 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10281), .S(n4855), .Z(
        P1_U3499) );
  MUX2_X1 U10926 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10282), .S(n4855), .Z(
        P1_U3496) );
  MUX2_X1 U10927 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10283), .S(n4855), .Z(
        P1_U3493) );
  MUX2_X1 U10928 ( .A(P1_D_REG_0__SCAN_IN), .B(n10284), .S(n10295), .Z(
        P1_U3440) );
  NAND3_X1 U10929 ( .A1(n5329), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n10287) );
  OAI22_X1 U10930 ( .A1(n10285), .A2(n10287), .B1(n6694), .B2(n10286), .ZN(
        n10288) );
  AOI21_X1 U10931 ( .B1(n10290), .B2(n10289), .A(n10288), .ZN(n10291) );
  INV_X1 U10932 ( .A(n10291), .ZN(P1_U3322) );
  MUX2_X1 U10933 ( .A(n10293), .B(n10292), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3353) );
  NAND2_X1 U10934 ( .A1(n10295), .A2(n10294), .ZN(n10296) );
  AND2_X1 U10935 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10296), .ZN(P1_U3321) );
  AND2_X1 U10936 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10296), .ZN(P1_U3320) );
  AND2_X1 U10937 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10296), .ZN(P1_U3319) );
  AND2_X1 U10938 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10296), .ZN(P1_U3318) );
  AND2_X1 U10939 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10296), .ZN(P1_U3317) );
  AND2_X1 U10940 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10296), .ZN(P1_U3316) );
  AND2_X1 U10941 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10296), .ZN(P1_U3315) );
  AND2_X1 U10942 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10296), .ZN(P1_U3314) );
  AND2_X1 U10943 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10296), .ZN(P1_U3313) );
  AND2_X1 U10944 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10296), .ZN(P1_U3312) );
  AND2_X1 U10945 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10296), .ZN(P1_U3311) );
  AND2_X1 U10946 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10296), .ZN(P1_U3310) );
  AND2_X1 U10947 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10296), .ZN(P1_U3309) );
  AND2_X1 U10948 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10296), .ZN(P1_U3308) );
  AND2_X1 U10949 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10296), .ZN(P1_U3307) );
  AND2_X1 U10950 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10296), .ZN(P1_U3306) );
  AND2_X1 U10951 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10296), .ZN(P1_U3305) );
  AND2_X1 U10952 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10296), .ZN(P1_U3304) );
  AND2_X1 U10953 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10296), .ZN(P1_U3303) );
  AND2_X1 U10954 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10296), .ZN(P1_U3302) );
  AND2_X1 U10955 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10296), .ZN(P1_U3301) );
  AND2_X1 U10956 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10296), .ZN(P1_U3300) );
  AND2_X1 U10957 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10296), .ZN(P1_U3299) );
  AND2_X1 U10958 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10296), .ZN(P1_U3298) );
  AND2_X1 U10959 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10296), .ZN(P1_U3297) );
  AND2_X1 U10960 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10296), .ZN(P1_U3296) );
  AND2_X1 U10961 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10296), .ZN(P1_U3295) );
  AND2_X1 U10962 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10296), .ZN(P1_U3294) );
  AND2_X1 U10963 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10296), .ZN(P1_U3293) );
  AND2_X1 U10964 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10296), .ZN(P1_U3292) );
  INV_X1 U10965 ( .A(n10297), .ZN(n10298) );
  NAND2_X1 U10966 ( .A1(n10299), .A2(n10298), .ZN(n10421) );
  AOI22_X1 U10967 ( .A1(n10301), .A2(n10423), .B1(n10300), .B2(n10421), .ZN(
        P2_U3438) );
  AND2_X1 U10968 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10421), .ZN(P2_U3326) );
  AND2_X1 U10969 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10421), .ZN(P2_U3325) );
  AND2_X1 U10970 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10421), .ZN(P2_U3324) );
  AND2_X1 U10971 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10421), .ZN(P2_U3323) );
  AND2_X1 U10972 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10421), .ZN(P2_U3322) );
  AND2_X1 U10973 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10421), .ZN(P2_U3321) );
  AND2_X1 U10974 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10421), .ZN(P2_U3320) );
  AND2_X1 U10975 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10421), .ZN(P2_U3319) );
  AND2_X1 U10976 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10421), .ZN(P2_U3318) );
  AND2_X1 U10977 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10421), .ZN(P2_U3317) );
  AND2_X1 U10978 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10421), .ZN(P2_U3316) );
  AND2_X1 U10979 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10421), .ZN(P2_U3315) );
  AND2_X1 U10980 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10421), .ZN(P2_U3314) );
  AND2_X1 U10981 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10421), .ZN(P2_U3313) );
  AND2_X1 U10982 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10421), .ZN(P2_U3312) );
  AND2_X1 U10983 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10421), .ZN(P2_U3311) );
  AND2_X1 U10984 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10421), .ZN(P2_U3310) );
  AND2_X1 U10985 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10421), .ZN(P2_U3309) );
  AND2_X1 U10986 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10421), .ZN(P2_U3308) );
  AND2_X1 U10987 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10421), .ZN(P2_U3307) );
  AND2_X1 U10988 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10421), .ZN(P2_U3306) );
  AND2_X1 U10989 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10421), .ZN(P2_U3305) );
  AND2_X1 U10990 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10421), .ZN(P2_U3304) );
  AND2_X1 U10991 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10421), .ZN(P2_U3303) );
  AND2_X1 U10992 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10421), .ZN(P2_U3302) );
  AND2_X1 U10993 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10421), .ZN(P2_U3301) );
  AND2_X1 U10994 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10421), .ZN(P2_U3300) );
  AND2_X1 U10995 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10421), .ZN(P2_U3299) );
  AND2_X1 U10996 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10421), .ZN(P2_U3298) );
  AND2_X1 U10997 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10421), .ZN(P2_U3297) );
  XOR2_X1 U10998 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  NAND3_X1 U10999 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10304) );
  AOI21_X1 U11000 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10306) );
  INV_X1 U11001 ( .A(n10306), .ZN(n10302) );
  NAND2_X1 U11002 ( .A1(n10304), .A2(n10302), .ZN(n10303) );
  XNOR2_X1 U11003 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10303), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11004 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10308) );
  INV_X1 U11005 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10305) );
  OAI21_X1 U11006 ( .B1(n10306), .B2(n10305), .A(n10304), .ZN(n10307) );
  XOR2_X1 U11007 ( .A(n10308), .B(n10307), .Z(ADD_1071_U54) );
  XOR2_X1 U11008 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10312) );
  NAND2_X1 U11009 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10310) );
  NAND2_X1 U11010 ( .A1(n10308), .A2(n10307), .ZN(n10309) );
  NAND2_X1 U11011 ( .A1(n10310), .A2(n10309), .ZN(n10311) );
  XOR2_X1 U11012 ( .A(n10312), .B(n10311), .Z(ADD_1071_U53) );
  XNOR2_X1 U11013 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10316) );
  NAND2_X1 U11014 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10314) );
  NAND2_X1 U11015 ( .A1(n10312), .A2(n10311), .ZN(n10313) );
  NAND2_X1 U11016 ( .A1(n10314), .A2(n10313), .ZN(n10315) );
  XNOR2_X1 U11017 ( .A(n10316), .B(n10315), .ZN(ADD_1071_U52) );
  NOR2_X1 U11018 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10318) );
  NOR2_X1 U11019 ( .A1(n10316), .A2(n10315), .ZN(n10317) );
  NOR2_X1 U11020 ( .A1(n10318), .A2(n10317), .ZN(n10319) );
  NOR2_X1 U11021 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10319), .ZN(n10323) );
  AND2_X1 U11022 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10319), .ZN(n10321) );
  NOR2_X1 U11023 ( .A1(n10323), .A2(n10321), .ZN(n10320) );
  XOR2_X1 U11024 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10320), .Z(ADD_1071_U51) );
  NOR2_X1 U11025 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10321), .ZN(n10322) );
  NOR2_X1 U11026 ( .A1(n10323), .A2(n10322), .ZN(n10324) );
  XOR2_X1 U11027 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10324), .Z(n10325) );
  XOR2_X1 U11028 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10325), .Z(ADD_1071_U50) );
  NAND2_X1 U11029 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10324), .ZN(n10327) );
  NAND2_X1 U11030 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10325), .ZN(n10326) );
  NAND2_X1 U11031 ( .A1(n10327), .A2(n10326), .ZN(n10328) );
  XOR2_X1 U11032 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10328), .Z(n10329) );
  XOR2_X1 U11033 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10329), .Z(ADD_1071_U49) );
  NAND2_X1 U11034 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10328), .ZN(n10331) );
  NAND2_X1 U11035 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10329), .ZN(n10330) );
  NAND2_X1 U11036 ( .A1(n10331), .A2(n10330), .ZN(n10332) );
  XOR2_X1 U11037 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10332), .Z(n10333) );
  XOR2_X1 U11038 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10333), .Z(ADD_1071_U48) );
  NAND2_X1 U11039 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10332), .ZN(n10335) );
  NAND2_X1 U11040 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10333), .ZN(n10334) );
  NAND2_X1 U11041 ( .A1(n10335), .A2(n10334), .ZN(n10336) );
  XOR2_X1 U11042 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n10336), .Z(n10337) );
  XOR2_X1 U11043 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10337), .Z(ADD_1071_U47) );
  XOR2_X1 U11044 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10341) );
  NAND2_X1 U11045 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n10336), .ZN(n10339) );
  NAND2_X1 U11046 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10337), .ZN(n10338) );
  NAND2_X1 U11047 ( .A1(n10339), .A2(n10338), .ZN(n10340) );
  XOR2_X1 U11048 ( .A(n10341), .B(n10340), .Z(ADD_1071_U63) );
  XOR2_X1 U11049 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10345) );
  NAND2_X1 U11050 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10343) );
  NAND2_X1 U11051 ( .A1(n10341), .A2(n10340), .ZN(n10342) );
  NAND2_X1 U11052 ( .A1(n10343), .A2(n10342), .ZN(n10344) );
  XOR2_X1 U11053 ( .A(n10345), .B(n10344), .Z(ADD_1071_U62) );
  NAND2_X1 U11054 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10347) );
  NAND2_X1 U11055 ( .A1(n10345), .A2(n10344), .ZN(n10346) );
  NAND2_X1 U11056 ( .A1(n10347), .A2(n10346), .ZN(n10349) );
  XNOR2_X1 U11057 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10348) );
  XNOR2_X1 U11058 ( .A(n10349), .B(n10348), .ZN(ADD_1071_U61) );
  NOR2_X1 U11059 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10351) );
  NOR2_X1 U11060 ( .A1(n10349), .A2(n10348), .ZN(n10350) );
  NOR2_X1 U11061 ( .A1(n10351), .A2(n10350), .ZN(n10353) );
  XNOR2_X1 U11062 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10352) );
  XNOR2_X1 U11063 ( .A(n10353), .B(n10352), .ZN(ADD_1071_U60) );
  NOR2_X1 U11064 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10355) );
  NOR2_X1 U11065 ( .A1(n10353), .A2(n10352), .ZN(n10354) );
  NOR2_X1 U11066 ( .A1(n10355), .A2(n10354), .ZN(n10357) );
  XNOR2_X1 U11067 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10356) );
  XNOR2_X1 U11068 ( .A(n10357), .B(n10356), .ZN(ADD_1071_U59) );
  NOR2_X1 U11069 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10359) );
  NOR2_X1 U11070 ( .A1(n10357), .A2(n10356), .ZN(n10358) );
  NOR2_X1 U11071 ( .A1(n10359), .A2(n10358), .ZN(n10361) );
  XNOR2_X1 U11072 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10360) );
  XNOR2_X1 U11073 ( .A(n10361), .B(n10360), .ZN(ADD_1071_U58) );
  NOR2_X1 U11074 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10363) );
  NOR2_X1 U11075 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  NOR2_X1 U11076 ( .A1(n10363), .A2(n10362), .ZN(n10365) );
  XNOR2_X1 U11077 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10364) );
  XNOR2_X1 U11078 ( .A(n10365), .B(n10364), .ZN(ADD_1071_U57) );
  NOR2_X1 U11079 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10367) );
  NOR2_X1 U11080 ( .A1(n10365), .A2(n10364), .ZN(n10366) );
  NOR2_X1 U11081 ( .A1(n10367), .A2(n10366), .ZN(n10369) );
  XNOR2_X1 U11082 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10368) );
  XNOR2_X1 U11083 ( .A(n10369), .B(n10368), .ZN(ADD_1071_U56) );
  NOR2_X1 U11084 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10371) );
  NOR2_X1 U11085 ( .A1(n10369), .A2(n10368), .ZN(n10370) );
  NOR2_X1 U11086 ( .A1(n10371), .A2(n10370), .ZN(n10372) );
  NOR2_X1 U11087 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10372), .ZN(n10375) );
  AND2_X1 U11088 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10372), .ZN(n10374) );
  NOR2_X1 U11089 ( .A1(n10375), .A2(n10374), .ZN(n10373) );
  XOR2_X1 U11090 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10373), .Z(ADD_1071_U55)
         );
  NOR2_X1 U11091 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10374), .ZN(n10376) );
  NOR2_X1 U11092 ( .A1(n10376), .A2(n10375), .ZN(n10378) );
  XNOR2_X1 U11093 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10377) );
  XNOR2_X1 U11094 ( .A(n10378), .B(n10377), .ZN(ADD_1071_U4) );
  AOI22_X1 U11095 ( .A1(n10407), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n10406), 
        .B2(n10379), .ZN(n10390) );
  INV_X1 U11096 ( .A(n10380), .ZN(n10389) );
  OAI211_X1 U11097 ( .C1(n10383), .C2(n10382), .A(n10398), .B(n10381), .ZN(
        n10388) );
  OAI211_X1 U11098 ( .C1(n10386), .C2(n10385), .A(n10414), .B(n10384), .ZN(
        n10387) );
  NAND4_X1 U11099 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        P1_U3247) );
  AOI22_X1 U11100 ( .A1(n10407), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n10406), 
        .B2(n10391), .ZN(n10404) );
  AOI21_X1 U11101 ( .B1(n10394), .B2(n10393), .A(n10392), .ZN(n10396) );
  OR2_X1 U11102 ( .A1(n10396), .A2(n10395), .ZN(n10402) );
  OAI211_X1 U11103 ( .C1(n10400), .C2(n10399), .A(n10398), .B(n10397), .ZN(
        n10401) );
  NAND4_X1 U11104 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        P1_U3251) );
  AOI22_X1 U11105 ( .A1(n10407), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n10406), 
        .B2(n10405), .ZN(n10420) );
  AOI21_X1 U11106 ( .B1(n10410), .B2(n10409), .A(n10408), .ZN(n10411) );
  OR2_X1 U11107 ( .A1(n10412), .A2(n10411), .ZN(n10418) );
  OAI211_X1 U11108 ( .C1(n10416), .C2(n10415), .A(n10414), .B(n10413), .ZN(
        n10417) );
  NAND4_X1 U11109 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        P1_U3246) );
  AOI22_X1 U11110 ( .A1(n10424), .A2(n10423), .B1(n10422), .B2(n10421), .ZN(
        P2_U3437) );
  AOI22_X1 U11111 ( .A1(n10425), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10457), .ZN(n10432) );
  AOI22_X1 U11112 ( .A1(n10448), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10431) );
  OAI21_X1 U11113 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10427), .A(n10426), .ZN(
        n10429) );
  NOR2_X1 U11114 ( .A1(n10449), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10428) );
  OAI21_X1 U11115 ( .B1(n10429), .B2(n10428), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10430) );
  OAI211_X1 U11116 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10432), .A(n10431), .B(
        n10430), .ZN(P2_U3245) );
  NAND2_X1 U11117 ( .A1(n10434), .A2(n10433), .ZN(n10437) );
  INV_X1 U11118 ( .A(n10435), .ZN(n10436) );
  NAND2_X1 U11119 ( .A1(n10437), .A2(n10436), .ZN(n10441) );
  NAND2_X1 U11120 ( .A1(n10455), .A2(n10438), .ZN(n10440) );
  AOI22_X1 U11121 ( .A1(n10448), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10439) );
  OAI211_X1 U11122 ( .C1(n10441), .C2(n10449), .A(n10440), .B(n10439), .ZN(
        n10442) );
  INV_X1 U11123 ( .A(n10442), .ZN(n10447) );
  AND2_X1 U11124 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10445) );
  OAI211_X1 U11125 ( .C1(n10445), .C2(n10444), .A(n10457), .B(n10443), .ZN(
        n10446) );
  NAND2_X1 U11126 ( .A1(n10447), .A2(n10446), .ZN(P2_U3246) );
  AOI22_X1 U11127 ( .A1(n10448), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10462) );
  AOI211_X1 U11128 ( .C1(n10452), .C2(n10451), .A(n10450), .B(n10449), .ZN(
        n10453) );
  AOI21_X1 U11129 ( .B1(n10455), .B2(n10454), .A(n10453), .ZN(n10461) );
  OAI211_X1 U11130 ( .C1(n10459), .C2(n10458), .A(n10457), .B(n10456), .ZN(
        n10460) );
  NAND3_X1 U11131 ( .A1(n10462), .A2(n10461), .A3(n10460), .ZN(P2_U3247) );
  XNOR2_X1 U11132 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U11133 ( .A1(n10463), .A2(n10666), .ZN(n10466) );
  INV_X1 U11134 ( .A(n10464), .ZN(n10465) );
  AOI211_X1 U11135 ( .C1(n10468), .C2(n10467), .A(n10466), .B(n10465), .ZN(
        n10469) );
  AOI22_X1 U11136 ( .A1(n10685), .A2(n10469), .B1(n6044), .B2(n10684), .ZN(
        P2_U3520) );
  AOI22_X1 U11137 ( .A1(n10689), .A2(n10469), .B1(n6043), .B2(n10686), .ZN(
        P2_U3451) );
  INV_X1 U11138 ( .A(n10470), .ZN(n10475) );
  OAI21_X1 U11139 ( .B1(n10472), .B2(n10651), .A(n10471), .ZN(n10474) );
  AOI211_X1 U11140 ( .C1(n10490), .C2(n10475), .A(n10474), .B(n10473), .ZN(
        n10476) );
  AOI22_X1 U11141 ( .A1(n10656), .A2(n10476), .B1(n6671), .B2(n10655), .ZN(
        P1_U3524) );
  AOI22_X1 U11142 ( .A1(n4855), .A2(n10476), .B1(n5340), .B2(n10657), .ZN(
        P1_U3457) );
  INV_X1 U11143 ( .A(n10477), .ZN(n10593) );
  OAI22_X1 U11144 ( .A1(n10479), .A2(n10678), .B1(n10478), .B2(n10676), .ZN(
        n10482) );
  INV_X1 U11145 ( .A(n10480), .ZN(n10481) );
  AOI211_X1 U11146 ( .C1(n10593), .C2(n10483), .A(n10482), .B(n10481), .ZN(
        n10484) );
  AOI22_X1 U11147 ( .A1(n10685), .A2(n10484), .B1(n7069), .B2(n10684), .ZN(
        P2_U3522) );
  AOI22_X1 U11148 ( .A1(n10689), .A2(n10484), .B1(n6058), .B2(n10686), .ZN(
        P2_U3457) );
  OAI22_X1 U11149 ( .A1(n10486), .A2(n10633), .B1(n10485), .B2(n10651), .ZN(
        n10488) );
  AOI211_X1 U11150 ( .C1(n10490), .C2(n10489), .A(n10488), .B(n10487), .ZN(
        n10492) );
  AOI22_X1 U11151 ( .A1(n10656), .A2(n10492), .B1(n6676), .B2(n10655), .ZN(
        P1_U3526) );
  INV_X1 U11152 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U11153 ( .A1(n4855), .A2(n10492), .B1(n10491), .B2(n10657), .ZN(
        P1_U3463) );
  NAND3_X1 U11154 ( .A1(n10560), .A2(n10493), .A3(n6947), .ZN(n10498) );
  OAI21_X1 U11155 ( .B1(n10495), .B2(n10494), .A(n10561), .ZN(n10497) );
  AOI21_X1 U11156 ( .B1(n10498), .B2(n10497), .A(n10496), .ZN(n10505) );
  OAI22_X1 U11157 ( .A1(n10500), .A2(n6948), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10499), .ZN(n10504) );
  OAI22_X1 U11158 ( .A1(n6546), .A2(n10502), .B1(n10501), .B2(n10611), .ZN(
        n10503) );
  NOR3_X1 U11159 ( .A1(n10505), .A2(n10504), .A3(n10503), .ZN(n10506) );
  OAI21_X1 U11160 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n10623), .A(n10506), .ZN(
        P2_U3220) );
  OAI22_X1 U11161 ( .A1(n10508), .A2(n10678), .B1(n10507), .B2(n10676), .ZN(
        n10510) );
  AOI211_X1 U11162 ( .C1(n10682), .C2(n10511), .A(n10510), .B(n10509), .ZN(
        n10512) );
  AOI22_X1 U11163 ( .A1(n10685), .A2(n10512), .B1(n6092), .B2(n10684), .ZN(
        P2_U3524) );
  AOI22_X1 U11164 ( .A1(n10689), .A2(n10512), .B1(n6094), .B2(n10686), .ZN(
        P2_U3463) );
  AOI21_X1 U11165 ( .B1(n10597), .B2(n10514), .A(n10513), .ZN(n10515) );
  OAI211_X1 U11166 ( .C1(n10580), .C2(n10517), .A(n10516), .B(n10515), .ZN(
        n10518) );
  INV_X1 U11167 ( .A(n10518), .ZN(n10519) );
  AOI22_X1 U11168 ( .A1(n10656), .A2(n10519), .B1(n6670), .B2(n10655), .ZN(
        P1_U3528) );
  AOI22_X1 U11169 ( .A1(n4855), .A2(n10519), .B1(n5446), .B2(n10657), .ZN(
        P1_U3469) );
  AND2_X1 U11170 ( .A1(n10520), .A2(n10682), .ZN(n10524) );
  OAI21_X1 U11171 ( .B1(n10522), .B2(n10676), .A(n10521), .ZN(n10523) );
  NOR3_X1 U11172 ( .A1(n10525), .A2(n10524), .A3(n10523), .ZN(n10526) );
  AOI22_X1 U11173 ( .A1(n10685), .A2(n10526), .B1(n6108), .B2(n10684), .ZN(
        P2_U3525) );
  AOI22_X1 U11174 ( .A1(n10689), .A2(n10526), .B1(n6114), .B2(n10686), .ZN(
        P2_U3466) );
  AOI22_X1 U11175 ( .A1(n10529), .A2(n10528), .B1(n10554), .B2(n10527), .ZN(
        n10533) );
  NAND3_X1 U11176 ( .A1(n10531), .A2(n10530), .A3(n10682), .ZN(n10532) );
  AND3_X1 U11177 ( .A1(n10534), .A2(n10533), .A3(n10532), .ZN(n10535) );
  AOI22_X1 U11178 ( .A1(n10685), .A2(n10535), .B1(n6127), .B2(n10684), .ZN(
        P2_U3526) );
  AOI22_X1 U11179 ( .A1(n10689), .A2(n10535), .B1(n6129), .B2(n10686), .ZN(
        P2_U3469) );
  AOI22_X1 U11180 ( .A1(n10609), .A2(n10536), .B1(P2_U3152), .B2(
        P2_REG3_REG_7__SCAN_IN), .ZN(n10537) );
  OAI21_X1 U11181 ( .B1(n10538), .B2(n10611), .A(n10537), .ZN(n10543) );
  INV_X1 U11182 ( .A(n10539), .ZN(n10563) );
  AOI211_X1 U11183 ( .C1(n10541), .C2(n10540), .A(n10615), .B(n10563), .ZN(
        n10542) );
  AOI211_X1 U11184 ( .C1(n10621), .C2(n10544), .A(n10543), .B(n10542), .ZN(
        n10545) );
  OAI21_X1 U11185 ( .B1(n10546), .B2(n10623), .A(n10545), .ZN(P2_U3215) );
  OAI22_X1 U11186 ( .A1(n10548), .A2(n10678), .B1(n10547), .B2(n10676), .ZN(
        n10549) );
  AOI21_X1 U11187 ( .B1(n10550), .B2(n10682), .A(n10549), .ZN(n10551) );
  AND2_X1 U11188 ( .A1(n10552), .A2(n10551), .ZN(n10553) );
  AOI22_X1 U11189 ( .A1(n10685), .A2(n10553), .B1(n7151), .B2(n10684), .ZN(
        P2_U3527) );
  AOI22_X1 U11190 ( .A1(n10689), .A2(n10553), .B1(n6143), .B2(n10686), .ZN(
        P2_U3472) );
  NAND2_X1 U11191 ( .A1(n10555), .A2(n10554), .ZN(n10576) );
  INV_X1 U11192 ( .A(n10576), .ZN(n10569) );
  AOI22_X1 U11193 ( .A1(n10609), .A2(n10558), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10556) );
  OAI21_X1 U11194 ( .B1(n10557), .B2(n10611), .A(n10556), .ZN(n10568) );
  NAND3_X1 U11195 ( .A1(n10560), .A2(n10559), .A3(n10558), .ZN(n10566) );
  OAI21_X1 U11196 ( .B1(n10563), .B2(n10562), .A(n10561), .ZN(n10565) );
  AOI21_X1 U11197 ( .B1(n10566), .B2(n10565), .A(n10564), .ZN(n10567) );
  AOI211_X1 U11198 ( .C1(n10570), .C2(n10569), .A(n10568), .B(n10567), .ZN(
        n10571) );
  OAI21_X1 U11199 ( .B1(n10572), .B2(n10623), .A(n10571), .ZN(P2_U3223) );
  NAND3_X1 U11200 ( .A1(n7586), .A2(n10573), .A3(n10682), .ZN(n10574) );
  AND4_X1 U11201 ( .A1(n10577), .A2(n10576), .A3(n10575), .A4(n10574), .ZN(
        n10579) );
  AOI22_X1 U11202 ( .A1(n10685), .A2(n10579), .B1(n10578), .B2(n10684), .ZN(
        P2_U3528) );
  AOI22_X1 U11203 ( .A1(n10689), .A2(n10579), .B1(n6163), .B2(n10686), .ZN(
        P2_U3475) );
  OAI21_X1 U11204 ( .B1(n5181), .B2(n10651), .A(n10582), .ZN(n10584) );
  AOI211_X1 U11205 ( .C1(n10585), .C2(n5960), .A(n10584), .B(n10583), .ZN(
        n10587) );
  AOI22_X1 U11206 ( .A1(n10656), .A2(n10587), .B1(n5517), .B2(n10655), .ZN(
        P1_U3532) );
  INV_X1 U11207 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U11208 ( .A1(n4855), .A2(n10587), .B1(n10586), .B2(n10657), .ZN(
        P1_U3481) );
  OAI22_X1 U11209 ( .A1(n10589), .A2(n10678), .B1(n5018), .B2(n10676), .ZN(
        n10591) );
  AOI211_X1 U11210 ( .C1(n10593), .C2(n10592), .A(n10591), .B(n10590), .ZN(
        n10594) );
  AOI22_X1 U11211 ( .A1(n10685), .A2(n10594), .B1(n7155), .B2(n10684), .ZN(
        P2_U3529) );
  AOI22_X1 U11212 ( .A1(n10689), .A2(n10594), .B1(n6177), .B2(n10686), .ZN(
        P2_U3478) );
  AOI21_X1 U11213 ( .B1(n10597), .B2(n10596), .A(n10595), .ZN(n10598) );
  OAI211_X1 U11214 ( .C1(n10601), .C2(n10600), .A(n10599), .B(n10598), .ZN(
        n10602) );
  AOI21_X1 U11215 ( .B1(n10604), .B2(n10603), .A(n10602), .ZN(n10606) );
  AOI22_X1 U11216 ( .A1(n10656), .A2(n10606), .B1(n6811), .B2(n10655), .ZN(
        P1_U3533) );
  INV_X1 U11217 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U11218 ( .A1(n4855), .A2(n10606), .B1(n10605), .B2(n10657), .ZN(
        P1_U3484) );
  AOI22_X1 U11219 ( .A1(n10609), .A2(n10608), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10610) );
  OAI21_X1 U11220 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(n10619) );
  INV_X1 U11221 ( .A(n10613), .ZN(n10614) );
  AOI211_X1 U11222 ( .C1(n10617), .C2(n10616), .A(n10615), .B(n10614), .ZN(
        n10618) );
  AOI211_X1 U11223 ( .C1(n10621), .C2(n10620), .A(n10619), .B(n10618), .ZN(
        n10622) );
  OAI21_X1 U11224 ( .B1(n10624), .B2(n10623), .A(n10622), .ZN(P2_U3219) );
  NOR2_X1 U11225 ( .A1(n10625), .A2(n10666), .ZN(n10630) );
  OAI22_X1 U11226 ( .A1(n10627), .A2(n10678), .B1(n10626), .B2(n10676), .ZN(
        n10629) );
  AOI211_X1 U11227 ( .C1(n10630), .C2(n7716), .A(n10629), .B(n10628), .ZN(
        n10631) );
  AOI22_X1 U11228 ( .A1(n10685), .A2(n10631), .B1(n7142), .B2(n10684), .ZN(
        P2_U3530) );
  AOI22_X1 U11229 ( .A1(n10689), .A2(n10631), .B1(n6199), .B2(n10686), .ZN(
        P2_U3481) );
  OAI22_X1 U11230 ( .A1(n10634), .A2(n10633), .B1(n10632), .B2(n10651), .ZN(
        n10636) );
  AOI211_X1 U11231 ( .C1(n5960), .C2(n10637), .A(n10636), .B(n10635), .ZN(
        n10639) );
  AOI22_X1 U11232 ( .A1(n10656), .A2(n10639), .B1(n5557), .B2(n10655), .ZN(
        P1_U3534) );
  INV_X1 U11233 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U11234 ( .A1(n4855), .A2(n10639), .B1(n10638), .B2(n10657), .ZN(
        P1_U3487) );
  OAI211_X1 U11235 ( .C1(n10642), .C2(n10676), .A(n10641), .B(n10640), .ZN(
        n10643) );
  AOI21_X1 U11236 ( .B1(n10644), .B2(n10682), .A(n10643), .ZN(n10646) );
  AOI22_X1 U11237 ( .A1(n10685), .A2(n10646), .B1(n7141), .B2(n10684), .ZN(
        P2_U3531) );
  INV_X1 U11238 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U11239 ( .A1(n10689), .A2(n10646), .B1(n10645), .B2(n10686), .ZN(
        P2_U3484) );
  NAND3_X1 U11240 ( .A1(n10648), .A2(n10647), .A3(n5960), .ZN(n10650) );
  OAI211_X1 U11241 ( .C1(n10652), .C2(n10651), .A(n10650), .B(n10649), .ZN(
        n10653) );
  NOR2_X1 U11242 ( .A1(n10654), .A2(n10653), .ZN(n10659) );
  AOI22_X1 U11243 ( .A1(n10656), .A2(n10659), .B1(n6989), .B2(n10655), .ZN(
        P1_U3535) );
  INV_X1 U11244 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U11245 ( .A1(n4855), .A2(n10659), .B1(n10658), .B2(n10657), .ZN(
        P1_U3490) );
  OAI22_X1 U11246 ( .A1(n10661), .A2(n10678), .B1(n10660), .B2(n10676), .ZN(
        n10663) );
  AOI211_X1 U11247 ( .C1(n10682), .C2(n10664), .A(n10663), .B(n10662), .ZN(
        n10665) );
  AOI22_X1 U11248 ( .A1(n10685), .A2(n10665), .B1(n7158), .B2(n10684), .ZN(
        P2_U3532) );
  AOI22_X1 U11249 ( .A1(n10689), .A2(n10665), .B1(n6248), .B2(n10686), .ZN(
        P2_U3487) );
  NOR2_X1 U11250 ( .A1(n10667), .A2(n10666), .ZN(n10672) );
  OAI22_X1 U11251 ( .A1(n10669), .A2(n10678), .B1(n10668), .B2(n10676), .ZN(
        n10671) );
  AOI211_X1 U11252 ( .C1(n10672), .C2(n7973), .A(n10671), .B(n10670), .ZN(
        n10674) );
  AOI22_X1 U11253 ( .A1(n10685), .A2(n10674), .B1(n6233), .B2(n10684), .ZN(
        P2_U3533) );
  INV_X1 U11254 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U11255 ( .A1(n10689), .A2(n10674), .B1(n10673), .B2(n10686), .ZN(
        P2_U3490) );
  INV_X1 U11256 ( .A(n10675), .ZN(n10683) );
  OAI22_X1 U11257 ( .A1(n10679), .A2(n10678), .B1(n10677), .B2(n10676), .ZN(
        n10680) );
  AOI211_X1 U11258 ( .C1(n10683), .C2(n10682), .A(n10681), .B(n10680), .ZN(
        n10688) );
  AOI22_X1 U11259 ( .A1(n10685), .A2(n10688), .B1(n6278), .B2(n10684), .ZN(
        P2_U3534) );
  INV_X1 U11260 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U11261 ( .A1(n10689), .A2(n10688), .B1(n10687), .B2(n10686), .ZN(
        P2_U3493) );
  XNOR2_X1 U11262 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  NAND2_X2 U5007 ( .A1(n6038), .A2(n6037), .ZN(n6448) );
  XNOR2_X1 U4949 ( .A(n6031), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6038) );
  CLKBUF_X1 U4931 ( .A(n6093), .Z(n6692) );
  NAND2_X2 U4964 ( .A1(n6547), .A2(n7063), .ZN(n7074) );
endmodule

