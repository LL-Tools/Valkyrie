

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157;

  NOR2_X1 U5182 ( .A1(n9358), .A2(n8600), .ZN(n9357) );
  CLKBUF_X2 U5183 ( .A(n7117), .Z(n7072) );
  OAI21_X1 U5184 ( .B1(n7421), .B2(n7546), .A(n7532), .ZN(n7422) );
  CLKBUF_X2 U5185 ( .A(n6900), .Z(n7117) );
  INV_X1 U5186 ( .A(n6789), .ZN(n9311) );
  CLKBUF_X3 U5188 ( .A(n6601), .Z(n5121) );
  INV_X1 U5189 ( .A(n8818), .ZN(n6310) );
  NAND2_X1 U5190 ( .A1(n5745), .A2(n5354), .ZN(n5353) );
  INV_X1 U5191 ( .A(n8635), .ZN(n6373) );
  CLKBUF_X2 U5192 ( .A(n6887), .Z(n7123) );
  AND2_X1 U5193 ( .A1(n5912), .A2(n5897), .ZN(n5713) );
  INV_X1 U5194 ( .A(n8996), .ZN(n6377) );
  OAI21_X1 U5195 ( .B1(n7536), .B2(n5459), .A(n5458), .ZN(n7517) );
  INV_X1 U5196 ( .A(n7059), .ZN(n7118) );
  INV_X1 U5197 ( .A(n6784), .ZN(n6733) );
  OR2_X1 U5198 ( .A1(n8497), .A2(n8496), .ZN(n8575) );
  OR2_X1 U5199 ( .A1(n9236), .A2(n9235), .ZN(n9925) );
  INV_X1 U5200 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6521) );
  INV_X1 U5201 ( .A(n6274), .ZN(n8852) );
  NOR2_X1 U5203 ( .A1(n6314), .A2(n10932), .ZN(n7448) );
  NAND2_X2 U5204 ( .A1(n6789), .A2(n6788), .ZN(n7153) );
  XNOR2_X1 U5205 ( .A(n6383), .B(n6382), .ZN(n6788) );
  XNOR2_X1 U5206 ( .A(n8575), .B(n8498), .ZN(n8499) );
  MUX2_X1 U5207 ( .A(n8628), .B(n8627), .S(n9417), .Z(n8631) );
  NAND2_X1 U5208 ( .A1(n6120), .A2(n6119), .ZN(n10572) );
  NAND2_X1 U5209 ( .A1(n6136), .A2(n6135), .ZN(n10568) );
  NAND2_X1 U5210 ( .A1(n6158), .A2(n6157), .ZN(n10405) );
  XNOR2_X1 U5211 ( .A(n5744), .B(n5743), .ZN(n6311) );
  CLKBUF_X3 U5212 ( .A(n7155), .Z(n5120) );
  AOI211_X1 U5213 ( .C1(n8632), .C2(n9429), .A(n8631), .B(n8630), .ZN(n8633)
         );
  AND2_X2 U5214 ( .A1(n5572), .A2(n5571), .ZN(n10173) );
  BUF_X4 U5216 ( .A(n7121), .Z(n5119) );
  NAND2_X2 U5217 ( .A1(n6854), .A2(n6853), .ZN(n7121) );
  NOR3_X2 U5218 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n6366) );
  NAND2_X2 U5219 ( .A1(n10052), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6368) );
  INV_X1 U5220 ( .A(n5785), .ZN(n7155) );
  NOR2_X2 U5221 ( .A1(n6689), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6699) );
  NAND2_X2 U5222 ( .A1(n6847), .A2(n6846), .ZN(n7060) );
  OAI222_X1 U5223 ( .A1(n10659), .A2(n8240), .B1(n7742), .B2(n8239), .C1(
        P1_U3086), .C2(n6274), .ZN(P1_U3333) );
  NAND2_X2 U5224 ( .A1(n7321), .A2(n6397), .ZN(n7416) );
  INV_X4 U5225 ( .A(n9311), .ZN(n9412) );
  NAND2_X2 U5226 ( .A1(n6918), .A2(n7504), .ZN(n10161) );
  NOR2_X2 U5227 ( .A1(n8185), .A2(n8184), .ZN(n8187) );
  XNOR2_X2 U5228 ( .A(n8586), .B(n8605), .ZN(n8504) );
  AND2_X2 U5229 ( .A1(n8503), .A2(n8502), .ZN(n8586) );
  AOI21_X1 U5230 ( .B1(n9912), .B2(n6708), .A(n6707), .ZN(n9900) );
  NAND2_X1 U5231 ( .A1(n10012), .A2(n6773), .ZN(n9115) );
  NAND2_X1 U5232 ( .A1(n7713), .A2(n7712), .ZN(n7711) );
  INV_X1 U5233 ( .A(n7550), .ZN(n8959) );
  INV_X1 U5234 ( .A(n7773), .ZN(n7489) );
  INV_X1 U5235 ( .A(n10211), .ZN(n7462) );
  INV_X2 U5236 ( .A(n8815), .ZN(n8782) );
  INV_X2 U5237 ( .A(n6408), .ZN(n6399) );
  NAND4_X1 U5238 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n10213)
         );
  INV_X8 U5239 ( .A(n6017), .ZN(n8647) );
  NAND2_X1 U5240 ( .A1(n8635), .A2(n6377), .ZN(n6477) );
  CLKBUF_X2 U5241 ( .A(n6311), .Z(n5123) );
  NAND2_X1 U5242 ( .A1(n5120), .A2(P1_U3086), .ZN(n10659) );
  NOR2_X1 U5243 ( .A1(n10173), .A2(n5570), .ZN(n7128) );
  NAND2_X1 U5244 ( .A1(n5288), .A2(n9307), .ZN(n5287) );
  OR2_X1 U5245 ( .A1(n8934), .A2(n6261), .ZN(n10333) );
  AOI21_X1 U5246 ( .B1(n9444), .B2(n10935), .A(n9443), .ZN(n9994) );
  AOI21_X1 U5247 ( .B1(n5202), .B2(n10935), .A(n5200), .ZN(n10002) );
  AND2_X1 U5248 ( .A1(n5466), .A2(n5136), .ZN(n9407) );
  NAND2_X1 U5249 ( .A1(n7000), .A2(n6999), .ZN(n10185) );
  NAND2_X1 U5250 ( .A1(n8615), .A2(n8614), .ZN(n9393) );
  OR2_X1 U5251 ( .A1(n9391), .A2(n5468), .ZN(n5466) );
  AND2_X1 U5252 ( .A1(n9976), .A2(n6654), .ZN(n9960) );
  NOR2_X1 U5253 ( .A1(n5297), .A2(n5295), .ZN(n5294) );
  NAND2_X1 U5254 ( .A1(n9362), .A2(n8610), .ZN(n9383) );
  XNOR2_X1 U5255 ( .A(n8582), .B(n8618), .ZN(n9391) );
  NOR2_X1 U5256 ( .A1(n9261), .A2(n9262), .ZN(n5295) );
  NAND2_X1 U5257 ( .A1(n10908), .A2(n5187), .ZN(n8441) );
  NAND2_X1 U5258 ( .A1(n6174), .A2(n6173), .ZN(n10558) );
  NAND2_X1 U5259 ( .A1(n8107), .A2(n8108), .ZN(n8195) );
  NAND4_X1 U5260 ( .A1(n6737), .A2(n6736), .A3(n6735), .A4(n6734), .ZN(n9874)
         );
  NOR2_X1 U5261 ( .A1(n5531), .A2(n8800), .ZN(n5530) );
  AND4_X1 U5262 ( .A1(n6718), .A2(n6717), .A3(n6716), .A4(n6715), .ZN(n8971)
         );
  AND4_X1 U5263 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n9251)
         );
  NAND2_X1 U5264 ( .A1(n5975), .A2(n5974), .ZN(n8214) );
  AND4_X1 U5265 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n9230)
         );
  NAND2_X2 U5266 ( .A1(n7568), .A2(n11012), .ZN(n11015) );
  AND2_X1 U5267 ( .A1(n6762), .A2(n6761), .ZN(n7877) );
  NAND2_X1 U5268 ( .A1(n5915), .A2(n5914), .ZN(n8175) );
  NAND2_X1 U5269 ( .A1(n5328), .A2(n7489), .ZN(n7599) );
  INV_X1 U5270 ( .A(n7704), .ZN(n7335) );
  NAND2_X1 U5271 ( .A1(n9133), .A2(n9132), .ZN(n9272) );
  NAND2_X1 U5272 ( .A1(n5839), .A2(n5838), .ZN(n5854) );
  NAND4_X1 U5273 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n10211)
         );
  XNOR2_X1 U5274 ( .A(n6757), .B(n6756), .ZN(n9268) );
  NAND2_X1 U5275 ( .A1(n6324), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6325) );
  CLKBUF_X1 U5276 ( .A(n6275), .Z(n8259) );
  NAND4_X2 U5277 ( .A1(n6425), .A2(n6424), .A3(n6423), .A4(n6422), .ZN(n9334)
         );
  INV_X2 U5278 ( .A(n6065), .ZN(n8653) );
  NAND4_X1 U5279 ( .A1(n6412), .A2(n6411), .A3(n6410), .A4(n6409), .ZN(n9335)
         );
  XNOR2_X1 U5280 ( .A(n6269), .B(n9627), .ZN(n8818) );
  INV_X2 U5281 ( .A(n5789), .ZN(n5807) );
  NAND2_X1 U5282 ( .A1(n5123), .A2(n5349), .ZN(n5348) );
  AOI21_X1 U5283 ( .B1(n5713), .B2(n5621), .A(n5620), .ZN(n5619) );
  OR2_X2 U5284 ( .A1(n8645), .A2(n5736), .ZN(n6301) );
  NAND2_X1 U5285 ( .A1(n5326), .A2(n5746), .ZN(n5352) );
  NAND2_X1 U5286 ( .A1(n8645), .A2(n5736), .ZN(n6017) );
  INV_X1 U5287 ( .A(n5353), .ZN(n5349) );
  NAND2_X1 U5288 ( .A1(n6816), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6387) );
  AND2_X1 U5290 ( .A1(n10872), .A2(n10873), .ZN(n10875) );
  XNOR2_X1 U5291 ( .A(n5731), .B(n10658), .ZN(n8645) );
  NAND2_X1 U5292 ( .A1(n5745), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5326) );
  OR2_X1 U5293 ( .A1(n6369), .A2(n6521), .ZN(n6371) );
  XNOR2_X1 U5294 ( .A(n5734), .B(n5733), .ZN(n5736) );
  NAND2_X1 U5295 ( .A1(n10657), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5731) );
  OR2_X1 U5296 ( .A1(n6525), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6537) );
  AND2_X1 U5297 ( .A1(n6270), .A2(n6272), .ZN(n6267) );
  NOR2_X1 U5298 ( .A1(n5496), .A2(n6367), .ZN(n6369) );
  NAND3_X1 U5299 ( .A1(n6413), .A2(n6415), .A3(n5451), .ZN(n10886) );
  AND2_X1 U5300 ( .A1(n6364), .A2(n6382), .ZN(n5497) );
  INV_X1 U5301 ( .A(n5971), .ZN(n5726) );
  NOR2_X1 U5302 ( .A1(n6363), .A2(n6624), .ZN(n6364) );
  AND2_X1 U5303 ( .A1(n5708), .A2(n5746), .ZN(n5547) );
  AND2_X1 U5304 ( .A1(n6358), .A2(n6359), .ZN(n5701) );
  AND4_X2 U5305 ( .A1(n9627), .A2(n6272), .A3(n6263), .A4(n6343), .ZN(n5706)
         );
  AND2_X1 U5306 ( .A1(n6414), .A2(n6356), .ZN(n5658) );
  NOR2_X2 U5307 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6395) );
  INV_X1 U5308 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6453) );
  INV_X1 U5309 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6414) );
  INV_X1 U5310 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6753) );
  INV_X1 U5311 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6263) );
  INV_X1 U5312 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6272) );
  INV_X1 U5313 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6031) );
  INV_X1 U5314 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6386) );
  INV_X1 U5315 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6593) );
  INV_X1 U5316 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6581) );
  INV_X1 U5317 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6358) );
  INV_X1 U5318 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6484) );
  OAI21_X2 U5319 ( .B1(n9926), .B2(n5485), .A(n5169), .ZN(n9896) );
  AND2_X1 U5320 ( .A1(n11110), .A2(n7849), .ZN(n5329) );
  NOR2_X4 U5321 ( .A1(n7746), .A2(n7866), .ZN(n7849) );
  OAI21_X2 U5322 ( .B1(n7064), .B2(n7063), .A(n10057), .ZN(n10124) );
  CLKBUF_X1 U5323 ( .A(n6314), .Z(n5122) );
  OAI211_X1 U5324 ( .C1(n5777), .C2(n7231), .A(n5760), .B(n5759), .ZN(n6314)
         );
  OAI21_X2 U5325 ( .B1(n5947), .B2(n5946), .A(n5945), .ZN(n5970) );
  NOR2_X1 U5326 ( .A1(n7531), .A2(n6421), .ZN(n7530) );
  NOR2_X2 U5327 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(n6631), .ZN(n6646) );
  AOI21_X2 U5328 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n9380), .A(n9374), .ZN(
        n8593) );
  NAND2_X4 U5329 ( .A1(n6373), .A2(n6377), .ZN(n6701) );
  AND2_X1 U5330 ( .A1(n8996), .A2(n8635), .ZN(n6601) );
  NAND2_X1 U5331 ( .A1(n10748), .A2(n6311), .ZN(n5777) );
  OR2_X1 U5332 ( .A1(n8777), .A2(n5628), .ZN(n5759) );
  NOR2_X2 U5333 ( .A1(n6561), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6571) );
  NOR2_X2 U5334 ( .A1(n6537), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6548) );
  OR2_X1 U5335 ( .A1(n8739), .A2(n8738), .ZN(n8746) );
  OR2_X1 U5336 ( .A1(n7339), .A2(n7761), .ZN(n7141) );
  INV_X1 U5337 ( .A(n6813), .ZN(n6803) );
  OR2_X1 U5338 ( .A1(n10612), .A2(n8303), .ZN(n8663) );
  AOI21_X1 U5339 ( .B1(n5125), .B2(n5145), .A(n5218), .ZN(n5217) );
  INV_X1 U5340 ( .A(n8345), .ZN(n5218) );
  AND4_X1 U5341 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(n8542)
         );
  INV_X1 U5342 ( .A(n6065), .ZN(n6305) );
  INV_X1 U5343 ( .A(n5903), .ZN(n6065) );
  OAI21_X1 U5344 ( .B1(n7949), .B2(n5529), .A(n5527), .ZN(n8318) );
  AOI21_X1 U5345 ( .B1(n5530), .B2(n5528), .A(n5157), .ZN(n5527) );
  INV_X1 U5346 ( .A(n5530), .ZN(n5529) );
  AND2_X1 U5347 ( .A1(n8749), .A2(n5362), .ZN(n5361) );
  NAND2_X1 U5348 ( .A1(n5363), .A2(n8744), .ZN(n5362) );
  NAND2_X1 U5349 ( .A1(n8756), .A2(n8815), .ZN(n5381) );
  INV_X1 U5350 ( .A(n6282), .ZN(n8690) );
  AOI21_X1 U5351 ( .B1(n7376), .B2(n8667), .A(n6290), .ZN(n8669) );
  INV_X1 U5352 ( .A(SI_15_), .ZN(n9656) );
  NAND2_X1 U5353 ( .A1(n5969), .A2(n5968), .ZN(n5305) );
  AND2_X1 U5354 ( .A1(n5130), .A2(n5311), .ZN(n5312) );
  INV_X1 U5355 ( .A(n5856), .ZN(n5245) );
  OR2_X1 U5356 ( .A1(n9906), .A2(n9914), .ZN(n5435) );
  OR2_X1 U5357 ( .A1(n10032), .A2(n8950), .ZN(n9118) );
  INV_X1 U5358 ( .A(n5420), .ZN(n5417) );
  NAND2_X1 U5359 ( .A1(n9268), .A2(n9409), .ZN(n7344) );
  AND2_X1 U5360 ( .A1(n6357), .A2(n6395), .ZN(n5231) );
  AND2_X1 U5361 ( .A1(n7055), .A2(n7061), .ZN(n5587) );
  INV_X1 U5362 ( .A(n5515), .ZN(n5512) );
  NOR2_X1 U5363 ( .A1(n10197), .A2(n10598), .ZN(n5334) );
  NAND2_X1 U5364 ( .A1(n5239), .A2(n5240), .ZN(n5237) );
  NOR2_X1 U5365 ( .A1(n8175), .A2(n7946), .ZN(n5331) );
  NOR2_X1 U5366 ( .A1(n5541), .A2(n5538), .ZN(n5539) );
  AND2_X1 U5367 ( .A1(n8687), .A2(n5501), .ZN(n5128) );
  NAND2_X1 U5368 ( .A1(n5502), .A2(n5869), .ZN(n5501) );
  INV_X1 U5369 ( .A(n8680), .ZN(n5502) );
  INV_X1 U5370 ( .A(n5869), .ZN(n5503) );
  NAND2_X1 U5371 ( .A1(n6134), .A2(n6133), .ZN(n6148) );
  OR2_X1 U5372 ( .A1(n5970), .A2(n5304), .ZN(n5300) );
  NAND2_X1 U5373 ( .A1(n5221), .A2(n8281), .ZN(n5220) );
  NOR2_X1 U5374 ( .A1(n8341), .A2(n8288), .ZN(n8342) );
  INV_X1 U5375 ( .A(n8343), .ZN(n5221) );
  NAND2_X1 U5376 ( .A1(n9016), .A2(n5235), .ZN(n5234) );
  INV_X1 U5377 ( .A(n8952), .ZN(n5235) );
  INV_X1 U5378 ( .A(n9034), .ZN(n5228) );
  NAND2_X1 U5379 ( .A1(n5289), .A2(n9268), .ZN(n5288) );
  INV_X1 U5380 ( .A(n9269), .ZN(n5290) );
  AND4_X1 U5381 ( .A1(n6674), .A2(n6673), .A3(n6672), .A4(n6671), .ZN(n9068)
         );
  NAND2_X1 U5382 ( .A1(n6395), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U5383 ( .A1(n5473), .A2(n5472), .ZN(n5471) );
  INV_X1 U5384 ( .A(n9339), .ZN(n5472) );
  NAND2_X1 U5385 ( .A1(n9103), .A2(n9102), .ZN(n9306) );
  NAND2_X1 U5386 ( .A1(n9892), .A2(n5431), .ZN(n9891) );
  OR2_X1 U5387 ( .A1(n5485), .A2(n9115), .ZN(n5484) );
  NAND2_X1 U5388 ( .A1(n5486), .A2(n9240), .ZN(n5485) );
  OR2_X1 U5389 ( .A1(n10020), .A2(n9068), .ZN(n9226) );
  NAND2_X1 U5390 ( .A1(n6770), .A2(n5494), .ZN(n5493) );
  NOR2_X1 U5391 ( .A1(n5495), .A2(n6771), .ZN(n5494) );
  INV_X1 U5392 ( .A(n9205), .ZN(n5495) );
  AND2_X1 U5393 ( .A1(n9118), .A2(n9116), .ZN(n9296) );
  OR2_X1 U5394 ( .A1(n11144), .A2(n8539), .ZN(n9205) );
  NAND2_X1 U5395 ( .A1(n7970), .A2(n7896), .ZN(n9165) );
  INV_X1 U5396 ( .A(n9101), .ZN(n6642) );
  INV_X1 U5397 ( .A(n7153), .ZN(n6641) );
  AND2_X1 U5398 ( .A1(n5410), .A2(n9278), .ZN(n5409) );
  NAND2_X1 U5399 ( .A1(n7153), .A2(n5120), .ZN(n6466) );
  AND2_X1 U5400 ( .A1(n6838), .A2(n5703), .ZN(n5702) );
  XNOR2_X1 U5401 ( .A(n9992), .B(n9874), .ZN(n9448) );
  NAND2_X1 U5402 ( .A1(n9120), .A2(n8237), .ZN(n11127) );
  NAND2_X1 U5403 ( .A1(n6818), .A2(n6838), .ZN(n6822) );
  NAND2_X1 U5404 ( .A1(n6805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6807) );
  INV_X1 U5405 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6806) );
  AND2_X1 U5406 ( .A1(n6852), .A2(n7577), .ZN(n6853) );
  NOR2_X1 U5407 ( .A1(n10174), .A2(n10175), .ZN(n5571) );
  OR2_X1 U5408 ( .A1(n8784), .A2(n5341), .ZN(n8817) );
  NOR3_X1 U5409 ( .A1(n8783), .A2(n10620), .A3(n8810), .ZN(n8784) );
  OAI21_X1 U5410 ( .B1(n5346), .B2(n5342), .A(n8842), .ZN(n5341) );
  NOR2_X1 U5411 ( .A1(n6259), .A2(n5525), .ZN(n5524) );
  INV_X1 U5412 ( .A(n6244), .ZN(n5525) );
  INV_X1 U5413 ( .A(n5204), .ZN(n6250) );
  NAND2_X1 U5414 ( .A1(n10352), .A2(n10628), .ZN(n10341) );
  OAI22_X1 U5415 ( .A1(n10387), .A2(n6183), .B1(n10416), .B2(n10558), .ZN(
        n10369) );
  NAND2_X1 U5416 ( .A1(n10462), .A2(n5309), .ZN(n8831) );
  NOR2_X1 U5417 ( .A1(n8742), .A2(n5310), .ZN(n5309) );
  INV_X1 U5418 ( .A(n8740), .ZN(n5310) );
  OR2_X1 U5419 ( .A1(n10578), .A2(n10081), .ZN(n8740) );
  AOI21_X1 U5420 ( .B1(n8803), .B2(n5507), .A(n5143), .ZN(n5506) );
  INV_X1 U5421 ( .A(n6022), .ZN(n5507) );
  INV_X1 U5422 ( .A(n8803), .ZN(n5508) );
  NAND2_X1 U5423 ( .A1(n8380), .A2(n8893), .ZN(n5398) );
  INV_X1 U5424 ( .A(n5535), .ZN(n5531) );
  NAND2_X1 U5425 ( .A1(n7949), .A2(n5533), .ZN(n5532) );
  NAND2_X1 U5426 ( .A1(n6300), .A2(n6299), .ZN(n10512) );
  INV_X1 U5427 ( .A(n10539), .ZN(n5197) );
  OAI21_X1 U5428 ( .B1(n6101), .B2(n6100), .A(n6099), .ZN(n6117) );
  AND2_X1 U5429 ( .A1(n6118), .A2(n6104), .ZN(n6116) );
  NAND2_X1 U5430 ( .A1(n6256), .A2(n6255), .ZN(n10338) );
  NAND2_X1 U5431 ( .A1(n9198), .A2(n5281), .ZN(n5280) );
  INV_X1 U5432 ( .A(n5282), .ZN(n5281) );
  OAI21_X1 U5433 ( .B1(n6579), .B2(n9199), .A(n9197), .ZN(n5282) );
  OR2_X1 U5434 ( .A1(n8891), .A2(n8815), .ZN(n5396) );
  INV_X1 U5435 ( .A(n5396), .ZN(n5392) );
  NAND2_X1 U5436 ( .A1(n5285), .A2(n5283), .ZN(n9198) );
  AND2_X1 U5437 ( .A1(n9289), .A2(n5284), .ZN(n5283) );
  NAND2_X1 U5438 ( .A1(n9188), .A2(n9187), .ZN(n5285) );
  NAND2_X1 U5439 ( .A1(n9119), .A2(n9244), .ZN(n5284) );
  NAND2_X1 U5440 ( .A1(n5272), .A2(n5277), .ZN(n5269) );
  NAND2_X1 U5441 ( .A1(n5273), .A2(n5153), .ZN(n5272) );
  AND2_X1 U5442 ( .A1(n9234), .A2(n9233), .ZN(n5277) );
  NOR2_X1 U5443 ( .A1(n9229), .A2(n5276), .ZN(n5275) );
  NOR2_X1 U5444 ( .A1(n5367), .A2(n5366), .ZN(n5365) );
  INV_X1 U5445 ( .A(n8751), .ZN(n5367) );
  INV_X1 U5446 ( .A(n5361), .ZN(n5360) );
  AND2_X1 U5447 ( .A1(n9262), .A2(n9261), .ZN(n5296) );
  INV_X1 U5448 ( .A(n6684), .ZN(n5448) );
  NAND2_X1 U5449 ( .A1(n6992), .A2(n5558), .ZN(n5557) );
  INV_X1 U5450 ( .A(n6990), .ZN(n5558) );
  INV_X1 U5451 ( .A(n8389), .ZN(n5559) );
  AND2_X1 U5452 ( .A1(n5177), .A2(n6980), .ZN(n5553) );
  NAND2_X1 U5453 ( .A1(n5378), .A2(n10336), .ZN(n5377) );
  NAND2_X1 U5454 ( .A1(n5379), .A2(n8760), .ZN(n5378) );
  NAND2_X1 U5455 ( .A1(n8701), .A2(n7840), .ZN(n6282) );
  INV_X1 U5456 ( .A(n6245), .ZN(n5614) );
  INV_X1 U5457 ( .A(n5314), .ZN(n5313) );
  INV_X1 U5458 ( .A(SI_10_), .ZN(n9698) );
  NAND2_X1 U5459 ( .A1(n5622), .A2(n5893), .ZN(n5268) );
  AND2_X1 U5460 ( .A1(n7342), .A2(n9313), .ZN(n5127) );
  NAND2_X1 U5461 ( .A1(n8958), .A2(n9946), .ZN(n5670) );
  NAND2_X1 U5462 ( .A1(n10886), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7406) );
  NOR2_X1 U5463 ( .A1(n7512), .A2(n5596), .ZN(n7692) );
  NOR2_X1 U5464 ( .A1(n7410), .A2(n6434), .ZN(n5596) );
  NOR2_X1 U5465 ( .A1(n8097), .A2(n8096), .ZN(n8188) );
  AND2_X1 U5466 ( .A1(n8103), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8096) );
  AND2_X1 U5467 ( .A1(n5434), .A2(n5435), .ZN(n5429) );
  OR2_X1 U5468 ( .A1(n10028), .A2(n8954), .ZN(n9221) );
  OR2_X1 U5469 ( .A1(n11138), .A2(n8467), .ZN(n9201) );
  AND2_X1 U5470 ( .A1(n9195), .A2(n5142), .ZN(n5489) );
  NAND2_X1 U5471 ( .A1(n5261), .A2(n5260), .ZN(n9154) );
  NOR2_X1 U5472 ( .A1(n9332), .A2(n7617), .ZN(n5416) );
  NOR2_X1 U5473 ( .A1(n5421), .A2(n6444), .ZN(n5420) );
  INV_X1 U5474 ( .A(n6432), .ZN(n5421) );
  OR2_X1 U5475 ( .A1(n7342), .A2(n9268), .ZN(n9271) );
  AOI21_X1 U5476 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_20__SCAN_IN), .ZN(n5686) );
  XNOR2_X1 U5477 ( .A(n6869), .B(n5119), .ZN(n6872) );
  NOR2_X1 U5478 ( .A1(n6036), .A2(n8022), .ZN(n5206) );
  NOR2_X1 U5479 ( .A1(n5976), .A2(n8301), .ZN(n5205) );
  INV_X1 U5480 ( .A(n8877), .ZN(n8793) );
  NAND2_X1 U5481 ( .A1(n8785), .A2(n5144), .ZN(n8789) );
  INV_X1 U5482 ( .A(n8781), .ZN(n5347) );
  NAND2_X1 U5483 ( .A1(n5345), .A2(n5343), .ZN(n5342) );
  AOI21_X1 U5484 ( .B1(n10320), .B2(n8815), .A(n5344), .ZN(n5343) );
  AND2_X1 U5485 ( .A1(n10201), .A2(n10313), .ZN(n5344) );
  NOR2_X1 U5486 ( .A1(n8939), .A2(n5403), .ZN(n5402) );
  NOR2_X1 U5487 ( .A1(n8809), .A2(n8834), .ZN(n5404) );
  NOR2_X1 U5488 ( .A1(n6233), .A2(n6232), .ZN(n5204) );
  NOR2_X1 U5489 ( .A1(n6108), .A2(n6107), .ZN(n5207) );
  INV_X1 U5490 ( .A(n5325), .ZN(n5248) );
  NAND2_X1 U5491 ( .A1(n5206), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6063) );
  INV_X1 U5492 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6062) );
  NOR2_X1 U5493 ( .A1(n5984), .A2(n5534), .ZN(n5533) );
  INV_X1 U5494 ( .A(n5964), .ZN(n5534) );
  AND2_X1 U5495 ( .A1(n6292), .A2(n5132), .ZN(n5239) );
  NAND2_X1 U5496 ( .A1(n5253), .A2(n10207), .ZN(n7840) );
  NOR2_X1 U5497 ( .A1(n6289), .A2(n5376), .ZN(n5375) );
  INV_X1 U5498 ( .A(n8868), .ZN(n5376) );
  NAND2_X1 U5499 ( .A1(n5371), .A2(n5141), .ZN(n8870) );
  INV_X1 U5500 ( .A(n7303), .ZN(n5371) );
  NAND2_X1 U5501 ( .A1(n6858), .A2(n10932), .ZN(n5542) );
  NAND2_X1 U5502 ( .A1(n5327), .A2(n5546), .ZN(n5745) );
  INV_X1 U5503 ( .A(n6266), .ZN(n5327) );
  NAND2_X1 U5504 ( .A1(n5643), .A2(n6221), .ZN(n6228) );
  NAND2_X1 U5505 ( .A1(n5640), .A2(n5638), .ZN(n5643) );
  NOR2_X1 U5506 ( .A1(n6222), .A2(n5639), .ZN(n5638) );
  INV_X1 U5507 ( .A(n6204), .ZN(n5639) );
  NOR2_X1 U5508 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6317) );
  OAI21_X1 U5509 ( .B1(n6148), .B2(n5647), .A(n5645), .ZN(n6185) );
  AOI21_X1 U5510 ( .B1(n6146), .B2(n5648), .A(n5646), .ZN(n5645) );
  INV_X1 U5511 ( .A(n5648), .ZN(n5647) );
  INV_X1 U5512 ( .A(n6168), .ZN(n5646) );
  AND2_X1 U5513 ( .A1(n6186), .A2(n6172), .ZN(n6184) );
  INV_X1 U5514 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6264) );
  OAI21_X1 U5515 ( .B1(n6008), .B2(n5654), .A(n5652), .ZN(n6055) );
  INV_X1 U5516 ( .A(n5653), .ZN(n5652) );
  OAI21_X1 U5517 ( .B1(n5656), .B2(n5654), .A(n6040), .ZN(n5653) );
  NAND2_X1 U5518 ( .A1(n5655), .A2(n6027), .ZN(n5654) );
  AND2_X1 U5519 ( .A1(n6056), .A2(n6045), .ZN(n6054) );
  AOI21_X1 U5520 ( .B1(n5303), .B2(n5302), .A(n5170), .ZN(n5301) );
  INV_X1 U5521 ( .A(n5968), .ZN(n5302) );
  INV_X1 U5522 ( .A(n5912), .ZN(n5620) );
  NOR2_X2 U5523 ( .A1(n5891), .A2(n5315), .ZN(n5314) );
  INV_X1 U5524 ( .A(n5874), .ZN(n5315) );
  OAI211_X1 U5525 ( .C1(n5245), .C2(n5853), .A(n5241), .B(n5871), .ZN(n5316)
         );
  NAND2_X1 U5526 ( .A1(n5839), .A2(n5242), .ZN(n5241) );
  NOR2_X1 U5527 ( .A1(n5245), .A2(n5243), .ZN(n5242) );
  NAND2_X1 U5528 ( .A1(n5627), .A2(n5626), .ZN(n5770) );
  OAI21_X1 U5529 ( .B1(n5629), .B2(n5628), .A(n5624), .ZN(n5623) );
  NAND2_X1 U5530 ( .A1(n5677), .A2(n5676), .ZN(n7816) );
  NOR2_X1 U5531 ( .A1(n7731), .A2(n5672), .ZN(n5677) );
  INV_X1 U5532 ( .A(n7733), .ZN(n5672) );
  OR2_X1 U5533 ( .A1(n5667), .A2(n9052), .ZN(n5666) );
  INV_X1 U5534 ( .A(n5670), .ZN(n5667) );
  OR2_X1 U5535 ( .A1(n8965), .A2(n8964), .ZN(n8966) );
  OR2_X1 U5536 ( .A1(n8955), .A2(n8954), .ZN(n8956) );
  OR2_X1 U5537 ( .A1(n8567), .A2(n5695), .ZN(n5694) );
  OR2_X1 U5538 ( .A1(n8567), .A2(n5189), .ZN(n5690) );
  INV_X1 U5539 ( .A(n8554), .ZN(n5691) );
  INV_X1 U5540 ( .A(n5694), .ZN(n5692) );
  NAND2_X1 U5541 ( .A1(n8564), .A2(n5697), .ZN(n5695) );
  AND2_X1 U5542 ( .A1(n8966), .A2(n8968), .ZN(n5698) );
  INV_X1 U5543 ( .A(n9044), .ZN(n8968) );
  INV_X1 U5544 ( .A(n8469), .ZN(n5214) );
  INV_X1 U5545 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U5546 ( .A1(n6365), .A2(n6364), .ZN(n6813) );
  OR2_X1 U5547 ( .A1(n7405), .A2(n7404), .ZN(n10873) );
  OR2_X1 U5548 ( .A1(n10880), .A2(n7395), .ZN(n5590) );
  INV_X1 U5549 ( .A(n7394), .ZN(n7395) );
  NAND2_X1 U5550 ( .A1(n5462), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5459) );
  XNOR2_X1 U5551 ( .A(n7692), .B(n7693), .ZN(n7513) );
  NOR2_X1 U5552 ( .A1(n7513), .A2(n6445), .ZN(n7694) );
  XNOR2_X1 U5553 ( .A(n8188), .B(n8193), .ZN(n8098) );
  AND2_X1 U5554 ( .A1(n5209), .A2(n5208), .ZN(n8183) );
  NAND2_X1 U5555 ( .A1(n8103), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5208) );
  INV_X1 U5556 ( .A(n8094), .ZN(n5209) );
  AND2_X1 U5557 ( .A1(n5593), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U5558 ( .A1(n10909), .A2(n10910), .ZN(n10908) );
  INV_X1 U5559 ( .A(n5456), .ZN(n5455) );
  NAND2_X1 U5560 ( .A1(n9363), .A2(n9364), .ZN(n9362) );
  OR2_X1 U5561 ( .A1(n9359), .A2(n8599), .ZN(n5600) );
  AOI21_X1 U5562 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9380), .A(n9376), .ZN(
        n8582) );
  NAND2_X1 U5563 ( .A1(n9900), .A2(n5429), .ZN(n5422) );
  NAND2_X1 U5564 ( .A1(n5428), .A2(n5434), .ZN(n5427) );
  INV_X1 U5565 ( .A(n5430), .ZN(n5428) );
  AOI21_X1 U5566 ( .B1(n9899), .B2(n5435), .A(n5431), .ZN(n5430) );
  OAI21_X1 U5567 ( .B1(n9900), .B2(n5426), .A(n5423), .ZN(n9872) );
  AOI21_X1 U5568 ( .B1(n5427), .B2(n5425), .A(n5424), .ZN(n5423) );
  INV_X1 U5569 ( .A(n5427), .ZN(n5426) );
  INV_X1 U5570 ( .A(n5429), .ZN(n5425) );
  NAND2_X1 U5571 ( .A1(n6774), .A2(n9899), .ZN(n9898) );
  NAND2_X1 U5572 ( .A1(n5479), .A2(n5481), .ZN(n9938) );
  NOR2_X1 U5573 ( .A1(n9932), .A2(n5482), .ZN(n5481) );
  NOR2_X1 U5574 ( .A1(n9952), .A2(n5483), .ZN(n5482) );
  AOI21_X1 U5575 ( .B1(n5440), .B2(n5442), .A(n5164), .ZN(n5439) );
  INV_X1 U5576 ( .A(n9944), .ZN(n9952) );
  NAND2_X1 U5577 ( .A1(n6772), .A2(n9223), .ZN(n9953) );
  NAND2_X1 U5578 ( .A1(n9953), .A2(n9952), .ZN(n9951) );
  NAND2_X1 U5579 ( .A1(n9960), .A2(n6664), .ZN(n9959) );
  AND4_X1 U5580 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n8539)
         );
  AND4_X1 U5581 ( .A1(n6565), .A2(n6564), .A3(n6563), .A4(n6562), .ZN(n8414)
         );
  INV_X1 U5582 ( .A(n9326), .ZN(n8331) );
  NOR2_X1 U5583 ( .A1(n9279), .A2(n9157), .ZN(n5478) );
  AND2_X1 U5584 ( .A1(n6491), .A2(n6490), .ZN(n7732) );
  NOR2_X1 U5585 ( .A1(n6458), .A2(n5419), .ZN(n5418) );
  INV_X1 U5586 ( .A(n6443), .ZN(n5419) );
  AOI21_X1 U5587 ( .B1(n5418), .B2(n5417), .A(n5416), .ZN(n5412) );
  NAND2_X1 U5588 ( .A1(n6433), .A2(n5420), .ZN(n5415) );
  OR2_X1 U5589 ( .A1(n9244), .A2(n9875), .ZN(n8523) );
  OR2_X1 U5590 ( .A1(n9244), .A2(n9902), .ZN(n8524) );
  AND2_X1 U5591 ( .A1(n6782), .A2(n7139), .ZN(n8157) );
  NOR2_X1 U5592 ( .A1(n11127), .A2(n7361), .ZN(n7363) );
  INV_X1 U5593 ( .A(n7143), .ZN(n7766) );
  NAND2_X1 U5594 ( .A1(n9872), .A2(n5432), .ZN(n9440) );
  NAND2_X1 U5595 ( .A1(n9996), .A2(n5433), .ZN(n5432) );
  NAND2_X1 U5596 ( .A1(n6687), .A2(n6686), .ZN(n10012) );
  OR2_X1 U5597 ( .A1(n9101), .A2(n7160), .ZN(n6417) );
  NOR2_X1 U5598 ( .A1(n7141), .A2(n7140), .ZN(n7362) );
  INV_X1 U5599 ( .A(n7192), .ZN(n7361) );
  INV_X1 U5600 ( .A(n5199), .ZN(n6367) );
  INV_X1 U5601 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6370) );
  OAI21_X1 U5602 ( .B1(n6640), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U5603 ( .A1(n6545), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6557) );
  AOI21_X1 U5604 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(n5700), .A(
        P2_IR_REG_11__SCAN_IN), .ZN(n5699) );
  INV_X1 U5605 ( .A(n5701), .ZN(n5700) );
  INV_X1 U5606 ( .A(n6395), .ZN(n7321) );
  NAND2_X1 U5607 ( .A1(n5205), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6014) );
  INV_X1 U5608 ( .A(n10069), .ZN(n5548) );
  NAND2_X1 U5609 ( .A1(n7001), .A2(n10185), .ZN(n10097) );
  NAND2_X1 U5610 ( .A1(n10097), .A2(n10098), .ZN(n10096) );
  INV_X1 U5611 ( .A(n5562), .ZN(n5561) );
  OAI21_X1 U5612 ( .B1(n10098), .B2(n5563), .A(n10109), .ZN(n5562) );
  NOR2_X1 U5613 ( .A1(n5589), .A2(n10143), .ZN(n5585) );
  NAND2_X1 U5614 ( .A1(n5584), .A2(n5589), .ZN(n5583) );
  OR2_X1 U5615 ( .A1(n5568), .A2(n10163), .ZN(n5567) );
  NOR2_X1 U5616 ( .A1(n5159), .A2(n5565), .ZN(n5564) );
  OR2_X1 U5617 ( .A1(n6847), .A2(n10749), .ZN(n5707) );
  NAND2_X1 U5618 ( .A1(n10079), .A2(n5587), .ZN(n10140) );
  NAND2_X1 U5619 ( .A1(n5580), .A2(n5589), .ZN(n5588) );
  NAND2_X1 U5620 ( .A1(n10079), .A2(n7055), .ZN(n5580) );
  INV_X1 U5621 ( .A(n8169), .ZN(n5577) );
  AND2_X1 U5622 ( .A1(n6958), .A2(n5577), .ZN(n5576) );
  XNOR2_X1 U5623 ( .A(n6879), .B(n7089), .ZN(n6884) );
  XNOR2_X1 U5624 ( .A(n6273), .B(n6272), .ZN(n8921) );
  AND2_X1 U5625 ( .A1(n6275), .A2(n8921), .ZN(n8919) );
  NAND2_X1 U5626 ( .A1(n5545), .A2(n8645), .ZN(n5789) );
  NAND3_X1 U5627 ( .A1(n5752), .A2(n5751), .A3(n5750), .ZN(n5541) );
  OAI21_X1 U5628 ( .B1(n6301), .B2(n5737), .A(n5544), .ZN(n5551) );
  NAND2_X1 U5629 ( .A1(n8764), .A2(n8763), .ZN(n10538) );
  OR2_X1 U5630 ( .A1(n10334), .A2(n10336), .ZN(n5526) );
  NAND2_X1 U5631 ( .A1(n10335), .A2(n5404), .ZN(n5308) );
  AND2_X1 U5632 ( .A1(n8809), .A2(n5252), .ZN(n5251) );
  NAND2_X1 U5633 ( .A1(n5403), .A2(n6298), .ZN(n5252) );
  NOR2_X1 U5634 ( .A1(n10370), .A2(n10353), .ZN(n10352) );
  NAND2_X1 U5635 ( .A1(n10394), .A2(n10636), .ZN(n10370) );
  INV_X1 U5636 ( .A(n6190), .ZN(n6191) );
  OAI21_X1 U5637 ( .B1(n10401), .B2(n6166), .A(n6167), .ZN(n10387) );
  NAND2_X1 U5638 ( .A1(n8831), .A2(n5156), .ZN(n10432) );
  NAND2_X1 U5639 ( .A1(n10471), .A2(n8899), .ZN(n10462) );
  AOI21_X1 U5640 ( .B1(n8733), .B2(n5516), .A(n5160), .ZN(n5515) );
  INV_X1 U5641 ( .A(n6073), .ZN(n5516) );
  AND2_X1 U5642 ( .A1(n8740), .A2(n10438), .ZN(n10463) );
  NAND2_X1 U5643 ( .A1(n10486), .A2(n6072), .ZN(n6074) );
  NAND2_X1 U5644 ( .A1(n10472), .A2(n5517), .ZN(n10471) );
  NAND2_X1 U5645 ( .A1(n5505), .A2(n5504), .ZN(n10513) );
  AOI21_X1 U5646 ( .B1(n5506), .B2(n5508), .A(n8804), .ZN(n5504) );
  NAND2_X1 U5647 ( .A1(n8321), .A2(n6294), .ZN(n8380) );
  AND2_X1 U5648 ( .A1(n5536), .A2(n5983), .ZN(n5535) );
  OR2_X1 U5649 ( .A1(n5537), .A2(n5984), .ZN(n5536) );
  NAND2_X1 U5650 ( .A1(n5965), .A2(n5964), .ZN(n5537) );
  AND2_X1 U5651 ( .A1(n8663), .A2(n8664), .ZN(n8800) );
  NAND2_X1 U5652 ( .A1(n5954), .A2(n5953), .ZN(n7956) );
  NAND2_X1 U5653 ( .A1(n5944), .A2(n5943), .ZN(n7949) );
  AOI21_X1 U5654 ( .B1(n5520), .B2(n5522), .A(n5152), .ZN(n5518) );
  NAND2_X1 U5655 ( .A1(n7849), .A2(n5331), .ZN(n7920) );
  NAND2_X1 U5656 ( .A1(n5500), .A2(n5499), .ZN(n7848) );
  AOI21_X1 U5657 ( .B1(n5128), .B2(n5503), .A(n5162), .ZN(n5499) );
  NAND2_X1 U5658 ( .A1(n7745), .A2(n8680), .ZN(n7744) );
  NAND2_X1 U5659 ( .A1(n8870), .A2(n8868), .ZN(n8665) );
  XNOR2_X1 U5660 ( .A(n10213), .B(n7335), .ZN(n8786) );
  INV_X1 U5661 ( .A(n8944), .ZN(n10509) );
  NAND2_X1 U5662 ( .A1(n10538), .A2(n10996), .ZN(n5338) );
  NAND2_X1 U5663 ( .A1(n6231), .A2(n6230), .ZN(n10344) );
  NAND2_X1 U5664 ( .A1(n5306), .A2(n6035), .ZN(n10598) );
  NAND2_X1 U5665 ( .A1(n7629), .A2(n5948), .ZN(n5306) );
  AND2_X1 U5666 ( .A1(n10933), .A2(n8921), .ZN(n10599) );
  INV_X1 U5667 ( .A(n10599), .ZN(n11049) );
  AND2_X1 U5668 ( .A1(n8359), .A2(n10616), .ZN(n11000) );
  AND2_X1 U5669 ( .A1(n6327), .A2(n6326), .ZN(n7182) );
  NAND2_X1 U5670 ( .A1(n6847), .A2(n7190), .ZN(n8851) );
  NAND2_X1 U5671 ( .A1(n8640), .A2(n8639), .ZN(n8656) );
  OR2_X1 U5672 ( .A1(n8638), .A2(n8637), .ZN(n8639) );
  OR2_X1 U5673 ( .A1(n8636), .A2(n9661), .ZN(n8640) );
  XNOR2_X1 U5674 ( .A(n8656), .B(n8655), .ZN(n9097) );
  NOR2_X1 U5675 ( .A1(n6154), .A2(n5649), .ZN(n5648) );
  INV_X1 U5676 ( .A(n6150), .ZN(n5649) );
  NAND2_X1 U5677 ( .A1(n6148), .A2(n6147), .ZN(n5650) );
  NAND2_X1 U5678 ( .A1(n5644), .A2(n6118), .ZN(n6130) );
  XNOR2_X1 U5679 ( .A(n6042), .B(n6041), .ZN(n7629) );
  NAND2_X1 U5680 ( .A1(n5651), .A2(n6027), .ZN(n6042) );
  NAND2_X1 U5681 ( .A1(n6008), .A2(n5656), .ZN(n5651) );
  NAND2_X1 U5682 ( .A1(n6008), .A2(n6007), .ZN(n6025) );
  INV_X1 U5683 ( .A(n6823), .ZN(n6840) );
  XNOR2_X1 U5684 ( .A(n8963), .B(n8964), .ZN(n9009) );
  NAND2_X1 U5685 ( .A1(n9009), .A2(n9934), .ZN(n9008) );
  OR2_X1 U5686 ( .A1(n8953), .A2(n5234), .ZN(n9015) );
  AOI21_X1 U5687 ( .B1(n5680), .B2(n5682), .A(n8977), .ZN(n5679) );
  NAND2_X1 U5688 ( .A1(n6729), .A2(n6728), .ZN(n9992) );
  NAND2_X1 U5689 ( .A1(n6710), .A2(n6709), .ZN(n9906) );
  AND4_X1 U5690 ( .A1(n6498), .A2(n6497), .A3(n6496), .A4(n6495), .ZN(n7896)
         );
  INV_X1 U5691 ( .A(n9972), .ZN(n10024) );
  NAND2_X1 U5692 ( .A1(n5233), .A2(n5155), .ZN(n9063) );
  NAND2_X1 U5693 ( .A1(n8953), .A2(n5661), .ZN(n5233) );
  AOI21_X1 U5694 ( .B1(n5661), .B2(n5663), .A(n5660), .ZN(n5659) );
  NAND2_X1 U5695 ( .A1(n9306), .A2(n9435), .ZN(n5286) );
  INV_X1 U5696 ( .A(n8971), .ZN(n9914) );
  OAI21_X1 U5697 ( .B1(n7681), .B2(n5464), .A(n5463), .ZN(n8094) );
  NAND2_X1 U5698 ( .A1(n5465), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U5699 ( .A1(n7987), .A2(n5465), .ZN(n5463) );
  INV_X1 U5700 ( .A(n7989), .ZN(n5465) );
  XNOR2_X1 U5701 ( .A(n8183), .B(n8193), .ZN(n8095) );
  OR2_X1 U5702 ( .A1(n8577), .A2(n8578), .ZN(n5473) );
  INV_X1 U5703 ( .A(n5471), .ZN(n9338) );
  NAND2_X1 U5704 ( .A1(n6720), .A2(n6719), .ZN(n10000) );
  AND2_X1 U5705 ( .A1(n9296), .A2(n9213), .ZN(n5492) );
  NAND2_X1 U5706 ( .A1(n6798), .A2(n5710), .ZN(n5475) );
  OR2_X1 U5707 ( .A1(n8992), .A2(n11127), .ZN(n5710) );
  NAND2_X1 U5708 ( .A1(n6825), .A2(n6824), .ZN(n7761) );
  INV_X1 U5709 ( .A(n10441), .ZN(n10082) );
  OR2_X1 U5710 ( .A1(n7094), .A2(n7095), .ZN(n5570) );
  AND2_X1 U5711 ( .A1(n7127), .A2(n11097), .ZN(n5569) );
  NAND2_X1 U5712 ( .A1(n7197), .A2(n5948), .ZN(n5901) );
  NAND2_X1 U5713 ( .A1(n6106), .A2(n6105), .ZN(n10578) );
  AND2_X1 U5714 ( .A1(n7100), .A2(n7101), .ZN(n11097) );
  INV_X1 U5715 ( .A(n10183), .ZN(n11088) );
  INV_X1 U5716 ( .A(n8259), .ZN(n8923) );
  NAND2_X1 U5717 ( .A1(n6241), .A2(n6240), .ZN(n10363) );
  AOI21_X1 U5718 ( .B1(n8947), .B2(n10512), .A(n5184), .ZN(n10539) );
  XNOR2_X1 U5719 ( .A(n5339), .B(n8940), .ZN(n10540) );
  AOI21_X1 U5720 ( .B1(n5524), .B2(n10336), .A(n5172), .ZN(n5523) );
  NAND2_X1 U5721 ( .A1(n5524), .A2(n10334), .ZN(n5340) );
  AND2_X1 U5722 ( .A1(n8661), .A2(n8660), .ZN(n10620) );
  NAND2_X1 U5723 ( .A1(n6248), .A2(n6247), .ZN(n10325) );
  NAND2_X1 U5724 ( .A1(n5255), .A2(n5321), .ZN(n6355) );
  NOR2_X1 U5725 ( .A1(n10330), .A2(n10329), .ZN(n5255) );
  INV_X1 U5726 ( .A(n5322), .ZN(n5321) );
  NOR2_X1 U5727 ( .A1(n10333), .A2(n11000), .ZN(n5322) );
  INV_X1 U5728 ( .A(n10344), .ZN(n10628) );
  CLKBUF_X1 U5729 ( .A(n6342), .Z(n6326) );
  AND2_X1 U5730 ( .A1(n7195), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7190) );
  NAND2_X1 U5731 ( .A1(n9153), .A2(n9154), .ZN(n5259) );
  NAND2_X1 U5732 ( .A1(n8693), .A2(n8692), .ZN(n8697) );
  NAND2_X1 U5733 ( .A1(n5258), .A2(n5256), .ZN(n9171) );
  INV_X1 U5734 ( .A(n5257), .ZN(n5256) );
  NAND2_X1 U5735 ( .A1(n5259), .A2(n5127), .ZN(n5258) );
  AOI21_X1 U5736 ( .B1(n9167), .B2(n9165), .A(n5127), .ZN(n5257) );
  OAI21_X1 U5737 ( .B1(n8725), .B2(n8891), .A(n8815), .ZN(n5393) );
  NAND2_X1 U5738 ( .A1(n5279), .A2(n5278), .ZN(n9210) );
  NAND2_X1 U5739 ( .A1(n9200), .A2(n5127), .ZN(n5278) );
  NAND2_X1 U5740 ( .A1(n5280), .A2(n9244), .ZN(n5279) );
  AND2_X1 U5741 ( .A1(n8723), .A2(n5384), .ZN(n5390) );
  NOR2_X1 U5742 ( .A1(n5393), .A2(n8815), .ZN(n5384) );
  OAI21_X1 U5743 ( .B1(n5396), .B2(n8893), .A(n5388), .ZN(n5387) );
  NAND2_X1 U5744 ( .A1(n5389), .A2(n5394), .ZN(n5388) );
  NAND2_X1 U5745 ( .A1(n8724), .A2(n8726), .ZN(n5394) );
  AND2_X1 U5746 ( .A1(n8722), .A2(n8815), .ZN(n5395) );
  INV_X1 U5747 ( .A(n5393), .ZN(n5389) );
  AND2_X1 U5748 ( .A1(n5383), .A2(n5382), .ZN(n5391) );
  NAND2_X1 U5749 ( .A1(n5274), .A2(n9222), .ZN(n5273) );
  INV_X1 U5750 ( .A(n5364), .ZN(n5363) );
  OAI21_X1 U5751 ( .B1(n8745), .B2(n8744), .A(n5368), .ZN(n5364) );
  INV_X1 U5752 ( .A(n10389), .ZN(n5366) );
  OAI211_X1 U5753 ( .C1(n5271), .C2(n5270), .A(n5269), .B(n9238), .ZN(n9241)
         );
  AOI21_X1 U5754 ( .B1(n5358), .B2(n5360), .A(n5357), .ZN(n5356) );
  AOI21_X1 U5755 ( .B1(n8755), .B2(n8782), .A(n10358), .ZN(n5380) );
  OAI21_X1 U5756 ( .B1(n8746), .B2(n5360), .A(n5358), .ZN(n8754) );
  INV_X1 U5757 ( .A(SI_17_), .ZN(n9478) );
  INV_X1 U5758 ( .A(SI_16_), .ZN(n9652) );
  INV_X1 U5759 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9583) );
  INV_X1 U5760 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9805) );
  INV_X1 U5761 ( .A(SI_11_), .ZN(n9694) );
  NOR2_X1 U5762 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .ZN(
        n5740) );
  INV_X1 U5763 ( .A(SI_21_), .ZN(n9467) );
  INV_X1 U5764 ( .A(SI_19_), .ZN(n9474) );
  INV_X1 U5765 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6262) );
  INV_X1 U5766 ( .A(n6041), .ZN(n5655) );
  OAI21_X1 U5767 ( .B1(n7159), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n5195), .ZN(
        n5875) );
  NAND2_X1 U5768 ( .A1(n7159), .A2(n9810), .ZN(n5195) );
  AND2_X1 U5769 ( .A1(n5666), .A2(n5180), .ZN(n5664) );
  AOI21_X1 U5770 ( .B1(n9263), .B2(n5294), .A(n5292), .ZN(n5291) );
  NAND2_X1 U5771 ( .A1(n5293), .A2(n9267), .ZN(n5292) );
  NAND2_X1 U5772 ( .A1(n5294), .A2(n5296), .ZN(n5293) );
  NAND2_X1 U5773 ( .A1(n5634), .A2(n5633), .ZN(n5632) );
  INV_X1 U5774 ( .A(n9304), .ZN(n5634) );
  AND2_X1 U5775 ( .A1(n5637), .A2(n5127), .ZN(n5633) );
  AOI21_X1 U5776 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n10903), .A(n10894), .ZN(
        n8000) );
  NAND2_X1 U5777 ( .A1(n8195), .A2(n8196), .ZN(n8198) );
  INV_X1 U5778 ( .A(n8584), .ZN(n5469) );
  OR2_X1 U5779 ( .A1(n9906), .A2(n8971), .ZN(n9246) );
  INV_X1 U5780 ( .A(n9226), .ZN(n5483) );
  NOR2_X1 U5781 ( .A1(n5483), .A2(n5276), .ZN(n5480) );
  INV_X1 U5782 ( .A(n5441), .ZN(n5440) );
  OAI21_X1 U5783 ( .B1(n6664), .B2(n5442), .A(n9944), .ZN(n5441) );
  INV_X1 U5784 ( .A(n6665), .ZN(n5442) );
  NOR2_X1 U5785 ( .A1(n6617), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U5786 ( .A1(n8042), .A2(n9281), .ZN(n5450) );
  OR2_X1 U5787 ( .A1(n5418), .A2(n5416), .ZN(n5410) );
  NOR2_X1 U5788 ( .A1(n5417), .A2(n5416), .ZN(n5414) );
  NOR2_X1 U5789 ( .A1(n5150), .A2(n5448), .ZN(n5447) );
  OR2_X1 U5790 ( .A1(n6822), .A2(n6836), .ZN(n7145) );
  AND2_X1 U5791 ( .A1(n6364), .A2(n6802), .ZN(n5704) );
  INV_X1 U5792 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6842) );
  INV_X1 U5793 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6359) );
  INV_X1 U5794 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U5795 ( .A1(n6427), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6454) );
  INV_X1 U5796 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5625) );
  NAND2_X1 U5797 ( .A1(n5740), .A2(n9421), .ZN(n5630) );
  INV_X1 U5798 ( .A(n7055), .ZN(n5584) );
  OR2_X1 U5799 ( .A1(n5587), .A2(n5582), .ZN(n5581) );
  INV_X1 U5800 ( .A(n10143), .ZN(n5582) );
  AND2_X1 U5801 ( .A1(n5566), .A2(n6942), .ZN(n5565) );
  NAND2_X1 U5802 ( .A1(n5552), .A2(n5555), .ZN(n6997) );
  INV_X1 U5803 ( .A(n5556), .ZN(n5555) );
  OAI21_X1 U5804 ( .B1(n6987), .B2(n5559), .A(n5557), .ZN(n5556) );
  AOI21_X1 U5805 ( .B1(n5377), .B2(n8771), .A(n8770), .ZN(n8776) );
  OR2_X1 U5806 ( .A1(n10538), .A2(n8765), .ZN(n8772) );
  NOR2_X1 U5807 ( .A1(n6175), .A2(n10125), .ZN(n6190) );
  OR2_X1 U5808 ( .A1(n10558), .A2(n10091), .ZN(n8825) );
  OR2_X1 U5809 ( .A1(n10405), .A2(n10147), .ZN(n8750) );
  OR2_X1 U5810 ( .A1(n10568), .A2(n10082), .ZN(n10410) );
  INV_X1 U5811 ( .A(n5533), .ZN(n5528) );
  NAND2_X1 U5812 ( .A1(n8690), .A2(n5154), .ZN(n8877) );
  NOR2_X1 U5813 ( .A1(n5904), .A2(n7247), .ZN(n5917) );
  INV_X1 U5814 ( .A(n5352), .ZN(n5351) );
  AND2_X1 U5815 ( .A1(n10652), .A2(n5131), .ZN(n5332) );
  AND2_X1 U5816 ( .A1(n8676), .A2(n8790), .ZN(n8674) );
  OAI21_X1 U5817 ( .B1(n6246), .B2(n5615), .A(n5613), .ZN(n8638) );
  AOI21_X1 U5818 ( .B1(n6738), .B2(n5614), .A(n5190), .ZN(n5613) );
  INV_X1 U5819 ( .A(n6738), .ZN(n5615) );
  XNOR2_X1 U5820 ( .A(n8638), .B(n8637), .ZN(n8636) );
  INV_X1 U5821 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5725) );
  INV_X1 U5822 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5724) );
  INV_X1 U5823 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5723) );
  AND2_X1 U5824 ( .A1(n6245), .A2(n6226), .ZN(n6227) );
  NOR2_X1 U5825 ( .A1(n6201), .A2(n5642), .ZN(n5641) );
  NAND2_X1 U5826 ( .A1(n6117), .A2(n6116), .ZN(n5644) );
  NOR2_X1 U5827 ( .A1(n6024), .A2(n5657), .ZN(n5656) );
  INV_X1 U5828 ( .A(n6007), .ZN(n5657) );
  NAND2_X1 U5829 ( .A1(n5300), .A2(n5149), .ZN(n6008) );
  INV_X1 U5830 ( .A(n6005), .ZN(n5299) );
  INV_X1 U5831 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5721) );
  INV_X1 U5832 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U5833 ( .A1(n5617), .A2(n5616), .ZN(n5947) );
  AOI21_X1 U5834 ( .B1(n5130), .B2(n5622), .A(n5171), .ZN(n5616) );
  OR2_X1 U5835 ( .A1(n5898), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5913) );
  NOR2_X1 U5836 ( .A1(n5268), .A2(n5870), .ZN(n5264) );
  OR2_X1 U5837 ( .A1(n5314), .A2(n5268), .ZN(n5262) );
  NAND2_X1 U5838 ( .A1(n5244), .A2(n5856), .ZN(n5872) );
  NAND2_X1 U5839 ( .A1(n5854), .A2(n5853), .ZN(n5244) );
  INV_X1 U5840 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U5841 ( .A1(n6514), .A2(n9744), .ZN(n6525) );
  AND2_X1 U5842 ( .A1(n5681), .A2(n9001), .ZN(n5680) );
  OR2_X1 U5843 ( .A1(n9078), .A2(n5682), .ZN(n5681) );
  INV_X1 U5844 ( .A(n8975), .ZN(n5682) );
  NAND2_X1 U5845 ( .A1(n9381), .A2(n6598), .ZN(n6617) );
  NAND2_X1 U5846 ( .A1(n7547), .A2(n7554), .ZN(n7605) );
  XNOR2_X1 U5847 ( .A(n10963), .B(n7550), .ZN(n7608) );
  NAND2_X1 U5848 ( .A1(n7733), .A2(n7890), .ZN(n5673) );
  INV_X1 U5849 ( .A(n9064), .ZN(n5660) );
  NAND2_X1 U5850 ( .A1(n5661), .A2(n5234), .ZN(n5232) );
  INV_X1 U5851 ( .A(n5664), .ZN(n5663) );
  AOI21_X1 U5852 ( .B1(n5664), .B2(n5669), .A(n5662), .ZN(n5661) );
  INV_X1 U5853 ( .A(n9023), .ZN(n5662) );
  XNOR2_X1 U5854 ( .A(n7550), .B(n8073), .ZN(n7348) );
  INV_X1 U5855 ( .A(n7608), .ZN(n7547) );
  NOR2_X1 U5856 ( .A1(n8553), .A2(n8554), .ZN(n8552) );
  INV_X1 U5857 ( .A(n9320), .ZN(n8950) );
  OR2_X1 U5858 ( .A1(n9244), .A2(n7344), .ZN(n7139) );
  OR2_X1 U5859 ( .A1(n6701), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6422) );
  AND2_X1 U5860 ( .A1(n7402), .A2(n7406), .ZN(n10872) );
  INV_X1 U5861 ( .A(n5461), .ZN(n7537) );
  OR2_X1 U5862 ( .A1(n7536), .A2(n7538), .ZN(n5461) );
  NOR2_X1 U5863 ( .A1(n7397), .A2(n7530), .ZN(n7399) );
  INV_X1 U5864 ( .A(n5590), .ZN(n7396) );
  AOI21_X1 U5865 ( .B1(n7521), .B2(n7520), .A(n7519), .ZN(n7522) );
  NOR2_X1 U5866 ( .A1(n7694), .A2(n7695), .ZN(n10896) );
  AOI21_X1 U5867 ( .B1(n7684), .B2(n7683), .A(n7682), .ZN(n10889) );
  NOR2_X1 U5868 ( .A1(n10891), .A2(n7680), .ZN(n7985) );
  OAI21_X1 U5869 ( .B1(n8098), .B2(n5603), .A(n5602), .ZN(n8426) );
  NAND2_X1 U5870 ( .A1(n5604), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5603) );
  INV_X1 U5871 ( .A(n8191), .ZN(n5604) );
  NOR2_X1 U5872 ( .A1(n8098), .A2(n8100), .ZN(n8189) );
  INV_X1 U5873 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U5874 ( .A1(n5607), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U5875 ( .A1(n8588), .A2(n5607), .ZN(n5605) );
  INV_X1 U5876 ( .A(n9342), .ZN(n5607) );
  NOR2_X1 U5877 ( .A1(n8504), .A2(n8506), .ZN(n8587) );
  NAND2_X1 U5878 ( .A1(n9347), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5470) );
  OAI21_X1 U5879 ( .B1(n9395), .B2(n5609), .A(n5608), .ZN(n9408) );
  NAND2_X1 U5880 ( .A1(n5612), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5609) );
  INV_X1 U5881 ( .A(n8596), .ZN(n5612) );
  NAND2_X1 U5882 ( .A1(n5469), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5468) );
  INV_X1 U5883 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n9421) );
  AND2_X1 U5884 ( .A1(n9240), .A2(n9239), .ZN(n9913) );
  INV_X1 U5885 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9540) );
  AND2_X1 U5886 ( .A1(n6699), .A2(n9540), .ZN(n6712) );
  OR2_X1 U5887 ( .A1(n6678), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U5888 ( .A1(n6669), .A2(n9027), .ZN(n6678) );
  AND2_X1 U5889 ( .A1(n6658), .A2(n9535), .ZN(n6669) );
  AND2_X1 U5890 ( .A1(n6646), .A2(n9518), .ZN(n6658) );
  INV_X1 U5891 ( .A(n6616), .ZN(n6631) );
  NOR2_X1 U5892 ( .A1(n6586), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U5893 ( .A1(n9348), .A2(n6571), .ZN(n6586) );
  INV_X1 U5894 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9348) );
  AND4_X1 U5895 ( .A1(n6590), .A2(n6589), .A3(n6588), .A4(n6587), .ZN(n8467)
         );
  NAND2_X1 U5896 ( .A1(n8329), .A2(n8335), .ZN(n5437) );
  AND2_X1 U5897 ( .A1(n9189), .A2(n8398), .ZN(n9196) );
  NAND2_X1 U5898 ( .A1(n5174), .A2(n9195), .ZN(n5488) );
  NAND2_X1 U5899 ( .A1(n6374), .A2(n6548), .ZN(n6561) );
  INV_X1 U5900 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6374) );
  AND2_X1 U5901 ( .A1(n9177), .A2(n9166), .ZN(n9283) );
  NAND2_X1 U5902 ( .A1(n5450), .A2(n6520), .ZN(n8156) );
  INV_X1 U5903 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7817) );
  AND2_X1 U5904 ( .A1(n6493), .A2(n7817), .ZN(n6514) );
  OR2_X1 U5905 ( .A1(n6460), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6478) );
  NOR2_X1 U5906 ( .A1(n6478), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6493) );
  INV_X1 U5907 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7642) );
  NOR2_X1 U5908 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6446) );
  NOR2_X1 U5909 ( .A1(n5120), .A2(n5631), .ZN(n5446) );
  NOR2_X1 U5910 ( .A1(n7168), .A2(n7159), .ZN(n5445) );
  OR2_X1 U5911 ( .A1(n9244), .A2(n6799), .ZN(n7759) );
  OR2_X1 U5912 ( .A1(n9435), .A2(n9434), .ZN(n9990) );
  NAND2_X1 U5913 ( .A1(n6644), .A2(n6643), .ZN(n10028) );
  NAND2_X1 U5914 ( .A1(n7711), .A2(n9156), .ZN(n7902) );
  OR2_X1 U5915 ( .A1(n8157), .A2(n11008), .ZN(n11132) );
  AND2_X1 U5916 ( .A1(n6817), .A2(n6816), .ZN(n6838) );
  XNOR2_X1 U5917 ( .A(n6841), .B(n6842), .ZN(n8266) );
  AOI21_X1 U5918 ( .B1(n5686), .B2(n6521), .A(n6521), .ZN(n5684) );
  AND2_X1 U5919 ( .A1(n6500), .A2(n6489), .ZN(n8001) );
  NAND2_X1 U5920 ( .A1(n10152), .A2(n10155), .ZN(n5549) );
  INV_X1 U5921 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U5922 ( .A1(n6013), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6036) );
  INV_X1 U5923 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8022) );
  INV_X1 U5924 ( .A(n5206), .ZN(n6049) );
  XNOR2_X1 U5925 ( .A(n6899), .B(n7089), .ZN(n6904) );
  INV_X1 U5926 ( .A(n6091), .ZN(n6089) );
  OR2_X1 U5927 ( .A1(n5957), .A2(n5956), .ZN(n5976) );
  INV_X1 U5928 ( .A(n5205), .ZN(n5996) );
  OR2_X1 U5929 ( .A1(n7461), .A2(n7059), .ZN(n6881) );
  NAND2_X1 U5930 ( .A1(n7029), .A2(n7028), .ZN(n10153) );
  INV_X1 U5931 ( .A(n7026), .ZN(n7029) );
  INV_X1 U5932 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5844) );
  NOR2_X1 U5933 ( .A1(n5845), .A2(n5844), .ZN(n5861) );
  OR2_X1 U5934 ( .A1(n8653), .A2(n7216), .ZN(n5790) );
  NAND2_X1 U5935 ( .A1(n6258), .A2(n5401), .ZN(n5400) );
  INV_X1 U5936 ( .A(n5404), .ZN(n5401) );
  NAND2_X1 U5937 ( .A1(n5204), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8935) );
  AND2_X1 U5938 ( .A1(n6250), .A2(n6234), .ZN(n10345) );
  OR2_X1 U5939 ( .A1(n10359), .A2(n10358), .ZN(n10361) );
  NOR2_X1 U5940 ( .A1(n10403), .A2(n10558), .ZN(n10394) );
  AND2_X1 U5941 ( .A1(n8829), .A2(n8757), .ZN(n10379) );
  NAND2_X1 U5942 ( .A1(n10402), .A2(n6315), .ZN(n10403) );
  NAND2_X1 U5943 ( .A1(n10422), .A2(n6145), .ZN(n10401) );
  NAND2_X1 U5944 ( .A1(n5207), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6138) );
  INV_X1 U5945 ( .A(n5207), .ZN(n6122) );
  AOI21_X1 U5946 ( .B1(n5511), .B2(n5517), .A(n5165), .ZN(n5510) );
  NAND2_X1 U5947 ( .A1(n5247), .A2(n5246), .ZN(n10472) );
  NOR2_X1 U5948 ( .A1(n5133), .A2(n8728), .ZN(n5246) );
  NAND2_X1 U5949 ( .A1(n8380), .A2(n5248), .ZN(n5247) );
  NAND2_X1 U5950 ( .A1(n5398), .A2(n5397), .ZN(n10488) );
  NAND2_X1 U5951 ( .A1(n8363), .A2(n5334), .ZN(n10516) );
  NAND2_X1 U5952 ( .A1(n8363), .A2(n10606), .ZN(n8376) );
  NAND2_X1 U5953 ( .A1(n5238), .A2(n5236), .ZN(n8351) );
  AND2_X1 U5954 ( .A1(n5176), .A2(n5237), .ZN(n5236) );
  NAND2_X1 U5955 ( .A1(n7834), .A2(n5239), .ZN(n5238) );
  OAI21_X1 U5956 ( .B1(n7834), .B2(n5240), .A(n5239), .ZN(n8138) );
  NAND2_X1 U5957 ( .A1(n7834), .A2(n8881), .ZN(n7950) );
  AOI21_X1 U5958 ( .B1(n8794), .B2(n5521), .A(n5163), .ZN(n5520) );
  INV_X1 U5959 ( .A(n5911), .ZN(n5521) );
  OAI21_X1 U5960 ( .B1(n6288), .B2(n5370), .A(n5372), .ZN(n5369) );
  INV_X1 U5961 ( .A(n6288), .ZN(n5374) );
  INV_X1 U5962 ( .A(n10209), .ZN(n7751) );
  NAND2_X1 U5963 ( .A1(n5373), .A2(n6288), .ZN(n7590) );
  NAND2_X1 U5964 ( .A1(n8870), .A2(n5375), .ZN(n5373) );
  NAND2_X1 U5965 ( .A1(n7335), .A2(n7448), .ZN(n7468) );
  OR2_X1 U5966 ( .A1(n7193), .A2(n5123), .ZN(n8353) );
  OR2_X1 U5967 ( .A1(n7193), .A2(n7248), .ZN(n8944) );
  AOI21_X1 U5968 ( .B1(n7182), .B2(n7191), .A(n7189), .ZN(n7098) );
  NAND2_X1 U5969 ( .A1(n6209), .A2(n6208), .ZN(n10353) );
  OAI21_X1 U5970 ( .B1(n7745), .B2(n5503), .A(n5128), .ZN(n7794) );
  NAND2_X1 U5971 ( .A1(n7744), .A2(n5869), .ZN(n7795) );
  OR2_X1 U5972 ( .A1(n8815), .A2(n8856), .ZN(n10616) );
  NOR2_X1 U5973 ( .A1(n7446), .A2(n5188), .ZN(n7579) );
  INV_X1 U5974 ( .A(n5542), .ZN(n7447) );
  OR2_X1 U5975 ( .A1(n7112), .A2(n8919), .ZN(n11109) );
  NOR2_X1 U5976 ( .A1(n6350), .A2(n7564), .ZN(n6354) );
  INV_X1 U5977 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5733) );
  XNOR2_X1 U5978 ( .A(n8636), .B(SI_29_), .ZN(n8762) );
  XNOR2_X1 U5979 ( .A(n6739), .B(n6738), .ZN(n8532) );
  NAND2_X1 U5980 ( .A1(n6246), .A2(n6245), .ZN(n6739) );
  NOR2_X1 U5981 ( .A1(n5746), .A2(n5803), .ZN(n5354) );
  XNOR2_X1 U5982 ( .A(n6223), .B(n6222), .ZN(n8476) );
  NAND2_X1 U5983 ( .A1(n5640), .A2(n6204), .ZN(n6223) );
  INV_X1 U5984 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U5985 ( .A1(n6319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6320) );
  XNOR2_X1 U5986 ( .A(n6347), .B(n6346), .ZN(n7195) );
  INV_X1 U5987 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6346) );
  XNOR2_X1 U5988 ( .A(n6085), .B(n6264), .ZN(n6275) );
  NAND2_X1 U5989 ( .A1(n5300), .A2(n5301), .ZN(n6006) );
  CLKBUF_X1 U5990 ( .A(n5971), .Z(n5972) );
  NAND2_X1 U5991 ( .A1(n5618), .A2(n5619), .ZN(n5925) );
  OR2_X1 U5992 ( .A1(n5894), .A2(n5622), .ZN(n5618) );
  NAND2_X1 U5993 ( .A1(n5316), .A2(n5314), .ZN(n5894) );
  NAND2_X1 U5994 ( .A1(n5267), .A2(n5265), .ZN(n7197) );
  NAND2_X1 U5995 ( .A1(n5316), .A2(n5266), .ZN(n5265) );
  AND3_X1 U5996 ( .A1(n5263), .A2(n5262), .A3(n5161), .ZN(n5267) );
  AND2_X1 U5997 ( .A1(n5314), .A2(n5713), .ZN(n5266) );
  OR2_X1 U5998 ( .A1(n5825), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5951) );
  AOI21_X1 U5999 ( .B1(n5801), .B2(n5800), .A(n5140), .ZN(n5819) );
  XNOR2_X1 U6000 ( .A(n5770), .B(n5756), .ZN(n5768) );
  AND2_X1 U6001 ( .A1(n5676), .A2(n7730), .ZN(n7734) );
  NAND2_X1 U6002 ( .A1(n5215), .A2(n5217), .ZN(n8470) );
  NAND2_X1 U6003 ( .A1(n5216), .A2(n5125), .ZN(n5215) );
  NAND2_X1 U6004 ( .A1(n7816), .A2(n7815), .ZN(n7891) );
  NAND2_X1 U6005 ( .A1(n5665), .A2(n5666), .ZN(n9025) );
  NAND2_X1 U6006 ( .A1(n9015), .A2(n5668), .ZN(n5665) );
  OR2_X1 U6007 ( .A1(n9312), .A2(n7368), .ZN(n9019) );
  NAND2_X1 U6008 ( .A1(n9008), .A2(n8966), .ZN(n9043) );
  NAND2_X1 U6009 ( .A1(n6697), .A2(n6696), .ZN(n10008) );
  OAI21_X1 U6010 ( .B1(n7722), .B2(n5210), .A(n5671), .ZN(n7893) );
  NAND2_X1 U6011 ( .A1(n5674), .A2(n5714), .ZN(n5210) );
  OAI21_X1 U6012 ( .B1(n5673), .B2(n7731), .A(n5674), .ZN(n5671) );
  AOI21_X1 U6013 ( .B1(n5675), .B2(n7890), .A(n7889), .ZN(n5674) );
  NAND2_X1 U6014 ( .A1(n7893), .A2(n7892), .ZN(n8131) );
  NAND2_X1 U6015 ( .A1(n9015), .A2(n8956), .ZN(n9053) );
  OAI21_X1 U6016 ( .B1(n9015), .B2(n5663), .A(n5661), .ZN(n9065) );
  INV_X1 U6017 ( .A(n5689), .ZN(n5688) );
  OAI21_X1 U6018 ( .B1(n5694), .B2(n5691), .A(n5690), .ZN(n5689) );
  INV_X1 U6019 ( .A(n5693), .ZN(n8566) );
  OAI21_X1 U6020 ( .B1(n8552), .B2(n5695), .A(n5189), .ZN(n5693) );
  AND3_X1 U6021 ( .A1(n6472), .A2(n6471), .A3(n6470), .ZN(n7625) );
  NAND2_X1 U6022 ( .A1(n5224), .A2(n5227), .ZN(n9075) );
  NAND2_X1 U6023 ( .A1(n9041), .A2(n5229), .ZN(n5224) );
  NAND2_X1 U6024 ( .A1(n5223), .A2(n5225), .ZN(n9077) );
  AND2_X1 U6025 ( .A1(n5226), .A2(n9078), .ZN(n5225) );
  NAND2_X1 U6026 ( .A1(n5227), .A2(n5230), .ZN(n5226) );
  INV_X1 U6027 ( .A(n9061), .ZN(n9076) );
  AOI21_X1 U6028 ( .B1(n5213), .B2(n5219), .A(n5126), .ZN(n5212) );
  NAND2_X1 U6029 ( .A1(n7364), .A2(n10950), .ZN(n9059) );
  OAI21_X1 U6030 ( .B1(n6813), .B2(n6367), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6383) );
  OR2_X1 U6031 ( .A1(n7139), .A2(n7361), .ZN(n9312) );
  XNOR2_X1 U6032 ( .A(n6758), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9313) );
  INV_X1 U6033 ( .A(n9068), .ZN(n9963) );
  INV_X1 U6034 ( .A(n8954), .ZN(n9962) );
  INV_X1 U6035 ( .A(P2_U3893), .ZN(n9336) );
  OAI21_X1 U6036 ( .B1(n7416), .B2(n7315), .A(n7403), .ZN(n7316) );
  NOR2_X1 U6037 ( .A1(n10882), .A2(n10881), .ZN(n10880) );
  XNOR2_X1 U6038 ( .A(n5590), .B(n7546), .ZN(n7531) );
  INV_X1 U6039 ( .A(n7409), .ZN(n5460) );
  XNOR2_X1 U6040 ( .A(n7985), .B(n8001), .ZN(n7681) );
  NOR2_X1 U6041 ( .A1(n7681), .A2(n6476), .ZN(n7986) );
  NAND2_X1 U6042 ( .A1(n5594), .A2(n5595), .ZN(n10913) );
  NAND2_X1 U6043 ( .A1(n6533), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6544) );
  INV_X1 U6044 ( .A(n6365), .ZN(n6533) );
  INV_X1 U6045 ( .A(n5600), .ZN(n9361) );
  OAI21_X1 U6046 ( .B1(n9359), .B2(n5598), .A(n5597), .ZN(n9374) );
  NAND2_X1 U6047 ( .A1(n5601), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U6048 ( .A1(n8591), .A2(n5601), .ZN(n5597) );
  INV_X1 U6049 ( .A(n9375), .ZN(n5601) );
  INV_X1 U6050 ( .A(n8591), .ZN(n5599) );
  NOR2_X1 U6051 ( .A1(n9408), .A2(n5610), .ZN(n9410) );
  NOR2_X1 U6052 ( .A1(n8595), .A2(n5611), .ZN(n5610) );
  AND2_X1 U6053 ( .A1(n10865), .A2(n9412), .ZN(n9429) );
  OAI21_X1 U6054 ( .B1(n9079), .B2(n8524), .A(n9442), .ZN(n9443) );
  NAND2_X1 U6055 ( .A1(n9891), .A2(n6775), .ZN(n9882) );
  AND2_X1 U6056 ( .A1(n9877), .A2(n9876), .ZN(n9998) );
  NAND2_X1 U6057 ( .A1(n5422), .A2(n5427), .ZN(n9873) );
  INV_X1 U6058 ( .A(n5201), .ZN(n5200) );
  XNOR2_X1 U6059 ( .A(n9888), .B(n9887), .ZN(n5202) );
  AOI22_X1 U6060 ( .A1(n5433), .A2(n10944), .B1(n9961), .B2(n9914), .ZN(n5201)
         );
  NAND2_X1 U6061 ( .A1(n6685), .A2(n6684), .ZN(n9922) );
  NAND2_X1 U6062 ( .A1(n9951), .A2(n9226), .ZN(n9940) );
  NAND2_X1 U6063 ( .A1(n6676), .A2(n6675), .ZN(n10016) );
  NAND2_X1 U6064 ( .A1(n6667), .A2(n6666), .ZN(n10020) );
  NAND2_X1 U6065 ( .A1(n9959), .A2(n6665), .ZN(n9945) );
  AND2_X1 U6066 ( .A1(n6656), .A2(n6655), .ZN(n9972) );
  AND2_X1 U6067 ( .A1(n5493), .A2(n9213), .ZN(n8528) );
  NAND2_X1 U6068 ( .A1(n6629), .A2(n6628), .ZN(n10032) );
  NAND2_X1 U6069 ( .A1(n6770), .A2(n9205), .ZN(n8485) );
  NAND2_X1 U6070 ( .A1(n6614), .A2(n6613), .ZN(n11150) );
  NAND2_X1 U6071 ( .A1(n6597), .A2(n6596), .ZN(n11144) );
  NAND2_X1 U6072 ( .A1(n6585), .A2(n6584), .ZN(n11138) );
  NAND2_X1 U6073 ( .A1(n5490), .A2(n8286), .ZN(n8336) );
  NAND2_X1 U6074 ( .A1(n6766), .A2(n5142), .ZN(n5490) );
  NAND2_X1 U6075 ( .A1(n6766), .A2(n9180), .ZN(n8217) );
  NAND2_X1 U6076 ( .A1(n6547), .A2(n6546), .ZN(n11105) );
  NAND2_X1 U6077 ( .A1(n6764), .A2(n9165), .ZN(n8041) );
  NAND2_X1 U6078 ( .A1(n6503), .A2(n6504), .ZN(n7970) );
  OAI21_X1 U6079 ( .B1(n6433), .B2(n5413), .A(n5412), .ZN(n7714) );
  INV_X1 U6080 ( .A(n5418), .ZN(n5413) );
  NAND2_X1 U6081 ( .A1(n5415), .A2(n6443), .ZN(n8079) );
  NAND2_X1 U6082 ( .A1(n6433), .A2(n6432), .ZN(n7878) );
  INV_X1 U6083 ( .A(n9954), .ZN(n9987) );
  OR2_X1 U6084 ( .A1(n11127), .A2(n7766), .ZN(n10974) );
  INV_X1 U6085 ( .A(n10963), .ZN(n10977) );
  OR2_X1 U6086 ( .A1(n10941), .A2(n10974), .ZN(n9984) );
  NAND2_X1 U6087 ( .A1(n11048), .A2(n11036), .ZN(n9954) );
  NAND2_X1 U6088 ( .A1(n7363), .A2(n7766), .ZN(n10950) );
  INV_X1 U6089 ( .A(n5475), .ZN(n5477) );
  OR2_X1 U6090 ( .A1(n10007), .A2(n10006), .ZN(n10042) );
  INV_X2 U6091 ( .A(n11154), .ZN(n11157) );
  AND2_X1 U6092 ( .A1(n7365), .A2(n7259), .ZN(n7192) );
  NAND2_X1 U6093 ( .A1(n5173), .A2(n5198), .ZN(n10052) );
  AND2_X1 U6094 ( .A1(n6365), .A2(n5199), .ZN(n5198) );
  INV_X1 U6095 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U6096 ( .A1(n6808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6810) );
  INV_X1 U6097 ( .A(n9313), .ZN(n8237) );
  INV_X1 U6098 ( .A(n7342), .ZN(n9120) );
  INV_X1 U6099 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U6100 ( .A1(n5685), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6757) );
  INV_X1 U6101 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7912) );
  XNOR2_X1 U6102 ( .A(n6754), .B(n6753), .ZN(n9409) );
  INV_X1 U6103 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7631) );
  INV_X1 U6104 ( .A(n8613), .ZN(n9380) );
  INV_X1 U6105 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7311) );
  INV_X1 U6106 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7255) );
  XNOR2_X1 U6107 ( .A(n6502), .B(n6501), .ZN(n8103) );
  NAND2_X1 U6108 ( .A1(n8298), .A2(n6987), .ZN(n8386) );
  NAND2_X1 U6109 ( .A1(n5554), .A2(n6992), .ZN(n8387) );
  NAND2_X1 U6110 ( .A1(n8298), .A2(n6990), .ZN(n5554) );
  AND2_X1 U6111 ( .A1(n5588), .A2(n5586), .ZN(n10058) );
  NAND2_X1 U6112 ( .A1(n10140), .A2(n10143), .ZN(n5586) );
  OR2_X1 U6113 ( .A1(n5578), .A2(n6958), .ZN(n8168) );
  AND2_X1 U6114 ( .A1(n7936), .A2(n6953), .ZN(n5578) );
  CLKBUF_X1 U6115 ( .A(n7486), .Z(n7487) );
  NAND2_X1 U6116 ( .A1(n5549), .A2(n10153), .ZN(n10068) );
  NAND2_X1 U6117 ( .A1(n6088), .A2(n6087), .ZN(n10479) );
  CLKBUF_X1 U6118 ( .A(n7431), .Z(n7432) );
  CLKBUF_X1 U6119 ( .A(n10078), .Z(n10079) );
  INV_X1 U6120 ( .A(n7956), .ZN(n11110) );
  INV_X1 U6121 ( .A(n5572), .ZN(n10176) );
  NAND2_X1 U6122 ( .A1(n6189), .A2(n6188), .ZN(n10373) );
  NAND2_X1 U6123 ( .A1(n10096), .A2(n7011), .ZN(n10108) );
  NAND2_X1 U6124 ( .A1(n8297), .A2(n6980), .ZN(n8298) );
  INV_X1 U6125 ( .A(n5576), .ZN(n5574) );
  OAI22_X1 U6126 ( .A1(n5576), .A2(n6953), .B1(n5577), .B2(n6958), .ZN(n5573)
         );
  INV_X1 U6127 ( .A(n7916), .ZN(n11095) );
  INV_X1 U6128 ( .A(n11091), .ZN(n10194) );
  INV_X1 U6129 ( .A(n11097), .ZN(n10199) );
  AOI21_X1 U6130 ( .B1(n10197), .B2(n7072), .A(n6996), .ZN(n10186) );
  NAND2_X1 U6131 ( .A1(n8857), .A2(n5712), .ZN(n8858) );
  INV_X1 U6132 ( .A(n8847), .ZN(n8857) );
  NAND2_X1 U6133 ( .A1(n6218), .A2(n6217), .ZN(n10381) );
  NAND2_X1 U6134 ( .A1(n6182), .A2(n6181), .ZN(n10416) );
  INV_X1 U6135 ( .A(n5541), .ZN(n5540) );
  INV_X1 U6136 ( .A(n5551), .ZN(n5550) );
  NAND2_X1 U6137 ( .A1(n8779), .A2(n8778), .ZN(n10320) );
  AND2_X1 U6138 ( .A1(n5526), .A2(n5524), .ZN(n8934) );
  NAND2_X1 U6139 ( .A1(n5526), .A2(n6244), .ZN(n6260) );
  NAND2_X1 U6140 ( .A1(n5307), .A2(n10512), .ZN(n6313) );
  AND2_X1 U6141 ( .A1(n8831), .A2(n6296), .ZN(n5249) );
  NAND2_X1 U6142 ( .A1(n10462), .A2(n8740), .ZN(n10439) );
  NAND2_X1 U6143 ( .A1(n5513), .A2(n5515), .ZN(n10457) );
  NAND2_X1 U6144 ( .A1(n5514), .A2(n8733), .ZN(n5513) );
  INV_X1 U6145 ( .A(n6074), .ZN(n5514) );
  NAND2_X1 U6146 ( .A1(n6074), .A2(n6073), .ZN(n10470) );
  OAI21_X1 U6147 ( .B1(n8320), .B2(n5508), .A(n5506), .ZN(n10515) );
  AND2_X1 U6148 ( .A1(n5398), .A2(n8726), .ZN(n10506) );
  NAND2_X1 U6149 ( .A1(n8374), .A2(n8803), .ZN(n8373) );
  NAND2_X1 U6150 ( .A1(n8320), .A2(n6022), .ZN(n8374) );
  NAND2_X1 U6151 ( .A1(n5532), .A2(n5530), .ZN(n8358) );
  NAND2_X1 U6152 ( .A1(n5532), .A2(n5535), .ZN(n8356) );
  OAI21_X1 U6153 ( .B1(n7949), .B2(n5965), .A(n5964), .ZN(n8145) );
  NAND2_X1 U6154 ( .A1(n7826), .A2(n8794), .ZN(n7825) );
  NAND2_X1 U6155 ( .A1(n7846), .A2(n5911), .ZN(n7826) );
  NAND2_X1 U6156 ( .A1(n7849), .A2(n11065), .ZN(n7828) );
  OR2_X1 U6157 ( .A1(n10466), .A2(n7569), .ZN(n10525) );
  AND2_X1 U6158 ( .A1(n8368), .A2(n7587), .ZN(n10504) );
  OR2_X1 U6159 ( .A1(n10466), .A2(n8923), .ZN(n11021) );
  INV_X1 U6160 ( .A(n10525), .ZN(n11018) );
  INV_X1 U6161 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6162 ( .A1(n5336), .A2(n5196), .ZN(n5498) );
  INV_X1 U6163 ( .A(n5337), .ZN(n5336) );
  NOR2_X1 U6164 ( .A1(n5197), .A2(n10537), .ZN(n5196) );
  INV_X1 U6165 ( .A(n10353), .ZN(n10632) );
  INV_X1 U6166 ( .A(n10373), .ZN(n10636) );
  INV_X1 U6167 ( .A(n10405), .ZN(n6315) );
  NAND2_X1 U6168 ( .A1(n7184), .A2(n7183), .ZN(n10671) );
  XNOR2_X1 U6169 ( .A(n8659), .B(n8658), .ZN(n10664) );
  OAI21_X1 U6170 ( .B1(n8656), .B2(n8655), .A(n8654), .ZN(n8659) );
  INV_X1 U6171 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9569) );
  INV_X1 U6172 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9782) );
  NAND2_X1 U6173 ( .A1(n6169), .A2(n6156), .ZN(n8265) );
  NAND2_X1 U6174 ( .A1(n5650), .A2(n5648), .ZN(n6169) );
  NAND2_X1 U6175 ( .A1(n5650), .A2(n6150), .ZN(n6155) );
  NAND2_X1 U6176 ( .A1(n6268), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6269) );
  INV_X1 U6177 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9573) );
  INV_X1 U6178 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9793) );
  INV_X1 U6179 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9797) );
  INV_X1 U6180 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9810) );
  CLKBUF_X1 U6181 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n10752) );
  INV_X1 U6182 ( .A(n5473), .ZN(n9340) );
  NAND2_X1 U6183 ( .A1(n5475), .A2(n11153), .ZN(n5474) );
  OAI21_X1 U6184 ( .B1(n7128), .B2(n7099), .A(n11097), .ZN(n5203) );
  NAND2_X1 U6185 ( .A1(n7128), .A2(n5569), .ZN(n7136) );
  OAI21_X1 U6186 ( .B1(n10539), .B2(n10466), .A(n5406), .ZN(P1_U3356) );
  AND2_X1 U6187 ( .A1(n5408), .A2(n5407), .ZN(n5406) );
  OR2_X1 U6188 ( .A1(n10540), .A2(n10504), .ZN(n5408) );
  AOI21_X1 U6189 ( .B1(n10537), .B2(n10520), .A(n8948), .ZN(n5407) );
  NOR2_X1 U6190 ( .A1(n5181), .A2(n5318), .ZN(n5317) );
  NAND2_X1 U6191 ( .A1(n6355), .A2(n11116), .ZN(n5320) );
  OAI21_X1 U6192 ( .B1(n6355), .B2(n11117), .A(n5254), .ZN(n6353) );
  OR2_X1 U6193 ( .A1(n11120), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5254) );
  AND2_X1 U6194 ( .A1(n8342), .A2(n5220), .ZN(n5125) );
  INV_X2 U6195 ( .A(n7060), .ZN(n6900) );
  AND2_X1 U6196 ( .A1(n8468), .A2(n8463), .ZN(n5126) );
  INV_X1 U6197 ( .A(n8707), .ZN(n5240) );
  NAND2_X1 U6198 ( .A1(n6395), .A2(n6414), .ZN(n6413) );
  XOR2_X1 U6199 ( .A(n6752), .B(n6778), .Z(n5129) );
  INV_X1 U6200 ( .A(n8794), .ZN(n5522) );
  AND2_X1 U6201 ( .A1(n5619), .A2(n5923), .ZN(n5130) );
  INV_X1 U6202 ( .A(n7412), .ZN(n7546) );
  AND2_X1 U6203 ( .A1(n5334), .A2(n5333), .ZN(n5131) );
  OR2_X1 U6204 ( .A1(n8881), .A2(n5240), .ZN(n5132) );
  AND2_X1 U6205 ( .A1(n6298), .A2(n6243), .ZN(n10336) );
  INV_X1 U6206 ( .A(n10336), .ZN(n5403) );
  AND2_X1 U6207 ( .A1(n5298), .A2(n8862), .ZN(n5133) );
  AND4_X1 U6208 ( .A1(n6519), .A2(n6518), .A3(n6517), .A4(n6516), .ZN(n7203)
         );
  INV_X1 U6209 ( .A(n7203), .ZN(n5260) );
  AND2_X1 U6210 ( .A1(n5331), .A2(n5330), .ZN(n5134) );
  AND3_X1 U6211 ( .A1(n6484), .A2(n6453), .A3(n6467), .ZN(n5135) );
  AND2_X1 U6212 ( .A1(n5467), .A2(n9405), .ZN(n5136) );
  AND2_X1 U6213 ( .A1(n6765), .A2(n9165), .ZN(n5137) );
  INV_X1 U6214 ( .A(n9079), .ZN(n5433) );
  NAND2_X1 U6215 ( .A1(n7618), .A2(n5714), .ZN(n5676) );
  NOR2_X1 U6216 ( .A1(n8422), .A2(n8438), .ZN(n5138) );
  INV_X2 U6217 ( .A(n5857), .ZN(n5948) );
  XNOR2_X1 U6218 ( .A(n6807), .B(n6806), .ZN(n6819) );
  INV_X1 U6219 ( .A(n9887), .ZN(n5431) );
  INV_X1 U6220 ( .A(n6778), .ZN(n5297) );
  INV_X1 U6221 ( .A(n8733), .ZN(n5517) );
  NAND2_X1 U6222 ( .A1(n8972), .A2(n8971), .ZN(n5139) );
  NOR2_X1 U6223 ( .A1(n5799), .A2(n5798), .ZN(n5140) );
  OR2_X1 U6224 ( .A1(n10213), .A2(n7335), .ZN(n5141) );
  NAND2_X1 U6225 ( .A1(n9041), .A2(n8970), .ZN(n9033) );
  INV_X1 U6226 ( .A(n9223), .ZN(n5276) );
  INV_X1 U6227 ( .A(n9119), .ZN(n5491) );
  AND2_X1 U6228 ( .A1(n5491), .A2(n9180), .ZN(n5142) );
  INV_X1 U6229 ( .A(n5298), .ZN(n5397) );
  NAND2_X1 U6230 ( .A1(n8726), .A2(n8894), .ZN(n5298) );
  INV_X1 U6231 ( .A(n7410), .ZN(n7520) );
  AND2_X1 U6232 ( .A1(n10598), .A2(n10508), .ZN(n5143) );
  INV_X1 U6233 ( .A(n9883), .ZN(n5424) );
  INV_X1 U6234 ( .A(n10423), .ZN(n5368) );
  AND3_X1 U6235 ( .A1(n6286), .A2(n8818), .A3(n10928), .ZN(n5144) );
  OR2_X1 U6236 ( .A1(n5222), .A2(n8343), .ZN(n5145) );
  INV_X1 U6237 ( .A(n8822), .ZN(n5357) );
  AND2_X1 U6238 ( .A1(n5392), .A2(n8815), .ZN(n5146) );
  AND3_X1 U6239 ( .A1(n10059), .A2(n5583), .A3(n5581), .ZN(n5147) );
  NAND2_X1 U6240 ( .A1(n9077), .A2(n8975), .ZN(n8999) );
  NAND2_X1 U6241 ( .A1(n10598), .A2(n10195), .ZN(n8726) );
  AND2_X1 U6242 ( .A1(n5452), .A2(n5456), .ZN(n5148) );
  NAND2_X1 U6243 ( .A1(n6012), .A2(n6011), .ZN(n10197) );
  AND2_X1 U6244 ( .A1(n5301), .A2(n5299), .ZN(n5149) );
  NOR2_X1 U6245 ( .A1(n10012), .A2(n9934), .ZN(n5150) );
  NOR2_X1 U6246 ( .A1(n7153), .A2(n7416), .ZN(n5151) );
  AND2_X1 U6247 ( .A1(n11089), .A2(n10205), .ZN(n5152) );
  NAND2_X1 U6248 ( .A1(n5901), .A2(n5900), .ZN(n7946) );
  AND2_X1 U6249 ( .A1(n9939), .A2(n9228), .ZN(n5153) );
  AND2_X1 U6250 ( .A1(n8683), .A2(n8676), .ZN(n5154) );
  AND2_X1 U6251 ( .A1(n5659), .A2(n5232), .ZN(n5155) );
  AND2_X1 U6252 ( .A1(n5368), .A2(n6296), .ZN(n5156) );
  INV_X1 U6253 ( .A(n5669), .ZN(n5668) );
  NAND2_X1 U6254 ( .A1(n5670), .A2(n8956), .ZN(n5669) );
  AND2_X1 U6255 ( .A1(n10612), .A2(n10203), .ZN(n5157) );
  AND2_X1 U6256 ( .A1(n10325), .A2(n6257), .ZN(n8939) );
  AND2_X1 U6257 ( .A1(n5600), .A2(n5599), .ZN(n5158) );
  NAND2_X1 U6258 ( .A1(n6938), .A2(n6937), .ZN(n5159) );
  INV_X1 U6259 ( .A(n5125), .ZN(n5219) );
  AND2_X1 U6260 ( .A1(n10479), .A2(n10493), .ZN(n5160) );
  NAND2_X1 U6261 ( .A1(n5713), .A2(n5621), .ZN(n5161) );
  NOR2_X1 U6262 ( .A1(n7866), .A2(n10207), .ZN(n5162) );
  NOR2_X1 U6263 ( .A1(n8175), .A2(n7916), .ZN(n5163) );
  INV_X1 U6264 ( .A(n5230), .ZN(n5229) );
  NAND2_X1 U6265 ( .A1(n5139), .A2(n8970), .ZN(n5230) );
  NOR2_X1 U6266 ( .A1(n10020), .A2(n9963), .ZN(n5164) );
  NOR2_X1 U6267 ( .A1(n10578), .A2(n10474), .ZN(n5165) );
  AND2_X1 U6268 ( .A1(n9308), .A2(n9309), .ZN(n5166) );
  AND2_X1 U6269 ( .A1(n10012), .A2(n9934), .ZN(n5167) );
  INV_X1 U6270 ( .A(n5697), .ZN(n5696) );
  NAND2_X1 U6271 ( .A1(n8541), .A2(n9322), .ZN(n5697) );
  OR2_X1 U6272 ( .A1(n6017), .A2(n5735), .ZN(n5168) );
  INV_X1 U6273 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5803) );
  AND2_X1 U6274 ( .A1(n8840), .A2(n8780), .ZN(n8814) );
  AND2_X1 U6275 ( .A1(n5484), .A2(n9239), .ZN(n5169) );
  AND2_X1 U6276 ( .A1(n5988), .A2(SI_13_), .ZN(n5170) );
  AND2_X1 U6277 ( .A1(n5924), .A2(SI_10_), .ZN(n5171) );
  INV_X1 U6278 ( .A(n5713), .ZN(n5622) );
  INV_X1 U6279 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5746) );
  AND2_X1 U6280 ( .A1(n10620), .A2(n10313), .ZN(n8916) );
  INV_X1 U6281 ( .A(n8916), .ZN(n5345) );
  AND2_X1 U6282 ( .A1(n10338), .A2(n10325), .ZN(n5172) );
  AND2_X1 U6283 ( .A1(n5497), .A2(n6370), .ZN(n5173) );
  OR2_X1 U6284 ( .A1(n8335), .A2(n9194), .ZN(n5174) );
  OR2_X1 U6285 ( .A1(n9331), .A2(n7625), .ZN(n9156) );
  AND3_X1 U6286 ( .A1(n5135), .A2(n5658), .A3(n5701), .ZN(n5175) );
  AND2_X1 U6287 ( .A1(n8799), .A2(n8713), .ZN(n5176) );
  OR2_X1 U6288 ( .A1(n6992), .A2(n8389), .ZN(n5177) );
  INV_X1 U6289 ( .A(n7011), .ZN(n5563) );
  NOR2_X1 U6290 ( .A1(n10463), .A2(n5512), .ZN(n5511) );
  OR2_X1 U6291 ( .A1(n5445), .A2(n5446), .ZN(n5178) );
  AND2_X1 U6292 ( .A1(n5424), .A2(n6775), .ZN(n5179) );
  INV_X1 U6293 ( .A(n10498), .ZN(n10652) );
  NAND2_X1 U6294 ( .A1(n6061), .A2(n6060), .ZN(n10498) );
  NAND2_X1 U6295 ( .A1(n5228), .A2(n5139), .ZN(n5227) );
  AND2_X1 U6296 ( .A1(n5217), .A2(n5214), .ZN(n5213) );
  INV_X1 U6297 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5743) );
  INV_X1 U6298 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5631) );
  INV_X1 U6299 ( .A(n8666), .ZN(n5370) );
  INV_X2 U6300 ( .A(n5127), .ZN(n9244) );
  INV_X1 U6301 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5628) );
  AND2_X1 U6302 ( .A1(n6508), .A2(n6358), .ZN(n6510) );
  OR2_X1 U6303 ( .A1(n8960), .A2(n9963), .ZN(n5180) );
  AND2_X1 U6304 ( .A1(n10325), .A2(n8211), .ZN(n5181) );
  AND2_X1 U6305 ( .A1(n9246), .A2(n9245), .ZN(n9899) );
  INV_X1 U6306 ( .A(n9899), .ZN(n5436) );
  NAND2_X1 U6307 ( .A1(n5578), .A2(n6958), .ZN(n8167) );
  AND4_X1 U6308 ( .A1(n6578), .A2(n6577), .A3(n6576), .A4(n6575), .ZN(n8463)
         );
  NOR2_X1 U6309 ( .A1(n8587), .A2(n8588), .ZN(n5182) );
  INV_X1 U6310 ( .A(n10402), .ZN(n10426) );
  NOR2_X1 U6311 ( .A1(n10446), .A2(n10568), .ZN(n10402) );
  NAND2_X1 U6312 ( .A1(n8363), .A2(n5131), .ZN(n5335) );
  NOR2_X1 U6313 ( .A1(n8953), .A2(n8952), .ZN(n5183) );
  NAND2_X1 U6314 ( .A1(n6390), .A2(n6389), .ZN(n9996) );
  INV_X1 U6315 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U6316 ( .A1(n8946), .A2(n8945), .ZN(n5184) );
  AND2_X1 U6317 ( .A1(n6131), .A2(n6118), .ZN(n5185) );
  AND4_X2 U6318 ( .A1(n6844), .A2(n7764), .A3(n7763), .A4(n10942), .ZN(n11153)
         );
  INV_X1 U6319 ( .A(n11153), .ZN(n5476) );
  NAND2_X1 U6320 ( .A1(n6804), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U6321 ( .A1(n7711), .A2(n5478), .ZN(n7900) );
  XNOR2_X1 U6322 ( .A(n6320), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6351) );
  XNOR2_X1 U6323 ( .A(n6810), .B(n6809), .ZN(n6823) );
  NAND2_X1 U6324 ( .A1(n6047), .A2(n6046), .ZN(n10594) );
  INV_X1 U6325 ( .A(n10594), .ZN(n5333) );
  INV_X1 U6326 ( .A(n10162), .ZN(n5566) );
  NAND2_X1 U6327 ( .A1(n5579), .A2(n6896), .ZN(n7495) );
  OAI21_X1 U6328 ( .B1(n10161), .B2(n5567), .A(n5564), .ZN(n7858) );
  INV_X1 U6329 ( .A(n10905), .ZN(n8438) );
  NOR2_X1 U6330 ( .A1(n8189), .A2(n8190), .ZN(n5186) );
  OR2_X1 U6331 ( .A1(n8439), .A2(n8438), .ZN(n5187) );
  AND2_X1 U6332 ( .A1(n6286), .A2(n7447), .ZN(n5188) );
  NAND2_X1 U6333 ( .A1(n8543), .A2(n8542), .ZN(n5189) );
  AND2_X1 U6334 ( .A1(n6741), .A2(n9662), .ZN(n5190) );
  AOI22_X1 U6335 ( .A1(n7729), .A2(n7728), .B1(n7727), .B2(n9331), .ZN(n7730)
         );
  AND2_X1 U6336 ( .A1(n8429), .A2(n10905), .ZN(n5191) );
  NAND2_X1 U6337 ( .A1(n5882), .A2(n5881), .ZN(n7866) );
  INV_X1 U6338 ( .A(n7866), .ZN(n5253) );
  AND2_X2 U6339 ( .A1(n6354), .A2(n7567), .ZN(n11120) );
  AND2_X2 U6340 ( .A1(n6354), .A2(n7098), .ZN(n11116) );
  INV_X1 U6341 ( .A(n6858), .ZN(n6861) );
  NAND2_X1 U6342 ( .A1(n5934), .A2(n5933), .ZN(n11089) );
  INV_X1 U6343 ( .A(n11089), .ZN(n5330) );
  NAND2_X1 U6344 ( .A1(n6513), .A2(n6512), .ZN(n8048) );
  INV_X1 U6345 ( .A(n8048), .ZN(n5261) );
  AND2_X1 U6346 ( .A1(n9104), .A2(n7138), .ZN(n10967) );
  INV_X1 U6347 ( .A(n10967), .ZN(n10935) );
  NOR2_X1 U6348 ( .A1(n7986), .A2(n7987), .ZN(n5192) );
  AND2_X1 U6349 ( .A1(n5461), .A2(n5460), .ZN(n5193) );
  OR2_X1 U6350 ( .A1(n11153), .A2(n6845), .ZN(n5194) );
  INV_X1 U6351 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5324) );
  INV_X1 U6352 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n5611) );
  NOR2_X4 U6353 ( .A1(n7108), .A2(n5124), .ZN(n10189) );
  INV_X1 U6354 ( .A(n6942), .ZN(n5568) );
  AND2_X2 U6355 ( .A1(n5231), .A2(n5175), .ZN(n6365) );
  NOR2_X2 U6356 ( .A1(n7415), .A2(n7401), .ZN(n7420) );
  NAND2_X1 U6357 ( .A1(n5381), .A2(n5380), .ZN(n5379) );
  INV_X1 U6358 ( .A(n5893), .ZN(n5621) );
  OAI21_X1 U6359 ( .B1(n5872), .B2(n5313), .A(n5312), .ZN(n5617) );
  NAND2_X1 U6360 ( .A1(n6057), .A2(n6056), .ZN(n6079) );
  NAND2_X1 U6361 ( .A1(n5361), .A2(n5364), .ZN(n5359) );
  INV_X1 U6362 ( .A(n8817), .ZN(n8813) );
  NAND2_X1 U6363 ( .A1(n5523), .A2(n5340), .ZN(n5339) );
  OAI21_X1 U6364 ( .B1(n10540), .B2(n11000), .A(n5338), .ZN(n5337) );
  OAI211_X2 U6365 ( .C1(n5857), .C2(n7169), .A(n5775), .B(n5774), .ZN(n7704)
         );
  NAND2_X1 U6366 ( .A1(n5437), .A2(n6566), .ZN(n8412) );
  NOR2_X2 U6367 ( .A1(n6384), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5199) );
  OAI21_X1 U6368 ( .B1(n8218), .B2(n8284), .A(n6555), .ZN(n8329) );
  NAND3_X1 U6369 ( .A1(n6859), .A2(n6860), .A3(n5707), .ZN(n7284) );
  NAND3_X1 U6370 ( .A1(n5203), .A2(n5709), .A3(n7116), .ZN(P1_U3214) );
  NAND2_X1 U6371 ( .A1(n7486), .A2(n7488), .ZN(n5579) );
  NAND2_X1 U6372 ( .A1(n5935), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5957) );
  NOR2_X1 U6373 ( .A1(n8499), .A2(n8507), .ZN(n8577) );
  XNOR2_X1 U6374 ( .A(n7676), .B(n7693), .ZN(n7518) );
  NOR2_X2 U6375 ( .A1(n9357), .A2(n8581), .ZN(n9378) );
  NOR2_X1 U6376 ( .A1(n10916), .A2(n5148), .ZN(n8425) );
  NOR2_X1 U6377 ( .A1(n10893), .A2(n10892), .ZN(n10891) );
  NOR2_X1 U6378 ( .A1(n9390), .A2(n8583), .ZN(n8585) );
  INV_X1 U6379 ( .A(n8283), .ZN(n5216) );
  NAND2_X1 U6380 ( .A1(n5211), .A2(n5212), .ZN(n8471) );
  NAND2_X1 U6381 ( .A1(n8283), .A2(n5213), .ZN(n5211) );
  AOI21_X1 U6382 ( .B1(n8283), .B2(n8282), .A(n8281), .ZN(n8344) );
  INV_X1 U6383 ( .A(n8282), .ZN(n5222) );
  NAND2_X1 U6384 ( .A1(n5698), .A2(n9008), .ZN(n9041) );
  NAND3_X1 U6385 ( .A1(n5698), .A2(n5227), .A3(n9008), .ZN(n5223) );
  AND3_X1 U6386 ( .A1(n5135), .A2(n5231), .A3(n5658), .ZN(n6508) );
  NAND2_X1 U6387 ( .A1(n5658), .A2(n6395), .ZN(n6427) );
  NAND2_X2 U6388 ( .A1(n7153), .A2(n7159), .ZN(n9101) );
  XNOR2_X2 U6389 ( .A(n6387), .B(n6386), .ZN(n6789) );
  NAND3_X1 U6390 ( .A1(n5625), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5629) );
  INV_X1 U6391 ( .A(n5838), .ZN(n5243) );
  OAI211_X1 U6392 ( .C1(n5249), .C2(n5368), .A(n10432), .B(n10512), .ZN(n10435) );
  NAND2_X1 U6393 ( .A1(n10337), .A2(n10336), .ZN(n10335) );
  NAND2_X1 U6394 ( .A1(n5308), .A2(n5250), .ZN(n5307) );
  OAI21_X1 U6395 ( .B1(n10337), .B2(n8834), .A(n5251), .ZN(n5250) );
  NAND2_X1 U6396 ( .A1(n5872), .A2(n5264), .ZN(n5263) );
  NAND3_X1 U6397 ( .A1(n9234), .A2(n5275), .A3(n9233), .ZN(n5270) );
  INV_X1 U6398 ( .A(n9224), .ZN(n5271) );
  INV_X1 U6399 ( .A(n9229), .ZN(n5274) );
  AOI21_X2 U6400 ( .B1(n5287), .B2(n5286), .A(n5166), .ZN(n9310) );
  NAND3_X1 U6401 ( .A1(n5632), .A2(n5635), .A3(n5290), .ZN(n5289) );
  OAI21_X1 U6402 ( .B1(n9263), .B2(n5296), .A(n5294), .ZN(n5637) );
  INV_X1 U6403 ( .A(n5291), .ZN(n5636) );
  NAND2_X2 U6404 ( .A1(n5629), .A2(n5630), .ZN(n5785) );
  NAND3_X1 U6405 ( .A1(n5630), .A2(n5629), .A3(n5757), .ZN(n6406) );
  OAI21_X1 U6406 ( .B1(n5970), .B2(n5969), .A(n5968), .ZN(n5987) );
  INV_X1 U6407 ( .A(n5304), .ZN(n5303) );
  NAND2_X1 U6408 ( .A1(n5305), .A2(n5986), .ZN(n5304) );
  NAND2_X1 U6409 ( .A1(n5870), .A2(n5314), .ZN(n5311) );
  NAND2_X1 U6410 ( .A1(n5316), .A2(n5874), .ZN(n5892) );
  NAND2_X1 U6411 ( .A1(n5320), .A2(n5317), .ZN(P1_U3550) );
  NOR2_X1 U6412 ( .A1(n11116), .A2(n5319), .ZN(n5318) );
  NAND2_X1 U6413 ( .A1(n5120), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5323) );
  OAI21_X1 U6414 ( .B1(n5120), .B2(n5324), .A(n5323), .ZN(n5820) );
  NAND2_X2 U6415 ( .A1(n7159), .A2(P2_U3151), .ZN(n8985) );
  MUX2_X1 U6416 ( .A(n9797), .B(n7631), .S(n5120), .Z(n6028) );
  MUX2_X1 U6417 ( .A(n9583), .B(n7311), .S(n5120), .Z(n5989) );
  MUX2_X1 U6418 ( .A(n9573), .B(n7912), .S(n5120), .Z(n6080) );
  MUX2_X1 U6419 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n5120), .Z(n6203) );
  MUX2_X1 U6420 ( .A(n9764), .B(n9098), .S(n5120), .Z(n8642) );
  MUX2_X1 U6421 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5120), .Z(n8657) );
  OAI21_X1 U6422 ( .B1(n5298), .B2(n8893), .A(n8862), .ZN(n5325) );
  NOR2_X2 U6423 ( .A1(n7599), .A2(n10995), .ZN(n7598) );
  INV_X1 U6424 ( .A(n7468), .ZN(n5328) );
  NAND2_X1 U6425 ( .A1(n5134), .A2(n5329), .ZN(n8147) );
  AND2_X1 U6426 ( .A1(n5134), .A2(n7849), .ZN(n7954) );
  NAND2_X1 U6427 ( .A1(n5332), .A2(n8363), .ZN(n10496) );
  INV_X1 U6428 ( .A(n5335), .ZN(n10519) );
  OAI21_X1 U6429 ( .B1(n6286), .B2(n7451), .A(n7450), .ZN(n7454) );
  NAND2_X1 U6430 ( .A1(n6286), .A2(n7451), .ZN(n7450) );
  NOR2_X1 U6431 ( .A1(n5347), .A2(n10320), .ZN(n5346) );
  NAND3_X4 U6432 ( .A1(n5350), .A2(n5120), .A3(n5348), .ZN(n8777) );
  NAND2_X1 U6433 ( .A1(n5351), .A2(n5124), .ZN(n5350) );
  NAND2_X2 U6434 ( .A1(n5352), .A2(n5353), .ZN(n10748) );
  NAND2_X1 U6435 ( .A1(n8746), .A2(n5358), .ZN(n5355) );
  NAND2_X1 U6436 ( .A1(n5355), .A2(n5356), .ZN(n8752) );
  AND2_X1 U6437 ( .A1(n5359), .A2(n5365), .ZN(n5358) );
  OAI21_X1 U6438 ( .B1(n5374), .B2(n8870), .A(n5369), .ZN(n7376) );
  NAND2_X1 U6439 ( .A1(n5375), .A2(n8666), .ZN(n5372) );
  NAND3_X1 U6440 ( .A1(n8723), .A2(n5392), .A3(n8782), .ZN(n5382) );
  NAND2_X1 U6441 ( .A1(n8722), .A2(n5146), .ZN(n5383) );
  NAND3_X1 U6442 ( .A1(n5391), .A2(n5386), .A3(n5385), .ZN(n8727) );
  NAND2_X1 U6443 ( .A1(n5395), .A2(n5389), .ZN(n5385) );
  NOR2_X1 U6444 ( .A1(n5390), .A2(n5387), .ZN(n5386) );
  NAND2_X1 U6445 ( .A1(n10337), .A2(n5402), .ZN(n5399) );
  NAND2_X1 U6446 ( .A1(n5399), .A2(n5400), .ZN(n8941) );
  NAND2_X1 U6447 ( .A1(n5785), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5405) );
  OAI21_X1 U6448 ( .B1(n5785), .B2(n7162), .A(n5405), .ZN(n5795) );
  NAND2_X1 U6449 ( .A1(n5411), .A2(n5409), .ZN(n6474) );
  NAND2_X1 U6450 ( .A1(n6433), .A2(n5414), .ZN(n5411) );
  OAI21_X1 U6451 ( .B1(n9900), .B2(n9899), .A(n5435), .ZN(n9888) );
  NAND2_X1 U6452 ( .A1(n9089), .A2(n9251), .ZN(n5434) );
  NAND2_X1 U6453 ( .A1(n9960), .A2(n5440), .ZN(n5438) );
  NAND2_X1 U6454 ( .A1(n5438), .A2(n5439), .ZN(n9933) );
  NAND2_X1 U6455 ( .A1(n5443), .A2(n11157), .ZN(n7150) );
  NAND2_X1 U6456 ( .A1(n8989), .A2(n5477), .ZN(n5443) );
  AOI21_X2 U6457 ( .B1(n5129), .B2(n10935), .A(n6796), .ZN(n8989) );
  AND2_X1 U6458 ( .A1(n7153), .A2(n5178), .ZN(n5444) );
  NOR2_X2 U6459 ( .A1(n5151), .A2(n5444), .ZN(n8073) );
  AOI21_X2 U6460 ( .B1(n6685), .B2(n5447), .A(n5167), .ZN(n9912) );
  NAND2_X1 U6461 ( .A1(n5450), .A2(n5449), .ZN(n6532) );
  AND2_X1 U6462 ( .A1(n5705), .A2(n6520), .ZN(n5449) );
  NAND3_X1 U6463 ( .A1(n7321), .A2(P2_IR_REG_2__SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n5451) );
  NOR2_X1 U6464 ( .A1(n8187), .A2(n8186), .ZN(n8423) );
  NAND2_X1 U6465 ( .A1(n8187), .A2(n5457), .ZN(n5452) );
  OAI211_X1 U6466 ( .C1(n8187), .C2(n5455), .A(n5454), .B(n5453), .ZN(n10917)
         );
  AOI22_X1 U6467 ( .A1(n5456), .A2(n8422), .B1(n8186), .B2(n5138), .ZN(n5453)
         );
  NAND2_X1 U6468 ( .A1(n8187), .A2(n5138), .ZN(n5454) );
  AOI21_X1 U6469 ( .B1(n8186), .B2(n5457), .A(n10905), .ZN(n5456) );
  INV_X1 U6470 ( .A(n8422), .ZN(n5457) );
  NAND2_X1 U6471 ( .A1(n5462), .A2(n7409), .ZN(n5458) );
  INV_X1 U6472 ( .A(n7411), .ZN(n5462) );
  XNOR2_X1 U6473 ( .A(n7408), .B(n7412), .ZN(n7536) );
  NAND2_X1 U6474 ( .A1(n8583), .A2(n5469), .ZN(n5467) );
  NOR2_X1 U6475 ( .A1(n9391), .A2(n6615), .ZN(n9390) );
  NAND2_X1 U6476 ( .A1(n5466), .A2(n5467), .ZN(n9406) );
  AND2_X2 U6478 ( .A1(n5471), .A2(n5470), .ZN(n8580) );
  NOR2_X1 U6479 ( .A1(n7678), .A2(n7677), .ZN(n10893) );
  NOR2_X1 U6480 ( .A1(n6448), .A2(n7518), .ZN(n7677) );
  INV_X1 U6481 ( .A(n8696), .ZN(n8706) );
  OAI211_X1 U6482 ( .C1(n8989), .C2(n5476), .A(n5474), .B(n5194), .ZN(P2_U3488) );
  NAND2_X1 U6483 ( .A1(n6772), .A2(n5480), .ZN(n5479) );
  NAND2_X1 U6484 ( .A1(n9891), .A2(n5179), .ZN(n9880) );
  NAND2_X1 U6485 ( .A1(n6764), .A2(n5137), .ZN(n8039) );
  NAND2_X1 U6486 ( .A1(n8039), .A2(n9169), .ZN(n8061) );
  OAI21_X1 U6487 ( .B1(n9926), .B2(n9236), .A(n9115), .ZN(n9911) );
  NAND2_X1 U6488 ( .A1(n9236), .A2(n9115), .ZN(n5486) );
  INV_X1 U6489 ( .A(n9896), .ZN(n6774) );
  NAND2_X1 U6490 ( .A1(n6766), .A2(n5489), .ZN(n5487) );
  NAND2_X1 U6491 ( .A1(n5487), .A2(n5488), .ZN(n8418) );
  NAND2_X1 U6492 ( .A1(n5493), .A2(n5492), .ZN(n8529) );
  NAND2_X1 U6493 ( .A1(n6365), .A2(n5497), .ZN(n5496) );
  MUX2_X1 U6494 ( .A(n5498), .B(P1_REG1_REG_29__SCAN_IN), .S(n11115), .Z(
        P1_U3551) );
  MUX2_X1 U6495 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n5498), .S(n11120), .Z(
        P1_U3519) );
  NAND2_X1 U6496 ( .A1(n7745), .A2(n5128), .ZN(n5500) );
  NAND2_X1 U6497 ( .A1(n8320), .A2(n5506), .ZN(n5505) );
  NAND2_X1 U6498 ( .A1(n6074), .A2(n5511), .ZN(n5509) );
  NAND2_X1 U6499 ( .A1(n5509), .A2(n5510), .ZN(n10445) );
  OAI21_X1 U6500 ( .B1(n7846), .B2(n5522), .A(n5520), .ZN(n7919) );
  NAND2_X1 U6501 ( .A1(n5519), .A2(n5518), .ZN(n5944) );
  NAND2_X1 U6502 ( .A1(n7846), .A2(n5520), .ZN(n5519) );
  INV_X1 U6503 ( .A(n5753), .ZN(n5538) );
  XNOR2_X1 U6504 ( .A(n5539), .B(n5122), .ZN(n5543) );
  NAND2_X1 U6505 ( .A1(n5540), .A2(n5753), .ZN(n10214) );
  INV_X1 U6506 ( .A(n5543), .ZN(n6286) );
  NAND2_X1 U6507 ( .A1(n5543), .A2(n5542), .ZN(n7445) );
  NAND3_X1 U6508 ( .A1(n5545), .A2(n8645), .A3(P1_REG1_REG_0__SCAN_IN), .ZN(
        n5544) );
  INV_X1 U6509 ( .A(n8645), .ZN(n5738) );
  INV_X1 U6510 ( .A(n5736), .ZN(n5545) );
  INV_X1 U6511 ( .A(n5730), .ZN(n5546) );
  NAND2_X1 U6512 ( .A1(n5726), .A2(n5708), .ZN(n6266) );
  NAND3_X1 U6513 ( .A1(n5547), .A2(n5546), .A3(n5726), .ZN(n5742) );
  AND4_X2 U6514 ( .A1(n5546), .A2(n5726), .A3(n5547), .A4(n5743), .ZN(n5732)
         );
  NAND3_X1 U6515 ( .A1(n5549), .A2(n10153), .A3(n5548), .ZN(n10066) );
  NAND3_X1 U6516 ( .A1(n5168), .A2(n5739), .A3(n5550), .ZN(n6858) );
  NAND2_X1 U6517 ( .A1(n8269), .A2(n5553), .ZN(n5552) );
  NAND2_X1 U6518 ( .A1(n5560), .A2(n5561), .ZN(n10107) );
  NAND3_X1 U6519 ( .A1(n7001), .A2(n7011), .A3(n10185), .ZN(n5560) );
  OAI21_X2 U6520 ( .B1(n10161), .B2(n10163), .A(n10162), .ZN(n7670) );
  OR2_X2 U6521 ( .A1(n10088), .A2(n10087), .ZN(n5572) );
  INV_X1 U6522 ( .A(n7935), .ZN(n5575) );
  AOI21_X2 U6523 ( .B1(n5575), .B2(n5574), .A(n5573), .ZN(n11084) );
  NAND3_X1 U6524 ( .A1(n5579), .A2(n6896), .A3(n6903), .ZN(n7496) );
  OAI21_X2 U6525 ( .B1(n10078), .B2(n5585), .A(n5147), .ZN(n10057) );
  INV_X1 U6526 ( .A(n5588), .ZN(n10142) );
  INV_X1 U6527 ( .A(n7061), .ZN(n5589) );
  NAND2_X1 U6528 ( .A1(n8430), .A2(n5191), .ZN(n5595) );
  OAI211_X1 U6529 ( .C1(n8430), .C2(n10905), .A(n5592), .B(n5595), .ZN(n10911)
         );
  NAND2_X1 U6530 ( .A1(n5591), .A2(n8438), .ZN(n5594) );
  NAND2_X1 U6531 ( .A1(n8430), .A2(n8429), .ZN(n5591) );
  OR2_X1 U6532 ( .A1(n8429), .A2(n10905), .ZN(n5593) );
  NAND2_X1 U6533 ( .A1(n10911), .A2(n5594), .ZN(n8431) );
  XNOR2_X1 U6534 ( .A(n8590), .B(n9371), .ZN(n9359) );
  NAND2_X1 U6535 ( .A1(n8190), .A2(n5604), .ZN(n5602) );
  OAI21_X1 U6536 ( .B1(n8504), .B2(n5606), .A(n5605), .ZN(n9341) );
  NAND2_X1 U6537 ( .A1(n8594), .A2(n5612), .ZN(n5608) );
  NOR2_X1 U6538 ( .A1(n9395), .A2(n11152), .ZN(n9394) );
  NOR2_X1 U6539 ( .A1(n9394), .A2(n8594), .ZN(n8597) );
  INV_X1 U6540 ( .A(n5623), .ZN(n5627) );
  NAND3_X1 U6541 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n5740), .A3(n9421), .ZN(
        n5624) );
  NAND3_X1 U6542 ( .A1(n5630), .A2(n5629), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n5626) );
  NAND3_X1 U6543 ( .A1(n9266), .A2(n9244), .A3(n5636), .ZN(n5635) );
  NAND2_X1 U6544 ( .A1(n6187), .A2(n5641), .ZN(n5640) );
  NAND2_X1 U6545 ( .A1(n6187), .A2(n6186), .ZN(n6202) );
  INV_X1 U6546 ( .A(n6186), .ZN(n5642) );
  NAND2_X1 U6547 ( .A1(n5644), .A2(n5185), .ZN(n6134) );
  INV_X1 U6548 ( .A(n7815), .ZN(n5675) );
  NAND2_X1 U6549 ( .A1(n5678), .A2(n5679), .ZN(n8979) );
  NAND2_X1 U6550 ( .A1(n9075), .A2(n5680), .ZN(n5678) );
  OAI21_X1 U6551 ( .B1(n9075), .B2(n5682), .A(n5680), .ZN(n9000) );
  NAND2_X1 U6552 ( .A1(n5683), .A2(n5684), .ZN(n6755) );
  NAND2_X1 U6553 ( .A1(n6754), .A2(n5686), .ZN(n5683) );
  NAND2_X1 U6554 ( .A1(n6754), .A2(n6753), .ZN(n5685) );
  NAND2_X1 U6555 ( .A1(n5687), .A2(n5688), .ZN(n8953) );
  NAND2_X1 U6556 ( .A1(n8553), .A2(n5692), .ZN(n5687) );
  NOR2_X1 U6557 ( .A1(n8552), .A2(n5696), .ZN(n8565) );
  OAI21_X1 U6558 ( .B1(n6508), .B2(n6521), .A(n5699), .ZN(n6545) );
  NAND2_X1 U6559 ( .A1(n6818), .A2(n5702), .ZN(n6820) );
  INV_X1 U6560 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U6561 ( .A1(n6365), .A2(n5704), .ZN(n6804) );
  OR2_X1 U6562 ( .A1(n10324), .A2(n6301), .ZN(n6256) );
  OR2_X1 U6563 ( .A1(n10355), .A2(n6301), .ZN(n6218) );
  AOI21_X2 U6564 ( .B1(n7964), .B2(n6507), .A(n5711), .ZN(n8042) );
  NAND2_X2 U6565 ( .A1(n5118), .A2(n7059), .ZN(n6887) );
  CLKBUF_X1 U6566 ( .A(n7935), .Z(n7936) );
  NAND2_X1 U6567 ( .A1(n9142), .A2(n9149), .ZN(n7975) );
  AND3_X1 U6568 ( .A1(n5721), .A2(n5720), .A3(n5823), .ZN(n5722) );
  CLKBUF_X1 U6569 ( .A(n8269), .Z(n8297) );
  INV_X1 U6570 ( .A(n6997), .ZN(n7000) );
  INV_X1 U6571 ( .A(n6872), .ZN(n6875) );
  OR2_X1 U6572 ( .A1(n5732), .A2(n5803), .ZN(n5734) );
  OR2_X1 U6573 ( .A1(n9271), .A2(n7138), .ZN(n7353) );
  XNOR2_X1 U6574 ( .A(n6890), .B(n5119), .ZN(n6893) );
  NAND2_X1 U6575 ( .A1(n6626), .A2(n6625), .ZN(n6640) );
  NAND2_X1 U6576 ( .A1(n6558), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6626) );
  XNOR2_X1 U6577 ( .A(n9440), .B(n9448), .ZN(n9444) );
  INV_X1 U6578 ( .A(n9306), .ZN(n9989) );
  AOI21_X1 U6579 ( .B1(n8860), .B2(n8859), .A(n8858), .ZN(n8930) );
  NAND2_X1 U6580 ( .A1(n8817), .A2(n8816), .ZN(n8860) );
  NAND2_X1 U6581 ( .A1(n8647), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5793) );
  XNOR2_X1 U6582 ( .A(n8226), .B(n8227), .ZN(n8228) );
  NAND2_X1 U6583 ( .A1(n9063), .A2(n8962), .ZN(n8963) );
  OR2_X1 U6584 ( .A1(n11075), .A2(n9328), .ZN(n5705) );
  INV_X1 U6585 ( .A(n11015), .ZN(n10466) );
  INV_X1 U6586 ( .A(n11015), .ZN(n10529) );
  INV_X1 U6587 ( .A(n7696), .ZN(n10903) );
  INV_X1 U6588 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7679) );
  INV_X1 U6589 ( .A(n8524), .ZN(n9961) );
  INV_X1 U6590 ( .A(n8001), .ZN(n7990) );
  AND4_X1 U6591 ( .A1(n5725), .A2(n5724), .A3(n5723), .A4(n6031), .ZN(n5708)
         );
  OR2_X1 U6592 ( .A1(n10628), .A2(n10183), .ZN(n5709) );
  NOR2_X1 U6593 ( .A1(n6506), .A2(n7965), .ZN(n5711) );
  AND2_X1 U6594 ( .A1(n8922), .A2(n8856), .ZN(n5712) );
  INV_X1 U6595 ( .A(n8102), .ZN(n8193) );
  AND4_X1 U6596 ( .A1(n6381), .A2(n6380), .A3(n6379), .A4(n6378), .ZN(n9079)
         );
  INV_X1 U6597 ( .A(n8940), .ZN(n8769) );
  INV_X1 U6598 ( .A(n8335), .ZN(n6768) );
  OR2_X1 U6599 ( .A1(n11124), .A2(n8414), .ZN(n9195) );
  AND2_X1 U6600 ( .A1(n7729), .A2(n7723), .ZN(n5714) );
  XNOR2_X1 U6601 ( .A(n7348), .B(n6399), .ZN(n7480) );
  NAND2_X1 U6602 ( .A1(n9270), .A2(n8069), .ZN(n8068) );
  OR2_X1 U6603 ( .A1(n10341), .A2(n10325), .ZN(n5715) );
  OAI22_X1 U6604 ( .A1(n8228), .A2(n9328), .B1(n8227), .B2(n8226), .ZN(n8283)
         );
  INV_X1 U6605 ( .A(n9196), .ZN(n6579) );
  AND2_X1 U6606 ( .A1(n9223), .A2(n9225), .ZN(n9969) );
  INV_X1 U6607 ( .A(n9969), .ZN(n6664) );
  NAND2_X1 U6608 ( .A1(n8703), .A2(n8782), .ZN(n8704) );
  OAI211_X1 U6609 ( .C1(n8706), .C2(n8782), .A(n8705), .B(n8704), .ZN(n8712)
         );
  INV_X1 U6610 ( .A(n8767), .ZN(n8768) );
  INV_X1 U6611 ( .A(n7406), .ZN(n7407) );
  NAND2_X1 U6612 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  NAND2_X1 U6613 ( .A1(n7608), .A2(n9335), .ZN(n7606) );
  INV_X1 U6614 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6802) );
  AND2_X1 U6615 ( .A1(n7344), .A2(n7343), .ZN(n7345) );
  NOR2_X1 U6616 ( .A1(n7410), .A2(n6436), .ZN(n7516) );
  INV_X1 U6617 ( .A(n9281), .ZN(n6765) );
  OR2_X1 U6618 ( .A1(n9091), .A2(n7323), .ZN(n6392) );
  NAND2_X1 U6619 ( .A1(n6744), .A2(n6743), .ZN(n6797) );
  OR2_X1 U6620 ( .A1(n6722), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6375) );
  INV_X1 U6621 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9027) );
  INV_X1 U6622 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U6623 ( .A1(n6580), .A2(n6579), .ZN(n8410) );
  INV_X1 U6624 ( .A(n8073), .ZN(n6398) );
  INV_X1 U6625 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6467) );
  INV_X1 U6626 ( .A(n7939), .ZN(n6949) );
  INV_X1 U6627 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5884) );
  INV_X1 U6628 ( .A(SI_23_), .ZN(n9674) );
  INV_X1 U6629 ( .A(SI_14_), .ZN(n9689) );
  INV_X1 U6630 ( .A(SI_9_), .ZN(n9699) );
  INV_X1 U6631 ( .A(n7730), .ZN(n7731) );
  OR2_X1 U6632 ( .A1(n8961), .A2(n9230), .ZN(n8962) );
  AND2_X1 U6633 ( .A1(n8280), .A2(n8279), .ZN(n8281) );
  INV_X1 U6634 ( .A(n6701), .ZN(n6600) );
  NOR2_X1 U6635 ( .A1(n8003), .A2(n8002), .ZN(n8006) );
  NOR2_X1 U6636 ( .A1(n8501), .A2(n8222), .ZN(n8496) );
  INV_X1 U6637 ( .A(n8575), .ZN(n8576) );
  AND2_X1 U6638 ( .A1(n6731), .A2(n9522), .ZN(n9433) );
  NOR2_X1 U6639 ( .A1(n6375), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6731) );
  NAND2_X1 U6640 ( .A1(n6712), .A2(n9735), .ZN(n6722) );
  INV_X1 U6641 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9535) );
  INV_X1 U6642 ( .A(n9409), .ZN(n9424) );
  INV_X1 U6643 ( .A(n9195), .ZN(n6767) );
  INV_X1 U6644 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6567) );
  INV_X1 U6645 ( .A(n7498), .ZN(n6903) );
  NAND2_X1 U6646 ( .A1(n6858), .A2(n6862), .ZN(n6865) );
  NAND2_X1 U6647 ( .A1(n6089), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6108) );
  OR2_X1 U6648 ( .A1(n6063), .A2(n6062), .ZN(n6091) );
  AND2_X1 U6649 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5830) );
  NAND2_X1 U6650 ( .A1(n6190), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6212) );
  OR2_X1 U6651 ( .A1(n6159), .A2(n10061), .ZN(n6175) );
  NAND2_X1 U6652 ( .A1(n6137), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6159) );
  INV_X1 U6653 ( .A(n8728), .ZN(n8895) );
  OR2_X1 U6654 ( .A1(n5885), .A2(n5884), .ZN(n5904) );
  INV_X1 U6655 ( .A(n10352), .ZN(n10343) );
  AOI21_X1 U6656 ( .B1(n7182), .B2(n7188), .A(n6328), .ZN(n7565) );
  INV_X1 U6657 ( .A(SI_18_), .ZN(n9655) );
  INV_X1 U6658 ( .A(SI_12_), .ZN(n9693) );
  INV_X1 U6659 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9518) );
  INV_X1 U6660 ( .A(n7614), .ZN(n7634) );
  INV_X1 U6661 ( .A(n6477), .ZN(n6784) );
  INV_X1 U6662 ( .A(n8605), .ZN(n8498) );
  INV_X1 U6663 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9381) );
  OR2_X1 U6664 ( .A1(P2_U3150), .A2(n7314), .ZN(n9422) );
  XNOR2_X1 U6665 ( .A(n6790), .B(n9412), .ZN(n9875) );
  AND2_X1 U6666 ( .A1(n9180), .A2(n9178), .ZN(n9285) );
  INV_X1 U6667 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U6668 ( .A1(n6763), .A2(n9146), .ZN(n8082) );
  NAND2_X1 U6669 ( .A1(n6521), .A2(n6414), .ZN(n6415) );
  AND2_X1 U6670 ( .A1(n7086), .A2(n7085), .ZN(n7095) );
  AND2_X1 U6671 ( .A1(n5917), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5935) );
  AND2_X1 U6672 ( .A1(n6309), .A2(n6308), .ZN(n8765) );
  INV_X1 U6673 ( .A(n6301), .ZN(n6235) );
  INV_X1 U6674 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7247) );
  INV_X1 U6675 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8301) );
  OR2_X1 U6676 ( .A1(n10756), .A2(n7248), .ZN(n10829) );
  OAI21_X1 U6677 ( .B1(n10369), .B2(n6199), .A(n6198), .ZN(n10351) );
  INV_X1 U6678 ( .A(n8804), .ZN(n10514) );
  AND2_X1 U6679 ( .A1(n8662), .A2(n8715), .ZN(n8799) );
  INV_X1 U6680 ( .A(n11109), .ZN(n10996) );
  INV_X1 U6681 ( .A(n10512), .ZN(n10929) );
  AND2_X1 U6682 ( .A1(n6838), .A2(n6837), .ZN(n6839) );
  INV_X1 U6683 ( .A(n9019), .ZN(n8568) );
  INV_X1 U6684 ( .A(n9067), .ZN(n9085) );
  AND4_X1 U6685 ( .A1(n6653), .A2(n6652), .A3(n6651), .A4(n6650), .ZN(n8954)
         );
  AND2_X1 U6686 ( .A1(n7317), .A2(n8533), .ZN(n10865) );
  INV_X1 U6687 ( .A(n9422), .ZN(n10907) );
  INV_X1 U6688 ( .A(n9426), .ZN(n10923) );
  INV_X1 U6689 ( .A(n8523), .ZN(n10944) );
  INV_X1 U6690 ( .A(n9185), .ZN(n9290) );
  INV_X1 U6691 ( .A(n9984), .ZN(n11043) );
  INV_X1 U6692 ( .A(n10950), .ZN(n11041) );
  AND2_X1 U6693 ( .A1(n7141), .A2(n6843), .ZN(n7764) );
  INV_X1 U6694 ( .A(n11132), .ZN(n11146) );
  INV_X1 U6695 ( .A(n11127), .ZN(n11151) );
  INV_X1 U6696 ( .A(n11071), .ZN(n11008) );
  INV_X1 U6697 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n10050) );
  AOI21_X1 U6698 ( .B1(n8175), .B2(n7072), .A(n6957), .ZN(n8169) );
  OR2_X1 U6699 ( .A1(n8851), .A2(n7114), .ZN(n11012) );
  INV_X1 U6700 ( .A(n8765), .ZN(n7886) );
  OR2_X1 U6701 ( .A1(n10375), .A2(n6301), .ZN(n6197) );
  INV_X1 U6702 ( .A(n10851), .ZN(n10794) );
  INV_X1 U6703 ( .A(n10829), .ZN(n10858) );
  INV_X1 U6704 ( .A(n10847), .ZN(n10822) );
  AND2_X1 U6705 ( .A1(n8825), .A2(n8822), .ZN(n10389) );
  INV_X1 U6706 ( .A(n8353), .ZN(n10507) );
  INV_X1 U6707 ( .A(n11021), .ZN(n10520) );
  INV_X1 U6708 ( .A(n10504), .ZN(n11023) );
  AND2_X1 U6709 ( .A1(n11116), .A2(n10996), .ZN(n8211) );
  AND2_X1 U6710 ( .A1(n11120), .A2(n10996), .ZN(n8213) );
  INV_X1 U6711 ( .A(n11000), .ZN(n11113) );
  NAND2_X1 U6712 ( .A1(n6840), .A2(n6839), .ZN(n7365) );
  AND2_X1 U6713 ( .A1(n7371), .A2(n7370), .ZN(n9082) );
  OR3_X1 U6714 ( .A1(n7367), .A2(n7361), .A3(n7358), .ZN(n9061) );
  AND4_X1 U6715 ( .A1(n9096), .A2(n6787), .A3(n6786), .A4(n6785), .ZN(n9106)
         );
  INV_X1 U6716 ( .A(n9230), .ZN(n9947) );
  INV_X1 U6717 ( .A(n7896), .ZN(n9329) );
  INV_X1 U6718 ( .A(n10906), .ZN(n10904) );
  INV_X1 U6719 ( .A(n9429), .ZN(n10915) );
  OR2_X1 U6720 ( .A1(n7318), .A2(n9412), .ZN(n10918) );
  AND2_X1 U6721 ( .A1(n9979), .A2(n9978), .ZN(n10030) );
  INV_X1 U6722 ( .A(n10981), .ZN(n11046) );
  NAND2_X1 U6723 ( .A1(n10941), .A2(n10950), .ZN(n11048) );
  INV_X1 U6724 ( .A(n11048), .ZN(n10981) );
  AND2_X1 U6725 ( .A1(n7148), .A2(n7147), .ZN(n11154) );
  NAND2_X1 U6726 ( .A1(n6822), .A2(n7192), .ZN(n7256) );
  AND2_X1 U6727 ( .A1(n8266), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7259) );
  INV_X1 U6728 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8268) );
  INV_X1 U6729 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7651) );
  AND2_X1 U6730 ( .A1(n7107), .A2(n7289), .ZN(n11101) );
  AND2_X1 U6731 ( .A1(n7115), .A2(n11012), .ZN(n10183) );
  NAND2_X1 U6732 ( .A1(n6197), .A2(n6196), .ZN(n10391) );
  OR2_X1 U6733 ( .A1(n6004), .A2(n6003), .ZN(n10203) );
  INV_X1 U6734 ( .A(n10754), .ZN(n10862) );
  OR2_X1 U6735 ( .A1(n10529), .A2(n7578), .ZN(n8368) );
  INV_X1 U6736 ( .A(n8211), .ZN(n10592) );
  INV_X1 U6737 ( .A(n11116), .ZN(n11115) );
  INV_X1 U6738 ( .A(n10320), .ZN(n10624) );
  INV_X1 U6739 ( .A(n8213), .ZN(n10651) );
  INV_X1 U6740 ( .A(n11120), .ZN(n11117) );
  AND2_X1 U6741 ( .A1(n8479), .A2(n6340), .ZN(n7189) );
  INV_X1 U6742 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9764) );
  INV_X1 U6743 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9788) );
  INV_X1 U6744 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9591) );
  NOR2_X2 U6745 ( .A1(n7365), .A2(n7151), .ZN(P2_U3893) );
  INV_X1 U6746 ( .A(n10215), .ZN(P1_U3973) );
  NAND2_X1 U6747 ( .A1(n6353), .A2(n6352), .ZN(P1_U3518) );
  NOR2_X2 U6748 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5718) );
  NOR2_X2 U6749 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5717) );
  NOR2_X2 U6750 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5716) );
  AND3_X2 U6751 ( .A1(n5718), .A2(n5717), .A3(n5716), .ZN(n5949) );
  NOR2_X1 U6752 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5719) );
  NOR2_X2 U6753 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5773) );
  AND2_X2 U6754 ( .A1(n5719), .A2(n5773), .ZN(n5802) );
  NAND3_X1 U6755 ( .A1(n5949), .A2(n5802), .A3(n5722), .ZN(n5971) );
  INV_X2 U6756 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9627) );
  INV_X2 U6757 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6343) );
  NOR2_X1 U6758 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5729) );
  NOR2_X1 U6759 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5728) );
  NOR2_X1 U6760 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5727) );
  NAND4_X1 U6761 ( .A1(n5706), .A2(n5729), .A3(n5728), .A4(n5727), .ZN(n5730)
         );
  NAND2_X1 U6762 ( .A1(n5732), .A2(n5733), .ZN(n10657) );
  INV_X1 U6763 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10658) );
  INV_X1 U6764 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5735) );
  INV_X1 U6765 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10749) );
  INV_X1 U6766 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U6767 ( .A1(n5738), .A2(n5736), .ZN(n5903) );
  INV_X1 U6768 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10750) );
  OR2_X1 U6769 ( .A1(n5903), .A2(n10750), .ZN(n5739) );
  INV_X8 U6770 ( .A(n7155), .ZN(n7159) );
  NAND2_X1 U6771 ( .A1(n7159), .A2(SI_0_), .ZN(n5741) );
  XNOR2_X1 U6772 ( .A(n5741), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10666) );
  NAND2_X1 U6773 ( .A1(n5742), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5744) );
  MUX2_X1 U6774 ( .A(n10752), .B(n10666), .S(n5777), .Z(n10932) );
  INV_X1 U6775 ( .A(n10932), .ZN(n7570) );
  NAND2_X1 U6776 ( .A1(n5807), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5753) );
  INV_X1 U6777 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5747) );
  OR2_X1 U6778 ( .A1(n6017), .A2(n5747), .ZN(n5752) );
  INV_X1 U6779 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5748) );
  OR2_X1 U6780 ( .A1(n6301), .A2(n5748), .ZN(n5751) );
  INV_X1 U6781 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5749) );
  OR2_X1 U6782 ( .A1(n5903), .A2(n5749), .ZN(n5750) );
  INV_X1 U6783 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U6784 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n10752), .ZN(n5754) );
  XNOR2_X1 U6785 ( .A(n5755), .B(n5754), .ZN(n7231) );
  NAND2_X2 U6786 ( .A1(n5777), .A2(n7159), .ZN(n5857) );
  INV_X1 U6787 ( .A(SI_1_), .ZN(n5756) );
  NAND3_X1 U6788 ( .A1(n5785), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n5758) );
  AND2_X1 U6789 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6790 ( .A1(n5758), .A2(n6406), .ZN(n5769) );
  XNOR2_X1 U6791 ( .A(n5768), .B(n5769), .ZN(n7168) );
  OR2_X1 U6792 ( .A1(n5857), .A2(n7168), .ZN(n5760) );
  OR2_X1 U6793 ( .A1(n10214), .A2(n5122), .ZN(n5761) );
  NAND2_X1 U6794 ( .A1(n7445), .A2(n5761), .ZN(n7299) );
  NAND2_X1 U6795 ( .A1(n8647), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5767) );
  INV_X1 U6796 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10234) );
  OR2_X1 U6797 ( .A1(n6301), .A2(n10234), .ZN(n5766) );
  INV_X1 U6798 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5762) );
  OR2_X1 U6799 ( .A1(n5903), .A2(n5762), .ZN(n5765) );
  INV_X1 U6800 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5763) );
  OR2_X1 U6801 ( .A1(n5789), .A2(n5763), .ZN(n5764) );
  NAND2_X1 U6802 ( .A1(n5769), .A2(n5768), .ZN(n5772) );
  NAND2_X1 U6803 ( .A1(n5770), .A2(SI_1_), .ZN(n5771) );
  NAND2_X1 U6804 ( .A1(n5772), .A2(n5771), .ZN(n5783) );
  MUX2_X1 U6805 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5785), .Z(n5784) );
  INV_X1 U6806 ( .A(SI_2_), .ZN(n9502) );
  XNOR2_X1 U6807 ( .A(n5784), .B(n9502), .ZN(n5782) );
  XNOR2_X1 U6808 ( .A(n5783), .B(n5782), .ZN(n7169) );
  INV_X1 U6809 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7170) );
  OR2_X1 U6810 ( .A1(n8777), .A2(n7170), .ZN(n5775) );
  OR2_X1 U6811 ( .A1(n5773), .A2(n5803), .ZN(n5779) );
  INV_X1 U6812 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5778) );
  XNOR2_X1 U6813 ( .A(n5779), .B(n5778), .ZN(n7230) );
  OR2_X1 U6814 ( .A1(n5777), .A2(n7230), .ZN(n5774) );
  NAND2_X1 U6815 ( .A1(n7299), .A2(n8786), .ZN(n7298) );
  OR2_X1 U6816 ( .A1(n10213), .A2(n7704), .ZN(n5776) );
  NAND2_X1 U6817 ( .A1(n7298), .A2(n5776), .ZN(n7460) );
  INV_X2 U6818 ( .A(n8777), .ZN(n6086) );
  INV_X2 U6819 ( .A(n5777), .ZN(n7194) );
  NAND2_X1 U6820 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  NAND2_X1 U6821 ( .A1(n5780), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5781) );
  XNOR2_X1 U6822 ( .A(n5781), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U6823 ( .A1(n6086), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n7194), .B2(
        n10250), .ZN(n5788) );
  NAND2_X1 U6824 ( .A1(n5783), .A2(n5782), .ZN(n5801) );
  NAND2_X1 U6825 ( .A1(n5784), .A2(SI_2_), .ZN(n5796) );
  NAND2_X1 U6826 ( .A1(n5801), .A2(n5796), .ZN(n5786) );
  INV_X1 U6827 ( .A(SI_3_), .ZN(n9709) );
  XNOR2_X1 U6828 ( .A(n5795), .B(n9709), .ZN(n5798) );
  XNOR2_X1 U6829 ( .A(n5786), .B(n5798), .ZN(n7161) );
  OR2_X1 U6830 ( .A1(n7161), .A2(n5857), .ZN(n5787) );
  NAND2_X1 U6831 ( .A1(n5788), .A2(n5787), .ZN(n7773) );
  INV_X1 U6832 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7234) );
  OR2_X1 U6833 ( .A1(n8649), .A2(n7234), .ZN(n5792) );
  OR2_X1 U6834 ( .A1(n6301), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5791) );
  INV_X1 U6835 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7216) );
  NAND4_X2 U6836 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n10212)
         );
  OR2_X1 U6837 ( .A1(n7489), .A2(n10212), .ZN(n8871) );
  AND2_X1 U6838 ( .A1(n10212), .A2(n7489), .ZN(n6289) );
  INV_X1 U6839 ( .A(n6289), .ZN(n8867) );
  NAND2_X1 U6840 ( .A1(n8871), .A2(n8867), .ZN(n7464) );
  NAND2_X1 U6841 ( .A1(n7460), .A2(n7464), .ZN(n7459) );
  OR2_X1 U6842 ( .A1(n10212), .A2(n7773), .ZN(n5794) );
  NAND2_X1 U6843 ( .A1(n7459), .A2(n5794), .ZN(n7588) );
  NAND2_X1 U6844 ( .A1(n5795), .A2(SI_3_), .ZN(n5797) );
  AND2_X1 U6845 ( .A1(n5796), .A2(n5797), .ZN(n5800) );
  INV_X1 U6846 ( .A(n5797), .ZN(n5799) );
  INV_X1 U6847 ( .A(SI_4_), .ZN(n9708) );
  XNOR2_X1 U6848 ( .A(n5820), .B(n9708), .ZN(n5818) );
  XNOR2_X1 U6849 ( .A(n5819), .B(n5818), .ZN(n7171) );
  OR2_X1 U6850 ( .A1(n7171), .A2(n5857), .ZN(n5806) );
  OR2_X1 U6851 ( .A1(n5802), .A2(n5803), .ZN(n5804) );
  XNOR2_X1 U6852 ( .A(n5804), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7236) );
  AOI22_X1 U6853 ( .A1(n6086), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n7194), .B2(
        n7236), .ZN(n5805) );
  NAND2_X1 U6854 ( .A1(n5806), .A2(n5805), .ZN(n10995) );
  NAND2_X1 U6855 ( .A1(n5807), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5815) );
  INV_X1 U6856 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5808) );
  OR2_X1 U6857 ( .A1(n6017), .A2(n5808), .ZN(n5814) );
  INV_X1 U6858 ( .A(n5830), .ZN(n5811) );
  INV_X1 U6859 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7774) );
  INV_X1 U6860 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U6861 ( .A1(n7774), .A2(n5809), .ZN(n5810) );
  NAND2_X1 U6862 ( .A1(n5811), .A2(n5810), .ZN(n7600) );
  OR2_X1 U6863 ( .A1(n6301), .A2(n7600), .ZN(n5813) );
  INV_X1 U6864 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7597) );
  OR2_X1 U6865 ( .A1(n8653), .A2(n7597), .ZN(n5812) );
  NOR2_X1 U6866 ( .A1(n10995), .A2(n10211), .ZN(n5817) );
  NAND2_X1 U6867 ( .A1(n10211), .A2(n10995), .ZN(n5816) );
  OAI21_X1 U6868 ( .B1(n7588), .B2(n5817), .A(n5816), .ZN(n7375) );
  NAND2_X1 U6869 ( .A1(n5819), .A2(n5818), .ZN(n5822) );
  NAND2_X1 U6870 ( .A1(n5820), .A2(SI_4_), .ZN(n5821) );
  NAND2_X1 U6871 ( .A1(n5822), .A2(n5821), .ZN(n5836) );
  MUX2_X1 U6872 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7159), .Z(n5837) );
  INV_X1 U6873 ( .A(SI_5_), .ZN(n9497) );
  XNOR2_X1 U6874 ( .A(n5837), .B(n9497), .ZN(n5835) );
  XNOR2_X1 U6875 ( .A(n5836), .B(n5835), .ZN(n7163) );
  OR2_X1 U6876 ( .A1(n7163), .A2(n5857), .ZN(n5828) );
  NAND2_X1 U6877 ( .A1(n5802), .A2(n5823), .ZN(n5825) );
  NAND2_X1 U6878 ( .A1(n5825), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5824) );
  MUX2_X1 U6879 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5824), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5826) );
  AND2_X1 U6880 ( .A1(n5826), .A2(n5951), .ZN(n10276) );
  AOI22_X1 U6881 ( .A1(n6086), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7194), .B2(
        n10276), .ZN(n5827) );
  NAND2_X1 U6882 ( .A1(n5828), .A2(n5827), .ZN(n11017) );
  NAND2_X1 U6883 ( .A1(n5807), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5834) );
  INV_X1 U6884 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5829) );
  OR2_X1 U6885 ( .A1(n6017), .A2(n5829), .ZN(n5833) );
  NAND2_X1 U6886 ( .A1(n5830), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5845) );
  OAI21_X1 U6887 ( .B1(n5830), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5845), .ZN(
        n11013) );
  OR2_X1 U6888 ( .A1(n6301), .A2(n11013), .ZN(n5832) );
  INV_X1 U6889 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11014) );
  OR2_X1 U6890 ( .A1(n8653), .A2(n11014), .ZN(n5831) );
  NAND4_X1 U6891 ( .A1(n5834), .A2(n5833), .A3(n5832), .A4(n5831), .ZN(n10210)
         );
  INV_X1 U6892 ( .A(n10210), .ZN(n7589) );
  OR2_X1 U6893 ( .A1(n11017), .A2(n7589), .ZN(n8873) );
  NAND2_X1 U6894 ( .A1(n11017), .A2(n7589), .ZN(n8672) );
  NAND2_X1 U6895 ( .A1(n8873), .A2(n8672), .ZN(n8788) );
  INV_X1 U6896 ( .A(n8788), .ZN(n8667) );
  OAI22_X1 U6897 ( .A1(n7375), .A2(n8667), .B1(n11017), .B2(n10210), .ZN(n7653) );
  NAND2_X1 U6898 ( .A1(n5836), .A2(n5835), .ZN(n5839) );
  NAND2_X1 U6899 ( .A1(n5837), .A2(SI_5_), .ZN(n5838) );
  MUX2_X1 U6900 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7159), .Z(n5855) );
  INV_X1 U6901 ( .A(SI_6_), .ZN(n9493) );
  XNOR2_X1 U6902 ( .A(n5855), .B(n9493), .ZN(n5853) );
  XNOR2_X1 U6903 ( .A(n5854), .B(n5853), .ZN(n7166) );
  OR2_X1 U6904 ( .A1(n7166), .A2(n5857), .ZN(n5842) );
  NAND2_X1 U6905 ( .A1(n5951), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U6906 ( .A(n5840), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U6907 ( .A1(n6086), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7194), .B2(
        n10289), .ZN(n5841) );
  NAND2_X1 U6908 ( .A1(n5842), .A2(n5841), .ZN(n10166) );
  NAND2_X1 U6909 ( .A1(n5807), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5851) );
  INV_X1 U6910 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5843) );
  OR2_X1 U6911 ( .A1(n6017), .A2(n5843), .ZN(n5850) );
  AND2_X1 U6912 ( .A1(n5845), .A2(n5844), .ZN(n5846) );
  OR2_X1 U6913 ( .A1(n5846), .A2(n5861), .ZN(n10168) );
  OR2_X1 U6914 ( .A1(n6301), .A2(n10168), .ZN(n5849) );
  INV_X1 U6915 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5847) );
  OR2_X1 U6916 ( .A1(n8653), .A2(n5847), .ZN(n5848) );
  NAND4_X1 U6917 ( .A1(n5851), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(n10209)
         );
  OR2_X1 U6918 ( .A1(n10166), .A2(n7751), .ZN(n8676) );
  NAND2_X1 U6919 ( .A1(n10166), .A2(n7751), .ZN(n8790) );
  INV_X1 U6920 ( .A(n8674), .ZN(n7652) );
  NAND2_X1 U6921 ( .A1(n7653), .A2(n7652), .ZN(n7655) );
  OR2_X1 U6922 ( .A1(n10166), .A2(n10209), .ZN(n5852) );
  NAND2_X1 U6923 ( .A1(n7655), .A2(n5852), .ZN(n7745) );
  NAND2_X1 U6924 ( .A1(n5855), .A2(SI_6_), .ZN(n5856) );
  MUX2_X1 U6925 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7159), .Z(n5873) );
  XNOR2_X1 U6926 ( .A(n5873), .B(SI_7_), .ZN(n5870) );
  XNOR2_X1 U6927 ( .A(n5872), .B(n5870), .ZN(n7172) );
  NAND2_X1 U6928 ( .A1(n7172), .A2(n5948), .ZN(n5860) );
  NOR2_X1 U6929 ( .A1(n5951), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5879) );
  OR2_X1 U6930 ( .A1(n5879), .A2(n5803), .ZN(n5858) );
  XNOR2_X1 U6931 ( .A(n5858), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U6932 ( .A1(n6086), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7194), .B2(
        n10302), .ZN(n5859) );
  NAND2_X1 U6933 ( .A1(n5860), .A2(n5859), .ZN(n7784) );
  NAND2_X1 U6934 ( .A1(n8647), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5867) );
  INV_X1 U6935 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7221) );
  OR2_X1 U6936 ( .A1(n5903), .A2(n7221), .ZN(n5866) );
  NAND2_X1 U6937 ( .A1(n5861), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5885) );
  OR2_X1 U6938 ( .A1(n5861), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U6939 ( .A1(n5885), .A2(n5862), .ZN(n7671) );
  OR2_X1 U6940 ( .A1(n6301), .A2(n7671), .ZN(n5865) );
  INV_X1 U6941 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5863) );
  OR2_X1 U6942 ( .A1(n8649), .A2(n5863), .ZN(n5864) );
  NAND4_X1 U6943 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n10208)
         );
  INV_X1 U6944 ( .A(n10208), .ZN(n5868) );
  OR2_X1 U6945 ( .A1(n7784), .A2(n5868), .ZN(n8683) );
  NAND2_X1 U6946 ( .A1(n7784), .A2(n5868), .ZN(n7797) );
  NAND2_X1 U6947 ( .A1(n8683), .A2(n7797), .ZN(n8680) );
  OR2_X1 U6948 ( .A1(n7784), .A2(n10208), .ZN(n5869) );
  INV_X1 U6949 ( .A(n5870), .ZN(n5871) );
  NAND2_X1 U6950 ( .A1(n5873), .A2(SI_7_), .ZN(n5874) );
  INV_X1 U6951 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7177) );
  INV_X1 U6952 ( .A(SI_8_), .ZN(n9700) );
  NAND2_X1 U6953 ( .A1(n5875), .A2(n9700), .ZN(n5893) );
  INV_X1 U6954 ( .A(n5875), .ZN(n5876) );
  NAND2_X1 U6955 ( .A1(n5876), .A2(SI_8_), .ZN(n5877) );
  NAND2_X1 U6956 ( .A1(n5893), .A2(n5877), .ZN(n5891) );
  XNOR2_X1 U6957 ( .A(n5892), .B(n5891), .ZN(n7176) );
  NAND2_X1 U6958 ( .A1(n7176), .A2(n5948), .ZN(n5882) );
  INV_X1 U6959 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U6960 ( .A1(n5879), .A2(n5878), .ZN(n5898) );
  NAND2_X1 U6961 ( .A1(n5898), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5880) );
  XNOR2_X1 U6962 ( .A(n5880), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7242) );
  AOI22_X1 U6963 ( .A1(n6086), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7194), .B2(
        n7242), .ZN(n5881) );
  NAND2_X1 U6964 ( .A1(n8647), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5890) );
  INV_X1 U6965 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5883) );
  OR2_X1 U6966 ( .A1(n8649), .A2(n5883), .ZN(n5889) );
  NAND2_X1 U6967 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  NAND2_X1 U6968 ( .A1(n5904), .A2(n5886), .ZN(n7862) );
  OR2_X1 U6969 ( .A1(n6301), .A2(n7862), .ZN(n5888) );
  INV_X1 U6970 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7804) );
  OR2_X1 U6971 ( .A1(n8653), .A2(n7804), .ZN(n5887) );
  NAND4_X1 U6972 ( .A1(n5890), .A2(n5889), .A3(n5888), .A4(n5887), .ZN(n10207)
         );
  INV_X1 U6973 ( .A(n10207), .ZN(n7752) );
  NAND2_X1 U6974 ( .A1(n7866), .A2(n7752), .ZN(n6280) );
  NAND2_X1 U6975 ( .A1(n7840), .A2(n6280), .ZN(n8687) );
  INV_X1 U6976 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7198) );
  MUX2_X1 U6977 ( .A(n7198), .B(n9591), .S(n7159), .Z(n5895) );
  NAND2_X1 U6978 ( .A1(n5895), .A2(n9699), .ZN(n5912) );
  INV_X1 U6979 ( .A(n5895), .ZN(n5896) );
  NAND2_X1 U6980 ( .A1(n5896), .A2(SI_9_), .ZN(n5897) );
  NAND2_X1 U6981 ( .A1(n5913), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5899) );
  XNOR2_X1 U6982 ( .A(n5899), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7271) );
  AOI22_X1 U6983 ( .A1(n6086), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7194), .B2(
        n7271), .ZN(n5900) );
  NAND2_X1 U6984 ( .A1(n8647), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5910) );
  INV_X1 U6985 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5902) );
  OR2_X1 U6986 ( .A1(n5903), .A2(n5902), .ZN(n5909) );
  AND2_X1 U6987 ( .A1(n5904), .A2(n7247), .ZN(n5905) );
  OR2_X1 U6988 ( .A1(n5905), .A2(n5917), .ZN(n7940) );
  OR2_X1 U6989 ( .A1(n6301), .A2(n7940), .ZN(n5908) );
  INV_X1 U6990 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5906) );
  OR2_X1 U6991 ( .A1(n8649), .A2(n5906), .ZN(n5907) );
  NAND4_X1 U6992 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n10206)
         );
  INV_X1 U6993 ( .A(n10206), .ZN(n7863) );
  OR2_X1 U6994 ( .A1(n7946), .A2(n7863), .ZN(n8701) );
  NAND2_X1 U6995 ( .A1(n7946), .A2(n7863), .ZN(n8694) );
  NAND2_X1 U6996 ( .A1(n8701), .A2(n8694), .ZN(n7847) );
  NAND2_X1 U6997 ( .A1(n7848), .A2(n7847), .ZN(n7846) );
  OR2_X1 U6998 ( .A1(n7946), .A2(n10206), .ZN(n5911) );
  MUX2_X1 U6999 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7159), .Z(n5924) );
  XNOR2_X1 U7000 ( .A(n5924), .B(n9698), .ZN(n5923) );
  XNOR2_X1 U7001 ( .A(n5925), .B(n5923), .ZN(n7200) );
  NAND2_X1 U7002 ( .A1(n7200), .A2(n5948), .ZN(n5915) );
  OAI21_X1 U7003 ( .B1(n5913), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U7004 ( .A(n5930), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U7005 ( .A1(n6086), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10857), 
        .B2(n7194), .ZN(n5914) );
  NAND2_X1 U7006 ( .A1(n5807), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5922) );
  INV_X1 U7007 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5916) );
  OR2_X1 U7008 ( .A1(n6017), .A2(n5916), .ZN(n5921) );
  NOR2_X1 U7009 ( .A1(n5917), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5918) );
  OR2_X1 U7010 ( .A1(n5935), .A2(n5918), .ZN(n8171) );
  OR2_X1 U7011 ( .A1(n6301), .A2(n8171), .ZN(n5920) );
  INV_X1 U7012 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7830) );
  OR2_X1 U7013 ( .A1(n8653), .A2(n7830), .ZN(n5919) );
  NAND4_X1 U7014 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n5919), .ZN(n7916)
         );
  OR2_X1 U7015 ( .A1(n8175), .A2(n11095), .ZN(n8878) );
  NAND2_X1 U7016 ( .A1(n8175), .A2(n11095), .ZN(n8698) );
  NAND2_X1 U7017 ( .A1(n8878), .A2(n8698), .ZN(n8794) );
  MUX2_X1 U7018 ( .A(n7255), .B(n9805), .S(n7159), .Z(n5926) );
  NAND2_X1 U7019 ( .A1(n5926), .A2(n9694), .ZN(n5945) );
  INV_X1 U7020 ( .A(n5926), .ZN(n5927) );
  NAND2_X1 U7021 ( .A1(n5927), .A2(SI_11_), .ZN(n5928) );
  NAND2_X1 U7022 ( .A1(n5945), .A2(n5928), .ZN(n5946) );
  XNOR2_X1 U7023 ( .A(n5947), .B(n5946), .ZN(n7212) );
  NAND2_X1 U7024 ( .A1(n7212), .A2(n5948), .ZN(n5934) );
  INV_X1 U7025 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7026 ( .A1(n5930), .A2(n5929), .ZN(n5931) );
  NAND2_X1 U7027 ( .A1(n5931), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5932) );
  XNOR2_X1 U7028 ( .A(n5932), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U7029 ( .A1(n10773), .A2(n7194), .B1(n6086), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7030 ( .A1(n8647), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5942) );
  INV_X1 U7031 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7272) );
  OR2_X1 U7032 ( .A1(n8649), .A2(n7272), .ZN(n5941) );
  INV_X1 U7033 ( .A(n5935), .ZN(n5937) );
  INV_X1 U7034 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7035 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  NAND2_X1 U7036 ( .A1(n5957), .A2(n5938), .ZN(n11100) );
  OR2_X1 U7037 ( .A1(n6301), .A2(n11100), .ZN(n5940) );
  INV_X1 U7038 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7921) );
  OR2_X1 U7039 ( .A1(n8653), .A2(n7921), .ZN(n5939) );
  NAND4_X1 U7040 ( .A1(n5942), .A2(n5941), .A3(n5940), .A4(n5939), .ZN(n10205)
         );
  OR2_X1 U7041 ( .A1(n11089), .A2(n10205), .ZN(n5943) );
  MUX2_X1 U7042 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7159), .Z(n5967) );
  XNOR2_X1 U7043 ( .A(n5967), .B(n9693), .ZN(n5966) );
  XNOR2_X1 U7044 ( .A(n5970), .B(n5966), .ZN(n7260) );
  NAND2_X1 U7045 ( .A1(n7260), .A2(n5948), .ZN(n5954) );
  INV_X1 U7046 ( .A(n5949), .ZN(n5950) );
  OAI21_X1 U7047 ( .B1(n5951), .B2(n5950), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5952) );
  XNOR2_X1 U7048 ( .A(n5952), .B(P1_IR_REG_12__SCAN_IN), .ZN(n8026) );
  AOI22_X1 U7049 ( .A1(n6086), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7194), .B2(
        n8026), .ZN(n5953) );
  NAND2_X1 U7050 ( .A1(n8647), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5963) );
  INV_X1 U7051 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5955) );
  OR2_X1 U7052 ( .A1(n8653), .A2(n5955), .ZN(n5962) );
  NAND2_X1 U7053 ( .A1(n5957), .A2(n5956), .ZN(n5958) );
  NAND2_X1 U7054 ( .A1(n5976), .A2(n5958), .ZN(n8274) );
  OR2_X1 U7055 ( .A1(n6301), .A2(n8274), .ZN(n5961) );
  INV_X1 U7056 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7057 ( .A1(n8649), .A2(n5959), .ZN(n5960) );
  NAND4_X1 U7058 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(n11090)
         );
  NOR2_X1 U7059 ( .A1(n7956), .A2(n11090), .ZN(n5965) );
  NAND2_X1 U7060 ( .A1(n7956), .A2(n11090), .ZN(n5964) );
  INV_X1 U7061 ( .A(n5966), .ZN(n5969) );
  NAND2_X1 U7062 ( .A1(n5967), .A2(SI_12_), .ZN(n5968) );
  MUX2_X1 U7063 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7159), .Z(n5988) );
  XNOR2_X1 U7064 ( .A(n5988), .B(SI_13_), .ZN(n5985) );
  XNOR2_X1 U7065 ( .A(n5987), .B(n5985), .ZN(n7282) );
  NAND2_X1 U7066 ( .A1(n7282), .A2(n5948), .ZN(n5975) );
  NAND2_X1 U7067 ( .A1(n5972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5973) );
  XNOR2_X1 U7068 ( .A(n5973), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U7069 ( .A1(n6086), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7194), .B2(
        n10842), .ZN(n5974) );
  NAND2_X1 U7070 ( .A1(n5807), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7071 ( .A1(n5976), .A2(n8301), .ZN(n5977) );
  NAND2_X1 U7072 ( .A1(n5996), .A2(n5977), .ZN(n8302) );
  OR2_X1 U7073 ( .A1(n8302), .A2(n6301), .ZN(n5981) );
  INV_X1 U7074 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5978) );
  OR2_X1 U7075 ( .A1(n6017), .A2(n5978), .ZN(n5980) );
  INV_X1 U7076 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8148) );
  OR2_X1 U7077 ( .A1(n8653), .A2(n8148), .ZN(n5979) );
  NAND4_X1 U7078 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n10204)
         );
  AND2_X1 U7079 ( .A1(n8214), .A2(n10204), .ZN(n5984) );
  OR2_X1 U7080 ( .A1(n8214), .A2(n10204), .ZN(n5983) );
  INV_X1 U7081 ( .A(n5985), .ZN(n5986) );
  NAND2_X1 U7082 ( .A1(n5989), .A2(n9689), .ZN(n6007) );
  INV_X1 U7083 ( .A(n5989), .ZN(n5990) );
  NAND2_X1 U7084 ( .A1(n5990), .A2(SI_14_), .ZN(n5991) );
  NAND2_X1 U7085 ( .A1(n6007), .A2(n5991), .ZN(n6005) );
  XNOR2_X1 U7086 ( .A(n6006), .B(n6005), .ZN(n7295) );
  NAND2_X1 U7087 ( .A1(n7295), .A2(n5948), .ZN(n5994) );
  OR2_X1 U7088 ( .A1(n5972), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7089 ( .A1(n6009), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U7090 ( .A(n5992), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U7091 ( .A1(n6086), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7194), .B2(
        n10789), .ZN(n5993) );
  NAND2_X2 U7092 ( .A1(n5994), .A2(n5993), .ZN(n10612) );
  INV_X1 U7093 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7094 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  NAND2_X1 U7095 ( .A1(n6014), .A2(n5997), .ZN(n8393) );
  INV_X1 U7096 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5998) );
  OR2_X1 U7097 ( .A1(n8653), .A2(n5998), .ZN(n5999) );
  OAI21_X1 U7098 ( .B1(n8393), .B2(n6301), .A(n5999), .ZN(n6004) );
  INV_X1 U7099 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6002) );
  INV_X1 U7100 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6000) );
  OR2_X1 U7101 ( .A1(n6017), .A2(n6000), .ZN(n6001) );
  OAI21_X1 U7102 ( .B1(n8649), .B2(n6002), .A(n6001), .ZN(n6003) );
  INV_X1 U7103 ( .A(n10203), .ZN(n8303) );
  AND2_X1 U7104 ( .A1(n10612), .A2(n8303), .ZN(n8717) );
  INV_X1 U7105 ( .A(n8717), .ZN(n8664) );
  MUX2_X1 U7106 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7159), .Z(n6026) );
  XNOR2_X1 U7107 ( .A(n6026), .B(n9656), .ZN(n6023) );
  XNOR2_X1 U7108 ( .A(n6025), .B(n6023), .ZN(n7388) );
  NAND2_X1 U7109 ( .A1(n7388), .A2(n5948), .ZN(n6012) );
  NOR2_X1 U7110 ( .A1(n6009), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6032) );
  OR2_X1 U7111 ( .A1(n6032), .A2(n5803), .ZN(n6010) );
  XNOR2_X1 U7112 ( .A(n6010), .B(n6031), .ZN(n8029) );
  INV_X1 U7113 ( .A(n8029), .ZN(n10814) );
  AOI22_X1 U7114 ( .A1(n6086), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7194), .B2(
        n10814), .ZN(n6011) );
  INV_X1 U7115 ( .A(n6014), .ZN(n6013) );
  INV_X1 U7116 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U7117 ( .A1(n6014), .A2(n10192), .ZN(n6015) );
  NAND2_X1 U7118 ( .A1(n6036), .A2(n6015), .ZN(n10188) );
  OR2_X1 U7119 ( .A1(n10188), .A2(n6301), .ZN(n6021) );
  INV_X1 U7120 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10807) );
  OR2_X1 U7121 ( .A1(n8649), .A2(n10807), .ZN(n6019) );
  INV_X1 U7122 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7123 ( .A1(n6017), .A2(n6016), .ZN(n6018) );
  AND2_X1 U7124 ( .A1(n6019), .A2(n6018), .ZN(n6020) );
  OAI211_X1 U7125 ( .C1(n8653), .C2(n10810), .A(n6021), .B(n6020), .ZN(n10202)
         );
  INV_X1 U7126 ( .A(n10202), .ZN(n8355) );
  NOR2_X1 U7127 ( .A1(n10197), .A2(n8355), .ZN(n8720) );
  INV_X1 U7128 ( .A(n8720), .ZN(n8379) );
  NAND2_X1 U7129 ( .A1(n10197), .A2(n8355), .ZN(n8724) );
  NAND2_X1 U7130 ( .A1(n8379), .A2(n8724), .ZN(n8802) );
  NAND2_X1 U7131 ( .A1(n8318), .A2(n8802), .ZN(n8320) );
  NAND2_X1 U7132 ( .A1(n10197), .A2(n10202), .ZN(n6022) );
  INV_X1 U7133 ( .A(n6023), .ZN(n6024) );
  NAND2_X1 U7134 ( .A1(n6026), .A2(SI_15_), .ZN(n6027) );
  NAND2_X1 U7135 ( .A1(n6028), .A2(n9652), .ZN(n6040) );
  INV_X1 U7136 ( .A(n6028), .ZN(n6029) );
  NAND2_X1 U7137 ( .A1(n6029), .A2(SI_16_), .ZN(n6030) );
  NAND2_X1 U7138 ( .A1(n6040), .A2(n6030), .ZN(n6041) );
  NAND2_X1 U7139 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  NAND2_X1 U7140 ( .A1(n6033), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6034) );
  XNOR2_X1 U7141 ( .A(n6034), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8120) );
  AOI22_X1 U7142 ( .A1(n6086), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7194), .B2(
        n8120), .ZN(n6035) );
  NAND2_X1 U7143 ( .A1(n6036), .A2(n8022), .ZN(n6037) );
  NAND2_X1 U7144 ( .A1(n6049), .A2(n6037), .ZN(n10101) );
  AOI22_X1 U7145 ( .A1(n6065), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8647), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n6039) );
  INV_X1 U7146 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8019) );
  OR2_X1 U7147 ( .A1(n8649), .A2(n8019), .ZN(n6038) );
  OAI211_X1 U7148 ( .C1(n10101), .C2(n6301), .A(n6039), .B(n6038), .ZN(n10508)
         );
  INV_X1 U7149 ( .A(n10508), .ZN(n10195) );
  OR2_X1 U7150 ( .A1(n10598), .A2(n10195), .ZN(n8725) );
  NAND2_X1 U7151 ( .A1(n8725), .A2(n8726), .ZN(n8803) );
  MUX2_X1 U7152 ( .A(n7651), .B(n9793), .S(n7159), .Z(n6043) );
  NAND2_X1 U7153 ( .A1(n6043), .A2(n9478), .ZN(n6056) );
  INV_X1 U7154 ( .A(n6043), .ZN(n6044) );
  NAND2_X1 U7155 ( .A1(n6044), .A2(SI_17_), .ZN(n6045) );
  XNOR2_X1 U7156 ( .A(n6055), .B(n6054), .ZN(n7649) );
  NAND2_X1 U7157 ( .A1(n7649), .A2(n5948), .ZN(n6047) );
  NAND2_X1 U7158 ( .A1(n6266), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6058) );
  XNOR2_X1 U7159 ( .A(n6058), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8249) );
  AOI22_X1 U7160 ( .A1(n6086), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7194), .B2(
        n8249), .ZN(n6046) );
  INV_X1 U7161 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8117) );
  INV_X1 U7162 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7163 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  NAND2_X1 U7164 ( .A1(n6063), .A2(n6050), .ZN(n10113) );
  OR2_X1 U7165 ( .A1(n10113), .A2(n6301), .ZN(n6052) );
  AOI22_X1 U7166 ( .A1(n5807), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n8647), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n6051) );
  OAI211_X1 U7167 ( .C1(n8653), .C2(n8117), .A(n6052), .B(n6051), .ZN(n10492)
         );
  XNOR2_X1 U7168 ( .A(n10594), .B(n10492), .ZN(n8804) );
  NAND2_X1 U7169 ( .A1(n10594), .A2(n10492), .ZN(n6053) );
  NAND2_X1 U7170 ( .A1(n10513), .A2(n6053), .ZN(n10486) );
  NAND2_X1 U7171 ( .A1(n6055), .A2(n6054), .ZN(n6057) );
  MUX2_X1 U7172 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7159), .Z(n6076) );
  XNOR2_X1 U7173 ( .A(n6076), .B(n9655), .ZN(n6075) );
  XNOR2_X1 U7174 ( .A(n6079), .B(n6075), .ZN(n7741) );
  NAND2_X1 U7175 ( .A1(n7741), .A2(n5948), .ZN(n6061) );
  NAND2_X1 U7176 ( .A1(n6058), .A2(n6262), .ZN(n6059) );
  NAND2_X1 U7177 ( .A1(n6059), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6083) );
  XNOR2_X1 U7178 ( .A(n6083), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8253) );
  AOI22_X1 U7179 ( .A1(n6086), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7194), .B2(
        n8253), .ZN(n6060) );
  NAND2_X1 U7180 ( .A1(n6063), .A2(n6062), .ZN(n6064) );
  AND2_X1 U7181 ( .A1(n6091), .A2(n6064), .ZN(n10499) );
  NAND2_X1 U7182 ( .A1(n10499), .A2(n6235), .ZN(n6071) );
  INV_X1 U7183 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7184 ( .A1(n5807), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7185 ( .A1(n8647), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6066) );
  OAI211_X1 U7186 ( .C1(n6068), .C2(n6305), .A(n6067), .B(n6066), .ZN(n6069)
         );
  INV_X1 U7187 ( .A(n6069), .ZN(n6070) );
  NAND2_X1 U7188 ( .A1(n6071), .A2(n6070), .ZN(n10510) );
  OR2_X1 U7189 ( .A1(n10498), .A2(n10510), .ZN(n6072) );
  NAND2_X1 U7190 ( .A1(n10498), .A2(n10510), .ZN(n6073) );
  INV_X1 U7191 ( .A(n6075), .ZN(n6078) );
  NAND2_X1 U7192 ( .A1(n6076), .A2(SI_18_), .ZN(n6077) );
  OAI21_X2 U7193 ( .B1(n6079), .B2(n6078), .A(n6077), .ZN(n6101) );
  NAND2_X1 U7194 ( .A1(n6080), .A2(n9474), .ZN(n6099) );
  INV_X1 U7195 ( .A(n6080), .ZN(n6081) );
  NAND2_X1 U7196 ( .A1(n6081), .A2(SI_19_), .ZN(n6082) );
  NAND2_X1 U7197 ( .A1(n6099), .A2(n6082), .ZN(n6100) );
  XNOR2_X1 U7198 ( .A(n6101), .B(n6100), .ZN(n7911) );
  NAND2_X1 U7199 ( .A1(n7911), .A2(n5948), .ZN(n6088) );
  NAND2_X1 U7200 ( .A1(n6083), .A2(n6263), .ZN(n6084) );
  NAND2_X1 U7201 ( .A1(n6084), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6085) );
  AOI22_X1 U7202 ( .A1(n6086), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8923), .B2(
        n7194), .ZN(n6087) );
  INV_X1 U7203 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7204 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  NAND2_X1 U7205 ( .A1(n6108), .A2(n6092), .ZN(n10070) );
  OR2_X1 U7206 ( .A1(n10070), .A2(n6301), .ZN(n6098) );
  INV_X1 U7207 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7208 ( .A1(n5807), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7209 ( .A1(n8647), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6093) );
  OAI211_X1 U7210 ( .C1(n6095), .C2(n6305), .A(n6094), .B(n6093), .ZN(n6096)
         );
  INV_X1 U7211 ( .A(n6096), .ZN(n6097) );
  NAND2_X1 U7212 ( .A1(n6098), .A2(n6097), .ZN(n10493) );
  INV_X1 U7213 ( .A(n10493), .ZN(n10157) );
  OR2_X1 U7214 ( .A1(n10479), .A2(n10157), .ZN(n8730) );
  NAND2_X1 U7215 ( .A1(n10479), .A2(n10157), .ZN(n8899) );
  NAND2_X1 U7216 ( .A1(n8730), .A2(n8899), .ZN(n8733) );
  MUX2_X1 U7217 ( .A(n8014), .B(n9788), .S(n7159), .Z(n6102) );
  INV_X1 U7218 ( .A(SI_20_), .ZN(n9675) );
  NAND2_X1 U7219 ( .A1(n6102), .A2(n9675), .ZN(n6118) );
  INV_X1 U7220 ( .A(n6102), .ZN(n6103) );
  NAND2_X1 U7221 ( .A1(n6103), .A2(SI_20_), .ZN(n6104) );
  XNOR2_X1 U7222 ( .A(n6117), .B(n6116), .ZN(n8013) );
  NAND2_X1 U7223 ( .A1(n8013), .A2(n5948), .ZN(n6106) );
  OR2_X1 U7224 ( .A1(n8777), .A2(n9788), .ZN(n6105) );
  INV_X1 U7225 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7226 ( .A1(n6108), .A2(n6107), .ZN(n6109) );
  AND2_X1 U7227 ( .A1(n6122), .A2(n6109), .ZN(n10459) );
  NAND2_X1 U7228 ( .A1(n10459), .A2(n6235), .ZN(n6115) );
  INV_X1 U7229 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7230 ( .A1(n5807), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7231 ( .A1(n8647), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6110) );
  OAI211_X1 U7232 ( .C1(n6112), .C2(n6305), .A(n6111), .B(n6110), .ZN(n6113)
         );
  INV_X1 U7233 ( .A(n6113), .ZN(n6114) );
  NAND2_X1 U7234 ( .A1(n6115), .A2(n6114), .ZN(n10474) );
  INV_X1 U7235 ( .A(n10474), .ZN(n10081) );
  NAND2_X1 U7236 ( .A1(n10578), .A2(n10081), .ZN(n10438) );
  MUX2_X1 U7237 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7159), .Z(n6132) );
  XNOR2_X1 U7238 ( .A(n6132), .B(n9467), .ZN(n6131) );
  XNOR2_X1 U7239 ( .A(n6130), .B(n6131), .ZN(n8179) );
  NAND2_X1 U7240 ( .A1(n8179), .A2(n5948), .ZN(n6120) );
  INV_X1 U7241 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8180) );
  OR2_X1 U7242 ( .A1(n8777), .A2(n8180), .ZN(n6119) );
  INV_X1 U7243 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7244 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  NAND2_X1 U7245 ( .A1(n6138), .A2(n6123), .ZN(n10450) );
  OR2_X1 U7246 ( .A1(n10450), .A2(n6301), .ZN(n6128) );
  INV_X1 U7247 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n10451) );
  NAND2_X1 U7248 ( .A1(n5807), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7249 ( .A1(n8647), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6124) );
  OAI211_X1 U7250 ( .C1(n10451), .C2(n6305), .A(n6125), .B(n6124), .ZN(n6126)
         );
  INV_X1 U7251 ( .A(n6126), .ZN(n6127) );
  NAND2_X1 U7252 ( .A1(n6128), .A2(n6127), .ZN(n10464) );
  INV_X1 U7253 ( .A(n10464), .ZN(n10146) );
  NOR2_X1 U7254 ( .A1(n10572), .A2(n10146), .ZN(n8742) );
  INV_X1 U7255 ( .A(n8742), .ZN(n8903) );
  AND2_X1 U7256 ( .A1(n10572), .A2(n10146), .ZN(n8743) );
  INV_X1 U7257 ( .A(n8743), .ZN(n6278) );
  NAND2_X1 U7258 ( .A1(n8903), .A2(n6278), .ZN(n10444) );
  NAND2_X1 U7259 ( .A1(n10445), .A2(n10444), .ZN(n10443) );
  OR2_X1 U7260 ( .A1(n10572), .A2(n10464), .ZN(n6129) );
  NAND2_X1 U7261 ( .A1(n10443), .A2(n6129), .ZN(n10424) );
  NAND2_X1 U7262 ( .A1(n6132), .A2(SI_21_), .ZN(n6133) );
  MUX2_X1 U7263 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n7159), .Z(n6149) );
  XNOR2_X1 U7264 ( .A(n6149), .B(SI_22_), .ZN(n6146) );
  XNOR2_X1 U7265 ( .A(n6148), .B(n6146), .ZN(n8236) );
  NAND2_X1 U7266 ( .A1(n8236), .A2(n5948), .ZN(n6136) );
  INV_X1 U7267 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8240) );
  OR2_X1 U7268 ( .A1(n8777), .A2(n8240), .ZN(n6135) );
  INV_X1 U7269 ( .A(n6138), .ZN(n6137) );
  INV_X1 U7270 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U7271 ( .A1(n6138), .A2(n10145), .ZN(n6139) );
  NAND2_X1 U7272 ( .A1(n6159), .A2(n6139), .ZN(n10429) );
  OR2_X1 U7273 ( .A1(n10429), .A2(n6301), .ZN(n6144) );
  INV_X1 U7274 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10428) );
  NAND2_X1 U7275 ( .A1(n8647), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7276 ( .A1(n5807), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6140) );
  OAI211_X1 U7277 ( .C1(n10428), .C2(n6305), .A(n6141), .B(n6140), .ZN(n6142)
         );
  INV_X1 U7278 ( .A(n6142), .ZN(n6143) );
  NAND2_X1 U7279 ( .A1(n6144), .A2(n6143), .ZN(n10441) );
  NAND2_X1 U7280 ( .A1(n10568), .A2(n10082), .ZN(n8747) );
  NAND2_X1 U7281 ( .A1(n10410), .A2(n8747), .ZN(n10423) );
  NAND2_X1 U7282 ( .A1(n10424), .A2(n10423), .ZN(n10422) );
  OR2_X1 U7283 ( .A1(n10568), .A2(n10441), .ZN(n6145) );
  INV_X1 U7284 ( .A(n6146), .ZN(n6147) );
  NAND2_X1 U7285 ( .A1(n6149), .A2(SI_22_), .ZN(n6150) );
  MUX2_X1 U7286 ( .A(n8268), .B(n9782), .S(n7159), .Z(n6151) );
  NAND2_X1 U7287 ( .A1(n6151), .A2(n9674), .ZN(n6168) );
  INV_X1 U7288 ( .A(n6151), .ZN(n6152) );
  NAND2_X1 U7289 ( .A1(n6152), .A2(SI_23_), .ZN(n6153) );
  NAND2_X1 U7290 ( .A1(n6168), .A2(n6153), .ZN(n6154) );
  NAND2_X1 U7291 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  NAND2_X1 U7292 ( .A1(n8265), .A2(n5948), .ZN(n6158) );
  OR2_X1 U7293 ( .A1(n8777), .A2(n9782), .ZN(n6157) );
  INV_X1 U7294 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U7295 ( .A1(n6159), .A2(n10061), .ZN(n6160) );
  NAND2_X1 U7296 ( .A1(n6175), .A2(n6160), .ZN(n10407) );
  OR2_X1 U7297 ( .A1(n10407), .A2(n6301), .ZN(n6165) );
  INV_X1 U7298 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n10406) );
  NAND2_X1 U7299 ( .A1(n5807), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7300 ( .A1(n8647), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6161) );
  OAI211_X1 U7301 ( .C1(n10406), .C2(n6305), .A(n6162), .B(n6161), .ZN(n6163)
         );
  INV_X1 U7302 ( .A(n6163), .ZN(n6164) );
  NAND2_X1 U7303 ( .A1(n6165), .A2(n6164), .ZN(n10433) );
  NOR2_X1 U7304 ( .A1(n10405), .A2(n10433), .ZN(n6166) );
  NAND2_X1 U7305 ( .A1(n10405), .A2(n10433), .ZN(n6167) );
  INV_X1 U7306 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8986) );
  MUX2_X1 U7307 ( .A(n8986), .B(n9569), .S(n7159), .Z(n6170) );
  INV_X1 U7308 ( .A(SI_24_), .ZN(n9667) );
  NAND2_X1 U7309 ( .A1(n6170), .A2(n9667), .ZN(n6186) );
  INV_X1 U7310 ( .A(n6170), .ZN(n6171) );
  NAND2_X1 U7311 ( .A1(n6171), .A2(SI_24_), .ZN(n6172) );
  XNOR2_X1 U7312 ( .A(n6185), .B(n6184), .ZN(n8372) );
  NAND2_X1 U7313 ( .A1(n8372), .A2(n5948), .ZN(n6174) );
  OR2_X1 U7314 ( .A1(n8777), .A2(n9569), .ZN(n6173) );
  INV_X1 U7315 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U7316 ( .A1(n6175), .A2(n10125), .ZN(n6176) );
  AND2_X1 U7317 ( .A1(n6191), .A2(n6176), .ZN(n10395) );
  NAND2_X1 U7318 ( .A1(n10395), .A2(n6235), .ZN(n6182) );
  INV_X1 U7319 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7320 ( .A1(n8647), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7321 ( .A1(n5807), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6177) );
  OAI211_X1 U7322 ( .C1(n6179), .C2(n6305), .A(n6178), .B(n6177), .ZN(n6180)
         );
  INV_X1 U7323 ( .A(n6180), .ZN(n6181) );
  AND2_X1 U7324 ( .A1(n10558), .A2(n10416), .ZN(n6183) );
  NAND2_X1 U7325 ( .A1(n6185), .A2(n6184), .ZN(n6187) );
  INV_X1 U7326 ( .A(SI_25_), .ZN(n9460) );
  XNOR2_X1 U7327 ( .A(n6203), .B(n9460), .ZN(n6200) );
  XNOR2_X1 U7328 ( .A(n6202), .B(n6200), .ZN(n8450) );
  NAND2_X1 U7329 ( .A1(n8450), .A2(n5948), .ZN(n6189) );
  INV_X1 U7330 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8451) );
  OR2_X1 U7331 ( .A1(n8777), .A2(n8451), .ZN(n6188) );
  INV_X1 U7332 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U7333 ( .A1(n6191), .A2(n10089), .ZN(n6192) );
  NAND2_X1 U7334 ( .A1(n6212), .A2(n6192), .ZN(n10375) );
  INV_X1 U7335 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10374) );
  NAND2_X1 U7336 ( .A1(n5807), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7337 ( .A1(n8647), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6193) );
  OAI211_X1 U7338 ( .C1(n10374), .C2(n6305), .A(n6194), .B(n6193), .ZN(n6195)
         );
  INV_X1 U7339 ( .A(n6195), .ZN(n6196) );
  NOR2_X1 U7340 ( .A1(n10373), .A2(n10391), .ZN(n6199) );
  NAND2_X1 U7341 ( .A1(n10373), .A2(n10391), .ZN(n6198) );
  INV_X1 U7342 ( .A(n6200), .ZN(n6201) );
  NAND2_X1 U7343 ( .A1(n6203), .A2(SI_25_), .ZN(n6204) );
  INV_X1 U7344 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8478) );
  INV_X1 U7345 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8481) );
  MUX2_X1 U7346 ( .A(n8478), .B(n8481), .S(n7159), .Z(n6205) );
  INV_X1 U7347 ( .A(SI_26_), .ZN(n9666) );
  NAND2_X1 U7348 ( .A1(n6205), .A2(n9666), .ZN(n6221) );
  INV_X1 U7349 ( .A(n6205), .ZN(n6206) );
  NAND2_X1 U7350 ( .A1(n6206), .A2(SI_26_), .ZN(n6207) );
  NAND2_X1 U7351 ( .A1(n6221), .A2(n6207), .ZN(n6222) );
  NAND2_X1 U7352 ( .A1(n8476), .A2(n5948), .ZN(n6209) );
  OR2_X1 U7353 ( .A1(n8777), .A2(n8481), .ZN(n6208) );
  INV_X1 U7354 ( .A(n6212), .ZN(n6210) );
  NAND2_X1 U7355 ( .A1(n6210), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6233) );
  INV_X1 U7356 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7357 ( .A1(n6212), .A2(n6211), .ZN(n6213) );
  NAND2_X1 U7358 ( .A1(n6233), .A2(n6213), .ZN(n10355) );
  INV_X1 U7359 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U7360 ( .A1(n8647), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7361 ( .A1(n5807), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6214) );
  OAI211_X1 U7362 ( .C1(n10354), .C2(n6305), .A(n6215), .B(n6214), .ZN(n6216)
         );
  INV_X1 U7363 ( .A(n6216), .ZN(n6217) );
  INV_X1 U7364 ( .A(n10381), .ZN(n10090) );
  OR2_X1 U7365 ( .A1(n10353), .A2(n10090), .ZN(n8832) );
  NAND2_X1 U7366 ( .A1(n10353), .A2(n10090), .ZN(n8758) );
  NAND2_X1 U7367 ( .A1(n8832), .A2(n8758), .ZN(n10358) );
  NAND2_X1 U7368 ( .A1(n10351), .A2(n10358), .ZN(n6220) );
  NAND2_X1 U7369 ( .A1(n10353), .A2(n10381), .ZN(n6219) );
  NAND2_X1 U7370 ( .A1(n6220), .A2(n6219), .ZN(n10334) );
  INV_X1 U7371 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6388) );
  INV_X1 U7372 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9774) );
  MUX2_X1 U7373 ( .A(n6388), .B(n9774), .S(n7159), .Z(n6224) );
  INV_X1 U7374 ( .A(SI_27_), .ZN(n9459) );
  NAND2_X1 U7375 ( .A1(n6224), .A2(n9459), .ZN(n6245) );
  INV_X1 U7376 ( .A(n6224), .ZN(n6225) );
  NAND2_X1 U7377 ( .A1(n6225), .A2(SI_27_), .ZN(n6226) );
  NAND2_X1 U7378 ( .A1(n6228), .A2(n6227), .ZN(n6246) );
  OR2_X1 U7379 ( .A1(n6228), .A2(n6227), .ZN(n6229) );
  NAND2_X1 U7380 ( .A1(n6246), .A2(n6229), .ZN(n8482) );
  NAND2_X1 U7381 ( .A1(n8482), .A2(n5948), .ZN(n6231) );
  OR2_X1 U7382 ( .A1(n8777), .A2(n9774), .ZN(n6230) );
  INV_X1 U7383 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7384 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  NAND2_X1 U7385 ( .A1(n10345), .A2(n6235), .ZN(n6241) );
  INV_X1 U7386 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7387 ( .A1(n5807), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7388 ( .A1(n8647), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6236) );
  OAI211_X1 U7389 ( .C1(n6238), .C2(n6305), .A(n6237), .B(n6236), .ZN(n6239)
         );
  INV_X1 U7390 ( .A(n6239), .ZN(n6240) );
  INV_X1 U7391 ( .A(n10363), .ZN(n6242) );
  NOR2_X1 U7392 ( .A1(n10344), .A2(n6242), .ZN(n8834) );
  INV_X1 U7393 ( .A(n8834), .ZN(n6298) );
  AND2_X1 U7394 ( .A1(n10344), .A2(n6242), .ZN(n8821) );
  INV_X1 U7395 ( .A(n8821), .ZN(n6243) );
  OR2_X1 U7396 ( .A1(n10344), .A2(n10363), .ZN(n6244) );
  MUX2_X1 U7397 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7159), .Z(n6740) );
  INV_X1 U7398 ( .A(SI_28_), .ZN(n9662) );
  XNOR2_X1 U7399 ( .A(n6740), .B(n9662), .ZN(n6738) );
  NAND2_X1 U7400 ( .A1(n8532), .A2(n5948), .ZN(n6248) );
  INV_X1 U7401 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8563) );
  OR2_X1 U7402 ( .A1(n8777), .A2(n8563), .ZN(n6247) );
  INV_X1 U7403 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7404 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  NAND2_X1 U7405 ( .A1(n8935), .A2(n6251), .ZN(n10324) );
  INV_X1 U7406 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10323) );
  NAND2_X1 U7407 ( .A1(n5807), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7408 ( .A1(n8647), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6252) );
  OAI211_X1 U7409 ( .C1(n10323), .C2(n6305), .A(n6253), .B(n6252), .ZN(n6254)
         );
  INV_X1 U7410 ( .A(n6254), .ZN(n6255) );
  INV_X1 U7411 ( .A(n10338), .ZN(n6257) );
  NOR2_X1 U7412 ( .A1(n10325), .A2(n6257), .ZN(n8766) );
  INV_X1 U7413 ( .A(n8766), .ZN(n8836) );
  INV_X1 U7414 ( .A(n8939), .ZN(n6258) );
  NAND2_X1 U7415 ( .A1(n8836), .A2(n6258), .ZN(n8809) );
  INV_X1 U7416 ( .A(n8809), .ZN(n6259) );
  AND2_X1 U7417 ( .A1(n6260), .A2(n6259), .ZN(n6261) );
  NAND3_X1 U7418 ( .A1(n6264), .A2(n6263), .A3(n6262), .ZN(n6265) );
  NOR2_X2 U7419 ( .A1(n6266), .A2(n6265), .ZN(n6270) );
  AND2_X2 U7420 ( .A1(n6267), .A2(n9627), .ZN(n6318) );
  OR2_X1 U7421 ( .A1(n6318), .A2(n5803), .ZN(n6344) );
  XNOR2_X2 U7422 ( .A(n6344), .B(n6343), .ZN(n6274) );
  NAND2_X2 U7423 ( .A1(n8852), .A2(n6275), .ZN(n6852) );
  INV_X1 U7424 ( .A(n6267), .ZN(n6268) );
  INV_X1 U7425 ( .A(n6270), .ZN(n6271) );
  NAND2_X1 U7426 ( .A1(n6271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7427 ( .A1(n6310), .A2(n8921), .ZN(n7577) );
  OR2_X1 U7428 ( .A1(n6852), .A2(n7577), .ZN(n7571) );
  NAND2_X1 U7429 ( .A1(n6274), .A2(n8818), .ZN(n7112) );
  INV_X1 U7430 ( .A(n8919), .ZN(n6848) );
  NAND2_X1 U7431 ( .A1(n6848), .A2(n6852), .ZN(n6276) );
  NAND3_X1 U7432 ( .A1(n7571), .A2(n7112), .A3(n6276), .ZN(n8359) );
  NAND2_X1 U7433 ( .A1(n6274), .A2(n8923), .ZN(n8815) );
  INV_X1 U7434 ( .A(n8921), .ZN(n8856) );
  INV_X1 U7435 ( .A(n10433), .ZN(n10147) );
  NAND2_X1 U7436 ( .A1(n10405), .A2(n10147), .ZN(n8828) );
  NAND2_X1 U7437 ( .A1(n8750), .A2(n8828), .ZN(n10411) );
  INV_X1 U7438 ( .A(n10411), .ZN(n6297) );
  INV_X1 U7439 ( .A(n10438), .ZN(n6277) );
  NAND2_X1 U7440 ( .A1(n8903), .A2(n6277), .ZN(n6279) );
  NAND2_X1 U7441 ( .A1(n6279), .A2(n6278), .ZN(n8823) );
  INV_X1 U7442 ( .A(n8823), .ZN(n6296) );
  INV_X1 U7443 ( .A(n10510), .ZN(n10116) );
  OR2_X1 U7444 ( .A1(n10498), .A2(n10116), .ZN(n8896) );
  INV_X1 U7445 ( .A(n10492), .ZN(n6295) );
  OR2_X1 U7446 ( .A1(n10594), .A2(n6295), .ZN(n10487) );
  AND2_X1 U7447 ( .A1(n8896), .A2(n10487), .ZN(n8862) );
  AND2_X1 U7448 ( .A1(n8725), .A2(n8379), .ZN(n8893) );
  INV_X1 U7449 ( .A(n8802), .ZN(n6294) );
  INV_X1 U7450 ( .A(n10204), .ZN(n8354) );
  OR2_X1 U7451 ( .A1(n8214), .A2(n8354), .ZN(n8662) );
  NAND2_X1 U7452 ( .A1(n8214), .A2(n8354), .ZN(n8715) );
  AND2_X1 U7453 ( .A1(n8694), .A2(n6280), .ZN(n8699) );
  INV_X1 U7454 ( .A(n8699), .ZN(n6281) );
  INV_X1 U7455 ( .A(n7797), .ZN(n8685) );
  NOR2_X1 U7456 ( .A1(n6281), .A2(n8685), .ZN(n8792) );
  INV_X1 U7457 ( .A(n8792), .ZN(n6284) );
  NAND2_X1 U7458 ( .A1(n6282), .A2(n8694), .ZN(n6283) );
  NAND2_X1 U7459 ( .A1(n6284), .A2(n6283), .ZN(n6285) );
  OAI21_X1 U7460 ( .B1(n8877), .B2(n8790), .A(n6285), .ZN(n8880) );
  AND2_X1 U7461 ( .A1(n6861), .A2(n10932), .ZN(n7451) );
  INV_X1 U7462 ( .A(n5122), .ZN(n8864) );
  OR2_X1 U7463 ( .A1(n10214), .A2(n8864), .ZN(n6287) );
  NAND2_X1 U7464 ( .A1(n7450), .A2(n6287), .ZN(n7303) );
  NAND2_X1 U7465 ( .A1(n10213), .A2(n7335), .ZN(n8868) );
  NAND2_X1 U7466 ( .A1(n7462), .A2(n10995), .ZN(n8671) );
  AND2_X1 U7467 ( .A1(n8671), .A2(n8871), .ZN(n6288) );
  INV_X1 U7468 ( .A(n10995), .ZN(n7601) );
  NAND2_X1 U7469 ( .A1(n7601), .A2(n10211), .ZN(n8666) );
  INV_X1 U7470 ( .A(n8873), .ZN(n6290) );
  INV_X1 U7471 ( .A(n8669), .ZN(n7748) );
  NOR2_X1 U7472 ( .A1(n7748), .A2(n8877), .ZN(n6291) );
  OR2_X1 U7473 ( .A1(n8880), .A2(n6291), .ZN(n7833) );
  NAND2_X1 U7474 ( .A1(n7833), .A2(n5522), .ZN(n7834) );
  INV_X1 U7475 ( .A(n10205), .ZN(n8172) );
  NAND2_X1 U7476 ( .A1(n11089), .A2(n8172), .ZN(n8708) );
  AND2_X1 U7477 ( .A1(n8708), .A2(n8698), .ZN(n8881) );
  OR2_X1 U7478 ( .A1(n11089), .A2(n8172), .ZN(n8707) );
  INV_X1 U7479 ( .A(n11090), .ZN(n6966) );
  OR2_X1 U7480 ( .A1(n7956), .A2(n6966), .ZN(n8713) );
  NAND2_X1 U7481 ( .A1(n7956), .A2(n6966), .ZN(n8883) );
  NAND2_X1 U7482 ( .A1(n8713), .A2(n8883), .ZN(n8797) );
  INV_X1 U7483 ( .A(n8797), .ZN(n6292) );
  NAND3_X1 U7484 ( .A1(n8800), .A2(n8351), .A3(n8715), .ZN(n6293) );
  NAND2_X1 U7485 ( .A1(n6293), .A2(n8663), .ZN(n8321) );
  INV_X1 U7486 ( .A(n8726), .ZN(n8891) );
  NAND2_X1 U7487 ( .A1(n10594), .A2(n6295), .ZN(n8894) );
  AND2_X1 U7488 ( .A1(n10498), .A2(n10116), .ZN(n8728) );
  NAND3_X1 U7489 ( .A1(n6297), .A2(n10410), .A3(n10432), .ZN(n10414) );
  AND2_X1 U7490 ( .A1(n10414), .A2(n8828), .ZN(n10390) );
  INV_X1 U7491 ( .A(n10416), .ZN(n10091) );
  NAND2_X1 U7492 ( .A1(n10558), .A2(n10091), .ZN(n8822) );
  NAND2_X1 U7493 ( .A1(n10390), .A2(n10389), .ZN(n10388) );
  NAND2_X1 U7494 ( .A1(n10388), .A2(n8825), .ZN(n10380) );
  INV_X1 U7495 ( .A(n10391), .ZN(n10126) );
  OR2_X1 U7496 ( .A1(n10373), .A2(n10126), .ZN(n8829) );
  NAND2_X1 U7497 ( .A1(n10373), .A2(n10126), .ZN(n8757) );
  NAND2_X1 U7498 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  NAND2_X1 U7499 ( .A1(n10378), .A2(n8829), .ZN(n10359) );
  AND2_X1 U7500 ( .A1(n10361), .A2(n8758), .ZN(n10337) );
  OR2_X1 U7501 ( .A1(n6274), .A2(n8259), .ZN(n6300) );
  OR2_X1 U7502 ( .A1(n8818), .A2(n8921), .ZN(n6299) );
  OR2_X1 U7503 ( .A1(n8935), .A2(n6301), .ZN(n6309) );
  INV_X1 U7504 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7505 ( .A1(n8647), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6304) );
  INV_X1 U7506 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6302) );
  OR2_X1 U7507 ( .A1(n8649), .A2(n6302), .ZN(n6303) );
  OAI211_X1 U7508 ( .C1(n6306), .C2(n6305), .A(n6304), .B(n6303), .ZN(n6307)
         );
  INV_X1 U7509 ( .A(n6307), .ZN(n6308) );
  NAND2_X1 U7510 ( .A1(n8852), .A2(n6310), .ZN(n7193) );
  INV_X1 U7511 ( .A(n5124), .ZN(n7248) );
  AOI22_X1 U7512 ( .A1(n7886), .A2(n10509), .B1(n10507), .B2(n10363), .ZN(
        n6312) );
  NAND2_X1 U7513 ( .A1(n6313), .A2(n6312), .ZN(n10330) );
  INV_X1 U7514 ( .A(n10572), .ZN(n10449) );
  INV_X1 U7515 ( .A(n10197), .ZN(n10606) );
  INV_X1 U7516 ( .A(n11017), .ZN(n7384) );
  AND2_X1 U7517 ( .A1(n7598), .A2(n7384), .ZN(n7381) );
  INV_X1 U7518 ( .A(n10166), .ZN(n11029) );
  NAND2_X1 U7519 ( .A1(n7381), .A2(n11029), .ZN(n7747) );
  OR2_X1 U7520 ( .A1(n7747), .A2(n7784), .ZN(n7746) );
  INV_X1 U7521 ( .A(n7946), .ZN(n11065) );
  OR2_X2 U7522 ( .A1(n8214), .A2(n8147), .ZN(n8364) );
  NOR2_X2 U7523 ( .A1(n10612), .A2(n8364), .ZN(n8363) );
  OR2_X2 U7524 ( .A1(n10496), .A2(n10479), .ZN(n10477) );
  NOR2_X2 U7525 ( .A1(n10578), .A2(n10477), .ZN(n10458) );
  NAND2_X1 U7526 ( .A1(n10449), .A2(n10458), .ZN(n10446) );
  INV_X1 U7527 ( .A(n7112), .ZN(n10933) );
  AOI21_X1 U7528 ( .B1(n10325), .B2(n10341), .A(n11049), .ZN(n6316) );
  AND2_X1 U7529 ( .A1(n6316), .A2(n5715), .ZN(n10329) );
  NAND2_X2 U7530 ( .A1(n6318), .A2(n6317), .ZN(n6319) );
  OAI21_X4 U7531 ( .B1(n6319), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6323) );
  XNOR2_X2 U7532 ( .A(n6323), .B(n6322), .ZN(n8452) );
  NAND2_X1 U7533 ( .A1(n8452), .A2(P1_B_REG_SCAN_IN), .ZN(n6321) );
  MUX2_X1 U7534 ( .A(n6321), .B(P1_B_REG_SCAN_IN), .S(n6351), .Z(n6327) );
  NAND2_X1 U7535 ( .A1(n6323), .A2(n6322), .ZN(n6324) );
  XNOR2_X2 U7536 ( .A(n6325), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6342) );
  INV_X1 U7537 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7188) );
  INV_X1 U7538 ( .A(n6326), .ZN(n8479) );
  AND2_X1 U7539 ( .A1(n8479), .A2(n8452), .ZN(n6328) );
  NAND2_X1 U7540 ( .A1(n10599), .A2(n8923), .ZN(n7114) );
  INV_X1 U7541 ( .A(n7114), .ZN(n6329) );
  OR2_X1 U7542 ( .A1(n7565), .A2(n6329), .ZN(n6350) );
  NOR2_X1 U7543 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .ZN(
        n6333) );
  NOR4_X1 U7544 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6332) );
  NOR4_X1 U7545 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6331) );
  NOR4_X1 U7546 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6330) );
  NAND4_X1 U7547 ( .A1(n6333), .A2(n6332), .A3(n6331), .A4(n6330), .ZN(n6339)
         );
  NOR4_X1 U7548 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6337) );
  NOR4_X1 U7549 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6336) );
  NOR4_X1 U7550 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6335) );
  NOR4_X1 U7551 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6334) );
  NAND4_X1 U7552 ( .A1(n6337), .A2(n6336), .A3(n6335), .A4(n6334), .ZN(n6338)
         );
  OAI21_X1 U7553 ( .B1(n6339), .B2(n6338), .A(n7182), .ZN(n7097) );
  INV_X1 U7554 ( .A(n6351), .ZN(n6340) );
  NOR2_X2 U7555 ( .A1(n8452), .A2(n6340), .ZN(n6341) );
  NAND2_X2 U7556 ( .A1(n6341), .A2(n6342), .ZN(n6854) );
  NAND2_X1 U7557 ( .A1(n6344), .A2(n6343), .ZN(n6345) );
  NAND2_X1 U7558 ( .A1(n6345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6347) );
  OR2_X1 U7559 ( .A1(n7193), .A2(n8919), .ZN(n7102) );
  INV_X1 U7560 ( .A(n7102), .ZN(n6348) );
  NOR2_X1 U7561 ( .A1(n8851), .A2(n6348), .ZN(n6349) );
  NAND2_X1 U7562 ( .A1(n7097), .A2(n6349), .ZN(n7564) );
  INV_X1 U7563 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7191) );
  INV_X1 U7564 ( .A(n7098), .ZN(n7567) );
  NAND2_X1 U7565 ( .A1(n10325), .A2(n8213), .ZN(n6352) );
  NOR2_X1 U7566 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6357) );
  NOR2_X1 U7567 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6361) );
  NOR2_X1 U7568 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6360) );
  NAND4_X1 U7569 ( .A1(n6361), .A2(n6360), .A3(n6753), .A4(n6756), .ZN(n6363)
         );
  NOR2_X1 U7570 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6362) );
  NAND4_X1 U7571 ( .A1(n6362), .A2(n6593), .A3(n6581), .A4(n6567), .ZN(n6624)
         );
  NAND2_X1 U7572 ( .A1(n6802), .A2(n6366), .ZN(n6812) );
  OR2_X2 U7573 ( .A1(n6812), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6384) );
  XNOR2_X2 U7574 ( .A(n6368), .B(n10050), .ZN(n8996) );
  XNOR2_X2 U7575 ( .A(n6371), .B(n6370), .ZN(n8635) );
  NAND2_X1 U7576 ( .A1(n5121), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6381) );
  NAND2_X4 U7577 ( .A1(n6373), .A2(n8996), .ZN(n9091) );
  INV_X1 U7578 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6372) );
  OR2_X1 U7579 ( .A1(n9091), .A2(n6372), .ZN(n6380) );
  NAND2_X1 U7580 ( .A1(n6446), .A2(n7642), .ZN(n6460) );
  INV_X1 U7581 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9735) );
  AND2_X1 U7582 ( .A1(n6375), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6376) );
  NOR2_X1 U7583 ( .A1(n6731), .A2(n6376), .ZN(n9878) );
  OR2_X1 U7584 ( .A1(n6701), .A2(n9878), .ZN(n6379) );
  INV_X1 U7585 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9879) );
  OR2_X1 U7586 ( .A1(n6733), .A2(n9879), .ZN(n6378) );
  INV_X1 U7587 ( .A(n6384), .ZN(n6385) );
  NAND2_X1 U7588 ( .A1(n6803), .A2(n6385), .ZN(n6816) );
  INV_X2 U7589 ( .A(n6466), .ZN(n6499) );
  NAND2_X1 U7590 ( .A1(n8482), .A2(n6499), .ZN(n6390) );
  OR2_X1 U7591 ( .A1(n9101), .A2(n6388), .ZN(n6389) );
  INV_X1 U7592 ( .A(n9996), .ZN(n9007) );
  NAND2_X1 U7593 ( .A1(n6601), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6394) );
  INV_X1 U7594 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8072) );
  OR2_X1 U7595 ( .A1(n6701), .A2(n8072), .ZN(n6393) );
  INV_X1 U7596 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7323) );
  INV_X1 U7597 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7324) );
  OR2_X1 U7598 ( .A1(n6477), .A2(n7324), .ZN(n6391) );
  NAND4_X2 U7599 ( .A1(n6394), .A2(n6393), .A3(n6392), .A4(n6391), .ZN(n6408)
         );
  NAND2_X1 U7600 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6396) );
  MUX2_X1 U7601 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6396), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6397) );
  NAND2_X2 U7602 ( .A1(n6399), .A2(n6398), .ZN(n9125) );
  NAND2_X1 U7603 ( .A1(n6408), .A2(n8073), .ZN(n9127) );
  NAND2_X2 U7604 ( .A1(n9125), .A2(n9127), .ZN(n9270) );
  NAND2_X1 U7605 ( .A1(n5121), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6403) );
  INV_X1 U7606 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10951) );
  OR2_X1 U7607 ( .A1(n6701), .A2(n10951), .ZN(n6402) );
  INV_X1 U7608 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7320) );
  OR2_X1 U7609 ( .A1(n9091), .A2(n7320), .ZN(n6401) );
  INV_X1 U7610 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10947) );
  OR2_X1 U7611 ( .A1(n6477), .A2(n10947), .ZN(n6400) );
  NAND4_X1 U7612 ( .A1(n6403), .A2(n6402), .A3(n6401), .A4(n6400), .ZN(n9337)
         );
  INV_X1 U7613 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7319) );
  NAND2_X1 U7614 ( .A1(n5120), .A2(SI_0_), .ZN(n6405) );
  INV_X1 U7615 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U7616 ( .A1(n6405), .A2(n6404), .ZN(n6407) );
  AND2_X1 U7617 ( .A1(n6407), .A2(n6406), .ZN(n10056) );
  MUX2_X1 U7618 ( .A(P2_IR_REG_0__SCAN_IN), .B(n10056), .S(n7153), .Z(n10938)
         );
  NAND2_X1 U7619 ( .A1(n9337), .A2(n10938), .ZN(n8069) );
  OR2_X1 U7620 ( .A1(n6408), .A2(n6398), .ZN(n10965) );
  NAND2_X1 U7621 ( .A1(n8068), .A2(n10965), .ZN(n6419) );
  NAND2_X1 U7622 ( .A1(n5121), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6412) );
  INV_X1 U7623 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10876) );
  OR2_X1 U7624 ( .A1(n6701), .A2(n10876), .ZN(n6411) );
  INV_X1 U7625 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7413) );
  OR2_X1 U7626 ( .A1(n9091), .A2(n7413), .ZN(n6410) );
  INV_X1 U7627 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7414) );
  OR2_X1 U7628 ( .A1(n6477), .A2(n7414), .ZN(n6409) );
  OR2_X1 U7629 ( .A1(n6466), .A2(n7169), .ZN(n6418) );
  INV_X1 U7630 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7160) );
  OR2_X1 U7631 ( .A1(n7153), .A2(n10886), .ZN(n6416) );
  AND3_X2 U7632 ( .A1(n6418), .A2(n6417), .A3(n6416), .ZN(n10963) );
  OR2_X2 U7633 ( .A1(n9335), .A2(n10963), .ZN(n9133) );
  NAND2_X1 U7634 ( .A1(n9335), .A2(n10963), .ZN(n9132) );
  NAND2_X1 U7635 ( .A1(n6419), .A2(n9272), .ZN(n10964) );
  OR2_X1 U7636 ( .A1(n9335), .A2(n10977), .ZN(n6420) );
  NAND2_X1 U7637 ( .A1(n10964), .A2(n6420), .ZN(n7976) );
  NAND2_X1 U7638 ( .A1(n5121), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6425) );
  INV_X1 U7639 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6421) );
  OR2_X1 U7640 ( .A1(n9091), .A2(n6421), .ZN(n6424) );
  OR2_X1 U7641 ( .A1(n6477), .A2(n7538), .ZN(n6423) );
  OR2_X1 U7642 ( .A1(n6466), .A2(n7161), .ZN(n6431) );
  INV_X1 U7643 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7162) );
  OR2_X1 U7644 ( .A1(n9101), .A2(n7162), .ZN(n6430) );
  NAND2_X1 U7645 ( .A1(n6413), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6426) );
  MUX2_X1 U7646 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6426), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6428) );
  AND2_X1 U7647 ( .A1(n6428), .A2(n6427), .ZN(n7412) );
  OR2_X1 U7648 ( .A1(n7153), .A2(n7546), .ZN(n6429) );
  AND3_X2 U7649 ( .A1(n6431), .A2(n6430), .A3(n6429), .ZN(n10982) );
  OR2_X1 U7650 ( .A1(n9334), .A2(n10982), .ZN(n9142) );
  NAND2_X1 U7651 ( .A1(n9334), .A2(n10982), .ZN(n9149) );
  NAND2_X1 U7652 ( .A1(n7976), .A2(n7975), .ZN(n6433) );
  INV_X1 U7653 ( .A(n10982), .ZN(n7557) );
  OR2_X1 U7654 ( .A1(n9334), .A2(n7557), .ZN(n6432) );
  NAND2_X1 U7655 ( .A1(n5121), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6440) );
  INV_X1 U7656 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6434) );
  OR2_X1 U7657 ( .A1(n9091), .A2(n6434), .ZN(n6439) );
  AND2_X1 U7658 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6435) );
  NOR2_X1 U7659 ( .A1(n6446), .A2(n6435), .ZN(n7882) );
  OR2_X1 U7660 ( .A1(n6701), .A2(n7882), .ZN(n6438) );
  INV_X1 U7661 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6436) );
  OR2_X1 U7662 ( .A1(n6477), .A2(n6436), .ZN(n6437) );
  NAND4_X1 U7663 ( .A1(n6440), .A2(n6439), .A3(n6438), .A4(n6437), .ZN(n9333)
         );
  XNOR2_X1 U7664 ( .A(n6454), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7410) );
  OR2_X1 U7665 ( .A1(n6466), .A2(n7171), .ZN(n6442) );
  INV_X1 U7666 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7165) );
  OR2_X1 U7667 ( .A1(n9101), .A2(n7165), .ZN(n6441) );
  OAI211_X1 U7668 ( .C1(n7153), .C2(n7520), .A(n6442), .B(n6441), .ZN(n7635)
         );
  NOR2_X1 U7669 ( .A1(n9333), .A2(n7635), .ZN(n6444) );
  NAND2_X1 U7670 ( .A1(n9333), .A2(n7635), .ZN(n6443) );
  NAND2_X1 U7671 ( .A1(n5121), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6452) );
  INV_X1 U7672 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6445) );
  OR2_X1 U7673 ( .A1(n9091), .A2(n6445), .ZN(n6451) );
  OR2_X1 U7674 ( .A1(n6446), .A2(n7642), .ZN(n6447) );
  AND2_X1 U7675 ( .A1(n6460), .A2(n6447), .ZN(n8089) );
  OR2_X1 U7676 ( .A1(n6701), .A2(n8089), .ZN(n6450) );
  INV_X1 U7677 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6448) );
  OR2_X1 U7678 ( .A1(n6477), .A2(n6448), .ZN(n6449) );
  NAND4_X1 U7679 ( .A1(n6452), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(n9332)
         );
  NAND2_X1 U7680 ( .A1(n6454), .A2(n6453), .ZN(n6455) );
  NAND2_X1 U7681 ( .A1(n6455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6468) );
  XNOR2_X1 U7682 ( .A(n6468), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7693) );
  INV_X1 U7683 ( .A(n7693), .ZN(n7683) );
  OR2_X1 U7684 ( .A1(n6466), .A2(n7163), .ZN(n6457) );
  INV_X1 U7685 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7164) );
  OR2_X1 U7686 ( .A1(n9101), .A2(n7164), .ZN(n6456) );
  OAI211_X1 U7687 ( .C1(n7153), .C2(n7683), .A(n6457), .B(n6456), .ZN(n7617)
         );
  AND2_X1 U7688 ( .A1(n9332), .A2(n7617), .ZN(n6458) );
  NAND2_X1 U7689 ( .A1(n5121), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6465) );
  INV_X1 U7690 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6459) );
  OR2_X1 U7691 ( .A1(n9091), .A2(n6459), .ZN(n6464) );
  NAND2_X1 U7692 ( .A1(n6460), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6461) );
  AND2_X1 U7693 ( .A1(n6478), .A2(n6461), .ZN(n7621) );
  OR2_X1 U7694 ( .A1(n6701), .A2(n7621), .ZN(n6463) );
  OR2_X1 U7695 ( .A1(n6477), .A2(n7679), .ZN(n6462) );
  NAND4_X1 U7696 ( .A1(n6465), .A2(n6464), .A3(n6463), .A4(n6462), .ZN(n9331)
         );
  OR2_X1 U7697 ( .A1(n6466), .A2(n7166), .ZN(n6472) );
  INV_X1 U7698 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7167) );
  OR2_X1 U7699 ( .A1(n9101), .A2(n7167), .ZN(n6471) );
  NAND2_X1 U7700 ( .A1(n6468), .A2(n6467), .ZN(n6469) );
  NAND2_X1 U7701 ( .A1(n6469), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6485) );
  XNOR2_X1 U7702 ( .A(n6485), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7696) );
  OR2_X1 U7703 ( .A1(n7153), .A2(n10903), .ZN(n6470) );
  NAND2_X1 U7704 ( .A1(n9331), .A2(n7625), .ZN(n9155) );
  NAND2_X1 U7705 ( .A1(n9156), .A2(n9155), .ZN(n9278) );
  INV_X1 U7706 ( .A(n7625), .ZN(n7769) );
  OR2_X1 U7707 ( .A1(n9331), .A2(n7769), .ZN(n6473) );
  NAND2_X1 U7708 ( .A1(n6474), .A2(n6473), .ZN(n7903) );
  NAND2_X1 U7709 ( .A1(n5121), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6483) );
  INV_X1 U7710 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6475) );
  OR2_X1 U7711 ( .A1(n9091), .A2(n6475), .ZN(n6482) );
  INV_X1 U7712 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6476) );
  OR2_X1 U7713 ( .A1(n6477), .A2(n6476), .ZN(n6481) );
  AND2_X1 U7714 ( .A1(n6478), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6479) );
  NOR2_X1 U7715 ( .A1(n6493), .A2(n6479), .ZN(n11040) );
  OR2_X1 U7716 ( .A1(n6701), .A2(n11040), .ZN(n6480) );
  NAND4_X1 U7717 ( .A1(n6483), .A2(n6482), .A3(n6481), .A4(n6480), .ZN(n9330)
         );
  NAND2_X1 U7718 ( .A1(n6485), .A2(n6484), .ZN(n6486) );
  NAND2_X1 U7719 ( .A1(n6486), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6488) );
  INV_X1 U7720 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7721 ( .A1(n6488), .A2(n6487), .ZN(n6500) );
  OR2_X1 U7722 ( .A1(n6488), .A2(n6487), .ZN(n6489) );
  AOI22_X1 U7723 ( .A1(n6642), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6641), .B2(
        n8001), .ZN(n6491) );
  NAND2_X1 U7724 ( .A1(n7172), .A2(n6499), .ZN(n6490) );
  OR2_X1 U7725 ( .A1(n9330), .A2(n7732), .ZN(n9164) );
  NAND2_X1 U7726 ( .A1(n9330), .A2(n7732), .ZN(n7961) );
  NAND2_X1 U7727 ( .A1(n9164), .A2(n7961), .ZN(n9279) );
  NAND2_X1 U7728 ( .A1(n7903), .A2(n9279), .ZN(n7964) );
  INV_X1 U7729 ( .A(n7732), .ZN(n11044) );
  OR2_X1 U7730 ( .A1(n9330), .A2(n11044), .ZN(n7963) );
  NAND2_X1 U7731 ( .A1(n5121), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6498) );
  INV_X1 U7732 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6492) );
  OR2_X1 U7733 ( .A1(n9091), .A2(n6492), .ZN(n6497) );
  NOR2_X1 U7734 ( .A1(n6493), .A2(n7817), .ZN(n6494) );
  OR2_X1 U7735 ( .A1(n6514), .A2(n6494), .ZN(n7969) );
  INV_X1 U7736 ( .A(n7969), .ZN(n7821) );
  OR2_X1 U7737 ( .A1(n6701), .A2(n7821), .ZN(n6496) );
  INV_X1 U7738 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7968) );
  OR2_X1 U7739 ( .A1(n6733), .A2(n7968), .ZN(n6495) );
  NAND2_X1 U7740 ( .A1(n7176), .A2(n6499), .ZN(n6504) );
  NAND2_X1 U7741 ( .A1(n6500), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6502) );
  INV_X1 U7742 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6501) );
  INV_X1 U7743 ( .A(n8103), .ZN(n8010) );
  AOI22_X1 U7744 ( .A1(n6642), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6641), .B2(
        n8010), .ZN(n6503) );
  OR2_X1 U7745 ( .A1(n9329), .A2(n7970), .ZN(n6505) );
  AND2_X1 U7746 ( .A1(n7963), .A2(n6505), .ZN(n6507) );
  INV_X1 U7747 ( .A(n6505), .ZN(n6506) );
  INV_X1 U7748 ( .A(n7970), .ZN(n11059) );
  NAND2_X1 U7749 ( .A1(n11059), .A2(n9329), .ZN(n9153) );
  NAND2_X1 U7750 ( .A1(n9165), .A2(n9153), .ZN(n7965) );
  NAND2_X1 U7751 ( .A1(n7197), .A2(n6499), .ZN(n6513) );
  NOR2_X1 U7752 ( .A1(n6508), .A2(n6521), .ZN(n6509) );
  MUX2_X1 U7753 ( .A(n6521), .B(n6509), .S(P2_IR_REG_9__SCAN_IN), .Z(n6511) );
  OR2_X1 U7754 ( .A1(n6511), .A2(n6510), .ZN(n8102) );
  AOI22_X1 U7755 ( .A1(n6642), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6641), .B2(
        n8193), .ZN(n6512) );
  NAND2_X1 U7756 ( .A1(n5121), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6519) );
  INV_X1 U7757 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8100) );
  OR2_X1 U7758 ( .A1(n9091), .A2(n8100), .ZN(n6518) );
  INV_X1 U7759 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8101) );
  OR2_X1 U7760 ( .A1(n6733), .A2(n8101), .ZN(n6517) );
  OR2_X1 U7761 ( .A1(n6514), .A2(n9744), .ZN(n6515) );
  AND2_X1 U7762 ( .A1(n6525), .A2(n6515), .ZN(n7894) );
  OR2_X1 U7763 ( .A1(n6701), .A2(n7894), .ZN(n6516) );
  NAND2_X1 U7764 ( .A1(n8048), .A2(n7203), .ZN(n9167) );
  NAND2_X1 U7765 ( .A1(n9154), .A2(n9167), .ZN(n9281) );
  OR2_X1 U7766 ( .A1(n8048), .A2(n5260), .ZN(n6520) );
  NAND2_X1 U7767 ( .A1(n7200), .A2(n6499), .ZN(n6524) );
  OR2_X1 U7768 ( .A1(n6510), .A2(n6521), .ZN(n6522) );
  XNOR2_X1 U7769 ( .A(n6522), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8428) );
  AOI22_X1 U7770 ( .A1(n6642), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6641), .B2(
        n8428), .ZN(n6523) );
  NAND2_X1 U7771 ( .A1(n6524), .A2(n6523), .ZN(n11075) );
  NAND2_X1 U7772 ( .A1(n5121), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6530) );
  INV_X1 U7773 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8427) );
  OR2_X1 U7774 ( .A1(n9091), .A2(n8427), .ZN(n6529) );
  NAND2_X1 U7775 ( .A1(n6525), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6526) );
  AND2_X1 U7776 ( .A1(n6537), .A2(n6526), .ZN(n8162) );
  OR2_X1 U7777 ( .A1(n6701), .A2(n8162), .ZN(n6528) );
  INV_X1 U7778 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8421) );
  OR2_X1 U7779 ( .A1(n6733), .A2(n8421), .ZN(n6527) );
  NAND4_X1 U7780 ( .A1(n6530), .A2(n6529), .A3(n6528), .A4(n6527), .ZN(n9328)
         );
  NAND2_X1 U7781 ( .A1(n11075), .A2(n9328), .ZN(n6531) );
  NAND2_X1 U7782 ( .A1(n6532), .A2(n6531), .ZN(n8056) );
  NAND2_X1 U7783 ( .A1(n7212), .A2(n6499), .ZN(n6535) );
  XNOR2_X1 U7784 ( .A(n6544), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U7785 ( .A1(n6642), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6641), .B2(
        n10905), .ZN(n6534) );
  NAND2_X1 U7786 ( .A1(n6535), .A2(n6534), .ZN(n11078) );
  NAND2_X1 U7787 ( .A1(n5121), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6542) );
  INV_X1 U7788 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6536) );
  OR2_X1 U7789 ( .A1(n9091), .A2(n6536), .ZN(n6541) );
  AOI21_X1 U7790 ( .B1(n6537), .B2(P2_REG3_REG_11__SCAN_IN), .A(n6548), .ZN(
        n8232) );
  OR2_X1 U7791 ( .A1(n6701), .A2(n8232), .ZN(n6540) );
  INV_X1 U7792 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6538) );
  OR2_X1 U7793 ( .A1(n6733), .A2(n6538), .ZN(n6539) );
  NAND4_X1 U7794 ( .A1(n6542), .A2(n6541), .A3(n6540), .A4(n6539), .ZN(n9327)
         );
  AND2_X1 U7795 ( .A1(n11078), .A2(n9327), .ZN(n6543) );
  OAI22_X1 U7796 ( .A1(n8056), .A2(n6543), .B1(n9327), .B2(n11078), .ZN(n8218)
         );
  NAND2_X1 U7797 ( .A1(n7260), .A2(n6499), .ZN(n6547) );
  XNOR2_X1 U7798 ( .A(n6557), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8501) );
  AOI22_X1 U7799 ( .A1(n6642), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6641), .B2(
        n8501), .ZN(n6546) );
  NAND2_X1 U7800 ( .A1(n5121), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6554) );
  INV_X1 U7801 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8500) );
  OR2_X1 U7802 ( .A1(n9091), .A2(n8500), .ZN(n6553) );
  INV_X1 U7803 ( .A(n6548), .ZN(n6550) );
  INV_X1 U7804 ( .A(n6561), .ZN(n6549) );
  AOI21_X1 U7805 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(n6550), .A(n6549), .ZN(
        n8291) );
  OR2_X1 U7806 ( .A1(n6701), .A2(n8291), .ZN(n6552) );
  OR2_X1 U7807 ( .A1(n6733), .A2(n8222), .ZN(n6551) );
  NAND4_X1 U7808 ( .A1(n6554), .A2(n6553), .A3(n6552), .A4(n6551), .ZN(n9326)
         );
  NOR2_X1 U7809 ( .A1(n11105), .A2(n9326), .ZN(n8284) );
  NAND2_X1 U7810 ( .A1(n11105), .A2(n9326), .ZN(n6555) );
  NAND2_X1 U7811 ( .A1(n7282), .A2(n6499), .ZN(n6560) );
  NAND2_X1 U7812 ( .A1(n6557), .A2(n6556), .ZN(n6558) );
  XNOR2_X1 U7813 ( .A(n6626), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8605) );
  AOI22_X1 U7814 ( .A1(n6642), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6641), .B2(
        n8605), .ZN(n6559) );
  NAND2_X1 U7815 ( .A1(n6560), .A2(n6559), .ZN(n11124) );
  NAND2_X1 U7816 ( .A1(n5121), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6565) );
  INV_X1 U7817 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8506) );
  OR2_X1 U7818 ( .A1(n9091), .A2(n8506), .ZN(n6564) );
  AOI21_X1 U7819 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(n6561), .A(n6571), .ZN(
        n8332) );
  OR2_X1 U7820 ( .A1(n6701), .A2(n8332), .ZN(n6563) );
  INV_X1 U7821 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8507) );
  OR2_X1 U7822 ( .A1(n6733), .A2(n8507), .ZN(n6562) );
  NAND2_X1 U7823 ( .A1(n11124), .A2(n8414), .ZN(n9199) );
  NAND2_X1 U7824 ( .A1(n9195), .A2(n9199), .ZN(n8335) );
  INV_X1 U7825 ( .A(n8414), .ZN(n9325) );
  NAND2_X1 U7826 ( .A1(n11124), .A2(n9325), .ZN(n6566) );
  INV_X1 U7827 ( .A(n8412), .ZN(n6580) );
  NAND2_X1 U7828 ( .A1(n7295), .A2(n6499), .ZN(n6570) );
  NAND2_X1 U7829 ( .A1(n6626), .A2(n6567), .ZN(n6568) );
  NAND2_X1 U7830 ( .A1(n6568), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6582) );
  XNOR2_X1 U7831 ( .A(n6582), .B(n6581), .ZN(n9347) );
  INV_X1 U7832 ( .A(n9347), .ZN(n8603) );
  AOI22_X1 U7833 ( .A1(n6642), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6641), .B2(
        n8603), .ZN(n6569) );
  NAND2_X1 U7834 ( .A1(n6570), .A2(n6569), .ZN(n8415) );
  NAND2_X1 U7835 ( .A1(n5121), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6578) );
  OAI21_X1 U7836 ( .B1(n9348), .B2(n6571), .A(n6586), .ZN(n6572) );
  INV_X1 U7837 ( .A(n6572), .ZN(n8416) );
  OR2_X1 U7838 ( .A1(n6701), .A2(n8416), .ZN(n6577) );
  INV_X1 U7839 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6573) );
  OR2_X1 U7840 ( .A1(n9091), .A2(n6573), .ZN(n6576) );
  INV_X1 U7841 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6574) );
  OR2_X1 U7842 ( .A1(n6733), .A2(n6574), .ZN(n6575) );
  OR2_X1 U7843 ( .A1(n8415), .A2(n8463), .ZN(n9189) );
  NAND2_X1 U7844 ( .A1(n8415), .A2(n8463), .ZN(n8398) );
  NAND2_X1 U7845 ( .A1(n7388), .A2(n6499), .ZN(n6585) );
  NAND2_X1 U7846 ( .A1(n6582), .A2(n6581), .ZN(n6583) );
  NAND2_X1 U7847 ( .A1(n6583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6594) );
  XNOR2_X1 U7848 ( .A(n6594), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9371) );
  AOI22_X1 U7849 ( .A1(n6642), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6641), .B2(
        n9371), .ZN(n6584) );
  NAND2_X1 U7850 ( .A1(n5121), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6590) );
  INV_X1 U7851 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8599) );
  OR2_X1 U7852 ( .A1(n9091), .A2(n8599), .ZN(n6589) );
  INV_X1 U7853 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8600) );
  OR2_X1 U7854 ( .A1(n6733), .A2(n8600), .ZN(n6588) );
  AOI21_X1 U7855 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(n6586), .A(n6598), .ZN(
        n8466) );
  OR2_X1 U7856 ( .A1(n6701), .A2(n8466), .ZN(n6587) );
  NAND2_X1 U7857 ( .A1(n11138), .A2(n8467), .ZN(n9203) );
  NAND2_X1 U7858 ( .A1(n9201), .A2(n9203), .ZN(n9191) );
  INV_X1 U7859 ( .A(n8463), .ZN(n9324) );
  OR2_X1 U7860 ( .A1(n8415), .A2(n9324), .ZN(n8400) );
  AND2_X1 U7861 ( .A1(n9191), .A2(n8400), .ZN(n6591) );
  NAND2_X1 U7862 ( .A1(n8410), .A2(n6591), .ZN(n8402) );
  INV_X1 U7863 ( .A(n8467), .ZN(n9323) );
  NAND2_X1 U7864 ( .A1(n11138), .A2(n9323), .ZN(n6592) );
  NAND2_X1 U7865 ( .A1(n8402), .A2(n6592), .ZN(n8454) );
  NAND2_X1 U7866 ( .A1(n7629), .A2(n6499), .ZN(n6597) );
  NAND2_X1 U7867 ( .A1(n6594), .A2(n6593), .ZN(n6595) );
  NAND2_X1 U7868 ( .A1(n6595), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6610) );
  XNOR2_X1 U7869 ( .A(n6610), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8613) );
  AOI22_X1 U7870 ( .A1(n6642), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8613), .B2(
        n6641), .ZN(n6596) );
  OR2_X1 U7871 ( .A1(n6598), .A2(n9381), .ZN(n6599) );
  NAND2_X1 U7872 ( .A1(n6599), .A2(n6617), .ZN(n8558) );
  NAND2_X1 U7873 ( .A1(n6600), .A2(n8558), .ZN(n6606) );
  INV_X1 U7874 ( .A(n5121), .ZN(n6748) );
  INV_X1 U7875 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6602) );
  OR2_X1 U7876 ( .A1(n6748), .A2(n6602), .ZN(n6605) );
  INV_X1 U7877 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8592) );
  OR2_X1 U7878 ( .A1(n9091), .A2(n8592), .ZN(n6604) );
  INV_X1 U7879 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8459) );
  OR2_X1 U7880 ( .A1(n6733), .A2(n8459), .ZN(n6603) );
  NAND2_X1 U7881 ( .A1(n11144), .A2(n8539), .ZN(n9204) );
  NAND2_X1 U7882 ( .A1(n9205), .A2(n9204), .ZN(n9292) );
  NAND2_X1 U7883 ( .A1(n8454), .A2(n9292), .ZN(n6608) );
  INV_X1 U7884 ( .A(n8539), .ZN(n9322) );
  NAND2_X1 U7885 ( .A1(n11144), .A2(n9322), .ZN(n6607) );
  NAND2_X1 U7886 ( .A1(n6608), .A2(n6607), .ZN(n8486) );
  NAND2_X1 U7887 ( .A1(n7649), .A2(n6499), .ZN(n6614) );
  INV_X1 U7888 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U7889 ( .A1(n6610), .A2(n6609), .ZN(n6611) );
  NAND2_X1 U7890 ( .A1(n6611), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6612) );
  XNOR2_X1 U7891 ( .A(n6612), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8618) );
  AOI22_X1 U7892 ( .A1(n8618), .A2(n6641), .B1(n6642), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6613) );
  NAND2_X1 U7893 ( .A1(n5121), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6621) );
  OR2_X1 U7894 ( .A1(n9091), .A2(n11152), .ZN(n6620) );
  INV_X1 U7895 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n6615) );
  OR2_X1 U7896 ( .A1(n6733), .A2(n6615), .ZN(n6619) );
  AOI21_X1 U7897 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n6617), .A(n6616), .ZN(
        n8546) );
  OR2_X1 U7898 ( .A1(n6701), .A2(n8546), .ZN(n6618) );
  OR2_X1 U7899 ( .A1(n11150), .A2(n8542), .ZN(n9214) );
  NAND2_X1 U7900 ( .A1(n11150), .A2(n8542), .ZN(n9213) );
  NAND2_X1 U7901 ( .A1(n9214), .A2(n9213), .ZN(n8487) );
  NAND2_X1 U7902 ( .A1(n8486), .A2(n8487), .ZN(n6623) );
  INV_X1 U7903 ( .A(n8542), .ZN(n9321) );
  NAND2_X1 U7904 ( .A1(n11150), .A2(n9321), .ZN(n6622) );
  NAND2_X1 U7905 ( .A1(n6623), .A2(n6622), .ZN(n8522) );
  NAND2_X1 U7906 ( .A1(n7741), .A2(n6499), .ZN(n6629) );
  NAND2_X1 U7907 ( .A1(n6624), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6625) );
  INV_X1 U7908 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6627) );
  XNOR2_X1 U7909 ( .A(n6640), .B(n6627), .ZN(n8595) );
  AOI22_X1 U7910 ( .A1(n6642), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6641), .B2(
        n8595), .ZN(n6628) );
  INV_X1 U7911 ( .A(n9091), .ZN(n6783) );
  NAND2_X1 U7912 ( .A1(n6783), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6636) );
  INV_X1 U7913 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6630) );
  OR2_X1 U7914 ( .A1(n6748), .A2(n6630), .ZN(n6635) );
  AND2_X1 U7915 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(n6631), .ZN(n6632) );
  NOR2_X1 U7916 ( .A1(n6646), .A2(n6632), .ZN(n8571) );
  OR2_X1 U7917 ( .A1(n6701), .A2(n8571), .ZN(n6634) );
  INV_X1 U7918 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8526) );
  OR2_X1 U7919 ( .A1(n6733), .A2(n8526), .ZN(n6633) );
  NAND4_X1 U7920 ( .A1(n6636), .A2(n6635), .A3(n6634), .A4(n6633), .ZN(n9320)
         );
  OR2_X1 U7921 ( .A1(n10032), .A2(n9320), .ZN(n6637) );
  NAND2_X1 U7922 ( .A1(n8522), .A2(n6637), .ZN(n6639) );
  NAND2_X1 U7923 ( .A1(n10032), .A2(n9320), .ZN(n6638) );
  NAND2_X1 U7924 ( .A1(n6639), .A2(n6638), .ZN(n9977) );
  NAND2_X1 U7925 ( .A1(n7911), .A2(n6499), .ZN(n6644) );
  AOI22_X1 U7926 ( .A1(n6642), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9424), .B2(
        n6641), .ZN(n6643) );
  NAND2_X1 U7927 ( .A1(n5121), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6653) );
  INV_X1 U7928 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n6645) );
  OR2_X1 U7929 ( .A1(n9091), .A2(n6645), .ZN(n6652) );
  NOR2_X1 U7930 ( .A1(n6646), .A2(n9518), .ZN(n6647) );
  OR2_X1 U7931 ( .A1(n6658), .A2(n6647), .ZN(n9982) );
  INV_X1 U7932 ( .A(n9982), .ZN(n6648) );
  OR2_X1 U7933 ( .A1(n6701), .A2(n6648), .ZN(n6651) );
  INV_X1 U7934 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6649) );
  OR2_X1 U7935 ( .A1(n6733), .A2(n6649), .ZN(n6650) );
  NAND2_X1 U7936 ( .A1(n10028), .A2(n8954), .ZN(n9967) );
  NAND2_X1 U7937 ( .A1(n9221), .A2(n9967), .ZN(n9980) );
  NAND2_X1 U7938 ( .A1(n9977), .A2(n9980), .ZN(n9976) );
  NAND2_X1 U7939 ( .A1(n10028), .A2(n9962), .ZN(n6654) );
  NAND2_X1 U7940 ( .A1(n8013), .A2(n6499), .ZN(n6656) );
  OR2_X1 U7941 ( .A1(n9101), .A2(n8014), .ZN(n6655) );
  NAND2_X1 U7942 ( .A1(n5121), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6663) );
  INV_X1 U7943 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6657) );
  OR2_X1 U7944 ( .A1(n9091), .A2(n6657), .ZN(n6662) );
  NOR2_X1 U7945 ( .A1(n6658), .A2(n9535), .ZN(n6659) );
  OR2_X1 U7946 ( .A1(n6669), .A2(n6659), .ZN(n9966) );
  INV_X1 U7947 ( .A(n9966), .ZN(n9057) );
  OR2_X1 U7948 ( .A1(n6701), .A2(n9057), .ZN(n6661) );
  INV_X1 U7949 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9971) );
  OR2_X1 U7950 ( .A1(n6733), .A2(n9971), .ZN(n6660) );
  NAND4_X1 U7951 ( .A1(n6663), .A2(n6662), .A3(n6661), .A4(n6660), .ZN(n9946)
         );
  NAND2_X1 U7952 ( .A1(n9972), .A2(n9946), .ZN(n9223) );
  INV_X1 U7953 ( .A(n9946), .ZN(n8957) );
  NAND2_X1 U7954 ( .A1(n10024), .A2(n8957), .ZN(n9225) );
  NAND2_X1 U7955 ( .A1(n9972), .A2(n8957), .ZN(n6665) );
  NAND2_X1 U7956 ( .A1(n8179), .A2(n6499), .ZN(n6667) );
  INV_X1 U7957 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8181) );
  OR2_X1 U7958 ( .A1(n9101), .A2(n8181), .ZN(n6666) );
  NAND2_X1 U7959 ( .A1(n6783), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6674) );
  INV_X1 U7960 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6668) );
  OR2_X1 U7961 ( .A1(n6748), .A2(n6668), .ZN(n6673) );
  OR2_X1 U7962 ( .A1(n6669), .A2(n9027), .ZN(n6670) );
  AND2_X1 U7963 ( .A1(n6670), .A2(n6678), .ZN(n9949) );
  OR2_X1 U7964 ( .A1(n6701), .A2(n9949), .ZN(n6672) );
  INV_X1 U7965 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9950) );
  OR2_X1 U7966 ( .A1(n6733), .A2(n9950), .ZN(n6671) );
  NAND2_X1 U7967 ( .A1(n10020), .A2(n9068), .ZN(n9227) );
  NAND2_X1 U7968 ( .A1(n9226), .A2(n9227), .ZN(n9944) );
  NAND2_X1 U7969 ( .A1(n8236), .A2(n6499), .ZN(n6676) );
  INV_X1 U7970 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8238) );
  OR2_X1 U7971 ( .A1(n9101), .A2(n8238), .ZN(n6675) );
  NAND2_X1 U7972 ( .A1(n5121), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6683) );
  INV_X1 U7973 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6677) );
  OR2_X1 U7974 ( .A1(n9091), .A2(n6677), .ZN(n6682) );
  NAND2_X1 U7975 ( .A1(n6678), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6679) );
  AND2_X1 U7976 ( .A1(n6689), .A2(n6679), .ZN(n9936) );
  OR2_X1 U7977 ( .A1(n6701), .A2(n9936), .ZN(n6681) );
  INV_X1 U7978 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9937) );
  OR2_X1 U7979 ( .A1(n6733), .A2(n9937), .ZN(n6680) );
  XNOR2_X1 U7980 ( .A(n10016), .B(n9230), .ZN(n9932) );
  NAND2_X1 U7981 ( .A1(n9933), .A2(n9932), .ZN(n6685) );
  OR2_X1 U7982 ( .A1(n10016), .A2(n9947), .ZN(n6684) );
  NAND2_X1 U7983 ( .A1(n8265), .A2(n6499), .ZN(n6687) );
  OR2_X1 U7984 ( .A1(n9101), .A2(n8268), .ZN(n6686) );
  NAND2_X1 U7985 ( .A1(n5121), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6695) );
  INV_X1 U7986 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6688) );
  OR2_X1 U7987 ( .A1(n9091), .A2(n6688), .ZN(n6694) );
  AND2_X1 U7988 ( .A1(n6689), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6690) );
  NOR2_X1 U7989 ( .A1(n6699), .A2(n6690), .ZN(n9010) );
  OR2_X1 U7990 ( .A1(n6701), .A2(n9010), .ZN(n6693) );
  INV_X1 U7991 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n6691) );
  OR2_X1 U7992 ( .A1(n6733), .A2(n6691), .ZN(n6692) );
  NAND4_X2 U7993 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n9934)
         );
  NAND2_X1 U7994 ( .A1(n8372), .A2(n6499), .ZN(n6697) );
  OR2_X1 U7995 ( .A1(n9101), .A2(n8986), .ZN(n6696) );
  NAND2_X1 U7996 ( .A1(n5121), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6706) );
  INV_X1 U7997 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6698) );
  OR2_X1 U7998 ( .A1(n9091), .A2(n6698), .ZN(n6705) );
  NOR2_X1 U7999 ( .A1(n6699), .A2(n9540), .ZN(n6700) );
  OR2_X1 U8000 ( .A1(n6712), .A2(n6700), .ZN(n9918) );
  INV_X1 U8001 ( .A(n9918), .ZN(n9048) );
  OR2_X1 U8002 ( .A1(n6701), .A2(n9048), .ZN(n6704) );
  INV_X1 U8003 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6702) );
  OR2_X1 U8004 ( .A1(n6733), .A2(n6702), .ZN(n6703) );
  NAND4_X1 U8005 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .ZN(n9923)
         );
  NAND2_X1 U8006 ( .A1(n10008), .A2(n9923), .ZN(n6708) );
  NOR2_X1 U8007 ( .A1(n10008), .A2(n9923), .ZN(n6707) );
  NAND2_X1 U8008 ( .A1(n8450), .A2(n6499), .ZN(n6710) );
  INV_X1 U8009 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8932) );
  OR2_X1 U8010 ( .A1(n9101), .A2(n8932), .ZN(n6709) );
  NAND2_X1 U8011 ( .A1(n5121), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6718) );
  INV_X1 U8012 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6711) );
  OR2_X1 U8013 ( .A1(n9091), .A2(n6711), .ZN(n6717) );
  OR2_X1 U8014 ( .A1(n6712), .A2(n9735), .ZN(n6713) );
  AND2_X1 U8015 ( .A1(n6722), .A2(n6713), .ZN(n9907) );
  OR2_X1 U8016 ( .A1(n6701), .A2(n9907), .ZN(n6716) );
  INV_X1 U8017 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6714) );
  OR2_X1 U8018 ( .A1(n6733), .A2(n6714), .ZN(n6715) );
  NAND2_X1 U8019 ( .A1(n9906), .A2(n8971), .ZN(n9245) );
  NAND2_X1 U8020 ( .A1(n8476), .A2(n6499), .ZN(n6720) );
  OR2_X1 U8021 ( .A1(n9101), .A2(n8478), .ZN(n6719) );
  NAND2_X1 U8022 ( .A1(n5121), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6726) );
  INV_X1 U8023 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6721) );
  OR2_X1 U8024 ( .A1(n9091), .A2(n6721), .ZN(n6725) );
  INV_X1 U8025 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9762) );
  XNOR2_X1 U8026 ( .A(n6722), .B(n9762), .ZN(n9889) );
  OR2_X1 U8027 ( .A1(n6701), .A2(n9889), .ZN(n6724) );
  INV_X1 U8028 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9890) );
  OR2_X1 U8029 ( .A1(n6733), .A2(n9890), .ZN(n6723) );
  XNOR2_X1 U8030 ( .A(n10000), .B(n9251), .ZN(n9887) );
  INV_X1 U8031 ( .A(n10000), .ZN(n9089) );
  OR2_X1 U8032 ( .A1(n9996), .A2(n9079), .ZN(n9259) );
  NAND2_X1 U8033 ( .A1(n9996), .A2(n9079), .ZN(n9254) );
  NAND2_X1 U8034 ( .A1(n9259), .A2(n9254), .ZN(n9883) );
  NAND2_X1 U8035 ( .A1(n8532), .A2(n6499), .ZN(n6729) );
  INV_X1 U8036 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6727) );
  OR2_X1 U8037 ( .A1(n9101), .A2(n6727), .ZN(n6728) );
  NAND2_X1 U8038 ( .A1(n6783), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6737) );
  INV_X1 U8039 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6730) );
  OR2_X1 U8040 ( .A1(n6748), .A2(n6730), .ZN(n6736) );
  INV_X1 U8041 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9522) );
  NOR2_X1 U8042 ( .A1(n6731), .A2(n9522), .ZN(n6732) );
  NOR2_X1 U8043 ( .A1(n9433), .A2(n6732), .ZN(n9445) );
  OR2_X1 U8044 ( .A1(n6701), .A2(n9445), .ZN(n6735) );
  INV_X1 U8045 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9446) );
  OR2_X1 U8046 ( .A1(n6733), .A2(n9446), .ZN(n6734) );
  OAI22_X1 U8047 ( .A1(n9440), .A2(n9448), .B1(n9874), .B2(n9992), .ZN(n6752)
         );
  INV_X1 U8048 ( .A(n6740), .ZN(n6741) );
  INV_X1 U8049 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6742) );
  INV_X1 U8050 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9760) );
  MUX2_X1 U8051 ( .A(n6742), .B(n9760), .S(n7159), .Z(n8637) );
  NAND2_X1 U8052 ( .A1(n8762), .A2(n6499), .ZN(n6744) );
  OR2_X1 U8053 ( .A1(n9101), .A2(n6742), .ZN(n6743) );
  INV_X1 U8054 ( .A(n9433), .ZN(n6745) );
  OR2_X1 U8055 ( .A1(n6701), .A2(n6745), .ZN(n9096) );
  NAND2_X1 U8056 ( .A1(n6783), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6751) );
  INV_X1 U8057 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6746) );
  OR2_X1 U8058 ( .A1(n6733), .A2(n6746), .ZN(n6750) );
  INV_X1 U8059 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6747) );
  OR2_X1 U8060 ( .A1(n6748), .A2(n6747), .ZN(n6749) );
  NAND4_X1 U8061 ( .A1(n9096), .A2(n6751), .A3(n6750), .A4(n6749), .ZN(n9441)
         );
  XNOR2_X1 U8062 ( .A(n6797), .B(n9441), .ZN(n6778) );
  XNOR2_X1 U8063 ( .A(n6755), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7342) );
  INV_X1 U8064 ( .A(n9268), .ZN(n6800) );
  NAND2_X1 U8065 ( .A1(n7342), .A2(n6800), .ZN(n9104) );
  NAND2_X1 U8066 ( .A1(n6813), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U8067 ( .A1(n9424), .A2(n9313), .ZN(n7138) );
  INV_X1 U8068 ( .A(n9270), .ZN(n8067) );
  INV_X1 U8069 ( .A(n10938), .ZN(n7560) );
  OR2_X1 U8070 ( .A1(n9337), .A2(n7560), .ZN(n9121) );
  INV_X1 U8071 ( .A(n9121), .ZN(n8066) );
  NAND2_X1 U8072 ( .A1(n8067), .A2(n8066), .ZN(n8065) );
  NAND2_X1 U8073 ( .A1(n8065), .A2(n9125), .ZN(n10962) );
  INV_X1 U8074 ( .A(n9272), .ZN(n10966) );
  NAND2_X1 U8075 ( .A1(n10962), .A2(n10966), .ZN(n7973) );
  AND2_X1 U8076 ( .A1(n9133), .A2(n9142), .ZN(n6759) );
  NAND2_X1 U8077 ( .A1(n7973), .A2(n6759), .ZN(n6762) );
  INV_X1 U8078 ( .A(n9142), .ZN(n6760) );
  INV_X1 U8079 ( .A(n7975), .ZN(n9275) );
  OR2_X1 U8080 ( .A1(n6760), .A2(n9275), .ZN(n6761) );
  INV_X1 U8081 ( .A(n7635), .ZN(n10988) );
  NAND2_X1 U8082 ( .A1(n9333), .A2(n10988), .ZN(n9140) );
  NAND2_X1 U8083 ( .A1(n7877), .A2(n9140), .ZN(n6763) );
  OR2_X1 U8084 ( .A1(n9333), .A2(n10988), .ZN(n9146) );
  INV_X1 U8085 ( .A(n7617), .ZN(n11004) );
  OR2_X1 U8086 ( .A1(n9332), .A2(n11004), .ZN(n9147) );
  NAND2_X1 U8087 ( .A1(n9332), .A2(n11004), .ZN(n9143) );
  NAND2_X1 U8088 ( .A1(n9147), .A2(n9143), .ZN(n9277) );
  INV_X1 U8089 ( .A(n9277), .ZN(n8081) );
  NAND2_X1 U8090 ( .A1(n8082), .A2(n8081), .ZN(n8080) );
  NAND2_X1 U8091 ( .A1(n8080), .A2(n9147), .ZN(n7713) );
  INV_X1 U8092 ( .A(n9278), .ZN(n7712) );
  AND2_X1 U8093 ( .A1(n9153), .A2(n7961), .ZN(n9170) );
  NAND2_X1 U8094 ( .A1(n7900), .A2(n9170), .ZN(n6764) );
  INV_X1 U8095 ( .A(n9328), .ZN(n8132) );
  OR2_X1 U8096 ( .A1(n11075), .A2(n8132), .ZN(n9177) );
  AND2_X1 U8097 ( .A1(n9177), .A2(n9154), .ZN(n9169) );
  INV_X1 U8098 ( .A(n9327), .ZN(n8279) );
  NAND2_X1 U8099 ( .A1(n11078), .A2(n8279), .ZN(n9178) );
  NAND2_X1 U8100 ( .A1(n11075), .A2(n8132), .ZN(n9166) );
  AND2_X1 U8101 ( .A1(n9178), .A2(n9166), .ZN(n9182) );
  NAND2_X1 U8102 ( .A1(n8061), .A2(n9182), .ZN(n6766) );
  OR2_X1 U8103 ( .A1(n11078), .A2(n8279), .ZN(n9180) );
  NOR2_X1 U8104 ( .A1(n11105), .A2(n8331), .ZN(n9119) );
  NAND2_X1 U8105 ( .A1(n11105), .A2(n8331), .ZN(n8286) );
  NAND2_X1 U8106 ( .A1(n8418), .A2(n9196), .ZN(n8397) );
  AND2_X1 U8107 ( .A1(n9203), .A2(n8398), .ZN(n9197) );
  NAND2_X1 U8108 ( .A1(n8397), .A2(n9197), .ZN(n6769) );
  NAND2_X1 U8109 ( .A1(n6769), .A2(n9201), .ZN(n8453) );
  INV_X1 U8110 ( .A(n9292), .ZN(n9193) );
  NAND2_X1 U8111 ( .A1(n8453), .A2(n9193), .ZN(n6770) );
  INV_X1 U8112 ( .A(n9214), .ZN(n6771) );
  NAND2_X1 U8113 ( .A1(n10032), .A2(n8950), .ZN(n9116) );
  AND2_X2 U8114 ( .A1(n8529), .A2(n9118), .ZN(n9981) );
  NAND2_X1 U8115 ( .A1(n9981), .A2(n9221), .ZN(n9968) );
  AND2_X1 U8116 ( .A1(n9225), .A2(n9967), .ZN(n9220) );
  NAND2_X1 U8117 ( .A1(n9968), .A2(n9220), .ZN(n6772) );
  INV_X1 U8118 ( .A(n9932), .ZN(n9939) );
  OR2_X1 U8119 ( .A1(n10016), .A2(n9230), .ZN(n9232) );
  NAND2_X1 U8120 ( .A1(n9938), .A2(n9232), .ZN(n9926) );
  INV_X1 U8121 ( .A(n9934), .ZN(n6773) );
  NOR2_X1 U8122 ( .A1(n10012), .A2(n6773), .ZN(n9236) );
  INV_X1 U8123 ( .A(n9923), .ZN(n8967) );
  OR2_X1 U8124 ( .A1(n10008), .A2(n8967), .ZN(n9240) );
  NAND2_X1 U8125 ( .A1(n10008), .A2(n8967), .ZN(n9239) );
  NAND2_X1 U8126 ( .A1(n9898), .A2(n9246), .ZN(n9892) );
  OR2_X1 U8127 ( .A1(n10000), .A2(n9251), .ZN(n6775) );
  AND2_X2 U8128 ( .A1(n9880), .A2(n9254), .ZN(n9449) );
  NAND2_X1 U8129 ( .A1(n9449), .A2(n9448), .ZN(n9447) );
  INV_X1 U8130 ( .A(n9874), .ZN(n6792) );
  OR2_X1 U8131 ( .A1(n9992), .A2(n6792), .ZN(n6776) );
  NAND2_X1 U8132 ( .A1(n9447), .A2(n6776), .ZN(n6779) );
  INV_X1 U8133 ( .A(n6779), .ZN(n6777) );
  NAND2_X1 U8134 ( .A1(n6777), .A2(n6778), .ZN(n9112) );
  NAND2_X1 U8135 ( .A1(n6779), .A2(n5297), .ZN(n6780) );
  NAND2_X1 U8136 ( .A1(n9112), .A2(n6780), .ZN(n8990) );
  AOI21_X1 U8137 ( .B1(n6800), .B2(n8237), .A(n9424), .ZN(n6781) );
  AND2_X1 U8138 ( .A1(n11127), .A2(n6781), .ZN(n6782) );
  NAND2_X1 U8139 ( .A1(n8990), .A2(n8157), .ZN(n6795) );
  NAND2_X1 U8140 ( .A1(n5121), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6787) );
  NAND2_X1 U8141 ( .A1(n6783), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8142 ( .A1(n6784), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6785) );
  INV_X1 U8143 ( .A(n6788), .ZN(n6790) );
  AND2_X1 U8144 ( .A1(n7153), .A2(P2_B_REG_SCAN_IN), .ZN(n6791) );
  OR2_X1 U8145 ( .A1(n8523), .A2(n6791), .ZN(n9434) );
  INV_X1 U8146 ( .A(n9875), .ZN(n9902) );
  OAI22_X1 U8147 ( .A1(n9106), .A2(n9434), .B1(n6792), .B2(n8524), .ZN(n6793)
         );
  INV_X1 U8148 ( .A(n6793), .ZN(n6794) );
  NAND2_X1 U8149 ( .A1(n6795), .A2(n6794), .ZN(n6796) );
  NAND2_X1 U8150 ( .A1(n9268), .A2(n9424), .ZN(n7143) );
  OR2_X1 U8151 ( .A1(n7143), .A2(n9313), .ZN(n11071) );
  NAND2_X1 U8152 ( .A1(n8990), .A2(n11008), .ZN(n6798) );
  INV_X1 U8153 ( .A(n6797), .ZN(n8992) );
  INV_X1 U8154 ( .A(n7344), .ZN(n6799) );
  NAND3_X1 U8155 ( .A1(n6800), .A2(n9313), .A3(n9409), .ZN(n6801) );
  NAND2_X1 U8156 ( .A1(n9244), .A2(n6801), .ZN(n7760) );
  NAND2_X1 U8157 ( .A1(n7759), .A2(n7760), .ZN(n6821) );
  NAND2_X1 U8158 ( .A1(n6841), .A2(n6842), .ZN(n6805) );
  XNOR2_X1 U8159 ( .A(n6819), .B(P2_B_REG_SCAN_IN), .ZN(n6811) );
  NAND2_X1 U8160 ( .A1(n6807), .A2(n6806), .ZN(n6808) );
  NAND2_X1 U8161 ( .A1(n6811), .A2(n6823), .ZN(n6818) );
  OR2_X1 U8162 ( .A1(n6813), .A2(n6812), .ZN(n6814) );
  NAND2_X1 U8163 ( .A1(n6814), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6815) );
  MUX2_X1 U8164 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6815), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6817) );
  INV_X1 U8165 ( .A(n6838), .ZN(n8477) );
  NAND2_X1 U8166 ( .A1(n6819), .A2(n8477), .ZN(n7257) );
  NAND2_X1 U8167 ( .A1(n6820), .A2(n7257), .ZN(n7339) );
  NAND2_X1 U8168 ( .A1(n6821), .A2(n7339), .ZN(n6844) );
  OR2_X1 U8169 ( .A1(n6822), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U8170 ( .A1(n6823), .A2(n8477), .ZN(n6824) );
  NOR2_X1 U8171 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6829) );
  NOR4_X1 U8172 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6828) );
  NOR4_X1 U8173 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6827) );
  NOR4_X1 U8174 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6826) );
  NAND4_X1 U8175 ( .A1(n6829), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(n6835)
         );
  NOR4_X1 U8176 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6833) );
  NOR4_X1 U8177 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6832) );
  NOR4_X1 U8178 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6831) );
  NOR4_X1 U8179 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6830) );
  NAND4_X1 U8180 ( .A1(n6833), .A2(n6832), .A3(n6831), .A4(n6830), .ZN(n6834)
         );
  NOR2_X1 U8181 ( .A1(n6835), .A2(n6834), .ZN(n6836) );
  INV_X1 U8182 ( .A(n6819), .ZN(n6837) );
  AND2_X1 U8183 ( .A1(n7145), .A2(n7192), .ZN(n6843) );
  NAND2_X1 U8184 ( .A1(n7760), .A2(n7761), .ZN(n7763) );
  OR2_X1 U8185 ( .A1(n11071), .A2(n7342), .ZN(n10942) );
  INV_X2 U8186 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U8187 ( .A(n7577), .ZN(n6846) );
  NAND2_X1 U8188 ( .A1(n6848), .A2(n7577), .ZN(n6849) );
  NAND2_X1 U8189 ( .A1(n6852), .A2(n6849), .ZN(n6850) );
  NAND2_X2 U8190 ( .A1(n6854), .A2(n6850), .ZN(n7059) );
  AND2_X1 U8191 ( .A1(n10433), .A2(n7118), .ZN(n6851) );
  AOI21_X1 U8192 ( .B1(n10405), .B2(n7072), .A(n6851), .ZN(n7062) );
  INV_X1 U8193 ( .A(n7062), .ZN(n7064) );
  NAND2_X1 U8194 ( .A1(n10405), .A2(n7123), .ZN(n6856) );
  NAND2_X1 U8195 ( .A1(n10433), .A2(n7117), .ZN(n6855) );
  NAND2_X1 U8196 ( .A1(n6856), .A2(n6855), .ZN(n6857) );
  XNOR2_X1 U8197 ( .A(n6857), .B(n5119), .ZN(n7063) );
  NAND2_X1 U8198 ( .A1(n6900), .A2(n6858), .ZN(n6860) );
  NAND2_X1 U8199 ( .A1(n6887), .A2(n10932), .ZN(n6859) );
  INV_X1 U8200 ( .A(n7059), .ZN(n6862) );
  INV_X1 U8201 ( .A(n6847), .ZN(n6863) );
  NAND2_X1 U8202 ( .A1(n6863), .A2(n10752), .ZN(n6864) );
  OAI211_X1 U8203 ( .C1(n7060), .C2(n7570), .A(n6865), .B(n6864), .ZN(n7285)
         );
  NAND2_X1 U8204 ( .A1(n7284), .A2(n7285), .ZN(n7287) );
  OR2_X1 U8205 ( .A1(n5119), .A2(n10932), .ZN(n6866) );
  NAND2_X1 U8206 ( .A1(n7287), .A2(n6866), .ZN(n6873) );
  NAND2_X1 U8207 ( .A1(n6887), .A2(n5122), .ZN(n6868) );
  NAND2_X1 U8208 ( .A1(n6900), .A2(n10214), .ZN(n6867) );
  NAND2_X1 U8209 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  NAND2_X1 U8210 ( .A1(n6873), .A2(n6872), .ZN(n7431) );
  INV_X1 U8211 ( .A(n10214), .ZN(n7304) );
  OR2_X1 U8212 ( .A1(n7304), .A2(n7059), .ZN(n6871) );
  OR2_X1 U8213 ( .A1(n7060), .A2(n8864), .ZN(n6870) );
  AND2_X1 U8214 ( .A1(n6871), .A2(n6870), .ZN(n7434) );
  NAND2_X1 U8215 ( .A1(n7431), .A2(n7434), .ZN(n6876) );
  INV_X1 U8216 ( .A(n6873), .ZN(n6874) );
  NAND2_X1 U8217 ( .A1(n6875), .A2(n6874), .ZN(n7433) );
  NAND2_X1 U8218 ( .A1(n6876), .A2(n7433), .ZN(n7439) );
  NAND2_X1 U8219 ( .A1(n6887), .A2(n7704), .ZN(n6878) );
  NAND2_X1 U8220 ( .A1(n6900), .A2(n10213), .ZN(n6877) );
  NAND2_X1 U8221 ( .A1(n6878), .A2(n6877), .ZN(n6879) );
  INV_X4 U8222 ( .A(n5119), .ZN(n7089) );
  INV_X1 U8223 ( .A(n10213), .ZN(n7461) );
  OR2_X1 U8224 ( .A1(n7060), .A2(n7335), .ZN(n6880) );
  NAND2_X1 U8225 ( .A1(n6881), .A2(n6880), .ZN(n6882) );
  XNOR2_X1 U8226 ( .A(n6884), .B(n6882), .ZN(n7440) );
  NAND2_X1 U8227 ( .A1(n7439), .A2(n7440), .ZN(n6886) );
  INV_X1 U8228 ( .A(n6882), .ZN(n6883) );
  NAND2_X1 U8229 ( .A1(n6884), .A2(n6883), .ZN(n6885) );
  NAND2_X1 U8230 ( .A1(n6886), .A2(n6885), .ZN(n7486) );
  NAND2_X1 U8231 ( .A1(n6887), .A2(n7773), .ZN(n6889) );
  NAND2_X1 U8232 ( .A1(n6900), .A2(n10212), .ZN(n6888) );
  NAND2_X1 U8233 ( .A1(n6889), .A2(n6888), .ZN(n6890) );
  NAND2_X1 U8234 ( .A1(n7118), .A2(n10212), .ZN(n6892) );
  NAND2_X1 U8235 ( .A1(n6900), .A2(n7773), .ZN(n6891) );
  AND2_X1 U8236 ( .A1(n6892), .A2(n6891), .ZN(n6894) );
  XNOR2_X1 U8237 ( .A(n6893), .B(n6894), .ZN(n7488) );
  INV_X1 U8238 ( .A(n6893), .ZN(n6895) );
  NAND2_X1 U8239 ( .A1(n6895), .A2(n6894), .ZN(n6896) );
  NAND2_X1 U8240 ( .A1(n6887), .A2(n10995), .ZN(n6898) );
  NAND2_X1 U8241 ( .A1(n6900), .A2(n10211), .ZN(n6897) );
  NAND2_X1 U8242 ( .A1(n6898), .A2(n6897), .ZN(n6899) );
  NAND2_X1 U8243 ( .A1(n7118), .A2(n10211), .ZN(n6902) );
  NAND2_X1 U8244 ( .A1(n6900), .A2(n10995), .ZN(n6901) );
  AND2_X1 U8245 ( .A1(n6902), .A2(n6901), .ZN(n6905) );
  XNOR2_X1 U8246 ( .A(n6904), .B(n6905), .ZN(n7498) );
  INV_X1 U8247 ( .A(n6904), .ZN(n6907) );
  INV_X1 U8248 ( .A(n6905), .ZN(n6906) );
  NAND2_X1 U8249 ( .A1(n6907), .A2(n6906), .ZN(n6908) );
  NAND2_X1 U8250 ( .A1(n7496), .A2(n6908), .ZN(n6914) );
  NAND2_X1 U8251 ( .A1(n7123), .A2(n11017), .ZN(n6910) );
  NAND2_X1 U8252 ( .A1(n7117), .A2(n10210), .ZN(n6909) );
  NAND2_X1 U8253 ( .A1(n6910), .A2(n6909), .ZN(n6911) );
  XNOR2_X1 U8254 ( .A(n6911), .B(n5119), .ZN(n6915) );
  NAND2_X1 U8255 ( .A1(n6914), .A2(n6915), .ZN(n7503) );
  NAND2_X1 U8256 ( .A1(n11017), .A2(n7117), .ZN(n6913) );
  NAND2_X1 U8257 ( .A1(n7118), .A2(n10210), .ZN(n6912) );
  AND2_X1 U8258 ( .A1(n6913), .A2(n6912), .ZN(n7505) );
  NAND2_X1 U8259 ( .A1(n7503), .A2(n7505), .ZN(n6918) );
  INV_X1 U8260 ( .A(n6914), .ZN(n6917) );
  INV_X1 U8261 ( .A(n6915), .ZN(n6916) );
  NAND2_X1 U8262 ( .A1(n6917), .A2(n6916), .ZN(n7504) );
  NAND2_X1 U8263 ( .A1(n10166), .A2(n7123), .ZN(n6920) );
  NAND2_X1 U8264 ( .A1(n7117), .A2(n10209), .ZN(n6919) );
  NAND2_X1 U8265 ( .A1(n6920), .A2(n6919), .ZN(n6921) );
  XNOR2_X1 U8266 ( .A(n6921), .B(n7089), .ZN(n6923) );
  NOR2_X1 U8267 ( .A1(n7751), .A2(n7059), .ZN(n6922) );
  AOI21_X1 U8268 ( .B1(n10166), .B2(n7117), .A(n6922), .ZN(n6924) );
  AND2_X1 U8269 ( .A1(n6923), .A2(n6924), .ZN(n10163) );
  INV_X1 U8270 ( .A(n6923), .ZN(n6926) );
  INV_X1 U8271 ( .A(n6924), .ZN(n6925) );
  NAND2_X1 U8272 ( .A1(n6926), .A2(n6925), .ZN(n10162) );
  NAND2_X1 U8273 ( .A1(n7784), .A2(n6887), .ZN(n6928) );
  NAND2_X1 U8274 ( .A1(n7117), .A2(n10208), .ZN(n6927) );
  NAND2_X1 U8275 ( .A1(n6928), .A2(n6927), .ZN(n6929) );
  XNOR2_X1 U8276 ( .A(n6929), .B(n5119), .ZN(n7668) );
  INV_X1 U8277 ( .A(n7668), .ZN(n6932) );
  NAND2_X1 U8278 ( .A1(n7784), .A2(n7117), .ZN(n6931) );
  NAND2_X1 U8279 ( .A1(n7118), .A2(n10208), .ZN(n6930) );
  NAND2_X1 U8280 ( .A1(n6931), .A2(n6930), .ZN(n6936) );
  INV_X1 U8281 ( .A(n6936), .ZN(n7667) );
  NAND2_X1 U8282 ( .A1(n6932), .A2(n7667), .ZN(n6942) );
  NAND2_X1 U8283 ( .A1(n7866), .A2(n7123), .ZN(n6934) );
  NAND2_X1 U8284 ( .A1(n7117), .A2(n10207), .ZN(n6933) );
  NAND2_X1 U8285 ( .A1(n6934), .A2(n6933), .ZN(n6935) );
  XNOR2_X1 U8286 ( .A(n6935), .B(n5119), .ZN(n6941) );
  INV_X1 U8287 ( .A(n6941), .ZN(n6938) );
  AND2_X1 U8288 ( .A1(n7668), .A2(n6936), .ZN(n6943) );
  INV_X1 U8289 ( .A(n6943), .ZN(n6937) );
  NAND2_X1 U8290 ( .A1(n7866), .A2(n7117), .ZN(n6940) );
  NAND2_X1 U8291 ( .A1(n7118), .A2(n10207), .ZN(n6939) );
  NAND2_X1 U8292 ( .A1(n6940), .A2(n6939), .ZN(n7861) );
  NAND2_X1 U8293 ( .A1(n7858), .A2(n7861), .ZN(n6944) );
  OAI211_X2 U8294 ( .C1(n7670), .C2(n6943), .A(n6942), .B(n6941), .ZN(n7859)
         );
  NAND2_X1 U8295 ( .A1(n6944), .A2(n7859), .ZN(n7938) );
  INV_X1 U8296 ( .A(n7938), .ZN(n6950) );
  NAND2_X1 U8297 ( .A1(n7946), .A2(n7123), .ZN(n6946) );
  NAND2_X1 U8298 ( .A1(n7072), .A2(n10206), .ZN(n6945) );
  NAND2_X1 U8299 ( .A1(n6946), .A2(n6945), .ZN(n6947) );
  XNOR2_X1 U8300 ( .A(n6947), .B(n7089), .ZN(n6952) );
  NOR2_X1 U8301 ( .A1(n7863), .A2(n7059), .ZN(n6948) );
  AOI21_X1 U8302 ( .B1(n7946), .B2(n7072), .A(n6948), .ZN(n6951) );
  XNOR2_X1 U8303 ( .A(n6952), .B(n6951), .ZN(n7939) );
  NAND2_X1 U8304 ( .A1(n6950), .A2(n6949), .ZN(n7935) );
  NAND2_X1 U8305 ( .A1(n6952), .A2(n6951), .ZN(n6953) );
  NAND2_X1 U8306 ( .A1(n8175), .A2(n7123), .ZN(n6955) );
  NAND2_X1 U8307 ( .A1(n7072), .A2(n7916), .ZN(n6954) );
  NAND2_X1 U8308 ( .A1(n6955), .A2(n6954), .ZN(n6956) );
  XNOR2_X1 U8309 ( .A(n6956), .B(n5119), .ZN(n6958) );
  NOR2_X1 U8310 ( .A1(n11095), .A2(n7059), .ZN(n6957) );
  NAND2_X1 U8311 ( .A1(n11089), .A2(n7123), .ZN(n6960) );
  NAND2_X1 U8312 ( .A1(n7072), .A2(n10205), .ZN(n6959) );
  NAND2_X1 U8313 ( .A1(n6960), .A2(n6959), .ZN(n6961) );
  XNOR2_X1 U8314 ( .A(n6961), .B(n7089), .ZN(n6968) );
  NOR2_X1 U8315 ( .A1(n8172), .A2(n7059), .ZN(n6962) );
  AOI21_X1 U8316 ( .B1(n11089), .B2(n7072), .A(n6962), .ZN(n6969) );
  NAND2_X1 U8317 ( .A1(n6968), .A2(n6969), .ZN(n11085) );
  NAND2_X1 U8318 ( .A1(n11084), .A2(n11085), .ZN(n8270) );
  NAND2_X1 U8319 ( .A1(n7956), .A2(n7123), .ZN(n6964) );
  NAND2_X1 U8320 ( .A1(n7072), .A2(n11090), .ZN(n6963) );
  NAND2_X1 U8321 ( .A1(n6964), .A2(n6963), .ZN(n6965) );
  XNOR2_X1 U8322 ( .A(n6965), .B(n5119), .ZN(n6977) );
  NOR2_X1 U8323 ( .A1(n6966), .A2(n7059), .ZN(n6967) );
  AOI21_X1 U8324 ( .B1(n7956), .B2(n7072), .A(n6967), .ZN(n6978) );
  XNOR2_X1 U8325 ( .A(n6977), .B(n6978), .ZN(n8271) );
  INV_X1 U8326 ( .A(n6968), .ZN(n6971) );
  INV_X1 U8327 ( .A(n6969), .ZN(n6970) );
  NAND2_X1 U8328 ( .A1(n6971), .A2(n6970), .ZN(n11086) );
  AND2_X1 U8329 ( .A1(n8271), .A2(n11086), .ZN(n6972) );
  NAND2_X1 U8330 ( .A1(n8270), .A2(n6972), .ZN(n8269) );
  NAND2_X1 U8331 ( .A1(n8214), .A2(n7123), .ZN(n6974) );
  NAND2_X1 U8332 ( .A1(n7072), .A2(n10204), .ZN(n6973) );
  NAND2_X1 U8333 ( .A1(n6974), .A2(n6973), .ZN(n6975) );
  XNOR2_X1 U8334 ( .A(n6975), .B(n5119), .ZN(n6986) );
  NOR2_X1 U8335 ( .A1(n8354), .A2(n7059), .ZN(n6976) );
  AOI21_X1 U8336 ( .B1(n8214), .B2(n7072), .A(n6976), .ZN(n6984) );
  XNOR2_X1 U8337 ( .A(n6986), .B(n6984), .ZN(n8299) );
  INV_X1 U8338 ( .A(n6977), .ZN(n6979) );
  NAND2_X1 U8339 ( .A1(n6979), .A2(n6978), .ZN(n8296) );
  AND2_X1 U8340 ( .A1(n8299), .A2(n8296), .ZN(n6980) );
  NAND2_X1 U8341 ( .A1(n10612), .A2(n7123), .ZN(n6982) );
  NAND2_X1 U8342 ( .A1(n7072), .A2(n10203), .ZN(n6981) );
  NAND2_X1 U8343 ( .A1(n6982), .A2(n6981), .ZN(n6983) );
  XNOR2_X1 U8344 ( .A(n6983), .B(n7089), .ZN(n6991) );
  INV_X1 U8345 ( .A(n6984), .ZN(n6985) );
  NAND2_X1 U8346 ( .A1(n6986), .A2(n6985), .ZN(n6990) );
  AND2_X1 U8347 ( .A1(n6991), .A2(n6990), .ZN(n6987) );
  NAND2_X1 U8348 ( .A1(n10612), .A2(n7072), .ZN(n6989) );
  NAND2_X1 U8349 ( .A1(n7118), .A2(n10203), .ZN(n6988) );
  NAND2_X1 U8350 ( .A1(n6989), .A2(n6988), .ZN(n8389) );
  INV_X1 U8351 ( .A(n6991), .ZN(n6992) );
  NAND2_X1 U8352 ( .A1(n10197), .A2(n7123), .ZN(n6994) );
  NAND2_X1 U8353 ( .A1(n7072), .A2(n10202), .ZN(n6993) );
  NAND2_X1 U8354 ( .A1(n6994), .A2(n6993), .ZN(n6995) );
  XNOR2_X1 U8355 ( .A(n6995), .B(n5119), .ZN(n6998) );
  NAND2_X1 U8356 ( .A1(n6997), .A2(n6998), .ZN(n10184) );
  AND2_X1 U8357 ( .A1(n7118), .A2(n10202), .ZN(n6996) );
  NAND2_X1 U8358 ( .A1(n10184), .A2(n10186), .ZN(n7001) );
  INV_X1 U8359 ( .A(n6998), .ZN(n6999) );
  NAND2_X1 U8360 ( .A1(n10598), .A2(n7123), .ZN(n7003) );
  NAND2_X1 U8361 ( .A1(n10508), .A2(n7117), .ZN(n7002) );
  NAND2_X1 U8362 ( .A1(n7003), .A2(n7002), .ZN(n7004) );
  XNOR2_X1 U8363 ( .A(n7004), .B(n7089), .ZN(n7006) );
  AND2_X1 U8364 ( .A1(n10508), .A2(n7118), .ZN(n7005) );
  AOI21_X1 U8365 ( .B1(n10598), .B2(n7072), .A(n7005), .ZN(n7007) );
  NAND2_X1 U8366 ( .A1(n7006), .A2(n7007), .ZN(n7011) );
  INV_X1 U8367 ( .A(n7006), .ZN(n7009) );
  INV_X1 U8368 ( .A(n7007), .ZN(n7008) );
  NAND2_X1 U8369 ( .A1(n7009), .A2(n7008), .ZN(n7010) );
  AND2_X1 U8370 ( .A1(n7011), .A2(n7010), .ZN(n10098) );
  NAND2_X1 U8371 ( .A1(n10594), .A2(n7123), .ZN(n7013) );
  NAND2_X1 U8372 ( .A1(n10492), .A2(n7117), .ZN(n7012) );
  NAND2_X1 U8373 ( .A1(n7013), .A2(n7012), .ZN(n7014) );
  XNOR2_X1 U8374 ( .A(n7014), .B(n5119), .ZN(n7017) );
  NAND2_X1 U8375 ( .A1(n10594), .A2(n7117), .ZN(n7016) );
  NAND2_X1 U8376 ( .A1(n10492), .A2(n7118), .ZN(n7015) );
  NAND2_X1 U8377 ( .A1(n7016), .A2(n7015), .ZN(n7018) );
  NAND2_X1 U8378 ( .A1(n7017), .A2(n7018), .ZN(n10109) );
  INV_X1 U8379 ( .A(n7017), .ZN(n7020) );
  INV_X1 U8380 ( .A(n7018), .ZN(n7019) );
  NAND2_X1 U8381 ( .A1(n7020), .A2(n7019), .ZN(n10111) );
  NAND2_X1 U8382 ( .A1(n10107), .A2(n10111), .ZN(n7026) );
  NAND2_X1 U8383 ( .A1(n10498), .A2(n7123), .ZN(n7022) );
  NAND2_X1 U8384 ( .A1(n10510), .A2(n7117), .ZN(n7021) );
  NAND2_X1 U8385 ( .A1(n7022), .A2(n7021), .ZN(n7023) );
  XNOR2_X1 U8386 ( .A(n7023), .B(n7089), .ZN(n7027) );
  NAND2_X1 U8387 ( .A1(n7026), .A2(n7027), .ZN(n10152) );
  NAND2_X1 U8388 ( .A1(n10498), .A2(n7072), .ZN(n7025) );
  NAND2_X1 U8389 ( .A1(n10510), .A2(n7118), .ZN(n7024) );
  NAND2_X1 U8390 ( .A1(n7025), .A2(n7024), .ZN(n10155) );
  INV_X1 U8391 ( .A(n7027), .ZN(n7028) );
  NAND2_X1 U8392 ( .A1(n10479), .A2(n7123), .ZN(n7031) );
  NAND2_X1 U8393 ( .A1(n10493), .A2(n7117), .ZN(n7030) );
  NAND2_X1 U8394 ( .A1(n7031), .A2(n7030), .ZN(n7032) );
  XNOR2_X1 U8395 ( .A(n7032), .B(n7089), .ZN(n7035) );
  AND2_X1 U8396 ( .A1(n10493), .A2(n7118), .ZN(n7033) );
  AOI21_X1 U8397 ( .B1(n10479), .B2(n7072), .A(n7033), .ZN(n7034) );
  XNOR2_X1 U8398 ( .A(n7035), .B(n7034), .ZN(n10069) );
  NAND2_X1 U8399 ( .A1(n7035), .A2(n7034), .ZN(n7036) );
  NAND2_X1 U8400 ( .A1(n10066), .A2(n7036), .ZN(n10133) );
  NAND2_X1 U8401 ( .A1(n10578), .A2(n7123), .ZN(n7038) );
  NAND2_X1 U8402 ( .A1(n10474), .A2(n7117), .ZN(n7037) );
  NAND2_X1 U8403 ( .A1(n7038), .A2(n7037), .ZN(n7039) );
  XNOR2_X1 U8404 ( .A(n7039), .B(n5119), .ZN(n7041) );
  AND2_X1 U8405 ( .A1(n10474), .A2(n7118), .ZN(n7040) );
  AOI21_X1 U8406 ( .B1(n10578), .B2(n7072), .A(n7040), .ZN(n7042) );
  XNOR2_X1 U8407 ( .A(n7041), .B(n7042), .ZN(n10134) );
  NAND2_X1 U8408 ( .A1(n10133), .A2(n10134), .ZN(n10132) );
  INV_X1 U8409 ( .A(n7041), .ZN(n7043) );
  NAND2_X1 U8410 ( .A1(n7043), .A2(n7042), .ZN(n7044) );
  NAND2_X1 U8411 ( .A1(n10132), .A2(n7044), .ZN(n10076) );
  INV_X1 U8412 ( .A(n10076), .ZN(n7050) );
  NAND2_X1 U8413 ( .A1(n10572), .A2(n7123), .ZN(n7046) );
  NAND2_X1 U8414 ( .A1(n10464), .A2(n7072), .ZN(n7045) );
  NAND2_X1 U8415 ( .A1(n7046), .A2(n7045), .ZN(n7047) );
  XNOR2_X1 U8416 ( .A(n7047), .B(n7089), .ZN(n7051) );
  AND2_X1 U8417 ( .A1(n10464), .A2(n7118), .ZN(n7048) );
  AOI21_X1 U8418 ( .B1(n10572), .B2(n7072), .A(n7048), .ZN(n7052) );
  XNOR2_X1 U8419 ( .A(n7051), .B(n7052), .ZN(n10077) );
  INV_X1 U8420 ( .A(n10077), .ZN(n7049) );
  NAND2_X1 U8421 ( .A1(n7050), .A2(n7049), .ZN(n10078) );
  INV_X1 U8422 ( .A(n7051), .ZN(n7054) );
  INV_X1 U8423 ( .A(n7052), .ZN(n7053) );
  NAND2_X1 U8424 ( .A1(n7054), .A2(n7053), .ZN(n7055) );
  NAND2_X1 U8425 ( .A1(n10568), .A2(n7123), .ZN(n7057) );
  NAND2_X1 U8426 ( .A1(n10441), .A2(n7072), .ZN(n7056) );
  NAND2_X1 U8427 ( .A1(n7057), .A2(n7056), .ZN(n7058) );
  XNOR2_X1 U8428 ( .A(n7058), .B(n7089), .ZN(n7061) );
  INV_X1 U8429 ( .A(n10568), .ZN(n10427) );
  OAI22_X1 U8430 ( .A1(n10427), .A2(n7060), .B1(n10082), .B2(n7059), .ZN(
        n10143) );
  XNOR2_X1 U8431 ( .A(n7063), .B(n7062), .ZN(n10059) );
  NAND2_X1 U8432 ( .A1(n10558), .A2(n7123), .ZN(n7066) );
  NAND2_X1 U8433 ( .A1(n10416), .A2(n7072), .ZN(n7065) );
  NAND2_X1 U8434 ( .A1(n7066), .A2(n7065), .ZN(n7067) );
  XNOR2_X1 U8435 ( .A(n7067), .B(n5119), .ZN(n7071) );
  NAND2_X1 U8436 ( .A1(n10558), .A2(n7072), .ZN(n7069) );
  NAND2_X1 U8437 ( .A1(n10416), .A2(n7118), .ZN(n7068) );
  NAND2_X1 U8438 ( .A1(n7069), .A2(n7068), .ZN(n7070) );
  NAND2_X1 U8439 ( .A1(n7071), .A2(n7070), .ZN(n10121) );
  NOR2_X1 U8440 ( .A1(n7071), .A2(n7070), .ZN(n10120) );
  AOI21_X2 U8441 ( .B1(n10124), .B2(n10121), .A(n10120), .ZN(n10088) );
  AOI22_X1 U8442 ( .A1(n10373), .A2(n7072), .B1(n7118), .B2(n10391), .ZN(n7076) );
  NAND2_X1 U8443 ( .A1(n10373), .A2(n7123), .ZN(n7074) );
  NAND2_X1 U8444 ( .A1(n10391), .A2(n7072), .ZN(n7073) );
  NAND2_X1 U8445 ( .A1(n7074), .A2(n7073), .ZN(n7075) );
  XNOR2_X1 U8446 ( .A(n7075), .B(n5119), .ZN(n7078) );
  XOR2_X1 U8447 ( .A(n7076), .B(n7078), .Z(n10087) );
  INV_X1 U8448 ( .A(n7076), .ZN(n7077) );
  NOR2_X1 U8449 ( .A1(n7078), .A2(n7077), .ZN(n10175) );
  NAND2_X1 U8450 ( .A1(n10353), .A2(n7123), .ZN(n7080) );
  NAND2_X1 U8451 ( .A1(n10381), .A2(n7117), .ZN(n7079) );
  NAND2_X1 U8452 ( .A1(n7080), .A2(n7079), .ZN(n7081) );
  XNOR2_X1 U8453 ( .A(n7081), .B(n7089), .ZN(n7083) );
  AND2_X1 U8454 ( .A1(n10381), .A2(n7118), .ZN(n7082) );
  AOI21_X1 U8455 ( .B1(n10353), .B2(n7072), .A(n7082), .ZN(n7084) );
  XNOR2_X1 U8456 ( .A(n7083), .B(n7084), .ZN(n10174) );
  INV_X1 U8457 ( .A(n7083), .ZN(n7086) );
  INV_X1 U8458 ( .A(n7084), .ZN(n7085) );
  NAND2_X1 U8459 ( .A1(n10344), .A2(n7123), .ZN(n7088) );
  NAND2_X1 U8460 ( .A1(n10363), .A2(n7072), .ZN(n7087) );
  NAND2_X1 U8461 ( .A1(n7088), .A2(n7087), .ZN(n7090) );
  XNOR2_X1 U8462 ( .A(n7090), .B(n7089), .ZN(n7093) );
  AND2_X1 U8463 ( .A1(n10363), .A2(n7118), .ZN(n7091) );
  AOI21_X1 U8464 ( .B1(n10344), .B2(n7072), .A(n7091), .ZN(n7092) );
  NAND2_X1 U8465 ( .A1(n7093), .A2(n7092), .ZN(n7131) );
  OAI21_X1 U8466 ( .B1(n7093), .B2(n7092), .A(n7131), .ZN(n7094) );
  OAI21_X1 U8467 ( .B1(n10173), .B2(n7095), .A(n7094), .ZN(n7096) );
  INV_X1 U8468 ( .A(n7096), .ZN(n7099) );
  NAND3_X1 U8469 ( .A1(n7098), .A2(n7565), .A3(n7097), .ZN(n7106) );
  NOR2_X1 U8470 ( .A1(n7106), .A2(n8851), .ZN(n7100) );
  AND2_X1 U8471 ( .A1(n11109), .A2(n7193), .ZN(n7101) );
  INV_X1 U8472 ( .A(n7100), .ZN(n7113) );
  OR2_X1 U8473 ( .A1(n7113), .A2(n7571), .ZN(n7108) );
  NOR2_X2 U8474 ( .A1(n7108), .A2(n7248), .ZN(n11091) );
  NAND2_X1 U8475 ( .A1(n7106), .A2(n7101), .ZN(n7104) );
  AND3_X1 U8476 ( .A1(n6847), .A2(n7195), .A3(n7102), .ZN(n7103) );
  NAND2_X1 U8477 ( .A1(n7104), .A2(n7103), .ZN(n7288) );
  NAND2_X1 U8478 ( .A1(n7288), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7107) );
  NAND2_X1 U8479 ( .A1(n8856), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7983) );
  OAI21_X1 U8480 ( .B1(n8851), .B2(n7571), .A(n7983), .ZN(n7105) );
  NAND2_X1 U8481 ( .A1(n7106), .A2(n7105), .ZN(n7289) );
  INV_X1 U8482 ( .A(n10345), .ZN(n7110) );
  AOI22_X1 U8483 ( .A1(n10381), .A2(n10189), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n7109) );
  OAI21_X1 U8484 ( .B1(n11101), .B2(n7110), .A(n7109), .ZN(n7111) );
  AOI21_X1 U8485 ( .B1(n11091), .B2(n10338), .A(n7111), .ZN(n7116) );
  OR2_X1 U8486 ( .A1(n7112), .A2(n8921), .ZN(n7569) );
  OR2_X1 U8487 ( .A1(n7113), .A2(n7569), .ZN(n7115) );
  NAND2_X1 U8488 ( .A1(n10325), .A2(n7117), .ZN(n7120) );
  NAND2_X1 U8489 ( .A1(n10338), .A2(n7118), .ZN(n7119) );
  NAND2_X1 U8490 ( .A1(n7120), .A2(n7119), .ZN(n7122) );
  XNOR2_X1 U8491 ( .A(n7122), .B(n5119), .ZN(n7125) );
  AOI22_X1 U8492 ( .A1(n10325), .A2(n7123), .B1(n7072), .B2(n10338), .ZN(n7124) );
  XNOR2_X1 U8493 ( .A(n7125), .B(n7124), .ZN(n7127) );
  INV_X1 U8494 ( .A(n7127), .ZN(n7132) );
  NAND3_X1 U8495 ( .A1(n7132), .A2(n11097), .A3(n7131), .ZN(n7126) );
  OR2_X2 U8496 ( .A1(n7128), .A2(n7126), .ZN(n7137) );
  AOI22_X1 U8497 ( .A1(n7886), .A2(n11091), .B1(n10189), .B2(n10363), .ZN(
        n7130) );
  NAND2_X1 U8498 ( .A1(P1_U3086), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7129) );
  OAI211_X1 U8499 ( .C1(n11101), .C2(n10324), .A(n7130), .B(n7129), .ZN(n7134)
         );
  NOR3_X1 U8500 ( .A1(n7132), .A2(n10199), .A3(n7131), .ZN(n7133) );
  AOI211_X1 U8501 ( .C1(n10325), .C2(n11088), .A(n7134), .B(n7133), .ZN(n7135)
         );
  NAND3_X1 U8502 ( .A1(n7137), .A2(n7136), .A3(n7135), .ZN(P1_U3220) );
  OAI21_X1 U8503 ( .B1(n7361), .B2(n7353), .A(n9312), .ZN(n7142) );
  INV_X1 U8504 ( .A(n7145), .ZN(n7140) );
  NAND2_X1 U8505 ( .A1(n7142), .A2(n7362), .ZN(n7148) );
  AND2_X1 U8506 ( .A1(n9244), .A2(n11127), .ZN(n7357) );
  NAND2_X1 U8507 ( .A1(n7357), .A2(n7353), .ZN(n7144) );
  NAND2_X1 U8508 ( .A1(n7144), .A2(n10974), .ZN(n7351) );
  NAND3_X1 U8509 ( .A1(n7339), .A2(n7761), .A3(n7145), .ZN(n7368) );
  NOR2_X1 U8510 ( .A1(n7368), .A2(n7361), .ZN(n7146) );
  NAND2_X1 U8511 ( .A1(n7351), .A2(n7146), .ZN(n7147) );
  OR2_X1 U8512 ( .A1(n11157), .A2(n6747), .ZN(n7149) );
  NAND2_X1 U8513 ( .A1(n7150), .A2(n7149), .ZN(P2_U3456) );
  INV_X1 U8514 ( .A(n7190), .ZN(n7186) );
  OR2_X2 U8515 ( .A1(n6847), .A2(n7186), .ZN(n10215) );
  INV_X1 U8516 ( .A(n7259), .ZN(n7151) );
  NAND2_X1 U8517 ( .A1(n9244), .A2(n7365), .ZN(n7152) );
  NAND2_X1 U8518 ( .A1(n7152), .A2(n8266), .ZN(n7317) );
  NAND2_X1 U8519 ( .A1(n7317), .A2(n7153), .ZN(n7154) );
  NAND2_X1 U8520 ( .A1(n7154), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X2 U8521 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  AND2_X1 U8522 ( .A1(n7159), .A2(P1_U3086), .ZN(n10663) );
  INV_X2 U8523 ( .A(n10663), .ZN(n7742) );
  INV_X1 U8524 ( .A(n10659), .ZN(n7296) );
  AOI22_X1 U8525 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n7296), .B1(n10250), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n7156) );
  OAI21_X1 U8526 ( .B1(n7161), .B2(n7742), .A(n7156), .ZN(P1_U3352) );
  OAI222_X1 U8527 ( .A1(n10659), .A2(n5628), .B1(n7742), .B2(n7168), .C1(
        P1_U3086), .C2(n7231), .ZN(P1_U3354) );
  AOI22_X1 U8528 ( .A1(n10276), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n7296), .ZN(n7157) );
  OAI21_X1 U8529 ( .B1(n7163), .B2(n7742), .A(n7157), .ZN(P1_U3350) );
  AOI22_X1 U8530 ( .A1(n10289), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n7296), .ZN(n7158) );
  OAI21_X1 U8531 ( .B1(n7166), .B2(n7742), .A(n7158), .ZN(P1_U3349) );
  INV_X1 U8532 ( .A(n8985), .ZN(n8534) );
  NOR2_X1 U8533 ( .A1(n7159), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10054) );
  INV_X2 U8534 ( .A(n10054), .ZN(n8998) );
  OAI222_X1 U8535 ( .A1(n8985), .A2(n7160), .B1(n8998), .B2(n7169), .C1(
        P2_U3151), .C2(n10886), .ZN(P2_U3293) );
  OAI222_X1 U8536 ( .A1(n8985), .A2(n7162), .B1(n8998), .B2(n7161), .C1(
        P2_U3151), .C2(n7546), .ZN(P2_U3292) );
  OAI222_X1 U8537 ( .A1(n8985), .A2(n7164), .B1(n8998), .B2(n7163), .C1(
        P2_U3151), .C2(n7683), .ZN(P2_U3290) );
  OAI222_X1 U8538 ( .A1(n8985), .A2(n7165), .B1(n8998), .B2(n7171), .C1(
        P2_U3151), .C2(n7520), .ZN(P2_U3291) );
  OAI222_X1 U8539 ( .A1(n8985), .A2(n7167), .B1(n8998), .B2(n7166), .C1(
        P2_U3151), .C2(n10903), .ZN(P2_U3289) );
  OAI222_X1 U8540 ( .A1(P2_U3151), .A2(n7416), .B1(n8998), .B2(n7168), .C1(
        n5631), .C2(n8985), .ZN(P2_U3294) );
  OAI222_X1 U8541 ( .A1(n10659), .A2(n7170), .B1(n7742), .B2(n7169), .C1(
        P1_U3086), .C2(n7230), .ZN(P1_U3353) );
  INV_X1 U8542 ( .A(n7236), .ZN(n10260) );
  OAI222_X1 U8543 ( .A1(n10659), .A2(n5324), .B1(n7742), .B2(n7171), .C1(
        P1_U3086), .C2(n10260), .ZN(P1_U3351) );
  INV_X1 U8544 ( .A(n7172), .ZN(n7174) );
  AOI22_X1 U8545 ( .A1(n10302), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7296), .ZN(n7173) );
  OAI21_X1 U8546 ( .B1(n7174), .B2(n7742), .A(n7173), .ZN(P1_U3348) );
  INV_X1 U8547 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7175) );
  OAI222_X1 U8548 ( .A1(n8985), .A2(n7175), .B1(n8998), .B2(n7174), .C1(
        P2_U3151), .C2(n7990), .ZN(P2_U3288) );
  INV_X1 U8549 ( .A(n7176), .ZN(n7178) );
  OAI222_X1 U8550 ( .A1(n8985), .A2(n7177), .B1(n8998), .B2(n7178), .C1(
        P2_U3151), .C2(n8103), .ZN(P2_U3287) );
  INV_X1 U8551 ( .A(n7242), .ZN(n10768) );
  OAI222_X1 U8552 ( .A1(n10659), .A2(n9810), .B1(n7742), .B2(n7178), .C1(
        P1_U3086), .C2(n10768), .ZN(P1_U3347) );
  INV_X1 U8553 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7181) );
  INV_X1 U8554 ( .A(n7761), .ZN(n7179) );
  NAND2_X1 U8555 ( .A1(n7179), .A2(n7192), .ZN(n7180) );
  OAI21_X1 U8556 ( .B1(n7192), .B2(n7181), .A(n7180), .ZN(P2_U3377) );
  INV_X1 U8557 ( .A(n7182), .ZN(n7184) );
  INV_X1 U8558 ( .A(n8851), .ZN(n7183) );
  INV_X1 U8559 ( .A(n8452), .ZN(n7185) );
  NOR3_X1 U8560 ( .A1(n6326), .A2(n7186), .A3(n7185), .ZN(n7187) );
  AOI21_X1 U8561 ( .B1(n10671), .B2(n7188), .A(n7187), .ZN(P1_U3440) );
  AOI22_X1 U8562 ( .A1(n10671), .A2(n7191), .B1(n7190), .B2(n7189), .ZN(
        P1_U3439) );
  AND2_X1 U8563 ( .A1(n7256), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8564 ( .A1(n7256), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8565 ( .A1(n7256), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8566 ( .A1(n7256), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8567 ( .A1(n7256), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8568 ( .A1(n7256), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8569 ( .A1(n7256), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8570 ( .A1(n7256), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8571 ( .A1(n7256), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8572 ( .A1(n7256), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8573 ( .A1(n7256), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  OR2_X1 U8574 ( .A1(n7195), .A2(P1_U3086), .ZN(n8861) );
  NAND2_X1 U8575 ( .A1(n8851), .A2(n8861), .ZN(n7229) );
  INV_X1 U8576 ( .A(n7193), .ZN(n8843) );
  AOI21_X1 U8577 ( .B1(n8843), .B2(n7195), .A(n7194), .ZN(n7228) );
  INV_X1 U8578 ( .A(n7228), .ZN(n7196) );
  AND2_X1 U8579 ( .A1(n7229), .A2(n7196), .ZN(n10754) );
  NOR2_X1 U8580 ( .A1(n10754), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8581 ( .A(n7197), .ZN(n7199) );
  OAI222_X1 U8582 ( .A1(n8985), .A2(n7198), .B1(n8998), .B2(n7199), .C1(n8102), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8583 ( .A(n7271), .ZN(n7249) );
  OAI222_X1 U8584 ( .A1(n10659), .A2(n9591), .B1(n7742), .B2(n7199), .C1(n7249), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8585 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7201) );
  INV_X1 U8586 ( .A(n7200), .ZN(n7202) );
  INV_X1 U8587 ( .A(n10857), .ZN(n7263) );
  OAI222_X1 U8588 ( .A1(n10659), .A2(n7201), .B1(n7742), .B2(n7202), .C1(n7263), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8589 ( .A(n8428), .ZN(n8434) );
  INV_X1 U8590 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7206) );
  OAI222_X1 U8591 ( .A1(P2_U3151), .A2(n8434), .B1(n8985), .B2(n7206), .C1(
        n7202), .C2(n8998), .ZN(P2_U3285) );
  MUX2_X1 U8592 ( .A(n9591), .B(n7203), .S(P2_U3893), .Z(n7204) );
  INV_X1 U8593 ( .A(n7204), .ZN(P2_U3500) );
  NAND2_X1 U8594 ( .A1(P1_U3973), .A2(n7916), .ZN(n7205) );
  OAI21_X1 U8595 ( .B1(P1_U3973), .B2(n7206), .A(n7205), .ZN(P1_U3564) );
  INV_X1 U8596 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7211) );
  INV_X1 U8597 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n7209) );
  NAND2_X1 U8598 ( .A1(n8647), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7208) );
  INV_X1 U8599 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10532) );
  OR2_X1 U8600 ( .A1(n8649), .A2(n10532), .ZN(n7207) );
  OAI211_X1 U8601 ( .C1(n8653), .C2(n7209), .A(n7208), .B(n7207), .ZN(n10313)
         );
  NAND2_X1 U8602 ( .A1(P1_U3973), .A2(n10313), .ZN(n7210) );
  OAI21_X1 U8603 ( .B1(P1_U3973), .B2(n7211), .A(n7210), .ZN(P1_U3585) );
  INV_X1 U8604 ( .A(n7212), .ZN(n7254) );
  AOI22_X1 U8605 ( .A1(n10773), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n7296), .ZN(n7213) );
  OAI21_X1 U8606 ( .B1(n7254), .B2(n7742), .A(n7213), .ZN(P1_U3344) );
  AOI22_X1 U8607 ( .A1(n7271), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n5902), .B2(
        n7249), .ZN(n7226) );
  XNOR2_X1 U8608 ( .A(n7230), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n10240) );
  XNOR2_X1 U8609 ( .A(n7231), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U8610 ( .A1(n10752), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10229) );
  INV_X1 U8611 ( .A(n10229), .ZN(n10217) );
  NAND2_X1 U8612 ( .A1(n10218), .A2(n10217), .ZN(n10216) );
  INV_X1 U8613 ( .A(n7231), .ZN(n10222) );
  NAND2_X1 U8614 ( .A1(n10222), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U8615 ( .A1(n10216), .A2(n7214), .ZN(n10239) );
  NAND2_X1 U8616 ( .A1(n10240), .A2(n10239), .ZN(n10238) );
  INV_X1 U8617 ( .A(n7230), .ZN(n10237) );
  NAND2_X1 U8618 ( .A1(n10237), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7215) );
  NAND2_X1 U8619 ( .A1(n10238), .A2(n7215), .ZN(n10252) );
  XNOR2_X1 U8620 ( .A(n10250), .B(n7216), .ZN(n10253) );
  NAND2_X1 U8621 ( .A1(n10252), .A2(n10253), .ZN(n10251) );
  NAND2_X1 U8622 ( .A1(n10250), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7217) );
  NAND2_X1 U8623 ( .A1(n10251), .A2(n7217), .ZN(n10267) );
  MUX2_X1 U8624 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7597), .S(n7236), .Z(n10268)
         );
  NAND2_X1 U8625 ( .A1(n10267), .A2(n10268), .ZN(n10266) );
  NAND2_X1 U8626 ( .A1(n7236), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7218) );
  NAND2_X1 U8627 ( .A1(n10266), .A2(n7218), .ZN(n10278) );
  XNOR2_X1 U8628 ( .A(n10276), .B(n11014), .ZN(n10279) );
  NAND2_X1 U8629 ( .A1(n10278), .A2(n10279), .ZN(n10277) );
  NAND2_X1 U8630 ( .A1(n10276), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7219) );
  NAND2_X1 U8631 ( .A1(n10277), .A2(n7219), .ZN(n10291) );
  MUX2_X1 U8632 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n5847), .S(n10289), .Z(n10292) );
  NAND2_X1 U8633 ( .A1(n10291), .A2(n10292), .ZN(n10290) );
  NAND2_X1 U8634 ( .A1(n10289), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7220) );
  NAND2_X1 U8635 ( .A1(n10290), .A2(n7220), .ZN(n10304) );
  XNOR2_X1 U8636 ( .A(n10302), .B(n7221), .ZN(n10305) );
  NAND2_X1 U8637 ( .A1(n10304), .A2(n10305), .ZN(n10303) );
  NAND2_X1 U8638 ( .A1(n10302), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7222) );
  NAND2_X1 U8639 ( .A1(n10303), .A2(n7222), .ZN(n10760) );
  OR2_X1 U8640 ( .A1(n7242), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7224) );
  NAND2_X1 U8641 ( .A1(n7242), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7223) );
  AND2_X1 U8642 ( .A1(n7224), .A2(n7223), .ZN(n10761) );
  AND2_X1 U8643 ( .A1(n10760), .A2(n10761), .ZN(n10758) );
  AOI21_X1 U8644 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7242), .A(n10758), .ZN(
        n7225) );
  NAND2_X1 U8645 ( .A1(n7226), .A2(n7225), .ZN(n7262) );
  OAI21_X1 U8646 ( .B1(n7226), .B2(n7225), .A(n7262), .ZN(n7227) );
  INV_X1 U8647 ( .A(n7227), .ZN(n7253) );
  NAND2_X1 U8648 ( .A1(n7229), .A2(n7228), .ZN(n10756) );
  OR2_X1 U8649 ( .A1(n5123), .A2(n10748), .ZN(n8848) );
  OR2_X1 U8650 ( .A1(n10756), .A2(n8848), .ZN(n10851) );
  AOI22_X1 U8651 ( .A1(n7271), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n5906), .B2(
        n7249), .ZN(n7244) );
  XNOR2_X1 U8652 ( .A(n7230), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n10243) );
  XNOR2_X1 U8653 ( .A(n7231), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n10221) );
  AND2_X1 U8654 ( .A1(n10752), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10220) );
  NAND2_X1 U8655 ( .A1(n10221), .A2(n10220), .ZN(n10219) );
  NAND2_X1 U8656 ( .A1(n10222), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7232) );
  NAND2_X1 U8657 ( .A1(n10219), .A2(n7232), .ZN(n10242) );
  NAND2_X1 U8658 ( .A1(n10243), .A2(n10242), .ZN(n10241) );
  NAND2_X1 U8659 ( .A1(n10237), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7233) );
  NAND2_X1 U8660 ( .A1(n10241), .A2(n7233), .ZN(n10255) );
  XNOR2_X1 U8661 ( .A(n10250), .B(n7234), .ZN(n10256) );
  NAND2_X1 U8662 ( .A1(n10255), .A2(n10256), .ZN(n10254) );
  NAND2_X1 U8663 ( .A1(n10250), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7235) );
  NAND2_X1 U8664 ( .A1(n10254), .A2(n7235), .ZN(n10264) );
  INV_X1 U8665 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n11002) );
  MUX2_X1 U8666 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n11002), .S(n7236), .Z(n10265) );
  NAND2_X1 U8667 ( .A1(n10264), .A2(n10265), .ZN(n10263) );
  NAND2_X1 U8668 ( .A1(n7236), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7237) );
  NAND2_X1 U8669 ( .A1(n10263), .A2(n7237), .ZN(n10281) );
  INV_X1 U8670 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7238) );
  XNOR2_X1 U8671 ( .A(n10276), .B(n7238), .ZN(n10282) );
  NAND2_X1 U8672 ( .A1(n10281), .A2(n10282), .ZN(n10280) );
  NAND2_X1 U8673 ( .A1(n10276), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7239) );
  NAND2_X1 U8674 ( .A1(n10280), .A2(n7239), .ZN(n10294) );
  INV_X1 U8675 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11033) );
  MUX2_X1 U8676 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n11033), .S(n10289), .Z(
        n10295) );
  NAND2_X1 U8677 ( .A1(n10294), .A2(n10295), .ZN(n10293) );
  NAND2_X1 U8678 ( .A1(n10289), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7240) );
  NAND2_X1 U8679 ( .A1(n10293), .A2(n7240), .ZN(n10307) );
  MUX2_X1 U8680 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n5863), .S(n10302), .Z(n10308) );
  NAND2_X1 U8681 ( .A1(n10307), .A2(n10308), .ZN(n10306) );
  NAND2_X1 U8682 ( .A1(n10302), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7241) );
  NAND2_X1 U8683 ( .A1(n10306), .A2(n7241), .ZN(n10764) );
  MUX2_X1 U8684 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n5883), .S(n7242), .Z(n10765)
         );
  AND2_X1 U8685 ( .A1(n10764), .A2(n10765), .ZN(n10762) );
  AOI21_X1 U8686 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7242), .A(n10762), .ZN(
        n7243) );
  NAND2_X1 U8687 ( .A1(n7244), .A2(n7243), .ZN(n7270) );
  OAI21_X1 U8688 ( .B1(n7244), .B2(n7243), .A(n7270), .ZN(n7246) );
  INV_X1 U8689 ( .A(n10748), .ZN(n7245) );
  OR2_X1 U8690 ( .A1(n10756), .A2(n7245), .ZN(n10847) );
  NAND2_X1 U8691 ( .A1(n7246), .A2(n10822), .ZN(n7252) );
  NOR2_X1 U8692 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7247), .ZN(n7942) );
  NOR2_X1 U8693 ( .A1(n10829), .A2(n7249), .ZN(n7250) );
  AOI211_X1 U8694 ( .C1(n10754), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7942), .B(
        n7250), .ZN(n7251) );
  OAI211_X1 U8695 ( .C1(n7253), .C2(n10851), .A(n7252), .B(n7251), .ZN(
        P1_U3252) );
  OAI222_X1 U8696 ( .A1(n8985), .A2(n7255), .B1(n8998), .B2(n7254), .C1(
        P2_U3151), .C2(n8438), .ZN(P2_U3284) );
  INV_X1 U8697 ( .A(n7257), .ZN(n7258) );
  AOI22_X1 U8698 ( .A1(n7256), .A2(n5703), .B1(n7259), .B2(n7258), .ZN(
        P2_U3376) );
  AND2_X1 U8699 ( .A1(n7256), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8700 ( .A1(n7256), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8701 ( .A1(n7256), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8702 ( .A1(n7256), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8703 ( .A1(n7256), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8704 ( .A1(n7256), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8705 ( .A1(n7256), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8706 ( .A1(n7256), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8707 ( .A1(n7256), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8708 ( .A1(n7256), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8709 ( .A1(n7256), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8710 ( .A1(n7256), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8711 ( .A1(n7256), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8712 ( .A1(n7256), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8713 ( .A1(n7256), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8714 ( .A1(n7256), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8715 ( .A1(n7256), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8716 ( .A1(n7256), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8717 ( .A1(n7256), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  INV_X1 U8718 ( .A(n7260), .ZN(n7280) );
  AOI22_X1 U8719 ( .A1(n8501), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8534), .ZN(n7261) );
  OAI21_X1 U8720 ( .B1(n7280), .B2(n8998), .A(n7261), .ZN(P2_U3283) );
  INV_X1 U8721 ( .A(n8026), .ZN(n7279) );
  AOI22_X1 U8722 ( .A1(n8026), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n5955), .B2(
        n7279), .ZN(n7266) );
  OAI21_X1 U8723 ( .B1(n7271), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7262), .ZN(
        n10854) );
  AOI22_X1 U8724 ( .A1(n10857), .A2(n7830), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n7263), .ZN(n10853) );
  NOR2_X1 U8725 ( .A1(n10854), .A2(n10853), .ZN(n10852) );
  AOI21_X1 U8726 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n10857), .A(n10852), .ZN(
        n10775) );
  NAND2_X1 U8727 ( .A1(n10773), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7264) );
  OAI21_X1 U8728 ( .B1(n10773), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7264), .ZN(
        n10776) );
  NOR2_X1 U8729 ( .A1(n10775), .A2(n10776), .ZN(n10774) );
  AOI21_X1 U8730 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10773), .A(n10774), .ZN(
        n7265) );
  NAND2_X1 U8731 ( .A1(n7266), .A2(n7265), .ZN(n8025) );
  OAI21_X1 U8732 ( .B1(n7266), .B2(n7265), .A(n8025), .ZN(n7267) );
  INV_X1 U8733 ( .A(n7267), .ZN(n7278) );
  AND2_X1 U8734 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8276) );
  NOR2_X1 U8735 ( .A1(n10829), .A2(n7279), .ZN(n7268) );
  AOI211_X1 U8736 ( .C1(n10754), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n8276), .B(
        n7268), .ZN(n7277) );
  AOI22_X1 U8737 ( .A1(n8026), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5959), .B2(
        n7279), .ZN(n7274) );
  INV_X1 U8738 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7269) );
  MUX2_X1 U8739 ( .A(n7269), .B(P1_REG1_REG_10__SCAN_IN), .S(n10857), .Z(
        n10849) );
  OAI21_X1 U8740 ( .B1(n7271), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7270), .ZN(
        n10850) );
  NOR2_X1 U8741 ( .A1(n10849), .A2(n10850), .ZN(n10848) );
  AOI21_X1 U8742 ( .B1(n10857), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10848), .ZN(
        n10779) );
  MUX2_X1 U8743 ( .A(n7272), .B(P1_REG1_REG_11__SCAN_IN), .S(n10773), .Z(
        n10780) );
  NOR2_X1 U8744 ( .A1(n10779), .A2(n10780), .ZN(n10778) );
  AOI21_X1 U8745 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n10773), .A(n10778), .ZN(
        n7273) );
  NAND2_X1 U8746 ( .A1(n7274), .A2(n7273), .ZN(n8016) );
  OAI21_X1 U8747 ( .B1(n7274), .B2(n7273), .A(n8016), .ZN(n7275) );
  NAND2_X1 U8748 ( .A1(n7275), .A2(n10822), .ZN(n7276) );
  OAI211_X1 U8749 ( .C1(n7278), .C2(n10851), .A(n7277), .B(n7276), .ZN(
        P1_U3255) );
  INV_X1 U8750 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7281) );
  OAI222_X1 U8751 ( .A1(n10659), .A2(n7281), .B1(n7742), .B2(n7280), .C1(n7279), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8752 ( .A(n7282), .ZN(n7293) );
  AOI22_X1 U8753 ( .A1(n10842), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7296), .ZN(n7283) );
  OAI21_X1 U8754 ( .B1(n7293), .B2(n7742), .A(n7283), .ZN(P1_U3342) );
  OR2_X1 U8755 ( .A1(n7285), .A2(n7284), .ZN(n7286) );
  NAND2_X1 U8756 ( .A1(n7287), .A2(n7286), .ZN(n10227) );
  AOI22_X1 U8757 ( .A1(n10932), .A2(n11088), .B1(n11091), .B2(n10214), .ZN(
        n7292) );
  INV_X1 U8758 ( .A(n7288), .ZN(n7290) );
  NAND3_X1 U8759 ( .A1(n7290), .A2(P1_STATE_REG_SCAN_IN), .A3(n7289), .ZN(
        n7441) );
  NAND2_X1 U8760 ( .A1(n7441), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7291) );
  OAI211_X1 U8761 ( .C1(n10227), .C2(n10199), .A(n7292), .B(n7291), .ZN(
        P1_U3232) );
  INV_X1 U8762 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7294) );
  OAI222_X1 U8763 ( .A1(n8985), .A2(n7294), .B1(n8998), .B2(n7293), .C1(
        P2_U3151), .C2(n8498), .ZN(P2_U3282) );
  INV_X1 U8764 ( .A(n7295), .ZN(n7310) );
  AOI22_X1 U8765 ( .A1(n10789), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7296), .ZN(n7297) );
  OAI21_X1 U8766 ( .B1(n7310), .B2(n7742), .A(n7297), .ZN(P1_U3341) );
  OAI21_X1 U8767 ( .B1(n7299), .B2(n8786), .A(n7298), .ZN(n7708) );
  INV_X1 U8768 ( .A(n10212), .ZN(n7300) );
  NOR2_X1 U8769 ( .A1(n7300), .A2(n8944), .ZN(n7703) );
  INV_X1 U8770 ( .A(n7703), .ZN(n7302) );
  XNOR2_X1 U8771 ( .A(n7448), .B(n7704), .ZN(n7301) );
  NAND2_X1 U8772 ( .A1(n7301), .A2(n10599), .ZN(n7706) );
  NAND2_X1 U8773 ( .A1(n7302), .A2(n7706), .ZN(n7306) );
  XNOR2_X1 U8774 ( .A(n7303), .B(n8786), .ZN(n7305) );
  OAI22_X1 U8775 ( .A1(n7305), .A2(n10929), .B1(n7304), .B2(n8353), .ZN(n7702)
         );
  AOI211_X1 U8776 ( .C1(n11113), .C2(n7708), .A(n7306), .B(n7702), .ZN(n7338)
         );
  INV_X1 U8777 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7307) );
  OAI22_X1 U8778 ( .A1(n10651), .A2(n7335), .B1(n11120), .B2(n7307), .ZN(n7308) );
  INV_X1 U8779 ( .A(n7308), .ZN(n7309) );
  OAI21_X1 U8780 ( .B1(n7338), .B2(n11117), .A(n7309), .ZN(P1_U3459) );
  OAI222_X1 U8781 ( .A1(n8985), .A2(n7311), .B1(n8998), .B2(n7310), .C1(
        P2_U3151), .C2(n9347), .ZN(P2_U3281) );
  NOR2_X1 U8782 ( .A1(n9412), .A2(P2_U3151), .ZN(n8483) );
  AND2_X1 U8783 ( .A1(n7317), .A2(n8483), .ZN(n7312) );
  MUX2_X1 U8784 ( .A(P2_U3893), .B(n7312), .S(n6788), .Z(n10906) );
  INV_X1 U8785 ( .A(n8266), .ZN(n7313) );
  NOR2_X1 U8786 ( .A1(n7365), .A2(n7313), .ZN(n7314) );
  AND2_X1 U8787 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n7319), .ZN(n7315) );
  NOR2_X1 U8788 ( .A1(n7316), .A2(n7324), .ZN(n7405) );
  AOI21_X1 U8789 ( .B1(n7324), .B2(n7316), .A(n7405), .ZN(n7331) );
  NOR2_X1 U8790 ( .A1(n6788), .A2(P2_U3151), .ZN(n8533) );
  INV_X1 U8791 ( .A(n10865), .ZN(n7318) );
  AOI21_X1 U8792 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n7319), .A(n7416), .ZN(
        n7322) );
  NOR2_X1 U8793 ( .A1(n7321), .A2(n7320), .ZN(n7392) );
  NOR2_X1 U8794 ( .A1(n7322), .A2(n7392), .ZN(n7393) );
  XOR2_X1 U8795 ( .A(n7323), .B(n7393), .Z(n7329) );
  MUX2_X1 U8796 ( .A(n7324), .B(n7323), .S(n6789), .Z(n7418) );
  XNOR2_X1 U8797 ( .A(n7418), .B(n7416), .ZN(n7326) );
  MUX2_X1 U8798 ( .A(n10947), .B(n7320), .S(n9412), .Z(n10863) );
  NAND2_X1 U8799 ( .A1(n10863), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7325) );
  NAND2_X1 U8800 ( .A1(n7326), .A2(n7325), .ZN(n7417) );
  NAND2_X1 U8801 ( .A1(P2_U3893), .A2(n6788), .ZN(n9426) );
  OAI211_X1 U8802 ( .C1(n7326), .C2(n7325), .A(n7417), .B(n10923), .ZN(n7327)
         );
  OAI21_X1 U8803 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n8072), .A(n7327), .ZN(n7328) );
  AOI21_X1 U8804 ( .B1(n9429), .B2(n7329), .A(n7328), .ZN(n7330) );
  OAI21_X1 U8805 ( .B1(n7331), .B2(n10918), .A(n7330), .ZN(n7332) );
  AOI21_X1 U8806 ( .B1(n10907), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n7332), .ZN(
        n7333) );
  OAI21_X1 U8807 ( .B1(n7416), .B2(n10904), .A(n7333), .ZN(P2_U3183) );
  NAND2_X1 U8808 ( .A1(n10433), .A2(P1_U3973), .ZN(n7334) );
  OAI21_X1 U8809 ( .B1(P1_U3973), .B2(n8268), .A(n7334), .ZN(P1_U3577) );
  OAI22_X1 U8810 ( .A1(n10592), .A2(n7335), .B1(n11116), .B2(n5763), .ZN(n7336) );
  INV_X1 U8811 ( .A(n7336), .ZN(n7337) );
  OAI21_X1 U8812 ( .B1(n7338), .B2(n11115), .A(n7337), .ZN(P1_U3524) );
  INV_X1 U8813 ( .A(n7339), .ZN(n7341) );
  INV_X1 U8814 ( .A(n9271), .ZN(n7340) );
  NAND2_X1 U8815 ( .A1(n7341), .A2(n7340), .ZN(n7346) );
  NAND2_X1 U8816 ( .A1(n7342), .A2(n9268), .ZN(n7343) );
  NAND2_X2 U8817 ( .A1(n7346), .A2(n7345), .ZN(n7550) );
  NAND2_X1 U8818 ( .A1(n8959), .A2(n7560), .ZN(n7347) );
  NAND2_X1 U8819 ( .A1(n9121), .A2(n7347), .ZN(n7482) );
  NAND2_X1 U8820 ( .A1(n7480), .A2(n7482), .ZN(n7481) );
  INV_X1 U8821 ( .A(n7348), .ZN(n7349) );
  NAND2_X1 U8822 ( .A1(n7349), .A2(n6399), .ZN(n7350) );
  NAND2_X1 U8823 ( .A1(n7481), .A2(n7350), .ZN(n7612) );
  INV_X1 U8824 ( .A(n9335), .ZN(n7554) );
  XNOR2_X1 U8825 ( .A(n7547), .B(n7554), .ZN(n7548) );
  XNOR2_X1 U8826 ( .A(n7612), .B(n7548), .ZN(n7374) );
  INV_X1 U8827 ( .A(n7362), .ZN(n7352) );
  NAND2_X1 U8828 ( .A1(n7352), .A2(n7351), .ZN(n7356) );
  INV_X1 U8829 ( .A(n7353), .ZN(n7354) );
  NAND2_X1 U8830 ( .A1(n7354), .A2(n7368), .ZN(n7355) );
  NAND2_X1 U8831 ( .A1(n7356), .A2(n7355), .ZN(n7367) );
  INV_X1 U8832 ( .A(n7357), .ZN(n7358) );
  NAND2_X1 U8833 ( .A1(n9334), .A2(n10944), .ZN(n7360) );
  NAND2_X1 U8834 ( .A1(n6408), .A2(n9961), .ZN(n7359) );
  NAND2_X1 U8835 ( .A1(n7360), .A2(n7359), .ZN(n10969) );
  NAND2_X1 U8836 ( .A1(n7362), .A2(n7363), .ZN(n7364) );
  AOI22_X1 U8837 ( .A1(n8568), .A2(n10969), .B1(n9059), .B2(n10977), .ZN(n7373) );
  NAND3_X1 U8838 ( .A1(n7759), .A2(n8266), .A3(n7365), .ZN(n7366) );
  OAI21_X1 U8839 ( .B1(n7367), .B2(n7366), .A(P2_STATE_REG_SCAN_IN), .ZN(n7371) );
  INV_X1 U8840 ( .A(n7368), .ZN(n7369) );
  OR2_X1 U8841 ( .A1(n9312), .A2(n7369), .ZN(n7370) );
  NAND2_X1 U8842 ( .A1(n9082), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7477) );
  NAND2_X1 U8843 ( .A1(n7477), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7372) );
  OAI211_X1 U8844 ( .C1(n7374), .C2(n9061), .A(n7373), .B(n7372), .ZN(P2_U3177) );
  XNOR2_X1 U8845 ( .A(n7375), .B(n8788), .ZN(n11011) );
  NAND2_X1 U8846 ( .A1(n7376), .A2(n8667), .ZN(n7380) );
  NOR2_X1 U8847 ( .A1(n8667), .A2(n5370), .ZN(n7377) );
  AOI21_X1 U8848 ( .B1(n7590), .B2(n7377), .A(n10929), .ZN(n7379) );
  OAI22_X1 U8849 ( .A1(n7751), .A2(n8944), .B1(n7462), .B2(n8353), .ZN(n7378)
         );
  AOI21_X1 U8850 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n11026) );
  INV_X1 U8851 ( .A(n7381), .ZN(n7662) );
  OAI211_X1 U8852 ( .C1(n7384), .C2(n7598), .A(n7662), .B(n10599), .ZN(n11020)
         );
  OAI211_X1 U8853 ( .C1(n11011), .C2(n11000), .A(n11026), .B(n11020), .ZN(
        n7386) );
  NAND2_X1 U8854 ( .A1(n7386), .A2(n11120), .ZN(n7383) );
  NAND2_X1 U8855 ( .A1(n8213), .A2(n11017), .ZN(n7382) );
  OAI211_X1 U8856 ( .C1(n11120), .C2(n5829), .A(n7383), .B(n7382), .ZN(
        P1_U3468) );
  OAI22_X1 U8857 ( .A1(n10592), .A2(n7384), .B1(n11116), .B2(n7238), .ZN(n7385) );
  AOI21_X1 U8858 ( .B1(n7386), .B2(n11116), .A(n7385), .ZN(n7387) );
  INV_X1 U8859 ( .A(n7387), .ZN(P1_U3527) );
  INV_X1 U8860 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7389) );
  INV_X1 U8861 ( .A(n7388), .ZN(n7390) );
  INV_X1 U8862 ( .A(n9371), .ZN(n8601) );
  OAI222_X1 U8863 ( .A1(n8985), .A2(n7389), .B1(n8998), .B2(n7390), .C1(n8601), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  INV_X1 U8864 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7391) );
  OAI222_X1 U8865 ( .A1(n10659), .A2(n7391), .B1(n7742), .B2(n7390), .C1(n8029), .C2(P1_U3086), .ZN(P1_U3340) );
  AOI21_X1 U8866 ( .B1(n7393), .B2(P2_REG1_REG_1__SCAN_IN), .A(n7392), .ZN(
        n10882) );
  NAND2_X1 U8867 ( .A1(P2_REG1_REG_2__SCAN_IN), .A2(n10886), .ZN(n7394) );
  OAI21_X1 U8868 ( .B1(n10886), .B2(P2_REG1_REG_2__SCAN_IN), .A(n7394), .ZN(
        n10881) );
  NOR2_X1 U8869 ( .A1(n7412), .A2(n7396), .ZN(n7397) );
  AOI22_X1 U8870 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n7410), .B1(n7520), .B2(
        n6434), .ZN(n7398) );
  NOR2_X1 U8871 ( .A1(n7399), .A2(n7398), .ZN(n7512) );
  AOI21_X1 U8872 ( .B1(n7399), .B2(n7398), .A(n7512), .ZN(n7400) );
  NOR2_X1 U8873 ( .A1(n10915), .A2(n7400), .ZN(n7429) );
  INV_X1 U8874 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7538) );
  INV_X1 U8875 ( .A(n10886), .ZN(n7401) );
  NAND2_X1 U8876 ( .A1(n7401), .A2(n7414), .ZN(n7402) );
  INV_X1 U8877 ( .A(n7403), .ZN(n7404) );
  NOR2_X2 U8878 ( .A1(n10875), .A2(n7407), .ZN(n7408) );
  NOR2_X1 U8879 ( .A1(n7412), .A2(n7408), .ZN(n7409) );
  AOI22_X1 U8880 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n7410), .B1(n7520), .B2(
        n6436), .ZN(n7411) );
  AOI21_X1 U8881 ( .B1(n5193), .B2(n7411), .A(n7517), .ZN(n7427) );
  MUX2_X1 U8882 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9412), .Z(n7521) );
  XNOR2_X1 U8883 ( .A(n7521), .B(n7520), .ZN(n7423) );
  MUX2_X1 U8884 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9412), .Z(n7421) );
  XNOR2_X1 U8885 ( .A(n7421), .B(n7412), .ZN(n7534) );
  MUX2_X1 U8886 ( .A(n7414), .B(n7413), .S(n9412), .Z(n7415) );
  AOI21_X1 U8887 ( .B1(n7401), .B2(n7415), .A(n7420), .ZN(n10869) );
  INV_X1 U8888 ( .A(n7416), .ZN(n7419) );
  OAI21_X1 U8889 ( .B1(n7419), .B2(n7418), .A(n7417), .ZN(n10868) );
  AND2_X1 U8890 ( .A1(n10869), .A2(n10868), .ZN(n10870) );
  NOR2_X1 U8891 ( .A1(n7420), .A2(n10870), .ZN(n7533) );
  NAND2_X1 U8892 ( .A1(n7534), .A2(n7533), .ZN(n7532) );
  NOR2_X1 U8893 ( .A1(n7423), .A2(n7422), .ZN(n7519) );
  AOI211_X1 U8894 ( .C1(n7423), .C2(n7422), .A(n9426), .B(n7519), .ZN(n7424)
         );
  INV_X1 U8895 ( .A(n7424), .ZN(n7426) );
  NAND2_X1 U8896 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3151), .ZN(n7425) );
  OAI211_X1 U8897 ( .C1(n7427), .C2(n10918), .A(n7426), .B(n7425), .ZN(n7428)
         );
  AOI211_X1 U8898 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10907), .A(n7429), .B(
        n7428), .ZN(n7430) );
  OAI21_X1 U8899 ( .B1(n7520), .B2(n10904), .A(n7430), .ZN(P2_U3186) );
  NAND2_X1 U8900 ( .A1(n7433), .A2(n7432), .ZN(n7435) );
  XNOR2_X1 U8901 ( .A(n7435), .B(n7434), .ZN(n7438) );
  AOI22_X1 U8902 ( .A1(n10189), .A2(n6858), .B1(n11091), .B2(n10213), .ZN(
        n7437) );
  AOI22_X1 U8903 ( .A1(n11088), .A2(n5122), .B1(n7441), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7436) );
  OAI211_X1 U8904 ( .C1(n7438), .C2(n10199), .A(n7437), .B(n7436), .ZN(
        P1_U3222) );
  XOR2_X1 U8905 ( .A(n7440), .B(n7439), .Z(n7444) );
  AOI22_X1 U8906 ( .A1(n10189), .A2(n10214), .B1(n11091), .B2(n10212), .ZN(
        n7443) );
  AOI22_X1 U8907 ( .A1(n11088), .A2(n7704), .B1(n7441), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7442) );
  OAI211_X1 U8908 ( .C1(n7444), .C2(n10199), .A(n7443), .B(n7442), .ZN(
        P1_U3237) );
  INV_X1 U8909 ( .A(n10616), .ZN(n11054) );
  INV_X1 U8910 ( .A(n7445), .ZN(n7446) );
  INV_X1 U8911 ( .A(n7579), .ZN(n7457) );
  INV_X1 U8912 ( .A(n7448), .ZN(n7583) );
  NAND2_X1 U8913 ( .A1(n5122), .A2(n10932), .ZN(n7582) );
  NAND3_X1 U8914 ( .A1(n7583), .A2(n10599), .A3(n7582), .ZN(n7449) );
  OAI21_X1 U8915 ( .B1(n8864), .B2(n11109), .A(n7449), .ZN(n7456) );
  OAI22_X1 U8916 ( .A1(n7461), .A2(n8944), .B1(n6861), .B2(n8353), .ZN(n7453)
         );
  NOR2_X1 U8917 ( .A1(n7579), .A2(n8359), .ZN(n7452) );
  AOI211_X1 U8918 ( .C1(n10512), .C2(n7454), .A(n7453), .B(n7452), .ZN(n7586)
         );
  INV_X1 U8919 ( .A(n7586), .ZN(n7455) );
  AOI211_X1 U8920 ( .C1(n11054), .C2(n7457), .A(n7456), .B(n7455), .ZN(n10961)
         );
  NAND2_X1 U8921 ( .A1(n11115), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7458) );
  OAI21_X1 U8922 ( .B1(n10961), .B2(n11115), .A(n7458), .ZN(P1_U3523) );
  INV_X1 U8923 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7473) );
  OAI21_X1 U8924 ( .B1(n7460), .B2(n7464), .A(n7459), .ZN(n7779) );
  INV_X1 U8925 ( .A(n7779), .ZN(n7470) );
  INV_X1 U8926 ( .A(n8359), .ZN(n7656) );
  OAI22_X1 U8927 ( .A1(n7462), .A2(n8944), .B1(n7461), .B2(n8353), .ZN(n7467)
         );
  INV_X1 U8928 ( .A(n8665), .ZN(n7463) );
  INV_X1 U8929 ( .A(n7464), .ZN(n8785) );
  NAND2_X1 U8930 ( .A1(n7463), .A2(n8785), .ZN(n7592) );
  NAND2_X1 U8931 ( .A1(n8665), .A2(n7464), .ZN(n7465) );
  AOI21_X1 U8932 ( .B1(n7592), .B2(n7465), .A(n10929), .ZN(n7466) );
  AOI211_X1 U8933 ( .C1(n7656), .C2(n7779), .A(n7467), .B(n7466), .ZN(n7782)
         );
  AOI21_X1 U8934 ( .B1(n7468), .B2(n7773), .A(n11049), .ZN(n7469) );
  NAND2_X1 U8935 ( .A1(n7469), .A2(n7599), .ZN(n7777) );
  OAI211_X1 U8936 ( .C1(n7470), .C2(n10616), .A(n7782), .B(n7777), .ZN(n7475)
         );
  NAND2_X1 U8937 ( .A1(n7475), .A2(n11120), .ZN(n7472) );
  NAND2_X1 U8938 ( .A1(n8213), .A2(n7773), .ZN(n7471) );
  OAI211_X1 U8939 ( .C1(n11120), .C2(n7473), .A(n7472), .B(n7471), .ZN(
        P1_U3462) );
  OAI22_X1 U8940 ( .A1(n10592), .A2(n7489), .B1(n11116), .B2(n7234), .ZN(n7474) );
  AOI21_X1 U8941 ( .B1(n7475), .B2(n11116), .A(n7474), .ZN(n7476) );
  INV_X1 U8942 ( .A(n7476), .ZN(P1_U3525) );
  INV_X1 U8943 ( .A(n7477), .ZN(n7563) );
  NAND2_X1 U8944 ( .A1(n9335), .A2(n10944), .ZN(n7479) );
  NAND2_X1 U8945 ( .A1(n9337), .A2(n9961), .ZN(n7478) );
  NAND2_X1 U8946 ( .A1(n7479), .A2(n7478), .ZN(n8070) );
  AOI22_X1 U8947 ( .A1(n8568), .A2(n8070), .B1(n9059), .B2(n6398), .ZN(n7485)
         );
  OAI21_X1 U8948 ( .B1(n7480), .B2(n7482), .A(n7481), .ZN(n7483) );
  NAND2_X1 U8949 ( .A1(n7483), .A2(n9076), .ZN(n7484) );
  OAI211_X1 U8950 ( .C1(n7563), .C2(n8072), .A(n7485), .B(n7484), .ZN(P2_U3162) );
  XOR2_X1 U8951 ( .A(n7488), .B(n7487), .Z(n7494) );
  INV_X1 U8952 ( .A(n11101), .ZN(n10190) );
  NAND2_X1 U8953 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10247) );
  INV_X1 U8954 ( .A(n10247), .ZN(n7491) );
  NOR2_X1 U8955 ( .A1(n10183), .A2(n7489), .ZN(n7490) );
  AOI211_X1 U8956 ( .C1(n7774), .C2(n10190), .A(n7491), .B(n7490), .ZN(n7493)
         );
  AOI22_X1 U8957 ( .A1(n11091), .A2(n10211), .B1(n10189), .B2(n10213), .ZN(
        n7492) );
  OAI211_X1 U8958 ( .C1(n10199), .C2(n7494), .A(n7493), .B(n7492), .ZN(
        P1_U3218) );
  INV_X1 U8959 ( .A(n7496), .ZN(n7497) );
  AOI211_X1 U8960 ( .C1(n7498), .C2(n7495), .A(n10199), .B(n7497), .ZN(n7502)
         );
  AOI22_X1 U8961 ( .A1(n10189), .A2(n10212), .B1(n11091), .B2(n10210), .ZN(
        n7500) );
  AND2_X1 U8962 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10262) );
  AOI21_X1 U8963 ( .B1(n11088), .B2(n10995), .A(n10262), .ZN(n7499) );
  OAI211_X1 U8964 ( .C1(n11101), .C2(n7600), .A(n7500), .B(n7499), .ZN(n7501)
         );
  OR2_X1 U8965 ( .A1(n7502), .A2(n7501), .ZN(P1_U3230) );
  NAND2_X1 U8966 ( .A1(n7504), .A2(n7503), .ZN(n7506) );
  XNOR2_X1 U8967 ( .A(n7506), .B(n7505), .ZN(n7511) );
  AOI22_X1 U8968 ( .A1(n11091), .A2(n10209), .B1(n10189), .B2(n10211), .ZN(
        n7510) );
  NAND2_X1 U8969 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10273) );
  INV_X1 U8970 ( .A(n10273), .ZN(n7508) );
  NOR2_X1 U8971 ( .A1(n11101), .A2(n11013), .ZN(n7507) );
  AOI211_X1 U8972 ( .C1(n11017), .C2(n11088), .A(n7508), .B(n7507), .ZN(n7509)
         );
  OAI211_X1 U8973 ( .C1(n7511), .C2(n10199), .A(n7510), .B(n7509), .ZN(
        P1_U3227) );
  AOI21_X1 U8974 ( .B1(n6445), .B2(n7513), .A(n7694), .ZN(n7515) );
  NAND2_X1 U8975 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3151), .ZN(n7514) );
  OAI21_X1 U8976 ( .B1(n7515), .B2(n10915), .A(n7514), .ZN(n7528) );
  NOR2_X2 U8977 ( .A1(n7517), .A2(n7516), .ZN(n7676) );
  AOI21_X1 U8978 ( .B1(n6448), .B2(n7518), .A(n7677), .ZN(n7526) );
  MUX2_X1 U8979 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n9412), .Z(n7684) );
  XNOR2_X1 U8980 ( .A(n7684), .B(n7683), .ZN(n7523) );
  NOR2_X1 U8981 ( .A1(n7522), .A2(n7523), .ZN(n7682) );
  AOI211_X1 U8982 ( .C1(n7523), .C2(n7522), .A(n9426), .B(n7682), .ZN(n7524)
         );
  INV_X1 U8983 ( .A(n7524), .ZN(n7525) );
  OAI21_X1 U8984 ( .B1(n7526), .B2(n10918), .A(n7525), .ZN(n7527) );
  AOI211_X1 U8985 ( .C1(n10907), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7528), .B(
        n7527), .ZN(n7529) );
  OAI21_X1 U8986 ( .B1(n7683), .B2(n10904), .A(n7529), .ZN(P2_U3187) );
  AOI21_X1 U8987 ( .B1(n7531), .B2(n6421), .A(n7530), .ZN(n7543) );
  OAI21_X1 U8988 ( .B1(n7534), .B2(n7533), .A(n7532), .ZN(n7541) );
  INV_X1 U8989 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7535) );
  NOR2_X1 U8990 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7535), .ZN(n7556) );
  AOI21_X1 U8991 ( .B1(n7538), .B2(n7536), .A(n7537), .ZN(n7539) );
  NOR2_X1 U8992 ( .A1(n10918), .A2(n7539), .ZN(n7540) );
  AOI211_X1 U8993 ( .C1(n10923), .C2(n7541), .A(n7556), .B(n7540), .ZN(n7542)
         );
  OAI21_X1 U8994 ( .B1(n7543), .B2(n10915), .A(n7542), .ZN(n7544) );
  AOI21_X1 U8995 ( .B1(n10907), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7544), .ZN(
        n7545) );
  OAI21_X1 U8996 ( .B1(n7546), .B2(n10904), .A(n7545), .ZN(P2_U3185) );
  INV_X1 U8997 ( .A(n7612), .ZN(n7549) );
  OAI21_X1 U8998 ( .B1(n7549), .B2(n7548), .A(n7605), .ZN(n7552) );
  XNOR2_X1 U8999 ( .A(n7550), .B(n10982), .ZN(n7609) );
  INV_X1 U9000 ( .A(n9334), .ZN(n7880) );
  XNOR2_X1 U9001 ( .A(n7609), .B(n7880), .ZN(n7551) );
  XNOR2_X1 U9002 ( .A(n7552), .B(n7551), .ZN(n7553) );
  NAND2_X1 U9003 ( .A1(n7553), .A2(n9076), .ZN(n7559) );
  NOR2_X2 U9004 ( .A1(n9019), .A2(n9875), .ZN(n9080) );
  INV_X1 U9005 ( .A(n9080), .ZN(n7643) );
  INV_X1 U9006 ( .A(n9333), .ZN(n8084) );
  NAND2_X1 U9007 ( .A1(n8568), .A2(n9875), .ZN(n9067) );
  OAI22_X1 U9008 ( .A1(n7643), .A2(n8084), .B1(n7554), .B2(n9067), .ZN(n7555)
         );
  AOI211_X1 U9009 ( .C1(n7557), .C2(n9059), .A(n7556), .B(n7555), .ZN(n7558)
         );
  OAI211_X1 U9010 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9082), .A(n7559), .B(
        n7558), .ZN(P2_U3158) );
  NAND2_X1 U9011 ( .A1(n9337), .A2(n7560), .ZN(n9124) );
  NAND2_X1 U9012 ( .A1(n9121), .A2(n9124), .ZN(n10937) );
  INV_X1 U9013 ( .A(n9059), .ZN(n9088) );
  OAI22_X1 U9014 ( .A1(n7643), .A2(n6399), .B1(n9088), .B2(n7560), .ZN(n7561)
         );
  AOI21_X1 U9015 ( .B1(n9076), .B2(n10937), .A(n7561), .ZN(n7562) );
  OAI21_X1 U9016 ( .B1(n7563), .B2(n10951), .A(n7562), .ZN(P2_U3172) );
  INV_X1 U9017 ( .A(n7564), .ZN(n7566) );
  NAND3_X1 U9018 ( .A1(n7567), .A2(n7566), .A3(n7565), .ZN(n7568) );
  NOR2_X1 U9019 ( .A1(n11021), .A2(n11049), .ZN(n10454) );
  OAI21_X1 U9020 ( .B1(n10454), .B2(n11018), .A(n10932), .ZN(n7575) );
  XNOR2_X1 U9021 ( .A(n6861), .B(n7570), .ZN(n10928) );
  INV_X1 U9022 ( .A(n7571), .ZN(n8849) );
  OR3_X1 U9023 ( .A1(n10928), .A2(n8849), .A3(n10933), .ZN(n7572) );
  NAND2_X1 U9024 ( .A1(n10214), .A2(n10509), .ZN(n10927) );
  OAI211_X1 U9025 ( .C1(n5737), .C2(n11012), .A(n7572), .B(n10927), .ZN(n7573)
         );
  NAND2_X1 U9026 ( .A1(n11015), .A2(n7573), .ZN(n7574) );
  OAI211_X1 U9027 ( .C1(n10750), .C2(n11015), .A(n7575), .B(n7574), .ZN(
        P1_U3293) );
  NAND2_X1 U9028 ( .A1(n10529), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7576) );
  OAI21_X1 U9029 ( .B1(n5748), .B2(n11012), .A(n7576), .ZN(n7581) );
  OR2_X1 U9030 ( .A1(n7577), .A2(n8259), .ZN(n7578) );
  NOR2_X1 U9031 ( .A1(n8368), .A2(n7579), .ZN(n7580) );
  AOI211_X1 U9032 ( .C1(n11018), .C2(n5122), .A(n7581), .B(n7580), .ZN(n7585)
         );
  NAND3_X1 U9033 ( .A1(n10454), .A2(n7583), .A3(n7582), .ZN(n7584) );
  OAI211_X1 U9034 ( .C1(n7586), .C2(n10466), .A(n7585), .B(n7584), .ZN(
        P1_U3292) );
  OR2_X1 U9035 ( .A1(n10529), .A2(n8359), .ZN(n7587) );
  NAND2_X1 U9036 ( .A1(n8666), .A2(n8671), .ZN(n8787) );
  XOR2_X1 U9037 ( .A(n8787), .B(n7588), .Z(n10999) );
  NOR2_X1 U9038 ( .A1(n7589), .A2(n8944), .ZN(n7596) );
  INV_X1 U9039 ( .A(n7590), .ZN(n7594) );
  INV_X1 U9040 ( .A(n8787), .ZN(n7591) );
  AOI21_X1 U9041 ( .B1(n7592), .B2(n8871), .A(n7591), .ZN(n7593) );
  AOI211_X1 U9042 ( .C1(n7594), .C2(n8666), .A(n10929), .B(n7593), .ZN(n7595)
         );
  AOI211_X1 U9043 ( .C1(n10507), .C2(n10212), .A(n7596), .B(n7595), .ZN(n10998) );
  MUX2_X1 U9044 ( .A(n7597), .B(n10998), .S(n11015), .Z(n7604) );
  AOI211_X1 U9045 ( .C1(n10995), .C2(n7599), .A(n11049), .B(n7598), .ZN(n10994) );
  OAI22_X1 U9046 ( .A1(n10525), .A2(n7601), .B1(n7600), .B2(n11012), .ZN(n7602) );
  AOI21_X1 U9047 ( .B1(n10520), .B2(n10994), .A(n7602), .ZN(n7603) );
  OAI211_X1 U9048 ( .C1(n10504), .C2(n10999), .A(n7604), .B(n7603), .ZN(
        P1_U3289) );
  OAI21_X1 U9049 ( .B1(n7609), .B2(n9334), .A(n7605), .ZN(n7613) );
  NAND2_X1 U9050 ( .A1(n7606), .A2(n7880), .ZN(n7610) );
  AND2_X1 U9051 ( .A1(n9334), .A2(n9335), .ZN(n7607) );
  AOI22_X1 U9052 ( .A1(n7610), .A2(n7609), .B1(n7608), .B2(n7607), .ZN(n7611)
         );
  OAI21_X1 U9053 ( .B1(n7613), .B2(n7612), .A(n7611), .ZN(n7614) );
  XNOR2_X1 U9054 ( .A(n7550), .B(n7635), .ZN(n7615) );
  XNOR2_X1 U9055 ( .A(n7615), .B(n9333), .ZN(n7633) );
  NAND2_X1 U9056 ( .A1(n7634), .A2(n7633), .ZN(n7632) );
  NAND2_X1 U9057 ( .A1(n7615), .A2(n8084), .ZN(n7616) );
  NAND2_X1 U9058 ( .A1(n7632), .A2(n7616), .ZN(n7722) );
  INV_X1 U9059 ( .A(n7722), .ZN(n7618) );
  XNOR2_X1 U9060 ( .A(n7550), .B(n7617), .ZN(n7724) );
  INV_X1 U9061 ( .A(n9332), .ZN(n7881) );
  XNOR2_X1 U9062 ( .A(n7724), .B(n7881), .ZN(n7641) );
  NAND2_X1 U9063 ( .A1(n7724), .A2(n7881), .ZN(n7723) );
  OAI21_X1 U9064 ( .B1(n7618), .B2(n7641), .A(n7723), .ZN(n7620) );
  XNOR2_X1 U9065 ( .A(n7769), .B(n7550), .ZN(n7726) );
  INV_X1 U9066 ( .A(n9331), .ZN(n8083) );
  XNOR2_X1 U9067 ( .A(n7726), .B(n8083), .ZN(n7619) );
  XNOR2_X1 U9068 ( .A(n7620), .B(n7619), .ZN(n7628) );
  INV_X1 U9069 ( .A(n9082), .ZN(n9071) );
  INV_X1 U9070 ( .A(n7621), .ZN(n7768) );
  NAND2_X1 U9071 ( .A1(n9330), .A2(n10944), .ZN(n7623) );
  NAND2_X1 U9072 ( .A1(n9332), .A2(n9961), .ZN(n7622) );
  NAND2_X1 U9073 ( .A1(n7623), .A2(n7622), .ZN(n7715) );
  AOI22_X1 U9074 ( .A1(n7715), .A2(n8568), .B1(P2_REG3_REG_6__SCAN_IN), .B2(
        P2_U3151), .ZN(n7624) );
  OAI21_X1 U9075 ( .B1(n7625), .B2(n9088), .A(n7624), .ZN(n7626) );
  AOI21_X1 U9076 ( .B1(n9071), .B2(n7768), .A(n7626), .ZN(n7627) );
  OAI21_X1 U9077 ( .B1(n7628), .B2(n9061), .A(n7627), .ZN(P2_U3179) );
  INV_X1 U9078 ( .A(n7629), .ZN(n7630) );
  INV_X1 U9079 ( .A(n8120), .ZN(n8024) );
  OAI222_X1 U9080 ( .A1(n10659), .A2(n9797), .B1(n7742), .B2(n7630), .C1(
        P1_U3086), .C2(n8024), .ZN(P1_U3339) );
  OAI222_X1 U9081 ( .A1(n8985), .A2(n7631), .B1(n8998), .B2(n7630), .C1(
        P2_U3151), .C2(n9380), .ZN(P2_U3279) );
  OAI21_X1 U9082 ( .B1(n7634), .B2(n7633), .A(n7632), .ZN(n7639) );
  AOI22_X1 U9083 ( .A1(n9059), .A2(n7635), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3151), .ZN(n7637) );
  AOI22_X1 U9084 ( .A1(n9085), .A2(n9334), .B1(n9080), .B2(n9332), .ZN(n7636)
         );
  OAI211_X1 U9085 ( .C1(n9082), .C2(n7882), .A(n7637), .B(n7636), .ZN(n7638)
         );
  AOI21_X1 U9086 ( .B1(n7639), .B2(n9076), .A(n7638), .ZN(n7640) );
  INV_X1 U9087 ( .A(n7640), .ZN(P2_U3170) );
  XNOR2_X1 U9088 ( .A(n7722), .B(n7641), .ZN(n7648) );
  INV_X1 U9089 ( .A(n8089), .ZN(n7646) );
  OAI22_X1 U9090 ( .A1(n9088), .A2(n11004), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7642), .ZN(n7645) );
  OAI22_X1 U9091 ( .A1(n7643), .A2(n8083), .B1(n8084), .B2(n9067), .ZN(n7644)
         );
  AOI211_X1 U9092 ( .C1(n9071), .C2(n7646), .A(n7645), .B(n7644), .ZN(n7647)
         );
  OAI21_X1 U9093 ( .B1(n7648), .B2(n9061), .A(n7647), .ZN(P2_U3167) );
  INV_X1 U9094 ( .A(n7649), .ZN(n7650) );
  INV_X1 U9095 ( .A(n8249), .ZN(n8123) );
  OAI222_X1 U9096 ( .A1(n10659), .A2(n9793), .B1(n7742), .B2(n7650), .C1(n8123), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U9097 ( .A(n8618), .ZN(n9396) );
  OAI222_X1 U9098 ( .A1(n8985), .A2(n7651), .B1(n8998), .B2(n7650), .C1(n9396), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  OR2_X1 U9099 ( .A1(n7653), .A2(n7652), .ZN(n7654) );
  NAND2_X1 U9100 ( .A1(n7655), .A2(n7654), .ZN(n11032) );
  INV_X1 U9101 ( .A(n11032), .ZN(n7666) );
  XNOR2_X1 U9102 ( .A(n7748), .B(n8674), .ZN(n7659) );
  NAND2_X1 U9103 ( .A1(n11032), .A2(n7656), .ZN(n7658) );
  AOI22_X1 U9104 ( .A1(n10509), .A2(n10208), .B1(n10210), .B2(n10507), .ZN(
        n7657) );
  OAI211_X1 U9105 ( .C1(n10929), .C2(n7659), .A(n7658), .B(n7657), .ZN(n11030)
         );
  MUX2_X1 U9106 ( .A(n11030), .B(P1_REG2_REG_6__SCAN_IN), .S(n10529), .Z(n7660) );
  INV_X1 U9107 ( .A(n7660), .ZN(n7665) );
  INV_X1 U9108 ( .A(n7747), .ZN(n7661) );
  AOI211_X1 U9109 ( .C1(n10166), .C2(n7662), .A(n11049), .B(n7661), .ZN(n11027) );
  OAI22_X1 U9110 ( .A1(n10525), .A2(n11029), .B1(n10168), .B2(n11012), .ZN(
        n7663) );
  AOI21_X1 U9111 ( .B1(n11027), .B2(n10520), .A(n7663), .ZN(n7664) );
  OAI211_X1 U9112 ( .C1(n7666), .C2(n8368), .A(n7665), .B(n7664), .ZN(P1_U3287) );
  XNOR2_X1 U9113 ( .A(n7668), .B(n7667), .ZN(n7669) );
  XNOR2_X1 U9114 ( .A(n7670), .B(n7669), .ZN(n7675) );
  INV_X1 U9115 ( .A(n7671), .ZN(n7786) );
  AOI22_X1 U9116 ( .A1(n7786), .A2(n10190), .B1(n10189), .B2(n10209), .ZN(
        n7672) );
  NAND2_X1 U9117 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10299) );
  OAI211_X1 U9118 ( .C1(n7752), .C2(n10194), .A(n7672), .B(n10299), .ZN(n7673)
         );
  AOI21_X1 U9119 ( .B1(n7784), .B2(n11088), .A(n7673), .ZN(n7674) );
  OAI21_X1 U9120 ( .B1(n7675), .B2(n10199), .A(n7674), .ZN(P1_U3213) );
  NOR2_X1 U9121 ( .A1(n7693), .A2(n7676), .ZN(n7678) );
  AOI22_X1 U9122 ( .A1(n7696), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7679), .B2(
        n10903), .ZN(n10892) );
  NOR2_X1 U9123 ( .A1(n7696), .A2(n7679), .ZN(n7680) );
  AOI21_X1 U9124 ( .B1(n6476), .B2(n7681), .A(n7986), .ZN(n7701) );
  MUX2_X1 U9125 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n9412), .Z(n7685) );
  XNOR2_X1 U9126 ( .A(n7685), .B(n7696), .ZN(n10888) );
  NAND2_X1 U9127 ( .A1(n10889), .A2(n10888), .ZN(n10887) );
  OAI21_X1 U9128 ( .B1(n7685), .B2(n10903), .A(n10887), .ZN(n7687) );
  MUX2_X1 U9129 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n9412), .Z(n7991) );
  XNOR2_X1 U9130 ( .A(n7991), .B(n8001), .ZN(n7686) );
  NAND2_X1 U9131 ( .A1(n7687), .A2(n7686), .ZN(n7992) );
  OAI21_X1 U9132 ( .B1(n7687), .B2(n7686), .A(n7992), .ZN(n7691) );
  INV_X1 U9133 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7736) );
  OAI22_X1 U9134 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7736), .B1(n10904), .B2(
        n7990), .ZN(n7690) );
  INV_X1 U9135 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7688) );
  NOR2_X1 U9136 ( .A1(n9422), .A2(n7688), .ZN(n7689) );
  AOI211_X1 U9137 ( .C1(n7691), .C2(n10923), .A(n7690), .B(n7689), .ZN(n7700)
         );
  NOR2_X1 U9138 ( .A1(n7693), .A2(n7692), .ZN(n7695) );
  AOI22_X1 U9139 ( .A1(n7696), .A2(P2_REG1_REG_6__SCAN_IN), .B1(n6459), .B2(
        n10903), .ZN(n10895) );
  NOR2_X1 U9140 ( .A1(n10896), .A2(n10895), .ZN(n10894) );
  XNOR2_X1 U9141 ( .A(n8000), .B(n8001), .ZN(n7697) );
  NOR2_X1 U9142 ( .A1(n6475), .A2(n7697), .ZN(n8002) );
  AOI21_X1 U9143 ( .B1(n7697), .B2(n6475), .A(n8002), .ZN(n7698) );
  OR2_X1 U9144 ( .A1(n7698), .A2(n10915), .ZN(n7699) );
  OAI211_X1 U9145 ( .C1(n7701), .C2(n10918), .A(n7700), .B(n7699), .ZN(
        P2_U3189) );
  INV_X1 U9146 ( .A(n11012), .ZN(n10521) );
  AOI211_X1 U9147 ( .C1(n10521), .C2(P1_REG3_REG_2__SCAN_IN), .A(n7703), .B(
        n7702), .ZN(n7710) );
  AOI22_X1 U9148 ( .A1(n11018), .A2(n7704), .B1(n10529), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n7705) );
  OAI21_X1 U9149 ( .B1(n11021), .B2(n7706), .A(n7705), .ZN(n7707) );
  AOI21_X1 U9150 ( .B1(n11023), .B2(n7708), .A(n7707), .ZN(n7709) );
  OAI21_X1 U9151 ( .B1(n10529), .B2(n7710), .A(n7709), .ZN(P1_U3291) );
  INV_X1 U9152 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7719) );
  OAI21_X1 U9153 ( .B1(n7713), .B2(n7712), .A(n7711), .ZN(n7758) );
  AOI22_X1 U9154 ( .A1(n7758), .A2(n11132), .B1(n11151), .B2(n7769), .ZN(n7717) );
  XNOR2_X1 U9155 ( .A(n7714), .B(n9278), .ZN(n7716) );
  AOI21_X1 U9156 ( .B1(n7716), .B2(n10935), .A(n7715), .ZN(n7767) );
  NAND2_X1 U9157 ( .A1(n7717), .A2(n7767), .ZN(n7720) );
  NAND2_X1 U9158 ( .A1(n7720), .A2(n11157), .ZN(n7718) );
  OAI21_X1 U9159 ( .B1(n7719), .B2(n11157), .A(n7718), .ZN(P2_U3408) );
  NAND2_X1 U9160 ( .A1(n7720), .A2(n11153), .ZN(n7721) );
  OAI21_X1 U9161 ( .B1(n11153), .B2(n6459), .A(n7721), .ZN(P2_U3465) );
  NAND2_X1 U9162 ( .A1(n7726), .A2(n8083), .ZN(n7729) );
  INV_X1 U9163 ( .A(n7724), .ZN(n7725) );
  AND2_X1 U9164 ( .A1(n7725), .A2(n9332), .ZN(n7728) );
  INV_X1 U9165 ( .A(n7726), .ZN(n7727) );
  XNOR2_X1 U9166 ( .A(n7732), .B(n7550), .ZN(n7813) );
  INV_X1 U9167 ( .A(n9330), .ZN(n7818) );
  XNOR2_X1 U9168 ( .A(n7813), .B(n7818), .ZN(n7733) );
  OAI21_X1 U9169 ( .B1(n7734), .B2(n7733), .A(n7816), .ZN(n7735) );
  NAND2_X1 U9170 ( .A1(n7735), .A2(n9076), .ZN(n7740) );
  OAI22_X1 U9171 ( .A1(n8083), .A2(n8524), .B1(n7896), .B2(n8523), .ZN(n7904)
         );
  INV_X1 U9172 ( .A(n7904), .ZN(n7737) );
  OAI22_X1 U9173 ( .A1(n7737), .A2(n9019), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7736), .ZN(n7738) );
  AOI21_X1 U9174 ( .B1(n11044), .B2(n9059), .A(n7738), .ZN(n7739) );
  OAI211_X1 U9175 ( .C1(n11040), .C2(n9082), .A(n7740), .B(n7739), .ZN(
        P2_U3153) );
  INV_X1 U9176 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7743) );
  INV_X1 U9177 ( .A(n7741), .ZN(n7756) );
  INV_X1 U9178 ( .A(n8253), .ZN(n10828) );
  OAI222_X1 U9179 ( .A1(n10659), .A2(n7743), .B1(n7742), .B2(n7756), .C1(
        n10828), .C2(P1_U3086), .ZN(P1_U3337) );
  OAI21_X1 U9180 ( .B1(n7745), .B2(n8680), .A(n7744), .ZN(n7791) );
  INV_X1 U9181 ( .A(n7746), .ZN(n7806) );
  AOI211_X1 U9182 ( .C1(n7784), .C2(n7747), .A(n11049), .B(n7806), .ZN(n7785)
         );
  NAND2_X1 U9183 ( .A1(n7748), .A2(n8790), .ZN(n7749) );
  NAND2_X1 U9184 ( .A1(n7749), .A2(n8676), .ZN(n7796) );
  XOR2_X1 U9185 ( .A(n8680), .B(n7796), .Z(n7750) );
  OAI222_X1 U9186 ( .A1(n8944), .A2(n7752), .B1(n8353), .B2(n7751), .C1(n10929), .C2(n7750), .ZN(n7783) );
  AOI211_X1 U9187 ( .C1(n11113), .C2(n7791), .A(n7785), .B(n7783), .ZN(n7755)
         );
  AOI22_X1 U9188 ( .A1(n8213), .A2(n7784), .B1(n11117), .B2(
        P1_REG0_REG_7__SCAN_IN), .ZN(n7753) );
  OAI21_X1 U9189 ( .B1(n7755), .B2(n11117), .A(n7753), .ZN(P1_U3474) );
  AOI22_X1 U9190 ( .A1(n8211), .A2(n7784), .B1(n11115), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7754) );
  OAI21_X1 U9191 ( .B1(n7755), .B2(n11115), .A(n7754), .ZN(P1_U3529) );
  INV_X1 U9192 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7757) );
  INV_X1 U9193 ( .A(n8595), .ZN(n9417) );
  OAI222_X1 U9194 ( .A1(n8985), .A2(n7757), .B1(P2_U3151), .B2(n9417), .C1(
        n7756), .C2(n8998), .ZN(P2_U3277) );
  INV_X1 U9195 ( .A(n7758), .ZN(n7772) );
  NAND2_X1 U9196 ( .A1(n7759), .A2(n7341), .ZN(n7762) );
  OAI22_X1 U9197 ( .A1(n7763), .A2(n7762), .B1(n7761), .B2(n7760), .ZN(n7765)
         );
  NAND2_X1 U9198 ( .A1(n7765), .A2(n7764), .ZN(n10941) );
  AND2_X1 U9199 ( .A1(n7766), .A2(n7342), .ZN(n8088) );
  OR2_X1 U9200 ( .A1(n8157), .A2(n8088), .ZN(n11036) );
  MUX2_X1 U9201 ( .A(n7679), .B(n7767), .S(n11048), .Z(n7771) );
  AOI22_X1 U9202 ( .A1(n11043), .A2(n7769), .B1(n11041), .B2(n7768), .ZN(n7770) );
  OAI211_X1 U9203 ( .C1(n7772), .C2(n9954), .A(n7771), .B(n7770), .ZN(P2_U3227) );
  INV_X1 U9204 ( .A(n8368), .ZN(n7780) );
  NAND2_X1 U9205 ( .A1(n11018), .A2(n7773), .ZN(n7776) );
  AOI22_X1 U9206 ( .A1(n10466), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10521), .B2(
        n7774), .ZN(n7775) );
  OAI211_X1 U9207 ( .C1(n7777), .C2(n11021), .A(n7776), .B(n7775), .ZN(n7778)
         );
  AOI21_X1 U9208 ( .B1(n7780), .B2(n7779), .A(n7778), .ZN(n7781) );
  OAI21_X1 U9209 ( .B1(n7782), .B2(n10466), .A(n7781), .ZN(P1_U3290) );
  INV_X1 U9210 ( .A(n7783), .ZN(n7793) );
  INV_X1 U9211 ( .A(n7784), .ZN(n7789) );
  NAND2_X1 U9212 ( .A1(n7785), .A2(n10520), .ZN(n7788) );
  AOI22_X1 U9213 ( .A1(n10529), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7786), .B2(
        n10521), .ZN(n7787) );
  OAI211_X1 U9214 ( .C1(n7789), .C2(n10525), .A(n7788), .B(n7787), .ZN(n7790)
         );
  AOI21_X1 U9215 ( .B1(n7791), .B2(n11023), .A(n7790), .ZN(n7792) );
  OAI21_X1 U9216 ( .B1(n7793), .B2(n10466), .A(n7792), .ZN(P1_U3286) );
  OAI21_X1 U9217 ( .B1(n7795), .B2(n8687), .A(n7794), .ZN(n11053) );
  INV_X1 U9218 ( .A(n11053), .ZN(n7812) );
  AOI22_X1 U9219 ( .A1(n10507), .A2(n10208), .B1(n10206), .B2(n10509), .ZN(
        n7803) );
  OR2_X1 U9220 ( .A1(n7796), .A2(n8680), .ZN(n7798) );
  NAND2_X1 U9221 ( .A1(n7798), .A2(n7797), .ZN(n7799) );
  INV_X1 U9222 ( .A(n7799), .ZN(n7801) );
  INV_X1 U9223 ( .A(n8687), .ZN(n7800) );
  OR2_X1 U9224 ( .A1(n7799), .A2(n8687), .ZN(n7841) );
  OAI211_X1 U9225 ( .C1(n7801), .C2(n7800), .A(n7841), .B(n10512), .ZN(n7802)
         );
  OAI211_X1 U9226 ( .C1(n7812), .C2(n8359), .A(n7803), .B(n7802), .ZN(n11051)
         );
  NAND2_X1 U9227 ( .A1(n11051), .A2(n11015), .ZN(n7811) );
  OAI22_X1 U9228 ( .A1(n11015), .A2(n7804), .B1(n7862), .B2(n11012), .ZN(n7809) );
  INV_X1 U9229 ( .A(n7849), .ZN(n7805) );
  OAI21_X1 U9230 ( .B1(n5253), .B2(n7806), .A(n7805), .ZN(n11050) );
  INV_X1 U9231 ( .A(n10454), .ZN(n7807) );
  NOR2_X1 U9232 ( .A1(n11050), .A2(n7807), .ZN(n7808) );
  AOI211_X1 U9233 ( .C1(n11018), .C2(n7866), .A(n7809), .B(n7808), .ZN(n7810)
         );
  OAI211_X1 U9234 ( .C1(n7812), .C2(n8368), .A(n7811), .B(n7810), .ZN(P1_U3285) );
  XNOR2_X1 U9235 ( .A(n7970), .B(n7550), .ZN(n7888) );
  XNOR2_X1 U9236 ( .A(n7888), .B(n9329), .ZN(n7890) );
  INV_X1 U9237 ( .A(n7813), .ZN(n7814) );
  NAND2_X1 U9238 ( .A1(n7814), .A2(n7818), .ZN(n7815) );
  XOR2_X1 U9239 ( .A(n7890), .B(n7891), .Z(n7824) );
  NOR2_X1 U9240 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7817), .ZN(n7996) );
  NOR2_X1 U9241 ( .A1(n9067), .A2(n7818), .ZN(n7819) );
  AOI211_X1 U9242 ( .C1(n9080), .C2(n5260), .A(n7996), .B(n7819), .ZN(n7820)
         );
  OAI21_X1 U9243 ( .B1(n7821), .B2(n9082), .A(n7820), .ZN(n7822) );
  AOI21_X1 U9244 ( .B1(n7970), .B2(n9059), .A(n7822), .ZN(n7823) );
  OAI21_X1 U9245 ( .B1(n7824), .B2(n9061), .A(n7823), .ZN(P2_U3161) );
  OAI21_X1 U9246 ( .B1(n7826), .B2(n8794), .A(n7825), .ZN(n7872) );
  INV_X1 U9247 ( .A(n7872), .ZN(n7839) );
  INV_X1 U9248 ( .A(n7920), .ZN(n7827) );
  AOI211_X1 U9249 ( .C1(n8175), .C2(n7828), .A(n11049), .B(n7827), .ZN(n7871)
         );
  INV_X1 U9250 ( .A(n8175), .ZN(n7829) );
  NOR2_X1 U9251 ( .A1(n7829), .A2(n10525), .ZN(n7832) );
  OAI22_X1 U9252 ( .A1(n11015), .A2(n7830), .B1(n8171), .B2(n11012), .ZN(n7831) );
  AOI211_X1 U9253 ( .C1(n7871), .C2(n10520), .A(n7832), .B(n7831), .ZN(n7838)
         );
  INV_X1 U9254 ( .A(n7833), .ZN(n7835) );
  INV_X1 U9255 ( .A(n7834), .ZN(n7914) );
  AOI21_X1 U9256 ( .B1(n7835), .B2(n8794), .A(n7914), .ZN(n7836) );
  OAI222_X1 U9257 ( .A1(n8944), .A2(n8172), .B1(n8353), .B2(n7863), .C1(n10929), .C2(n7836), .ZN(n7870) );
  NAND2_X1 U9258 ( .A1(n7870), .A2(n11015), .ZN(n7837) );
  OAI211_X1 U9259 ( .C1(n7839), .C2(n10504), .A(n7838), .B(n7837), .ZN(
        P1_U3283) );
  NAND2_X1 U9260 ( .A1(n7841), .A2(n7840), .ZN(n7842) );
  XNOR2_X1 U9261 ( .A(n7842), .B(n7847), .ZN(n7843) );
  NAND2_X1 U9262 ( .A1(n7843), .A2(n10512), .ZN(n7845) );
  NAND2_X1 U9263 ( .A1(n10207), .A2(n10507), .ZN(n7844) );
  NAND2_X1 U9264 ( .A1(n7845), .A2(n7844), .ZN(n11066) );
  INV_X1 U9265 ( .A(n11066), .ZN(n7856) );
  OAI21_X1 U9266 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(n11068) );
  XNOR2_X1 U9267 ( .A(n7849), .B(n7946), .ZN(n7851) );
  AND2_X1 U9268 ( .A1(n7916), .A2(n10509), .ZN(n7850) );
  AOI21_X1 U9269 ( .B1(n7851), .B2(n10599), .A(n7850), .ZN(n11064) );
  OAI22_X1 U9270 ( .A1(n11015), .A2(n5902), .B1(n7940), .B2(n11012), .ZN(n7852) );
  AOI21_X1 U9271 ( .B1(n11018), .B2(n7946), .A(n7852), .ZN(n7853) );
  OAI21_X1 U9272 ( .B1(n11064), .B2(n11021), .A(n7853), .ZN(n7854) );
  AOI21_X1 U9273 ( .B1(n11068), .B2(n11023), .A(n7854), .ZN(n7855) );
  OAI21_X1 U9274 ( .B1(n10529), .B2(n7856), .A(n7855), .ZN(P1_U3284) );
  NAND2_X1 U9275 ( .A1(n9336), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7857) );
  OAI21_X1 U9276 ( .B1(n9106), .B2(n9336), .A(n7857), .ZN(P2_U3521) );
  NAND2_X1 U9277 ( .A1(n7859), .A2(n7858), .ZN(n7860) );
  XOR2_X1 U9278 ( .A(n7861), .B(n7860), .Z(n7869) );
  NAND2_X1 U9279 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10770) );
  INV_X1 U9280 ( .A(n10770), .ZN(n7865) );
  OAI22_X1 U9281 ( .A1(n10194), .A2(n7863), .B1(n11101), .B2(n7862), .ZN(n7864) );
  AOI211_X1 U9282 ( .C1(n10189), .C2(n10208), .A(n7865), .B(n7864), .ZN(n7868)
         );
  NAND2_X1 U9283 ( .A1(n11088), .A2(n7866), .ZN(n7867) );
  OAI211_X1 U9284 ( .C1(n7869), .C2(n10199), .A(n7868), .B(n7867), .ZN(
        P1_U3221) );
  AOI211_X1 U9285 ( .C1(n11113), .C2(n7872), .A(n7871), .B(n7870), .ZN(n7876)
         );
  NOR2_X1 U9286 ( .A1(n11120), .A2(n5916), .ZN(n7873) );
  AOI21_X1 U9287 ( .B1(n8175), .B2(n8213), .A(n7873), .ZN(n7874) );
  OAI21_X1 U9288 ( .B1(n7876), .B2(n11117), .A(n7874), .ZN(P1_U3483) );
  AOI22_X1 U9289 ( .A1(n8175), .A2(n8211), .B1(n11115), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7875) );
  OAI21_X1 U9290 ( .B1(n7876), .B2(n11115), .A(n7875), .ZN(P1_U3532) );
  NAND2_X1 U9291 ( .A1(n9146), .A2(n9140), .ZN(n9137) );
  XNOR2_X1 U9292 ( .A(n7877), .B(n9137), .ZN(n10989) );
  INV_X1 U9293 ( .A(n9137), .ZN(n9273) );
  XNOR2_X1 U9294 ( .A(n7878), .B(n9273), .ZN(n7879) );
  OAI222_X1 U9295 ( .A1(n8523), .A2(n7881), .B1(n8524), .B2(n7880), .C1(n10967), .C2(n7879), .ZN(n10991) );
  NAND2_X1 U9296 ( .A1(n10991), .A2(n11048), .ZN(n7885) );
  OAI22_X1 U9297 ( .A1(n9984), .A2(n10988), .B1(n7882), .B2(n10950), .ZN(n7883) );
  AOI21_X1 U9298 ( .B1(n10981), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7883), .ZN(
        n7884) );
  OAI211_X1 U9299 ( .C1(n10989), .C2(n9954), .A(n7885), .B(n7884), .ZN(
        P2_U3229) );
  NAND2_X1 U9300 ( .A1(n7886), .A2(P1_U3973), .ZN(n7887) );
  OAI21_X1 U9301 ( .B1(n6742), .B2(P1_U3973), .A(n7887), .ZN(P1_U3583) );
  AND2_X1 U9302 ( .A1(n7888), .A2(n7896), .ZN(n7889) );
  XNOR2_X1 U9303 ( .A(n8048), .B(n7550), .ZN(n8128) );
  XNOR2_X1 U9304 ( .A(n8128), .B(n5260), .ZN(n7892) );
  OAI211_X1 U9305 ( .C1(n7893), .C2(n7892), .A(n8131), .B(n9076), .ZN(n7899)
         );
  INV_X1 U9306 ( .A(n7894), .ZN(n8044) );
  NOR2_X1 U9307 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9744), .ZN(n8109) );
  AOI21_X1 U9308 ( .B1(n9080), .B2(n9328), .A(n8109), .ZN(n7895) );
  OAI21_X1 U9309 ( .B1(n7896), .B2(n9067), .A(n7895), .ZN(n7897) );
  AOI21_X1 U9310 ( .B1(n9071), .B2(n8044), .A(n7897), .ZN(n7898) );
  OAI211_X1 U9311 ( .C1(n5261), .C2(n9088), .A(n7899), .B(n7898), .ZN(P2_U3171) );
  INV_X1 U9312 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7908) );
  INV_X1 U9313 ( .A(n7900), .ZN(n7901) );
  AOI21_X1 U9314 ( .B1(n9279), .B2(n7902), .A(n7901), .ZN(n11035) );
  AOI22_X1 U9315 ( .A1(n11035), .A2(n11132), .B1(n11151), .B2(n11044), .ZN(
        n7906) );
  XNOR2_X1 U9316 ( .A(n7903), .B(n9279), .ZN(n7905) );
  AOI21_X1 U9317 ( .B1(n7905), .B2(n10935), .A(n7904), .ZN(n11037) );
  NAND2_X1 U9318 ( .A1(n7906), .A2(n11037), .ZN(n7909) );
  NAND2_X1 U9319 ( .A1(n7909), .A2(n11157), .ZN(n7907) );
  OAI21_X1 U9320 ( .B1(n7908), .B2(n11157), .A(n7907), .ZN(P2_U3411) );
  NAND2_X1 U9321 ( .A1(n7909), .A2(n11153), .ZN(n7910) );
  OAI21_X1 U9322 ( .B1(n11153), .B2(n6475), .A(n7910), .ZN(P2_U3466) );
  INV_X1 U9323 ( .A(n7911), .ZN(n7913) );
  OAI222_X1 U9324 ( .A1(n8985), .A2(n7912), .B1(n8998), .B2(n7913), .C1(n9409), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U9325 ( .A1(n10659), .A2(n9573), .B1(n7742), .B2(n7913), .C1(
        P1_U3086), .C2(n8259), .ZN(P1_U3336) );
  INV_X1 U9326 ( .A(n8698), .ZN(n8702) );
  NAND2_X1 U9327 ( .A1(n8707), .A2(n8708), .ZN(n8796) );
  OAI21_X1 U9328 ( .B1(n7914), .B2(n8702), .A(n8796), .ZN(n7915) );
  OAI211_X1 U9329 ( .C1(n5240), .C2(n7950), .A(n7915), .B(n10512), .ZN(n7918)
         );
  AOI22_X1 U9330 ( .A1(n10507), .A2(n7916), .B1(n11090), .B2(n10509), .ZN(
        n7917) );
  NAND2_X1 U9331 ( .A1(n7918), .A2(n7917), .ZN(n7927) );
  INV_X1 U9332 ( .A(n7927), .ZN(n7926) );
  XNOR2_X1 U9333 ( .A(n7919), .B(n8796), .ZN(n7929) );
  NAND2_X1 U9334 ( .A1(n7929), .A2(n11023), .ZN(n7925) );
  AOI211_X1 U9335 ( .C1(n11089), .C2(n7920), .A(n11049), .B(n7954), .ZN(n7928)
         );
  NOR2_X1 U9336 ( .A1(n5330), .A2(n10525), .ZN(n7923) );
  OAI22_X1 U9337 ( .A1(n11015), .A2(n7921), .B1(n11100), .B2(n11012), .ZN(
        n7922) );
  AOI211_X1 U9338 ( .C1(n7928), .C2(n10520), .A(n7923), .B(n7922), .ZN(n7924)
         );
  OAI211_X1 U9339 ( .C1(n10529), .C2(n7926), .A(n7925), .B(n7924), .ZN(
        P1_U3282) );
  AOI211_X1 U9340 ( .C1(n7929), .C2(n11113), .A(n7928), .B(n7927), .ZN(n7934)
         );
  AOI22_X1 U9341 ( .A1(n11089), .A2(n8211), .B1(n11115), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7930) );
  OAI21_X1 U9342 ( .B1(n7934), .B2(n11115), .A(n7930), .ZN(P1_U3533) );
  INV_X1 U9343 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7931) );
  NOR2_X1 U9344 ( .A1(n11120), .A2(n7931), .ZN(n7932) );
  AOI21_X1 U9345 ( .B1(n11089), .B2(n8213), .A(n7932), .ZN(n7933) );
  OAI21_X1 U9346 ( .B1(n7934), .B2(n11117), .A(n7933), .ZN(P1_U3486) );
  INV_X1 U9347 ( .A(n7936), .ZN(n7937) );
  AOI21_X1 U9348 ( .B1(n7939), .B2(n7938), .A(n7937), .ZN(n7948) );
  INV_X1 U9349 ( .A(n7940), .ZN(n7941) );
  AOI22_X1 U9350 ( .A1(n7941), .A2(n10190), .B1(n10189), .B2(n10207), .ZN(
        n7944) );
  INV_X1 U9351 ( .A(n7942), .ZN(n7943) );
  OAI211_X1 U9352 ( .C1(n11095), .C2(n10194), .A(n7944), .B(n7943), .ZN(n7945)
         );
  AOI21_X1 U9353 ( .B1(n7946), .B2(n11088), .A(n7945), .ZN(n7947) );
  OAI21_X1 U9354 ( .B1(n7948), .B2(n10199), .A(n7947), .ZN(P1_U3231) );
  XNOR2_X1 U9355 ( .A(n7949), .B(n8797), .ZN(n11114) );
  INV_X1 U9356 ( .A(n11114), .ZN(n7960) );
  NAND3_X1 U9357 ( .A1(n7950), .A2(n8707), .A3(n8797), .ZN(n7951) );
  NAND3_X1 U9358 ( .A1(n8138), .A2(n10512), .A3(n7951), .ZN(n7953) );
  AOI22_X1 U9359 ( .A1(n10509), .A2(n10204), .B1(n10205), .B2(n10507), .ZN(
        n7952) );
  NAND2_X1 U9360 ( .A1(n7953), .A2(n7952), .ZN(n11112) );
  OAI211_X1 U9361 ( .C1(n11110), .C2(n7954), .A(n10599), .B(n8147), .ZN(n11108) );
  OAI22_X1 U9362 ( .A1(n11015), .A2(n5955), .B1(n8274), .B2(n11012), .ZN(n7955) );
  AOI21_X1 U9363 ( .B1(n7956), .B2(n11018), .A(n7955), .ZN(n7957) );
  OAI21_X1 U9364 ( .B1(n11108), .B2(n11021), .A(n7957), .ZN(n7958) );
  AOI21_X1 U9365 ( .B1(n11112), .B2(n11015), .A(n7958), .ZN(n7959) );
  OAI21_X1 U9366 ( .B1(n7960), .B2(n10504), .A(n7959), .ZN(P1_U3281) );
  NAND2_X1 U9367 ( .A1(n7900), .A2(n7961), .ZN(n7962) );
  INV_X1 U9368 ( .A(n7965), .ZN(n9282) );
  XNOR2_X1 U9369 ( .A(n7962), .B(n9282), .ZN(n11057) );
  NAND2_X1 U9370 ( .A1(n7964), .A2(n7963), .ZN(n7966) );
  XNOR2_X1 U9371 ( .A(n7966), .B(n7965), .ZN(n7967) );
  AOI222_X1 U9372 ( .A1(n10935), .A2(n7967), .B1(n5260), .B2(n10944), .C1(
        n9330), .C2(n9961), .ZN(n11058) );
  MUX2_X1 U9373 ( .A(n7968), .B(n11058), .S(n11048), .Z(n7972) );
  AOI22_X1 U9374 ( .A1(n11043), .A2(n7970), .B1(n11041), .B2(n7969), .ZN(n7971) );
  OAI211_X1 U9375 ( .C1(n11057), .C2(n9954), .A(n7972), .B(n7971), .ZN(
        P2_U3225) );
  NAND2_X1 U9376 ( .A1(n7973), .A2(n9133), .ZN(n7974) );
  XNOR2_X1 U9377 ( .A(n9275), .B(n7974), .ZN(n10985) );
  OAI22_X1 U9378 ( .A1(n9984), .A2(n10982), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10950), .ZN(n7981) );
  XNOR2_X1 U9379 ( .A(n7976), .B(n7975), .ZN(n7977) );
  NAND2_X1 U9380 ( .A1(n7977), .A2(n10935), .ZN(n7979) );
  AOI22_X1 U9381 ( .A1(n9961), .A2(n9335), .B1(n9333), .B2(n10944), .ZN(n7978)
         );
  NAND2_X1 U9382 ( .A1(n7979), .A2(n7978), .ZN(n10983) );
  MUX2_X1 U9383 ( .A(n10983), .B(P2_REG2_REG_3__SCAN_IN), .S(n10981), .Z(n7980) );
  AOI211_X1 U9384 ( .C1(n9987), .C2(n10985), .A(n7981), .B(n7980), .ZN(n7982)
         );
  INV_X1 U9385 ( .A(n7982), .ZN(P2_U3230) );
  NAND2_X1 U9386 ( .A1(n8013), .A2(n10663), .ZN(n7984) );
  OAI211_X1 U9387 ( .C1(n9788), .C2(n10659), .A(n7984), .B(n7983), .ZN(
        P1_U3335) );
  NOR2_X1 U9388 ( .A1(n8001), .A2(n7985), .ZN(n7987) );
  NAND2_X1 U9389 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n8103), .ZN(n7988) );
  OAI21_X1 U9390 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n8103), .A(n7988), .ZN(
        n7989) );
  AOI21_X1 U9391 ( .B1(n5192), .B2(n7989), .A(n8094), .ZN(n8012) );
  INV_X1 U9392 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7999) );
  MUX2_X1 U9393 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n9412), .Z(n8104) );
  XNOR2_X1 U9394 ( .A(n8104), .B(n8010), .ZN(n7995) );
  OR2_X1 U9395 ( .A1(n7991), .A2(n7990), .ZN(n7993) );
  NAND2_X1 U9396 ( .A1(n7993), .A2(n7992), .ZN(n7994) );
  NAND2_X1 U9397 ( .A1(n7995), .A2(n7994), .ZN(n8105) );
  OAI21_X1 U9398 ( .B1(n7995), .B2(n7994), .A(n8105), .ZN(n7997) );
  AOI21_X1 U9399 ( .B1(n7997), .B2(n10923), .A(n7996), .ZN(n7998) );
  OAI21_X1 U9400 ( .B1(n9422), .B2(n7999), .A(n7998), .ZN(n8009) );
  NOR2_X1 U9401 ( .A1(n8001), .A2(n8000), .ZN(n8003) );
  NAND2_X1 U9402 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n8103), .ZN(n8004) );
  OAI21_X1 U9403 ( .B1(n8103), .B2(P2_REG1_REG_8__SCAN_IN), .A(n8004), .ZN(
        n8005) );
  NOR2_X1 U9404 ( .A1(n8006), .A2(n8005), .ZN(n8097) );
  AOI21_X1 U9405 ( .B1(n8006), .B2(n8005), .A(n8097), .ZN(n8007) );
  NOR2_X1 U9406 ( .A1(n8007), .A2(n10915), .ZN(n8008) );
  AOI211_X1 U9407 ( .C1(n10906), .C2(n8010), .A(n8009), .B(n8008), .ZN(n8011)
         );
  OAI21_X1 U9408 ( .B1(n8012), .B2(n10918), .A(n8011), .ZN(P2_U3190) );
  INV_X1 U9409 ( .A(n8013), .ZN(n8015) );
  OAI222_X1 U9410 ( .A1(P2_U3151), .A2(n9268), .B1(n8998), .B2(n8015), .C1(
        n8014), .C2(n8985), .ZN(P2_U3275) );
  XNOR2_X1 U9411 ( .A(n10842), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10835) );
  OAI21_X1 U9412 ( .B1(n8026), .B2(P1_REG1_REG_12__SCAN_IN), .A(n8016), .ZN(
        n10836) );
  NOR2_X1 U9413 ( .A1(n10835), .A2(n10836), .ZN(n10834) );
  AOI21_X1 U9414 ( .B1(n10842), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10834), .ZN(
        n10796) );
  XNOR2_X1 U9415 ( .A(n10789), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10797) );
  NOR2_X1 U9416 ( .A1(n10796), .A2(n10797), .ZN(n10795) );
  AOI21_X1 U9417 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n10789), .A(n10795), .ZN(
        n8017) );
  NOR2_X1 U9418 ( .A1(n8017), .A2(n8029), .ZN(n8018) );
  XNOR2_X1 U9419 ( .A(n8029), .B(n8017), .ZN(n10808) );
  NOR2_X1 U9420 ( .A1(n10807), .A2(n10808), .ZN(n10806) );
  NOR2_X1 U9421 ( .A1(n8018), .A2(n10806), .ZN(n8021) );
  AOI22_X1 U9422 ( .A1(n8120), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8019), .B2(
        n8024), .ZN(n8020) );
  NAND2_X1 U9423 ( .A1(n8020), .A2(n8021), .ZN(n8119) );
  OAI21_X1 U9424 ( .B1(n8021), .B2(n8020), .A(n8119), .ZN(n8037) );
  NOR2_X1 U9425 ( .A1(n8022), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10103) );
  AOI21_X1 U9426 ( .B1(n10754), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10103), .ZN(
        n8023) );
  OAI21_X1 U9427 ( .B1(n10829), .B2(n8024), .A(n8023), .ZN(n8036) );
  OAI21_X1 U9428 ( .B1(n8026), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8025), .ZN(
        n10839) );
  NAND2_X1 U9429 ( .A1(n10842), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8027) );
  OAI21_X1 U9430 ( .B1(n10842), .B2(P1_REG2_REG_13__SCAN_IN), .A(n8027), .ZN(
        n10838) );
  NOR2_X1 U9431 ( .A1(n10839), .A2(n10838), .ZN(n10837) );
  AOI21_X1 U9432 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10842), .A(n10837), .ZN(
        n10791) );
  NAND2_X1 U9433 ( .A1(n10789), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8028) );
  OAI21_X1 U9434 ( .B1(n10789), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8028), .ZN(
        n10792) );
  NOR2_X1 U9435 ( .A1(n10791), .A2(n10792), .ZN(n10790) );
  AOI21_X1 U9436 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n10789), .A(n10790), .ZN(
        n8030) );
  NOR2_X1 U9437 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  INV_X1 U9438 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10810) );
  XNOR2_X1 U9439 ( .A(n8030), .B(n8029), .ZN(n10811) );
  NOR2_X1 U9440 ( .A1(n10810), .A2(n10811), .ZN(n10809) );
  NOR2_X1 U9441 ( .A1(n8031), .A2(n10809), .ZN(n8034) );
  NAND2_X1 U9442 ( .A1(n8120), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8032) );
  OAI21_X1 U9443 ( .B1(n8120), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8032), .ZN(
        n8033) );
  NOR2_X1 U9444 ( .A1(n8034), .A2(n8033), .ZN(n8118) );
  AOI211_X1 U9445 ( .C1(n8034), .C2(n8033), .A(n8118), .B(n10851), .ZN(n8035)
         );
  AOI211_X1 U9446 ( .C1(n10822), .C2(n8037), .A(n8036), .B(n8035), .ZN(n8038)
         );
  INV_X1 U9447 ( .A(n8038), .ZN(P1_U3259) );
  INV_X1 U9448 ( .A(n8039), .ZN(n8040) );
  AOI21_X1 U9449 ( .B1(n9281), .B2(n8041), .A(n8040), .ZN(n8049) );
  INV_X1 U9450 ( .A(n8049), .ZN(n8047) );
  XNOR2_X1 U9451 ( .A(n8042), .B(n9281), .ZN(n8043) );
  AOI222_X1 U9452 ( .A1(n10935), .A2(n8043), .B1(n9329), .B2(n9961), .C1(n9328), .C2(n10944), .ZN(n8050) );
  MUX2_X1 U9453 ( .A(n8101), .B(n8050), .S(n11048), .Z(n8046) );
  AOI22_X1 U9454 ( .A1(n11043), .A2(n8048), .B1(n11041), .B2(n8044), .ZN(n8045) );
  OAI211_X1 U9455 ( .C1(n9954), .C2(n8047), .A(n8046), .B(n8045), .ZN(P2_U3224) );
  INV_X1 U9456 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8053) );
  AOI22_X1 U9457 ( .A1(n8049), .A2(n11132), .B1(n11151), .B2(n8048), .ZN(n8051) );
  NAND2_X1 U9458 ( .A1(n8051), .A2(n8050), .ZN(n8054) );
  NAND2_X1 U9459 ( .A1(n8054), .A2(n11157), .ZN(n8052) );
  OAI21_X1 U9460 ( .B1(n8053), .B2(n11157), .A(n8052), .ZN(P2_U3417) );
  NAND2_X1 U9461 ( .A1(n8054), .A2(n11153), .ZN(n8055) );
  OAI21_X1 U9462 ( .B1(n11153), .B2(n8100), .A(n8055), .ZN(P2_U3468) );
  XNOR2_X1 U9463 ( .A(n8056), .B(n9285), .ZN(n8059) );
  NAND2_X1 U9464 ( .A1(n9326), .A2(n10944), .ZN(n8058) );
  NAND2_X1 U9465 ( .A1(n9328), .A2(n9961), .ZN(n8057) );
  NAND2_X1 U9466 ( .A1(n8058), .A2(n8057), .ZN(n8229) );
  AOI21_X1 U9467 ( .B1(n8059), .B2(n10935), .A(n8229), .ZN(n11081) );
  OAI22_X1 U9468 ( .A1(n11048), .A2(n6538), .B1(n8232), .B2(n10950), .ZN(n8060) );
  AOI21_X1 U9469 ( .B1(n11078), .B2(n11043), .A(n8060), .ZN(n8064) );
  NAND2_X1 U9470 ( .A1(n8061), .A2(n9166), .ZN(n8062) );
  XNOR2_X1 U9471 ( .A(n8062), .B(n9285), .ZN(n11079) );
  NAND2_X1 U9472 ( .A1(n11079), .A2(n9987), .ZN(n8063) );
  OAI211_X1 U9473 ( .C1(n11081), .C2(n10981), .A(n8064), .B(n8063), .ZN(
        P2_U3222) );
  OAI21_X1 U9474 ( .B1(n8067), .B2(n8066), .A(n8065), .ZN(n10956) );
  INV_X1 U9475 ( .A(n10956), .ZN(n8078) );
  OAI21_X1 U9476 ( .B1(n8069), .B2(n9270), .A(n8068), .ZN(n8071) );
  AOI21_X1 U9477 ( .B1(n8071), .B2(n10935), .A(n8070), .ZN(n10957) );
  INV_X1 U9478 ( .A(n10957), .ZN(n8076) );
  NOR2_X1 U9479 ( .A1(n11046), .A2(n7324), .ZN(n8075) );
  OAI22_X1 U9480 ( .A1(n9984), .A2(n8073), .B1(n8072), .B2(n10950), .ZN(n8074)
         );
  AOI211_X1 U9481 ( .C1(n8076), .C2(n11046), .A(n8075), .B(n8074), .ZN(n8077)
         );
  OAI21_X1 U9482 ( .B1(n8078), .B2(n9954), .A(n8077), .ZN(P2_U3232) );
  XNOR2_X1 U9483 ( .A(n8079), .B(n9277), .ZN(n8087) );
  OAI21_X1 U9484 ( .B1(n8082), .B2(n8081), .A(n8080), .ZN(n11007) );
  OAI22_X1 U9485 ( .A1(n8084), .A2(n8524), .B1(n8083), .B2(n8523), .ZN(n8085)
         );
  AOI21_X1 U9486 ( .B1(n11007), .B2(n8157), .A(n8085), .ZN(n8086) );
  OAI21_X1 U9487 ( .B1(n10967), .B2(n8087), .A(n8086), .ZN(n11005) );
  INV_X1 U9488 ( .A(n11005), .ZN(n8093) );
  INV_X1 U9489 ( .A(n11048), .ZN(n9958) );
  AND2_X1 U9490 ( .A1(n11048), .A2(n8088), .ZN(n8994) );
  NOR2_X1 U9491 ( .A1(n11046), .A2(n6448), .ZN(n8091) );
  OAI22_X1 U9492 ( .A1(n9984), .A2(n11004), .B1(n8089), .B2(n10950), .ZN(n8090) );
  AOI211_X1 U9493 ( .C1(n11007), .C2(n8994), .A(n8091), .B(n8090), .ZN(n8092)
         );
  OAI21_X1 U9494 ( .B1(n8093), .B2(n9958), .A(n8092), .ZN(P2_U3228) );
  NOR2_X1 U9495 ( .A1(n8101), .A2(n8095), .ZN(n8184) );
  AOI21_X1 U9496 ( .B1(n8101), .B2(n8095), .A(n8184), .ZN(n8116) );
  INV_X1 U9497 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8113) );
  AND2_X1 U9498 ( .A1(n8098), .A2(n8100), .ZN(n8099) );
  OAI21_X1 U9499 ( .B1(n8189), .B2(n8099), .A(n9429), .ZN(n8112) );
  MUX2_X1 U9500 ( .A(n8101), .B(n8100), .S(n9412), .Z(n8194) );
  XNOR2_X1 U9501 ( .A(n8194), .B(n8102), .ZN(n8108) );
  OR2_X1 U9502 ( .A1(n8104), .A2(n8103), .ZN(n8106) );
  NAND2_X1 U9503 ( .A1(n8106), .A2(n8105), .ZN(n8107) );
  OAI21_X1 U9504 ( .B1(n8108), .B2(n8107), .A(n8195), .ZN(n8110) );
  AOI21_X1 U9505 ( .B1(n8110), .B2(n10923), .A(n8109), .ZN(n8111) );
  OAI211_X1 U9506 ( .C1(n8113), .C2(n9422), .A(n8112), .B(n8111), .ZN(n8114)
         );
  AOI21_X1 U9507 ( .B1(n8193), .B2(n10906), .A(n8114), .ZN(n8115) );
  OAI21_X1 U9508 ( .B1(n8116), .B2(n10918), .A(n8115), .ZN(P2_U3191) );
  XNOR2_X1 U9509 ( .A(n8249), .B(n8117), .ZN(n8242) );
  AOI21_X1 U9510 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n8120), .A(n8118), .ZN(
        n8243) );
  XOR2_X1 U9511 ( .A(n8242), .B(n8243), .Z(n8127) );
  OAI21_X1 U9512 ( .B1(n8120), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8119), .ZN(
        n8252) );
  INV_X1 U9513 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8121) );
  XNOR2_X1 U9514 ( .A(n8249), .B(n8121), .ZN(n8251) );
  XNOR2_X1 U9515 ( .A(n8252), .B(n8251), .ZN(n8125) );
  NAND2_X1 U9516 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10114) );
  NAND2_X1 U9517 ( .A1(n10754), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n8122) );
  OAI211_X1 U9518 ( .C1(n10829), .C2(n8123), .A(n10114), .B(n8122), .ZN(n8124)
         );
  AOI21_X1 U9519 ( .B1(n8125), .B2(n10822), .A(n8124), .ZN(n8126) );
  OAI21_X1 U9520 ( .B1(n8127), .B2(n10851), .A(n8126), .ZN(P1_U3260) );
  INV_X1 U9521 ( .A(n8128), .ZN(n8129) );
  NAND2_X1 U9522 ( .A1(n8129), .A2(n5260), .ZN(n8130) );
  NAND2_X1 U9523 ( .A1(n8131), .A2(n8130), .ZN(n8226) );
  XOR2_X1 U9524 ( .A(n7550), .B(n11075), .Z(n8227) );
  XNOR2_X1 U9525 ( .A(n8228), .B(n8132), .ZN(n8137) );
  AOI22_X1 U9526 ( .A1(n9080), .A2(n9327), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3151), .ZN(n8134) );
  NAND2_X1 U9527 ( .A1(n9085), .A2(n5260), .ZN(n8133) );
  OAI211_X1 U9528 ( .C1(n9082), .C2(n8162), .A(n8134), .B(n8133), .ZN(n8135)
         );
  AOI21_X1 U9529 ( .B1(n11075), .B2(n9059), .A(n8135), .ZN(n8136) );
  OAI21_X1 U9530 ( .B1(n8137), .B2(n9061), .A(n8136), .ZN(P2_U3157) );
  INV_X1 U9531 ( .A(n8799), .ZN(n8140) );
  NAND2_X1 U9532 ( .A1(n8138), .A2(n8713), .ZN(n8139) );
  NAND2_X1 U9533 ( .A1(n8140), .A2(n8139), .ZN(n8141) );
  NAND2_X1 U9534 ( .A1(n8141), .A2(n8351), .ZN(n8142) );
  NAND2_X1 U9535 ( .A1(n8142), .A2(n10512), .ZN(n8144) );
  AOI22_X1 U9536 ( .A1(n10509), .A2(n10203), .B1(n11090), .B2(n10507), .ZN(
        n8143) );
  NAND2_X1 U9537 ( .A1(n8144), .A2(n8143), .ZN(n8208) );
  INV_X1 U9538 ( .A(n8208), .ZN(n8153) );
  XNOR2_X1 U9539 ( .A(n8145), .B(n8799), .ZN(n8210) );
  NAND2_X1 U9540 ( .A1(n8210), .A2(n11023), .ZN(n8152) );
  INV_X1 U9541 ( .A(n8364), .ZN(n8146) );
  AOI211_X1 U9542 ( .C1(n8214), .C2(n8147), .A(n11049), .B(n8146), .ZN(n8209)
         );
  INV_X1 U9543 ( .A(n8214), .ZN(n8307) );
  NOR2_X1 U9544 ( .A1(n8307), .A2(n10525), .ZN(n8150) );
  OAI22_X1 U9545 ( .A1(n11015), .A2(n8148), .B1(n8302), .B2(n11012), .ZN(n8149) );
  AOI211_X1 U9546 ( .C1(n8209), .C2(n10520), .A(n8150), .B(n8149), .ZN(n8151)
         );
  OAI211_X1 U9547 ( .C1(n10529), .C2(n8153), .A(n8152), .B(n8151), .ZN(
        P1_U3280) );
  NAND2_X1 U9548 ( .A1(n8039), .A2(n9154), .ZN(n8155) );
  INV_X1 U9549 ( .A(n9283), .ZN(n8154) );
  XNOR2_X1 U9550 ( .A(n8155), .B(n8154), .ZN(n8158) );
  INV_X1 U9551 ( .A(n8158), .ZN(n11072) );
  INV_X1 U9552 ( .A(n8994), .ZN(n8166) );
  XNOR2_X1 U9553 ( .A(n8156), .B(n9283), .ZN(n8161) );
  NAND2_X1 U9554 ( .A1(n8158), .A2(n8157), .ZN(n8160) );
  AOI22_X1 U9555 ( .A1(n5260), .A2(n9961), .B1(n10944), .B2(n9327), .ZN(n8159)
         );
  OAI211_X1 U9556 ( .C1(n10967), .C2(n8161), .A(n8160), .B(n8159), .ZN(n11073)
         );
  NAND2_X1 U9557 ( .A1(n11073), .A2(n11046), .ZN(n8165) );
  OAI22_X1 U9558 ( .A1(n11048), .A2(n8421), .B1(n8162), .B2(n10950), .ZN(n8163) );
  AOI21_X1 U9559 ( .B1(n11043), .B2(n11075), .A(n8163), .ZN(n8164) );
  OAI211_X1 U9560 ( .C1(n11072), .C2(n8166), .A(n8165), .B(n8164), .ZN(
        P2_U3223) );
  NAND2_X1 U9561 ( .A1(n8167), .A2(n8168), .ZN(n8170) );
  XNOR2_X1 U9562 ( .A(n8170), .B(n8169), .ZN(n8178) );
  NAND2_X1 U9563 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10859) );
  INV_X1 U9564 ( .A(n10859), .ZN(n8174) );
  OAI22_X1 U9565 ( .A1(n10194), .A2(n8172), .B1(n11101), .B2(n8171), .ZN(n8173) );
  AOI211_X1 U9566 ( .C1(n10189), .C2(n10206), .A(n8174), .B(n8173), .ZN(n8177)
         );
  NAND2_X1 U9567 ( .A1(n8175), .A2(n11088), .ZN(n8176) );
  OAI211_X1 U9568 ( .C1(n8178), .C2(n10199), .A(n8177), .B(n8176), .ZN(
        P1_U3217) );
  INV_X1 U9569 ( .A(n8179), .ZN(n8182) );
  OAI222_X1 U9570 ( .A1(n10659), .A2(n8180), .B1(n7742), .B2(n8182), .C1(n8818), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI222_X1 U9571 ( .A1(P2_U3151), .A2(n9120), .B1(n8998), .B2(n8182), .C1(
        n8181), .C2(n8985), .ZN(P2_U3274) );
  NOR2_X1 U9572 ( .A1(n8193), .A2(n8183), .ZN(n8185) );
  AOI22_X1 U9573 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n8428), .B1(n8434), .B2(
        n8421), .ZN(n8186) );
  AOI21_X1 U9574 ( .B1(n8187), .B2(n8186), .A(n8423), .ZN(n8207) );
  NOR2_X1 U9575 ( .A1(n8193), .A2(n8188), .ZN(n8190) );
  MUX2_X1 U9576 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n8427), .S(n8428), .Z(n8191)
         );
  AOI21_X1 U9577 ( .B1(n5186), .B2(n8191), .A(n8426), .ZN(n8192) );
  NOR2_X1 U9578 ( .A1(n8192), .A2(n10915), .ZN(n8205) );
  INV_X1 U9579 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U9580 ( .A1(n8194), .A2(n8193), .ZN(n8196) );
  MUX2_X1 U9581 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n9412), .Z(n8435) );
  XNOR2_X1 U9582 ( .A(n8435), .B(n8428), .ZN(n8197) );
  NAND2_X1 U9583 ( .A1(n8197), .A2(n8198), .ZN(n8436) );
  OAI21_X1 U9584 ( .B1(n8198), .B2(n8197), .A(n8436), .ZN(n8201) );
  INV_X1 U9585 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8199) );
  OAI22_X1 U9586 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8199), .B1(n10904), .B2(
        n8434), .ZN(n8200) );
  AOI21_X1 U9587 ( .B1(n8201), .B2(n10923), .A(n8200), .ZN(n8202) );
  OAI21_X1 U9588 ( .B1(n9422), .B2(n8203), .A(n8202), .ZN(n8204) );
  NOR2_X1 U9589 ( .A1(n8205), .A2(n8204), .ZN(n8206) );
  OAI21_X1 U9590 ( .B1(n8207), .B2(n10918), .A(n8206), .ZN(P2_U3192) );
  AOI211_X1 U9591 ( .C1(n8210), .C2(n11113), .A(n8209), .B(n8208), .ZN(n8216)
         );
  AOI22_X1 U9592 ( .A1(n8214), .A2(n8211), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n11115), .ZN(n8212) );
  OAI21_X1 U9593 ( .B1(n8216), .B2(n11115), .A(n8212), .ZN(P1_U3535) );
  AOI22_X1 U9594 ( .A1(n8214), .A2(n8213), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n11117), .ZN(n8215) );
  OAI21_X1 U9595 ( .B1(n8216), .B2(n11117), .A(n8215), .ZN(P1_U3492) );
  INV_X1 U9596 ( .A(n8286), .ZN(n9194) );
  OR2_X1 U9597 ( .A1(n9194), .A2(n9119), .ZN(n9185) );
  XNOR2_X1 U9598 ( .A(n8217), .B(n9290), .ZN(n11102) );
  XNOR2_X1 U9599 ( .A(n8218), .B(n9290), .ZN(n8221) );
  OR2_X1 U9600 ( .A1(n8414), .A2(n8523), .ZN(n8220) );
  NAND2_X1 U9601 ( .A1(n9327), .A2(n9961), .ZN(n8219) );
  AND2_X1 U9602 ( .A1(n8220), .A2(n8219), .ZN(n8290) );
  OAI21_X1 U9603 ( .B1(n8221), .B2(n10967), .A(n8290), .ZN(n11103) );
  NAND2_X1 U9604 ( .A1(n11103), .A2(n11046), .ZN(n8225) );
  INV_X1 U9605 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8222) );
  OAI22_X1 U9606 ( .A1(n11048), .A2(n8222), .B1(n8291), .B2(n10950), .ZN(n8223) );
  AOI21_X1 U9607 ( .B1(n11105), .B2(n11043), .A(n8223), .ZN(n8224) );
  OAI211_X1 U9608 ( .C1(n11102), .C2(n9954), .A(n8225), .B(n8224), .ZN(
        P2_U3221) );
  XNOR2_X1 U9609 ( .A(n11078), .B(n7550), .ZN(n8280) );
  XNOR2_X1 U9610 ( .A(n8280), .B(n9327), .ZN(n8282) );
  XNOR2_X1 U9611 ( .A(n8283), .B(n8282), .ZN(n8234) );
  AOI22_X1 U9612 ( .A1(n8229), .A2(n8568), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3151), .ZN(n8231) );
  NAND2_X1 U9613 ( .A1(n11078), .A2(n9059), .ZN(n8230) );
  OAI211_X1 U9614 ( .C1(n9082), .C2(n8232), .A(n8231), .B(n8230), .ZN(n8233)
         );
  AOI21_X1 U9615 ( .B1(n8234), .B2(n9076), .A(n8233), .ZN(n8235) );
  INV_X1 U9616 ( .A(n8235), .ZN(P2_U3176) );
  INV_X1 U9617 ( .A(n8236), .ZN(n8239) );
  OAI222_X1 U9618 ( .A1(n8985), .A2(n8238), .B1(n8998), .B2(n8239), .C1(
        P2_U3151), .C2(n8237), .ZN(P2_U3273) );
  NOR2_X1 U9619 ( .A1(n8249), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8241) );
  AOI21_X1 U9620 ( .B1(n8243), .B2(n8242), .A(n8241), .ZN(n10819) );
  OR2_X1 U9621 ( .A1(n8253), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U9622 ( .A1(n8253), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8245) );
  AND2_X1 U9623 ( .A1(n8244), .A2(n8245), .ZN(n10818) );
  AND2_X1 U9624 ( .A1(n10819), .A2(n10818), .ZN(n10821) );
  INV_X1 U9625 ( .A(n8245), .ZN(n8246) );
  NOR2_X1 U9626 ( .A1(n10821), .A2(n8246), .ZN(n8248) );
  MUX2_X1 U9627 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n6095), .S(n8259), .Z(n8247)
         );
  XNOR2_X1 U9628 ( .A(n8248), .B(n8247), .ZN(n8263) );
  NOR2_X1 U9629 ( .A1(n8249), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8250) );
  AOI21_X1 U9630 ( .B1(n8252), .B2(n8251), .A(n8250), .ZN(n10825) );
  OR2_X1 U9631 ( .A1(n8253), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U9632 ( .A1(n8253), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8255) );
  AND2_X1 U9633 ( .A1(n8254), .A2(n8255), .ZN(n10824) );
  NAND2_X1 U9634 ( .A1(n10825), .A2(n10824), .ZN(n10823) );
  NAND2_X1 U9635 ( .A1(n10823), .A2(n8255), .ZN(n8257) );
  INV_X1 U9636 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10585) );
  XNOR2_X1 U9637 ( .A(n8259), .B(n10585), .ZN(n8256) );
  XNOR2_X1 U9638 ( .A(n8257), .B(n8256), .ZN(n8261) );
  NAND2_X1 U9639 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U9640 ( .A1(n10754), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n8258) );
  OAI211_X1 U9641 ( .C1(n10829), .C2(n8259), .A(n10071), .B(n8258), .ZN(n8260)
         );
  AOI21_X1 U9642 ( .B1(n8261), .B2(n10822), .A(n8260), .ZN(n8262) );
  OAI21_X1 U9643 ( .B1(n8263), .B2(n10851), .A(n8262), .ZN(P1_U3262) );
  NAND2_X1 U9644 ( .A1(n8265), .A2(n10663), .ZN(n8264) );
  OAI211_X1 U9645 ( .C1(n9782), .C2(n10659), .A(n8264), .B(n8861), .ZN(
        P1_U3332) );
  NAND2_X1 U9646 ( .A1(n8265), .A2(n10054), .ZN(n8267) );
  OR2_X1 U9647 ( .A1(n8266), .A2(P2_U3151), .ZN(n9316) );
  OAI211_X1 U9648 ( .C1(n8268), .C2(n8985), .A(n8267), .B(n9316), .ZN(P2_U3272) );
  INV_X1 U9649 ( .A(n8297), .ZN(n8273) );
  AOI21_X1 U9650 ( .B1(n8270), .B2(n11086), .A(n8271), .ZN(n8272) );
  OAI21_X1 U9651 ( .B1(n8273), .B2(n8272), .A(n11097), .ZN(n8278) );
  OAI22_X1 U9652 ( .A1(n10194), .A2(n8354), .B1(n11101), .B2(n8274), .ZN(n8275) );
  AOI211_X1 U9653 ( .C1(n10189), .C2(n10205), .A(n8276), .B(n8275), .ZN(n8277)
         );
  OAI211_X1 U9654 ( .C1(n11110), .C2(n10183), .A(n8278), .B(n8277), .ZN(
        P1_U3224) );
  INV_X1 U9655 ( .A(n8284), .ZN(n8285) );
  MUX2_X1 U9656 ( .A(n8286), .B(n8285), .S(n8959), .Z(n8340) );
  INV_X1 U9657 ( .A(n8340), .ZN(n8288) );
  XNOR2_X1 U9658 ( .A(n11105), .B(n7550), .ZN(n8287) );
  NOR2_X1 U9659 ( .A1(n8287), .A2(n8331), .ZN(n8343) );
  NOR2_X1 U9660 ( .A1(n8288), .A2(n8343), .ZN(n8289) );
  XNOR2_X1 U9661 ( .A(n8344), .B(n8289), .ZN(n8295) );
  NAND2_X1 U9662 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8442) );
  OAI21_X1 U9663 ( .B1(n8290), .B2(n9019), .A(n8442), .ZN(n8293) );
  NOR2_X1 U9664 ( .A1(n9082), .A2(n8291), .ZN(n8292) );
  AOI211_X1 U9665 ( .C1(n11105), .C2(n9059), .A(n8293), .B(n8292), .ZN(n8294)
         );
  OAI21_X1 U9666 ( .B1(n8295), .B2(n9061), .A(n8294), .ZN(P2_U3164) );
  AND2_X1 U9667 ( .A1(n8297), .A2(n8296), .ZN(n8300) );
  OAI211_X1 U9668 ( .C1(n8300), .C2(n8299), .A(n11097), .B(n8298), .ZN(n8306)
         );
  NOR2_X1 U9669 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8301), .ZN(n10843) );
  OAI22_X1 U9670 ( .A1(n10194), .A2(n8303), .B1(n11101), .B2(n8302), .ZN(n8304) );
  AOI211_X1 U9671 ( .C1(n10189), .C2(n11090), .A(n10843), .B(n8304), .ZN(n8305) );
  OAI211_X1 U9672 ( .C1(n8307), .C2(n10183), .A(n8306), .B(n8305), .ZN(
        P1_U3234) );
  AOI21_X1 U9673 ( .B1(n8344), .B2(n8340), .A(n8343), .ZN(n8311) );
  XNOR2_X1 U9674 ( .A(n11124), .B(n7550), .ZN(n8309) );
  INV_X1 U9675 ( .A(n8309), .ZN(n8308) );
  NAND2_X1 U9676 ( .A1(n8308), .A2(n9325), .ZN(n8345) );
  NAND2_X1 U9677 ( .A1(n8309), .A2(n8414), .ZN(n8339) );
  NAND2_X1 U9678 ( .A1(n8345), .A2(n8339), .ZN(n8310) );
  XNOR2_X1 U9679 ( .A(n8311), .B(n8310), .ZN(n8317) );
  INV_X1 U9680 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8312) );
  NOR2_X1 U9681 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8312), .ZN(n8514) );
  NOR2_X1 U9682 ( .A1(n9067), .A2(n8331), .ZN(n8313) );
  AOI211_X1 U9683 ( .C1(n9080), .C2(n9324), .A(n8514), .B(n8313), .ZN(n8314)
         );
  OAI21_X1 U9684 ( .B1(n8332), .B2(n9082), .A(n8314), .ZN(n8315) );
  AOI21_X1 U9685 ( .B1(n11124), .B2(n9059), .A(n8315), .ZN(n8316) );
  OAI21_X1 U9686 ( .B1(n8317), .B2(n9061), .A(n8316), .ZN(P2_U3174) );
  OR2_X1 U9687 ( .A1(n8318), .A2(n8802), .ZN(n8319) );
  NAND2_X1 U9688 ( .A1(n8320), .A2(n8319), .ZN(n10604) );
  XNOR2_X1 U9689 ( .A(n8321), .B(n8802), .ZN(n8322) );
  NAND2_X1 U9690 ( .A1(n8322), .A2(n10512), .ZN(n8324) );
  AOI22_X1 U9691 ( .A1(n10508), .A2(n10509), .B1(n10507), .B2(n10203), .ZN(
        n8323) );
  NAND2_X1 U9692 ( .A1(n8324), .A2(n8323), .ZN(n10608) );
  OAI211_X1 U9693 ( .C1(n10606), .C2(n8363), .A(n10599), .B(n8376), .ZN(n10605) );
  OAI22_X1 U9694 ( .A1(n11015), .A2(n10810), .B1(n10188), .B2(n11012), .ZN(
        n8325) );
  AOI21_X1 U9695 ( .B1(n10197), .B2(n11018), .A(n8325), .ZN(n8326) );
  OAI21_X1 U9696 ( .B1(n10605), .B2(n11021), .A(n8326), .ZN(n8327) );
  AOI21_X1 U9697 ( .B1(n10608), .B2(n11015), .A(n8327), .ZN(n8328) );
  OAI21_X1 U9698 ( .B1(n10604), .B2(n10504), .A(n8328), .ZN(P1_U3278) );
  XNOR2_X1 U9699 ( .A(n8329), .B(n8335), .ZN(n8330) );
  OAI222_X1 U9700 ( .A1(n8523), .A2(n8463), .B1(n8524), .B2(n8331), .C1(n8330), 
        .C2(n10967), .ZN(n11122) );
  INV_X1 U9701 ( .A(n11124), .ZN(n8333) );
  OAI22_X1 U9702 ( .A1(n8333), .A2(n10974), .B1(n8332), .B2(n10950), .ZN(n8334) );
  OAI21_X1 U9703 ( .B1(n11122), .B2(n8334), .A(n11046), .ZN(n8338) );
  XNOR2_X1 U9704 ( .A(n8336), .B(n6768), .ZN(n11121) );
  NAND2_X1 U9705 ( .A1(n11121), .A2(n9987), .ZN(n8337) );
  OAI211_X1 U9706 ( .C1(n8507), .C2(n11046), .A(n8338), .B(n8337), .ZN(
        P2_U3220) );
  XNOR2_X1 U9707 ( .A(n8415), .B(n7550), .ZN(n8468) );
  XNOR2_X1 U9708 ( .A(n8468), .B(n8463), .ZN(n8469) );
  INV_X1 U9709 ( .A(n8339), .ZN(n8341) );
  XOR2_X1 U9710 ( .A(n8469), .B(n8470), .Z(n8350) );
  AOI22_X1 U9711 ( .A1(n9080), .A2(n9323), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8347) );
  NAND2_X1 U9712 ( .A1(n9085), .A2(n9325), .ZN(n8346) );
  OAI211_X1 U9713 ( .C1(n9082), .C2(n8416), .A(n8347), .B(n8346), .ZN(n8348)
         );
  AOI21_X1 U9714 ( .B1(n8415), .B2(n9059), .A(n8348), .ZN(n8349) );
  OAI21_X1 U9715 ( .B1(n8350), .B2(n9061), .A(n8349), .ZN(P2_U3155) );
  NAND2_X1 U9716 ( .A1(n8351), .A2(n8715), .ZN(n8352) );
  XNOR2_X1 U9717 ( .A(n8352), .B(n8800), .ZN(n8362) );
  OAI22_X1 U9718 ( .A1(n8355), .A2(n8944), .B1(n8354), .B2(n8353), .ZN(n8361)
         );
  NAND2_X1 U9719 ( .A1(n8356), .A2(n8800), .ZN(n8357) );
  NAND2_X1 U9720 ( .A1(n8358), .A2(n8357), .ZN(n10615) );
  NOR2_X1 U9721 ( .A1(n10615), .A2(n8359), .ZN(n8360) );
  AOI211_X1 U9722 ( .C1(n8362), .C2(n10512), .A(n8361), .B(n8360), .ZN(n10614)
         );
  AOI211_X1 U9723 ( .C1(n10612), .C2(n8364), .A(n11049), .B(n8363), .ZN(n10611) );
  INV_X1 U9724 ( .A(n10612), .ZN(n8367) );
  INV_X1 U9725 ( .A(n8393), .ZN(n8365) );
  AOI22_X1 U9726 ( .A1(n10529), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8365), .B2(
        n10521), .ZN(n8366) );
  OAI21_X1 U9727 ( .B1(n8367), .B2(n10525), .A(n8366), .ZN(n8370) );
  NOR2_X1 U9728 ( .A1(n10615), .A2(n8368), .ZN(n8369) );
  AOI211_X1 U9729 ( .C1(n10611), .C2(n10520), .A(n8370), .B(n8369), .ZN(n8371)
         );
  OAI21_X1 U9730 ( .B1(n10614), .B2(n10466), .A(n8371), .ZN(P1_U3279) );
  INV_X1 U9731 ( .A(n8372), .ZN(n8987) );
  OAI222_X1 U9732 ( .A1(P1_U3086), .A2(n6340), .B1(n7742), .B2(n8987), .C1(
        n9569), .C2(n10659), .ZN(P1_U3331) );
  OAI21_X1 U9733 ( .B1(n8374), .B2(n8803), .A(n8373), .ZN(n10603) );
  INV_X1 U9734 ( .A(n10516), .ZN(n8375) );
  AOI21_X1 U9735 ( .B1(n10598), .B2(n8376), .A(n8375), .ZN(n10600) );
  INV_X1 U9736 ( .A(n10598), .ZN(n10106) );
  INV_X1 U9737 ( .A(n10101), .ZN(n8377) );
  AOI22_X1 U9738 ( .A1(n10529), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8377), .B2(
        n10521), .ZN(n8378) );
  OAI21_X1 U9739 ( .B1(n10106), .B2(n10525), .A(n8378), .ZN(n8384) );
  NAND2_X1 U9740 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  XNOR2_X1 U9741 ( .A(n8381), .B(n8803), .ZN(n8382) );
  AOI222_X1 U9742 ( .A1(n10512), .A2(n8382), .B1(n10492), .B2(n10509), .C1(
        n10202), .C2(n10507), .ZN(n10602) );
  NOR2_X1 U9743 ( .A1(n10602), .A2(n10466), .ZN(n8383) );
  AOI211_X1 U9744 ( .C1(n10600), .C2(n10454), .A(n8384), .B(n8383), .ZN(n8385)
         );
  OAI21_X1 U9745 ( .B1(n10504), .B2(n10603), .A(n8385), .ZN(P1_U3277) );
  NAND2_X1 U9746 ( .A1(n8387), .A2(n8386), .ZN(n8388) );
  XOR2_X1 U9747 ( .A(n8389), .B(n8388), .Z(n8396) );
  NAND2_X1 U9748 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10803) );
  INV_X1 U9749 ( .A(n10803), .ZN(n8390) );
  AOI21_X1 U9750 ( .B1(n11091), .B2(n10202), .A(n8390), .ZN(n8392) );
  NAND2_X1 U9751 ( .A1(n10189), .A2(n10204), .ZN(n8391) );
  OAI211_X1 U9752 ( .C1(n11101), .C2(n8393), .A(n8392), .B(n8391), .ZN(n8394)
         );
  AOI21_X1 U9753 ( .B1(n10612), .B2(n11088), .A(n8394), .ZN(n8395) );
  OAI21_X1 U9754 ( .B1(n8396), .B2(n10199), .A(n8395), .ZN(P1_U3215) );
  NAND2_X1 U9755 ( .A1(n8397), .A2(n8398), .ZN(n8399) );
  XNOR2_X1 U9756 ( .A(n8399), .B(n9191), .ZN(n11135) );
  NAND2_X1 U9757 ( .A1(n8410), .A2(n8400), .ZN(n8401) );
  INV_X1 U9758 ( .A(n9191), .ZN(n9291) );
  NAND2_X1 U9759 ( .A1(n8401), .A2(n9291), .ZN(n8403) );
  NAND3_X1 U9760 ( .A1(n8403), .A2(n10935), .A3(n8402), .ZN(n8406) );
  OAI22_X1 U9761 ( .A1(n8463), .A2(n8524), .B1(n8539), .B2(n8523), .ZN(n8404)
         );
  INV_X1 U9762 ( .A(n8404), .ZN(n8405) );
  NAND2_X1 U9763 ( .A1(n8406), .A2(n8405), .ZN(n11137) );
  NOR2_X1 U9764 ( .A1(n10950), .A2(n8466), .ZN(n8407) );
  OAI21_X1 U9765 ( .B1(n11137), .B2(n8407), .A(n11046), .ZN(n8409) );
  AOI22_X1 U9766 ( .A1(n11138), .A2(n11043), .B1(n10981), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n8408) );
  OAI211_X1 U9767 ( .C1(n9954), .C2(n11135), .A(n8409), .B(n8408), .ZN(
        P2_U3218) );
  INV_X1 U9768 ( .A(n8410), .ZN(n8411) );
  AOI21_X1 U9769 ( .B1(n9196), .B2(n8412), .A(n8411), .ZN(n8413) );
  OAI222_X1 U9770 ( .A1(n8523), .A2(n8467), .B1(n8524), .B2(n8414), .C1(n10967), .C2(n8413), .ZN(n11129) );
  INV_X1 U9771 ( .A(n8415), .ZN(n11128) );
  OAI22_X1 U9772 ( .A1(n11128), .A2(n10974), .B1(n8416), .B2(n10950), .ZN(
        n8417) );
  OAI21_X1 U9773 ( .B1(n11129), .B2(n8417), .A(n11046), .ZN(n8420) );
  OAI21_X1 U9774 ( .B1(n8418), .B2(n9196), .A(n8397), .ZN(n11131) );
  AOI22_X1 U9775 ( .A1(n11131), .A2(n9987), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n10981), .ZN(n8419) );
  NAND2_X1 U9776 ( .A1(n8420), .A2(n8419), .ZN(P2_U3219) );
  INV_X1 U9777 ( .A(n8501), .ZN(n8508) );
  NOR2_X1 U9778 ( .A1(n8428), .A2(n8421), .ZN(n8422) );
  NOR2_X1 U9779 ( .A1(n10917), .A2(n6538), .ZN(n10916) );
  MUX2_X1 U9780 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8222), .S(n8501), .Z(n8424)
         );
  NOR2_X1 U9781 ( .A1(n8424), .A2(n8425), .ZN(n8497) );
  AOI21_X1 U9782 ( .B1(n8425), .B2(n8424), .A(n8497), .ZN(n8447) );
  MUX2_X1 U9783 ( .A(n8500), .B(P2_REG1_REG_12__SCAN_IN), .S(n8501), .Z(n8432)
         );
  INV_X1 U9784 ( .A(n8426), .ZN(n8430) );
  OR2_X1 U9785 ( .A1(n8428), .A2(n8427), .ZN(n8429) );
  NAND2_X1 U9786 ( .A1(n8432), .A2(n8431), .ZN(n8503) );
  OAI21_X1 U9787 ( .B1(n8432), .B2(n8431), .A(n8503), .ZN(n8433) );
  NAND2_X1 U9788 ( .A1(n9429), .A2(n8433), .ZN(n8446) );
  MUX2_X1 U9789 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9412), .Z(n8439) );
  XNOR2_X1 U9790 ( .A(n8439), .B(n10905), .ZN(n10910) );
  OR2_X1 U9791 ( .A1(n8435), .A2(n8434), .ZN(n8437) );
  NAND2_X1 U9792 ( .A1(n8437), .A2(n8436), .ZN(n10909) );
  MUX2_X1 U9793 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n9412), .Z(n8509) );
  XNOR2_X1 U9794 ( .A(n8509), .B(n8501), .ZN(n8440) );
  NAND2_X1 U9795 ( .A1(n8440), .A2(n8441), .ZN(n8510) );
  OAI21_X1 U9796 ( .B1(n8441), .B2(n8440), .A(n8510), .ZN(n8444) );
  INV_X1 U9797 ( .A(n8442), .ZN(n8443) );
  AOI21_X1 U9798 ( .B1(n8444), .B2(n10923), .A(n8443), .ZN(n8445) );
  OAI211_X1 U9799 ( .C1(n8447), .C2(n10918), .A(n8446), .B(n8445), .ZN(n8448)
         );
  AOI21_X1 U9800 ( .B1(n10907), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8448), .ZN(
        n8449) );
  OAI21_X1 U9801 ( .B1(n8508), .B2(n10904), .A(n8449), .ZN(P2_U3194) );
  INV_X1 U9802 ( .A(n8450), .ZN(n8933) );
  OAI222_X1 U9803 ( .A1(P1_U3086), .A2(n8452), .B1(n7742), .B2(n8933), .C1(
        n8451), .C2(n10659), .ZN(P1_U3330) );
  XNOR2_X1 U9804 ( .A(n8453), .B(n9193), .ZN(n11141) );
  XNOR2_X1 U9805 ( .A(n8454), .B(n9292), .ZN(n8457) );
  OR2_X1 U9806 ( .A1(n8542), .A2(n8523), .ZN(n8456) );
  OR2_X1 U9807 ( .A1(n8467), .A2(n8524), .ZN(n8455) );
  AND2_X1 U9808 ( .A1(n8456), .A2(n8455), .ZN(n8556) );
  OAI21_X1 U9809 ( .B1(n8457), .B2(n10967), .A(n8556), .ZN(n11142) );
  NAND2_X1 U9810 ( .A1(n11142), .A2(n11046), .ZN(n8462) );
  INV_X1 U9811 ( .A(n8558), .ZN(n8458) );
  OAI22_X1 U9812 ( .A1(n11048), .A2(n8459), .B1(n8458), .B2(n10950), .ZN(n8460) );
  AOI21_X1 U9813 ( .B1(n11144), .B2(n11043), .A(n8460), .ZN(n8461) );
  OAI211_X1 U9814 ( .C1(n11141), .C2(n9954), .A(n8462), .B(n8461), .ZN(
        P2_U3217) );
  AND2_X1 U9815 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9365) );
  NOR2_X1 U9816 ( .A1(n9067), .A2(n8463), .ZN(n8464) );
  AOI211_X1 U9817 ( .C1(n9080), .C2(n9322), .A(n9365), .B(n8464), .ZN(n8465)
         );
  OAI21_X1 U9818 ( .B1(n8466), .B2(n9082), .A(n8465), .ZN(n8474) );
  XNOR2_X1 U9819 ( .A(n11138), .B(n7550), .ZN(n8536) );
  XNOR2_X1 U9820 ( .A(n8536), .B(n8467), .ZN(n8472) );
  NOR2_X1 U9821 ( .A1(n8471), .A2(n8472), .ZN(n8537) );
  AOI211_X1 U9822 ( .C1(n8472), .C2(n8471), .A(n9061), .B(n8537), .ZN(n8473)
         );
  AOI211_X1 U9823 ( .C1(n11138), .C2(n9059), .A(n8474), .B(n8473), .ZN(n8475)
         );
  INV_X1 U9824 ( .A(n8475), .ZN(P2_U3181) );
  INV_X1 U9825 ( .A(n8476), .ZN(n8480) );
  OAI222_X1 U9826 ( .A1(n8985), .A2(n8478), .B1(n8998), .B2(n8480), .C1(n8477), 
        .C2(P2_U3151), .ZN(P2_U3269) );
  OAI222_X1 U9827 ( .A1(n10659), .A2(n8481), .B1(n7742), .B2(n8480), .C1(
        P1_U3086), .C2(n8479), .ZN(P1_U3329) );
  INV_X1 U9828 ( .A(n8482), .ZN(n8646) );
  AOI21_X1 U9829 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n8534), .A(n8483), .ZN(
        n8484) );
  OAI21_X1 U9830 ( .B1(n8646), .B2(n8998), .A(n8484), .ZN(P2_U3268) );
  INV_X1 U9831 ( .A(n8487), .ZN(n9295) );
  XNOR2_X1 U9832 ( .A(n8485), .B(n9295), .ZN(n11147) );
  XNOR2_X1 U9833 ( .A(n8486), .B(n8487), .ZN(n8490) );
  OR2_X1 U9834 ( .A1(n8539), .A2(n8524), .ZN(n8489) );
  NAND2_X1 U9835 ( .A1(n9320), .A2(n10944), .ZN(n8488) );
  AND2_X1 U9836 ( .A1(n8489), .A2(n8488), .ZN(n8547) );
  OAI21_X1 U9837 ( .B1(n8490), .B2(n10967), .A(n8547), .ZN(n11148) );
  NAND2_X1 U9838 ( .A1(n11148), .A2(n11046), .ZN(n8495) );
  INV_X1 U9839 ( .A(n8546), .ZN(n8491) );
  NAND2_X1 U9840 ( .A1(n11041), .A2(n8491), .ZN(n8492) );
  OAI21_X1 U9841 ( .B1(n11048), .B2(n6615), .A(n8492), .ZN(n8493) );
  AOI21_X1 U9842 ( .B1(n11150), .B2(n11043), .A(n8493), .ZN(n8494) );
  OAI211_X1 U9843 ( .C1(n11147), .C2(n9954), .A(n8495), .B(n8494), .ZN(
        P2_U3216) );
  AOI21_X1 U9844 ( .B1(n8507), .B2(n8499), .A(n8577), .ZN(n8521) );
  INV_X1 U9845 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8518) );
  OR2_X1 U9846 ( .A1(n8501), .A2(n8500), .ZN(n8502) );
  AND2_X1 U9847 ( .A1(n8504), .A2(n8506), .ZN(n8505) );
  OAI21_X1 U9848 ( .B1(n8587), .B2(n8505), .A(n9429), .ZN(n8517) );
  MUX2_X1 U9849 ( .A(n8507), .B(n8506), .S(n9412), .Z(n8606) );
  XNOR2_X1 U9850 ( .A(n8606), .B(n8498), .ZN(n8513) );
  OR2_X1 U9851 ( .A1(n8509), .A2(n8508), .ZN(n8511) );
  NAND2_X1 U9852 ( .A1(n8511), .A2(n8510), .ZN(n8512) );
  NAND2_X1 U9853 ( .A1(n8513), .A2(n8512), .ZN(n8607) );
  OAI21_X1 U9854 ( .B1(n8513), .B2(n8512), .A(n8607), .ZN(n8515) );
  AOI21_X1 U9855 ( .B1(n8515), .B2(n10923), .A(n8514), .ZN(n8516) );
  OAI211_X1 U9856 ( .C1(n8518), .C2(n9422), .A(n8517), .B(n8516), .ZN(n8519)
         );
  AOI21_X1 U9857 ( .B1(n8605), .B2(n10906), .A(n8519), .ZN(n8520) );
  OAI21_X1 U9858 ( .B1(n8521), .B2(n10918), .A(n8520), .ZN(P2_U3195) );
  XNOR2_X1 U9859 ( .A(n8522), .B(n9296), .ZN(n8525) );
  OAI22_X1 U9860 ( .A1(n8542), .A2(n8524), .B1(n8954), .B2(n8523), .ZN(n8569)
         );
  AOI21_X1 U9861 ( .B1(n8525), .B2(n10935), .A(n8569), .ZN(n10034) );
  OAI22_X1 U9862 ( .A1(n11048), .A2(n8526), .B1(n8571), .B2(n10950), .ZN(n8527) );
  AOI21_X1 U9863 ( .B1(n10032), .B2(n11043), .A(n8527), .ZN(n8531) );
  OR2_X1 U9864 ( .A1(n8528), .A2(n9296), .ZN(n10033) );
  NAND3_X1 U9865 ( .A1(n10033), .A2(n9987), .A3(n8529), .ZN(n8530) );
  OAI211_X1 U9866 ( .C1(n10034), .C2(n10981), .A(n8531), .B(n8530), .ZN(
        P2_U3215) );
  INV_X1 U9867 ( .A(n8532), .ZN(n8562) );
  AOI21_X1 U9868 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n8534), .A(n8533), .ZN(
        n8535) );
  OAI21_X1 U9869 ( .B1(n8562), .B2(n8998), .A(n8535), .ZN(P2_U3267) );
  XNOR2_X1 U9870 ( .A(n11144), .B(n7550), .ZN(n8540) );
  INV_X1 U9871 ( .A(n8540), .ZN(n8541) );
  INV_X1 U9872 ( .A(n8536), .ZN(n8538) );
  AOI21_X1 U9873 ( .B1(n8538), .B2(n9323), .A(n8537), .ZN(n8553) );
  XNOR2_X1 U9874 ( .A(n8540), .B(n8539), .ZN(n8554) );
  XNOR2_X1 U9875 ( .A(n11150), .B(n7550), .ZN(n8543) );
  INV_X1 U9876 ( .A(n8543), .ZN(n8544) );
  NAND2_X1 U9877 ( .A1(n8544), .A2(n9321), .ZN(n8564) );
  NAND2_X1 U9878 ( .A1(n5189), .A2(n8564), .ZN(n8545) );
  XNOR2_X1 U9879 ( .A(n8565), .B(n8545), .ZN(n8551) );
  NOR2_X1 U9880 ( .A1(n9082), .A2(n8546), .ZN(n8549) );
  INV_X1 U9881 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9397) );
  OAI22_X1 U9882 ( .A1(n8547), .A2(n9019), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9397), .ZN(n8548) );
  AOI211_X1 U9883 ( .C1(n11150), .C2(n9059), .A(n8549), .B(n8548), .ZN(n8550)
         );
  OAI21_X1 U9884 ( .B1(n8551), .B2(n9061), .A(n8550), .ZN(P2_U3168) );
  INV_X1 U9885 ( .A(n11144), .ZN(n8561) );
  AOI211_X1 U9886 ( .C1(n8554), .C2(n8553), .A(n9061), .B(n8552), .ZN(n8555)
         );
  INV_X1 U9887 ( .A(n8555), .ZN(n8560) );
  OAI22_X1 U9888 ( .A1(n8556), .A2(n9019), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9381), .ZN(n8557) );
  AOI21_X1 U9889 ( .B1(n9071), .B2(n8558), .A(n8557), .ZN(n8559) );
  OAI211_X1 U9890 ( .C1(n8561), .C2(n9088), .A(n8560), .B(n8559), .ZN(P2_U3166) );
  OAI222_X1 U9891 ( .A1(n10659), .A2(n8563), .B1(n7742), .B2(n8562), .C1(n5123), .C2(P1_U3086), .ZN(P1_U3327) );
  XNOR2_X1 U9892 ( .A(n10032), .B(n7550), .ZN(n8951) );
  XNOR2_X1 U9893 ( .A(n8951), .B(n8950), .ZN(n8567) );
  AOI21_X1 U9894 ( .B1(n8567), .B2(n8566), .A(n8953), .ZN(n8574) );
  NAND2_X1 U9895 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n8629) );
  NAND2_X1 U9896 ( .A1(n8569), .A2(n8568), .ZN(n8570) );
  OAI211_X1 U9897 ( .C1(n9082), .C2(n8571), .A(n8629), .B(n8570), .ZN(n8572)
         );
  AOI21_X1 U9898 ( .B1(n10032), .B2(n9059), .A(n8572), .ZN(n8573) );
  OAI21_X1 U9899 ( .B1(n8574), .B2(n9061), .A(n8573), .ZN(P2_U3178) );
  NOR2_X1 U9900 ( .A1(n8605), .A2(n8576), .ZN(n8578) );
  NAND2_X1 U9901 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9347), .ZN(n8579) );
  OAI21_X1 U9902 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9347), .A(n8579), .ZN(
        n9339) );
  NOR2_X1 U9903 ( .A1(n9371), .A2(n8580), .ZN(n8581) );
  AOI22_X1 U9904 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8613), .B1(n9380), .B2(
        n8459), .ZN(n9377) );
  NOR2_X1 U9905 ( .A1(n9378), .A2(n9377), .ZN(n9376) );
  NOR2_X1 U9906 ( .A1(n8618), .A2(n8582), .ZN(n8583) );
  NAND2_X1 U9907 ( .A1(n9417), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9405) );
  OAI21_X1 U9908 ( .B1(n9417), .B2(P2_REG2_REG_18__SCAN_IN), .A(n9405), .ZN(
        n8584) );
  AOI21_X1 U9909 ( .B1(n8585), .B2(n8584), .A(n9406), .ZN(n8634) );
  NOR2_X1 U9910 ( .A1(n8605), .A2(n8586), .ZN(n8588) );
  NAND2_X1 U9911 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9347), .ZN(n8589) );
  OAI21_X1 U9912 ( .B1(n9347), .B2(P2_REG1_REG_14__SCAN_IN), .A(n8589), .ZN(
        n9342) );
  AOI21_X1 U9913 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9347), .A(n9341), .ZN(
        n8590) );
  NOR2_X1 U9914 ( .A1(n9371), .A2(n8590), .ZN(n8591) );
  MUX2_X1 U9915 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8592), .S(n8613), .Z(n9375)
         );
  NOR2_X1 U9916 ( .A1(n8618), .A2(n8593), .ZN(n8594) );
  INV_X1 U9917 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11152) );
  XNOR2_X1 U9918 ( .A(n8618), .B(n8593), .ZN(n9395) );
  MUX2_X1 U9919 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n5611), .S(n8595), .Z(n8596)
         );
  AOI21_X1 U9920 ( .B1(n8597), .B2(n8596), .A(n9408), .ZN(n8598) );
  INV_X1 U9921 ( .A(n8598), .ZN(n8632) );
  MUX2_X1 U9922 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9412), .Z(n8611) );
  XNOR2_X1 U9923 ( .A(n8613), .B(n8611), .ZN(n9382) );
  MUX2_X1 U9924 ( .A(n8600), .B(n8599), .S(n9412), .Z(n8602) );
  NAND2_X1 U9925 ( .A1(n8602), .A2(n9371), .ZN(n8610) );
  XNOR2_X1 U9926 ( .A(n8602), .B(n8601), .ZN(n9364) );
  MUX2_X1 U9927 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n9412), .Z(n8604) );
  OR2_X1 U9928 ( .A1(n8604), .A2(n9347), .ZN(n8609) );
  XNOR2_X1 U9929 ( .A(n8604), .B(n8603), .ZN(n9345) );
  NAND2_X1 U9930 ( .A1(n8606), .A2(n8605), .ZN(n8608) );
  NAND2_X1 U9931 ( .A1(n8608), .A2(n8607), .ZN(n9346) );
  NAND2_X1 U9932 ( .A1(n9345), .A2(n9346), .ZN(n9344) );
  NAND2_X1 U9933 ( .A1(n8609), .A2(n9344), .ZN(n9363) );
  NAND2_X1 U9934 ( .A1(n9382), .A2(n9383), .ZN(n8615) );
  INV_X1 U9935 ( .A(n8611), .ZN(n8612) );
  NAND2_X1 U9936 ( .A1(n8613), .A2(n8612), .ZN(n8614) );
  MUX2_X1 U9937 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n9412), .Z(n8616) );
  XNOR2_X1 U9938 ( .A(n8618), .B(n8616), .ZN(n9392) );
  INV_X1 U9939 ( .A(n8616), .ZN(n8617) );
  AND2_X1 U9940 ( .A1(n8618), .A2(n8617), .ZN(n8619) );
  AOI21_X1 U9941 ( .B1(n9393), .B2(n9392), .A(n8619), .ZN(n8620) );
  MUX2_X1 U9942 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6789), .Z(n8621) );
  AND2_X1 U9943 ( .A1(n8620), .A2(n8621), .ZN(n9415) );
  INV_X1 U9944 ( .A(n8620), .ZN(n8623) );
  INV_X1 U9945 ( .A(n8621), .ZN(n8622) );
  NAND2_X1 U9946 ( .A1(n8623), .A2(n8622), .ZN(n9416) );
  INV_X1 U9947 ( .A(n9416), .ZN(n8624) );
  NOR2_X1 U9948 ( .A1(n9415), .A2(n8624), .ZN(n8626) );
  INV_X1 U9949 ( .A(n8626), .ZN(n8625) );
  OAI21_X1 U9950 ( .B1(n8625), .B2(n9336), .A(n10904), .ZN(n8628) );
  NOR2_X1 U9951 ( .A1(n8626), .A2(n9426), .ZN(n8627) );
  INV_X1 U9952 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10741) );
  OAI21_X1 U9953 ( .B1(n9422), .B2(n10741), .A(n8629), .ZN(n8630) );
  OAI21_X1 U9954 ( .B1(n8634), .B2(n10918), .A(n8633), .ZN(P2_U3200) );
  INV_X1 U9955 ( .A(n8762), .ZN(n8949) );
  OAI222_X1 U9956 ( .A1(n8998), .A2(n8949), .B1(n8985), .B2(n6742), .C1(n8635), 
        .C2(P2_U3151), .ZN(P2_U3266) );
  INV_X1 U9957 ( .A(SI_29_), .ZN(n9661) );
  INV_X1 U9958 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9098) );
  INV_X1 U9959 ( .A(SI_30_), .ZN(n8641) );
  NAND2_X1 U9960 ( .A1(n8642), .A2(n8641), .ZN(n8654) );
  INV_X1 U9961 ( .A(n8642), .ZN(n8643) );
  NAND2_X1 U9962 ( .A1(n8643), .A2(SI_30_), .ZN(n8644) );
  NAND2_X1 U9963 ( .A1(n8654), .A2(n8644), .ZN(n8655) );
  INV_X1 U9964 ( .A(n9097), .ZN(n8997) );
  OAI222_X1 U9965 ( .A1(n10659), .A2(n9764), .B1(n7742), .B2(n8997), .C1(
        P1_U3086), .C2(n8645), .ZN(P1_U3325) );
  OAI222_X1 U9966 ( .A1(n10659), .A2(n9774), .B1(n7742), .B2(n8646), .C1(
        P1_U3086), .C2(n10748), .ZN(P1_U3328) );
  INV_X1 U9967 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U9968 ( .A1(n8647), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8651) );
  INV_X1 U9969 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8648) );
  OR2_X1 U9970 ( .A1(n8649), .A2(n8648), .ZN(n8650) );
  OAI211_X1 U9971 ( .C1(n8653), .C2(n8652), .A(n8651), .B(n8650), .ZN(n10201)
         );
  INV_X1 U9972 ( .A(SI_31_), .ZN(n9657) );
  XNOR2_X1 U9973 ( .A(n8657), .B(n9657), .ZN(n8658) );
  NAND2_X1 U9974 ( .A1(n10664), .A2(n5948), .ZN(n8661) );
  INV_X1 U9975 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10660) );
  OR2_X1 U9976 ( .A1(n8777), .A2(n10660), .ZN(n8660) );
  AND2_X1 U9977 ( .A1(n8663), .A2(n8662), .ZN(n8718) );
  INV_X1 U9978 ( .A(n8718), .ZN(n8888) );
  OAI211_X1 U9979 ( .C1(n8888), .C2(n8715), .A(n8724), .B(n8664), .ZN(n8890)
         );
  INV_X1 U9980 ( .A(n8878), .ZN(n8695) );
  NAND2_X1 U9981 ( .A1(n8665), .A2(n8871), .ZN(n8668) );
  NAND4_X1 U9982 ( .A1(n8668), .A2(n8667), .A3(n8666), .A4(n8867), .ZN(n8670)
         );
  MUX2_X1 U9983 ( .A(n8670), .B(n8669), .S(n8782), .Z(n8675) );
  NAND2_X1 U9984 ( .A1(n8672), .A2(n8671), .ZN(n8874) );
  NAND3_X1 U9985 ( .A1(n8874), .A2(n8815), .A3(n8873), .ZN(n8673) );
  NAND3_X1 U9986 ( .A1(n8675), .A2(n8674), .A3(n8673), .ZN(n8682) );
  INV_X1 U9987 ( .A(n8790), .ZN(n8678) );
  INV_X1 U9988 ( .A(n8676), .ZN(n8677) );
  MUX2_X1 U9989 ( .A(n8678), .B(n8677), .S(n8815), .Z(n8679) );
  NOR2_X1 U9990 ( .A1(n8680), .A2(n8679), .ZN(n8681) );
  NAND2_X1 U9991 ( .A1(n8682), .A2(n8681), .ZN(n8689) );
  INV_X1 U9992 ( .A(n8683), .ZN(n8684) );
  MUX2_X1 U9993 ( .A(n8685), .B(n8684), .S(n8782), .Z(n8686) );
  NOR2_X1 U9994 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  NAND2_X1 U9995 ( .A1(n8689), .A2(n8688), .ZN(n8693) );
  NAND2_X1 U9996 ( .A1(n8878), .A2(n8690), .ZN(n8691) );
  NAND2_X1 U9997 ( .A1(n8691), .A2(n8815), .ZN(n8692) );
  OAI211_X1 U9998 ( .C1(n8695), .C2(n8694), .A(n8697), .B(n8881), .ZN(n8696)
         );
  INV_X1 U9999 ( .A(n8697), .ZN(n8700) );
  NAND3_X1 U10000 ( .A1(n8700), .A2(n8699), .A3(n8698), .ZN(n8705) );
  OAI211_X1 U10001 ( .C1(n8702), .C2(n8701), .A(n8707), .B(n8878), .ZN(n8703)
         );
  NAND2_X1 U10002 ( .A1(n8713), .A2(n8707), .ZN(n8863) );
  NAND2_X1 U10003 ( .A1(n8883), .A2(n8708), .ZN(n8709) );
  MUX2_X1 U10004 ( .A(n8863), .B(n8709), .S(n8782), .Z(n8710) );
  INV_X1 U10005 ( .A(n8710), .ZN(n8711) );
  NAND2_X1 U10006 ( .A1(n8712), .A2(n8711), .ZN(n8716) );
  AND3_X1 U10007 ( .A1(n8718), .A2(n8713), .A3(n8716), .ZN(n8714) );
  NOR2_X1 U10008 ( .A1(n8890), .A2(n8714), .ZN(n8723) );
  NAND3_X1 U10009 ( .A1(n8716), .A2(n8883), .A3(n8715), .ZN(n8719) );
  AOI21_X1 U10010 ( .B1(n8719), .B2(n8718), .A(n8717), .ZN(n8721) );
  NOR2_X1 U10011 ( .A1(n8721), .A2(n8720), .ZN(n8722) );
  NAND2_X1 U10012 ( .A1(n8727), .A2(n8804), .ZN(n8731) );
  AOI21_X1 U10013 ( .B1(n8731), .B2(n8862), .A(n8728), .ZN(n8729) );
  OAI21_X1 U10014 ( .B1(n8729), .B2(n8815), .A(n8899), .ZN(n8737) );
  AND2_X1 U10015 ( .A1(n8740), .A2(n8730), .ZN(n8904) );
  NAND4_X1 U10016 ( .A1(n8731), .A2(n8815), .A3(n8895), .A4(n8894), .ZN(n8735)
         );
  INV_X1 U10017 ( .A(n8896), .ZN(n8732) );
  OAI21_X1 U10018 ( .B1(n8733), .B2(n8732), .A(n8815), .ZN(n8734) );
  NAND3_X1 U10019 ( .A1(n8735), .A2(n10438), .A3(n8734), .ZN(n8736) );
  AOI21_X1 U10020 ( .B1(n8737), .B2(n8904), .A(n8736), .ZN(n8739) );
  AOI21_X1 U10021 ( .B1(n10438), .B2(n8899), .A(n8782), .ZN(n8738) );
  NOR2_X1 U10022 ( .A1(n8740), .A2(n8782), .ZN(n8741) );
  NOR2_X1 U10023 ( .A1(n10444), .A2(n8741), .ZN(n8745) );
  MUX2_X1 U10024 ( .A(n8743), .B(n8742), .S(n8782), .Z(n8744) );
  NAND2_X1 U10025 ( .A1(n8750), .A2(n10410), .ZN(n8827) );
  NAND2_X1 U10026 ( .A1(n8828), .A2(n8747), .ZN(n8824) );
  MUX2_X1 U10027 ( .A(n8827), .B(n8824), .S(n8815), .Z(n8748) );
  INV_X1 U10028 ( .A(n8748), .ZN(n8749) );
  MUX2_X1 U10029 ( .A(n8828), .B(n8750), .S(n8815), .Z(n8751) );
  NAND2_X1 U10030 ( .A1(n8752), .A2(n8829), .ZN(n8753) );
  NAND2_X1 U10031 ( .A1(n8753), .A2(n8757), .ZN(n8756) );
  NAND3_X1 U10032 ( .A1(n10379), .A2(n8825), .A3(n8754), .ZN(n8755) );
  NAND2_X1 U10033 ( .A1(n8758), .A2(n8757), .ZN(n8909) );
  NAND2_X1 U10034 ( .A1(n8909), .A2(n8782), .ZN(n8759) );
  MUX2_X1 U10035 ( .A(n8782), .B(n8759), .S(n8832), .Z(n8760) );
  MUX2_X1 U10036 ( .A(n8821), .B(n8834), .S(n8815), .Z(n8761) );
  NOR2_X1 U10037 ( .A1(n8809), .A2(n8761), .ZN(n8771) );
  NAND2_X1 U10038 ( .A1(n8762), .A2(n5948), .ZN(n8764) );
  OR2_X1 U10039 ( .A1(n8777), .A2(n9760), .ZN(n8763) );
  NAND2_X1 U10040 ( .A1(n10538), .A2(n8765), .ZN(n8819) );
  NAND2_X1 U10041 ( .A1(n8772), .A2(n8819), .ZN(n8940) );
  MUX2_X1 U10042 ( .A(n8766), .B(n8939), .S(n8815), .Z(n8767) );
  INV_X1 U10043 ( .A(n8819), .ZN(n8774) );
  INV_X1 U10044 ( .A(n8772), .ZN(n8773) );
  MUX2_X1 U10045 ( .A(n8774), .B(n8773), .S(n8815), .Z(n8775) );
  NOR2_X1 U10046 ( .A1(n8776), .A2(n8775), .ZN(n8781) );
  NAND2_X1 U10047 ( .A1(n9097), .A2(n5948), .ZN(n8779) );
  OR2_X1 U10048 ( .A1(n8777), .A2(n9764), .ZN(n8778) );
  INV_X1 U10049 ( .A(n10620), .ZN(n8840) );
  INV_X1 U10050 ( .A(n10313), .ZN(n8780) );
  MUX2_X1 U10051 ( .A(n8782), .B(n8781), .S(n10320), .Z(n8783) );
  INV_X1 U10052 ( .A(n10201), .ZN(n8810) );
  OAI21_X1 U10053 ( .B1(n8813), .B2(n6274), .A(n6310), .ZN(n8812) );
  NOR2_X1 U10054 ( .A1(n10320), .A2(n8810), .ZN(n8841) );
  NOR2_X1 U10055 ( .A1(n8814), .A2(n8841), .ZN(n8918) );
  NAND2_X1 U10056 ( .A1(n8896), .A2(n8895), .ZN(n10489) );
  NOR4_X1 U10057 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n8791)
         );
  NAND4_X1 U10058 ( .A1(n8793), .A2(n8792), .A3(n8791), .A4(n8790), .ZN(n8795)
         );
  NOR4_X1 U10059 ( .A1(n8797), .A2(n8796), .A3(n8795), .A4(n8794), .ZN(n8798)
         );
  NAND3_X1 U10060 ( .A1(n8800), .A2(n8799), .A3(n8798), .ZN(n8801) );
  NOR4_X1 U10061 ( .A1(n10489), .A2(n8803), .A3(n8802), .A4(n8801), .ZN(n8805)
         );
  NAND4_X1 U10062 ( .A1(n10463), .A2(n5517), .A3(n8805), .A4(n8804), .ZN(n8806) );
  NOR4_X1 U10063 ( .A1(n10411), .A2(n10423), .A3(n10444), .A4(n8806), .ZN(
        n8807) );
  NAND4_X1 U10064 ( .A1(n10336), .A2(n10389), .A3(n10379), .A4(n8807), .ZN(
        n8808) );
  NOR4_X1 U10065 ( .A1(n8940), .A2(n10358), .A3(n8809), .A4(n8808), .ZN(n8811)
         );
  NAND2_X1 U10066 ( .A1(n10320), .A2(n8810), .ZN(n8820) );
  NAND4_X1 U10067 ( .A1(n8918), .A2(n8811), .A3(n5345), .A4(n8820), .ZN(n8845)
         );
  NAND3_X1 U10068 ( .A1(n8812), .A2(n8923), .A3(n8845), .ZN(n8931) );
  INV_X1 U10069 ( .A(n8814), .ZN(n8842) );
  NAND2_X1 U10070 ( .A1(n8814), .A2(n8782), .ZN(n8816) );
  AOI211_X1 U10071 ( .C1(n8916), .C2(n8923), .A(n8852), .B(n8818), .ZN(n8859)
         );
  NAND2_X1 U10072 ( .A1(n8820), .A2(n8819), .ZN(n8914) );
  NOR2_X1 U10073 ( .A1(n8939), .A2(n8821), .ZN(n8913) );
  NOR3_X1 U10074 ( .A1(n5357), .A2(n8824), .A3(n8823), .ZN(n8907) );
  INV_X1 U10075 ( .A(n8825), .ZN(n8826) );
  AOI21_X1 U10076 ( .B1(n8828), .B2(n8827), .A(n8826), .ZN(n8830) );
  OAI21_X1 U10077 ( .B1(n8830), .B2(n5357), .A(n8829), .ZN(n8905) );
  AOI21_X1 U10078 ( .B1(n8907), .B2(n8831), .A(n8905), .ZN(n8835) );
  INV_X1 U10079 ( .A(n8832), .ZN(n8833) );
  NOR2_X1 U10080 ( .A1(n8834), .A2(n8833), .ZN(n8908) );
  OAI21_X1 U10081 ( .B1(n8835), .B2(n8909), .A(n8908), .ZN(n8837) );
  NAND2_X1 U10082 ( .A1(n8772), .A2(n8836), .ZN(n8911) );
  AOI21_X1 U10083 ( .B1(n8913), .B2(n8837), .A(n8911), .ZN(n8838) );
  AOI211_X1 U10084 ( .C1(n10620), .C2(n10320), .A(n8914), .B(n8838), .ZN(n8839) );
  AOI21_X1 U10085 ( .B1(n8841), .B2(n8840), .A(n8839), .ZN(n8844) );
  OAI211_X1 U10086 ( .C1(n8844), .C2(n8916), .A(n8843), .B(n8842), .ZN(n8846)
         );
  AOI21_X1 U10087 ( .B1(n8846), .B2(n8845), .A(n8923), .ZN(n8847) );
  INV_X1 U10088 ( .A(n8848), .ZN(n10231) );
  NAND2_X1 U10089 ( .A1(n8849), .A2(n10231), .ZN(n8850) );
  OR2_X1 U10090 ( .A1(n8851), .A2(n8850), .ZN(n8855) );
  OAI21_X1 U10091 ( .B1(n8861), .B2(n8852), .A(P1_B_REG_SCAN_IN), .ZN(n8853)
         );
  INV_X1 U10092 ( .A(n8853), .ZN(n8854) );
  NAND2_X1 U10093 ( .A1(n8855), .A2(n8854), .ZN(n8922) );
  INV_X1 U10094 ( .A(n8861), .ZN(n8928) );
  INV_X1 U10095 ( .A(n8922), .ZN(n8927) );
  INV_X1 U10096 ( .A(n8862), .ZN(n8901) );
  INV_X1 U10097 ( .A(n8863), .ZN(n8886) );
  NAND2_X1 U10098 ( .A1(n10214), .A2(n8864), .ZN(n8865) );
  OAI211_X1 U10099 ( .C1(n6861), .C2(n10932), .A(n6310), .B(n8865), .ZN(n8866)
         );
  INV_X1 U10100 ( .A(n8866), .ZN(n8869) );
  OAI211_X1 U10101 ( .C1(n8870), .C2(n8869), .A(n8868), .B(n8867), .ZN(n8872)
         );
  AOI21_X1 U10102 ( .B1(n8872), .B2(n8871), .A(n5370), .ZN(n8875) );
  OAI21_X1 U10103 ( .B1(n8875), .B2(n8874), .A(n8873), .ZN(n8876) );
  NOR2_X1 U10104 ( .A1(n8877), .A2(n8876), .ZN(n8879) );
  OAI21_X1 U10105 ( .B1(n8880), .B2(n8879), .A(n8878), .ZN(n8882) );
  NAND2_X1 U10106 ( .A1(n8882), .A2(n8881), .ZN(n8885) );
  INV_X1 U10107 ( .A(n8883), .ZN(n8884) );
  AOI21_X1 U10108 ( .B1(n8886), .B2(n8885), .A(n8884), .ZN(n8887) );
  NOR2_X1 U10109 ( .A1(n8888), .A2(n8887), .ZN(n8889) );
  OR2_X1 U10110 ( .A1(n8890), .A2(n8889), .ZN(n8892) );
  AOI21_X1 U10111 ( .B1(n8893), .B2(n8892), .A(n8891), .ZN(n8900) );
  NAND2_X1 U10112 ( .A1(n8895), .A2(n8894), .ZN(n8897) );
  NAND2_X1 U10113 ( .A1(n8897), .A2(n8896), .ZN(n8898) );
  OAI211_X1 U10114 ( .C1(n8901), .C2(n8900), .A(n8899), .B(n8898), .ZN(n8902)
         );
  NAND3_X1 U10115 ( .A1(n8904), .A2(n8903), .A3(n8902), .ZN(n8906) );
  AOI21_X1 U10116 ( .B1(n8907), .B2(n8906), .A(n8905), .ZN(n8910) );
  OAI21_X1 U10117 ( .B1(n8910), .B2(n8909), .A(n8908), .ZN(n8912) );
  AOI21_X1 U10118 ( .B1(n8913), .B2(n8912), .A(n8911), .ZN(n8915) );
  OR2_X1 U10119 ( .A1(n8915), .A2(n8914), .ZN(n8917) );
  AOI21_X1 U10120 ( .B1(n8918), .B2(n8917), .A(n8916), .ZN(n8920) );
  NAND3_X1 U10121 ( .A1(n8920), .A2(n8919), .A3(n8922), .ZN(n8926) );
  INV_X1 U10122 ( .A(n8920), .ZN(n8924) );
  NAND4_X1 U10123 ( .A1(n8924), .A2(n8923), .A3(n8922), .A4(n8921), .ZN(n8925)
         );
  OAI211_X1 U10124 ( .C1(n8928), .C2(n8927), .A(n8926), .B(n8925), .ZN(n8929)
         );
  AOI21_X1 U10125 ( .B1(n8931), .B2(n8930), .A(n8929), .ZN(P1_U3242) );
  OAI222_X1 U10126 ( .A1(n6823), .A2(P2_U3151), .B1(n8998), .B2(n8933), .C1(
        n8932), .C2(n8985), .ZN(P2_U3270) );
  NOR2_X2 U10127 ( .A1(n5715), .A2(n10538), .ZN(n10317) );
  AOI211_X1 U10128 ( .C1(n10538), .C2(n5715), .A(n11049), .B(n10317), .ZN(
        n10537) );
  INV_X1 U10129 ( .A(n10538), .ZN(n8938) );
  INV_X1 U10130 ( .A(n8935), .ZN(n8936) );
  AOI22_X1 U10131 ( .A1(n8936), .A2(n10521), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10466), .ZN(n8937) );
  OAI21_X1 U10132 ( .B1(n8938), .B2(n10525), .A(n8937), .ZN(n8948) );
  XNOR2_X1 U10133 ( .A(n8941), .B(n8940), .ZN(n8947) );
  NAND2_X1 U10134 ( .A1(n10338), .A2(n10507), .ZN(n8946) );
  INV_X1 U10135 ( .A(P1_B_REG_SCAN_IN), .ZN(n8942) );
  NOR2_X1 U10136 ( .A1(n10748), .A2(n8942), .ZN(n8943) );
  NOR2_X1 U10137 ( .A1(n8944), .A2(n8943), .ZN(n10312) );
  NAND2_X1 U10138 ( .A1(n10201), .A2(n10312), .ZN(n8945) );
  OAI222_X1 U10139 ( .A1(n10659), .A2(n9760), .B1(n7742), .B2(n8949), .C1(
        n5736), .C2(P1_U3086), .ZN(P1_U3326) );
  AND2_X1 U10140 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  XNOR2_X1 U10141 ( .A(n10028), .B(n7550), .ZN(n8955) );
  XNOR2_X1 U10142 ( .A(n8955), .B(n9962), .ZN(n9016) );
  XNOR2_X1 U10143 ( .A(n9972), .B(n7550), .ZN(n8958) );
  XNOR2_X1 U10144 ( .A(n8958), .B(n8957), .ZN(n9052) );
  XNOR2_X1 U10145 ( .A(n10020), .B(n8959), .ZN(n8960) );
  NAND2_X1 U10146 ( .A1(n8960), .A2(n9963), .ZN(n9023) );
  XNOR2_X1 U10147 ( .A(n10016), .B(n7550), .ZN(n8961) );
  XNOR2_X1 U10148 ( .A(n8961), .B(n9947), .ZN(n9064) );
  XNOR2_X1 U10149 ( .A(n10012), .B(n7550), .ZN(n8964) );
  INV_X1 U10150 ( .A(n8963), .ZN(n8965) );
  XNOR2_X1 U10151 ( .A(n10008), .B(n7550), .ZN(n8969) );
  XNOR2_X1 U10152 ( .A(n8969), .B(n8967), .ZN(n9044) );
  NAND2_X1 U10153 ( .A1(n8969), .A2(n8967), .ZN(n8970) );
  XNOR2_X1 U10154 ( .A(n9906), .B(n7550), .ZN(n8972) );
  XNOR2_X1 U10155 ( .A(n8972), .B(n9914), .ZN(n9034) );
  XNOR2_X1 U10156 ( .A(n10000), .B(n7550), .ZN(n8973) );
  XOR2_X1 U10157 ( .A(n9251), .B(n8973), .Z(n9078) );
  INV_X1 U10158 ( .A(n8973), .ZN(n8974) );
  INV_X1 U10159 ( .A(n9251), .ZN(n9319) );
  NAND2_X1 U10160 ( .A1(n8974), .A2(n9319), .ZN(n8975) );
  XNOR2_X1 U10161 ( .A(n9996), .B(n7550), .ZN(n8976) );
  NOR2_X1 U10162 ( .A1(n8976), .A2(n9079), .ZN(n8977) );
  AOI21_X1 U10163 ( .B1(n9079), .B2(n8976), .A(n8977), .ZN(n9001) );
  XNOR2_X1 U10164 ( .A(n9448), .B(n7550), .ZN(n8978) );
  XNOR2_X1 U10165 ( .A(n8979), .B(n8978), .ZN(n8984) );
  OAI22_X1 U10166 ( .A1(n9067), .A2(n9079), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9522), .ZN(n8980) );
  AOI21_X1 U10167 ( .B1(n9080), .B2(n9441), .A(n8980), .ZN(n8981) );
  OAI21_X1 U10168 ( .B1(n9082), .B2(n9445), .A(n8981), .ZN(n8982) );
  AOI21_X1 U10169 ( .B1(n9992), .B2(n9059), .A(n8982), .ZN(n8983) );
  OAI21_X1 U10170 ( .B1(n8984), .B2(n9061), .A(n8983), .ZN(P2_U3160) );
  OAI222_X1 U10171 ( .A1(n6819), .A2(P2_U3151), .B1(n8998), .B2(n8987), .C1(
        n8986), .C2(n8985), .ZN(P2_U3271) );
  AOI22_X1 U10172 ( .A1(n10981), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n9433), 
        .B2(n11041), .ZN(n8991) );
  OAI21_X1 U10173 ( .B1(n8992), .B2(n9984), .A(n8991), .ZN(n8993) );
  AOI21_X1 U10174 ( .B1(n8990), .B2(n8994), .A(n8993), .ZN(n8995) );
  OAI21_X1 U10175 ( .B1(n8989), .B2(n9958), .A(n8995), .ZN(P2_U3204) );
  OAI222_X1 U10176 ( .A1(n8985), .A2(n9098), .B1(n8998), .B2(n8997), .C1(n8996), .C2(P2_U3151), .ZN(P2_U3265) );
  OAI211_X1 U10177 ( .C1(n8999), .C2(n9001), .A(n9000), .B(n9076), .ZN(n9006)
         );
  INV_X1 U10178 ( .A(n9878), .ZN(n9004) );
  AOI22_X1 U10179 ( .A1(n9080), .A2(n9874), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n9002) );
  OAI21_X1 U10180 ( .B1(n9251), .B2(n9067), .A(n9002), .ZN(n9003) );
  AOI21_X1 U10181 ( .B1(n9071), .B2(n9004), .A(n9003), .ZN(n9005) );
  OAI211_X1 U10182 ( .C1(n9007), .C2(n9088), .A(n9006), .B(n9005), .ZN(
        P2_U3154) );
  INV_X1 U10183 ( .A(n10012), .ZN(n9929) );
  OAI211_X1 U10184 ( .C1(n9009), .C2(n9934), .A(n9008), .B(n9076), .ZN(n9014)
         );
  INV_X1 U10185 ( .A(n9010), .ZN(n9927) );
  AOI22_X1 U10186 ( .A1(n9080), .A2(n9923), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n9011) );
  OAI21_X1 U10187 ( .B1(n9230), .B2(n9067), .A(n9011), .ZN(n9012) );
  AOI21_X1 U10188 ( .B1(n9071), .B2(n9927), .A(n9012), .ZN(n9013) );
  OAI211_X1 U10189 ( .C1(n9929), .C2(n9088), .A(n9014), .B(n9013), .ZN(
        P2_U3156) );
  INV_X1 U10190 ( .A(n10028), .ZN(n9985) );
  OAI211_X1 U10191 ( .C1(n5183), .C2(n9016), .A(n9015), .B(n9076), .ZN(n9022)
         );
  NAND2_X1 U10192 ( .A1(n9946), .A2(n10944), .ZN(n9018) );
  NAND2_X1 U10193 ( .A1(n9320), .A2(n9961), .ZN(n9017) );
  AND2_X1 U10194 ( .A1(n9018), .A2(n9017), .ZN(n9978) );
  OAI22_X1 U10195 ( .A1(n9978), .A2(n9019), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9518), .ZN(n9020) );
  AOI21_X1 U10196 ( .B1(n9071), .B2(n9982), .A(n9020), .ZN(n9021) );
  OAI211_X1 U10197 ( .C1(n9985), .C2(n9088), .A(n9022), .B(n9021), .ZN(
        P2_U3159) );
  NAND2_X1 U10198 ( .A1(n5180), .A2(n9023), .ZN(n9024) );
  XNOR2_X1 U10199 ( .A(n9025), .B(n9024), .ZN(n9032) );
  NAND2_X1 U10200 ( .A1(n9080), .A2(n9947), .ZN(n9026) );
  OAI21_X1 U10201 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n9027), .A(n9026), .ZN(
        n9028) );
  AOI21_X1 U10202 ( .B1(n9085), .B2(n9946), .A(n9028), .ZN(n9029) );
  OAI21_X1 U10203 ( .B1(n9949), .B2(n9082), .A(n9029), .ZN(n9030) );
  AOI21_X1 U10204 ( .B1(n10020), .B2(n9059), .A(n9030), .ZN(n9031) );
  OAI21_X1 U10205 ( .B1(n9032), .B2(n9061), .A(n9031), .ZN(P2_U3163) );
  XOR2_X1 U10206 ( .A(n9034), .B(n9033), .Z(n9040) );
  NAND2_X1 U10207 ( .A1(n9080), .A2(n9319), .ZN(n9035) );
  OAI21_X1 U10208 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n9735), .A(n9035), .ZN(
        n9036) );
  AOI21_X1 U10209 ( .B1(n9085), .B2(n9923), .A(n9036), .ZN(n9037) );
  OAI21_X1 U10210 ( .B1(n9907), .B2(n9082), .A(n9037), .ZN(n9038) );
  AOI21_X1 U10211 ( .B1(n9906), .B2(n9059), .A(n9038), .ZN(n9039) );
  OAI21_X1 U10212 ( .B1(n9040), .B2(n9061), .A(n9039), .ZN(P2_U3165) );
  INV_X1 U10213 ( .A(n9041), .ZN(n9042) );
  AOI21_X1 U10214 ( .B1(n9044), .B2(n9043), .A(n9042), .ZN(n9051) );
  NAND2_X1 U10215 ( .A1(n9080), .A2(n9914), .ZN(n9045) );
  OAI21_X1 U10216 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n9540), .A(n9045), .ZN(
        n9046) );
  AOI21_X1 U10217 ( .B1(n9085), .B2(n9934), .A(n9046), .ZN(n9047) );
  OAI21_X1 U10218 ( .B1(n9048), .B2(n9082), .A(n9047), .ZN(n9049) );
  AOI21_X1 U10219 ( .B1(n10008), .B2(n9059), .A(n9049), .ZN(n9050) );
  OAI21_X1 U10220 ( .B1(n9051), .B2(n9061), .A(n9050), .ZN(P2_U3169) );
  XNOR2_X1 U10221 ( .A(n9053), .B(n9052), .ZN(n9062) );
  NAND2_X1 U10222 ( .A1(n9080), .A2(n9963), .ZN(n9054) );
  OAI21_X1 U10223 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n9535), .A(n9054), .ZN(
        n9055) );
  AOI21_X1 U10224 ( .B1(n9085), .B2(n9962), .A(n9055), .ZN(n9056) );
  OAI21_X1 U10225 ( .B1(n9057), .B2(n9082), .A(n9056), .ZN(n9058) );
  AOI21_X1 U10226 ( .B1(n10024), .B2(n9059), .A(n9058), .ZN(n9060) );
  OAI21_X1 U10227 ( .B1(n9062), .B2(n9061), .A(n9060), .ZN(P2_U3173) );
  INV_X1 U10228 ( .A(n10016), .ZN(n9074) );
  OAI211_X1 U10229 ( .C1(n9065), .C2(n9064), .A(n9063), .B(n9076), .ZN(n9073)
         );
  INV_X1 U10230 ( .A(n9936), .ZN(n9070) );
  AOI22_X1 U10231 ( .A1(n9080), .A2(n9934), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n9066) );
  OAI21_X1 U10232 ( .B1(n9068), .B2(n9067), .A(n9066), .ZN(n9069) );
  AOI21_X1 U10233 ( .B1(n9071), .B2(n9070), .A(n9069), .ZN(n9072) );
  OAI211_X1 U10234 ( .C1(n9074), .C2(n9088), .A(n9073), .B(n9072), .ZN(
        P2_U3175) );
  OAI211_X1 U10235 ( .C1(n9075), .C2(n9078), .A(n9077), .B(n9076), .ZN(n9087)
         );
  NAND2_X1 U10236 ( .A1(n9080), .A2(n5433), .ZN(n9081) );
  OAI21_X1 U10237 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n9762), .A(n9081), .ZN(
        n9084) );
  NOR2_X1 U10238 ( .A1(n9082), .A2(n9889), .ZN(n9083) );
  AOI211_X1 U10239 ( .C1(n9085), .C2(n9914), .A(n9084), .B(n9083), .ZN(n9086)
         );
  OAI211_X1 U10240 ( .C1(n9089), .C2(n9088), .A(n9087), .B(n9086), .ZN(
        P2_U3180) );
  NAND2_X1 U10241 ( .A1(n5121), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9095) );
  INV_X1 U10242 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9090) );
  OR2_X1 U10243 ( .A1(n9091), .A2(n9090), .ZN(n9094) );
  INV_X1 U10244 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9092) );
  OR2_X1 U10245 ( .A1(n6733), .A2(n9092), .ZN(n9093) );
  NAND4_X1 U10246 ( .A1(n9096), .A2(n9095), .A3(n9094), .A4(n9093), .ZN(n9318)
         );
  NAND2_X1 U10247 ( .A1(n9097), .A2(n6499), .ZN(n9100) );
  OR2_X1 U10248 ( .A1(n9101), .A2(n9098), .ZN(n9099) );
  NAND2_X1 U10249 ( .A1(n9100), .A2(n9099), .ZN(n9107) );
  OR2_X1 U10250 ( .A1(n9107), .A2(n9106), .ZN(n9266) );
  NAND2_X1 U10251 ( .A1(n10664), .A2(n6499), .ZN(n9103) );
  OR2_X1 U10252 ( .A1(n9101), .A2(n7211), .ZN(n9102) );
  AOI21_X1 U10253 ( .B1(n9318), .B2(n9266), .A(n9989), .ZN(n9105) );
  NOR2_X1 U10254 ( .A1(n9105), .A2(n9104), .ZN(n9309) );
  INV_X1 U10255 ( .A(n9107), .ZN(n9991) );
  INV_X1 U10256 ( .A(n9318), .ZN(n9435) );
  OR2_X1 U10257 ( .A1(n9306), .A2(n9435), .ZN(n9109) );
  NAND2_X1 U10258 ( .A1(n9107), .A2(n9106), .ZN(n9108) );
  NAND2_X1 U10259 ( .A1(n9109), .A2(n9108), .ZN(n9269) );
  INV_X1 U10260 ( .A(n9441), .ZN(n9264) );
  NAND2_X1 U10261 ( .A1(n6797), .A2(n9264), .ZN(n9267) );
  INV_X1 U10262 ( .A(n9267), .ZN(n9110) );
  OR2_X1 U10263 ( .A1(n9269), .A2(n9110), .ZN(n9305) );
  INV_X1 U10264 ( .A(n9305), .ZN(n9111) );
  OAI211_X1 U10265 ( .C1(n9991), .C2(n9306), .A(n9112), .B(n9111), .ZN(n9308)
         );
  OR2_X1 U10266 ( .A1(n9992), .A2(n9244), .ZN(n9114) );
  OR2_X1 U10267 ( .A1(n9874), .A2(n5127), .ZN(n9113) );
  NAND2_X1 U10268 ( .A1(n9114), .A2(n9113), .ZN(n9262) );
  MUX2_X1 U10269 ( .A(n9239), .B(n9240), .S(n9244), .Z(n9243) );
  INV_X1 U10270 ( .A(n9115), .ZN(n9235) );
  INV_X1 U10271 ( .A(n9925), .ZN(n9234) );
  AND2_X1 U10272 ( .A1(n9967), .A2(n9116), .ZN(n9117) );
  MUX2_X1 U10273 ( .A(n9118), .B(n9117), .S(n9244), .Z(n9218) );
  AND2_X1 U10274 ( .A1(n9196), .A2(n6768), .ZN(n9289) );
  NAND2_X1 U10275 ( .A1(n9121), .A2(n9120), .ZN(n9122) );
  NAND3_X1 U10276 ( .A1(n9122), .A2(n9127), .A3(n9124), .ZN(n9123) );
  NAND2_X1 U10277 ( .A1(n9123), .A2(n9125), .ZN(n9130) );
  INV_X1 U10278 ( .A(n9124), .ZN(n9126) );
  NAND2_X1 U10279 ( .A1(n9126), .A2(n9125), .ZN(n9128) );
  NAND2_X1 U10280 ( .A1(n9128), .A2(n9127), .ZN(n9129) );
  MUX2_X1 U10281 ( .A(n9130), .B(n9129), .S(n5127), .Z(n9131) );
  NAND2_X1 U10282 ( .A1(n9131), .A2(n10966), .ZN(n9139) );
  NAND2_X1 U10283 ( .A1(n9149), .A2(n9132), .ZN(n9135) );
  NAND2_X1 U10284 ( .A1(n9142), .A2(n9133), .ZN(n9134) );
  MUX2_X1 U10285 ( .A(n9135), .B(n9134), .S(n9244), .Z(n9136) );
  INV_X1 U10286 ( .A(n9136), .ZN(n9138) );
  AOI21_X1 U10287 ( .B1(n9139), .B2(n9138), .A(n9137), .ZN(n9150) );
  NAND2_X1 U10288 ( .A1(n9140), .A2(n9143), .ZN(n9141) );
  AOI21_X1 U10289 ( .B1(n9150), .B2(n9142), .A(n9141), .ZN(n9145) );
  NAND2_X1 U10290 ( .A1(n9155), .A2(n9143), .ZN(n9144) );
  MUX2_X1 U10291 ( .A(n9145), .B(n9144), .S(n9244), .Z(n9163) );
  NAND2_X1 U10292 ( .A1(n9156), .A2(n9147), .ZN(n9152) );
  NAND2_X1 U10293 ( .A1(n9147), .A2(n9146), .ZN(n9148) );
  AOI21_X1 U10294 ( .B1(n9150), .B2(n9149), .A(n9148), .ZN(n9151) );
  MUX2_X1 U10295 ( .A(n9152), .B(n9151), .S(n9244), .Z(n9162) );
  INV_X1 U10296 ( .A(n9171), .ZN(n9161) );
  INV_X1 U10297 ( .A(n9155), .ZN(n9158) );
  INV_X1 U10298 ( .A(n9156), .ZN(n9157) );
  MUX2_X1 U10299 ( .A(n9158), .B(n9157), .S(n9244), .Z(n9159) );
  NOR2_X1 U10300 ( .A1(n9159), .A2(n9279), .ZN(n9160) );
  OAI211_X1 U10301 ( .C1(n9163), .C2(n9162), .A(n9161), .B(n9160), .ZN(n9176)
         );
  AND2_X1 U10302 ( .A1(n9165), .A2(n9164), .ZN(n9168) );
  OAI211_X1 U10303 ( .C1(n9171), .C2(n9168), .A(n9167), .B(n9166), .ZN(n9173)
         );
  OAI21_X1 U10304 ( .B1(n9171), .B2(n9170), .A(n9169), .ZN(n9172) );
  MUX2_X1 U10305 ( .A(n9173), .B(n9172), .S(n9244), .Z(n9174) );
  INV_X1 U10306 ( .A(n9174), .ZN(n9175) );
  NAND3_X1 U10307 ( .A1(n9176), .A2(n9285), .A3(n9175), .ZN(n9188) );
  NAND2_X1 U10308 ( .A1(n9180), .A2(n9177), .ZN(n9179) );
  AND2_X1 U10309 ( .A1(n9179), .A2(n9178), .ZN(n9184) );
  INV_X1 U10310 ( .A(n9180), .ZN(n9181) );
  NOR2_X1 U10311 ( .A1(n9182), .A2(n9181), .ZN(n9183) );
  MUX2_X1 U10312 ( .A(n9184), .B(n9183), .S(n9244), .Z(n9186) );
  NOR2_X1 U10313 ( .A1(n9186), .A2(n9185), .ZN(n9187) );
  INV_X1 U10314 ( .A(n9189), .ZN(n9190) );
  OAI21_X1 U10315 ( .B1(n9191), .B2(n9190), .A(n5127), .ZN(n9192) );
  OAI211_X1 U10316 ( .C1(n9194), .C2(n9198), .A(n9193), .B(n9192), .ZN(n9211)
         );
  AND2_X1 U10317 ( .A1(n9196), .A2(n6767), .ZN(n9200) );
  NAND2_X1 U10318 ( .A1(n9205), .A2(n9201), .ZN(n9202) );
  NAND2_X1 U10319 ( .A1(n9202), .A2(n9204), .ZN(n9208) );
  NAND2_X1 U10320 ( .A1(n9204), .A2(n9203), .ZN(n9206) );
  NAND2_X1 U10321 ( .A1(n9206), .A2(n9205), .ZN(n9207) );
  MUX2_X1 U10322 ( .A(n9208), .B(n9207), .S(n5127), .Z(n9209) );
  OAI21_X1 U10323 ( .B1(n9211), .B2(n9210), .A(n9209), .ZN(n9212) );
  NAND2_X1 U10324 ( .A1(n9212), .A2(n9295), .ZN(n9216) );
  MUX2_X1 U10325 ( .A(n9214), .B(n9213), .S(n5127), .Z(n9215) );
  NAND3_X1 U10326 ( .A1(n9216), .A2(n9296), .A3(n9215), .ZN(n9217) );
  NAND3_X1 U10327 ( .A1(n9218), .A2(n9221), .A3(n9217), .ZN(n9219) );
  OAI21_X1 U10328 ( .B1(n9220), .B2(n9244), .A(n9219), .ZN(n9224) );
  AOI21_X1 U10329 ( .B1(n9223), .B2(n9221), .A(n5127), .ZN(n9222) );
  OAI21_X1 U10330 ( .B1(n5127), .B2(n9225), .A(n9952), .ZN(n9229) );
  MUX2_X1 U10331 ( .A(n9227), .B(n9226), .S(n9244), .Z(n9228) );
  NAND2_X1 U10332 ( .A1(n10016), .A2(n9230), .ZN(n9231) );
  MUX2_X1 U10333 ( .A(n9232), .B(n9231), .S(n9244), .Z(n9233) );
  MUX2_X1 U10334 ( .A(n9236), .B(n9235), .S(n5127), .Z(n9237) );
  INV_X1 U10335 ( .A(n9237), .ZN(n9238) );
  NAND2_X1 U10336 ( .A1(n9241), .A2(n9913), .ZN(n9242) );
  NAND3_X1 U10337 ( .A1(n9899), .A2(n9243), .A3(n9242), .ZN(n9248) );
  MUX2_X1 U10338 ( .A(n9246), .B(n9245), .S(n9244), .Z(n9247) );
  NAND2_X1 U10339 ( .A1(n9248), .A2(n9247), .ZN(n9256) );
  OAI21_X1 U10340 ( .B1(n9256), .B2(n9251), .A(n10000), .ZN(n9249) );
  NAND2_X1 U10341 ( .A1(n9249), .A2(n9254), .ZN(n9250) );
  NAND2_X1 U10342 ( .A1(n9250), .A2(n9244), .ZN(n9258) );
  NOR2_X1 U10343 ( .A1(n9251), .A2(n9244), .ZN(n9903) );
  NOR2_X1 U10344 ( .A1(n9251), .A2(n5127), .ZN(n9253) );
  NAND2_X1 U10345 ( .A1(n9256), .A2(n9903), .ZN(n9252) );
  OAI21_X1 U10346 ( .B1(n9253), .B2(n10000), .A(n9252), .ZN(n9255) );
  OAI211_X1 U10347 ( .C1(n9903), .C2(n9256), .A(n9255), .B(n9254), .ZN(n9257)
         );
  NAND2_X1 U10348 ( .A1(n9258), .A2(n9257), .ZN(n9260) );
  MUX2_X1 U10349 ( .A(n5127), .B(n9260), .S(n9259), .Z(n9263) );
  MUX2_X1 U10350 ( .A(n9874), .B(n9992), .S(n9244), .Z(n9261) );
  OR2_X1 U10351 ( .A1(n6797), .A2(n9264), .ZN(n9265) );
  NAND2_X1 U10352 ( .A1(n9266), .A2(n9265), .ZN(n9304) );
  NOR2_X1 U10353 ( .A1(n9270), .A2(n10937), .ZN(n9276) );
  NOR2_X1 U10354 ( .A1(n9272), .A2(n9271), .ZN(n9274) );
  NAND4_X1 U10355 ( .A1(n9276), .A2(n9275), .A3(n9274), .A4(n9273), .ZN(n9280)
         );
  NOR4_X1 U10356 ( .A1(n9280), .A2(n9279), .A3(n9278), .A4(n9277), .ZN(n9284)
         );
  NAND4_X1 U10357 ( .A1(n9284), .A2(n6765), .A3(n9283), .A4(n9282), .ZN(n9287)
         );
  INV_X1 U10358 ( .A(n9285), .ZN(n9286) );
  NOR2_X1 U10359 ( .A1(n9287), .A2(n9286), .ZN(n9288) );
  NAND4_X1 U10360 ( .A1(n9291), .A2(n9290), .A3(n9289), .A4(n9288), .ZN(n9293)
         );
  NOR2_X1 U10361 ( .A1(n9293), .A2(n9292), .ZN(n9294) );
  NAND3_X1 U10362 ( .A1(n9296), .A2(n9295), .A3(n9294), .ZN(n9297) );
  NOR2_X1 U10363 ( .A1(n9980), .A2(n9297), .ZN(n9298) );
  NAND3_X1 U10364 ( .A1(n9952), .A2(n9969), .A3(n9298), .ZN(n9299) );
  NOR3_X1 U10365 ( .A1(n9925), .A2(n9932), .A3(n9299), .ZN(n9300) );
  NAND3_X1 U10366 ( .A1(n9899), .A2(n9913), .A3(n9300), .ZN(n9301) );
  NOR3_X1 U10367 ( .A1(n9883), .A2(n9887), .A3(n9301), .ZN(n9302) );
  NAND2_X1 U10368 ( .A1(n9448), .A2(n9302), .ZN(n9303) );
  OR3_X1 U10369 ( .A1(n9305), .A2(n9304), .A3(n9303), .ZN(n9307) );
  XNOR2_X1 U10370 ( .A(n9310), .B(n9409), .ZN(n9317) );
  NOR3_X1 U10371 ( .A1(n9312), .A2(n9311), .A3(n6788), .ZN(n9315) );
  OAI21_X1 U10372 ( .B1(n9316), .B2(n9313), .A(P2_B_REG_SCAN_IN), .ZN(n9314)
         );
  OAI22_X1 U10373 ( .A1(n9317), .A2(n9316), .B1(n9315), .B2(n9314), .ZN(
        P2_U3296) );
  MUX2_X1 U10374 ( .A(n9318), .B(P2_DATAO_REG_31__SCAN_IN), .S(n9336), .Z(
        P2_U3522) );
  MUX2_X1 U10375 ( .A(n9441), .B(P2_DATAO_REG_29__SCAN_IN), .S(n9336), .Z(
        P2_U3520) );
  MUX2_X1 U10376 ( .A(n9874), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9336), .Z(
        P2_U3519) );
  MUX2_X1 U10377 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n5433), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10378 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9319), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10379 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9914), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10380 ( .A(n9923), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9336), .Z(
        P2_U3515) );
  MUX2_X1 U10381 ( .A(n9934), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9336), .Z(
        P2_U3514) );
  MUX2_X1 U10382 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9947), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10383 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9963), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10384 ( .A(n9946), .B(P2_DATAO_REG_20__SCAN_IN), .S(n9336), .Z(
        P2_U3511) );
  MUX2_X1 U10385 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9962), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10386 ( .A(n9320), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9336), .Z(
        P2_U3509) );
  MUX2_X1 U10387 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9321), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10388 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9322), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10389 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9323), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10390 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9324), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10391 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9325), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10392 ( .A(n9326), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9336), .Z(
        P2_U3503) );
  MUX2_X1 U10393 ( .A(n9327), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9336), .Z(
        P2_U3502) );
  MUX2_X1 U10394 ( .A(n9328), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9336), .Z(
        P2_U3501) );
  MUX2_X1 U10395 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n9329), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10396 ( .A(n9330), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9336), .Z(
        P2_U3498) );
  MUX2_X1 U10397 ( .A(n9331), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9336), .Z(
        P2_U3497) );
  MUX2_X1 U10398 ( .A(n9332), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9336), .Z(
        P2_U3496) );
  MUX2_X1 U10399 ( .A(n9333), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9336), .Z(
        P2_U3495) );
  MUX2_X1 U10400 ( .A(n9334), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9336), .Z(
        P2_U3494) );
  MUX2_X1 U10401 ( .A(n9335), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9336), .Z(
        P2_U3493) );
  MUX2_X1 U10402 ( .A(n6408), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9336), .Z(
        P2_U3492) );
  MUX2_X1 U10403 ( .A(n9337), .B(P2_DATAO_REG_0__SCAN_IN), .S(n9336), .Z(
        P2_U3491) );
  AOI21_X1 U10404 ( .B1(n9340), .B2(n9339), .A(n9338), .ZN(n9356) );
  AOI21_X1 U10405 ( .B1(n5182), .B2(n9342), .A(n9341), .ZN(n9343) );
  NOR2_X1 U10406 ( .A1(n9343), .A2(n10915), .ZN(n9354) );
  INV_X1 U10407 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9352) );
  OAI21_X1 U10408 ( .B1(n9346), .B2(n9345), .A(n9344), .ZN(n9350) );
  OAI22_X1 U10409 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9348), .B1(n10904), .B2(
        n9347), .ZN(n9349) );
  AOI21_X1 U10410 ( .B1(n9350), .B2(n10923), .A(n9349), .ZN(n9351) );
  OAI21_X1 U10411 ( .B1(n9422), .B2(n9352), .A(n9351), .ZN(n9353) );
  NOR2_X1 U10412 ( .A1(n9354), .A2(n9353), .ZN(n9355) );
  OAI21_X1 U10413 ( .B1(n9356), .B2(n10918), .A(n9355), .ZN(P2_U3196) );
  AOI21_X1 U10414 ( .B1(n8600), .B2(n9358), .A(n9357), .ZN(n9373) );
  INV_X1 U10415 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9369) );
  AND2_X1 U10416 ( .A1(n9359), .A2(n8599), .ZN(n9360) );
  OAI21_X1 U10417 ( .B1(n9361), .B2(n9360), .A(n9429), .ZN(n9368) );
  OAI21_X1 U10418 ( .B1(n9364), .B2(n9363), .A(n9362), .ZN(n9366) );
  AOI21_X1 U10419 ( .B1(n9366), .B2(n10923), .A(n9365), .ZN(n9367) );
  OAI211_X1 U10420 ( .C1(n9369), .C2(n9422), .A(n9368), .B(n9367), .ZN(n9370)
         );
  AOI21_X1 U10421 ( .B1(n9371), .B2(n10906), .A(n9370), .ZN(n9372) );
  OAI21_X1 U10422 ( .B1(n9373), .B2(n10918), .A(n9372), .ZN(P2_U3197) );
  AOI21_X1 U10423 ( .B1(n5158), .B2(n9375), .A(n9374), .ZN(n9389) );
  AOI21_X1 U10424 ( .B1(n9378), .B2(n9377), .A(n9376), .ZN(n9379) );
  OR2_X1 U10425 ( .A1(n9379), .A2(n10918), .ZN(n9388) );
  OAI22_X1 U10426 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9381), .B1(n10904), .B2(
        n9380), .ZN(n9386) );
  XOR2_X1 U10427 ( .A(n9383), .B(n9382), .Z(n9384) );
  NOR2_X1 U10428 ( .A1(n9384), .A2(n9426), .ZN(n9385) );
  AOI211_X1 U10429 ( .C1(n10907), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n9386), .B(
        n9385), .ZN(n9387) );
  OAI211_X1 U10430 ( .C1(n9389), .C2(n10915), .A(n9388), .B(n9387), .ZN(
        P2_U3198) );
  AOI21_X1 U10431 ( .B1(n6615), .B2(n9391), .A(n9390), .ZN(n9404) );
  XNOR2_X1 U10432 ( .A(n9393), .B(n9392), .ZN(n9402) );
  AOI21_X1 U10433 ( .B1(n9395), .B2(n11152), .A(n9394), .ZN(n9400) );
  OAI22_X1 U10434 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9397), .B1(n10904), .B2(
        n9396), .ZN(n9398) );
  AOI21_X1 U10435 ( .B1(n10907), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9398), .ZN(
        n9399) );
  OAI21_X1 U10436 ( .B1(n9400), .B2(n10915), .A(n9399), .ZN(n9401) );
  AOI21_X1 U10437 ( .B1(n10923), .B2(n9402), .A(n9401), .ZN(n9403) );
  OAI21_X1 U10438 ( .B1(n9404), .B2(n10918), .A(n9403), .ZN(P2_U3199) );
  MUX2_X1 U10439 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n6649), .S(n9409), .Z(n9413) );
  XNOR2_X1 U10440 ( .A(n9407), .B(n9413), .ZN(n9432) );
  XNOR2_X1 U10441 ( .A(n9409), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9411) );
  XNOR2_X1 U10442 ( .A(n9410), .B(n9411), .ZN(n9430) );
  INV_X1 U10443 ( .A(n9411), .ZN(n9414) );
  MUX2_X1 U10444 ( .A(n9414), .B(n9413), .S(n9311), .Z(n9419) );
  AOI21_X1 U10445 ( .B1(n9417), .B2(n9416), .A(n9415), .ZN(n9418) );
  XOR2_X1 U10446 ( .A(n9419), .B(n9418), .Z(n9427) );
  NAND2_X1 U10447 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n9420) );
  OAI21_X1 U10448 ( .B1(n9422), .B2(n9421), .A(n9420), .ZN(n9423) );
  AOI21_X1 U10449 ( .B1(n9424), .B2(n10906), .A(n9423), .ZN(n9425) );
  OAI21_X1 U10450 ( .B1(n9427), .B2(n9426), .A(n9425), .ZN(n9428) );
  AOI21_X1 U10451 ( .B1(n9430), .B2(n9429), .A(n9428), .ZN(n9431) );
  OAI21_X1 U10452 ( .B1(n10918), .B2(n9432), .A(n9431), .ZN(P2_U3201) );
  AOI21_X1 U10453 ( .B1(n11041), .B2(n9433), .A(n9958), .ZN(n9436) );
  NAND2_X1 U10454 ( .A1(n9436), .A2(n9990), .ZN(n9438) );
  OAI21_X1 U10455 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n11048), .A(n9438), .ZN(
        n9437) );
  OAI21_X1 U10456 ( .B1(n9989), .B2(n9984), .A(n9437), .ZN(P2_U3202) );
  OAI21_X1 U10457 ( .B1(P2_REG2_REG_30__SCAN_IN), .B2(n11048), .A(n9438), .ZN(
        n9439) );
  OAI21_X1 U10458 ( .B1(n9991), .B2(n9984), .A(n9439), .ZN(P2_U3203) );
  NAND2_X1 U10459 ( .A1(n9441), .A2(n10944), .ZN(n9442) );
  OAI22_X1 U10460 ( .A1(n11048), .A2(n9446), .B1(n9445), .B2(n10950), .ZN(
        n9451) );
  OAI21_X1 U10461 ( .B1(n9449), .B2(n9448), .A(n9447), .ZN(n9995) );
  NOR2_X1 U10462 ( .A1(n9995), .A2(n9954), .ZN(n9450) );
  AOI211_X1 U10463 ( .C1(n11043), .C2(n9992), .A(n9451), .B(n9450), .ZN(n9452)
         );
  OAI21_X1 U10464 ( .B1(n9994), .B2(n10981), .A(n9452), .ZN(n9871) );
  XOR2_X1 U10465 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n9455) );
  XNOR2_X1 U10466 ( .A(n9657), .B(keyinput_1), .ZN(n9454) );
  XNOR2_X1 U10467 ( .A(SI_30_), .B(keyinput_2), .ZN(n9453) );
  NAND3_X1 U10468 ( .A1(n9455), .A2(n9454), .A3(n9453), .ZN(n9458) );
  XNOR2_X1 U10469 ( .A(SI_29_), .B(keyinput_3), .ZN(n9457) );
  XNOR2_X1 U10470 ( .A(SI_28_), .B(keyinput_4), .ZN(n9456) );
  AOI21_X1 U10471 ( .B1(n9458), .B2(n9457), .A(n9456), .ZN(n9466) );
  XNOR2_X1 U10472 ( .A(n9459), .B(keyinput_5), .ZN(n9465) );
  XNOR2_X1 U10473 ( .A(n9666), .B(keyinput_6), .ZN(n9463) );
  XNOR2_X1 U10474 ( .A(n9460), .B(keyinput_7), .ZN(n9462) );
  XNOR2_X1 U10475 ( .A(SI_24_), .B(keyinput_8), .ZN(n9461) );
  NOR3_X1 U10476 ( .A1(n9463), .A2(n9462), .A3(n9461), .ZN(n9464) );
  OAI21_X1 U10477 ( .B1(n9466), .B2(n9465), .A(n9464), .ZN(n9473) );
  XNOR2_X1 U10478 ( .A(n9674), .B(keyinput_9), .ZN(n9472) );
  XNOR2_X1 U10479 ( .A(n9467), .B(keyinput_11), .ZN(n9470) );
  XNOR2_X1 U10480 ( .A(n9675), .B(keyinput_12), .ZN(n9469) );
  XNOR2_X1 U10481 ( .A(SI_22_), .B(keyinput_10), .ZN(n9468) );
  NAND3_X1 U10482 ( .A1(n9470), .A2(n9469), .A3(n9468), .ZN(n9471) );
  AOI21_X1 U10483 ( .B1(n9473), .B2(n9472), .A(n9471), .ZN(n9477) );
  XNOR2_X1 U10484 ( .A(n9474), .B(keyinput_13), .ZN(n9476) );
  XNOR2_X1 U10485 ( .A(n9655), .B(keyinput_14), .ZN(n9475) );
  OAI21_X1 U10486 ( .B1(n9477), .B2(n9476), .A(n9475), .ZN(n9481) );
  XNOR2_X1 U10487 ( .A(n9652), .B(keyinput_16), .ZN(n9480) );
  XNOR2_X1 U10488 ( .A(n9478), .B(keyinput_15), .ZN(n9479) );
  NAND3_X1 U10489 ( .A1(n9481), .A2(n9480), .A3(n9479), .ZN(n9485) );
  XNOR2_X1 U10490 ( .A(SI_15_), .B(keyinput_17), .ZN(n9484) );
  XNOR2_X1 U10491 ( .A(n9689), .B(keyinput_18), .ZN(n9483) );
  XOR2_X1 U10492 ( .A(SI_13_), .B(keyinput_19), .Z(n9482) );
  AOI211_X1 U10493 ( .C1(n9485), .C2(n9484), .A(n9483), .B(n9482), .ZN(n9488)
         );
  XNOR2_X1 U10494 ( .A(SI_12_), .B(keyinput_20), .ZN(n9487) );
  XNOR2_X1 U10495 ( .A(n9694), .B(keyinput_21), .ZN(n9486) );
  OAI21_X1 U10496 ( .B1(n9488), .B2(n9487), .A(n9486), .ZN(n9492) );
  XNOR2_X1 U10497 ( .A(n9698), .B(keyinput_22), .ZN(n9491) );
  XNOR2_X1 U10498 ( .A(n9699), .B(keyinput_23), .ZN(n9490) );
  XNOR2_X1 U10499 ( .A(SI_8_), .B(keyinput_24), .ZN(n9489) );
  AOI211_X1 U10500 ( .C1(n9492), .C2(n9491), .A(n9490), .B(n9489), .ZN(n9496)
         );
  XNOR2_X1 U10501 ( .A(n9493), .B(keyinput_26), .ZN(n9495) );
  XNOR2_X1 U10502 ( .A(SI_7_), .B(keyinput_25), .ZN(n9494) );
  NOR3_X1 U10503 ( .A1(n9496), .A2(n9495), .A3(n9494), .ZN(n9501) );
  XNOR2_X1 U10504 ( .A(n9497), .B(keyinput_27), .ZN(n9500) );
  XNOR2_X1 U10505 ( .A(n9709), .B(keyinput_29), .ZN(n9499) );
  XNOR2_X1 U10506 ( .A(SI_4_), .B(keyinput_28), .ZN(n9498) );
  OAI211_X1 U10507 ( .C1(n9501), .C2(n9500), .A(n9499), .B(n9498), .ZN(n9508)
         );
  XNOR2_X1 U10508 ( .A(n9502), .B(keyinput_30), .ZN(n9507) );
  XNOR2_X1 U10509 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n9505) );
  XNOR2_X1 U10510 ( .A(SI_0_), .B(keyinput_32), .ZN(n9504) );
  XNOR2_X1 U10511 ( .A(SI_1_), .B(keyinput_31), .ZN(n9503) );
  NAND3_X1 U10512 ( .A1(n9505), .A2(n9504), .A3(n9503), .ZN(n9506) );
  AOI21_X1 U10513 ( .B1(n9508), .B2(n9507), .A(n9506), .ZN(n9514) );
  XNOR2_X1 U10514 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_34), .ZN(n9513) );
  XOR2_X1 U10515 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .Z(n9511) );
  XOR2_X1 U10516 ( .A(keyinput_37), .B(P2_REG3_REG_14__SCAN_IN), .Z(n9510) );
  XOR2_X1 U10517 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .Z(n9509) );
  NOR3_X1 U10518 ( .A1(n9511), .A2(n9510), .A3(n9509), .ZN(n9512) );
  OAI21_X1 U10519 ( .B1(n9514), .B2(n9513), .A(n9512), .ZN(n9517) );
  XOR2_X1 U10520 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .Z(n9516) );
  XNOR2_X1 U10521 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n9515)
         );
  AOI21_X1 U10522 ( .B1(n9517), .B2(n9516), .A(n9515), .ZN(n9521) );
  XNOR2_X1 U10523 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n9520) );
  XNOR2_X1 U10524 ( .A(n9518), .B(keyinput_41), .ZN(n9519) );
  OAI21_X1 U10525 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(n9525) );
  XNOR2_X1 U10526 ( .A(n9522), .B(keyinput_42), .ZN(n9524) );
  XNOR2_X1 U10527 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_43), .ZN(n9523) );
  AOI21_X1 U10528 ( .B1(n9525), .B2(n9524), .A(n9523), .ZN(n9534) );
  XNOR2_X1 U10529 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n9533)
         );
  XNOR2_X1 U10530 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n9532)
         );
  INV_X1 U10531 ( .A(keyinput_44), .ZN(n9526) );
  XNOR2_X1 U10532 ( .A(n9526), .B(P2_REG3_REG_1__SCAN_IN), .ZN(n9530) );
  XNOR2_X1 U10533 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n9529)
         );
  XNOR2_X1 U10534 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n9528) );
  XNOR2_X1 U10535 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_48), .ZN(n9527)
         );
  NAND4_X1 U10536 ( .A1(n9530), .A2(n9529), .A3(n9528), .A4(n9527), .ZN(n9531)
         );
  NOR4_X1 U10537 ( .A1(n9534), .A2(n9533), .A3(n9532), .A4(n9531), .ZN(n9548)
         );
  XNOR2_X1 U10538 ( .A(keyinput_50), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n9547)
         );
  XOR2_X1 U10539 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_56), .Z(n9539) );
  XOR2_X1 U10540 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_57), .Z(n9538) );
  XOR2_X1 U10541 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n9537) );
  XNOR2_X1 U10542 ( .A(n9535), .B(keyinput_55), .ZN(n9536) );
  NOR4_X1 U10543 ( .A1(n9539), .A2(n9538), .A3(n9537), .A4(n9536), .ZN(n9546)
         );
  XOR2_X1 U10544 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .Z(n9544) );
  XNOR2_X1 U10545 ( .A(n9744), .B(keyinput_53), .ZN(n9543) );
  XNOR2_X1 U10546 ( .A(n9540), .B(keyinput_51), .ZN(n9542) );
  XNOR2_X1 U10547 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n9541)
         );
  NOR4_X1 U10548 ( .A1(n9544), .A2(n9543), .A3(n9542), .A4(n9541), .ZN(n9545)
         );
  OAI211_X1 U10549 ( .C1(n9548), .C2(n9547), .A(n9546), .B(n9545), .ZN(n9551)
         );
  XNOR2_X1 U10550 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n9550) );
  XNOR2_X1 U10551 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n9549)
         );
  NAND3_X1 U10552 ( .A1(n9551), .A2(n9550), .A3(n9549), .ZN(n9565) );
  XNOR2_X1 U10553 ( .A(n9762), .B(keyinput_62), .ZN(n9561) );
  INV_X1 U10554 ( .A(P2_B_REG_SCAN_IN), .ZN(n9763) );
  OAI22_X1 U10555 ( .A1(keyinput_64), .A2(n9763), .B1(n9764), .B2(keyinput_66), 
        .ZN(n9560) );
  INV_X1 U10556 ( .A(keyinput_67), .ZN(n9552) );
  NAND2_X1 U10557 ( .A1(n9552), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9557) );
  AOI22_X1 U10558 ( .A1(n9763), .A2(keyinput_64), .B1(n9760), .B2(keyinput_67), 
        .ZN(n9555) );
  AOI22_X1 U10559 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_65), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_63), .ZN(n9554) );
  AOI22_X1 U10560 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_61), .B1(n9764), 
        .B2(keyinput_66), .ZN(n9553) );
  AND3_X1 U10561 ( .A1(n9555), .A2(n9554), .A3(n9553), .ZN(n9556) );
  OAI211_X1 U10562 ( .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_61), .A(n9557), 
        .B(n9556), .ZN(n9559) );
  OAI22_X1 U10563 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_65), .B1(
        keyinput_63), .B2(P2_REG3_REG_15__SCAN_IN), .ZN(n9558) );
  NOR4_X1 U10564 ( .A1(n9561), .A2(n9560), .A3(n9559), .A4(n9558), .ZN(n9564)
         );
  XNOR2_X1 U10565 ( .A(n9774), .B(keyinput_69), .ZN(n9563) );
  XNOR2_X1 U10566 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .ZN(n9562)
         );
  AOI211_X1 U10567 ( .C1(n9565), .C2(n9564), .A(n9563), .B(n9562), .ZN(n9568)
         );
  XNOR2_X1 U10568 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .ZN(n9567)
         );
  XNOR2_X1 U10569 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n9566)
         );
  OAI21_X1 U10570 ( .B1(n9568), .B2(n9567), .A(n9566), .ZN(n9572) );
  XNOR2_X1 U10571 ( .A(n9569), .B(keyinput_72), .ZN(n9571) );
  XNOR2_X1 U10572 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n9570)
         );
  NAND3_X1 U10573 ( .A1(n9572), .A2(n9571), .A3(n9570), .ZN(n9579) );
  XOR2_X1 U10574 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .Z(n9578) );
  XNOR2_X1 U10575 ( .A(n9788), .B(keyinput_76), .ZN(n9576) );
  XNOR2_X1 U10576 ( .A(n9573), .B(keyinput_77), .ZN(n9575) );
  XNOR2_X1 U10577 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .ZN(n9574)
         );
  NAND3_X1 U10578 ( .A1(n9576), .A2(n9575), .A3(n9574), .ZN(n9577) );
  AOI21_X1 U10579 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9582) );
  XNOR2_X1 U10580 ( .A(n9793), .B(keyinput_79), .ZN(n9581) );
  XNOR2_X1 U10581 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .ZN(n9580)
         );
  NOR3_X1 U10582 ( .A1(n9582), .A2(n9581), .A3(n9580), .ZN(n9587) );
  XNOR2_X1 U10583 ( .A(n9797), .B(keyinput_80), .ZN(n9586) );
  XOR2_X1 U10584 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .Z(n9585) );
  XNOR2_X1 U10585 ( .A(n9583), .B(keyinput_82), .ZN(n9584) );
  OAI211_X1 U10586 ( .C1(n9587), .C2(n9586), .A(n9585), .B(n9584), .ZN(n9590)
         );
  XOR2_X1 U10587 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .Z(n9589) );
  XNOR2_X1 U10588 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n9588)
         );
  NAND3_X1 U10589 ( .A1(n9590), .A2(n9589), .A3(n9588), .ZN(n9595) );
  XNOR2_X1 U10590 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n9594)
         );
  XNOR2_X1 U10591 ( .A(n9591), .B(keyinput_87), .ZN(n9593) );
  XOR2_X1 U10592 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .Z(n9592) );
  AOI211_X1 U10593 ( .C1(n9595), .C2(n9594), .A(n9593), .B(n9592), .ZN(n9602)
         );
  XNOR2_X1 U10594 ( .A(n9810), .B(keyinput_88), .ZN(n9601) );
  XOR2_X1 U10595 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_92), .Z(n9599) );
  XNOR2_X1 U10596 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n9598)
         );
  XNOR2_X1 U10597 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_91), .ZN(n9597) );
  XNOR2_X1 U10598 ( .A(n10752), .B(keyinput_90), .ZN(n9596) );
  NOR4_X1 U10599 ( .A1(n9599), .A2(n9598), .A3(n9597), .A4(n9596), .ZN(n9600)
         );
  OAI21_X1 U10600 ( .B1(n9602), .B2(n9601), .A(n9600), .ZN(n9605) );
  XNOR2_X1 U10601 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n9604) );
  XNOR2_X1 U10602 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_94), .ZN(n9603) );
  NAND3_X1 U10603 ( .A1(n9605), .A2(n9604), .A3(n9603), .ZN(n9609) );
  XOR2_X1 U10604 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_97), .Z(n9608) );
  XOR2_X1 U10605 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_95), .Z(n9607) );
  XNOR2_X1 U10606 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_96), .ZN(n9606) );
  NAND4_X1 U10607 ( .A1(n9609), .A2(n9608), .A3(n9607), .A4(n9606), .ZN(n9613)
         );
  XOR2_X1 U10608 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_100), .Z(n9612) );
  XOR2_X1 U10609 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_99), .Z(n9611) );
  XNOR2_X1 U10610 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_98), .ZN(n9610) );
  NAND4_X1 U10611 ( .A1(n9613), .A2(n9612), .A3(n9611), .A4(n9610), .ZN(n9617)
         );
  XOR2_X1 U10612 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_101), .Z(n9616) );
  XOR2_X1 U10613 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_103), .Z(n9615) );
  XNOR2_X1 U10614 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_102), .ZN(n9614) );
  AOI211_X1 U10615 ( .C1(n9617), .C2(n9616), .A(n9615), .B(n9614), .ZN(n9624)
         );
  XOR2_X1 U10616 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_108), .Z(n9623) );
  XNOR2_X1 U10617 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_105), .ZN(n9622) );
  XOR2_X1 U10618 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_107), .Z(n9620) );
  XNOR2_X1 U10619 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_104), .ZN(n9619) );
  XNOR2_X1 U10620 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_106), .ZN(n9618) );
  NAND3_X1 U10621 ( .A1(n9620), .A2(n9619), .A3(n9618), .ZN(n9621) );
  NOR4_X1 U10622 ( .A1(n9624), .A2(n9623), .A3(n9622), .A4(n9621), .ZN(n9631)
         );
  XOR2_X1 U10623 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_109), .Z(n9630) );
  XOR2_X1 U10624 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_112), .Z(n9629) );
  OAI22_X1 U10625 ( .A1(n9627), .A2(keyinput_111), .B1(keyinput_110), .B2(
        P1_IR_REG_20__SCAN_IN), .ZN(n9626) );
  AND2_X1 U10626 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_110), .ZN(n9625)
         );
  AOI211_X1 U10627 ( .C1(keyinput_111), .C2(n9627), .A(n9626), .B(n9625), .ZN(
        n9628) );
  OAI211_X1 U10628 ( .C1(n9631), .C2(n9630), .A(n9629), .B(n9628), .ZN(n9634)
         );
  XOR2_X1 U10629 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_114), .Z(n9633) );
  XNOR2_X1 U10630 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_113), .ZN(n9632) );
  NAND3_X1 U10631 ( .A1(n9634), .A2(n9633), .A3(n9632), .ZN(n9637) );
  XOR2_X1 U10632 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_115), .Z(n9636) );
  XNOR2_X1 U10633 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_116), .ZN(n9635) );
  AOI21_X1 U10634 ( .B1(n9637), .B2(n9636), .A(n9635), .ZN(n9641) );
  XOR2_X1 U10635 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_117), .Z(n9640) );
  XNOR2_X1 U10636 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_119), .ZN(n9639) );
  XNOR2_X1 U10637 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_118), .ZN(n9638) );
  OAI211_X1 U10638 ( .C1(n9641), .C2(n9640), .A(n9639), .B(n9638), .ZN(n9644)
         );
  XOR2_X1 U10639 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_120), .Z(n9643) );
  XNOR2_X1 U10640 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_121), .ZN(n9642) );
  AOI21_X1 U10641 ( .B1(n9644), .B2(n9643), .A(n9642), .ZN(n9648) );
  XNOR2_X1 U10642 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_122), .ZN(n9647) );
  XNOR2_X1 U10643 ( .A(keyinput_124), .B(P1_D_REG_2__SCAN_IN), .ZN(n9646) );
  XNOR2_X1 U10644 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_123), .ZN(n9645) );
  OAI211_X1 U10645 ( .C1(n9648), .C2(n9647), .A(n9646), .B(n9645), .ZN(n9651)
         );
  INV_X1 U10646 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10668) );
  XNOR2_X1 U10647 ( .A(n10668), .B(keyinput_125), .ZN(n9650) );
  INV_X1 U10648 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10669) );
  XNOR2_X1 U10649 ( .A(n10669), .B(keyinput_126), .ZN(n9649) );
  AOI21_X1 U10650 ( .B1(n9651), .B2(n9650), .A(n9649), .ZN(n9869) );
  XOR2_X1 U10651 ( .A(keyinput_255), .B(keyinput_127), .Z(n9868) );
  XNOR2_X1 U10652 ( .A(n9652), .B(keyinput_144), .ZN(n9654) );
  XNOR2_X1 U10653 ( .A(SI_17_), .B(keyinput_143), .ZN(n9653) );
  NAND2_X1 U10654 ( .A1(n9654), .A2(n9653), .ZN(n9683) );
  INV_X1 U10655 ( .A(n9683), .ZN(n9688) );
  XNOR2_X1 U10656 ( .A(n9655), .B(keyinput_142), .ZN(n9687) );
  XNOR2_X1 U10657 ( .A(n9656), .B(keyinput_145), .ZN(n9686) );
  XOR2_X1 U10658 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n9660) );
  XNOR2_X1 U10659 ( .A(n9657), .B(keyinput_129), .ZN(n9659) );
  XNOR2_X1 U10660 ( .A(SI_30_), .B(keyinput_130), .ZN(n9658) );
  NAND3_X1 U10661 ( .A1(n9660), .A2(n9659), .A3(n9658), .ZN(n9665) );
  XNOR2_X1 U10662 ( .A(n9661), .B(keyinput_131), .ZN(n9664) );
  XNOR2_X1 U10663 ( .A(n9662), .B(keyinput_132), .ZN(n9663) );
  AOI21_X1 U10664 ( .B1(n9665), .B2(n9664), .A(n9663), .ZN(n9673) );
  XNOR2_X1 U10665 ( .A(SI_27_), .B(keyinput_133), .ZN(n9672) );
  XNOR2_X1 U10666 ( .A(n9666), .B(keyinput_134), .ZN(n9670) );
  XNOR2_X1 U10667 ( .A(n9667), .B(keyinput_136), .ZN(n9669) );
  XNOR2_X1 U10668 ( .A(SI_25_), .B(keyinput_135), .ZN(n9668) );
  NOR3_X1 U10669 ( .A1(n9670), .A2(n9669), .A3(n9668), .ZN(n9671) );
  OAI21_X1 U10670 ( .B1(n9673), .B2(n9672), .A(n9671), .ZN(n9681) );
  XNOR2_X1 U10671 ( .A(n9674), .B(keyinput_137), .ZN(n9680) );
  XOR2_X1 U10672 ( .A(SI_22_), .B(keyinput_138), .Z(n9678) );
  XNOR2_X1 U10673 ( .A(n9675), .B(keyinput_140), .ZN(n9677) );
  XNOR2_X1 U10674 ( .A(SI_21_), .B(keyinput_139), .ZN(n9676) );
  NAND3_X1 U10675 ( .A1(n9678), .A2(n9677), .A3(n9676), .ZN(n9679) );
  AOI21_X1 U10676 ( .B1(n9681), .B2(n9680), .A(n9679), .ZN(n9684) );
  XNOR2_X1 U10677 ( .A(SI_19_), .B(keyinput_141), .ZN(n9682) );
  NOR3_X1 U10678 ( .A1(n9684), .A2(n9683), .A3(n9682), .ZN(n9685) );
  AOI211_X1 U10679 ( .C1(n9688), .C2(n9687), .A(n9686), .B(n9685), .ZN(n9692)
         );
  XNOR2_X1 U10680 ( .A(n9689), .B(keyinput_146), .ZN(n9691) );
  XOR2_X1 U10681 ( .A(SI_13_), .B(keyinput_147), .Z(n9690) );
  NOR3_X1 U10682 ( .A1(n9692), .A2(n9691), .A3(n9690), .ZN(n9697) );
  XNOR2_X1 U10683 ( .A(n9693), .B(keyinput_148), .ZN(n9696) );
  XNOR2_X1 U10684 ( .A(n9694), .B(keyinput_149), .ZN(n9695) );
  OAI21_X1 U10685 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(n9704) );
  XNOR2_X1 U10686 ( .A(n9698), .B(keyinput_150), .ZN(n9703) );
  XNOR2_X1 U10687 ( .A(n9699), .B(keyinput_151), .ZN(n9702) );
  XNOR2_X1 U10688 ( .A(n9700), .B(keyinput_152), .ZN(n9701) );
  AOI211_X1 U10689 ( .C1(n9704), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9707)
         );
  XNOR2_X1 U10690 ( .A(SI_7_), .B(keyinput_153), .ZN(n9706) );
  XNOR2_X1 U10691 ( .A(SI_6_), .B(keyinput_154), .ZN(n9705) );
  NOR3_X1 U10692 ( .A1(n9707), .A2(n9706), .A3(n9705), .ZN(n9713) );
  XNOR2_X1 U10693 ( .A(SI_5_), .B(keyinput_155), .ZN(n9712) );
  XNOR2_X1 U10694 ( .A(n9708), .B(keyinput_156), .ZN(n9711) );
  XNOR2_X1 U10695 ( .A(n9709), .B(keyinput_157), .ZN(n9710) );
  OAI211_X1 U10696 ( .C1(n9713), .C2(n9712), .A(n9711), .B(n9710), .ZN(n9719)
         );
  XNOR2_X1 U10697 ( .A(SI_2_), .B(keyinput_158), .ZN(n9718) );
  XNOR2_X1 U10698 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_161), .ZN(n9717) );
  XNOR2_X1 U10699 ( .A(SI_0_), .B(keyinput_160), .ZN(n9715) );
  XNOR2_X1 U10700 ( .A(SI_1_), .B(keyinput_159), .ZN(n9714) );
  NAND2_X1 U10701 ( .A1(n9715), .A2(n9714), .ZN(n9716) );
  AOI211_X1 U10702 ( .C1(n9719), .C2(n9718), .A(n9717), .B(n9716), .ZN(n9725)
         );
  XNOR2_X1 U10703 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_162), .ZN(n9724) );
  XOR2_X1 U10704 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_163), .Z(n9722) );
  XOR2_X1 U10705 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .Z(n9721) );
  XNOR2_X1 U10706 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n9720)
         );
  NOR3_X1 U10707 ( .A1(n9722), .A2(n9721), .A3(n9720), .ZN(n9723) );
  OAI21_X1 U10708 ( .B1(n9725), .B2(n9724), .A(n9723), .ZN(n9728) );
  XNOR2_X1 U10709 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n9727)
         );
  XOR2_X1 U10710 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .Z(n9726) );
  AOI21_X1 U10711 ( .B1(n9728), .B2(n9727), .A(n9726), .ZN(n9731) );
  XOR2_X1 U10712 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .Z(n9730) );
  XNOR2_X1 U10713 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n9729)
         );
  OAI21_X1 U10714 ( .B1(n9731), .B2(n9730), .A(n9729), .ZN(n9734) );
  XNOR2_X1 U10715 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n9733)
         );
  XNOR2_X1 U10716 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n9732)
         );
  AOI21_X1 U10717 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(n9743) );
  XNOR2_X1 U10718 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n9742)
         );
  XNOR2_X1 U10719 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n9741)
         );
  XOR2_X1 U10720 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .Z(n9739) );
  XOR2_X1 U10721 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_174), .Z(n9738) );
  XNOR2_X1 U10722 ( .A(n9735), .B(keyinput_175), .ZN(n9737) );
  XNOR2_X1 U10723 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_177), .ZN(n9736)
         );
  NAND4_X1 U10724 ( .A1(n9739), .A2(n9738), .A3(n9737), .A4(n9736), .ZN(n9740)
         );
  NOR4_X1 U10725 ( .A1(n9743), .A2(n9742), .A3(n9741), .A4(n9740), .ZN(n9756)
         );
  XOR2_X1 U10726 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .Z(n9755) );
  XOR2_X1 U10727 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .Z(n9748) );
  XOR2_X1 U10728 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_184), .Z(n9747) );
  XOR2_X1 U10729 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .Z(n9746) );
  XNOR2_X1 U10730 ( .A(n9744), .B(keyinput_181), .ZN(n9745) );
  NOR4_X1 U10731 ( .A1(n9748), .A2(n9747), .A3(n9746), .A4(n9745), .ZN(n9754)
         );
  XOR2_X1 U10732 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_186), .Z(n9752) );
  XNOR2_X1 U10733 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_185), .ZN(n9751)
         );
  XNOR2_X1 U10734 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_179), .ZN(n9750)
         );
  XNOR2_X1 U10735 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_183), .ZN(n9749)
         );
  NOR4_X1 U10736 ( .A1(n9752), .A2(n9751), .A3(n9750), .A4(n9749), .ZN(n9753)
         );
  OAI211_X1 U10737 ( .C1(n9756), .C2(n9755), .A(n9754), .B(n9753), .ZN(n9759)
         );
  XOR2_X1 U10738 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n9758) );
  XNOR2_X1 U10739 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n9757)
         );
  NAND3_X1 U10740 ( .A1(n9759), .A2(n9758), .A3(n9757), .ZN(n9778) );
  XNOR2_X1 U10741 ( .A(n9760), .B(keyinput_195), .ZN(n9773) );
  OAI22_X1 U10742 ( .A1(keyinput_194), .A2(n9764), .B1(n9763), .B2(
        keyinput_192), .ZN(n9772) );
  INV_X1 U10743 ( .A(keyinput_190), .ZN(n9761) );
  NAND2_X1 U10744 ( .A1(n9761), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9769) );
  AOI22_X1 U10745 ( .A1(n9763), .A2(keyinput_192), .B1(n9762), .B2(
        keyinput_190), .ZN(n9767) );
  AOI22_X1 U10746 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_189), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_191), .ZN(n9766) );
  AOI22_X1 U10747 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_193), .B1(
        n9764), .B2(keyinput_194), .ZN(n9765) );
  AND3_X1 U10748 ( .A1(n9767), .A2(n9766), .A3(n9765), .ZN(n9768) );
  OAI211_X1 U10749 ( .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_189), .A(n9769), 
        .B(n9768), .ZN(n9771) );
  OAI22_X1 U10750 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_193), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_191), .ZN(n9770) );
  NOR4_X1 U10751 ( .A1(n9773), .A2(n9772), .A3(n9771), .A4(n9770), .ZN(n9777)
         );
  XNOR2_X1 U10752 ( .A(n9774), .B(keyinput_197), .ZN(n9776) );
  XNOR2_X1 U10753 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n9775)
         );
  AOI211_X1 U10754 ( .C1(n9778), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9781)
         );
  XNOR2_X1 U10755 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .ZN(n9780)
         );
  XOR2_X1 U10756 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .Z(n9779)
         );
  OAI21_X1 U10757 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9785) );
  XNOR2_X1 U10758 ( .A(n9782), .B(keyinput_201), .ZN(n9784) );
  XNOR2_X1 U10759 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .ZN(n9783)
         );
  NAND3_X1 U10760 ( .A1(n9785), .A2(n9784), .A3(n9783), .ZN(n9787) );
  XNOR2_X1 U10761 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n9786)
         );
  NAND2_X1 U10762 ( .A1(n9787), .A2(n9786), .ZN(n9792) );
  XNOR2_X1 U10763 ( .A(n9788), .B(keyinput_204), .ZN(n9791) );
  XOR2_X1 U10764 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n9790)
         );
  XNOR2_X1 U10765 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .ZN(n9789)
         );
  NAND4_X1 U10766 ( .A1(n9792), .A2(n9791), .A3(n9790), .A4(n9789), .ZN(n9796)
         );
  XNOR2_X1 U10767 ( .A(n9793), .B(keyinput_207), .ZN(n9795) );
  XOR2_X1 U10768 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .Z(n9794)
         );
  NAND3_X1 U10769 ( .A1(n9796), .A2(n9795), .A3(n9794), .ZN(n9801) );
  XNOR2_X1 U10770 ( .A(n9797), .B(keyinput_208), .ZN(n9800) );
  XNOR2_X1 U10771 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n9799)
         );
  XNOR2_X1 U10772 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .ZN(n9798)
         );
  AOI211_X1 U10773 ( .C1(n9801), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9804)
         );
  XNOR2_X1 U10774 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .ZN(n9803)
         );
  XNOR2_X1 U10775 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .ZN(n9802)
         );
  NOR3_X1 U10776 ( .A1(n9804), .A2(n9803), .A3(n9802), .ZN(n9809) );
  XNOR2_X1 U10777 ( .A(n9805), .B(keyinput_213), .ZN(n9808) );
  XNOR2_X1 U10778 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .ZN(n9807)
         );
  XNOR2_X1 U10779 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n9806)
         );
  OAI211_X1 U10780 ( .C1(n9809), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9817)
         );
  XNOR2_X1 U10781 ( .A(n9810), .B(keyinput_216), .ZN(n9816) );
  XOR2_X1 U10782 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_220), .Z(n9814) );
  XOR2_X1 U10783 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .Z(n9813) );
  XOR2_X1 U10784 ( .A(n10752), .B(keyinput_218), .Z(n9812) );
  XNOR2_X1 U10785 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_219), .ZN(n9811) );
  NAND4_X1 U10786 ( .A1(n9814), .A2(n9813), .A3(n9812), .A4(n9811), .ZN(n9815)
         );
  AOI21_X1 U10787 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9820) );
  XOR2_X1 U10788 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_222), .Z(n9819) );
  XOR2_X1 U10789 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_221), .Z(n9818) );
  NOR3_X1 U10790 ( .A1(n9820), .A2(n9819), .A3(n9818), .ZN(n9824) );
  XOR2_X1 U10791 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_225), .Z(n9823) );
  XOR2_X1 U10792 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_223), .Z(n9822) );
  XOR2_X1 U10793 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_224), .Z(n9821) );
  NOR4_X1 U10794 ( .A1(n9824), .A2(n9823), .A3(n9822), .A4(n9821), .ZN(n9828)
         );
  XOR2_X1 U10795 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_228), .Z(n9827) );
  XNOR2_X1 U10796 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_226), .ZN(n9826) );
  XNOR2_X1 U10797 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_227), .ZN(n9825) );
  NOR4_X1 U10798 ( .A1(n9828), .A2(n9827), .A3(n9826), .A4(n9825), .ZN(n9832)
         );
  XOR2_X1 U10799 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_229), .Z(n9831) );
  XNOR2_X1 U10800 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_231), .ZN(n9830) );
  XNOR2_X1 U10801 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_230), .ZN(n9829) );
  OAI211_X1 U10802 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9839)
         );
  XOR2_X1 U10803 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_234), .Z(n9835) );
  XOR2_X1 U10804 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_233), .Z(n9834) );
  XNOR2_X1 U10805 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_232), .ZN(n9833) );
  NOR3_X1 U10806 ( .A1(n9835), .A2(n9834), .A3(n9833), .ZN(n9838) );
  XNOR2_X1 U10807 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_235), .ZN(n9837) );
  XNOR2_X1 U10808 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_236), .ZN(n9836) );
  NAND4_X1 U10809 ( .A1(n9839), .A2(n9838), .A3(n9837), .A4(n9836), .ZN(n9845)
         );
  XOR2_X1 U10810 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_237), .Z(n9844) );
  XOR2_X1 U10811 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_240), .Z(n9842) );
  XNOR2_X1 U10812 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_239), .ZN(n9841) );
  XNOR2_X1 U10813 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_238), .ZN(n9840) );
  NAND3_X1 U10814 ( .A1(n9842), .A2(n9841), .A3(n9840), .ZN(n9843) );
  AOI21_X1 U10815 ( .B1(n9845), .B2(n9844), .A(n9843), .ZN(n9848) );
  XOR2_X1 U10816 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_241), .Z(n9847) );
  XNOR2_X1 U10817 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_242), .ZN(n9846) );
  NOR3_X1 U10818 ( .A1(n9848), .A2(n9847), .A3(n9846), .ZN(n9851) );
  XNOR2_X1 U10819 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_243), .ZN(n9850) );
  XOR2_X1 U10820 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_244), .Z(n9849) );
  OAI21_X1 U10821 ( .B1(n9851), .B2(n9850), .A(n9849), .ZN(n9855) );
  XOR2_X1 U10822 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_245), .Z(n9854) );
  XNOR2_X1 U10823 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_247), .ZN(n9853) );
  XNOR2_X1 U10824 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_246), .ZN(n9852) );
  AOI211_X1 U10825 ( .C1(n9855), .C2(n9854), .A(n9853), .B(n9852), .ZN(n9858)
         );
  XOR2_X1 U10826 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_248), .Z(n9857) );
  XOR2_X1 U10827 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_249), .Z(n9856) );
  OAI21_X1 U10828 ( .B1(n9858), .B2(n9857), .A(n9856), .ZN(n9862) );
  XOR2_X1 U10829 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_250), .Z(n9861) );
  INV_X1 U10830 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10667) );
  XNOR2_X1 U10831 ( .A(n10667), .B(keyinput_252), .ZN(n9860) );
  XOR2_X1 U10832 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_251), .Z(n9859) );
  AOI211_X1 U10833 ( .C1(n9862), .C2(n9861), .A(n9860), .B(n9859), .ZN(n9865)
         );
  XNOR2_X1 U10834 ( .A(n10668), .B(keyinput_253), .ZN(n9864) );
  XNOR2_X1 U10835 ( .A(n10669), .B(keyinput_254), .ZN(n9863) );
  OAI21_X1 U10836 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(n9867) );
  XNOR2_X1 U10837 ( .A(keyinput_255), .B(P1_D_REG_5__SCAN_IN), .ZN(n9866) );
  OAI211_X1 U10838 ( .C1(n9869), .C2(n9868), .A(n9867), .B(n9866), .ZN(n9870)
         );
  XNOR2_X1 U10839 ( .A(n9871), .B(n9870), .ZN(P2_U3205) );
  OAI211_X1 U10840 ( .C1(n9873), .C2(n9883), .A(n9872), .B(n10935), .ZN(n9877)
         );
  AOI22_X1 U10841 ( .A1(n9903), .A2(n9875), .B1(n10944), .B2(n9874), .ZN(n9876) );
  OAI22_X1 U10842 ( .A1(n11048), .A2(n9879), .B1(n9878), .B2(n10950), .ZN(
        n9885) );
  INV_X1 U10843 ( .A(n9880), .ZN(n9881) );
  AOI21_X1 U10844 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(n9999) );
  NOR2_X1 U10845 ( .A1(n9999), .A2(n9954), .ZN(n9884) );
  AOI211_X1 U10846 ( .C1(n11043), .C2(n9996), .A(n9885), .B(n9884), .ZN(n9886)
         );
  OAI21_X1 U10847 ( .B1(n10981), .B2(n9998), .A(n9886), .ZN(P2_U3206) );
  OAI22_X1 U10848 ( .A1(n11048), .A2(n9890), .B1(n9889), .B2(n10950), .ZN(
        n9894) );
  OAI21_X1 U10849 ( .B1(n9892), .B2(n5431), .A(n9891), .ZN(n10003) );
  NOR2_X1 U10850 ( .A1(n10003), .A2(n9954), .ZN(n9893) );
  AOI211_X1 U10851 ( .C1(n11043), .C2(n10000), .A(n9894), .B(n9893), .ZN(n9895) );
  OAI21_X1 U10852 ( .B1(n10002), .B2(n10981), .A(n9895), .ZN(P2_U3207) );
  NAND2_X1 U10853 ( .A1(n9896), .A2(n5436), .ZN(n9897) );
  NAND2_X1 U10854 ( .A1(n9898), .A2(n9897), .ZN(n10005) );
  XNOR2_X1 U10855 ( .A(n9900), .B(n9899), .ZN(n9901) );
  NAND2_X1 U10856 ( .A1(n9901), .A2(n10935), .ZN(n9905) );
  AOI22_X1 U10857 ( .A1(n9903), .A2(n9902), .B1(n9961), .B2(n9923), .ZN(n9904)
         );
  NAND2_X1 U10858 ( .A1(n9905), .A2(n9904), .ZN(n10007) );
  INV_X1 U10859 ( .A(n9906), .ZN(n10004) );
  OAI22_X1 U10860 ( .A1(n10004), .A2(n10974), .B1(n9907), .B2(n10950), .ZN(
        n9908) );
  OAI21_X1 U10861 ( .B1(n10007), .B2(n9908), .A(n11046), .ZN(n9910) );
  NAND2_X1 U10862 ( .A1(n10981), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9909) );
  OAI211_X1 U10863 ( .C1(n10005), .C2(n9954), .A(n9910), .B(n9909), .ZN(
        P2_U3208) );
  XNOR2_X1 U10864 ( .A(n9911), .B(n9913), .ZN(n10009) );
  INV_X1 U10865 ( .A(n10009), .ZN(n9921) );
  INV_X1 U10866 ( .A(n10008), .ZN(n9916) );
  XOR2_X1 U10867 ( .A(n9912), .B(n9913), .Z(n9915) );
  AOI222_X1 U10868 ( .A1(n10935), .A2(n9915), .B1(n9914), .B2(n10944), .C1(
        n9934), .C2(n9961), .ZN(n10011) );
  OAI21_X1 U10869 ( .B1(n9916), .B2(n10974), .A(n10011), .ZN(n9917) );
  NAND2_X1 U10870 ( .A1(n9917), .A2(n11046), .ZN(n9920) );
  AOI22_X1 U10871 ( .A1(n10981), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n11041), 
        .B2(n9918), .ZN(n9919) );
  OAI211_X1 U10872 ( .C1(n9921), .C2(n9954), .A(n9920), .B(n9919), .ZN(
        P2_U3209) );
  XNOR2_X1 U10873 ( .A(n9922), .B(n9925), .ZN(n9924) );
  AOI222_X1 U10874 ( .A1(n10935), .A2(n9924), .B1(n9923), .B2(n10944), .C1(
        n9947), .C2(n9961), .ZN(n10015) );
  XNOR2_X1 U10875 ( .A(n9926), .B(n9925), .ZN(n10013) );
  AOI22_X1 U10876 ( .A1(n10981), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n11041), 
        .B2(n9927), .ZN(n9928) );
  OAI21_X1 U10877 ( .B1(n9929), .B2(n9984), .A(n9928), .ZN(n9930) );
  AOI21_X1 U10878 ( .B1(n10013), .B2(n9987), .A(n9930), .ZN(n9931) );
  OAI21_X1 U10879 ( .B1(n10015), .B2(n10981), .A(n9931), .ZN(P2_U3210) );
  XNOR2_X1 U10880 ( .A(n9933), .B(n9932), .ZN(n9935) );
  AOI222_X1 U10881 ( .A1(n10935), .A2(n9935), .B1(n9934), .B2(n10944), .C1(
        n9963), .C2(n9961), .ZN(n10018) );
  OAI22_X1 U10882 ( .A1(n11048), .A2(n9937), .B1(n9936), .B2(n10950), .ZN(
        n9942) );
  OAI21_X1 U10883 ( .B1(n9940), .B2(n9939), .A(n9938), .ZN(n10019) );
  NOR2_X1 U10884 ( .A1(n10019), .A2(n9954), .ZN(n9941) );
  AOI211_X1 U10885 ( .C1(n11043), .C2(n10016), .A(n9942), .B(n9941), .ZN(n9943) );
  OAI21_X1 U10886 ( .B1(n10018), .B2(n10981), .A(n9943), .ZN(P2_U3211) );
  XNOR2_X1 U10887 ( .A(n9945), .B(n9944), .ZN(n9948) );
  AOI222_X1 U10888 ( .A1(n10935), .A2(n9948), .B1(n9947), .B2(n10944), .C1(
        n9946), .C2(n9961), .ZN(n10022) );
  OAI22_X1 U10889 ( .A1(n11048), .A2(n9950), .B1(n9949), .B2(n10950), .ZN(
        n9956) );
  OAI21_X1 U10890 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n10023) );
  NOR2_X1 U10891 ( .A1(n10023), .A2(n9954), .ZN(n9955) );
  AOI211_X1 U10892 ( .C1(n11043), .C2(n10020), .A(n9956), .B(n9955), .ZN(n9957) );
  OAI21_X1 U10893 ( .B1(n10022), .B2(n9958), .A(n9957), .ZN(P2_U3212) );
  OAI21_X1 U10894 ( .B1(n9960), .B2(n6664), .A(n9959), .ZN(n9964) );
  AOI222_X1 U10895 ( .A1(n10935), .A2(n9964), .B1(n9963), .B2(n10944), .C1(
        n9962), .C2(n9961), .ZN(n10027) );
  INV_X1 U10896 ( .A(n10027), .ZN(n9965) );
  AOI21_X1 U10897 ( .B1(n11041), .B2(n9966), .A(n9965), .ZN(n9975) );
  NAND2_X1 U10898 ( .A1(n9968), .A2(n9967), .ZN(n9970) );
  XNOR2_X1 U10899 ( .A(n9970), .B(n9969), .ZN(n10025) );
  OAI22_X1 U10900 ( .A1(n9972), .A2(n9984), .B1(n9971), .B2(n11046), .ZN(n9973) );
  AOI21_X1 U10901 ( .B1(n10025), .B2(n9987), .A(n9973), .ZN(n9974) );
  OAI21_X1 U10902 ( .B1(n9975), .B2(n10981), .A(n9974), .ZN(P2_U3213) );
  OAI211_X1 U10903 ( .C1(n9977), .C2(n9980), .A(n9976), .B(n10935), .ZN(n9979)
         );
  XOR2_X1 U10904 ( .A(n9981), .B(n9980), .Z(n10029) );
  AOI22_X1 U10905 ( .A1(n10981), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n11041), 
        .B2(n9982), .ZN(n9983) );
  OAI21_X1 U10906 ( .B1(n9985), .B2(n9984), .A(n9983), .ZN(n9986) );
  AOI21_X1 U10907 ( .B1(n10029), .B2(n9987), .A(n9986), .ZN(n9988) );
  OAI21_X1 U10908 ( .B1(n10981), .B2(n10030), .A(n9988), .ZN(P2_U3214) );
  OAI21_X1 U10909 ( .B1(n9989), .B2(n11127), .A(n9990), .ZN(n10037) );
  MUX2_X1 U10910 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n10037), .S(n11153), .Z(
        P2_U3490) );
  OAI21_X1 U10911 ( .B1(n9991), .B2(n11127), .A(n9990), .ZN(n10038) );
  MUX2_X1 U10912 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n10038), .S(n11153), .Z(
        P2_U3489) );
  NAND2_X1 U10913 ( .A1(n9992), .A2(n11151), .ZN(n9993) );
  OAI211_X1 U10914 ( .C1(n11146), .C2(n9995), .A(n9994), .B(n9993), .ZN(n10039) );
  MUX2_X1 U10915 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n10039), .S(n11153), .Z(
        P2_U3487) );
  NAND2_X1 U10916 ( .A1(n9996), .A2(n11151), .ZN(n9997) );
  OAI211_X1 U10917 ( .C1(n9999), .C2(n11146), .A(n9998), .B(n9997), .ZN(n10040) );
  MUX2_X1 U10918 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n10040), .S(n11153), .Z(
        P2_U3486) );
  NAND2_X1 U10919 ( .A1(n10000), .A2(n11151), .ZN(n10001) );
  OAI211_X1 U10920 ( .C1(n11146), .C2(n10003), .A(n10002), .B(n10001), .ZN(
        n10041) );
  MUX2_X1 U10921 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n10041), .S(n11153), .Z(
        P2_U3485) );
  OAI22_X1 U10922 ( .A1(n10005), .A2(n11146), .B1(n10004), .B2(n11127), .ZN(
        n10006) );
  MUX2_X1 U10923 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n10042), .S(n11153), .Z(
        P2_U3484) );
  AOI22_X1 U10924 ( .A1(n10009), .A2(n11132), .B1(n11151), .B2(n10008), .ZN(
        n10010) );
  NAND2_X1 U10925 ( .A1(n10011), .A2(n10010), .ZN(n10043) );
  MUX2_X1 U10926 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n10043), .S(n11153), .Z(
        P2_U3483) );
  AOI22_X1 U10927 ( .A1(n10013), .A2(n11132), .B1(n11151), .B2(n10012), .ZN(
        n10014) );
  NAND2_X1 U10928 ( .A1(n10015), .A2(n10014), .ZN(n10044) );
  MUX2_X1 U10929 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n10044), .S(n11153), .Z(
        P2_U3482) );
  NAND2_X1 U10930 ( .A1(n10016), .A2(n11151), .ZN(n10017) );
  OAI211_X1 U10931 ( .C1(n11146), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        n10045) );
  MUX2_X1 U10932 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n10045), .S(n11153), .Z(
        P2_U3481) );
  NAND2_X1 U10933 ( .A1(n10020), .A2(n11151), .ZN(n10021) );
  OAI211_X1 U10934 ( .C1(n11146), .C2(n10023), .A(n10022), .B(n10021), .ZN(
        n10046) );
  MUX2_X1 U10935 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n10046), .S(n11153), .Z(
        P2_U3480) );
  AOI22_X1 U10936 ( .A1(n10025), .A2(n11132), .B1(n11151), .B2(n10024), .ZN(
        n10026) );
  NAND2_X1 U10937 ( .A1(n10027), .A2(n10026), .ZN(n10047) );
  MUX2_X1 U10938 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n10047), .S(n11153), .Z(
        P2_U3479) );
  AOI22_X1 U10939 ( .A1(n10029), .A2(n11132), .B1(n11151), .B2(n10028), .ZN(
        n10031) );
  NAND2_X1 U10940 ( .A1(n10031), .A2(n10030), .ZN(n10048) );
  MUX2_X1 U10941 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n10048), .S(n11153), .Z(
        P2_U3478) );
  INV_X1 U10942 ( .A(n10032), .ZN(n10036) );
  NAND3_X1 U10943 ( .A1(n10033), .A2(n8529), .A3(n11132), .ZN(n10035) );
  OAI211_X1 U10944 ( .C1(n10036), .C2(n11127), .A(n10035), .B(n10034), .ZN(
        n10049) );
  MUX2_X1 U10945 ( .A(n10049), .B(P2_REG1_REG_18__SCAN_IN), .S(n5476), .Z(
        P2_U3477) );
  MUX2_X1 U10946 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n10037), .S(n11157), .Z(
        P2_U3458) );
  MUX2_X1 U10947 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n10038), .S(n11157), .Z(
        P2_U3457) );
  MUX2_X1 U10948 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n10039), .S(n11157), .Z(
        P2_U3455) );
  MUX2_X1 U10949 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n10040), .S(n11157), .Z(
        P2_U3454) );
  MUX2_X1 U10950 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n10041), .S(n11157), .Z(
        P2_U3453) );
  MUX2_X1 U10951 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n10042), .S(n11157), .Z(
        P2_U3452) );
  MUX2_X1 U10952 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n10043), .S(n11157), .Z(
        P2_U3451) );
  MUX2_X1 U10953 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n10044), .S(n11157), .Z(
        P2_U3450) );
  MUX2_X1 U10954 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n10045), .S(n11157), .Z(
        P2_U3449) );
  MUX2_X1 U10955 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n10046), .S(n11157), .Z(
        P2_U3448) );
  MUX2_X1 U10956 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n10047), .S(n11157), .Z(
        P2_U3447) );
  MUX2_X1 U10957 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n10048), .S(n11157), .Z(
        P2_U3446) );
  MUX2_X1 U10958 ( .A(n10049), .B(P2_REG0_REG_18__SCAN_IN), .S(n11154), .Z(
        P2_U3444) );
  NAND3_X1 U10959 ( .A1(n10050), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n10051) );
  OAI22_X1 U10960 ( .A1(n10052), .A2(n10051), .B1(n7211), .B2(n8985), .ZN(
        n10053) );
  AOI21_X1 U10961 ( .B1(n10664), .B2(n10054), .A(n10053), .ZN(n10055) );
  INV_X1 U10962 ( .A(n10055), .ZN(P2_U3264) );
  MUX2_X1 U10963 ( .A(n10056), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10964 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(n10060) );
  NAND2_X1 U10965 ( .A1(n10060), .A2(n11097), .ZN(n10065) );
  OAI22_X1 U10966 ( .A1(n10091), .A2(n10194), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10061), .ZN(n10063) );
  INV_X1 U10967 ( .A(n10189), .ZN(n11094) );
  OAI22_X1 U10968 ( .A1(n10082), .A2(n11094), .B1(n11101), .B2(n10407), .ZN(
        n10062) );
  AOI211_X1 U10969 ( .C1(n10405), .C2(n11088), .A(n10063), .B(n10062), .ZN(
        n10064) );
  NAND2_X1 U10970 ( .A1(n10065), .A2(n10064), .ZN(P1_U3216) );
  INV_X1 U10971 ( .A(n10066), .ZN(n10067) );
  AOI21_X1 U10972 ( .B1(n10069), .B2(n10068), .A(n10067), .ZN(n10075) );
  INV_X1 U10973 ( .A(n10070), .ZN(n10480) );
  AOI22_X1 U10974 ( .A1(n10480), .A2(n10190), .B1(n10189), .B2(n10510), .ZN(
        n10072) );
  OAI211_X1 U10975 ( .C1(n10081), .C2(n10194), .A(n10072), .B(n10071), .ZN(
        n10073) );
  AOI21_X1 U10976 ( .B1(n10479), .B2(n11088), .A(n10073), .ZN(n10074) );
  OAI21_X1 U10977 ( .B1(n10075), .B2(n10199), .A(n10074), .ZN(P1_U3219) );
  AOI21_X1 U10978 ( .B1(n10076), .B2(n10077), .A(n10199), .ZN(n10080) );
  NAND2_X1 U10979 ( .A1(n10080), .A2(n10079), .ZN(n10086) );
  NOR2_X1 U10980 ( .A1(n11094), .A2(n10081), .ZN(n10084) );
  OAI22_X1 U10981 ( .A1(n10082), .A2(n10194), .B1(n11101), .B2(n10450), .ZN(
        n10083) );
  AOI211_X1 U10982 ( .C1(P1_REG3_REG_21__SCAN_IN), .C2(P1_U3086), .A(n10084), 
        .B(n10083), .ZN(n10085) );
  OAI211_X1 U10983 ( .C1(n10449), .C2(n10183), .A(n10086), .B(n10085), .ZN(
        P1_U3223) );
  AOI21_X1 U10984 ( .B1(n10088), .B2(n10087), .A(n10176), .ZN(n10095) );
  OAI22_X1 U10985 ( .A1(n10090), .A2(n10194), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10089), .ZN(n10093) );
  OAI22_X1 U10986 ( .A1(n10091), .A2(n11094), .B1(n11101), .B2(n10375), .ZN(
        n10092) );
  AOI211_X1 U10987 ( .C1(n10373), .C2(n11088), .A(n10093), .B(n10092), .ZN(
        n10094) );
  OAI21_X1 U10988 ( .B1(n10095), .B2(n10199), .A(n10094), .ZN(P1_U3225) );
  OAI21_X1 U10989 ( .B1(n10098), .B2(n10097), .A(n10096), .ZN(n10099) );
  NAND2_X1 U10990 ( .A1(n10099), .A2(n11097), .ZN(n10105) );
  NAND2_X1 U10991 ( .A1(n10189), .A2(n10202), .ZN(n10100) );
  OAI21_X1 U10992 ( .B1(n11101), .B2(n10101), .A(n10100), .ZN(n10102) );
  AOI211_X1 U10993 ( .C1(n11091), .C2(n10492), .A(n10103), .B(n10102), .ZN(
        n10104) );
  OAI211_X1 U10994 ( .C1(n10106), .C2(n10183), .A(n10105), .B(n10104), .ZN(
        P1_U3226) );
  INV_X1 U10995 ( .A(n10107), .ZN(n10112) );
  AOI21_X1 U10996 ( .B1(n10111), .B2(n10109), .A(n10108), .ZN(n10110) );
  AOI21_X1 U10997 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(n10119) );
  INV_X1 U10998 ( .A(n10113), .ZN(n10522) );
  AOI22_X1 U10999 ( .A1(n10522), .A2(n10190), .B1(n10189), .B2(n10508), .ZN(
        n10115) );
  OAI211_X1 U11000 ( .C1(n10116), .C2(n10194), .A(n10115), .B(n10114), .ZN(
        n10117) );
  AOI21_X1 U11001 ( .B1(n10594), .B2(n11088), .A(n10117), .ZN(n10118) );
  OAI21_X1 U11002 ( .B1(n10119), .B2(n10199), .A(n10118), .ZN(P1_U3228) );
  INV_X1 U11003 ( .A(n10120), .ZN(n10122) );
  NAND2_X1 U11004 ( .A1(n10122), .A2(n10121), .ZN(n10123) );
  XNOR2_X1 U11005 ( .A(n10124), .B(n10123), .ZN(n10131) );
  OAI22_X1 U11006 ( .A1(n10126), .A2(n10194), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10125), .ZN(n10129) );
  INV_X1 U11007 ( .A(n10395), .ZN(n10127) );
  OAI22_X1 U11008 ( .A1(n10147), .A2(n11094), .B1(n10127), .B2(n11101), .ZN(
        n10128) );
  AOI211_X1 U11009 ( .C1(n10558), .C2(n11088), .A(n10129), .B(n10128), .ZN(
        n10130) );
  OAI21_X1 U11010 ( .B1(n10131), .B2(n10199), .A(n10130), .ZN(P1_U3229) );
  OAI21_X1 U11011 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(n10135) );
  NAND2_X1 U11012 ( .A1(n10135), .A2(n11097), .ZN(n10139) );
  AOI22_X1 U11013 ( .A1(n11091), .A2(n10464), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10138) );
  AOI22_X1 U11014 ( .A1(n10459), .A2(n10190), .B1(n10189), .B2(n10493), .ZN(
        n10137) );
  NAND2_X1 U11015 ( .A1(n10578), .A2(n11088), .ZN(n10136) );
  NAND4_X1 U11016 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        P1_U3233) );
  INV_X1 U11017 ( .A(n10140), .ZN(n10141) );
  NOR2_X1 U11018 ( .A1(n10142), .A2(n10141), .ZN(n10144) );
  XNOR2_X1 U11019 ( .A(n10144), .B(n10143), .ZN(n10151) );
  OAI22_X1 U11020 ( .A1(n11094), .A2(n10146), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10145), .ZN(n10149) );
  OAI22_X1 U11021 ( .A1(n10147), .A2(n10194), .B1(n11101), .B2(n10429), .ZN(
        n10148) );
  AOI211_X1 U11022 ( .C1(n10568), .C2(n11088), .A(n10149), .B(n10148), .ZN(
        n10150) );
  OAI21_X1 U11023 ( .B1(n10151), .B2(n10199), .A(n10150), .ZN(P1_U3235) );
  NAND2_X1 U11024 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  XOR2_X1 U11025 ( .A(n10155), .B(n10154), .Z(n10160) );
  AOI22_X1 U11026 ( .A1(n10499), .A2(n10190), .B1(n10189), .B2(n10492), .ZN(
        n10156) );
  NAND2_X1 U11027 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10831)
         );
  OAI211_X1 U11028 ( .C1(n10157), .C2(n10194), .A(n10156), .B(n10831), .ZN(
        n10158) );
  AOI21_X1 U11029 ( .B1(n10498), .B2(n11088), .A(n10158), .ZN(n10159) );
  OAI21_X1 U11030 ( .B1(n10160), .B2(n10199), .A(n10159), .ZN(P1_U3238) );
  NOR2_X1 U11031 ( .A1(n5566), .A2(n10163), .ZN(n10164) );
  XNOR2_X1 U11032 ( .A(n10161), .B(n10164), .ZN(n10165) );
  NAND2_X1 U11033 ( .A1(n10165), .A2(n11097), .ZN(n10172) );
  AOI22_X1 U11034 ( .A1(n10166), .A2(n11088), .B1(n11091), .B2(n10208), .ZN(
        n10171) );
  NAND2_X1 U11035 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10286) );
  INV_X1 U11036 ( .A(n10286), .ZN(n10167) );
  AOI21_X1 U11037 ( .B1(n10189), .B2(n10210), .A(n10167), .ZN(n10170) );
  OR2_X1 U11038 ( .A1(n11101), .A2(n10168), .ZN(n10169) );
  NAND4_X1 U11039 ( .A1(n10172), .A2(n10171), .A3(n10170), .A4(n10169), .ZN(
        P1_U3239) );
  INV_X1 U11040 ( .A(n10173), .ZN(n10178) );
  OAI21_X1 U11041 ( .B1(n10176), .B2(n10175), .A(n10174), .ZN(n10177) );
  NAND3_X1 U11042 ( .A1(n10178), .A2(n11097), .A3(n10177), .ZN(n10182) );
  AOI22_X1 U11043 ( .A1(n10391), .A2(n10189), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10179) );
  OAI21_X1 U11044 ( .B1(n11101), .B2(n10355), .A(n10179), .ZN(n10180) );
  AOI21_X1 U11045 ( .B1(n11091), .B2(n10363), .A(n10180), .ZN(n10181) );
  OAI211_X1 U11046 ( .C1(n10632), .C2(n10183), .A(n10182), .B(n10181), .ZN(
        P1_U3240) );
  NAND2_X1 U11047 ( .A1(n10185), .A2(n10184), .ZN(n10187) );
  XNOR2_X1 U11048 ( .A(n10187), .B(n10186), .ZN(n10200) );
  INV_X1 U11049 ( .A(n10188), .ZN(n10191) );
  AOI22_X1 U11050 ( .A1(n10191), .A2(n10190), .B1(n10189), .B2(n10203), .ZN(
        n10193) );
  OR2_X1 U11051 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10192), .ZN(n10815) );
  OAI211_X1 U11052 ( .C1(n10195), .C2(n10194), .A(n10193), .B(n10815), .ZN(
        n10196) );
  AOI21_X1 U11053 ( .B1(n10197), .B2(n11088), .A(n10196), .ZN(n10198) );
  OAI21_X1 U11054 ( .B1(n10200), .B2(n10199), .A(n10198), .ZN(P1_U3241) );
  MUX2_X1 U11055 ( .A(n10201), .B(P1_DATAO_REG_30__SCAN_IN), .S(n10215), .Z(
        P1_U3584) );
  MUX2_X1 U11056 ( .A(n10338), .B(P1_DATAO_REG_28__SCAN_IN), .S(n10215), .Z(
        P1_U3582) );
  MUX2_X1 U11057 ( .A(n10363), .B(P1_DATAO_REG_27__SCAN_IN), .S(n10215), .Z(
        P1_U3581) );
  MUX2_X1 U11058 ( .A(n10381), .B(P1_DATAO_REG_26__SCAN_IN), .S(n10215), .Z(
        P1_U3580) );
  MUX2_X1 U11059 ( .A(n10391), .B(P1_DATAO_REG_25__SCAN_IN), .S(n10215), .Z(
        P1_U3579) );
  MUX2_X1 U11060 ( .A(n10416), .B(P1_DATAO_REG_24__SCAN_IN), .S(n10215), .Z(
        P1_U3578) );
  MUX2_X1 U11061 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10441), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U11062 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10464), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U11063 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10474), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U11064 ( .A(n10493), .B(P1_DATAO_REG_19__SCAN_IN), .S(n10215), .Z(
        P1_U3573) );
  MUX2_X1 U11065 ( .A(n10510), .B(P1_DATAO_REG_18__SCAN_IN), .S(n10215), .Z(
        P1_U3572) );
  MUX2_X1 U11066 ( .A(n10492), .B(P1_DATAO_REG_17__SCAN_IN), .S(n10215), .Z(
        P1_U3571) );
  MUX2_X1 U11067 ( .A(n10508), .B(P1_DATAO_REG_16__SCAN_IN), .S(n10215), .Z(
        P1_U3570) );
  MUX2_X1 U11068 ( .A(n10202), .B(P1_DATAO_REG_15__SCAN_IN), .S(n10215), .Z(
        P1_U3569) );
  MUX2_X1 U11069 ( .A(n10203), .B(P1_DATAO_REG_14__SCAN_IN), .S(n10215), .Z(
        P1_U3568) );
  MUX2_X1 U11070 ( .A(n10204), .B(P1_DATAO_REG_13__SCAN_IN), .S(n10215), .Z(
        P1_U3567) );
  MUX2_X1 U11071 ( .A(n11090), .B(P1_DATAO_REG_12__SCAN_IN), .S(n10215), .Z(
        P1_U3566) );
  MUX2_X1 U11072 ( .A(n10205), .B(P1_DATAO_REG_11__SCAN_IN), .S(n10215), .Z(
        P1_U3565) );
  MUX2_X1 U11073 ( .A(n10206), .B(P1_DATAO_REG_9__SCAN_IN), .S(n10215), .Z(
        P1_U3563) );
  MUX2_X1 U11074 ( .A(n10207), .B(P1_DATAO_REG_8__SCAN_IN), .S(n10215), .Z(
        P1_U3562) );
  MUX2_X1 U11075 ( .A(n10208), .B(P1_DATAO_REG_7__SCAN_IN), .S(n10215), .Z(
        P1_U3561) );
  MUX2_X1 U11076 ( .A(n10209), .B(P1_DATAO_REG_6__SCAN_IN), .S(n10215), .Z(
        P1_U3560) );
  MUX2_X1 U11077 ( .A(n10210), .B(P1_DATAO_REG_5__SCAN_IN), .S(n10215), .Z(
        P1_U3559) );
  MUX2_X1 U11078 ( .A(n10211), .B(P1_DATAO_REG_4__SCAN_IN), .S(n10215), .Z(
        P1_U3558) );
  MUX2_X1 U11079 ( .A(n10212), .B(P1_DATAO_REG_3__SCAN_IN), .S(n10215), .Z(
        P1_U3557) );
  MUX2_X1 U11080 ( .A(n10213), .B(P1_DATAO_REG_2__SCAN_IN), .S(n10215), .Z(
        P1_U3556) );
  MUX2_X1 U11081 ( .A(n10214), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10215), .Z(
        P1_U3555) );
  MUX2_X1 U11082 ( .A(n6858), .B(P1_DATAO_REG_0__SCAN_IN), .S(n10215), .Z(
        P1_U3554) );
  OAI211_X1 U11083 ( .C1(n10218), .C2(n10217), .A(n10794), .B(n10216), .ZN(
        n10226) );
  OAI211_X1 U11084 ( .C1(n10221), .C2(n10220), .A(n10822), .B(n10219), .ZN(
        n10225) );
  AOI22_X1 U11085 ( .A1(n10754), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10224) );
  NAND2_X1 U11086 ( .A1(n10858), .A2(n10222), .ZN(n10223) );
  NAND4_X1 U11087 ( .A1(n10226), .A2(n10225), .A3(n10224), .A4(n10223), .ZN(
        P1_U3244) );
  NAND2_X1 U11088 ( .A1(n10227), .A2(n10748), .ZN(n10228) );
  MUX2_X1 U11089 ( .A(n10228), .B(n10752), .S(n5123), .Z(n10233) );
  OAI21_X1 U11090 ( .B1(n10752), .B2(P1_REG2_REG_0__SCAN_IN), .A(n10229), .ZN(
        n10230) );
  AOI21_X1 U11091 ( .B1(n10231), .B2(n10230), .A(n10215), .ZN(n10232) );
  NAND2_X1 U11092 ( .A1(n10233), .A2(n10232), .ZN(n10272) );
  INV_X1 U11093 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10235) );
  OAI22_X1 U11094 ( .A1(n10862), .A2(n10235), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10234), .ZN(n10236) );
  AOI21_X1 U11095 ( .B1(n10237), .B2(n10858), .A(n10236), .ZN(n10246) );
  OAI211_X1 U11096 ( .C1(n10240), .C2(n10239), .A(n10794), .B(n10238), .ZN(
        n10245) );
  OAI211_X1 U11097 ( .C1(n10243), .C2(n10242), .A(n10822), .B(n10241), .ZN(
        n10244) );
  NAND4_X1 U11098 ( .A1(n10272), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        P1_U3245) );
  INV_X1 U11099 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10248) );
  OAI21_X1 U11100 ( .B1(n10862), .B2(n10248), .A(n10247), .ZN(n10249) );
  AOI21_X1 U11101 ( .B1(n10250), .B2(n10858), .A(n10249), .ZN(n10259) );
  OAI211_X1 U11102 ( .C1(n10253), .C2(n10252), .A(n10794), .B(n10251), .ZN(
        n10258) );
  OAI211_X1 U11103 ( .C1(n10256), .C2(n10255), .A(n10822), .B(n10254), .ZN(
        n10257) );
  NAND3_X1 U11104 ( .A1(n10259), .A2(n10258), .A3(n10257), .ZN(P1_U3246) );
  NOR2_X1 U11105 ( .A1(n10829), .A2(n10260), .ZN(n10261) );
  AOI211_X1 U11106 ( .C1(n10754), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n10262), .B(
        n10261), .ZN(n10271) );
  OAI211_X1 U11107 ( .C1(n10265), .C2(n10264), .A(n10822), .B(n10263), .ZN(
        n10270) );
  OAI211_X1 U11108 ( .C1(n10268), .C2(n10267), .A(n10794), .B(n10266), .ZN(
        n10269) );
  NAND4_X1 U11109 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        P1_U3247) );
  INV_X1 U11110 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10274) );
  OAI21_X1 U11111 ( .B1(n10862), .B2(n10274), .A(n10273), .ZN(n10275) );
  AOI21_X1 U11112 ( .B1(n10276), .B2(n10858), .A(n10275), .ZN(n10285) );
  OAI211_X1 U11113 ( .C1(n10279), .C2(n10278), .A(n10794), .B(n10277), .ZN(
        n10284) );
  OAI211_X1 U11114 ( .C1(n10282), .C2(n10281), .A(n10822), .B(n10280), .ZN(
        n10283) );
  NAND3_X1 U11115 ( .A1(n10285), .A2(n10284), .A3(n10283), .ZN(P1_U3248) );
  INV_X1 U11116 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10287) );
  OAI21_X1 U11117 ( .B1(n10862), .B2(n10287), .A(n10286), .ZN(n10288) );
  AOI21_X1 U11118 ( .B1(n10289), .B2(n10858), .A(n10288), .ZN(n10298) );
  OAI211_X1 U11119 ( .C1(n10292), .C2(n10291), .A(n10794), .B(n10290), .ZN(
        n10297) );
  OAI211_X1 U11120 ( .C1(n10295), .C2(n10294), .A(n10822), .B(n10293), .ZN(
        n10296) );
  NAND3_X1 U11121 ( .A1(n10298), .A2(n10297), .A3(n10296), .ZN(P1_U3249) );
  INV_X1 U11122 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10300) );
  OAI21_X1 U11123 ( .B1(n10862), .B2(n10300), .A(n10299), .ZN(n10301) );
  AOI21_X1 U11124 ( .B1(n10302), .B2(n10858), .A(n10301), .ZN(n10311) );
  OAI211_X1 U11125 ( .C1(n10305), .C2(n10304), .A(n10794), .B(n10303), .ZN(
        n10310) );
  OAI211_X1 U11126 ( .C1(n10308), .C2(n10307), .A(n10822), .B(n10306), .ZN(
        n10309) );
  NAND3_X1 U11127 ( .A1(n10311), .A2(n10310), .A3(n10309), .ZN(P1_U3250) );
  NAND2_X1 U11128 ( .A1(n10624), .A2(n10317), .ZN(n10316) );
  XNOR2_X1 U11129 ( .A(n10620), .B(n10316), .ZN(n10531) );
  NAND2_X1 U11130 ( .A1(n10531), .A2(n10454), .ZN(n10315) );
  AND2_X1 U11131 ( .A1(n10313), .A2(n10312), .ZN(n10530) );
  INV_X1 U11132 ( .A(n10530), .ZN(n10534) );
  NOR2_X1 U11133 ( .A1(n10529), .A2(n10534), .ZN(n10319) );
  AOI21_X1 U11134 ( .B1(n10529), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10319), 
        .ZN(n10314) );
  OAI211_X1 U11135 ( .C1(n10620), .C2(n10525), .A(n10315), .B(n10314), .ZN(
        P1_U3263) );
  OAI211_X1 U11136 ( .C1(n10624), .C2(n10317), .A(n10599), .B(n10316), .ZN(
        n10535) );
  AND2_X1 U11137 ( .A1(n10529), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n10318) );
  NOR2_X1 U11138 ( .A1(n10319), .A2(n10318), .ZN(n10322) );
  NAND2_X1 U11139 ( .A1(n10320), .A2(n11018), .ZN(n10321) );
  OAI211_X1 U11140 ( .C1(n10535), .C2(n11021), .A(n10322), .B(n10321), .ZN(
        P1_U3264) );
  OAI22_X1 U11141 ( .A1(n10324), .A2(n11012), .B1(n10323), .B2(n11015), .ZN(
        n10328) );
  INV_X1 U11142 ( .A(n10325), .ZN(n10326) );
  NOR2_X1 U11143 ( .A1(n10326), .A2(n10525), .ZN(n10327) );
  AOI211_X1 U11144 ( .C1(n10520), .C2(n10329), .A(n10328), .B(n10327), .ZN(
        n10332) );
  NAND2_X1 U11145 ( .A1(n10330), .A2(n11015), .ZN(n10331) );
  OAI211_X1 U11146 ( .C1(n10333), .C2(n10504), .A(n10332), .B(n10331), .ZN(
        P1_U3265) );
  XNOR2_X1 U11147 ( .A(n10334), .B(n10336), .ZN(n10543) );
  INV_X1 U11148 ( .A(n10543), .ZN(n10350) );
  OAI211_X1 U11149 ( .C1(n10337), .C2(n10336), .A(n10335), .B(n10512), .ZN(
        n10340) );
  AOI22_X1 U11150 ( .A1(n10338), .A2(n10509), .B1(n10507), .B2(n10381), .ZN(
        n10339) );
  NAND2_X1 U11151 ( .A1(n10340), .A2(n10339), .ZN(n10541) );
  INV_X1 U11152 ( .A(n10341), .ZN(n10342) );
  AOI211_X1 U11153 ( .C1(n10344), .C2(n10343), .A(n11049), .B(n10342), .ZN(
        n10542) );
  NAND2_X1 U11154 ( .A1(n10542), .A2(n10520), .ZN(n10347) );
  AOI22_X1 U11155 ( .A1(n10345), .A2(n10521), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10466), .ZN(n10346) );
  OAI211_X1 U11156 ( .C1(n10628), .C2(n10525), .A(n10347), .B(n10346), .ZN(
        n10348) );
  AOI21_X1 U11157 ( .B1(n10541), .B2(n11015), .A(n10348), .ZN(n10349) );
  OAI21_X1 U11158 ( .B1(n10350), .B2(n10504), .A(n10349), .ZN(P1_U3266) );
  XOR2_X1 U11159 ( .A(n10351), .B(n10358), .Z(n10548) );
  INV_X1 U11160 ( .A(n10548), .ZN(n10368) );
  AOI211_X1 U11161 ( .C1(n10353), .C2(n10370), .A(n11049), .B(n10352), .ZN(
        n10547) );
  NOR2_X1 U11162 ( .A1(n10632), .A2(n10525), .ZN(n10357) );
  OAI22_X1 U11163 ( .A1(n10355), .A2(n11012), .B1(n10354), .B2(n11015), .ZN(
        n10356) );
  AOI211_X1 U11164 ( .C1(n10547), .C2(n10520), .A(n10357), .B(n10356), .ZN(
        n10367) );
  NAND2_X1 U11165 ( .A1(n10359), .A2(n10358), .ZN(n10360) );
  NAND2_X1 U11166 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  NAND2_X1 U11167 ( .A1(n10362), .A2(n10512), .ZN(n10365) );
  AOI22_X1 U11168 ( .A1(n10363), .A2(n10509), .B1(n10507), .B2(n10391), .ZN(
        n10364) );
  NAND2_X1 U11169 ( .A1(n10365), .A2(n10364), .ZN(n10546) );
  NAND2_X1 U11170 ( .A1(n10546), .A2(n11015), .ZN(n10366) );
  OAI211_X1 U11171 ( .C1(n10368), .C2(n10504), .A(n10367), .B(n10366), .ZN(
        P1_U3267) );
  XOR2_X1 U11172 ( .A(n10369), .B(n10379), .Z(n10553) );
  INV_X1 U11173 ( .A(n10553), .ZN(n10386) );
  INV_X1 U11174 ( .A(n10394), .ZN(n10372) );
  INV_X1 U11175 ( .A(n10370), .ZN(n10371) );
  AOI211_X1 U11176 ( .C1(n10373), .C2(n10372), .A(n11049), .B(n10371), .ZN(
        n10552) );
  NOR2_X1 U11177 ( .A1(n10636), .A2(n10525), .ZN(n10377) );
  OAI22_X1 U11178 ( .A1(n10375), .A2(n11012), .B1(n10374), .B2(n11015), .ZN(
        n10376) );
  AOI211_X1 U11179 ( .C1(n10552), .C2(n10520), .A(n10377), .B(n10376), .ZN(
        n10385) );
  OAI211_X1 U11180 ( .C1(n10380), .C2(n10379), .A(n10378), .B(n10512), .ZN(
        n10383) );
  AOI22_X1 U11181 ( .A1(n10381), .A2(n10509), .B1(n10507), .B2(n10416), .ZN(
        n10382) );
  NAND2_X1 U11182 ( .A1(n10383), .A2(n10382), .ZN(n10551) );
  NAND2_X1 U11183 ( .A1(n10551), .A2(n11015), .ZN(n10384) );
  OAI211_X1 U11184 ( .C1(n10386), .C2(n10504), .A(n10385), .B(n10384), .ZN(
        P1_U3268) );
  XOR2_X1 U11185 ( .A(n10387), .B(n10389), .Z(n10560) );
  OAI211_X1 U11186 ( .C1(n10390), .C2(n10389), .A(n10388), .B(n10512), .ZN(
        n10393) );
  AOI22_X1 U11187 ( .A1(n10391), .A2(n10509), .B1(n10507), .B2(n10433), .ZN(
        n10392) );
  NAND2_X1 U11188 ( .A1(n10393), .A2(n10392), .ZN(n10557) );
  INV_X1 U11189 ( .A(n10558), .ZN(n10398) );
  AOI211_X1 U11190 ( .C1(n10558), .C2(n10403), .A(n11049), .B(n10394), .ZN(
        n10556) );
  NAND2_X1 U11191 ( .A1(n10556), .A2(n10520), .ZN(n10397) );
  AOI22_X1 U11192 ( .A1(n10395), .A2(n10521), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10466), .ZN(n10396) );
  OAI211_X1 U11193 ( .C1(n10398), .C2(n10525), .A(n10397), .B(n10396), .ZN(
        n10399) );
  AOI21_X1 U11194 ( .B1(n11015), .B2(n10557), .A(n10399), .ZN(n10400) );
  OAI21_X1 U11195 ( .B1(n10560), .B2(n10504), .A(n10400), .ZN(P1_U3269) );
  XNOR2_X1 U11196 ( .A(n10401), .B(n10411), .ZN(n10563) );
  INV_X1 U11197 ( .A(n10563), .ZN(n10421) );
  INV_X1 U11198 ( .A(n10403), .ZN(n10404) );
  AOI211_X1 U11199 ( .C1(n10405), .C2(n10426), .A(n11049), .B(n10404), .ZN(
        n10562) );
  NOR2_X1 U11200 ( .A1(n6315), .A2(n10525), .ZN(n10409) );
  OAI22_X1 U11201 ( .A1(n10407), .A2(n11012), .B1(n10406), .B2(n11015), .ZN(
        n10408) );
  AOI211_X1 U11202 ( .C1(n10562), .C2(n10520), .A(n10409), .B(n10408), .ZN(
        n10420) );
  NAND2_X1 U11203 ( .A1(n10432), .A2(n10410), .ZN(n10412) );
  NAND2_X1 U11204 ( .A1(n10412), .A2(n10411), .ZN(n10413) );
  NAND2_X1 U11205 ( .A1(n10414), .A2(n10413), .ZN(n10415) );
  NAND2_X1 U11206 ( .A1(n10415), .A2(n10512), .ZN(n10418) );
  AOI22_X1 U11207 ( .A1(n10416), .A2(n10509), .B1(n10507), .B2(n10441), .ZN(
        n10417) );
  NAND2_X1 U11208 ( .A1(n10418), .A2(n10417), .ZN(n10561) );
  NAND2_X1 U11209 ( .A1(n10561), .A2(n11015), .ZN(n10419) );
  OAI211_X1 U11210 ( .C1(n10421), .C2(n10504), .A(n10420), .B(n10419), .ZN(
        P1_U3270) );
  OAI21_X1 U11211 ( .B1(n10424), .B2(n10423), .A(n10422), .ZN(n10425) );
  INV_X1 U11212 ( .A(n10425), .ZN(n10570) );
  AOI211_X1 U11213 ( .C1(n10568), .C2(n10446), .A(n11049), .B(n10402), .ZN(
        n10566) );
  NOR2_X1 U11214 ( .A1(n10427), .A2(n10525), .ZN(n10431) );
  OAI22_X1 U11215 ( .A1(n10429), .A2(n11012), .B1(n11015), .B2(n10428), .ZN(
        n10430) );
  AOI211_X1 U11216 ( .C1(n10566), .C2(n10520), .A(n10431), .B(n10430), .ZN(
        n10437) );
  AOI22_X1 U11217 ( .A1(n10433), .A2(n10509), .B1(n10507), .B2(n10464), .ZN(
        n10434) );
  NAND2_X1 U11218 ( .A1(n10435), .A2(n10434), .ZN(n10567) );
  NAND2_X1 U11219 ( .A1(n10567), .A2(n11015), .ZN(n10436) );
  OAI211_X1 U11220 ( .C1(n10570), .C2(n10504), .A(n10437), .B(n10436), .ZN(
        P1_U3271) );
  NAND2_X1 U11221 ( .A1(n10439), .A2(n10438), .ZN(n10440) );
  XOR2_X1 U11222 ( .A(n10444), .B(n10440), .Z(n10442) );
  AOI222_X1 U11223 ( .A1(n10512), .A2(n10442), .B1(n10441), .B2(n10509), .C1(
        n10474), .C2(n10507), .ZN(n10575) );
  OAI21_X1 U11224 ( .B1(n10445), .B2(n10444), .A(n10443), .ZN(n10571) );
  NAND2_X1 U11225 ( .A1(n10571), .A2(n11023), .ZN(n10456) );
  INV_X1 U11226 ( .A(n10458), .ZN(n10448) );
  INV_X1 U11227 ( .A(n10446), .ZN(n10447) );
  AOI21_X1 U11228 ( .B1(n10572), .B2(n10448), .A(n10447), .ZN(n10573) );
  NOR2_X1 U11229 ( .A1(n10449), .A2(n10525), .ZN(n10453) );
  OAI22_X1 U11230 ( .A1(n11015), .A2(n10451), .B1(n10450), .B2(n11012), .ZN(
        n10452) );
  AOI211_X1 U11231 ( .C1(n10573), .C2(n10454), .A(n10453), .B(n10452), .ZN(
        n10455) );
  OAI211_X1 U11232 ( .C1(n10529), .C2(n10575), .A(n10456), .B(n10455), .ZN(
        P1_U3272) );
  XOR2_X1 U11233 ( .A(n10463), .B(n10457), .Z(n10581) );
  AOI211_X1 U11234 ( .C1(n10578), .C2(n10477), .A(n11049), .B(n10458), .ZN(
        n10577) );
  INV_X1 U11235 ( .A(n10578), .ZN(n10461) );
  AOI22_X1 U11236 ( .A1(n10529), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10459), 
        .B2(n10521), .ZN(n10460) );
  OAI21_X1 U11237 ( .B1(n10461), .B2(n10525), .A(n10460), .ZN(n10468) );
  XNOR2_X1 U11238 ( .A(n10463), .B(n10462), .ZN(n10465) );
  AOI222_X1 U11239 ( .A1(n10512), .A2(n10465), .B1(n10493), .B2(n10507), .C1(
        n10464), .C2(n10509), .ZN(n10580) );
  NOR2_X1 U11240 ( .A1(n10580), .A2(n10466), .ZN(n10467) );
  AOI211_X1 U11241 ( .C1(n10577), .C2(n10520), .A(n10468), .B(n10467), .ZN(
        n10469) );
  OAI21_X1 U11242 ( .B1(n10504), .B2(n10581), .A(n10469), .ZN(P1_U3273) );
  XNOR2_X1 U11243 ( .A(n10470), .B(n5517), .ZN(n10584) );
  INV_X1 U11244 ( .A(n10584), .ZN(n10485) );
  OAI21_X1 U11245 ( .B1(n5517), .B2(n10472), .A(n10471), .ZN(n10473) );
  NAND2_X1 U11246 ( .A1(n10473), .A2(n10512), .ZN(n10476) );
  AOI22_X1 U11247 ( .A1(n10474), .A2(n10509), .B1(n10507), .B2(n10510), .ZN(
        n10475) );
  NAND2_X1 U11248 ( .A1(n10476), .A2(n10475), .ZN(n10582) );
  INV_X1 U11249 ( .A(n10479), .ZN(n10647) );
  INV_X1 U11250 ( .A(n10477), .ZN(n10478) );
  AOI211_X1 U11251 ( .C1(n10479), .C2(n10496), .A(n11049), .B(n10478), .ZN(
        n10583) );
  NAND2_X1 U11252 ( .A1(n10583), .A2(n10520), .ZN(n10482) );
  AOI22_X1 U11253 ( .A1(n10529), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10480), 
        .B2(n10521), .ZN(n10481) );
  OAI211_X1 U11254 ( .C1(n10647), .C2(n10525), .A(n10482), .B(n10481), .ZN(
        n10483) );
  AOI21_X1 U11255 ( .B1(n11015), .B2(n10582), .A(n10483), .ZN(n10484) );
  OAI21_X1 U11256 ( .B1(n10485), .B2(n10504), .A(n10484), .ZN(P1_U3274) );
  XOR2_X1 U11257 ( .A(n10489), .B(n10486), .Z(n10589) );
  INV_X1 U11258 ( .A(n10589), .ZN(n10505) );
  NAND2_X1 U11259 ( .A1(n10488), .A2(n10487), .ZN(n10490) );
  XNOR2_X1 U11260 ( .A(n10490), .B(n10489), .ZN(n10491) );
  NAND2_X1 U11261 ( .A1(n10491), .A2(n10512), .ZN(n10495) );
  AOI22_X1 U11262 ( .A1(n10493), .A2(n10509), .B1(n10507), .B2(n10492), .ZN(
        n10494) );
  NAND2_X1 U11263 ( .A1(n10495), .A2(n10494), .ZN(n10587) );
  INV_X1 U11264 ( .A(n10496), .ZN(n10497) );
  AOI211_X1 U11265 ( .C1(n10498), .C2(n5335), .A(n11049), .B(n10497), .ZN(
        n10588) );
  NAND2_X1 U11266 ( .A1(n10588), .A2(n10520), .ZN(n10501) );
  AOI22_X1 U11267 ( .A1(n10529), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10499), 
        .B2(n10521), .ZN(n10500) );
  OAI211_X1 U11268 ( .C1(n10652), .C2(n10525), .A(n10501), .B(n10500), .ZN(
        n10502) );
  AOI21_X1 U11269 ( .B1(n11015), .B2(n10587), .A(n10502), .ZN(n10503) );
  OAI21_X1 U11270 ( .B1(n10505), .B2(n10504), .A(n10503), .ZN(P1_U3275) );
  XNOR2_X1 U11271 ( .A(n10514), .B(n10506), .ZN(n10511) );
  AOI222_X1 U11272 ( .A1(n10512), .A2(n10511), .B1(n10510), .B2(n10509), .C1(
        n10508), .C2(n10507), .ZN(n10596) );
  OAI21_X1 U11273 ( .B1(n10515), .B2(n10514), .A(n10513), .ZN(n10597) );
  INV_X1 U11274 ( .A(n10597), .ZN(n10527) );
  NAND2_X1 U11275 ( .A1(n10594), .A2(n10516), .ZN(n10517) );
  NAND2_X1 U11276 ( .A1(n10517), .A2(n10599), .ZN(n10518) );
  NOR2_X1 U11277 ( .A1(n10519), .A2(n10518), .ZN(n10593) );
  NAND2_X1 U11278 ( .A1(n10593), .A2(n10520), .ZN(n10524) );
  AOI22_X1 U11279 ( .A1(n10466), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10522), 
        .B2(n10521), .ZN(n10523) );
  OAI211_X1 U11280 ( .C1(n5333), .C2(n10525), .A(n10524), .B(n10523), .ZN(
        n10526) );
  AOI21_X1 U11281 ( .B1(n10527), .B2(n11023), .A(n10526), .ZN(n10528) );
  OAI21_X1 U11282 ( .B1(n10529), .B2(n10596), .A(n10528), .ZN(P1_U3276) );
  AOI21_X1 U11283 ( .B1(n10531), .B2(n10599), .A(n10530), .ZN(n10617) );
  MUX2_X1 U11284 ( .A(n10532), .B(n10617), .S(n11116), .Z(n10533) );
  OAI21_X1 U11285 ( .B1(n10620), .B2(n10592), .A(n10533), .ZN(P1_U3553) );
  AND2_X1 U11286 ( .A1(n10535), .A2(n10534), .ZN(n10621) );
  MUX2_X1 U11287 ( .A(n8648), .B(n10621), .S(n11116), .Z(n10536) );
  OAI21_X1 U11288 ( .B1(n10624), .B2(n10592), .A(n10536), .ZN(P1_U3552) );
  INV_X1 U11289 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10544) );
  AOI211_X1 U11290 ( .C1(n10543), .C2(n11113), .A(n10542), .B(n10541), .ZN(
        n10625) );
  MUX2_X1 U11291 ( .A(n10544), .B(n10625), .S(n11116), .Z(n10545) );
  OAI21_X1 U11292 ( .B1(n10628), .B2(n10592), .A(n10545), .ZN(P1_U3549) );
  INV_X1 U11293 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10549) );
  AOI211_X1 U11294 ( .C1(n10548), .C2(n11113), .A(n10547), .B(n10546), .ZN(
        n10629) );
  MUX2_X1 U11295 ( .A(n10549), .B(n10629), .S(n11116), .Z(n10550) );
  OAI21_X1 U11296 ( .B1(n10632), .B2(n10592), .A(n10550), .ZN(P1_U3548) );
  INV_X1 U11297 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10554) );
  AOI211_X1 U11298 ( .C1(n10553), .C2(n11113), .A(n10552), .B(n10551), .ZN(
        n10633) );
  MUX2_X1 U11299 ( .A(n10554), .B(n10633), .S(n11116), .Z(n10555) );
  OAI21_X1 U11300 ( .B1(n10636), .B2(n10592), .A(n10555), .ZN(P1_U3547) );
  AOI211_X1 U11301 ( .C1(n10996), .C2(n10558), .A(n10557), .B(n10556), .ZN(
        n10559) );
  OAI21_X1 U11302 ( .B1(n10560), .B2(n11000), .A(n10559), .ZN(n10637) );
  MUX2_X1 U11303 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10637), .S(n11116), .Z(
        P1_U3546) );
  INV_X1 U11304 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10564) );
  AOI211_X1 U11305 ( .C1(n10563), .C2(n11113), .A(n10562), .B(n10561), .ZN(
        n10638) );
  MUX2_X1 U11306 ( .A(n10564), .B(n10638), .S(n11116), .Z(n10565) );
  OAI21_X1 U11307 ( .B1(n6315), .B2(n10592), .A(n10565), .ZN(P1_U3545) );
  AOI211_X1 U11308 ( .C1(n10996), .C2(n10568), .A(n10567), .B(n10566), .ZN(
        n10569) );
  OAI21_X1 U11309 ( .B1(n10570), .B2(n11000), .A(n10569), .ZN(n10641) );
  MUX2_X1 U11310 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10641), .S(n11116), .Z(
        P1_U3544) );
  INV_X1 U11311 ( .A(n10571), .ZN(n10576) );
  AOI22_X1 U11312 ( .A1(n10573), .A2(n10599), .B1(n10996), .B2(n10572), .ZN(
        n10574) );
  OAI211_X1 U11313 ( .C1(n10576), .C2(n11000), .A(n10575), .B(n10574), .ZN(
        n10642) );
  MUX2_X1 U11314 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10642), .S(n11116), .Z(
        P1_U3543) );
  AOI21_X1 U11315 ( .B1(n10996), .B2(n10578), .A(n10577), .ZN(n10579) );
  OAI211_X1 U11316 ( .C1(n10581), .C2(n11000), .A(n10580), .B(n10579), .ZN(
        n10643) );
  MUX2_X1 U11317 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10643), .S(n11116), .Z(
        P1_U3542) );
  AOI211_X1 U11318 ( .C1(n10584), .C2(n11113), .A(n10583), .B(n10582), .ZN(
        n10644) );
  MUX2_X1 U11319 ( .A(n10585), .B(n10644), .S(n11116), .Z(n10586) );
  OAI21_X1 U11320 ( .B1(n10647), .B2(n10592), .A(n10586), .ZN(P1_U3541) );
  INV_X1 U11321 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10590) );
  AOI211_X1 U11322 ( .C1(n10589), .C2(n11113), .A(n10588), .B(n10587), .ZN(
        n10648) );
  MUX2_X1 U11323 ( .A(n10590), .B(n10648), .S(n11116), .Z(n10591) );
  OAI21_X1 U11324 ( .B1(n10652), .B2(n10592), .A(n10591), .ZN(P1_U3540) );
  AOI21_X1 U11325 ( .B1(n10996), .B2(n10594), .A(n10593), .ZN(n10595) );
  OAI211_X1 U11326 ( .C1(n10597), .C2(n11000), .A(n10596), .B(n10595), .ZN(
        n10653) );
  MUX2_X1 U11327 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10653), .S(n11116), .Z(
        P1_U3539) );
  AOI22_X1 U11328 ( .A1(n10600), .A2(n10599), .B1(n10996), .B2(n10598), .ZN(
        n10601) );
  OAI211_X1 U11329 ( .C1(n10603), .C2(n11000), .A(n10602), .B(n10601), .ZN(
        n10654) );
  MUX2_X1 U11330 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10654), .S(n11116), .Z(
        P1_U3538) );
  OR2_X1 U11331 ( .A1(n10604), .A2(n11000), .ZN(n10610) );
  OAI21_X1 U11332 ( .B1(n10606), .B2(n11109), .A(n10605), .ZN(n10607) );
  NOR2_X1 U11333 ( .A1(n10608), .A2(n10607), .ZN(n10609) );
  NAND2_X1 U11334 ( .A1(n10610), .A2(n10609), .ZN(n10655) );
  MUX2_X1 U11335 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10655), .S(n11116), .Z(
        P1_U3537) );
  AOI21_X1 U11336 ( .B1(n10996), .B2(n10612), .A(n10611), .ZN(n10613) );
  OAI211_X1 U11337 ( .C1(n10616), .C2(n10615), .A(n10614), .B(n10613), .ZN(
        n10656) );
  MUX2_X1 U11338 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10656), .S(n11116), .Z(
        P1_U3536) );
  INV_X1 U11339 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10618) );
  MUX2_X1 U11340 ( .A(n10618), .B(n10617), .S(n11120), .Z(n10619) );
  OAI21_X1 U11341 ( .B1(n10620), .B2(n10651), .A(n10619), .ZN(P1_U3521) );
  INV_X1 U11342 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10622) );
  MUX2_X1 U11343 ( .A(n10622), .B(n10621), .S(n11120), .Z(n10623) );
  OAI21_X1 U11344 ( .B1(n10624), .B2(n10651), .A(n10623), .ZN(P1_U3520) );
  INV_X1 U11345 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10626) );
  MUX2_X1 U11346 ( .A(n10626), .B(n10625), .S(n11120), .Z(n10627) );
  OAI21_X1 U11347 ( .B1(n10628), .B2(n10651), .A(n10627), .ZN(P1_U3517) );
  INV_X1 U11348 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10630) );
  MUX2_X1 U11349 ( .A(n10630), .B(n10629), .S(n11120), .Z(n10631) );
  OAI21_X1 U11350 ( .B1(n10632), .B2(n10651), .A(n10631), .ZN(P1_U3516) );
  INV_X1 U11351 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10634) );
  MUX2_X1 U11352 ( .A(n10634), .B(n10633), .S(n11120), .Z(n10635) );
  OAI21_X1 U11353 ( .B1(n10636), .B2(n10651), .A(n10635), .ZN(P1_U3515) );
  MUX2_X1 U11354 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10637), .S(n11120), .Z(
        P1_U3514) );
  INV_X1 U11355 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10639) );
  MUX2_X1 U11356 ( .A(n10639), .B(n10638), .S(n11120), .Z(n10640) );
  OAI21_X1 U11357 ( .B1(n6315), .B2(n10651), .A(n10640), .ZN(P1_U3513) );
  MUX2_X1 U11358 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10641), .S(n11120), .Z(
        P1_U3512) );
  MUX2_X1 U11359 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10642), .S(n11120), .Z(
        P1_U3511) );
  MUX2_X1 U11360 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10643), .S(n11120), .Z(
        P1_U3510) );
  INV_X1 U11361 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10645) );
  MUX2_X1 U11362 ( .A(n10645), .B(n10644), .S(n11120), .Z(n10646) );
  OAI21_X1 U11363 ( .B1(n10647), .B2(n10651), .A(n10646), .ZN(P1_U3509) );
  INV_X1 U11364 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10649) );
  MUX2_X1 U11365 ( .A(n10649), .B(n10648), .S(n11120), .Z(n10650) );
  OAI21_X1 U11366 ( .B1(n10652), .B2(n10651), .A(n10650), .ZN(P1_U3507) );
  MUX2_X1 U11367 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10653), .S(n11120), .Z(
        P1_U3504) );
  MUX2_X1 U11368 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10654), .S(n11120), .Z(
        P1_U3501) );
  MUX2_X1 U11369 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10655), .S(n11120), .Z(
        P1_U3498) );
  MUX2_X1 U11370 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10656), .S(n11120), .Z(
        P1_U3495) );
  NAND3_X1 U11371 ( .A1(n10658), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n10661) );
  OAI22_X1 U11372 ( .A1(n10657), .A2(n10661), .B1(n10660), .B2(n10659), .ZN(
        n10662) );
  AOI21_X1 U11373 ( .B1(n10664), .B2(n10663), .A(n10662), .ZN(n10665) );
  INV_X1 U11374 ( .A(n10665), .ZN(P1_U3324) );
  MUX2_X1 U11375 ( .A(n10666), .B(n10752), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  INV_X1 U11376 ( .A(n10671), .ZN(n10670) );
  NOR2_X1 U11377 ( .A1(n10670), .A2(n10667), .ZN(P1_U3323) );
  NOR2_X1 U11378 ( .A1(n10670), .A2(n10668), .ZN(P1_U3322) );
  NOR2_X1 U11379 ( .A1(n10670), .A2(n10669), .ZN(P1_U3321) );
  AND2_X1 U11380 ( .A1(n10671), .A2(P1_D_REG_5__SCAN_IN), .ZN(P1_U3320) );
  AND2_X1 U11381 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10671), .ZN(P1_U3319) );
  AND2_X1 U11382 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10671), .ZN(P1_U3318) );
  AND2_X1 U11383 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10671), .ZN(P1_U3317) );
  AND2_X1 U11384 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10671), .ZN(P1_U3316) );
  AND2_X1 U11385 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10671), .ZN(P1_U3315) );
  AND2_X1 U11386 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10671), .ZN(P1_U3314) );
  AND2_X1 U11387 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10671), .ZN(P1_U3313) );
  AND2_X1 U11388 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10671), .ZN(P1_U3312) );
  AND2_X1 U11389 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10671), .ZN(P1_U3311) );
  AND2_X1 U11390 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10671), .ZN(P1_U3310) );
  AND2_X1 U11391 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10671), .ZN(P1_U3309) );
  AND2_X1 U11392 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10671), .ZN(P1_U3308) );
  AND2_X1 U11393 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10671), .ZN(P1_U3307) );
  AND2_X1 U11394 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10671), .ZN(P1_U3306) );
  AND2_X1 U11395 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10671), .ZN(P1_U3305) );
  AND2_X1 U11396 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10671), .ZN(P1_U3304) );
  AND2_X1 U11397 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10671), .ZN(P1_U3303) );
  AND2_X1 U11398 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10671), .ZN(P1_U3302) );
  AND2_X1 U11399 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10671), .ZN(P1_U3301) );
  AND2_X1 U11400 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10671), .ZN(P1_U3300) );
  AND2_X1 U11401 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10671), .ZN(P1_U3299) );
  AND2_X1 U11402 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10671), .ZN(P1_U3298) );
  AND2_X1 U11403 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10671), .ZN(P1_U3297) );
  AND2_X1 U11404 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10671), .ZN(P1_U3296) );
  AND2_X1 U11405 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10671), .ZN(P1_U3295) );
  AND2_X1 U11406 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10671), .ZN(P1_U3294) );
  NAND2_X1 U11407 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n10675) );
  OAI21_X1 U11408 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(n10675), .ZN(n10672) );
  INV_X1 U11409 ( .A(n10672), .ZN(ADD_1068_U46) );
  INV_X1 U11410 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10673) );
  NAND2_X1 U11411 ( .A1(n10673), .A2(n10675), .ZN(n10676) );
  OAI21_X1 U11412 ( .B1(n10673), .B2(n10675), .A(n10676), .ZN(n10674) );
  XNOR2_X1 U11413 ( .A(n10674), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1068_U5)
         );
  INV_X1 U11414 ( .A(n10675), .ZN(n10677) );
  AOI22_X1 U11415 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10677), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10676), .ZN(n10680) );
  NAND2_X1 U11416 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10678) );
  OAI21_X1 U11417 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10678), .ZN(n10679) );
  NOR2_X1 U11418 ( .A1(n10680), .A2(n10679), .ZN(n10681) );
  AOI21_X1 U11419 ( .B1(n10680), .B2(n10679), .A(n10681), .ZN(ADD_1068_U54) );
  AOI21_X1 U11420 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10681), .ZN(n10684) );
  NAND2_X1 U11421 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10682) );
  OAI21_X1 U11422 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10682), .ZN(n10683) );
  NOR2_X1 U11423 ( .A1(n10684), .A2(n10683), .ZN(n10685) );
  AOI21_X1 U11424 ( .B1(n10684), .B2(n10683), .A(n10685), .ZN(ADD_1068_U53) );
  AOI21_X1 U11425 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10685), .ZN(n10688) );
  NOR2_X1 U11426 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10686) );
  AOI21_X1 U11427 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10686), .ZN(n10687) );
  NAND2_X1 U11428 ( .A1(n10688), .A2(n10687), .ZN(n10690) );
  OAI21_X1 U11429 ( .B1(n10688), .B2(n10687), .A(n10690), .ZN(ADD_1068_U52) );
  NOR2_X1 U11430 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10689) );
  AOI21_X1 U11431 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10689), .ZN(n10692) );
  OAI21_X1 U11432 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10690), .ZN(n10691) );
  NAND2_X1 U11433 ( .A1(n10692), .A2(n10691), .ZN(n10694) );
  OAI21_X1 U11434 ( .B1(n10692), .B2(n10691), .A(n10694), .ZN(ADD_1068_U51) );
  NOR2_X1 U11435 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10693) );
  AOI21_X1 U11436 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10693), .ZN(n10696) );
  OAI21_X1 U11437 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10694), .ZN(n10695) );
  NAND2_X1 U11438 ( .A1(n10696), .A2(n10695), .ZN(n10698) );
  OAI21_X1 U11439 ( .B1(n10696), .B2(n10695), .A(n10698), .ZN(ADD_1068_U50) );
  NOR2_X1 U11440 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10697) );
  AOI21_X1 U11441 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10697), .ZN(n10700) );
  OAI21_X1 U11442 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10698), .ZN(n10699) );
  NAND2_X1 U11443 ( .A1(n10700), .A2(n10699), .ZN(n10702) );
  OAI21_X1 U11444 ( .B1(n10700), .B2(n10699), .A(n10702), .ZN(ADD_1068_U49) );
  NOR2_X1 U11445 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10701) );
  AOI21_X1 U11446 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10701), .ZN(n10704) );
  OAI21_X1 U11447 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10702), .ZN(n10703) );
  NAND2_X1 U11448 ( .A1(n10704), .A2(n10703), .ZN(n10706) );
  OAI21_X1 U11449 ( .B1(n10704), .B2(n10703), .A(n10706), .ZN(ADD_1068_U48) );
  NOR2_X1 U11450 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10705) );
  AOI21_X1 U11451 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10705), .ZN(n10708) );
  OAI21_X1 U11452 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10706), .ZN(n10707) );
  NAND2_X1 U11453 ( .A1(n10708), .A2(n10707), .ZN(n10710) );
  OAI21_X1 U11454 ( .B1(n10708), .B2(n10707), .A(n10710), .ZN(ADD_1068_U47) );
  NOR2_X1 U11455 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10709) );
  AOI21_X1 U11456 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10709), .ZN(n10712) );
  OAI21_X1 U11457 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10710), .ZN(n10711) );
  NAND2_X1 U11458 ( .A1(n10712), .A2(n10711), .ZN(n10714) );
  OAI21_X1 U11459 ( .B1(n10712), .B2(n10711), .A(n10714), .ZN(ADD_1068_U63) );
  NOR2_X1 U11460 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10713) );
  AOI21_X1 U11461 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10713), .ZN(n10716) );
  OAI21_X1 U11462 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10714), .ZN(n10715) );
  NAND2_X1 U11463 ( .A1(n10716), .A2(n10715), .ZN(n10718) );
  OAI21_X1 U11464 ( .B1(n10716), .B2(n10715), .A(n10718), .ZN(ADD_1068_U62) );
  NOR2_X1 U11465 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10717) );
  AOI21_X1 U11466 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10717), .ZN(n10720) );
  OAI21_X1 U11467 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10718), .ZN(n10719) );
  NAND2_X1 U11468 ( .A1(n10720), .A2(n10719), .ZN(n10722) );
  OAI21_X1 U11469 ( .B1(n10720), .B2(n10719), .A(n10722), .ZN(ADD_1068_U61) );
  NOR2_X1 U11470 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10721) );
  AOI21_X1 U11471 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10721), .ZN(n10724) );
  OAI21_X1 U11472 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10722), .ZN(n10723) );
  NAND2_X1 U11473 ( .A1(n10724), .A2(n10723), .ZN(n10726) );
  OAI21_X1 U11474 ( .B1(n10724), .B2(n10723), .A(n10726), .ZN(ADD_1068_U60) );
  NOR2_X1 U11475 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10725) );
  AOI21_X1 U11476 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10725), .ZN(n10728) );
  OAI21_X1 U11477 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10726), .ZN(n10727) );
  NAND2_X1 U11478 ( .A1(n10728), .A2(n10727), .ZN(n10730) );
  OAI21_X1 U11479 ( .B1(n10728), .B2(n10727), .A(n10730), .ZN(ADD_1068_U59) );
  NOR2_X1 U11480 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10729) );
  AOI21_X1 U11481 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10729), .ZN(n10732) );
  OAI21_X1 U11482 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10730), .ZN(n10731) );
  NAND2_X1 U11483 ( .A1(n10732), .A2(n10731), .ZN(n10734) );
  OAI21_X1 U11484 ( .B1(n10732), .B2(n10731), .A(n10734), .ZN(ADD_1068_U58) );
  NOR2_X1 U11485 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10733) );
  AOI21_X1 U11486 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10733), .ZN(n10736) );
  OAI21_X1 U11487 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10734), .ZN(n10735) );
  NAND2_X1 U11488 ( .A1(n10736), .A2(n10735), .ZN(n10738) );
  OAI21_X1 U11489 ( .B1(n10736), .B2(n10735), .A(n10738), .ZN(ADD_1068_U57) );
  NOR2_X1 U11490 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10737) );
  AOI21_X1 U11491 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10737), .ZN(n10740) );
  OAI21_X1 U11492 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10738), .ZN(n10739) );
  NAND2_X1 U11493 ( .A1(n10740), .A2(n10739), .ZN(n10742) );
  OAI21_X1 U11494 ( .B1(n10740), .B2(n10739), .A(n10742), .ZN(ADD_1068_U56) );
  INV_X1 U11495 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U11496 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .B1(n10833), .B2(n10741), .ZN(n10744) );
  OAI21_X1 U11497 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10742), .ZN(n10743) );
  NAND2_X1 U11498 ( .A1(n10744), .A2(n10743), .ZN(n10745) );
  OAI21_X1 U11499 ( .B1(n10744), .B2(n10743), .A(n10745), .ZN(ADD_1068_U55) );
  OAI21_X1 U11500 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10745), .ZN(n10747) );
  XOR2_X1 U11501 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n10746) );
  XNOR2_X1 U11502 ( .A(n10747), .B(n10746), .ZN(ADD_1068_U4) );
  MUX2_X1 U11503 ( .A(n10750), .B(n10749), .S(n10748), .Z(n10751) );
  NOR2_X1 U11504 ( .A1(n10751), .A2(n5124), .ZN(n10753) );
  XNOR2_X1 U11505 ( .A(n10753), .B(n10752), .ZN(n10757) );
  AOI22_X1 U11506 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10754), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10755) );
  OAI21_X1 U11507 ( .B1(n10757), .B2(n10756), .A(n10755), .ZN(P1_U3243) );
  INV_X1 U11508 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10772) );
  INV_X1 U11509 ( .A(n10758), .ZN(n10759) );
  OAI211_X1 U11510 ( .C1(n10761), .C2(n10760), .A(n10794), .B(n10759), .ZN(
        n10767) );
  INV_X1 U11511 ( .A(n10762), .ZN(n10763) );
  OAI211_X1 U11512 ( .C1(n10765), .C2(n10764), .A(n10822), .B(n10763), .ZN(
        n10766) );
  OAI211_X1 U11513 ( .C1(n10829), .C2(n10768), .A(n10767), .B(n10766), .ZN(
        n10769) );
  INV_X1 U11514 ( .A(n10769), .ZN(n10771) );
  OAI211_X1 U11515 ( .C1(n10862), .C2(n10772), .A(n10771), .B(n10770), .ZN(
        P1_U3251) );
  INV_X1 U11516 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10788) );
  INV_X1 U11517 ( .A(n10773), .ZN(n10784) );
  AOI21_X1 U11518 ( .B1(n10776), .B2(n10775), .A(n10774), .ZN(n10777) );
  NAND2_X1 U11519 ( .A1(n10794), .A2(n10777), .ZN(n10783) );
  AOI21_X1 U11520 ( .B1(n10780), .B2(n10779), .A(n10778), .ZN(n10781) );
  NAND2_X1 U11521 ( .A1(n10822), .A2(n10781), .ZN(n10782) );
  OAI211_X1 U11522 ( .C1(n10829), .C2(n10784), .A(n10783), .B(n10782), .ZN(
        n10785) );
  INV_X1 U11523 ( .A(n10785), .ZN(n10787) );
  NAND2_X1 U11524 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n10786)
         );
  OAI211_X1 U11525 ( .C1(n10862), .C2(n10788), .A(n10787), .B(n10786), .ZN(
        P1_U3254) );
  INV_X1 U11526 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10805) );
  INV_X1 U11527 ( .A(n10789), .ZN(n10801) );
  AOI21_X1 U11528 ( .B1(n10792), .B2(n10791), .A(n10790), .ZN(n10793) );
  NAND2_X1 U11529 ( .A1(n10794), .A2(n10793), .ZN(n10800) );
  AOI21_X1 U11530 ( .B1(n10797), .B2(n10796), .A(n10795), .ZN(n10798) );
  NAND2_X1 U11531 ( .A1(n10822), .A2(n10798), .ZN(n10799) );
  OAI211_X1 U11532 ( .C1(n10829), .C2(n10801), .A(n10800), .B(n10799), .ZN(
        n10802) );
  INV_X1 U11533 ( .A(n10802), .ZN(n10804) );
  OAI211_X1 U11534 ( .C1(n10862), .C2(n10805), .A(n10804), .B(n10803), .ZN(
        P1_U3257) );
  INV_X1 U11535 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10817) );
  AOI211_X1 U11536 ( .C1(n10808), .C2(n10807), .A(n10806), .B(n10847), .ZN(
        n10813) );
  AOI211_X1 U11537 ( .C1(n10811), .C2(n10810), .A(n10809), .B(n10851), .ZN(
        n10812) );
  AOI211_X1 U11538 ( .C1(n10858), .C2(n10814), .A(n10813), .B(n10812), .ZN(
        n10816) );
  OAI211_X1 U11539 ( .C1(n10862), .C2(n10817), .A(n10816), .B(n10815), .ZN(
        P1_U3258) );
  NOR2_X1 U11540 ( .A1(n10819), .A2(n10818), .ZN(n10820) );
  OR3_X1 U11541 ( .A1(n10821), .A2(n10820), .A3(n10851), .ZN(n10827) );
  OAI211_X1 U11542 ( .C1(n10825), .C2(n10824), .A(n10823), .B(n10822), .ZN(
        n10826) );
  OAI211_X1 U11543 ( .C1(n10829), .C2(n10828), .A(n10827), .B(n10826), .ZN(
        n10830) );
  INV_X1 U11544 ( .A(n10830), .ZN(n10832) );
  OAI211_X1 U11545 ( .C1(n10862), .C2(n10833), .A(n10832), .B(n10831), .ZN(
        P1_U3261) );
  INV_X1 U11546 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10846) );
  AOI211_X1 U11547 ( .C1(n10836), .C2(n10835), .A(n10834), .B(n10847), .ZN(
        n10841) );
  AOI211_X1 U11548 ( .C1(n10839), .C2(n10838), .A(n10837), .B(n10851), .ZN(
        n10840) );
  AOI211_X1 U11549 ( .C1(n10858), .C2(n10842), .A(n10841), .B(n10840), .ZN(
        n10845) );
  INV_X1 U11550 ( .A(n10843), .ZN(n10844) );
  OAI211_X1 U11551 ( .C1(n10862), .C2(n10846), .A(n10845), .B(n10844), .ZN(
        P1_U3256) );
  INV_X1 U11552 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10861) );
  AOI211_X1 U11553 ( .C1(n10850), .C2(n10849), .A(n10848), .B(n10847), .ZN(
        n10856) );
  AOI211_X1 U11554 ( .C1(n10854), .C2(n10853), .A(n10852), .B(n10851), .ZN(
        n10855) );
  AOI211_X1 U11555 ( .C1(n10858), .C2(n10857), .A(n10856), .B(n10855), .ZN(
        n10860) );
  OAI211_X1 U11556 ( .C1(n10862), .C2(n10861), .A(n10860), .B(n10859), .ZN(
        P1_U3253) );
  AOI22_X1 U11557 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n10906), .B1(n10907), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n10867) );
  XNOR2_X1 U11558 ( .A(n10863), .B(P2_IR_REG_0__SCAN_IN), .ZN(n10864) );
  OAI21_X1 U11559 ( .B1(n10865), .B2(n10923), .A(n10864), .ZN(n10866) );
  OAI211_X1 U11560 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10951), .A(n10867), .B(
        n10866), .ZN(P2_U3182) );
  OAI21_X1 U11561 ( .B1(n10869), .B2(n10868), .A(n10923), .ZN(n10871) );
  NOR2_X1 U11562 ( .A1(n10871), .A2(n10870), .ZN(n10879) );
  NOR2_X1 U11563 ( .A1(n10873), .A2(n10872), .ZN(n10874) );
  NOR2_X1 U11564 ( .A1(n10875), .A2(n10874), .ZN(n10877) );
  OAI22_X1 U11565 ( .A1(n10918), .A2(n10877), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10876), .ZN(n10878) );
  AOI211_X1 U11566 ( .C1(P2_ADDR_REG_2__SCAN_IN), .C2(n10907), .A(n10879), .B(
        n10878), .ZN(n10885) );
  AOI21_X1 U11567 ( .B1(n10882), .B2(n10881), .A(n10880), .ZN(n10883) );
  OR2_X1 U11568 ( .A1(n10915), .A2(n10883), .ZN(n10884) );
  OAI211_X1 U11569 ( .C1(n10904), .C2(n10886), .A(n10885), .B(n10884), .ZN(
        P2_U3184) );
  OAI21_X1 U11570 ( .B1(n10889), .B2(n10888), .A(n10887), .ZN(n10890) );
  AND2_X1 U11571 ( .A1(n10890), .A2(n10923), .ZN(n10900) );
  AOI21_X1 U11572 ( .B1(n10893), .B2(n10892), .A(n10891), .ZN(n10898) );
  AOI21_X1 U11573 ( .B1(n10896), .B2(n10895), .A(n10894), .ZN(n10897) );
  OAI22_X1 U11574 ( .A1(n10898), .A2(n10918), .B1(n10897), .B2(n10915), .ZN(
        n10899) );
  AOI211_X1 U11575 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n10907), .A(n10900), .B(
        n10899), .ZN(n10902) );
  NAND2_X1 U11576 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n10901) );
  OAI211_X1 U11577 ( .C1(n10904), .C2(n10903), .A(n10902), .B(n10901), .ZN(
        P2_U3188) );
  INV_X1 U11578 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U11579 ( .A1(n10907), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n10906), 
        .B2(n10905), .ZN(n10925) );
  OAI21_X1 U11580 ( .B1(n10910), .B2(n10909), .A(n10908), .ZN(n10922) );
  INV_X1 U11581 ( .A(n10911), .ZN(n10912) );
  AOI21_X1 U11582 ( .B1(n10913), .B2(n6536), .A(n10912), .ZN(n10914) );
  NOR2_X1 U11583 ( .A1(n10915), .A2(n10914), .ZN(n10921) );
  AOI21_X1 U11584 ( .B1(n10917), .B2(n6538), .A(n10916), .ZN(n10919) );
  NOR2_X1 U11585 ( .A1(n10919), .A2(n10918), .ZN(n10920) );
  AOI211_X1 U11586 ( .C1(n10923), .C2(n10922), .A(n10921), .B(n10920), .ZN(
        n10924) );
  OAI211_X1 U11587 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10926), .A(n10925), .B(
        n10924), .ZN(P2_U3193) );
  XNOR2_X1 U11588 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11589 ( .A(n10927), .ZN(n10931) );
  AOI21_X1 U11590 ( .B1(n11000), .B2(n10929), .A(n10928), .ZN(n10930) );
  AOI211_X1 U11591 ( .C1(n10933), .C2(n10932), .A(n10931), .B(n10930), .ZN(
        n10934) );
  AOI22_X1 U11592 ( .A1(n11116), .A2(n10934), .B1(n10749), .B2(n11115), .ZN(
        P1_U3522) );
  AOI22_X1 U11593 ( .A1(n11120), .A2(n10934), .B1(n5735), .B2(n11117), .ZN(
        P1_U3453) );
  OR2_X1 U11594 ( .A1(n11132), .A2(n10935), .ZN(n10936) );
  NAND2_X1 U11595 ( .A1(n10937), .A2(n10936), .ZN(n10940) );
  NAND2_X1 U11596 ( .A1(n11151), .A2(n10938), .ZN(n10939) );
  NAND2_X1 U11597 ( .A1(n10940), .A2(n10939), .ZN(n10953) );
  INV_X1 U11598 ( .A(n10941), .ZN(n10943) );
  NAND3_X1 U11599 ( .A1(n10953), .A2(n10943), .A3(n10942), .ZN(n10946) );
  AND2_X1 U11600 ( .A1(n6408), .A2(n10944), .ZN(n10952) );
  NAND2_X1 U11601 ( .A1(n11046), .A2(n10952), .ZN(n10945) );
  OAI211_X1 U11602 ( .C1(n11048), .C2(n10947), .A(n10946), .B(n10945), .ZN(
        n10948) );
  INV_X1 U11603 ( .A(n10948), .ZN(n10949) );
  OAI21_X1 U11604 ( .B1(n10951), .B2(n10950), .A(n10949), .ZN(P2_U3233) );
  NOR2_X1 U11605 ( .A1(n10953), .A2(n10952), .ZN(n10955) );
  AOI22_X1 U11606 ( .A1(n11153), .A2(n10955), .B1(n7320), .B2(n5476), .ZN(
        P2_U3459) );
  INV_X1 U11607 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U11608 ( .A1(n11157), .A2(n10955), .B1(n10954), .B2(n11154), .ZN(
        P2_U3390) );
  AOI22_X1 U11609 ( .A1(n10956), .A2(n11132), .B1(n11151), .B2(n6398), .ZN(
        n10958) );
  AND2_X1 U11610 ( .A1(n10958), .A2(n10957), .ZN(n10960) );
  AOI22_X1 U11611 ( .A1(n11153), .A2(n10960), .B1(n7323), .B2(n5476), .ZN(
        P2_U3460) );
  INV_X1 U11612 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U11613 ( .A1(n11157), .A2(n10960), .B1(n10959), .B2(n11154), .ZN(
        P2_U3393) );
  AOI22_X1 U11614 ( .A1(n11120), .A2(n10961), .B1(n5747), .B2(n11117), .ZN(
        P1_U3456) );
  XNOR2_X1 U11615 ( .A(n10962), .B(n10966), .ZN(n10975) );
  NOR2_X1 U11616 ( .A1(n10963), .A2(n11127), .ZN(n10971) );
  NAND3_X1 U11617 ( .A1(n8068), .A2(n10966), .A3(n10965), .ZN(n10968) );
  AOI21_X1 U11618 ( .B1(n10964), .B2(n10968), .A(n10967), .ZN(n10970) );
  OR2_X1 U11619 ( .A1(n10970), .A2(n10969), .ZN(n10978) );
  AOI211_X1 U11620 ( .C1(n10975), .C2(n11132), .A(n10971), .B(n10978), .ZN(
        n10973) );
  AOI22_X1 U11621 ( .A1(n11153), .A2(n10973), .B1(n7413), .B2(n5476), .ZN(
        P2_U3461) );
  INV_X1 U11622 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U11623 ( .A1(n11157), .A2(n10973), .B1(n10972), .B2(n11154), .ZN(
        P2_U3396) );
  INV_X1 U11624 ( .A(n10974), .ZN(n10976) );
  AOI222_X1 U11625 ( .A1(n10977), .A2(n10976), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n11041), .C1(n11036), .C2(n10975), .ZN(n10980) );
  NOR2_X1 U11626 ( .A1(n10981), .A2(n10978), .ZN(n10979) );
  AOI22_X1 U11627 ( .A1(n7414), .A2(n10981), .B1(n10980), .B2(n10979), .ZN(
        P2_U3231) );
  NOR2_X1 U11628 ( .A1(n10982), .A2(n11127), .ZN(n10984) );
  AOI211_X1 U11629 ( .C1(n10985), .C2(n11132), .A(n10984), .B(n10983), .ZN(
        n10987) );
  AOI22_X1 U11630 ( .A1(n11153), .A2(n10987), .B1(n6421), .B2(n5476), .ZN(
        P2_U3462) );
  INV_X1 U11631 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U11632 ( .A1(n11157), .A2(n10987), .B1(n10986), .B2(n11154), .ZN(
        P2_U3399) );
  OAI22_X1 U11633 ( .A1(n10989), .A2(n11146), .B1(n10988), .B2(n11127), .ZN(
        n10990) );
  NOR2_X1 U11634 ( .A1(n10991), .A2(n10990), .ZN(n10993) );
  AOI22_X1 U11635 ( .A1(n11153), .A2(n10993), .B1(n6434), .B2(n5476), .ZN(
        P2_U3463) );
  INV_X1 U11636 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U11637 ( .A1(n11157), .A2(n10993), .B1(n10992), .B2(n11154), .ZN(
        P2_U3402) );
  AOI21_X1 U11638 ( .B1(n10996), .B2(n10995), .A(n10994), .ZN(n10997) );
  OAI211_X1 U11639 ( .C1(n11000), .C2(n10999), .A(n10998), .B(n10997), .ZN(
        n11001) );
  INV_X1 U11640 ( .A(n11001), .ZN(n11003) );
  AOI22_X1 U11641 ( .A1(n11116), .A2(n11003), .B1(n11002), .B2(n11115), .ZN(
        P1_U3526) );
  AOI22_X1 U11642 ( .A1(n11120), .A2(n11003), .B1(n5808), .B2(n11117), .ZN(
        P1_U3465) );
  NOR2_X1 U11643 ( .A1(n11004), .A2(n11127), .ZN(n11006) );
  AOI211_X1 U11644 ( .C1(n11008), .C2(n11007), .A(n11006), .B(n11005), .ZN(
        n11010) );
  AOI22_X1 U11645 ( .A1(n11153), .A2(n11010), .B1(n6445), .B2(n5476), .ZN(
        P2_U3464) );
  INV_X1 U11646 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U11647 ( .A1(n11157), .A2(n11010), .B1(n11009), .B2(n11154), .ZN(
        P2_U3405) );
  INV_X1 U11648 ( .A(n11011), .ZN(n11024) );
  OAI22_X1 U11649 ( .A1(n11015), .A2(n11014), .B1(n11013), .B2(n11012), .ZN(
        n11016) );
  AOI21_X1 U11650 ( .B1(n11018), .B2(n11017), .A(n11016), .ZN(n11019) );
  OAI21_X1 U11651 ( .B1(n11021), .B2(n11020), .A(n11019), .ZN(n11022) );
  AOI21_X1 U11652 ( .B1(n11024), .B2(n11023), .A(n11022), .ZN(n11025) );
  OAI21_X1 U11653 ( .B1(n10529), .B2(n11026), .A(n11025), .ZN(P1_U3288) );
  INV_X1 U11654 ( .A(n11027), .ZN(n11028) );
  OAI21_X1 U11655 ( .B1(n11029), .B2(n11109), .A(n11028), .ZN(n11031) );
  AOI211_X1 U11656 ( .C1(n11054), .C2(n11032), .A(n11031), .B(n11030), .ZN(
        n11034) );
  AOI22_X1 U11657 ( .A1(n11116), .A2(n11034), .B1(n11033), .B2(n11115), .ZN(
        P1_U3528) );
  AOI22_X1 U11658 ( .A1(n11120), .A2(n11034), .B1(n5843), .B2(n11117), .ZN(
        P1_U3471) );
  INV_X1 U11659 ( .A(n11035), .ZN(n11039) );
  INV_X1 U11660 ( .A(n11036), .ZN(n11038) );
  OAI21_X1 U11661 ( .B1(n11039), .B2(n11038), .A(n11037), .ZN(n11045) );
  INV_X1 U11662 ( .A(n11040), .ZN(n11042) );
  AOI222_X1 U11663 ( .A1(n11046), .A2(n11045), .B1(n11044), .B2(n11043), .C1(
        n11042), .C2(n11041), .ZN(n11047) );
  OAI21_X1 U11664 ( .B1(n11048), .B2(n6476), .A(n11047), .ZN(P2_U3226) );
  OAI22_X1 U11665 ( .A1(n11050), .A2(n11049), .B1(n5253), .B2(n11109), .ZN(
        n11052) );
  AOI211_X1 U11666 ( .C1(n11054), .C2(n11053), .A(n11052), .B(n11051), .ZN(
        n11056) );
  AOI22_X1 U11667 ( .A1(n11116), .A2(n11056), .B1(n5883), .B2(n11115), .ZN(
        P1_U3530) );
  INV_X1 U11668 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U11669 ( .A1(n11120), .A2(n11056), .B1(n11055), .B2(n11117), .ZN(
        P1_U3477) );
  INV_X1 U11670 ( .A(n11057), .ZN(n11061) );
  OAI21_X1 U11671 ( .B1(n11059), .B2(n11127), .A(n11058), .ZN(n11060) );
  AOI21_X1 U11672 ( .B1(n11132), .B2(n11061), .A(n11060), .ZN(n11063) );
  AOI22_X1 U11673 ( .A1(n11153), .A2(n11063), .B1(n6492), .B2(n5476), .ZN(
        P2_U3467) );
  INV_X1 U11674 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U11675 ( .A1(n11157), .A2(n11063), .B1(n11062), .B2(n11154), .ZN(
        P2_U3414) );
  OAI21_X1 U11676 ( .B1(n11065), .B2(n11109), .A(n11064), .ZN(n11067) );
  AOI211_X1 U11677 ( .C1(n11113), .C2(n11068), .A(n11067), .B(n11066), .ZN(
        n11070) );
  AOI22_X1 U11678 ( .A1(n11116), .A2(n11070), .B1(n5906), .B2(n11115), .ZN(
        P1_U3531) );
  INV_X1 U11679 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U11680 ( .A1(n11120), .A2(n11070), .B1(n11069), .B2(n11117), .ZN(
        P1_U3480) );
  NOR2_X1 U11681 ( .A1(n11072), .A2(n11071), .ZN(n11074) );
  AOI211_X1 U11682 ( .C1(n11151), .C2(n11075), .A(n11074), .B(n11073), .ZN(
        n11077) );
  AOI22_X1 U11683 ( .A1(n11153), .A2(n11077), .B1(n8427), .B2(n5476), .ZN(
        P2_U3469) );
  INV_X1 U11684 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U11685 ( .A1(n11157), .A2(n11077), .B1(n11076), .B2(n11154), .ZN(
        P2_U3420) );
  AOI22_X1 U11686 ( .A1(n11079), .A2(n11132), .B1(n11151), .B2(n11078), .ZN(
        n11080) );
  AND2_X1 U11687 ( .A1(n11081), .A2(n11080), .ZN(n11083) );
  AOI22_X1 U11688 ( .A1(n11153), .A2(n11083), .B1(n6536), .B2(n5476), .ZN(
        P2_U3470) );
  INV_X1 U11689 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U11690 ( .A1(n11157), .A2(n11083), .B1(n11082), .B2(n11154), .ZN(
        P2_U3423) );
  NAND2_X1 U11691 ( .A1(n11086), .A2(n11085), .ZN(n11087) );
  XNOR2_X1 U11692 ( .A(n11084), .B(n11087), .ZN(n11098) );
  NAND2_X1 U11693 ( .A1(n11089), .A2(n11088), .ZN(n11093) );
  AOI22_X1 U11694 ( .A1(n11091), .A2(n11090), .B1(P1_REG3_REG_11__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11092) );
  OAI211_X1 U11695 ( .C1(n11095), .C2(n11094), .A(n11093), .B(n11092), .ZN(
        n11096) );
  AOI21_X1 U11696 ( .B1(n11098), .B2(n11097), .A(n11096), .ZN(n11099) );
  OAI21_X1 U11697 ( .B1(n11101), .B2(n11100), .A(n11099), .ZN(P1_U3236) );
  NOR2_X1 U11698 ( .A1(n11102), .A2(n11146), .ZN(n11104) );
  AOI211_X1 U11699 ( .C1(n11151), .C2(n11105), .A(n11104), .B(n11103), .ZN(
        n11107) );
  AOI22_X1 U11700 ( .A1(n11153), .A2(n11107), .B1(n8500), .B2(n5476), .ZN(
        P2_U3471) );
  INV_X1 U11701 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U11702 ( .A1(n11157), .A2(n11107), .B1(n11106), .B2(n11154), .ZN(
        P2_U3426) );
  OAI21_X1 U11703 ( .B1(n11110), .B2(n11109), .A(n11108), .ZN(n11111) );
  AOI211_X1 U11704 ( .C1(n11114), .C2(n11113), .A(n11112), .B(n11111), .ZN(
        n11119) );
  AOI22_X1 U11705 ( .A1(n11116), .A2(n11119), .B1(n5959), .B2(n11115), .ZN(
        P1_U3534) );
  INV_X1 U11706 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U11707 ( .A1(n11120), .A2(n11119), .B1(n11118), .B2(n11117), .ZN(
        P1_U3489) );
  AND2_X1 U11708 ( .A1(n11121), .A2(n11132), .ZN(n11123) );
  AOI211_X1 U11709 ( .C1(n11151), .C2(n11124), .A(n11123), .B(n11122), .ZN(
        n11126) );
  AOI22_X1 U11710 ( .A1(n11153), .A2(n11126), .B1(n8506), .B2(n5476), .ZN(
        P2_U3472) );
  INV_X1 U11711 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11125) );
  AOI22_X1 U11712 ( .A1(n11157), .A2(n11126), .B1(n11125), .B2(n11154), .ZN(
        P2_U3429) );
  NOR2_X1 U11713 ( .A1(n11128), .A2(n11127), .ZN(n11130) );
  AOI211_X1 U11714 ( .C1(n11132), .C2(n11131), .A(n11130), .B(n11129), .ZN(
        n11134) );
  AOI22_X1 U11715 ( .A1(n11153), .A2(n11134), .B1(n6573), .B2(n5476), .ZN(
        P2_U3473) );
  INV_X1 U11716 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U11717 ( .A1(n11157), .A2(n11134), .B1(n11133), .B2(n11154), .ZN(
        P2_U3432) );
  NOR2_X1 U11718 ( .A1(n11135), .A2(n11146), .ZN(n11136) );
  AOI211_X1 U11719 ( .C1(n11151), .C2(n11138), .A(n11137), .B(n11136), .ZN(
        n11140) );
  AOI22_X1 U11720 ( .A1(n11153), .A2(n11140), .B1(n8599), .B2(n5476), .ZN(
        P2_U3474) );
  INV_X1 U11721 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U11722 ( .A1(n11157), .A2(n11140), .B1(n11139), .B2(n11154), .ZN(
        P2_U3435) );
  NOR2_X1 U11723 ( .A1(n11141), .A2(n11146), .ZN(n11143) );
  AOI211_X1 U11724 ( .C1(n11151), .C2(n11144), .A(n11143), .B(n11142), .ZN(
        n11145) );
  AOI22_X1 U11725 ( .A1(n11153), .A2(n11145), .B1(n8592), .B2(n5476), .ZN(
        P2_U3475) );
  AOI22_X1 U11726 ( .A1(n11157), .A2(n11145), .B1(n6602), .B2(n11154), .ZN(
        P2_U3438) );
  NOR2_X1 U11727 ( .A1(n11147), .A2(n11146), .ZN(n11149) );
  AOI211_X1 U11728 ( .C1(n11151), .C2(n11150), .A(n11149), .B(n11148), .ZN(
        n11156) );
  AOI22_X1 U11729 ( .A1(n11153), .A2(n11156), .B1(n11152), .B2(n5476), .ZN(
        P2_U3476) );
  INV_X1 U11730 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n11155) );
  AOI22_X1 U11731 ( .A1(n11157), .A2(n11156), .B1(n11155), .B2(n11154), .ZN(
        P2_U3441) );
  XNOR2_X1 U11732 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X1 U5187 ( .A(n7121), .Z(n5118) );
  CLKBUF_X1 U5202 ( .A(n5789), .Z(n8649) );
  CLKBUF_X2 U5215 ( .A(n6311), .Z(n5124) );
  XNOR2_X1 U5289 ( .A(n8580), .B(n9371), .ZN(n9358) );
  CLKBUF_X3 U6477 ( .A(n6854), .Z(n6847) );
endmodule

