

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2971, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803;

  INV_X1 U3419 ( .A(n6311), .ZN(n6299) );
  INV_X1 U3420 ( .A(n5600), .ZN(n5565) );
  AND2_X1 U3421 ( .A1(n6096), .A2(n6075), .ZN(n6116) );
  OAI21_X1 U3422 ( .B1(n4496), .B2(n3919), .A(n4622), .ZN(n6452) );
  NAND2_X2 U3423 ( .A1(n3502), .A2(n3503), .ZN(n3535) );
  INV_X2 U3424 ( .A(n6802), .ZN(n5377) );
  CLKBUF_X2 U3426 ( .A(n3311), .Z(n4108) );
  CLKBUF_X2 U3427 ( .A(n3273), .Z(n4112) );
  INV_X2 U3428 ( .A(n2975), .ZN(n4561) );
  INV_X1 U3429 ( .A(n3289), .ZN(n3247) );
  AND2_X2 U3430 ( .A1(n3148), .A2(n4449), .ZN(n3339) );
  CLKBUF_X2 U3432 ( .A(n3326), .Z(n3494) );
  AND4_X1 U3433 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3371)
         );
  OR2_X1 U3434 ( .A1(n4244), .A2(n3282), .ZN(n4257) );
  NOR2_X1 U3435 ( .A1(n5565), .A2(n3074), .ZN(n5553) );
  OR2_X1 U3436 ( .A1(n6452), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3070)
         );
  INV_X1 U3438 ( .A(n4026), .ZN(n4081) );
  NOR2_X1 U3439 ( .A1(n5593), .A2(n5590), .ZN(n5579) );
  INV_X1 U3440 ( .A(n5214), .ZN(n5610) );
  INV_X1 U3441 ( .A(n6259), .ZN(n6303) );
  NAND2_X1 U3442 ( .A1(n3429), .A2(n3428), .ZN(n4316) );
  XNOR2_X1 U3443 ( .A(n4160), .B(n4159), .ZN(n5918) );
  NOR2_X1 U3444 ( .A1(n5938), .A2(n5912), .ZN(n5935) );
  INV_X1 U34450 ( .A(n6305), .ZN(n6260) );
  INV_X1 U34460 ( .A(n6266), .ZN(n6282) );
  XNOR2_X1 U34470 ( .A(n4152), .B(n4151), .ZN(n5254) );
  OR2_X1 U34480 ( .A1(n4392), .A2(n4964), .ZN(n6161) );
  NOR2_X4 U3449 ( .A1(n5307), .A2(n5309), .ZN(n5294) );
  NAND2_X2 U3450 ( .A1(n5360), .A2(n3132), .ZN(n5307) );
  NAND2_X2 U34510 ( .A1(n5029), .A2(n5200), .ZN(n5214) );
  AND2_X1 U34520 ( .A1(n4449), .A2(n3011), .ZN(n2971) );
  OAI21_X2 U34530 ( .B1(n4081), .B2(EBX_REG_1__SCAN_IN), .A(n4000), .ZN(n4001)
         );
  AND2_X4 U3454 ( .A1(n5190), .A2(n4451), .ZN(n3341) );
  AND2_X1 U34550 ( .A1(n3073), .A2(n2998), .ZN(n5552) );
  NAND2_X1 U34560 ( .A1(n5232), .A2(n5231), .ZN(n3045) );
  OR2_X1 U3457 ( .A1(n2983), .A2(n4131), .ZN(n4137) );
  NAND2_X1 U3458 ( .A1(n4316), .A2(n4317), .ZN(n4315) );
  INV_X1 U34590 ( .A(n3535), .ZN(n3047) );
  INV_X1 U34610 ( .A(n4077), .ZN(n4016) );
  INV_X1 U34620 ( .A(n3383), .ZN(n4535) );
  NAND2_X1 U34630 ( .A1(n3299), .A2(n3140), .ZN(n3384) );
  INV_X2 U34650 ( .A(n3288), .ZN(n3358) );
  NAND2_X2 U3466 ( .A1(n3356), .A2(n3355), .ZN(n3031) );
  NAND4_X1 U3467 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n3998)
         );
  AND4_X1 U34680 ( .A1(n3325), .A2(n3324), .A3(n3323), .A4(n3322), .ZN(n3337)
         );
  AND4_X1 U34690 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3336)
         );
  AND4_X1 U34700 ( .A1(n3321), .A2(n3320), .A3(n3319), .A4(n3318), .ZN(n3338)
         );
  BUF_X2 U34710 ( .A(n3340), .Z(n4109) );
  BUF_X2 U34720 ( .A(n3342), .Z(n3819) );
  BUF_X2 U34730 ( .A(n3343), .Z(n3818) );
  BUF_X2 U34740 ( .A(n3341), .Z(n3838) );
  BUF_X2 U3475 ( .A(n3431), .Z(n4110) );
  CLKBUF_X2 U3476 ( .A(n3349), .Z(n4103) );
  OAI21_X1 U3477 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5621), .A(n5611), 
        .ZN(n5612) );
  NOR2_X1 U3478 ( .A1(n5552), .A2(n3077), .ZN(n5237) );
  AND2_X1 U3479 ( .A1(n3073), .A2(n5236), .ZN(n2991) );
  NAND2_X1 U3480 ( .A1(n3010), .A2(n3081), .ZN(n5602) );
  NAND2_X1 U3481 ( .A1(n5825), .A2(n5824), .ZN(n5823) );
  NOR2_X1 U3482 ( .A1(n4147), .A2(n4146), .ZN(n4148) );
  AND2_X1 U3483 ( .A1(n3061), .A2(n3033), .ZN(n3032) );
  NAND2_X1 U3484 ( .A1(n3136), .A2(n3009), .ZN(n6425) );
  AOI21_X1 U3485 ( .B1(n3086), .B2(n3091), .A(n3082), .ZN(n3081) );
  NAND2_X1 U3486 ( .A1(n6435), .A2(n6434), .ZN(n3046) );
  OAI21_X1 U3487 ( .B1(n3067), .B2(n3056), .A(n2994), .ZN(n3062) );
  AND2_X1 U3488 ( .A1(n3087), .A2(n3089), .ZN(n3082) );
  NAND2_X1 U3489 ( .A1(n5019), .A2(n5018), .ZN(n6435) );
  AND2_X1 U3490 ( .A1(n2988), .A2(n5225), .ZN(n3066) );
  AOI21_X1 U3491 ( .B1(n6311), .B2(n5559), .A(n4096), .ZN(n4097) );
  XNOR2_X1 U3492 ( .A(n5214), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5832)
         );
  NAND2_X1 U3493 ( .A1(n3609), .A2(n3608), .ZN(n4798) );
  NAND2_X1 U3494 ( .A1(n4137), .A2(n5377), .ZN(n4157) );
  AND2_X2 U3495 ( .A1(n5248), .A2(n3997), .ZN(n6311) );
  XNOR2_X1 U3496 ( .A(n5029), .B(n3601), .ZN(n5201) );
  NAND2_X1 U3497 ( .A1(n4315), .A2(n3507), .ZN(n4428) );
  AND2_X1 U3498 ( .A1(n4626), .A2(n4625), .ZN(n6453) );
  CLKBUF_X1 U3499 ( .A(n4496), .Z(n6551) );
  NAND2_X1 U3500 ( .A1(n3019), .A2(n3534), .ZN(n4516) );
  NAND2_X1 U3501 ( .A1(n5349), .A2(n5350), .ZN(n5334) );
  NAND2_X1 U3502 ( .A1(n4343), .A2(n3471), .ZN(n4317) );
  CLKBUF_X1 U3503 ( .A(n5349), .Z(n5363) );
  AND2_X1 U3505 ( .A1(n3465), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4345) );
  CLKBUF_X1 U3506 ( .A(n4492), .Z(n4870) );
  NAND2_X1 U3507 ( .A1(n3528), .A2(n3527), .ZN(n4520) );
  NAND2_X1 U3508 ( .A1(n3464), .A2(n3463), .ZN(n4492) );
  NAND2_X1 U3509 ( .A1(n3460), .A2(n3418), .ZN(n3421) );
  OAI21_X1 U3510 ( .B1(n4460), .B2(STATE2_REG_0__SCAN_IN), .A(n3501), .ZN(
        n3503) );
  NAND2_X1 U3511 ( .A1(n3466), .A2(n4488), .ZN(n3460) );
  NOR2_X2 U3512 ( .A1(n4845), .A2(n5045), .ZN(n5174) );
  NOR2_X1 U3513 ( .A1(n6392), .A2(n4561), .ZN(n6359) );
  NAND2_X1 U3514 ( .A1(n3410), .A2(n3411), .ZN(n3485) );
  NAND2_X1 U3515 ( .A1(n3394), .A2(n3393), .ZN(n3410) );
  NAND2_X1 U3516 ( .A1(n3397), .A2(n3396), .ZN(n3411) );
  AOI22_X1 U3517 ( .A1(n5377), .A2(n5465), .B1(n4077), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4340) );
  NAND2_X1 U3518 ( .A1(n4077), .A2(n5377), .ZN(n4342) );
  NAND2_X1 U3519 ( .A1(n4240), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3370) );
  INV_X1 U3520 ( .A(n4509), .ZN(n4513) );
  AND2_X2 U3521 ( .A1(n3363), .A2(n4400), .ZN(n3921) );
  NAND2_X2 U3522 ( .A1(n4535), .A2(n2976), .ZN(n4077) );
  CLKBUF_X1 U3523 ( .A(n4087), .Z(n5216) );
  INV_X1 U3524 ( .A(n3031), .ZN(n3380) );
  INV_X2 U3525 ( .A(n3384), .ZN(n2974) );
  AND4_X1 U3526 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3299)
         );
  AND4_X1 U3527 ( .A1(n3354), .A2(n3353), .A3(n3352), .A4(n3351), .ZN(n3355)
         );
  BUF_X2 U3528 ( .A(n3350), .Z(n4102) );
  AND4_X1 U3529 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3335)
         );
  AND2_X1 U3530 ( .A1(n3022), .A2(n3021), .ZN(n3315) );
  AND4_X1 U3531 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3279)
         );
  AND4_X1 U3532 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3280)
         );
  AND4_X1 U3533 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3278)
         );
  AND4_X1 U3534 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3281)
         );
  AND4_X1 U3535 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(n3235)
         );
  AND2_X1 U3536 ( .A1(n3250), .A2(n3249), .ZN(n3251) );
  AND4_X1 U3537 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3236)
         );
  AND4_X1 U3538 ( .A1(n3348), .A2(n3347), .A3(n3346), .A4(n3345), .ZN(n3356)
         );
  BUF_X2 U3539 ( .A(n3344), .Z(n3448) );
  BUF_X2 U3540 ( .A(n3430), .Z(n4101) );
  BUF_X2 U3541 ( .A(n3339), .Z(n3836) );
  BUF_X2 U3542 ( .A(n4111), .Z(n3837) );
  OR2_X2 U3543 ( .A1(n6137), .A2(STATE_REG_2__SCAN_IN), .ZN(n4215) );
  AND2_X4 U3544 ( .A1(n4451), .A2(n4480), .ZN(n3349) );
  BUF_X2 U3545 ( .A(n3998), .Z(n2975) );
  BUF_X4 U3546 ( .A(n3998), .Z(n2976) );
  AND2_X4 U3547 ( .A1(n3011), .A2(n4480), .ZN(n3431) );
  NOR2_X1 U3548 ( .A1(n3048), .A2(n3535), .ZN(n3578) );
  OAI21_X2 U3549 ( .B1(n5269), .B2(n5271), .A(n5270), .ZN(n5571) );
  NAND3_X2 U3550 ( .A1(n4431), .A2(n3357), .A3(n4513), .ZN(n4269) );
  NOR2_X2 U3551 ( .A1(n5334), .A2(n5335), .ZN(n5322) );
  NOR2_X4 U3552 ( .A1(n4575), .A2(n3595), .ZN(n4760) );
  XNOR2_X1 U3553 ( .A(n4291), .B(n4290), .ZN(n4446) );
  AOI211_X2 U3554 ( .C1(n5939), .C2(n5570), .A(n5569), .B(n5568), .ZN(n5946)
         );
  AND2_X1 U3555 ( .A1(n3001), .A2(n5321), .ZN(n3132) );
  NAND2_X1 U3556 ( .A1(n5823), .A2(n5229), .ZN(n5232) );
  NAND2_X1 U3557 ( .A1(n4386), .A2(n6750), .ZN(n4392) );
  AND2_X1 U3558 ( .A1(n3590), .A2(n3589), .ZN(n3597) );
  NOR2_X1 U3559 ( .A1(n3123), .A2(n3122), .ZN(n3121) );
  INV_X1 U3560 ( .A(n5180), .ZN(n3120) );
  INV_X1 U3561 ( .A(n5512), .ZN(n3122) );
  NAND2_X1 U3562 ( .A1(n5600), .A2(n2980), .ZN(n3073) );
  NAND2_X1 U3563 ( .A1(n5297), .A2(n5284), .ZN(n3096) );
  NAND2_X1 U3564 ( .A1(n3093), .A2(n3080), .ZN(n3079) );
  NOR2_X1 U3565 ( .A1(n5620), .A2(n5910), .ZN(n3092) );
  AND3_X1 U3566 ( .A1(n2974), .A2(n4535), .A3(n3358), .ZN(n4319) );
  NAND2_X1 U3567 ( .A1(n3017), .A2(n3385), .ZN(n3969) );
  NAND2_X1 U3568 ( .A1(n6132), .A2(n4487), .ZN(n4529) );
  AND2_X1 U3569 ( .A1(n4475), .A2(n4474), .ZN(n4959) );
  NAND2_X1 U3570 ( .A1(n4278), .A2(n4277), .ZN(n4507) );
  OR2_X1 U3571 ( .A1(n4392), .A2(n3964), .ZN(n4298) );
  AND2_X1 U3572 ( .A1(n4686), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4149) );
  AND2_X1 U3573 ( .A1(n3126), .A2(n3128), .ZN(n3125) );
  INV_X1 U3574 ( .A(n3903), .ZN(n3126) );
  INV_X1 U3575 ( .A(n5374), .ZN(n3020) );
  NAND2_X1 U3576 ( .A1(n5647), .A2(n5606), .ZN(n3055) );
  NAND2_X1 U3577 ( .A1(n5657), .A2(n5653), .ZN(n5647) );
  INV_X1 U3578 ( .A(n3062), .ZN(n3061) );
  NAND2_X1 U3579 ( .A1(n3064), .A2(n3034), .ZN(n3033) );
  OR3_X1 U3580 ( .A1(n4392), .A2(n4391), .A3(n3384), .ZN(n4393) );
  NAND2_X1 U3581 ( .A1(n3023), .A2(n4432), .ZN(n3914) );
  NAND2_X1 U3582 ( .A1(n3954), .A2(n3031), .ZN(n3023) );
  AND2_X1 U3583 ( .A1(n2976), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3363) );
  AND2_X1 U3584 ( .A1(n6626), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3925)
         );
  AND2_X1 U3585 ( .A1(n5706), .A2(n3939), .ZN(n3941) );
  NAND2_X1 U3586 ( .A1(n3599), .A2(n3598), .ZN(n5029) );
  INV_X1 U3587 ( .A(n3597), .ZN(n3598) );
  OR2_X1 U3588 ( .A1(n3454), .A2(n3453), .ZN(n5215) );
  NAND2_X1 U3589 ( .A1(n3398), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3489) );
  OAI211_X1 U3590 ( .C1(n3969), .C2(n3014), .A(n3013), .B(n4401), .ZN(n3359)
         );
  NAND2_X1 U3591 ( .A1(n3044), .A2(n2990), .ZN(n3013) );
  AOI21_X1 U3592 ( .B1(n3379), .B2(n4257), .A(n4535), .ZN(n3391) );
  NOR2_X1 U3593 ( .A1(n3900), .A2(n5573), .ZN(n3028) );
  NAND2_X1 U3594 ( .A1(n3130), .A2(n5295), .ZN(n3129) );
  INV_X1 U3595 ( .A(n5282), .ZN(n3130) );
  NOR2_X1 U3596 ( .A1(n5348), .A2(n3134), .ZN(n3133) );
  INV_X1 U3597 ( .A(n5362), .ZN(n3134) );
  INV_X1 U3598 ( .A(n5173), .ZN(n3114) );
  AND2_X1 U3599 ( .A1(n3646), .A2(n3625), .ZN(n3115) );
  INV_X1 U3600 ( .A(n5043), .ZN(n3646) );
  INV_X1 U3601 ( .A(n4840), .ZN(n3625) );
  INV_X1 U3602 ( .A(n3602), .ZN(n3607) );
  AND2_X1 U3603 ( .A1(n4512), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3548) );
  NOR2_X1 U3604 ( .A1(n5610), .A2(n5939), .ZN(n3078) );
  AOI21_X1 U3605 ( .B1(n3090), .B2(n3088), .A(n5610), .ZN(n3086) );
  AOI21_X1 U3606 ( .B1(n5233), .B2(n3088), .A(n3005), .ZN(n3087) );
  INV_X1 U3607 ( .A(n5233), .ZN(n3089) );
  NAND2_X1 U3608 ( .A1(n3085), .A2(n3084), .ZN(n3083) );
  INV_X1 U3609 ( .A(n3087), .ZN(n3084) );
  INV_X1 U3610 ( .A(n3086), .ZN(n3085) );
  NOR2_X1 U3611 ( .A1(n3052), .A2(n3036), .ZN(n3035) );
  INV_X1 U3612 ( .A(n3053), .ZN(n3052) );
  INV_X1 U3613 ( .A(n5606), .ZN(n3051) );
  INV_X1 U3614 ( .A(n3106), .ZN(n3104) );
  INV_X1 U3615 ( .A(n4059), .ZN(n3105) );
  NOR2_X1 U3616 ( .A1(n5639), .A2(n3054), .ZN(n3053) );
  INV_X1 U3617 ( .A(n5608), .ZN(n3054) );
  NOR2_X1 U3618 ( .A1(n4305), .A2(n4256), .ZN(n4407) );
  INV_X1 U3619 ( .A(n5208), .ZN(n5210) );
  NOR2_X1 U3620 ( .A1(n6423), .A2(n3060), .ZN(n3059) );
  INV_X1 U3621 ( .A(n5028), .ZN(n3060) );
  INV_X1 U3622 ( .A(n5433), .ZN(n3099) );
  OR2_X1 U3623 ( .A1(n3408), .A2(n3407), .ZN(n4618) );
  INV_X1 U3624 ( .A(n4370), .ZN(n3514) );
  AND2_X1 U3625 ( .A1(n3007), .A2(n3484), .ZN(n3486) );
  NAND2_X1 U3626 ( .A1(n3029), .A2(n3485), .ZN(n3007) );
  NAND4_X1 U3627 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(n3301)
         );
  OR2_X1 U3628 ( .A1(n3462), .A2(n3461), .ZN(n3463) );
  NAND2_X1 U3629 ( .A1(n3460), .A2(n3459), .ZN(n3464) );
  INV_X1 U3630 ( .A(n5216), .ZN(n6796) );
  OR2_X1 U3631 ( .A1(n5435), .A2(n4088), .ZN(n4093) );
  OR2_X1 U3632 ( .A1(n6794), .A2(n3978), .ZN(n6233) );
  INV_X2 U3633 ( .A(n2984), .ZN(n4395) );
  AND2_X1 U3634 ( .A1(n3385), .A2(n3289), .ZN(n4512) );
  NAND2_X1 U3635 ( .A1(n3692), .A2(n3124), .ZN(n3123) );
  INV_X1 U3636 ( .A(n5548), .ZN(n3124) );
  NAND2_X1 U3637 ( .A1(n3028), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4126)
         );
  AND2_X1 U3638 ( .A1(n3117), .A2(n2982), .ZN(n3116) );
  INV_X1 U3639 ( .A(n5484), .ZN(n3117) );
  CLKBUF_X1 U3640 ( .A(n5360), .Z(n5361) );
  NAND2_X1 U3641 ( .A1(n3740), .A2(n3003), .ZN(n3785) );
  NOR2_X1 U3642 ( .A1(n3733), .A2(n6208), .ZN(n3740) );
  INV_X1 U3643 ( .A(n5689), .ZN(n3738) );
  NAND2_X1 U3644 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n3718), .ZN(n3733)
         );
  CLKBUF_X1 U3645 ( .A(n5510), .Z(n5511) );
  OR2_X1 U3646 ( .A1(n4344), .A2(n3976), .ZN(n3471) );
  INV_X1 U3647 ( .A(n5234), .ZN(n3076) );
  AND2_X1 U3648 ( .A1(n4076), .A2(n4075), .ZN(n5284) );
  NOR3_X1 U3649 ( .A1(n5323), .A2(n3096), .A3(n5311), .ZN(n5286) );
  NAND2_X1 U3650 ( .A1(n5600), .A2(n3079), .ZN(n5593) );
  NAND2_X1 U3651 ( .A1(n5322), .A2(n5324), .ZN(n5323) );
  NAND2_X1 U3652 ( .A1(n5487), .A2(n3107), .ZN(n3106) );
  INV_X1 U3653 ( .A(n5394), .ZN(n3107) );
  AND2_X1 U3654 ( .A1(n3039), .A2(n5233), .ZN(n3037) );
  INV_X1 U3655 ( .A(n4443), .ZN(n6081) );
  NAND2_X1 U3656 ( .A1(n2988), .A2(n3057), .ZN(n3067) );
  INV_X1 U3657 ( .A(n5227), .ZN(n3057) );
  NAND2_X1 U3658 ( .A1(n5222), .A2(n5221), .ZN(n5836) );
  NAND2_X1 U3659 ( .A1(n3008), .A2(n6453), .ZN(n3071) );
  NAND3_X1 U3660 ( .A1(n3069), .A2(n3068), .A3(n4641), .ZN(n3072) );
  NOR2_X1 U3661 ( .A1(n3969), .A2(n3968), .ZN(n4279) );
  OR2_X1 U3662 ( .A1(n3967), .A2(n3966), .ZN(n3968) );
  NOR2_X1 U3663 ( .A1(n4803), .A2(n4849), .ZN(n4807) );
  AND3_X1 U3664 ( .A1(n6780), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6627) );
  OR2_X1 U3665 ( .A1(n6551), .A2(n4520), .ZN(n4803) );
  AND2_X1 U3666 ( .A1(n4855), .A2(n4685), .ZN(n5056) );
  AND2_X1 U3667 ( .A1(n5050), .A2(n2977), .ZN(n6681) );
  OR2_X1 U3668 ( .A1(n4764), .A2(n4870), .ZN(n5047) );
  NOR2_X1 U3669 ( .A1(n6551), .A2(n4579), .ZN(n4584) );
  AND2_X1 U3670 ( .A1(n6550), .A2(n6774), .ZN(n4588) );
  INV_X1 U3671 ( .A(n6624), .ZN(n4765) );
  AND2_X1 U3672 ( .A1(n4529), .A2(n4488), .ZN(n4855) );
  AND2_X1 U3673 ( .A1(n4581), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4684)
         );
  OR2_X1 U3674 ( .A1(n6551), .A2(n4521), .ZN(n4531) );
  INV_X1 U3675 ( .A(n3011), .ZN(n4478) );
  NAND2_X1 U3676 ( .A1(n3961), .A2(n3960), .ZN(n3962) );
  AOI21_X1 U3677 ( .B1(n3949), .B2(n3948), .A(n3947), .ZN(n3958) );
  NAND2_X1 U3678 ( .A1(n6160), .A2(n4686), .ZN(n3976) );
  OR2_X1 U3679 ( .A1(n4269), .A2(n6796), .ZN(n4973) );
  INV_X1 U3680 ( .A(n4167), .ZN(n3101) );
  AND2_X1 U3681 ( .A1(n6233), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6306) );
  OAI21_X1 U3682 ( .B1(n4507), .B2(n4506), .A(n6750), .ZN(n4508) );
  INV_X1 U3683 ( .A(n6406), .ZN(n6409) );
  AOI22_X1 U3684 ( .A1(n4150), .A2(EAX_REG_31__SCAN_IN), .B1(n4149), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4151) );
  OAI21_X1 U3685 ( .B1(n4128), .B2(n4129), .A(n4152), .ZN(n5243) );
  AND2_X1 U3686 ( .A1(n6050), .A2(n6016), .ZN(n6033) );
  INV_X1 U3687 ( .A(n6534), .ZN(n6121) );
  INV_X1 U3688 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6626) );
  INV_X1 U3689 ( .A(n6778), .ZN(n6781) );
  NAND2_X1 U3690 ( .A1(n4807), .A2(n4870), .ZN(n6634) );
  NAND2_X1 U3691 ( .A1(n4727), .A2(n4870), .ZN(n5058) );
  NAND2_X1 U3692 ( .A1(n4584), .A2(n4870), .ZN(n4690) );
  INV_X1 U3693 ( .A(n3967), .ZN(n3016) );
  AOI22_X1 U3694 ( .A1(n3431), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3232) );
  AOI22_X1 U3695 ( .A1(n3339), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3228) );
  AND2_X1 U3696 ( .A1(n3556), .A2(n3577), .ZN(n3049) );
  OR2_X1 U3697 ( .A1(n3588), .A2(n3587), .ZN(n5203) );
  OR2_X1 U3698 ( .A1(n3567), .A2(n3566), .ZN(n5032) );
  OR2_X1 U3699 ( .A1(n3545), .A2(n3544), .ZN(n5021) );
  OR2_X1 U3700 ( .A1(n3500), .A2(n3499), .ZN(n4620) );
  NAND2_X1 U3701 ( .A1(n3415), .A2(n3031), .ZN(n3365) );
  OAI21_X1 U3702 ( .B1(n4244), .B2(n4400), .A(n3385), .ZN(n4249) );
  INV_X1 U3703 ( .A(n4246), .ZN(n3361) );
  CLKBUF_X1 U3704 ( .A(n4246), .Z(n4247) );
  AOI21_X1 U3705 ( .B1(n3350), .B2(INSTQUEUE_REG_2__2__SCAN_IN), .A(n3006), 
        .ZN(n3291) );
  AND2_X1 U3706 ( .A1(n3342), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3006) );
  NAND2_X1 U3707 ( .A1(n3350), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3022) );
  NAND2_X1 U3708 ( .A1(n3342), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3021) );
  AOI22_X1 U3709 ( .A1(n3349), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U3710 ( .A1(n3326), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3431), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U3711 ( .A1(n4111), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3244) );
  OR2_X1 U3712 ( .A1(n3526), .A2(n3525), .ZN(n4649) );
  AOI21_X1 U3713 ( .B1(n4243), .B2(n3913), .A(n3058), .ZN(n3912) );
  INV_X1 U3714 ( .A(n3363), .ZN(n3058) );
  NAND2_X1 U3715 ( .A1(n3302), .A2(n3398), .ZN(n4246) );
  NAND2_X1 U3716 ( .A1(n3953), .A2(n3952), .ZN(n3972) );
  AND2_X1 U3717 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6546), .ZN(n3950)
         );
  NAND2_X1 U3718 ( .A1(n3945), .A2(n3944), .ZN(n3974) );
  INV_X1 U3719 ( .A(n4269), .ZN(n3044) );
  NAND2_X1 U3720 ( .A1(n3350), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3322) );
  NAND2_X1 U3721 ( .A1(n3273), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U3722 ( .A1(n3342), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3254) );
  AND2_X1 U3723 ( .A1(n3477), .A2(n3476), .ZN(n3507) );
  AND2_X1 U3724 ( .A1(n3380), .A2(n2976), .ZN(n4087) );
  NOR2_X1 U3725 ( .A1(n3131), .A2(n3129), .ZN(n3128) );
  INV_X1 U3726 ( .A(n5271), .ZN(n3131) );
  OR2_X1 U3727 ( .A1(n3206), .A2(n3205), .ZN(n3884) );
  NOR2_X1 U3728 ( .A1(n3868), .A2(n5615), .ZN(n3027) );
  INV_X1 U3729 ( .A(n4124), .ZN(n3893) );
  INV_X1 U3730 ( .A(n5498), .ZN(n3119) );
  AND2_X1 U3731 ( .A1(n3693), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3718)
         );
  INV_X1 U3732 ( .A(n4839), .ZN(n3626) );
  XNOR2_X1 U3733 ( .A(n3557), .B(n3556), .ZN(n4648) );
  INV_X1 U3734 ( .A(n5221), .ZN(n3034) );
  INV_X1 U3735 ( .A(n5832), .ZN(n3056) );
  AND2_X1 U3736 ( .A1(n5199), .A2(n3920), .ZN(n5200) );
  NOR2_X1 U3737 ( .A1(n5517), .A2(n3109), .ZN(n3108) );
  INV_X1 U3738 ( .A(n3110), .ZN(n3109) );
  NOR2_X1 U3739 ( .A1(n3111), .A2(n5186), .ZN(n3110) );
  INV_X1 U3740 ( .A(n5175), .ZN(n3111) );
  NAND2_X1 U3741 ( .A1(n2984), .A2(n5377), .ZN(n4083) );
  OR2_X1 U3742 ( .A1(n3443), .A2(n3442), .ZN(n4619) );
  AND2_X1 U3743 ( .A1(n3457), .A2(n4618), .ZN(n3409) );
  AND2_X2 U3744 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U3745 ( .A1(n3483), .A2(n3482), .ZN(n3487) );
  AOI21_X1 U3746 ( .B1(n3478), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3373), 
        .ZN(n3041) );
  INV_X1 U3747 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4852) );
  INV_X1 U3748 ( .A(n5452), .ZN(n4722) );
  OR2_X1 U3749 ( .A1(n3933), .A2(n3932), .ZN(n3948) );
  AND2_X1 U3750 ( .A1(n3946), .A2(n3974), .ZN(n3947) );
  NAND2_X1 U3751 ( .A1(n3921), .A2(n3920), .ZN(n3959) );
  INV_X1 U3752 ( .A(n3959), .ZN(n3961) );
  INV_X1 U3753 ( .A(n3972), .ZN(n3960) );
  NOR2_X1 U3754 ( .A1(n3991), .A2(n6199), .ZN(n5382) );
  NOR2_X1 U3755 ( .A1(n6216), .A2(n6217), .ZN(n6192) );
  NAND2_X1 U3756 ( .A1(n6319), .A2(n3990), .ZN(n6216) );
  INV_X1 U3757 ( .A(n3395), .ZN(n3396) );
  INV_X1 U3758 ( .A(n3392), .ZN(n3393) );
  NAND2_X1 U3759 ( .A1(n3095), .A2(n5273), .ZN(n3094) );
  INV_X1 U3760 ( .A(n5311), .ZN(n3095) );
  OR2_X1 U3761 ( .A1(n2985), .A2(n5491), .ZN(n5493) );
  NAND2_X1 U3762 ( .A1(n4642), .A2(n3424), .ZN(n3019) );
  OR2_X1 U3763 ( .A1(n2987), .A2(n5583), .ZN(n3900) );
  INV_X1 U3764 ( .A(n3028), .ZN(n3904) );
  INV_X1 U3765 ( .A(n3129), .ZN(n3127) );
  NAND2_X1 U3766 ( .A1(n3027), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3882)
         );
  OR2_X1 U3767 ( .A1(n3856), .A2(n5626), .ZN(n3868) );
  INV_X1 U3768 ( .A(n3027), .ZN(n3879) );
  NOR2_X1 U3769 ( .A1(n3817), .A2(n5642), .ZN(n3851) );
  INV_X1 U3770 ( .A(n3855), .ZN(n5348) );
  INV_X1 U3771 ( .A(n3785), .ZN(n3286) );
  OR2_X1 U3772 ( .A1(n3801), .A2(n5650), .ZN(n3817) );
  AND2_X1 U3773 ( .A1(n3740), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3768)
         );
  AND2_X1 U3774 ( .A1(n3675), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3693)
         );
  AND2_X1 U3775 ( .A1(n3671), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3675)
         );
  AND2_X1 U3776 ( .A1(n3657), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3671)
         );
  AND3_X1 U3777 ( .A1(n3660), .A2(n3659), .A3(n3658), .ZN(n5173) );
  CLKBUF_X1 U3778 ( .A(n5171), .Z(n5172) );
  NAND2_X1 U3779 ( .A1(n3026), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3627)
         );
  INV_X1 U3780 ( .A(n3620), .ZN(n3026) );
  NOR2_X1 U3781 ( .A1(n3627), .A2(n5728), .ZN(n3657) );
  AND2_X1 U3782 ( .A1(n3645), .A2(n3644), .ZN(n5043) );
  AND3_X1 U3783 ( .A1(n3624), .A2(n3623), .A3(n3622), .ZN(n4840) );
  NOR2_X1 U3784 ( .A1(n3591), .A2(n3285), .ZN(n3603) );
  INV_X1 U3785 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3285) );
  NAND2_X1 U3786 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n3603), .ZN(n3620)
         );
  NOR2_X1 U3787 ( .A1(n3607), .A2(n3606), .ZN(n3608) );
  NOR2_X1 U3788 ( .A1(n3605), .A2(n3976), .ZN(n3606) );
  AND2_X1 U3789 ( .A1(n3529), .A2(n3024), .ZN(n3571) );
  NOR2_X1 U3790 ( .A1(n3025), .A2(n4657), .ZN(n3024) );
  INV_X1 U3791 ( .A(n3472), .ZN(n3529) );
  NAND2_X1 U3792 ( .A1(n3529), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3550)
         );
  NAND2_X1 U3793 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3472) );
  NOR2_X1 U3794 ( .A1(n3427), .A2(n3426), .ZN(n3428) );
  OAI21_X1 U3795 ( .B1(n4866), .B2(n3721), .A(n3470), .ZN(n4344) );
  NAND2_X1 U3796 ( .A1(n2980), .A2(n3078), .ZN(n3074) );
  OR2_X1 U3797 ( .A1(n5973), .A2(n5960), .ZN(n5938) );
  NAND2_X1 U3798 ( .A1(n5232), .A2(n3083), .ZN(n3010) );
  NAND2_X1 U3799 ( .A1(n2993), .A2(n3012), .ZN(n5621) );
  INV_X1 U3800 ( .A(n5630), .ZN(n3012) );
  AOI21_X1 U3801 ( .B1(n3053), .B2(n3051), .A(n2992), .ZN(n3050) );
  NAND2_X1 U3802 ( .A1(n5657), .A2(n3035), .ZN(n3038) );
  AND2_X1 U3803 ( .A1(n5174), .A2(n3108), .ZN(n6091) );
  OR2_X1 U3804 ( .A1(n6539), .A2(n6095), .ZN(n6108) );
  NAND2_X1 U3805 ( .A1(n5174), .A2(n5175), .ZN(n5185) );
  NAND2_X1 U3806 ( .A1(n3046), .A2(n3059), .ZN(n3009) );
  NAND2_X1 U3807 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  XNOR2_X1 U3808 ( .A(n5027), .B(n6502), .ZN(n6434) );
  INV_X1 U3809 ( .A(n4664), .ZN(n3098) );
  NAND2_X1 U3810 ( .A1(n4647), .A2(n6441), .ZN(n4655) );
  AND2_X1 U3811 ( .A1(n4423), .A2(n2979), .ZN(n5432) );
  INV_X1 U3812 ( .A(n6508), .ZN(n6531) );
  OR2_X1 U3813 ( .A1(n4411), .A2(n6508), .ZN(n4443) );
  NAND2_X1 U3814 ( .A1(n3516), .A2(n3515), .ZN(n4290) );
  INV_X1 U3815 ( .A(n4257), .ZN(n4948) );
  CLKBUF_X1 U3817 ( .A(n4460), .Z(n4461) );
  INV_X1 U3818 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4452) );
  AND2_X1 U3819 ( .A1(n4289), .A2(n4288), .ZN(n4954) );
  AOI21_X1 U3820 ( .B1(n4850), .B2(n6774), .A(n6776), .ZN(n4876) );
  AND2_X1 U3821 ( .A1(n4871), .A2(n4870), .ZN(n4983) );
  NAND2_X1 U3822 ( .A1(n4855), .A2(n4524), .ZN(n6558) );
  OR2_X1 U3823 ( .A1(n4642), .A2(n4848), .ZN(n6548) );
  INV_X1 U3824 ( .A(n4496), .ZN(n4848) );
  AND2_X1 U3825 ( .A1(n4804), .A2(n4831), .ZN(n4809) );
  NAND2_X1 U3826 ( .A1(n4642), .A2(n6551), .ZN(n6677) );
  OR2_X1 U3827 ( .A1(n4764), .A2(n4858), .ZN(n6547) );
  OR2_X1 U3828 ( .A1(n4461), .A2(n5452), .ZN(n6586) );
  XNOR2_X1 U3829 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U3830 ( .A1(n4529), .A2(n6766), .ZN(n4566) );
  OR2_X1 U3831 ( .A1(n6678), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4982) );
  INV_X1 U3832 ( .A(n6558), .ZN(n6687) );
  OR2_X1 U3833 ( .A1(n4282), .A2(n4243), .ZN(n4964) );
  AND2_X1 U3834 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n4490) );
  INV_X1 U3835 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4193) );
  INV_X1 U3836 ( .A(n5293), .ZN(n5278) );
  NAND2_X1 U3837 ( .A1(n5330), .A2(n3994), .ZN(n5293) );
  AND2_X1 U3838 ( .A1(n5358), .A2(n3993), .ZN(n5330) );
  AND2_X1 U3839 ( .A1(n5382), .A2(n3992), .ZN(n5358) );
  AND2_X1 U3840 ( .A1(n5391), .A2(n3983), .ZN(n5383) );
  INV_X1 U3841 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5728) );
  AOI21_X1 U3842 ( .B1(n5429), .B2(n4260), .A(n6266), .ZN(n6292) );
  INV_X1 U3843 ( .A(n5519), .ZN(n6331) );
  INV_X1 U3844 ( .A(n6335), .ZN(n5504) );
  AND2_X1 U3845 ( .A1(n4320), .A2(n6750), .ZN(n6335) );
  AND2_X1 U3846 ( .A1(n6354), .A2(n4513), .ZN(n6342) );
  NOR2_X1 U3847 ( .A1(n5180), .A2(n3123), .ZN(n5513) );
  INV_X1 U3848 ( .A(n6148), .ZN(n6351) );
  INV_X1 U3849 ( .A(n6354), .ZN(n6345) );
  OR2_X1 U3850 ( .A1(n6340), .A2(n6342), .ZN(n6350) );
  INV_X1 U3851 ( .A(n6350), .ZN(n6349) );
  NAND2_X2 U3852 ( .A1(n6354), .A2(n4511), .ZN(n6148) );
  NOR2_X1 U3853 ( .A1(n4950), .A2(n4302), .ZN(n4303) );
  OR2_X1 U3854 ( .A1(n4298), .A2(n4297), .ZN(n6406) );
  INV_X1 U3855 ( .A(n6418), .ZN(n6419) );
  XNOR2_X1 U3856 ( .A(n3907), .B(n3906), .ZN(n5248) );
  INV_X1 U3857 ( .A(n4126), .ZN(n3905) );
  INV_X1 U3858 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5626) );
  INV_X1 U3859 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U3860 ( .A1(n3118), .A2(n3116), .ZN(n5375) );
  AND2_X1 U3861 ( .A1(n3740), .A2(n3000), .ZN(n3770) );
  NAND2_X1 U3862 ( .A1(n4369), .A2(n6774), .ZN(n5886) );
  INV_X1 U3863 ( .A(n6161), .ZN(n6455) );
  INV_X1 U3864 ( .A(n5879), .ZN(n6450) );
  INV_X1 U3865 ( .A(n5886), .ZN(n6456) );
  NOR2_X1 U3866 ( .A1(n5565), .A2(n3075), .ZN(n3077) );
  NAND2_X1 U3867 ( .A1(n2980), .A2(n3002), .ZN(n3075) );
  INV_X1 U3868 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5939) );
  OR2_X1 U3869 ( .A1(n5286), .A2(n5285), .ZN(n5948) );
  NOR3_X1 U3870 ( .A1(n5393), .A2(n3106), .A3(n4059), .ZN(n5366) );
  NAND2_X1 U3871 ( .A1(n3055), .A2(n5608), .ZN(n5638) );
  NAND2_X1 U3872 ( .A1(n3045), .A2(n5233), .ZN(n5654) );
  NOR2_X1 U3873 ( .A1(n6067), .A2(n5908), .ZN(n6050) );
  NAND2_X1 U3874 ( .A1(n6464), .A2(n6055), .ZN(n6067) );
  NAND2_X1 U3875 ( .A1(n3063), .A2(n3067), .ZN(n5831) );
  NAND2_X1 U3876 ( .A1(n5836), .A2(n3066), .ZN(n3063) );
  INV_X1 U3877 ( .A(n6490), .ZN(n6120) );
  AND2_X2 U3878 ( .A1(n5260), .A2(n6748), .ZN(n6490) );
  INV_X1 U3879 ( .A(n3072), .ZN(n6444) );
  NAND2_X1 U3880 ( .A1(n3071), .A2(n3070), .ZN(n6443) );
  AND2_X1 U3881 ( .A1(n4410), .A2(n4402), .ZN(n6534) );
  INV_X1 U3882 ( .A(n3466), .ZN(n4866) );
  INV_X1 U3883 ( .A(n4870), .ZN(n4858) );
  INV_X1 U3885 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6160) );
  NAND2_X1 U3886 ( .A1(n6769), .A2(n4686), .ZN(n6678) );
  INV_X1 U3888 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6780) );
  INV_X1 U3889 ( .A(n4982), .ZN(n6776) );
  INV_X1 U3890 ( .A(n6678), .ZN(n6774) );
  INV_X1 U3891 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6546) );
  OR2_X1 U3892 ( .A1(n4489), .A2(n4855), .ZN(n6778) );
  INV_X1 U3893 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5264) );
  INV_X1 U3894 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4295) );
  AND2_X1 U3895 ( .A1(n4279), .A2(n3380), .ZN(n4482) );
  NOR2_X1 U3896 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5260) );
  OR2_X1 U3897 ( .A1(n4293), .A2(n6766), .ZN(n6135) );
  INV_X1 U3898 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4865) );
  INV_X1 U3899 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4918) );
  AND2_X1 U3900 ( .A1(n4871), .A2(n4858), .ZN(n4939) );
  NOR2_X2 U3901 ( .A1(n6548), .A2(n5047), .ZN(n6578) );
  NOR2_X2 U3902 ( .A1(n4806), .A2(n4870), .ZN(n6616) );
  NAND2_X1 U3903 ( .A1(n6633), .A2(n6632), .ZN(n6672) );
  AND2_X1 U3904 ( .A1(n4727), .A2(n4858), .ZN(n5125) );
  OAI211_X1 U3905 ( .C1(n5057), .C2(n6681), .A(n5056), .B(n5055), .ZN(n5080)
         );
  OR2_X1 U3906 ( .A1(n6677), .A2(n5047), .ZN(n6737) );
  INV_X1 U3907 ( .A(n6739), .ZN(n5123) );
  NOR2_X2 U3908 ( .A1(n4583), .A2(n4870), .ZN(n5120) );
  AOI22_X1 U3909 ( .A1(n4588), .A2(n4582), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5091), .ZN(n4615) );
  NAND2_X1 U3910 ( .A1(n4855), .A2(DATAI_1_), .ZN(n6699) );
  OR2_X1 U3911 ( .A1(n4566), .A2(n3380), .ZN(n5164) );
  NAND2_X1 U3912 ( .A1(n4855), .A2(DATAI_2_), .ZN(n6705) );
  OR2_X1 U3913 ( .A1(n4566), .A2(n2974), .ZN(n5137) );
  NAND2_X1 U3914 ( .A1(n4855), .A2(DATAI_3_), .ZN(n6711) );
  OR2_X1 U3915 ( .A1(n4566), .A2(n4535), .ZN(n5141) );
  NAND2_X1 U3916 ( .A1(n4855), .A2(DATAI_4_), .ZN(n6718) );
  OR2_X1 U3917 ( .A1(n4566), .A2(n3398), .ZN(n6712) );
  NAND2_X1 U3918 ( .A1(n4855), .A2(DATAI_6_), .ZN(n6733) );
  OR2_X1 U3919 ( .A1(n4566), .A2(n4541), .ZN(n5145) );
  NAND2_X1 U3920 ( .A1(n4855), .A2(DATAI_7_), .ZN(n6744) );
  OR2_X1 U3921 ( .A1(n4566), .A2(n5251), .ZN(n6735) );
  OAI21_X1 U3922 ( .B1(n4689), .B2(n4688), .A(n4687), .ZN(n4714) );
  INV_X1 U3923 ( .A(n4688), .ZN(n4721) );
  INV_X1 U3924 ( .A(n5158), .ZN(n6683) );
  NOR2_X2 U3925 ( .A1(n4531), .A2(n4858), .ZN(n4938) );
  NOR2_X1 U3926 ( .A1(n4531), .A2(n4870), .ZN(n4688) );
  NAND2_X1 U3927 ( .A1(n4386), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6132) );
  AND2_X1 U3928 ( .A1(n3963), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6750) );
  INV_X1 U3929 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6747) );
  NOR2_X1 U3930 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_0__SCAN_IN), .ZN(
        n6748) );
  INV_X1 U3931 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6769) );
  INV_X1 U3932 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4199) );
  OR2_X1 U3933 ( .A1(n6137), .A2(n4193), .ZN(n4203) );
  INV_X1 U3934 ( .A(n4203), .ZN(n4235) );
  OAI211_X1 U3935 ( .C1(n5254), .C2(n6282), .A(n3100), .B(n3102), .ZN(U2796)
         );
  NOR3_X1 U3936 ( .A1(n4163), .A2(n2989), .A3(n3101), .ZN(n3100) );
  NAND2_X1 U3937 ( .A1(n5918), .A2(n6305), .ZN(n3102) );
  NAND2_X1 U3938 ( .A1(n3139), .A2(n4145), .ZN(n4146) );
  INV_X1 U3939 ( .A(n3385), .ZN(n5251) );
  NAND2_X1 U3940 ( .A1(n3118), .A2(n2981), .ZN(n5389) );
  INV_X2 U3941 ( .A(n5610), .ZN(n3093) );
  NOR2_X1 U3942 ( .A1(n5180), .A2(n5516), .ZN(n2978) );
  AND2_X1 U3943 ( .A1(n5360), .A2(n3133), .ZN(n5332) );
  AND2_X1 U3944 ( .A1(n5360), .A2(n3001), .ZN(n5320) );
  NAND2_X1 U3945 ( .A1(n3626), .A2(n3115), .ZN(n5042) );
  NAND2_X1 U3946 ( .A1(n3626), .A2(n3625), .ZN(n4838) );
  INV_X1 U3947 ( .A(n5231), .ZN(n3088) );
  AND2_X1 U3948 ( .A1(n4422), .A2(n3099), .ZN(n2979) );
  AND2_X1 U3949 ( .A1(n4561), .A2(n3383), .ZN(n4254) );
  NAND2_X1 U3950 ( .A1(n3380), .A2(n4561), .ZN(n3910) );
  AND2_X1 U3951 ( .A1(n5294), .A2(n3125), .ZN(n4128) );
  AND2_X1 U3952 ( .A1(n3079), .A2(n3076), .ZN(n2980) );
  INV_X1 U3953 ( .A(n3301), .ZN(n3398) );
  INV_X1 U3954 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4657) );
  AND2_X1 U3955 ( .A1(n5390), .A2(n3119), .ZN(n2981) );
  AND2_X1 U3956 ( .A1(n3784), .A2(n2981), .ZN(n2982) );
  NAND2_X1 U3957 ( .A1(n5174), .A2(n3110), .ZN(n3112) );
  INV_X1 U3958 ( .A(n6229), .ZN(n6259) );
  OR3_X1 U3959 ( .A1(n5323), .A2(n3094), .A3(n3096), .ZN(n2983) );
  NAND2_X1 U3960 ( .A1(n3044), .A2(n2976), .ZN(n3964) );
  AND2_X4 U3961 ( .A1(n2976), .A2(n3031), .ZN(n2984) );
  INV_X1 U3962 ( .A(n3289), .ZN(n4541) );
  INV_X1 U3963 ( .A(n5499), .ZN(n3118) );
  OR2_X1 U3964 ( .A1(n5393), .A2(n5394), .ZN(n2985) );
  AND2_X1 U3965 ( .A1(n3118), .A2(n2982), .ZN(n2986) );
  NOR2_X1 U3966 ( .A1(n5323), .A2(n5311), .ZN(n5296) );
  NOR2_X1 U3967 ( .A1(n5506), .A2(n6064), .ZN(n5501) );
  NOR2_X1 U3968 ( .A1(n5499), .A2(n5498), .ZN(n5388) );
  OR2_X1 U3969 ( .A1(n3882), .A2(n3881), .ZN(n2987) );
  AND2_X2 U3970 ( .A1(n4451), .A2(n4449), .ZN(n3273) );
  OR2_X1 U3971 ( .A1(n5214), .A2(n6104), .ZN(n2988) );
  AND3_X1 U3972 ( .A1(n4164), .A2(REIP_REG_30__SCAN_IN), .A3(n4237), .ZN(n2989) );
  NAND2_X1 U3973 ( .A1(n5294), .A2(n3128), .ZN(n5270) );
  NAND2_X1 U3974 ( .A1(n5360), .A2(n5362), .ZN(n5346) );
  NAND2_X2 U3975 ( .A1(n5602), .A2(n5601), .ZN(n5600) );
  INV_X1 U3976 ( .A(n5322), .ZN(n5337) );
  AND2_X1 U3977 ( .A1(n3364), .A2(n2976), .ZN(n2990) );
  INV_X1 U3978 ( .A(n3091), .ZN(n3090) );
  NAND2_X1 U3979 ( .A1(n5233), .A2(n3092), .ZN(n3091) );
  AND2_X1 U3980 ( .A1(n3093), .A2(n6007), .ZN(n2992) );
  AND2_X1 U3981 ( .A1(n3055), .A2(n3053), .ZN(n2993) );
  INV_X1 U3982 ( .A(n3065), .ZN(n3064) );
  NAND2_X1 U3983 ( .A1(n3066), .A2(n5832), .ZN(n3065) );
  NAND2_X1 U3984 ( .A1(n5214), .A2(n6077), .ZN(n2994) );
  NOR3_X1 U3985 ( .A1(n5323), .A2(n5311), .A3(n3097), .ZN(n5283) );
  OR2_X1 U3986 ( .A1(n5393), .A2(n3106), .ZN(n2995) );
  NAND2_X1 U3987 ( .A1(n5171), .A2(n5181), .ZN(n5180) );
  AND2_X1 U3988 ( .A1(n3108), .A2(n6090), .ZN(n2996) );
  AND2_X1 U3989 ( .A1(n4616), .A2(n3098), .ZN(n2997) );
  AND2_X1 U3990 ( .A1(n5236), .A2(n5934), .ZN(n2998) );
  NAND2_X1 U3991 ( .A1(n3979), .A2(n4172), .ZN(n2999) );
  INV_X1 U3992 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n4488) );
  INV_X1 U3993 ( .A(n3467), .ZN(n3706) );
  INV_X1 U3994 ( .A(n3706), .ZN(n4150) );
  INV_X2 U3995 ( .A(n6332), .ZN(n5521) );
  NAND2_X1 U3996 ( .A1(n3511), .A2(n3510), .ZN(n4426) );
  AND3_X1 U3997 ( .A1(n4423), .A2(n2979), .A3(n2997), .ZN(n4662) );
  NAND2_X1 U3998 ( .A1(n4423), .A2(n4422), .ZN(n4424) );
  INV_X1 U3999 ( .A(n5653), .ZN(n3036) );
  AND2_X1 U4000 ( .A1(n5174), .A2(n2996), .ZN(n5507) );
  AND2_X1 U4001 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3000) );
  NAND2_X1 U4002 ( .A1(n3031), .A2(n3288), .ZN(n3919) );
  OR2_X1 U4003 ( .A1(n3289), .A2(n4686), .ZN(n3721) );
  AND2_X1 U4004 ( .A1(n3133), .A2(n3865), .ZN(n3001) );
  AND2_X1 U4005 ( .A1(n3078), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3002)
         );
  AND2_X1 U4006 ( .A1(n3000), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3003)
         );
  INV_X1 U4007 ( .A(n5297), .ZN(n3097) );
  NAND2_X1 U4008 ( .A1(n3116), .A2(n3020), .ZN(n3004) );
  NAND2_X1 U4009 ( .A1(n3115), .A2(n3114), .ZN(n3113) );
  INV_X1 U4010 ( .A(n3784), .ZN(n5490) );
  INV_X1 U4011 ( .A(n3910), .ZN(n4260) );
  INV_X1 U4012 ( .A(n5516), .ZN(n3692) );
  INV_X1 U4013 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3025) );
  NAND4_X1 U4014 ( .A1(n6022), .A2(n5978), .A3(n6007), .A4(n5997), .ZN(n3005)
         );
  AND2_X2 U4015 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3011) );
  INV_X1 U4016 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3080) );
  AND2_X2 U4017 ( .A1(n3150), .A2(n3148), .ZN(n3342) );
  AND2_X2 U4019 ( .A1(n3018), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3150)
         );
  NAND2_X1 U4020 ( .A1(n2974), .A2(n3383), .ZN(n3369) );
  NOR2_X1 U4021 ( .A1(n2974), .A2(n4541), .ZN(n3303) );
  NAND3_X1 U4022 ( .A1(n3007), .A2(n3484), .A3(n3487), .ZN(n4291) );
  NAND3_X1 U4023 ( .A1(n3071), .A2(n3070), .A3(n3072), .ZN(n6441) );
  NAND2_X1 U4024 ( .A1(n6452), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3008)
         );
  NAND2_X2 U4025 ( .A1(n3045), .A2(n3037), .ZN(n5657) );
  AND2_X2 U4026 ( .A1(n5190), .A2(n3011), .ZN(n3430) );
  AND2_X2 U4027 ( .A1(n3150), .A2(n3011), .ZN(n3326) );
  INV_X1 U4028 ( .A(n3415), .ZN(n3488) );
  NOR2_X1 U4029 ( .A1(n2975), .A2(n4488), .ZN(n3415) );
  AND2_X2 U4030 ( .A1(n3484), .A2(n3042), .ZN(n3029) );
  NAND2_X1 U4031 ( .A1(n3359), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3043) );
  NAND3_X1 U4032 ( .A1(n4260), .A2(n4319), .A3(n4512), .ZN(n4401) );
  NAND2_X1 U4033 ( .A1(n3016), .A2(n3015), .ZN(n3014) );
  AND2_X1 U4034 ( .A1(n3965), .A2(n3380), .ZN(n3015) );
  NAND2_X1 U4035 ( .A1(n3304), .A2(n3305), .ZN(n3017) );
  INV_X1 U4036 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3018) );
  XNOR2_X1 U4037 ( .A(n3535), .B(n4520), .ZN(n4642) );
  NOR2_X2 U4038 ( .A1(n5499), .A2(n3004), .ZN(n5360) );
  NOR2_X2 U4039 ( .A1(n4839), .A2(n3113), .ZN(n5171) );
  NAND2_X2 U4040 ( .A1(n3489), .A2(n3488), .ZN(n3954) );
  OAI21_X4 U4041 ( .B1(n3958), .B2(n3957), .A(n3962), .ZN(n4386) );
  INV_X2 U4042 ( .A(n6319), .ZN(n6289) );
  NOR2_X2 U4043 ( .A1(n5435), .A2(n3980), .ZN(n6319) );
  NAND4_X1 U4044 ( .A1(n3529), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .A3(
        PHYADDRPOINTER_REG_3__SCAN_IN), .A4(PHYADDRPOINTER_REG_4__SCAN_IN), 
        .ZN(n3591) );
  NOR2_X2 U4045 ( .A1(n5248), .A2(n3996), .ZN(n6266) );
  XNOR2_X1 U4046 ( .A(n3485), .B(n3029), .ZN(n4501) );
  NAND3_X1 U4047 ( .A1(n3356), .A2(n3355), .A3(n2999), .ZN(n3364) );
  NAND2_X1 U4048 ( .A1(n3031), .A2(n4380), .ZN(n4382) );
  NAND2_X1 U4049 ( .A1(n3031), .A2(n4179), .ZN(n4297) );
  NAND2_X1 U4050 ( .A1(n4561), .A2(n3031), .ZN(n5434) );
  AND2_X1 U4053 ( .A1(n4279), .A2(n3031), .ZN(n4950) );
  OAI21_X2 U4054 ( .B1(n5222), .B2(n3065), .A(n3032), .ZN(n5825) );
  NAND2_X1 U4055 ( .A1(n3038), .A2(n3050), .ZN(n5631) );
  INV_X1 U4056 ( .A(n5655), .ZN(n3039) );
  AND2_X2 U4057 ( .A1(n3150), .A2(n4451), .ZN(n3350) );
  NOR2_X4 U4058 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4451) );
  NAND3_X2 U4059 ( .A1(n3372), .A2(n3371), .A3(n3370), .ZN(n3478) );
  NAND2_X1 U4060 ( .A1(n3359), .A2(n3040), .ZN(n3042) );
  AND2_X1 U4061 ( .A1(n3360), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3040) );
  NAND2_X1 U4062 ( .A1(n3041), .A2(n3043), .ZN(n3484) );
  NAND2_X1 U4063 ( .A1(n3046), .A2(n5028), .ZN(n5212) );
  OAI21_X1 U4064 ( .B1(n6435), .B2(n6434), .A(n3046), .ZN(n6436) );
  NAND2_X1 U4065 ( .A1(n4520), .A2(n3556), .ZN(n3048) );
  NAND3_X1 U4066 ( .A1(n3047), .A2(n3049), .A3(n4520), .ZN(n3596) );
  NAND2_X1 U4067 ( .A1(n3047), .A2(n4520), .ZN(n3557) );
  NAND2_X1 U4068 ( .A1(n4632), .A2(n4520), .ZN(n3068) );
  NAND2_X1 U4069 ( .A1(n4639), .A2(n4638), .ZN(n3069) );
  NAND3_X1 U4070 ( .A1(n4423), .A2(n2979), .A3(n4616), .ZN(n4663) );
  NOR2_X2 U4071 ( .A1(n5393), .A2(n3103), .ZN(n5349) );
  NAND3_X1 U4072 ( .A1(n3105), .A2(n5365), .A3(n3104), .ZN(n3103) );
  INV_X1 U4073 ( .A(n3112), .ZN(n5184) );
  AND2_X2 U4074 ( .A1(n6802), .A2(n2984), .ZN(n4026) );
  NAND2_X1 U4075 ( .A1(n3120), .A2(n3121), .ZN(n5510) );
  AND2_X1 U4076 ( .A1(n5294), .A2(n3127), .ZN(n5269) );
  NAND2_X1 U4077 ( .A1(n5294), .A2(n5295), .ZN(n5281) );
  INV_X1 U4079 ( .A(n3381), .ZN(n3390) );
  OAI21_X1 U4080 ( .B1(n4100), .B2(n6282), .A(n4099), .ZN(U2798) );
  INV_X1 U4081 ( .A(n3410), .ZN(n3413) );
  AND2_X2 U4082 ( .A1(n3150), .A2(n3149), .ZN(n3340) );
  NAND2_X1 U4083 ( .A1(n3362), .A2(n4306), .ZN(n3381) );
  INV_X1 U4084 ( .A(n3504), .ZN(n3502) );
  NAND2_X1 U4085 ( .A1(n3419), .A2(n3421), .ZN(n3504) );
  NAND2_X1 U4086 ( .A1(n3594), .A2(n3593), .ZN(n4758) );
  AND2_X2 U4087 ( .A1(n3148), .A2(n5190), .ZN(n4111) );
  INV_X1 U4088 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4686) );
  NOR2_X1 U4089 ( .A1(n5501), .A2(n6065), .ZN(n3135) );
  AND2_X1 U4090 ( .A1(n6424), .A2(n5211), .ZN(n3136) );
  AND2_X1 U4091 ( .A1(n4541), .A2(n3385), .ZN(n3137) );
  AND2_X1 U4093 ( .A1(n4166), .A2(REIP_REG_30__SCAN_IN), .ZN(n3138) );
  AND2_X1 U4094 ( .A1(n4171), .A2(STATE_REG_1__SCAN_IN), .ZN(n4202) );
  OR2_X1 U4095 ( .A1(n6299), .A2(n5196), .ZN(n3139) );
  AND4_X1 U4096 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3140)
         );
  INV_X1 U4097 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5209) );
  INV_X1 U4098 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5787) );
  AND2_X1 U4099 ( .A1(n6392), .A2(n6791), .ZN(n6385) );
  AND3_X1 U4100 ( .A1(n3388), .A2(n6751), .A3(n4467), .ZN(n3389) );
  INV_X1 U4101 ( .A(n3577), .ZN(n3570) );
  OR2_X1 U4102 ( .A1(n3373), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3360)
         );
  NAND2_X1 U4103 ( .A1(n4400), .A2(n4541), .ZN(n3290) );
  OR2_X1 U4104 ( .A1(n3924), .A2(n3923), .ZN(n3931) );
  INV_X1 U4105 ( .A(n3411), .ZN(n3412) );
  INV_X1 U4106 ( .A(n3921), .ZN(n3946) );
  AOI22_X1 U4107 ( .A1(n3430), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3352) );
  INV_X1 U4108 ( .A(n3421), .ZN(n3422) );
  NAND2_X1 U4109 ( .A1(n3383), .A2(n4244), .ZN(n3382) );
  INV_X1 U4110 ( .A(n5333), .ZN(n3865) );
  NAND2_X1 U4111 ( .A1(n6780), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5706) );
  INV_X1 U4112 ( .A(n4576), .ZN(n3555) );
  OR2_X2 U4113 ( .A1(n3317), .A2(n3316), .ZN(n3383) );
  OR2_X1 U4114 ( .A1(n3951), .A2(n3950), .ZN(n3953) );
  OR3_X1 U4115 ( .A1(n3951), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6546), 
        .ZN(n3945) );
  NAND2_X1 U4116 ( .A1(n3286), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3801)
         );
  NAND2_X1 U4117 ( .A1(n3851), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3856)
         );
  AND2_X1 U4118 ( .A1(n4040), .A2(n4039), .ZN(n6090) );
  OR2_X1 U4119 ( .A1(n6588), .A2(n4866), .ZN(n4804) );
  INV_X1 U4120 ( .A(n6586), .ZN(n5094) );
  AND2_X1 U4121 ( .A1(n4279), .A2(n3975), .ZN(n4261) );
  AOI21_X1 U4122 ( .B1(n4164), .B2(n4222), .A(n3138), .ZN(n4145) );
  AND2_X1 U4123 ( .A1(n5300), .A2(n3989), .ZN(n5272) );
  INV_X1 U4124 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6208) );
  INV_X1 U4125 ( .A(n6306), .ZN(n6294) );
  NAND2_X1 U4126 ( .A1(n6233), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U4127 ( .A1(n4948), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4124) );
  INV_X1 U4128 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5615) );
  INV_X1 U4129 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5650) );
  AND3_X1 U4130 ( .A1(n3737), .A2(n3736), .A3(n3735), .ZN(n5689) );
  OR2_X1 U4131 ( .A1(n3093), .A2(n6032), .ZN(n5653) );
  NOR2_X1 U4132 ( .A1(n6548), .A2(n4849), .ZN(n4871) );
  AND2_X1 U4133 ( .A1(n3512), .A2(n4523), .ZN(n6585) );
  OR2_X1 U4134 ( .A1(n4461), .A2(n4722), .ZN(n6624) );
  NOR2_X1 U4135 ( .A1(n6677), .A2(n4849), .ZN(n4727) );
  AND2_X1 U4136 ( .A1(n4852), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6554)
         );
  INV_X1 U4137 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4580) );
  OR2_X1 U4138 ( .A1(n4566), .A2(n3358), .ZN(n6719) );
  AND2_X1 U4139 ( .A1(n6747), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3963) );
  NOR2_X1 U4140 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6797) );
  NOR2_X2 U4141 ( .A1(n4093), .A2(n4086), .ZN(n6305) );
  AND2_X1 U4142 ( .A1(n6354), .A2(n4512), .ZN(n6340) );
  INV_X1 U4143 ( .A(n4350), .ZN(n6416) );
  INV_X1 U4144 ( .A(n6461), .ZN(n5882) );
  NAND2_X1 U4145 ( .A1(n6161), .A2(n4371), .ZN(n5879) );
  OAI211_X1 U4146 ( .C1(n5557), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5556), .B(n6803), .ZN(n5558) );
  AND2_X1 U4147 ( .A1(n6033), .A2(n5909), .ZN(n5990) );
  INV_X1 U4148 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6007) );
  OR3_X1 U4149 ( .A1(n6110), .A2(n6100), .A3(n6082), .ZN(n6099) );
  NAND2_X1 U4150 ( .A1(n6108), .A2(n6079), .ZN(n6464) );
  AND2_X1 U4151 ( .A1(n4410), .A2(n4409), .ZN(n6508) );
  INV_X1 U4152 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6540) );
  INV_X1 U4153 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6074) );
  AND2_X1 U4154 ( .A1(n4410), .A2(n4399), .ZN(n6537) );
  OAI21_X1 U4155 ( .B1(n4876), .B2(n4875), .A(n4874), .ZN(n4899) );
  OAI211_X1 U4156 ( .C1(n4985), .C2(n4988), .A(n5056), .B(n5131), .ZN(n5010)
         );
  OAI21_X1 U4157 ( .B1(n6562), .B2(n6561), .A(n6560), .ZN(n6579) );
  INV_X1 U4158 ( .A(n6590), .ZN(n6614) );
  OAI211_X1 U4159 ( .C1(n6774), .C2(n6587), .A(n4810), .B(n6687), .ZN(n4833)
         );
  INV_X1 U4160 ( .A(n6634), .ZN(n6670) );
  OAI21_X1 U4161 ( .B1(n4770), .B2(n6627), .A(n6687), .ZN(n4794) );
  NOR2_X2 U4162 ( .A1(n4803), .A2(n6547), .ZN(n5167) );
  OAI211_X1 U4163 ( .C1(n6774), .C2(n5129), .A(n4731), .B(n6687), .ZN(n4754)
         );
  INV_X1 U4164 ( .A(n5058), .ZN(n5083) );
  INV_X1 U4165 ( .A(n6737), .ZN(n6729) );
  NOR2_X1 U4166 ( .A1(n6677), .A2(n6547), .ZN(n6739) );
  OAI211_X1 U4167 ( .C1(n6774), .C2(n5091), .A(n4589), .B(n6687), .ZN(n4612)
         );
  INV_X1 U4168 ( .A(DATAI_16_), .ZN(n5812) );
  INV_X1 U4169 ( .A(n4690), .ZN(n4718) );
  INV_X1 U4170 ( .A(n6641), .ZN(n6695) );
  INV_X1 U4171 ( .A(n6655), .ZN(n6715) );
  INV_X1 U4172 ( .A(n6676), .ZN(n6740) );
  INV_X1 U4173 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4171) );
  NAND2_X1 U4174 ( .A1(n4298), .A2(n4238), .ZN(n6794) );
  INV_X1 U4175 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6162) );
  NAND2_X1 U4176 ( .A1(n6406), .A2(n4508), .ZN(n6354) );
  NAND2_X1 U4177 ( .A1(n4490), .A2(n4488), .ZN(n6791) );
  INV_X1 U4178 ( .A(n6385), .ZN(n6369) );
  OR3_X1 U4179 ( .A1(n4392), .A2(n4303), .A3(n4380), .ZN(n6392) );
  OR2_X1 U4180 ( .A1(n4392), .A2(n4973), .ZN(n6418) );
  INV_X1 U4181 ( .A(n6420), .ZN(n4350) );
  NAND2_X1 U4182 ( .A1(n5879), .A2(n4656), .ZN(n6461) );
  INV_X1 U4183 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6063) );
  INV_X1 U4184 ( .A(n6537), .ZN(n6483) );
  NOR2_X1 U4185 ( .A1(n4857), .A2(n4856), .ZN(n4943) );
  AOI22_X1 U4186 ( .A1(n4869), .A2(n4875), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4868), .ZN(n4902) );
  INV_X1 U4187 ( .A(n4983), .ZN(n5016) );
  OR2_X1 U4188 ( .A1(n6548), .A2(n6547), .ZN(n6620) );
  AOI22_X1 U4189 ( .A1(n6589), .A2(n4805), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6587), .ZN(n4836) );
  OR2_X1 U4190 ( .A1(n4803), .A2(n5047), .ZN(n6675) );
  INV_X1 U4191 ( .A(n5125), .ZN(n5170) );
  AOI22_X1 U4192 ( .A1(n4730), .A2(n4726), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5129), .ZN(n4757) );
  AOI21_X1 U4193 ( .B1(n5053), .B2(n6681), .A(n5052), .ZN(n5086) );
  AOI22_X1 U4194 ( .A1(n6686), .A2(n6682), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6689), .ZN(n6745) );
  OR2_X1 U4195 ( .A1(n5886), .A2(n4536), .ZN(n6606) );
  NAND2_X1 U4196 ( .A1(n4855), .A2(DATAI_0_), .ZN(n6693) );
  NAND2_X1 U4197 ( .A1(n4855), .A2(DATAI_5_), .ZN(n6725) );
  OR2_X1 U4198 ( .A1(n5886), .A2(n4570), .ZN(n6641) );
  OR2_X1 U4199 ( .A1(n5886), .A2(n4543), .ZN(n6665) );
  AOI21_X1 U4200 ( .B1(n4526), .B2(n4528), .A(n4525), .ZN(n4574) );
  OR2_X1 U4201 ( .A1(n6158), .A2(n6769), .ZN(n4979) );
  INV_X1 U4202 ( .A(n6761), .ZN(n6765) );
  NAND2_X1 U4203 ( .A1(n4200), .A2(n6137), .ZN(n6761) );
  INV_X1 U4204 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6247) );
  OAI21_X1 U4205 ( .B1(n5243), .B2(n6282), .A(n4148), .ZN(U2797) );
  INV_X1 U4206 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3141) );
  AND2_X2 U4207 ( .A1(n3141), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3149)
         );
  INV_X1 U4208 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3142) );
  AND2_X2 U4209 ( .A1(n3142), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5190)
         );
  AND2_X2 U4210 ( .A1(n3149), .A2(n5190), .ZN(n3344) );
  INV_X1 U4211 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U4212 ( .A1(n3448), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3147) );
  AND2_X4 U4213 ( .A1(n3149), .A2(n4449), .ZN(n3436) );
  AOI22_X1 U4214 ( .A1(n3437), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3146) );
  NOR2_X4 U4215 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4480) );
  AOI22_X1 U4216 ( .A1(n3836), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4217 ( .A1(n3341), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3144) );
  NAND4_X1 U4218 ( .A1(n3147), .A2(n3146), .A3(n3145), .A4(n3144), .ZN(n3156)
         );
  AND2_X2 U4219 ( .A1(n3148), .A2(n4480), .ZN(n3343) );
  AOI22_X1 U4220 ( .A1(n4109), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4221 ( .A1(n4101), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3153) );
  AND2_X2 U4222 ( .A1(n3149), .A2(n4480), .ZN(n3311) );
  AOI22_X1 U4223 ( .A1(n4108), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4224 ( .A1(n3494), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3151) );
  NAND4_X1 U4225 ( .A1(n3154), .A2(n3153), .A3(n3152), .A4(n3151), .ZN(n3155)
         );
  NOR2_X1 U4226 ( .A1(n3156), .A2(n3155), .ZN(n3889) );
  AOI22_X1 U4227 ( .A1(n3837), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4228 ( .A1(n3494), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4229 ( .A1(n3448), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4230 ( .A1(n4103), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3157) );
  NAND4_X1 U4231 ( .A1(n3160), .A2(n3159), .A3(n3158), .A4(n3157), .ZN(n3166)
         );
  AOI22_X1 U4232 ( .A1(n3838), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4233 ( .A1(n4109), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4234 ( .A1(n3437), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4235 ( .A1(n3819), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3161) );
  NAND4_X1 U4236 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3165)
         );
  NOR2_X1 U4237 ( .A1(n3166), .A2(n3165), .ZN(n3875) );
  AOI22_X1 U4238 ( .A1(n3838), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4239 ( .A1(n3437), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4240 ( .A1(n3448), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4241 ( .A1(n3494), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3167) );
  NAND4_X1 U4242 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n3176)
         );
  AOI22_X1 U4243 ( .A1(n3837), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4244 ( .A1(n4109), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4245 ( .A1(n4101), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4246 ( .A1(n4112), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3171) );
  NAND4_X1 U4247 ( .A1(n3174), .A2(n3173), .A3(n3172), .A4(n3171), .ZN(n3175)
         );
  NOR2_X1 U4248 ( .A1(n3176), .A2(n3175), .ZN(n3858) );
  AOI22_X1 U4249 ( .A1(n4109), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4250 ( .A1(n3436), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4251 ( .A1(n3838), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4252 ( .A1(n3836), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3177) );
  NAND4_X1 U4253 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3186)
         );
  AOI22_X1 U4254 ( .A1(n3448), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4255 ( .A1(n4101), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4256 ( .A1(n3494), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4257 ( .A1(n4108), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3181) );
  NAND4_X1 U4258 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n3185)
         );
  NOR2_X1 U4259 ( .A1(n3186), .A2(n3185), .ZN(n3857) );
  OR2_X1 U4260 ( .A1(n3858), .A2(n3857), .ZN(n3867) );
  AOI22_X1 U4261 ( .A1(n3836), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3190) );
  INV_X1 U4262 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5810) );
  AOI22_X1 U4263 ( .A1(n3818), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3189) );
  AOI22_X1 U4264 ( .A1(n4101), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4265 ( .A1(n3837), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3187) );
  NAND4_X1 U4266 ( .A1(n3190), .A2(n3189), .A3(n3188), .A4(n3187), .ZN(n3196)
         );
  AOI22_X1 U4267 ( .A1(n3437), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4268 ( .A1(n3344), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4269 ( .A1(n4109), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U4270 ( .A1(n4112), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3191) );
  NAND4_X1 U4271 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .ZN(n3195)
         );
  NOR2_X1 U4272 ( .A1(n3196), .A2(n3195), .ZN(n3866) );
  OR2_X1 U4273 ( .A1(n3867), .A2(n3866), .ZN(n3874) );
  NOR2_X1 U4274 ( .A1(n3875), .A2(n3874), .ZN(n3885) );
  AOI22_X1 U4275 ( .A1(n3838), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4276 ( .A1(n4109), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4277 ( .A1(n3437), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U4278 ( .A1(n3819), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3197) );
  NAND4_X1 U4279 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n3197), .ZN(n3206)
         );
  AOI22_X1 U4280 ( .A1(n3837), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U4281 ( .A1(n3494), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3203) );
  AOI22_X1 U4282 ( .A1(n3448), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3202) );
  AOI22_X1 U4283 ( .A1(n4103), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3201) );
  NAND4_X1 U4284 ( .A1(n3204), .A2(n3203), .A3(n3202), .A4(n3201), .ZN(n3205)
         );
  NAND2_X1 U4285 ( .A1(n3885), .A2(n3884), .ZN(n3890) );
  NOR2_X1 U4286 ( .A1(n3889), .A2(n3890), .ZN(n3897) );
  AOI22_X1 U4287 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n3838), .B1(n4108), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4288 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n4109), .B1(n3818), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4289 ( .A1(n3437), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3208) );
  AOI22_X1 U4290 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n3819), .B1(n4102), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3207) );
  NAND4_X1 U4291 ( .A1(n3210), .A2(n3209), .A3(n3208), .A4(n3207), .ZN(n3216)
         );
  AOI22_X1 U4292 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n3837), .B1(n3836), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4293 ( .A1(n3494), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U4294 ( .A1(n3448), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4295 ( .A1(n4103), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3211) );
  NAND4_X1 U4296 ( .A1(n3214), .A2(n3213), .A3(n3212), .A4(n3211), .ZN(n3215)
         );
  OR2_X1 U4297 ( .A1(n3216), .A2(n3215), .ZN(n3896) );
  NAND2_X1 U4298 ( .A1(n3897), .A2(n3896), .ZN(n4119) );
  AOI22_X1 U4299 ( .A1(n4111), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4300 ( .A1(n3448), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4301 ( .A1(n3436), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4302 ( .A1(n3819), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3217) );
  NAND4_X1 U4303 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3226)
         );
  AOI22_X1 U4304 ( .A1(n4109), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3224) );
  AOI22_X1 U4305 ( .A1(n3494), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3223) );
  AOI22_X1 U4306 ( .A1(n3838), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3222) );
  AOI22_X1 U4307 ( .A1(n4112), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3221) );
  NAND4_X1 U4308 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .ZN(n3225)
         );
  NOR2_X1 U4309 ( .A1(n3226), .A2(n3225), .ZN(n4120) );
  XOR2_X1 U4310 ( .A(n4119), .B(n4120), .Z(n3284) );
  AOI22_X1 U4311 ( .A1(n3344), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4111), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3230) );
  AOI22_X1 U4312 ( .A1(n3436), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3229) );
  AOI22_X1 U4313 ( .A1(n3340), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U4314 ( .A1(n3342), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4315 ( .A1(n3341), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4316 ( .A1(n3343), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U4317 ( .A1(n3236), .A2(n3235), .ZN(n3288) );
  INV_X1 U4318 ( .A(n3358), .ZN(n3248) );
  AOI22_X1 U4319 ( .A1(n3341), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4320 ( .A1(n3340), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4321 ( .A1(n3436), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4322 ( .A1(n3342), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3237) );
  NAND4_X1 U4323 ( .A1(n3240), .A2(n3239), .A3(n3238), .A4(n3237), .ZN(n3246)
         );
  AOI22_X1 U4324 ( .A1(n3344), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3242) );
  NAND4_X1 U4325 ( .A1(n3244), .A2(n3243), .A3(n3242), .A4(n3241), .ZN(n3245)
         );
  NAND2_X4 U4327 ( .A1(n3248), .A2(n3247), .ZN(n4244) );
  AOI22_X1 U4328 ( .A1(n3436), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4329 ( .A1(n3344), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4111), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3252) );
  NAND2_X1 U4330 ( .A1(n3311), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3250) );
  NAND4_X1 U4331 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n3260)
         );
  AOI22_X1 U4332 ( .A1(n3341), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4333 ( .A1(n3326), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3431), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4334 ( .A1(n3340), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4335 ( .A1(n3339), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3255) );
  NAND4_X1 U4336 ( .A1(n3258), .A2(n3257), .A3(n3256), .A4(n3255), .ZN(n3259)
         );
  NAND2_X1 U4337 ( .A1(n3341), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3264) );
  NAND2_X1 U4338 ( .A1(n3311), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3263) );
  NAND2_X1 U4339 ( .A1(n3343), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3262) );
  NAND2_X1 U4340 ( .A1(n3340), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3261)
         );
  NAND2_X1 U4341 ( .A1(n3436), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3268)
         );
  NAND2_X1 U4342 ( .A1(n3430), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3267)
         );
  NAND2_X1 U4343 ( .A1(n3342), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U4344 ( .A1(n3350), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3265) );
  NAND2_X1 U4345 ( .A1(n4111), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3272) );
  NAND2_X1 U4346 ( .A1(n3339), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4347 ( .A1(n3326), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3270)
         );
  NAND2_X1 U4348 ( .A1(n3431), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3269)
         );
  NAND2_X1 U4349 ( .A1(n3344), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3277) );
  NAND2_X1 U4350 ( .A1(n3273), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4351 ( .A1(n3349), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4352 ( .A1(n3310), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3274)
         );
  NAND2_X1 U4353 ( .A1(n3385), .A2(n4400), .ZN(n3282) );
  NOR2_X2 U4354 ( .A1(n3385), .A2(n4686), .ZN(n3467) );
  INV_X1 U4355 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4363) );
  INV_X1 U4356 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5561) );
  OAI22_X1 U4357 ( .A1(n3706), .A2(n4363), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5561), .ZN(n3283) );
  AOI21_X1 U4358 ( .B1(n3284), .B2(n3893), .A(n3283), .ZN(n3287) );
  INV_X1 U4359 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3881) );
  INV_X1 U4360 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5583) );
  INV_X1 U4361 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5573) );
  XNOR2_X1 U4362 ( .A(n3904), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5559)
         );
  INV_X2 U4363 ( .A(n3976), .ZN(n3870) );
  MUX2_X1 U4364 ( .A(n3287), .B(n5559), .S(n3870), .Z(n3903) );
  NAND2_X1 U4365 ( .A1(n3358), .A2(n3289), .ZN(n3302) );
  NAND2_X1 U4366 ( .A1(n3290), .A2(n3302), .ZN(n3300) );
  AOI22_X1 U4367 ( .A1(n4111), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4368 ( .A1(n3430), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4369 ( .A1(n3339), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4370 ( .A1(n3340), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4371 ( .A1(n3344), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3431), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4372 ( .A1(n3436), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4373 ( .A1(n3273), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3295) );
  NAND2_X1 U4374 ( .A1(n3300), .A2(n2974), .ZN(n3305) );
  NAND2_X1 U4375 ( .A1(n3361), .A2(n3303), .ZN(n3304) );
  AOI22_X1 U4376 ( .A1(n3341), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4377 ( .A1(n3436), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4378 ( .A1(n3344), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4379 ( .A1(n3349), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3306) );
  NAND4_X1 U4380 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3317)
         );
  AOI22_X1 U4381 ( .A1(n4111), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4382 ( .A1(n3340), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4383 ( .A1(n3339), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3431), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3312) );
  NAND4_X1 U4384 ( .A1(n3315), .A2(n3314), .A3(n3313), .A4(n3312), .ZN(n3316)
         );
  NAND2_X1 U4385 ( .A1(n3382), .A2(n4432), .ZN(n3967) );
  NAND2_X1 U4386 ( .A1(n3311), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4387 ( .A1(n3341), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4388 ( .A1(n3343), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4389 ( .A1(n3340), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3318)
         );
  NAND2_X1 U4390 ( .A1(n3436), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3325)
         );
  NAND2_X1 U4391 ( .A1(n3430), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3324)
         );
  NAND2_X1 U4392 ( .A1(n3342), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3323) );
  NAND2_X1 U4393 ( .A1(n4111), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U4394 ( .A1(n3339), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3329) );
  NAND2_X1 U4395 ( .A1(n3326), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3328)
         );
  NAND2_X1 U4396 ( .A1(n3431), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3327)
         );
  NAND2_X1 U4397 ( .A1(n3273), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U4398 ( .A1(n3344), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4399 ( .A1(n3349), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4400 ( .A1(n2971), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3331)
         );
  NOR2_X1 U4401 ( .A1(n4400), .A2(n2976), .ZN(n3965) );
  AOI22_X1 U4402 ( .A1(n4111), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4403 ( .A1(n3340), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4404 ( .A1(n3343), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3342), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4405 ( .A1(n3344), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4406 ( .A1(n3349), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4407 ( .A1(n3436), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4408 ( .A1(n3326), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3431), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3351) );
  INV_X1 U4409 ( .A(n3369), .ZN(n4431) );
  INV_X1 U4410 ( .A(n4246), .ZN(n3357) );
  NAND2_X1 U4411 ( .A1(n3358), .A2(n3385), .ZN(n4509) );
  NAND2_X1 U4412 ( .A1(n4199), .A2(n4193), .ZN(n3979) );
  NAND2_X1 U4413 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n4172) );
  NAND2_X1 U4414 ( .A1(n5260), .A2(n4488), .ZN(n4370) );
  OAI22_X1 U4415 ( .A1(n4370), .A2(n5051), .B1(n3963), .B2(n4580), .ZN(n3373)
         );
  NAND2_X1 U4416 ( .A1(n3361), .A2(n3385), .ZN(n3379) );
  NAND2_X1 U4417 ( .A1(n3379), .A2(n4087), .ZN(n3362) );
  NOR2_X2 U4418 ( .A1(n3919), .A2(n4400), .ZN(n3376) );
  NAND2_X1 U4419 ( .A1(n3376), .A2(n3383), .ZN(n4306) );
  NAND2_X1 U4420 ( .A1(n3381), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3372) );
  NAND2_X1 U4421 ( .A1(n3921), .A2(n4244), .ZN(n3368) );
  NAND3_X1 U4422 ( .A1(n4254), .A2(STATE2_REG_0__SCAN_IN), .A3(n4244), .ZN(
        n3367) );
  NAND3_X1 U4423 ( .A1(n3364), .A2(n3358), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3366) );
  OR2_X2 U4424 ( .A1(n3369), .A2(n4249), .ZN(n4240) );
  NAND2_X1 U4425 ( .A1(n4254), .A2(n4244), .ZN(n3374) );
  NAND2_X1 U4426 ( .A1(n3374), .A2(n5434), .ZN(n3375) );
  AOI21_X1 U4427 ( .B1(n3969), .B2(n4561), .A(n3375), .ZN(n3378) );
  NAND2_X1 U4428 ( .A1(n3384), .A2(n2976), .ZN(n3377) );
  OAI21_X1 U4429 ( .B1(n3378), .B2(n3376), .A(n3377), .ZN(n4253) );
  INV_X1 U4430 ( .A(n4253), .ZN(n3394) );
  NAND2_X1 U4431 ( .A1(n3382), .A2(n4087), .ZN(n3388) );
  AND2_X1 U4432 ( .A1(n5260), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6751) );
  AND2_X1 U4433 ( .A1(n4561), .A2(n4400), .ZN(n3387) );
  NOR2_X1 U4434 ( .A1(n3384), .A2(n3383), .ZN(n3386) );
  NAND3_X1 U4435 ( .A1(n3387), .A2(n3386), .A3(n3137), .ZN(n4467) );
  OAI211_X1 U4436 ( .C1(n3391), .C2(n3380), .A(n3390), .B(n3389), .ZN(n3392)
         );
  NAND2_X1 U4437 ( .A1(n3478), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3397) );
  INV_X1 U4438 ( .A(n3963), .ZN(n3513) );
  MUX2_X1 U4439 ( .A(n3514), .B(n3513), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3395) );
  INV_X1 U4440 ( .A(n3489), .ZN(n3457) );
  AOI22_X1 U4441 ( .A1(n4101), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4442 ( .A1(n3437), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4443 ( .A1(n3494), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3431), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4444 ( .A1(n4108), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3399) );
  NAND4_X1 U4445 ( .A1(n3402), .A2(n3401), .A3(n3400), .A4(n3399), .ZN(n3408)
         );
  AOI22_X1 U4446 ( .A1(n3837), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4447 ( .A1(n4109), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4448 ( .A1(n3341), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4449 ( .A1(n3448), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3403) );
  NAND4_X1 U4450 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(n3407)
         );
  AOI21_X2 U4451 ( .B1(n4501), .B2(n4488), .A(n3409), .ZN(n3420) );
  INV_X1 U4452 ( .A(n3420), .ZN(n3419) );
  NAND2_X1 U4453 ( .A1(n3413), .A2(n3412), .ZN(n3414) );
  AND2_X2 U4454 ( .A1(n3485), .A2(n3414), .ZN(n3466) );
  NAND2_X1 U4455 ( .A1(n3415), .A2(n4618), .ZN(n3416) );
  OAI211_X1 U4456 ( .C1(n3946), .C2(n4918), .A(n3489), .B(n3416), .ZN(n3417)
         );
  INV_X1 U4457 ( .A(n3417), .ZN(n3418) );
  NAND2_X1 U4458 ( .A1(n3420), .A2(n3422), .ZN(n3423) );
  NAND2_X1 U4459 ( .A1(n3504), .A2(n3423), .ZN(n4495) );
  INV_X1 U4460 ( .A(n3721), .ZN(n3424) );
  NAND2_X1 U4461 ( .A1(n4849), .A2(n3424), .ZN(n3429) );
  AOI22_X1 U4462 ( .A1(n4150), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n4686), .ZN(n3425) );
  INV_X1 U4463 ( .A(n3425), .ZN(n3427) );
  INV_X1 U4464 ( .A(n3548), .ZN(n3532) );
  INV_X1 U4465 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5194) );
  NOR2_X1 U4466 ( .A1(n3532), .A2(n5194), .ZN(n3426) );
  AOI22_X1 U4467 ( .A1(n3838), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4468 ( .A1(n4101), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4469 ( .A1(n3494), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3431), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4470 ( .A1(n3836), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3432) );
  NAND4_X1 U4471 ( .A1(n3435), .A2(n3434), .A3(n3433), .A4(n3432), .ZN(n3443)
         );
  AOI22_X1 U4472 ( .A1(n3448), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4473 ( .A1(n4109), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4475 ( .A1(n3436), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4476 ( .A1(n3349), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3438) );
  NAND4_X1 U4477 ( .A1(n3441), .A2(n3440), .A3(n3439), .A4(n3438), .ZN(n3442)
         );
  AOI21_X1 U4478 ( .B1(n4561), .B2(n4619), .A(n4488), .ZN(n3455) );
  AOI22_X1 U4479 ( .A1(n3341), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4480 ( .A1(n4109), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4481 ( .A1(n3437), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4482 ( .A1(n3819), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3444) );
  NAND4_X1 U4483 ( .A1(n3447), .A2(n3446), .A3(n3445), .A4(n3444), .ZN(n3454)
         );
  AOI22_X1 U4484 ( .A1(n3837), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4485 ( .A1(n3494), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3431), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4486 ( .A1(n3448), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4487 ( .A1(n4103), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3449) );
  NAND4_X1 U4488 ( .A1(n3452), .A2(n3451), .A3(n3450), .A4(n3449), .ZN(n3453)
         );
  NAND2_X1 U4489 ( .A1(n3398), .A2(n5215), .ZN(n5198) );
  OAI211_X1 U4490 ( .C1(n3946), .C2(n4865), .A(n3455), .B(n5198), .ZN(n3462)
         );
  INV_X1 U4491 ( .A(n4619), .ZN(n3456) );
  XNOR2_X1 U4492 ( .A(n3456), .B(n5215), .ZN(n3458) );
  NAND2_X1 U4493 ( .A1(n3458), .A2(n3457), .ZN(n3461) );
  AND2_X1 U4494 ( .A1(n3462), .A2(n3461), .ZN(n3459) );
  OR2_X1 U4495 ( .A1(n4492), .A2(n3289), .ZN(n3465) );
  AOI22_X1 U4496 ( .A1(n3467), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4686), .ZN(n3469) );
  NAND2_X1 U4497 ( .A1(n3548), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3468) );
  AND2_X1 U4498 ( .A1(n3469), .A2(n3468), .ZN(n3470) );
  NAND2_X1 U4499 ( .A1(n4345), .A2(n4344), .ZN(n4343) );
  NAND2_X1 U4500 ( .A1(n3548), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3477) );
  OAI21_X1 U4501 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3472), .ZN(n6460) );
  NAND2_X1 U4502 ( .A1(n6460), .A2(n3870), .ZN(n3474) );
  NAND2_X1 U4503 ( .A1(n4149), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3473)
         );
  NAND2_X1 U4504 ( .A1(n3474), .A2(n3473), .ZN(n3475) );
  AOI21_X1 U4505 ( .B1(n4150), .B2(EAX_REG_2__SCAN_IN), .A(n3475), .ZN(n3476)
         );
  NAND2_X1 U4506 ( .A1(n3478), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3483) );
  NAND2_X1 U4507 ( .A1(n6554), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U4508 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3479) );
  NAND2_X1 U4509 ( .A1(n3479), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3480) );
  NAND2_X1 U4510 ( .A1(n3481), .A2(n3480), .ZN(n4691) );
  AOI22_X1 U4511 ( .A1(n4691), .A2(n3514), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3513), .ZN(n3482) );
  OAI21_X1 U4512 ( .B1(n3487), .B2(n3486), .A(n4291), .ZN(n4460) );
  AOI22_X1 U4513 ( .A1(n3838), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4514 ( .A1(n4109), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4515 ( .A1(n3437), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4516 ( .A1(n3819), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3490) );
  NAND4_X1 U4517 ( .A1(n3493), .A2(n3492), .A3(n3491), .A4(n3490), .ZN(n3500)
         );
  AOI22_X1 U4518 ( .A1(n3837), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4519 ( .A1(n3494), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3497) );
  AOI22_X1 U4520 ( .A1(n3448), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4521 ( .A1(n4103), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3495) );
  NAND4_X1 U4522 ( .A1(n3498), .A2(n3497), .A3(n3496), .A4(n3495), .ZN(n3499)
         );
  AOI22_X1 U4523 ( .A1(n3954), .A2(n4620), .B1(n3921), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3501) );
  INV_X1 U4524 ( .A(n3503), .ZN(n3505) );
  NAND2_X1 U4525 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  NAND2_X1 U4526 ( .A1(n3535), .A2(n3506), .ZN(n4496) );
  INV_X1 U4527 ( .A(n4149), .ZN(n3642) );
  OAI21_X1 U4528 ( .B1(n4496), .B2(n3721), .A(n3642), .ZN(n4429) );
  NAND2_X1 U4529 ( .A1(n4428), .A2(n4429), .ZN(n3511) );
  INV_X1 U4530 ( .A(n4315), .ZN(n3509) );
  INV_X1 U4531 ( .A(n3507), .ZN(n3508) );
  NAND2_X1 U4532 ( .A1(n3509), .A2(n3508), .ZN(n3510) );
  NAND2_X1 U4533 ( .A1(n3478), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3516) );
  NAND2_X1 U4534 ( .A1(n6627), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4791) );
  NAND2_X1 U4535 ( .A1(n4791), .A2(n6780), .ZN(n3512) );
  AND2_X1 U4536 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4581) );
  NAND2_X1 U4537 ( .A1(n4684), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U4538 ( .A1(n6585), .A2(n3514), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3513), .ZN(n3515) );
  NAND2_X1 U4539 ( .A1(n4446), .A2(n4488), .ZN(n3528) );
  AOI22_X1 U4540 ( .A1(n4109), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4541 ( .A1(n3437), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4542 ( .A1(n3819), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4543 ( .A1(n3494), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3517) );
  NAND4_X1 U4544 ( .A1(n3520), .A2(n3519), .A3(n3518), .A4(n3517), .ZN(n3526)
         );
  AOI22_X1 U4545 ( .A1(n3837), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4546 ( .A1(n4101), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4547 ( .A1(n3448), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4548 ( .A1(n4103), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3521) );
  NAND4_X1 U4549 ( .A1(n3524), .A2(n3523), .A3(n3522), .A4(n3521), .ZN(n3525)
         );
  AOI22_X1 U4550 ( .A1(n3954), .A2(n4649), .B1(n3921), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3527) );
  OAI21_X1 U4551 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3529), .A(n3550), 
        .ZN(n6448) );
  AOI22_X1 U4552 ( .A1(n3870), .A2(n6448), .B1(n4149), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U4553 ( .A1(n4150), .A2(EAX_REG_3__SCAN_IN), .ZN(n3530) );
  OAI211_X1 U4554 ( .C1(n3532), .C2(n4452), .A(n3531), .B(n3530), .ZN(n3533)
         );
  INV_X1 U4555 ( .A(n3533), .ZN(n3534) );
  NAND2_X1 U4556 ( .A1(n4426), .A2(n4516), .ZN(n4576) );
  AOI22_X1 U4557 ( .A1(n3838), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4558 ( .A1(n4109), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4559 ( .A1(n3437), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4560 ( .A1(n3819), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3536) );
  NAND4_X1 U4561 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3545)
         );
  AOI22_X1 U4562 ( .A1(n3837), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4563 ( .A1(n3494), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4564 ( .A1(n3448), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4565 ( .A1(n4103), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3540) );
  NAND4_X1 U4566 ( .A1(n3543), .A2(n3542), .A3(n3541), .A4(n3540), .ZN(n3544)
         );
  NAND2_X1 U4567 ( .A1(n3954), .A2(n5021), .ZN(n3547) );
  NAND2_X1 U4568 ( .A1(n3921), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3546) );
  NAND2_X1 U4569 ( .A1(n3547), .A2(n3546), .ZN(n3556) );
  NAND2_X1 U4570 ( .A1(n3548), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3552) );
  AOI21_X1 U4571 ( .B1(n4657), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3549) );
  AOI21_X1 U4572 ( .B1(n4150), .B2(EAX_REG_4__SCAN_IN), .A(n3549), .ZN(n3551)
         );
  AOI21_X1 U4573 ( .B1(n4657), .B2(n3550), .A(n3571), .ZN(n6312) );
  AOI22_X1 U4574 ( .A1(n3552), .A2(n3551), .B1(n3870), .B2(n6312), .ZN(n3553)
         );
  AOI21_X1 U4575 ( .B1(n4648), .B2(n3424), .A(n3553), .ZN(n4577) );
  INV_X1 U4576 ( .A(n4577), .ZN(n3554) );
  NAND2_X1 U4577 ( .A1(n3555), .A2(n3554), .ZN(n4575) );
  AOI22_X1 U4578 ( .A1(n3836), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4579 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4108), .B1(n4109), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4580 ( .A1(n3437), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4581 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4103), .B1(n4112), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U4582 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3567)
         );
  AOI22_X1 U4583 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n3818), .B1(n3838), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4584 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n3819), .B1(n4101), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4585 ( .A1(n3837), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4586 ( .A1(n3448), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3562) );
  NAND4_X1 U4587 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n3566)
         );
  NAND2_X1 U4588 ( .A1(n3954), .A2(n5032), .ZN(n3569) );
  NAND2_X1 U4589 ( .A1(n3921), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3568) );
  NAND2_X1 U4590 ( .A1(n3569), .A2(n3568), .ZN(n3577) );
  XNOR2_X1 U4591 ( .A(n3578), .B(n3570), .ZN(n5020) );
  NAND2_X1 U4592 ( .A1(n5020), .A2(n3424), .ZN(n3576) );
  OAI21_X1 U4593 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3571), .A(n3591), 
        .ZN(n6440) );
  NAND2_X1 U4594 ( .A1(n6440), .A2(n3870), .ZN(n3573) );
  NAND2_X1 U4595 ( .A1(n4149), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3572)
         );
  NAND2_X1 U4596 ( .A1(n3573), .A2(n3572), .ZN(n3574) );
  AOI21_X1 U4597 ( .B1(n3467), .B2(EAX_REG_5__SCAN_IN), .A(n3574), .ZN(n3575)
         );
  NAND2_X1 U4598 ( .A1(n3576), .A2(n3575), .ZN(n4661) );
  AOI22_X1 U4599 ( .A1(n3838), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4600 ( .A1(n4109), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4601 ( .A1(n3437), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4602 ( .A1(n3819), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3579) );
  NAND4_X1 U4603 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3588)
         );
  AOI22_X1 U4604 ( .A1(n3837), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4605 ( .A1(n3494), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4606 ( .A1(n3448), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4607 ( .A1(n4103), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3583) );
  NAND4_X1 U4608 ( .A1(n3586), .A2(n3585), .A3(n3584), .A4(n3583), .ZN(n3587)
         );
  NAND2_X1 U4609 ( .A1(n3954), .A2(n5203), .ZN(n3590) );
  NAND2_X1 U4610 ( .A1(n3921), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4611 ( .A1(n3596), .A2(n3597), .ZN(n5030) );
  NAND2_X1 U4612 ( .A1(n5030), .A2(n3424), .ZN(n3594) );
  XNOR2_X1 U4613 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3591), .ZN(n5038) );
  AOI22_X1 U4614 ( .A1(n4150), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n4686), .ZN(n3592) );
  MUX2_X1 U4615 ( .A(n5038), .B(n3592), .S(n3976), .Z(n3593) );
  NAND2_X1 U4616 ( .A1(n4661), .A2(n4758), .ZN(n3595) );
  INV_X1 U4617 ( .A(n3596), .ZN(n3599) );
  INV_X1 U4618 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U4619 ( .A1(n3954), .A2(n5215), .ZN(n3600) );
  OAI21_X1 U4620 ( .B1(n3946), .B2(n4933), .A(n3600), .ZN(n3601) );
  NAND2_X1 U4621 ( .A1(n5201), .A2(n3424), .ZN(n3609) );
  AOI22_X1 U4622 ( .A1(n3467), .A2(EAX_REG_7__SCAN_IN), .B1(n4149), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3602) );
  OR2_X1 U4623 ( .A1(n3603), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3604) );
  NAND2_X1 U4624 ( .A1(n3604), .A2(n3620), .ZN(n6433) );
  INV_X1 U4625 ( .A(n6433), .ZN(n3605) );
  NAND2_X1 U4626 ( .A1(n4760), .A2(n4798), .ZN(n4839) );
  NAND2_X1 U4627 ( .A1(n4150), .A2(EAX_REG_8__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4628 ( .A1(n4109), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4629 ( .A1(n4101), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4630 ( .A1(n3836), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4631 ( .A1(n3838), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3610) );
  NAND4_X1 U4632 ( .A1(n3613), .A2(n3612), .A3(n3611), .A4(n3610), .ZN(n3619)
         );
  AOI22_X1 U4633 ( .A1(n3837), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4634 ( .A1(n3436), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4635 ( .A1(n3448), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4636 ( .A1(n4108), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3614) );
  NAND4_X1 U4637 ( .A1(n3617), .A2(n3616), .A3(n3615), .A4(n3614), .ZN(n3618)
         );
  OAI21_X1 U4638 ( .B1(n3619), .B2(n3618), .A(n3424), .ZN(n3623) );
  XNOR2_X1 U4639 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3620), .ZN(n5881) );
  INV_X1 U4640 ( .A(n5881), .ZN(n3621) );
  AOI22_X1 U4641 ( .A1(n4149), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n3870), 
        .B2(n3621), .ZN(n3622) );
  NAND2_X1 U4642 ( .A1(n3627), .A2(n5728), .ZN(n3629) );
  INV_X1 U4643 ( .A(n3657), .ZN(n3628) );
  NAND2_X1 U4644 ( .A1(n3629), .A2(n3628), .ZN(n5869) );
  NAND2_X1 U4645 ( .A1(n5869), .A2(n3870), .ZN(n3645) );
  AOI22_X1 U4646 ( .A1(n3818), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4647 ( .A1(n4108), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4648 ( .A1(n3837), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4649 ( .A1(n3448), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3630) );
  NAND4_X1 U4650 ( .A1(n3633), .A2(n3632), .A3(n3631), .A4(n3630), .ZN(n3639)
         );
  AOI22_X1 U4651 ( .A1(n4109), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4652 ( .A1(n3437), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4653 ( .A1(n3836), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4654 ( .A1(n3341), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3634) );
  NAND4_X1 U4655 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3638)
         );
  OAI21_X1 U4656 ( .B1(n3639), .B2(n3638), .A(n3424), .ZN(n3641) );
  NAND2_X1 U4657 ( .A1(n4150), .A2(EAX_REG_9__SCAN_IN), .ZN(n3640) );
  OAI211_X1 U4658 ( .C1(n3642), .C2(n5728), .A(n3641), .B(n3640), .ZN(n3643)
         );
  INV_X1 U4659 ( .A(n3643), .ZN(n3644) );
  NAND2_X1 U4660 ( .A1(n3467), .A2(EAX_REG_10__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4661 ( .A1(n3838), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4662 ( .A1(n4109), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4663 ( .A1(n3494), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4664 ( .A1(n4103), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3647) );
  NAND4_X1 U4665 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(n3656)
         );
  AOI22_X1 U4666 ( .A1(n3837), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4667 ( .A1(n3437), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4668 ( .A1(n3819), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4669 ( .A1(n3448), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3651) );
  NAND4_X1 U4670 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), .ZN(n3655)
         );
  OAI21_X1 U4671 ( .B1(n3656), .B2(n3655), .A(n3424), .ZN(n3659) );
  XOR2_X1 U4672 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3657), .Z(n6264) );
  INV_X1 U4673 ( .A(n6264), .ZN(n5859) );
  AOI22_X1 U4674 ( .A1(n4149), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n3870), 
        .B2(n5859), .ZN(n3658) );
  AOI22_X1 U4675 ( .A1(n3448), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4676 ( .A1(n3818), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4677 ( .A1(n3494), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4678 ( .A1(n4108), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3661) );
  NAND4_X1 U4679 ( .A1(n3664), .A2(n3663), .A3(n3662), .A4(n3661), .ZN(n3670)
         );
  AOI22_X1 U4680 ( .A1(n4109), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4681 ( .A1(n3437), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4682 ( .A1(n3838), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4683 ( .A1(n3836), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3665) );
  NAND4_X1 U4684 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(n3669)
         );
  NOR2_X1 U4685 ( .A1(n3670), .A2(n3669), .ZN(n3674) );
  NAND2_X1 U4686 ( .A1(n3467), .A2(EAX_REG_11__SCAN_IN), .ZN(n3673) );
  XNOR2_X1 U4687 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3671), .ZN(n6252)
         );
  AOI22_X1 U4688 ( .A1(n3870), .A2(n6252), .B1(n4149), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3672) );
  OAI211_X1 U4689 ( .C1(n3674), .C2(n3721), .A(n3673), .B(n3672), .ZN(n5181)
         );
  XOR2_X1 U4690 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3675), .Z(n6242) );
  NAND2_X1 U4691 ( .A1(n6242), .A2(n3870), .ZN(n3691) );
  INV_X1 U4692 ( .A(EAX_REG_12__SCAN_IN), .ZN(n3677) );
  OAI21_X1 U4693 ( .B1(n6160), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n4686), 
        .ZN(n3676) );
  OAI21_X1 U4694 ( .B1(n3706), .B2(n3677), .A(n3676), .ZN(n3690) );
  AOI22_X1 U4695 ( .A1(n4109), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4696 ( .A1(n3818), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4697 ( .A1(n4110), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4698 ( .A1(n3838), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3678) );
  NAND4_X1 U4699 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3687)
         );
  AOI22_X1 U4700 ( .A1(n3448), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4701 ( .A1(n3836), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4702 ( .A1(n3437), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4703 ( .A1(n4101), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3682) );
  NAND4_X1 U4704 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3686)
         );
  NOR2_X1 U4705 ( .A1(n3687), .A2(n3686), .ZN(n3688) );
  NOR2_X1 U4706 ( .A1(n3721), .A2(n3688), .ZN(n3689) );
  AOI21_X1 U4707 ( .B1(n3691), .B2(n3690), .A(n3689), .ZN(n5516) );
  XNOR2_X1 U4708 ( .A(n3693), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6230)
         );
  INV_X1 U4709 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5551) );
  AOI22_X1 U4710 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n3837), .B1(n3836), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4711 ( .A1(n4109), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4712 ( .A1(n3494), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4713 ( .A1(n4103), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3694) );
  NAND4_X1 U4714 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3703)
         );
  AOI22_X1 U4715 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n4108), .B1(n3838), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4716 ( .A1(n4101), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4717 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n3819), .B1(n4102), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4718 ( .A1(n3448), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3698) );
  NAND4_X1 U4719 ( .A1(n3701), .A2(n3700), .A3(n3699), .A4(n3698), .ZN(n3702)
         );
  OAI21_X1 U4720 ( .B1(n3703), .B2(n3702), .A(n3424), .ZN(n3705) );
  NAND2_X1 U4721 ( .A1(n4149), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3704)
         );
  OAI211_X1 U4722 ( .C1(n3706), .C2(n5551), .A(n3705), .B(n3704), .ZN(n3707)
         );
  AOI21_X1 U4723 ( .B1(n6230), .B2(n3870), .A(n3707), .ZN(n5548) );
  AOI22_X1 U4724 ( .A1(n3448), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4725 ( .A1(n3437), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4726 ( .A1(n3836), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4727 ( .A1(n3818), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3708) );
  NAND4_X1 U4728 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3717)
         );
  AOI22_X1 U4729 ( .A1(n4109), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4730 ( .A1(n3819), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4731 ( .A1(n3494), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4732 ( .A1(n3838), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3712) );
  NAND4_X1 U4733 ( .A1(n3715), .A2(n3714), .A3(n3713), .A4(n3712), .ZN(n3716)
         );
  NOR2_X1 U4734 ( .A1(n3717), .A2(n3716), .ZN(n3722) );
  NAND2_X1 U4735 ( .A1(n3467), .A2(EAX_REG_14__SCAN_IN), .ZN(n3720) );
  XNOR2_X1 U4736 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3718), .ZN(n6221)
         );
  AOI22_X1 U4737 ( .A1(n3870), .A2(n6221), .B1(n4149), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3719) );
  OAI211_X1 U4738 ( .C1(n3722), .C2(n3721), .A(n3720), .B(n3719), .ZN(n5512)
         );
  INV_X1 U4739 ( .A(n5510), .ZN(n3739) );
  NAND2_X1 U4740 ( .A1(n3467), .A2(EAX_REG_15__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4741 ( .A1(n3818), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4742 ( .A1(n4101), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4743 ( .A1(n3836), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4744 ( .A1(n3838), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3723) );
  NAND4_X1 U4745 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3732)
         );
  AOI22_X1 U4746 ( .A1(n3448), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4747 ( .A1(n3436), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4748 ( .A1(n3494), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4749 ( .A1(n4109), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3727) );
  NAND4_X1 U4750 ( .A1(n3730), .A2(n3729), .A3(n3728), .A4(n3727), .ZN(n3731)
         );
  OAI21_X1 U4751 ( .B1(n3732), .B2(n3731), .A(n3424), .ZN(n3736) );
  INV_X1 U4752 ( .A(n3733), .ZN(n3734) );
  XNOR2_X1 U4753 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3734), .ZN(n6211)
         );
  AOI22_X1 U4754 ( .A1(n3870), .A2(n6211), .B1(n4149), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3735) );
  NAND2_X1 U4755 ( .A1(n3739), .A2(n3738), .ZN(n5499) );
  INV_X1 U4756 ( .A(n3768), .ZN(n3742) );
  OR2_X1 U4757 ( .A1(n3740), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3741)
         );
  NAND2_X1 U4758 ( .A1(n3742), .A2(n3741), .ZN(n6193) );
  AOI22_X1 U4759 ( .A1(n3437), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4760 ( .A1(n3836), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4761 ( .A1(n3838), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4762 ( .A1(n3448), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3743) );
  NAND4_X1 U4763 ( .A1(n3746), .A2(n3745), .A3(n3744), .A4(n3743), .ZN(n3752)
         );
  AOI22_X1 U4764 ( .A1(n4101), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4765 ( .A1(n3819), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4766 ( .A1(n3837), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4767 ( .A1(n4109), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3747) );
  NAND4_X1 U4768 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n3751)
         );
  NOR2_X1 U4769 ( .A1(n3752), .A2(n3751), .ZN(n3754) );
  AOI22_X1 U4770 ( .A1(n3467), .A2(EAX_REG_16__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n4149), .ZN(n3753) );
  OAI21_X1 U4771 ( .B1(n4124), .B2(n3754), .A(n3753), .ZN(n3755) );
  AOI21_X1 U4772 ( .B1(n6193), .B2(n3870), .A(n3755), .ZN(n5498) );
  AOI22_X1 U4773 ( .A1(n3837), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4774 ( .A1(n3818), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4775 ( .A1(n3436), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4776 ( .A1(n3448), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3756) );
  NAND4_X1 U4777 ( .A1(n3759), .A2(n3758), .A3(n3757), .A4(n3756), .ZN(n3765)
         );
  AOI22_X1 U4778 ( .A1(n4109), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4779 ( .A1(n4101), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4780 ( .A1(n3494), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4781 ( .A1(n4103), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U4782 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3764)
         );
  NOR2_X1 U4783 ( .A1(n3765), .A2(n3764), .ZN(n3767) );
  AOI22_X1 U4784 ( .A1(n3467), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4686), .ZN(n3766) );
  OAI21_X1 U4785 ( .B1(n4124), .B2(n3767), .A(n3766), .ZN(n3769) );
  XNOR2_X1 U4786 ( .A(n3768), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5675)
         );
  MUX2_X1 U4787 ( .A(n3769), .B(n5675), .S(n3870), .Z(n5390) );
  OAI21_X1 U4788 ( .B1(n3770), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n3785), 
        .ZN(n6186) );
  AOI22_X1 U4789 ( .A1(n3448), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4790 ( .A1(n4109), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4791 ( .A1(n3437), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4792 ( .A1(n3836), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3771) );
  NAND4_X1 U4793 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3780)
         );
  AOI22_X1 U4794 ( .A1(n3818), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4795 ( .A1(n3837), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4796 ( .A1(n3838), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4797 ( .A1(n4112), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4798 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3779)
         );
  NOR2_X1 U4799 ( .A1(n3780), .A2(n3779), .ZN(n3782) );
  AOI22_X1 U4800 ( .A1(n4150), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4686), .ZN(n3781) );
  OAI21_X1 U4801 ( .B1(n4124), .B2(n3782), .A(n3781), .ZN(n3783) );
  MUX2_X1 U4802 ( .A(n6186), .B(n3783), .S(n3976), .Z(n3784) );
  XNOR2_X1 U4803 ( .A(n3785), .B(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6142)
         );
  NAND2_X1 U4804 ( .A1(n6142), .A2(n3870), .ZN(n3800) );
  AOI22_X1 U4805 ( .A1(n3838), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4806 ( .A1(n4109), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4807 ( .A1(n3437), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4101), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4808 ( .A1(n3819), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4809 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3795)
         );
  AOI22_X1 U4810 ( .A1(n3837), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4811 ( .A1(n3494), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4812 ( .A1(n3448), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4813 ( .A1(n4103), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3790) );
  NAND4_X1 U4814 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3794)
         );
  NOR2_X1 U4815 ( .A1(n3795), .A2(n3794), .ZN(n3798) );
  INV_X1 U4816 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5659) );
  AOI21_X1 U4817 ( .B1(n5659), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3796) );
  AOI21_X1 U4818 ( .B1(n3467), .B2(EAX_REG_19__SCAN_IN), .A(n3796), .ZN(n3797)
         );
  OAI21_X1 U4819 ( .B1(n4124), .B2(n3798), .A(n3797), .ZN(n3799) );
  NAND2_X1 U4820 ( .A1(n3800), .A2(n3799), .ZN(n5484) );
  NAND2_X1 U4821 ( .A1(n3801), .A2(n5650), .ZN(n3802) );
  AND2_X1 U4822 ( .A1(n3817), .A2(n3802), .ZN(n5648) );
  AOI22_X1 U4823 ( .A1(n3448), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4824 ( .A1(n3818), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4825 ( .A1(n3436), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4826 ( .A1(n3836), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4827 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3812)
         );
  AOI22_X1 U4828 ( .A1(n4109), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4829 ( .A1(n4101), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4830 ( .A1(n4112), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4831 ( .A1(n4103), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4832 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3811)
         );
  OR2_X1 U4833 ( .A1(n3812), .A2(n3811), .ZN(n3815) );
  INV_X1 U4834 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3813) );
  OAI22_X1 U4835 ( .A1(n3706), .A2(n3813), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5650), .ZN(n3814) );
  AOI21_X1 U4836 ( .B1(n3893), .B2(n3815), .A(n3814), .ZN(n3816) );
  MUX2_X1 U4837 ( .A(n5648), .B(n3816), .S(n3976), .Z(n5374) );
  XNOR2_X1 U4838 ( .A(n3817), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5640)
         );
  AOI22_X1 U4839 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n4108), .B1(n3838), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4840 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n3818), .B1(n4109), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4841 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n3437), .B1(n4101), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4842 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n3819), .B1(n4102), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4843 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3830)
         );
  AOI22_X1 U4844 ( .A1(n3837), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4845 ( .A1(n3494), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4846 ( .A1(n3448), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4847 ( .A1(n4103), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3825) );
  NAND4_X1 U4848 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3829)
         );
  OR2_X1 U4849 ( .A1(n3830), .A2(n3829), .ZN(n3834) );
  INV_X1 U4850 ( .A(EAX_REG_21__SCAN_IN), .ZN(n3832) );
  OAI21_X1 U4851 ( .B1(n6160), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4686), 
        .ZN(n3831) );
  OAI21_X1 U4852 ( .B1(n3706), .B2(n3832), .A(n3831), .ZN(n3833) );
  AOI21_X1 U4853 ( .B1(n3893), .B2(n3834), .A(n3833), .ZN(n3835) );
  AOI21_X1 U4854 ( .B1(n5640), .B2(n3870), .A(n3835), .ZN(n5362) );
  AOI22_X1 U4855 ( .A1(n3837), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4856 ( .A1(n3448), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4857 ( .A1(n4101), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4858 ( .A1(n3436), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4859 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3848)
         );
  AOI22_X1 U4860 ( .A1(n3818), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4861 ( .A1(n3494), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4862 ( .A1(n4109), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4863 ( .A1(n4112), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4864 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3847)
         );
  NOR2_X1 U4865 ( .A1(n3848), .A2(n3847), .ZN(n3850) );
  AOI22_X1 U4866 ( .A1(n3467), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n4686), .ZN(n3849) );
  OAI21_X1 U4867 ( .B1(n4124), .B2(n3850), .A(n3849), .ZN(n3854) );
  INV_X1 U4868 ( .A(n3851), .ZN(n3852) );
  INV_X1 U4869 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U4870 ( .A1(n3852), .A2(n5351), .ZN(n3853) );
  NAND2_X1 U4871 ( .A1(n3856), .A2(n3853), .ZN(n5634) );
  MUX2_X1 U4872 ( .A(n3854), .B(n5634), .S(n3870), .Z(n3855) );
  XNOR2_X1 U4873 ( .A(n3856), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5624)
         );
  NAND2_X1 U4874 ( .A1(n5624), .A2(n3870), .ZN(n3864) );
  XOR2_X1 U4875 ( .A(n3858), .B(n3857), .Z(n3859) );
  NAND2_X1 U4876 ( .A1(n3859), .A2(n3893), .ZN(n3862) );
  AOI21_X1 U4877 ( .B1(n5626), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3860) );
  AOI21_X1 U4878 ( .B1(n3467), .B2(EAX_REG_23__SCAN_IN), .A(n3860), .ZN(n3861)
         );
  NAND2_X1 U4879 ( .A1(n3862), .A2(n3861), .ZN(n3863) );
  NAND2_X1 U4880 ( .A1(n3864), .A2(n3863), .ZN(n5333) );
  XNOR2_X1 U4881 ( .A(n3867), .B(n3866), .ZN(n3873) );
  NAND2_X1 U4882 ( .A1(n3868), .A2(n5615), .ZN(n3869) );
  NAND2_X1 U4883 ( .A1(n3879), .A2(n3869), .ZN(n5614) );
  NAND2_X1 U4884 ( .A1(n5614), .A2(n3870), .ZN(n3872) );
  AOI22_X1 U4885 ( .A1(n4150), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4149), .ZN(n3871) );
  OAI211_X1 U4886 ( .C1(n4124), .C2(n3873), .A(n3872), .B(n3871), .ZN(n5321)
         );
  XOR2_X1 U4887 ( .A(n3875), .B(n3874), .Z(n3878) );
  INV_X1 U4888 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3876) );
  INV_X1 U4889 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5597) );
  OAI22_X1 U4890 ( .A1(n3706), .A2(n3876), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5597), .ZN(n3877) );
  AOI21_X1 U4891 ( .B1(n3878), .B2(n3893), .A(n3877), .ZN(n3880) );
  XNOR2_X1 U4892 ( .A(n3879), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5599)
         );
  MUX2_X1 U4893 ( .A(n3880), .B(n5599), .S(n3870), .Z(n5309) );
  NAND2_X1 U4894 ( .A1(n3882), .A2(n3881), .ZN(n3883) );
  NAND2_X1 U4895 ( .A1(n2987), .A2(n3883), .ZN(n5587) );
  XNOR2_X1 U4896 ( .A(n3885), .B(n3884), .ZN(n3887) );
  AOI22_X1 U4897 ( .A1(n3467), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n4686), .ZN(n3886) );
  OAI21_X1 U4898 ( .B1(n3887), .B2(n4124), .A(n3886), .ZN(n3888) );
  MUX2_X1 U4899 ( .A(n5587), .B(n3888), .S(n3976), .Z(n5295) );
  XOR2_X1 U4900 ( .A(n3890), .B(n3889), .Z(n3894) );
  INV_X1 U4901 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3891) );
  OAI22_X1 U4902 ( .A1(n3706), .A2(n3891), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5583), .ZN(n3892) );
  AOI21_X1 U4903 ( .B1(n3894), .B2(n3893), .A(n3892), .ZN(n3895) );
  XNOR2_X1 U4904 ( .A(n2987), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5581)
         );
  MUX2_X1 U4905 ( .A(n3895), .B(n5581), .S(n3870), .Z(n5282) );
  XNOR2_X1 U4906 ( .A(n3897), .B(n3896), .ZN(n3899) );
  AOI22_X1 U4907 ( .A1(n4150), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n4686), .ZN(n3898) );
  OAI21_X1 U4908 ( .B1(n3899), .B2(n4124), .A(n3898), .ZN(n3902) );
  NAND2_X1 U4909 ( .A1(n3900), .A2(n5573), .ZN(n3901) );
  NAND2_X1 U4910 ( .A1(n3904), .A2(n3901), .ZN(n5572) );
  MUX2_X1 U4911 ( .A(n3902), .B(n5572), .S(n3870), .Z(n5271) );
  AOI21_X1 U4912 ( .B1(n3903), .B2(n5270), .A(n4128), .ZN(n5563) );
  INV_X1 U4913 ( .A(n5563), .ZN(n4100) );
  NAND2_X1 U4914 ( .A1(n3905), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3907)
         );
  INV_X1 U4915 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3906) );
  INV_X1 U4916 ( .A(n3925), .ZN(n3908) );
  XNOR2_X1 U4917 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3926) );
  XNOR2_X1 U4918 ( .A(n3908), .B(n3926), .ZN(n3970) );
  AND2_X1 U4919 ( .A1(n3970), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3915) );
  NAND2_X1 U4920 ( .A1(n3398), .A2(n4432), .ZN(n4243) );
  AND2_X1 U4921 ( .A1(n3018), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3909)
         );
  NOR2_X1 U4922 ( .A1(n3925), .A2(n3909), .ZN(n3913) );
  NAND2_X1 U4923 ( .A1(n3380), .A2(n4432), .ZN(n3911) );
  NAND2_X1 U4924 ( .A1(n3910), .A2(n3911), .ZN(n3929) );
  OAI22_X1 U4925 ( .A1(n3914), .A2(n3915), .B1(n3912), .B2(n3929), .ZN(n3922)
         );
  NAND2_X1 U4926 ( .A1(n3954), .A2(n3913), .ZN(n3918) );
  INV_X1 U4927 ( .A(n3914), .ZN(n3917) );
  INV_X1 U4928 ( .A(n3915), .ZN(n3916) );
  OAI22_X1 U4929 ( .A1(n3922), .A2(n3918), .B1(n3917), .B2(n3916), .ZN(n3924)
         );
  INV_X1 U4930 ( .A(n3919), .ZN(n3920) );
  AOI21_X1 U4931 ( .B1(n3922), .B2(n3970), .A(n3959), .ZN(n3923) );
  NAND2_X1 U4932 ( .A1(n3926), .A2(n3925), .ZN(n3928) );
  NAND2_X1 U4933 ( .A1(n4580), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3927) );
  NAND2_X1 U4934 ( .A1(n3928), .A2(n3927), .ZN(n3936) );
  XNOR2_X1 U4935 ( .A(n5264), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3934)
         );
  XNOR2_X1 U4936 ( .A(n3936), .B(n3934), .ZN(n3971) );
  NAND2_X1 U4937 ( .A1(n3954), .A2(n3971), .ZN(n3932) );
  INV_X1 U4938 ( .A(n3929), .ZN(n3933) );
  OAI211_X1 U4939 ( .C1(n3971), .C2(n3946), .A(n3932), .B(n3933), .ZN(n3930)
         );
  NAND2_X1 U4940 ( .A1(n3931), .A2(n3930), .ZN(n3949) );
  INV_X1 U4941 ( .A(n3934), .ZN(n3935) );
  NAND2_X1 U4942 ( .A1(n3936), .A2(n3935), .ZN(n3938) );
  NAND2_X1 U4943 ( .A1(n4852), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3937) );
  NAND2_X1 U4944 ( .A1(n3938), .A2(n3937), .ZN(n3943) );
  NAND2_X1 U4945 ( .A1(n4452), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3939) );
  NAND2_X1 U4946 ( .A1(n3943), .A2(n3941), .ZN(n3940) );
  NAND2_X1 U4947 ( .A1(n3940), .A2(n5706), .ZN(n3951) );
  INV_X1 U4948 ( .A(n3941), .ZN(n3942) );
  XNOR2_X1 U4949 ( .A(n3943), .B(n3942), .ZN(n3944) );
  INV_X1 U4950 ( .A(n3974), .ZN(n3956) );
  NAND2_X1 U4951 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4295), .ZN(n3952) );
  AOI22_X1 U4952 ( .A1(n3954), .A2(n3960), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4488), .ZN(n3955) );
  OAI21_X1 U4953 ( .B1(n3956), .B2(n3959), .A(n3955), .ZN(n3957) );
  INV_X1 U4954 ( .A(n3965), .ZN(n3966) );
  NAND2_X1 U4955 ( .A1(n3971), .A2(n3970), .ZN(n3973) );
  OAI21_X1 U4956 ( .B1(n3974), .B2(n3973), .A(n3972), .ZN(n4276) );
  INV_X1 U4957 ( .A(n4276), .ZN(n3975) );
  NAND2_X1 U4958 ( .A1(n4261), .A2(n6750), .ZN(n4238) );
  NAND2_X1 U4959 ( .A1(n4488), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4180) );
  NOR2_X1 U4960 ( .A1(n3976), .A2(n4180), .ZN(n6756) );
  INV_X1 U4961 ( .A(n6756), .ZN(n3977) );
  NAND2_X1 U4962 ( .A1(n6797), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6158) );
  NAND3_X1 U4963 ( .A1(n3977), .A2(n6120), .A3(n4979), .ZN(n3978) );
  NAND2_X1 U4964 ( .A1(n6233), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3996) );
  INV_X1 U4965 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6206) );
  INV_X1 U4966 ( .A(REIP_REG_9__SCAN_IN), .ZN(n4213) );
  INV_X1 U4967 ( .A(REIP_REG_7__SCAN_IN), .ZN(n4209) );
  INV_X1 U4968 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6287) );
  NAND4_X1 U4969 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .A4(REIP_REG_3__SCAN_IN), .ZN(n6288) );
  NOR2_X1 U4970 ( .A1(n6287), .A2(n6288), .ZN(n5419) );
  NAND2_X1 U4971 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5419), .ZN(n6275) );
  NOR2_X1 U4972 ( .A1(n4209), .A2(n6275), .ZN(n5414) );
  NAND2_X1 U4973 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5414), .ZN(n5404) );
  NOR2_X1 U4974 ( .A1(n4213), .A2(n5404), .ZN(n6269) );
  NAND2_X1 U4975 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6269), .ZN(n6248) );
  NOR2_X1 U4976 ( .A1(n6247), .A2(n6248), .ZN(n6241) );
  NAND2_X1 U4977 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6241), .ZN(n6227) );
  NOR2_X1 U4978 ( .A1(n5787), .A2(n6227), .ZN(n3990) );
  NAND3_X1 U4979 ( .A1(REIP_REG_14__SCAN_IN), .A2(n3990), .A3(n6233), .ZN(
        n6190) );
  NAND2_X1 U4980 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n3991) );
  NOR3_X1 U4981 ( .A1(n6206), .A2(n6190), .A3(n3991), .ZN(n3981) );
  NAND3_X1 U4982 ( .A1(n3979), .A2(n4171), .A3(n4172), .ZN(n4380) );
  NAND2_X1 U4983 ( .A1(n3380), .A2(n4380), .ZN(n4388) );
  NOR2_X1 U4984 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n4088) );
  NAND3_X1 U4985 ( .A1(n4388), .A2(n4088), .A3(n2976), .ZN(n3980) );
  NAND2_X1 U4986 ( .A1(n6289), .A2(n6233), .ZN(n6191) );
  INV_X1 U4987 ( .A(n6191), .ZN(n6232) );
  OR2_X1 U4988 ( .A1(n3981), .A2(n6232), .ZN(n5391) );
  AND3_X1 U4989 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_20__SCAN_IN), .ZN(n3992) );
  INV_X1 U4990 ( .A(n3992), .ZN(n3982) );
  NAND2_X1 U4991 ( .A1(n6191), .A2(n3982), .ZN(n3983) );
  NAND2_X1 U4992 ( .A1(REIP_REG_21__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .ZN(
        n5341) );
  INV_X1 U4993 ( .A(REIP_REG_23__SCAN_IN), .ZN(n3984) );
  NOR2_X1 U4994 ( .A1(n5341), .A2(n3984), .ZN(n3993) );
  INV_X1 U4995 ( .A(n3993), .ZN(n3985) );
  NAND2_X1 U4996 ( .A1(n6319), .A2(n3985), .ZN(n3986) );
  NAND2_X1 U4997 ( .A1(n5383), .A2(n3986), .ZN(n5342) );
  AND3_X1 U4998 ( .A1(REIP_REG_25__SCAN_IN), .A2(REIP_REG_24__SCAN_IN), .A3(
        REIP_REG_26__SCAN_IN), .ZN(n3994) );
  INV_X1 U4999 ( .A(n3994), .ZN(n3987) );
  AND2_X1 U5000 ( .A1(n6191), .A2(n3987), .ZN(n3988) );
  NOR2_X1 U5001 ( .A1(n5342), .A2(n3988), .ZN(n5300) );
  NAND2_X1 U5002 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4141) );
  NAND2_X1 U5003 ( .A1(n6319), .A2(n4141), .ZN(n3989) );
  INV_X1 U5004 ( .A(REIP_REG_29__SCAN_IN), .ZN(n4198) );
  INV_X1 U5005 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U5006 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6192), .ZN(n6199) );
  NOR2_X1 U5007 ( .A1(REIP_REG_29__SCAN_IN), .A2(n4141), .ZN(n3995) );
  NAND2_X1 U5008 ( .A1(n5278), .A2(n3995), .ZN(n4144) );
  INV_X1 U5009 ( .A(n3996), .ZN(n3997) );
  INV_X1 U5010 ( .A(EBX_REG_1__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U5011 ( .A1(n2984), .A2(n5456), .ZN(n3999) );
  OAI211_X1 U5012 ( .C1(n4016), .C2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n3999), 
        .B(n5377), .ZN(n4000) );
  INV_X1 U5013 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5465) );
  XNOR2_X1 U5014 ( .A(n4001), .B(n4340), .ZN(n4321) );
  NOR2_X1 U5015 ( .A1(n4321), .A2(n4395), .ZN(n4003) );
  INV_X1 U5016 ( .A(n4001), .ZN(n4002) );
  NOR2_X2 U5017 ( .A1(n4003), .A2(n4002), .ZN(n4423) );
  MUX2_X1 U5018 ( .A(n4081), .B(n4077), .S(EBX_REG_2__SCAN_IN), .Z(n4006) );
  NAND2_X1 U5019 ( .A1(n4395), .A2(n4016), .ZN(n4047) );
  NAND2_X1 U5020 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n4395), .ZN(n4004)
         );
  AND2_X1 U5021 ( .A1(n4047), .A2(n4004), .ZN(n4005) );
  NAND2_X1 U5022 ( .A1(n4006), .A2(n4005), .ZN(n4422) );
  INV_X1 U5023 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6527) );
  INV_X1 U5024 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U5025 ( .A1(n2984), .A2(n6334), .ZN(n4008) );
  OAI211_X1 U5026 ( .C1(n6802), .C2(n6527), .A(n4008), .B(n4077), .ZN(n4009)
         );
  OAI21_X1 U5027 ( .B1(n4083), .B2(EBX_REG_3__SCAN_IN), .A(n4009), .ZN(n5433)
         );
  MUX2_X1 U5028 ( .A(n4081), .B(n4077), .S(EBX_REG_4__SCAN_IN), .Z(n4012) );
  NAND2_X1 U5029 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n4395), .ZN(n4010)
         );
  AND2_X1 U5030 ( .A1(n4047), .A2(n4010), .ZN(n4011) );
  NAND2_X1 U5031 ( .A1(n4012), .A2(n4011), .ZN(n4616) );
  MUX2_X1 U5032 ( .A(n4083), .B(n5377), .S(EBX_REG_5__SCAN_IN), .Z(n4013) );
  OAI21_X1 U5033 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4342), .A(n4013), 
        .ZN(n4664) );
  INV_X1 U5034 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4014) );
  NAND2_X1 U5035 ( .A1(n2984), .A2(n4014), .ZN(n4015) );
  OAI211_X1 U5036 ( .C1(n4016), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4015), 
        .B(n5377), .ZN(n4017) );
  OAI21_X1 U5037 ( .B1(n4081), .B2(EBX_REG_6__SCAN_IN), .A(n4017), .ZN(n4762)
         );
  NAND2_X1 U5038 ( .A1(n4662), .A2(n4762), .ZN(n4799) );
  INV_X1 U5039 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6493) );
  INV_X1 U5040 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U5041 ( .A1(n2984), .A2(n5796), .ZN(n4018) );
  OAI211_X1 U5042 ( .C1(n6802), .C2(n6493), .A(n4018), .B(n4077), .ZN(n4019)
         );
  OAI21_X1 U5043 ( .B1(n4083), .B2(EBX_REG_7__SCAN_IN), .A(n4019), .ZN(n4801)
         );
  NOR2_X2 U5044 ( .A1(n4799), .A2(n4801), .ZN(n4843) );
  INV_X1 U5045 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4020) );
  NAND2_X1 U5046 ( .A1(n4026), .A2(n4020), .ZN(n4024) );
  INV_X1 U5047 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U5048 ( .A1(n4077), .A2(n6487), .ZN(n4022) );
  NAND2_X1 U5049 ( .A1(n2984), .A2(n4020), .ZN(n4021) );
  NAND3_X1 U5050 ( .A1(n4022), .A2(n5377), .A3(n4021), .ZN(n4023) );
  NAND2_X1 U5051 ( .A1(n4024), .A2(n4023), .ZN(n4844) );
  NAND2_X1 U5052 ( .A1(n4843), .A2(n4844), .ZN(n4845) );
  MUX2_X1 U5053 ( .A(n4083), .B(n5377), .S(EBX_REG_9__SCAN_IN), .Z(n4025) );
  OAI21_X1 U5054 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n4342), .A(n4025), 
        .ZN(n5045) );
  INV_X1 U5055 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U5056 ( .A1(n4026), .A2(n6258), .ZN(n4030) );
  INV_X1 U5057 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U5058 ( .A1(n4077), .A2(n5837), .ZN(n4028) );
  NAND2_X1 U5059 ( .A1(n2984), .A2(n6258), .ZN(n4027) );
  NAND3_X1 U5060 ( .A1(n4028), .A2(n5377), .A3(n4027), .ZN(n4029) );
  NAND2_X1 U5061 ( .A1(n4030), .A2(n4029), .ZN(n5175) );
  INV_X1 U5062 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6468) );
  INV_X1 U5063 ( .A(EBX_REG_11__SCAN_IN), .ZN(n4031) );
  NAND2_X1 U5064 ( .A1(n2984), .A2(n4031), .ZN(n4032) );
  OAI211_X1 U5065 ( .C1(n6802), .C2(n6468), .A(n4032), .B(n4077), .ZN(n4033)
         );
  OAI21_X1 U5066 ( .B1(n4083), .B2(EBX_REG_11__SCAN_IN), .A(n4033), .ZN(n5186)
         );
  MUX2_X1 U5067 ( .A(n4081), .B(n4077), .S(EBX_REG_12__SCAN_IN), .Z(n4036) );
  NAND2_X1 U5068 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4395), .ZN(n4034) );
  AND2_X1 U5069 ( .A1(n4047), .A2(n4034), .ZN(n4035) );
  AND2_X1 U5070 ( .A1(n4036), .A2(n4035), .ZN(n5517) );
  INV_X1 U5071 ( .A(n4083), .ZN(n4073) );
  INV_X1 U5072 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U5073 ( .A1(n4073), .A2(n6329), .ZN(n4040) );
  NAND2_X1 U5074 ( .A1(n2984), .A2(n6329), .ZN(n4038) );
  NAND2_X1 U5075 ( .A1(n5377), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4037) );
  NAND3_X1 U5076 ( .A1(n4038), .A2(n4077), .A3(n4037), .ZN(n4039) );
  MUX2_X1 U5077 ( .A(n4081), .B(n4077), .S(EBX_REG_14__SCAN_IN), .Z(n4043) );
  NAND2_X1 U5078 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4395), .ZN(n4041) );
  AND2_X1 U5079 ( .A1(n4047), .A2(n4041), .ZN(n4042) );
  NAND2_X1 U5080 ( .A1(n4043), .A2(n4042), .ZN(n5508) );
  NAND2_X1 U5081 ( .A1(n5507), .A2(n5508), .ZN(n5506) );
  INV_X1 U5082 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6068) );
  INV_X1 U5083 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U5084 ( .A1(n2984), .A2(n6325), .ZN(n4044) );
  OAI211_X1 U5085 ( .C1(n6802), .C2(n6068), .A(n4044), .B(n4077), .ZN(n4045)
         );
  OAI21_X1 U5086 ( .B1(n4083), .B2(EBX_REG_15__SCAN_IN), .A(n4045), .ZN(n6064)
         );
  MUX2_X1 U5087 ( .A(n4081), .B(n4077), .S(EBX_REG_16__SCAN_IN), .Z(n4049) );
  NAND2_X1 U5088 ( .A1(n4395), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4046) );
  AND2_X1 U5089 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  NAND2_X1 U5090 ( .A1(n4049), .A2(n4048), .ZN(n5502) );
  NAND2_X1 U5091 ( .A1(n5501), .A2(n5502), .ZN(n5393) );
  INV_X1 U5092 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6049) );
  INV_X1 U5093 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U5094 ( .A1(n2984), .A2(n5398), .ZN(n4050) );
  OAI211_X1 U5095 ( .C1(n6802), .C2(n6049), .A(n4050), .B(n4077), .ZN(n4051)
         );
  OAI21_X1 U5096 ( .B1(n4083), .B2(EBX_REG_17__SCAN_IN), .A(n4051), .ZN(n5394)
         );
  MUX2_X1 U5097 ( .A(n4081), .B(n4077), .S(EBX_REG_19__SCAN_IN), .Z(n4053) );
  NAND2_X1 U5098 ( .A1(n4395), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4052) );
  NAND2_X1 U5099 ( .A1(n4053), .A2(n4052), .ZN(n5487) );
  OR2_X1 U5100 ( .A1(n4342), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4055)
         );
  INV_X1 U5101 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U5102 ( .A1(n2984), .A2(n5482), .ZN(n4054) );
  AND2_X1 U5103 ( .A1(n4055), .A2(n4054), .ZN(n5379) );
  OR2_X1 U5104 ( .A1(n4342), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4056)
         );
  INV_X1 U5105 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U5106 ( .A1(n2984), .A2(n5494), .ZN(n5485) );
  NAND2_X1 U5107 ( .A1(n4056), .A2(n5485), .ZN(n5486) );
  NAND2_X1 U5108 ( .A1(n6802), .A2(EBX_REG_20__SCAN_IN), .ZN(n4058) );
  NAND2_X1 U5109 ( .A1(n5486), .A2(n5377), .ZN(n4057) );
  OAI211_X1 U5110 ( .C1(n5379), .C2(n5486), .A(n4058), .B(n4057), .ZN(n4059)
         );
  MUX2_X1 U5111 ( .A(n4083), .B(n5377), .S(EBX_REG_21__SCAN_IN), .Z(n4060) );
  OAI21_X1 U5112 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4342), .A(n4060), 
        .ZN(n4061) );
  INV_X1 U5113 ( .A(n4061), .ZN(n5365) );
  MUX2_X1 U5114 ( .A(n4081), .B(n4077), .S(EBX_REG_22__SCAN_IN), .Z(n4063) );
  NAND2_X1 U5115 ( .A1(n4395), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U5116 ( .A1(n4063), .A2(n4062), .ZN(n5350) );
  INV_X1 U5117 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U5118 ( .A1(n2984), .A2(n5479), .ZN(n4065) );
  NAND2_X1 U5119 ( .A1(n5377), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4064) );
  NAND3_X1 U5120 ( .A1(n4065), .A2(n4077), .A3(n4064), .ZN(n4066) );
  OAI21_X1 U5121 ( .B1(n4083), .B2(EBX_REG_23__SCAN_IN), .A(n4066), .ZN(n5335)
         );
  MUX2_X1 U5122 ( .A(n4081), .B(n4077), .S(EBX_REG_24__SCAN_IN), .Z(n4068) );
  NAND2_X1 U5123 ( .A1(n4395), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4067) );
  NAND2_X1 U5124 ( .A1(n4068), .A2(n4067), .ZN(n5324) );
  MUX2_X1 U5125 ( .A(n4083), .B(n5377), .S(EBX_REG_25__SCAN_IN), .Z(n4069) );
  OAI21_X1 U5126 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4342), .A(n4069), 
        .ZN(n5311) );
  INV_X1 U5127 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U5128 ( .A1(n4077), .A2(n5962), .ZN(n4071) );
  INV_X1 U5129 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U5130 ( .A1(n2984), .A2(n5476), .ZN(n4070) );
  NAND3_X1 U5131 ( .A1(n4071), .A2(n5377), .A3(n4070), .ZN(n4072) );
  OAI21_X1 U5132 ( .B1(n4081), .B2(EBX_REG_26__SCAN_IN), .A(n4072), .ZN(n5297)
         );
  INV_X1 U5133 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U5134 ( .A1(n4073), .A2(n5475), .ZN(n4076) );
  INV_X1 U5135 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U5136 ( .A1(n2984), .A2(n5475), .ZN(n4074) );
  OAI211_X1 U5137 ( .C1(n6802), .C2(n5952), .A(n4074), .B(n4077), .ZN(n4075)
         );
  NAND2_X1 U5138 ( .A1(n4077), .A2(n5939), .ZN(n4079) );
  INV_X1 U5139 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U5140 ( .A1(n2984), .A2(n5474), .ZN(n4078) );
  NAND3_X1 U5141 ( .A1(n4079), .A2(n5377), .A3(n4078), .ZN(n4080) );
  OAI21_X1 U5142 ( .B1(n4081), .B2(EBX_REG_28__SCAN_IN), .A(n4080), .ZN(n5273)
         );
  OR2_X1 U5143 ( .A1(n4342), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4130)
         );
  INV_X1 U5144 ( .A(n4130), .ZN(n4082) );
  MUX2_X1 U5145 ( .A(EBX_REG_29__SCAN_IN), .B(n4082), .S(n5377), .Z(n4085) );
  NOR2_X1 U5146 ( .A1(n4083), .A2(EBX_REG_29__SCAN_IN), .ZN(n4084) );
  NOR2_X1 U5147 ( .A1(n4085), .A2(n4084), .ZN(n4153) );
  XNOR2_X1 U5148 ( .A(n2983), .B(n4153), .ZN(n5472) );
  NAND2_X1 U5149 ( .A1(n2984), .A2(EBX_REG_31__SCAN_IN), .ZN(n4086) );
  NAND2_X1 U5150 ( .A1(n5472), .A2(n6305), .ZN(n4095) );
  INV_X1 U5151 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U5152 ( .A1(n2976), .A2(n5766), .ZN(n4092) );
  INV_X1 U5153 ( .A(n4088), .ZN(n4089) );
  OR2_X1 U5154 ( .A1(n4380), .A2(n4089), .ZN(n4974) );
  NAND2_X1 U5155 ( .A1(n5216), .A2(n4974), .ZN(n4090) );
  OR2_X1 U5156 ( .A1(n5435), .A2(n4090), .ZN(n4091) );
  OAI21_X1 U5157 ( .B1(n4093), .B2(n4092), .A(n4091), .ZN(n6229) );
  AOI22_X1 U5158 ( .A1(n6303), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6306), .ZN(n4094) );
  NAND2_X1 U5159 ( .A1(n4095), .A2(n4094), .ZN(n4096) );
  OAI211_X1 U5160 ( .C1(n5272), .C2(n4198), .A(n4144), .B(n4097), .ZN(n4098)
         );
  INV_X1 U5161 ( .A(n4098), .ZN(n4099) );
  AOI22_X1 U5162 ( .A1(n3836), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3494), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5163 ( .A1(n4101), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5164 ( .A1(n3819), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4102), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5165 ( .A1(n4103), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4104) );
  NAND4_X1 U5166 ( .A1(n4107), .A2(n4106), .A3(n4105), .A4(n4104), .ZN(n4118)
         );
  AOI22_X1 U5167 ( .A1(n3838), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5168 ( .A1(n4109), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5169 ( .A1(n4111), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4110), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5170 ( .A1(n3448), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4112), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4113) );
  NAND4_X1 U5171 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(n4117)
         );
  NOR2_X1 U5172 ( .A1(n4118), .A2(n4117), .ZN(n4122) );
  NOR2_X1 U5173 ( .A1(n4120), .A2(n4119), .ZN(n4121) );
  XOR2_X1 U5174 ( .A(n4122), .B(n4121), .Z(n4125) );
  AOI22_X1 U5175 ( .A1(n3467), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n4686), .ZN(n4123) );
  OAI21_X1 U5176 ( .B1(n4125), .B2(n4124), .A(n4123), .ZN(n4127) );
  XOR2_X1 U5177 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .B(n4126), .Z(n5196) );
  MUX2_X1 U5178 ( .A(n4127), .B(n5196), .S(n3870), .Z(n4129) );
  NAND2_X1 U5179 ( .A1(n4128), .A2(n4129), .ZN(n4152) );
  OAI21_X1 U5180 ( .B1(EBX_REG_29__SCAN_IN), .B2(n4395), .A(n4130), .ZN(n4131)
         );
  INV_X1 U5181 ( .A(n2983), .ZN(n4155) );
  NAND2_X1 U5182 ( .A1(n4137), .A2(n4155), .ZN(n4135) );
  NAND2_X1 U5183 ( .A1(n4342), .A2(EBX_REG_30__SCAN_IN), .ZN(n4133) );
  NAND2_X1 U5184 ( .A1(n4395), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4132) );
  AND2_X1 U5185 ( .A1(n4133), .A2(n4132), .ZN(n4154) );
  INV_X1 U5186 ( .A(n4154), .ZN(n4134) );
  NAND3_X1 U5187 ( .A1(n4157), .A2(n4135), .A3(n4134), .ZN(n4139) );
  NAND2_X1 U5188 ( .A1(n2983), .A2(n6802), .ZN(n4136) );
  NAND3_X1 U5189 ( .A1(n4137), .A2(n4154), .A3(n4136), .ZN(n4138) );
  NAND2_X1 U5190 ( .A1(n4139), .A2(n4138), .ZN(n5922) );
  AOI22_X1 U5191 ( .A1(n6303), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6306), .ZN(n4140) );
  OAI21_X1 U5192 ( .B1(n5922), .B2(n6260), .A(n4140), .ZN(n4147) );
  INV_X1 U5193 ( .A(n4141), .ZN(n4142) );
  NAND2_X1 U5194 ( .A1(REIP_REG_29__SCAN_IN), .A2(n4142), .ZN(n4143) );
  NOR2_X1 U5195 ( .A1(n5293), .A2(n4143), .ZN(n4164) );
  INV_X1 U5196 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4222) );
  NAND2_X1 U5197 ( .A1(n4144), .A2(n5272), .ZN(n4166) );
  NAND3_X1 U5198 ( .A1(n4155), .A2(n4154), .A3(n4153), .ZN(n4156) );
  NAND2_X1 U5199 ( .A1(n4157), .A2(n4156), .ZN(n4160) );
  INV_X1 U5200 ( .A(n4342), .ZN(n4158) );
  INV_X1 U5201 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5916) );
  AOI22_X1 U5202 ( .A1(n4158), .A2(n5916), .B1(n2984), .B2(n5766), .ZN(n4159)
         );
  NAND3_X1 U5203 ( .A1(n5216), .A2(EBX_REG_31__SCAN_IN), .A3(n4974), .ZN(n4162) );
  NAND2_X1 U5204 ( .A1(n6306), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4161)
         );
  OAI21_X1 U5205 ( .B1(n5435), .B2(n4162), .A(n4161), .ZN(n4163) );
  INV_X1 U5206 ( .A(REIP_REG_31__SCAN_IN), .ZN(n4237) );
  NOR2_X1 U5207 ( .A1(n6289), .A2(REIP_REG_30__SCAN_IN), .ZN(n4165) );
  OAI21_X1 U5208 ( .B1(n4166), .B2(n4165), .A(REIP_REG_31__SCAN_IN), .ZN(n4167) );
  INV_X1 U5209 ( .A(READY_N), .ZN(n4179) );
  AOI221_X1 U5210 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4179), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4168) );
  AOI221_X1 U5211 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n4168), .C2(HOLD), .A(n4171), .ZN(n4175) );
  AND2_X1 U5212 ( .A1(n4172), .A2(n4171), .ZN(n4170) );
  INV_X1 U5213 ( .A(NA_N), .ZN(n4173) );
  NAND2_X1 U5214 ( .A1(n4173), .A2(STATE_REG_2__SCAN_IN), .ZN(n4169) );
  AND2_X1 U5215 ( .A1(n4170), .A2(n4169), .ZN(n4186) );
  AOI22_X1 U5216 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n4190) );
  INV_X1 U5217 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4184) );
  NOR2_X1 U5218 ( .A1(n4171), .A2(n4184), .ZN(n4177) );
  INV_X1 U5219 ( .A(n4172), .ZN(n4189) );
  AOI21_X1 U5220 ( .B1(n4173), .B2(n4177), .A(n4189), .ZN(n4174) );
  OAI22_X1 U5221 ( .A1(n4175), .A2(n4186), .B1(n4190), .B2(n4174), .ZN(U3183)
         );
  AND2_X1 U5222 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n4185) );
  NAND2_X1 U5223 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4176) );
  OAI21_X1 U5224 ( .B1(n4177), .B2(n4185), .A(n4176), .ZN(n4178) );
  OAI211_X1 U5225 ( .C1(n4179), .C2(n4199), .A(n4178), .B(n4380), .ZN(U3182)
         );
  AOI211_X1 U5226 ( .C1(n4686), .C2(READY_N), .A(n6748), .B(n6797), .ZN(n4181)
         );
  NAND2_X1 U5227 ( .A1(n4490), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6767) );
  NOR2_X1 U5228 ( .A1(n4180), .A2(n6160), .ZN(n4369) );
  AOI21_X1 U5229 ( .B1(n4181), .B2(n6767), .A(n4369), .ZN(n4182) );
  INV_X1 U5230 ( .A(n4182), .ZN(U3150) );
  INV_X2 U5231 ( .A(n4202), .ZN(n6137) );
  NAND2_X1 U5232 ( .A1(n6137), .A2(W_R_N_REG_SCAN_IN), .ZN(n4183) );
  OAI21_X1 U5233 ( .B1(n6137), .B2(READREQUEST_REG_SCAN_IN), .A(n4183), .ZN(
        U3470) );
  OAI21_X1 U5234 ( .B1(n4185), .B2(n4184), .A(n6137), .ZN(n4188) );
  INV_X1 U5235 ( .A(n4186), .ZN(n4187) );
  OAI211_X1 U5236 ( .C1(n4190), .C2(n4189), .A(n4188), .B(n4187), .ZN(U3181)
         );
  NOR2_X1 U5237 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6159) );
  OAI21_X1 U5238 ( .B1(n6159), .B2(D_C_N_REG_SCAN_IN), .A(n6137), .ZN(n4191)
         );
  OAI21_X1 U5239 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6137), .A(n4191), .ZN(
        U2791) );
  INV_X1 U5240 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6790) );
  NAND2_X1 U5241 ( .A1(BE_N_REG_0__SCAN_IN), .A2(n6137), .ZN(n4192) );
  OAI21_X1 U5242 ( .B1(n6790), .B2(n6137), .A(n4192), .ZN(U3448) );
  INV_X1 U5243 ( .A(REIP_REG_24__SCAN_IN), .ZN(n5329) );
  INV_X1 U5244 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n4194) );
  OAI222_X1 U5245 ( .A1(n4215), .A2(n5329), .B1(n4194), .B2(n4202), .C1(n4203), 
        .C2(n3984), .ZN(U3206) );
  INV_X1 U5246 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n5737) );
  OAI222_X1 U5247 ( .A1(n4215), .A2(n6217), .B1(n4203), .B2(n5787), .C1(n5737), 
        .C2(n4202), .ZN(U3196) );
  INV_X1 U5248 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6138) );
  INV_X1 U5249 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n4195) );
  OAI222_X1 U5250 ( .A1(n4215), .A2(n6138), .B1(n4195), .B2(n4202), .C1(n4203), 
        .C2(n4230), .ZN(U3200) );
  INV_X1 U5251 ( .A(REIP_REG_20__SCAN_IN), .ZN(n4197) );
  INV_X1 U5252 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n4196) );
  INV_X1 U5253 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6139) );
  OAI222_X1 U5254 ( .A1(n4215), .A2(n4197), .B1(n4196), .B2(n4202), .C1(n4203), 
        .C2(n6139), .ZN(U3202) );
  INV_X1 U5255 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5352) );
  INV_X1 U5256 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n5798) );
  OAI222_X1 U5257 ( .A1(n4203), .A2(n5352), .B1(n4202), .B2(n5798), .C1(n4215), 
        .C2(n3984), .ZN(U3205) );
  INV_X1 U5258 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5793) );
  INV_X1 U5259 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n5782) );
  OAI222_X1 U5260 ( .A1(n4203), .A2(n5793), .B1(n4202), .B2(n5782), .C1(n4198), 
        .C2(n4215), .ZN(U3211) );
  INV_X1 U5261 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4201) );
  OAI21_X1 U5262 ( .B1(n4199), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n4200) );
  OAI21_X1 U5263 ( .B1(n4202), .B2(n4201), .A(n6761), .ZN(U2789) );
  INV_X1 U5264 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6270) );
  AOI22_X1 U5265 ( .A1(n4235), .A2(REIP_REG_9__SCAN_IN), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6137), .ZN(n4204) );
  OAI21_X1 U5266 ( .B1(n6270), .B2(n4215), .A(n4204), .ZN(U3192) );
  AOI22_X1 U5267 ( .A1(n4235), .A2(REIP_REG_4__SCAN_IN), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6137), .ZN(n4205) );
  OAI21_X1 U5268 ( .B1(n6287), .B2(n4215), .A(n4205), .ZN(U3187) );
  INV_X1 U5269 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U5270 ( .A1(n4235), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6137), .ZN(n4206) );
  OAI21_X1 U5271 ( .B1(n4207), .B2(n4215), .A(n4206), .ZN(U3185) );
  AOI22_X1 U5272 ( .A1(n4235), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6137), .ZN(n4208) );
  OAI21_X1 U5273 ( .B1(n4209), .B2(n4215), .A(n4208), .ZN(U3189) );
  INV_X1 U5274 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5877) );
  AOI22_X1 U5275 ( .A1(n4235), .A2(REIP_REG_7__SCAN_IN), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6137), .ZN(n4210) );
  OAI21_X1 U5276 ( .B1(n5877), .B2(n4215), .A(n4210), .ZN(U3190) );
  INV_X1 U5277 ( .A(REIP_REG_6__SCAN_IN), .ZN(n5422) );
  AOI22_X1 U5278 ( .A1(n4235), .A2(REIP_REG_5__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6137), .ZN(n4211) );
  OAI21_X1 U5279 ( .B1(n5422), .B2(n4215), .A(n4211), .ZN(U3188) );
  AOI22_X1 U5280 ( .A1(n4235), .A2(REIP_REG_8__SCAN_IN), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6137), .ZN(n4212) );
  OAI21_X1 U5281 ( .B1(n4213), .B2(n4215), .A(n4212), .ZN(U3191) );
  AOI22_X1 U5282 ( .A1(n4235), .A2(REIP_REG_10__SCAN_IN), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6137), .ZN(n4214) );
  OAI21_X1 U5283 ( .B1(n6247), .B2(n4215), .A(n4214), .ZN(U3193) );
  INV_X1 U5284 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6318) );
  AOI22_X1 U5285 ( .A1(n4235), .A2(REIP_REG_3__SCAN_IN), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6137), .ZN(n4216) );
  OAI21_X1 U5286 ( .B1(n6318), .B2(n4215), .A(n4216), .ZN(U3186) );
  AOI22_X1 U5287 ( .A1(n4235), .A2(REIP_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6137), .ZN(n4217) );
  OAI21_X1 U5288 ( .B1(n5787), .B2(n4215), .A(n4217), .ZN(U3195) );
  INV_X1 U5289 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6316) );
  AOI22_X1 U5290 ( .A1(n4235), .A2(REIP_REG_1__SCAN_IN), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6137), .ZN(n4218) );
  OAI21_X1 U5291 ( .B1(n6316), .B2(n4215), .A(n4218), .ZN(U3184) );
  INV_X1 U5292 ( .A(REIP_REG_25__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5293 ( .A1(n4235), .A2(REIP_REG_24__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6137), .ZN(n4219) );
  OAI21_X1 U5294 ( .B1(n4220), .B2(n4215), .A(n4219), .ZN(U3207) );
  AOI22_X1 U5295 ( .A1(n4235), .A2(REIP_REG_29__SCAN_IN), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6137), .ZN(n4221) );
  OAI21_X1 U5296 ( .B1(n4222), .B2(n4215), .A(n4221), .ZN(U3212) );
  INV_X1 U5297 ( .A(REIP_REG_12__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U5298 ( .A1(n4235), .A2(REIP_REG_11__SCAN_IN), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6137), .ZN(n4223) );
  OAI21_X1 U5299 ( .B1(n4224), .B2(n4215), .A(n4223), .ZN(U3194) );
  AOI22_X1 U5300 ( .A1(n4235), .A2(REIP_REG_18__SCAN_IN), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6137), .ZN(n4225) );
  OAI21_X1 U5301 ( .B1(n6139), .B2(n4215), .A(n4225), .ZN(U3201) );
  AOI22_X1 U5302 ( .A1(n4235), .A2(REIP_REG_14__SCAN_IN), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6137), .ZN(n4226) );
  OAI21_X1 U5303 ( .B1(n6206), .B2(n4215), .A(n4226), .ZN(U3197) );
  INV_X1 U5304 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6205) );
  AOI22_X1 U5305 ( .A1(n4235), .A2(REIP_REG_15__SCAN_IN), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6137), .ZN(n4227) );
  OAI21_X1 U5306 ( .B1(n6205), .B2(n4215), .A(n4227), .ZN(U3198) );
  AOI22_X1 U5307 ( .A1(n4235), .A2(REIP_REG_21__SCAN_IN), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6137), .ZN(n4228) );
  OAI21_X1 U5308 ( .B1(n5352), .B2(n4215), .A(n4228), .ZN(U3204) );
  INV_X1 U5309 ( .A(REIP_REG_17__SCAN_IN), .ZN(n4230) );
  AOI22_X1 U5310 ( .A1(n4235), .A2(REIP_REG_16__SCAN_IN), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6137), .ZN(n4229) );
  OAI21_X1 U5311 ( .B1(n4230), .B2(n4215), .A(n4229), .ZN(U3199) );
  INV_X1 U5312 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5301) );
  AOI22_X1 U5313 ( .A1(n4235), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6137), .ZN(n4231) );
  OAI21_X1 U5314 ( .B1(n5301), .B2(n4215), .A(n4231), .ZN(U3208) );
  INV_X1 U5315 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5288) );
  AOI22_X1 U5316 ( .A1(n4235), .A2(REIP_REG_26__SCAN_IN), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6137), .ZN(n4232) );
  OAI21_X1 U5317 ( .B1(n5288), .B2(n4215), .A(n4232), .ZN(U3209) );
  AOI22_X1 U5318 ( .A1(n4235), .A2(REIP_REG_27__SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6137), .ZN(n4233) );
  OAI21_X1 U5319 ( .B1(n5793), .B2(n4215), .A(n4233), .ZN(U3210) );
  INV_X1 U5320 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5369) );
  AOI22_X1 U5321 ( .A1(n4235), .A2(REIP_REG_20__SCAN_IN), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6137), .ZN(n4234) );
  OAI21_X1 U5322 ( .B1(n5369), .B2(n4215), .A(n4234), .ZN(U3203) );
  AOI22_X1 U5323 ( .A1(n4235), .A2(REIP_REG_30__SCAN_IN), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6137), .ZN(n4236) );
  OAI21_X1 U5324 ( .B1(n4237), .B2(n4215), .A(n4236), .ZN(U3213) );
  NOR2_X1 U5325 ( .A1(n6678), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5392) );
  INV_X1 U5326 ( .A(n4298), .ZN(n4296) );
  AOI211_X1 U5327 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4238), .A(n5392), .B(
        n4296), .ZN(n4239) );
  INV_X1 U5328 ( .A(n4239), .ZN(U2788) );
  INV_X1 U5329 ( .A(n4240), .ZN(n4242) );
  NAND2_X1 U5330 ( .A1(n4257), .A2(n4561), .ZN(n4241) );
  NAND2_X1 U5331 ( .A1(n4242), .A2(n4241), .ZN(n4282) );
  NOR2_X1 U5332 ( .A1(n4282), .A2(n3910), .ZN(n4275) );
  INV_X1 U5333 ( .A(n4275), .ZN(n4447) );
  NAND3_X1 U5334 ( .A1(n4447), .A2(n3964), .A3(n4964), .ZN(n4258) );
  NOR2_X1 U5335 ( .A1(n5434), .A2(n3384), .ZN(n4285) );
  OAI21_X1 U5336 ( .B1(n4285), .B2(n4342), .A(n3369), .ZN(n4251) );
  NAND2_X1 U5337 ( .A1(n4244), .A2(n2976), .ZN(n4245) );
  NAND2_X1 U5338 ( .A1(n6796), .A2(n4245), .ZN(n4248) );
  NAND2_X1 U5339 ( .A1(n4248), .A2(n4247), .ZN(n4280) );
  INV_X1 U5340 ( .A(n4249), .ZN(n4250) );
  NAND3_X1 U5341 ( .A1(n4251), .A2(n4280), .A3(n4250), .ZN(n4252) );
  OR2_X1 U5342 ( .A1(n4253), .A2(n4252), .ZN(n4305) );
  NAND2_X1 U5343 ( .A1(n3376), .A2(n4254), .ZN(n4255) );
  NAND2_X1 U5344 ( .A1(n4255), .A2(n4467), .ZN(n4256) );
  NOR2_X1 U5345 ( .A1(n4257), .A2(n3380), .ZN(n4379) );
  NAND2_X1 U5346 ( .A1(n4407), .A2(n4379), .ZN(n4448) );
  INV_X1 U5347 ( .A(n4448), .ZN(n4409) );
  MUX2_X1 U5348 ( .A(n4258), .B(n4409), .S(n4386), .Z(n4259) );
  AOI21_X1 U5349 ( .B1(n4276), .B2(n4279), .A(n4259), .ZN(n4965) );
  OR2_X1 U5350 ( .A1(n4386), .A2(n4260), .ZN(n4264) );
  INV_X1 U5351 ( .A(n4261), .ZN(n4262) );
  NAND2_X1 U5352 ( .A1(n4262), .A2(n3964), .ZN(n4263) );
  NAND2_X1 U5353 ( .A1(n4264), .A2(n4263), .ZN(n6156) );
  INV_X1 U5354 ( .A(n5434), .ZN(n4265) );
  OR2_X1 U5355 ( .A1(n5216), .A2(n4265), .ZN(n5266) );
  AOI21_X1 U5356 ( .B1(n5266), .B2(n4380), .A(READY_N), .ZN(n6795) );
  NOR2_X1 U5357 ( .A1(n6156), .A2(n6795), .ZN(n4962) );
  INV_X1 U5358 ( .A(n6750), .ZN(n6155) );
  OR2_X1 U5359 ( .A1(n4962), .A2(n6155), .ZN(n4268) );
  INV_X1 U5360 ( .A(n4268), .ZN(n6163) );
  INV_X1 U5361 ( .A(MORE_REG_SCAN_IN), .ZN(n4266) );
  OR2_X1 U5362 ( .A1(n6163), .A2(n4266), .ZN(n4267) );
  OAI21_X1 U5363 ( .B1(n4965), .B2(n4268), .A(n4267), .ZN(U3471) );
  INV_X1 U5364 ( .A(n4380), .ZN(n4270) );
  NOR2_X1 U5365 ( .A1(n2984), .A2(n4270), .ZN(n4272) );
  NAND2_X1 U5366 ( .A1(n4950), .A2(n4270), .ZN(n4271) );
  OAI21_X1 U5367 ( .B1(n4272), .B2(n4269), .A(n4271), .ZN(n4273) );
  NAND2_X1 U5368 ( .A1(n4273), .A2(n4179), .ZN(n4274) );
  MUX2_X1 U5369 ( .A(n4448), .B(n4274), .S(n4386), .Z(n4289) );
  NAND2_X1 U5370 ( .A1(n4386), .A2(n4275), .ZN(n4278) );
  NOR2_X1 U5371 ( .A1(READY_N), .A2(n4276), .ZN(n4381) );
  NAND2_X1 U5372 ( .A1(n4482), .A2(n4381), .ZN(n4277) );
  INV_X1 U5373 ( .A(n4279), .ZN(n4284) );
  INV_X1 U5374 ( .A(n4280), .ZN(n4281) );
  OR2_X1 U5375 ( .A1(n4282), .A2(n4281), .ZN(n4283) );
  NAND2_X1 U5376 ( .A1(n4284), .A2(n4283), .ZN(n4384) );
  INV_X1 U5377 ( .A(n4285), .ZN(n4286) );
  NAND2_X1 U5378 ( .A1(n4384), .A2(n4286), .ZN(n4287) );
  NOR2_X1 U5379 ( .A1(n4507), .A2(n4287), .ZN(n4288) );
  OAI22_X1 U5380 ( .A1(n4954), .A2(n6155), .B1(n6162), .B2(n6767), .ZN(n4293)
         );
  NOR2_X1 U5381 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6769), .ZN(n6766) );
  INV_X1 U5382 ( .A(n4290), .ZN(n5087) );
  OR2_X1 U5383 ( .A1(n4291), .A2(n5087), .ZN(n4292) );
  XNOR2_X1 U5384 ( .A(n4292), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6301)
         );
  NAND4_X1 U5385 ( .A1(n4293), .A2(n4482), .A3(n5260), .A4(n6301), .ZN(n4294)
         );
  OAI21_X1 U5386 ( .B1(n6135), .B2(n4295), .A(n4294), .ZN(U3455) );
  OAI21_X2 U5387 ( .B1(n5216), .B2(n4179), .A(n4296), .ZN(n6420) );
  INV_X1 U5388 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U5389 ( .A1(n6419), .A2(EAX_REG_29__SCAN_IN), .ZN(n4299) );
  NAND2_X1 U5390 ( .A1(n6409), .A2(DATAI_13_), .ZN(n4300) );
  OAI211_X1 U5391 ( .C1(n4350), .C2(n5801), .A(n4299), .B(n4300), .ZN(U2937)
         );
  INV_X1 U5392 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U5393 ( .A1(n6419), .A2(EAX_REG_13__SCAN_IN), .ZN(n4301) );
  OAI211_X1 U5394 ( .C1(n4350), .C2(n5769), .A(n4301), .B(n4300), .ZN(U2952)
         );
  INV_X1 U5395 ( .A(n4973), .ZN(n4302) );
  INV_X1 U5396 ( .A(n6392), .ZN(n6367) );
  INV_X2 U5397 ( .A(n6791), .ZN(n6390) );
  AOI222_X1 U5398 ( .A1(n6385), .A2(DATAO_REG_0__SCAN_IN), .B1(n6367), .B2(
        EAX_REG_0__SCAN_IN), .C1(n6390), .C2(LWORD_REG_0__SCAN_IN), .ZN(n4304)
         );
  INV_X1 U5399 ( .A(n4304), .ZN(U2923) );
  OAI21_X1 U5400 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6132), .A(n6135), 
        .ZN(n5188) );
  INV_X1 U5401 ( .A(n4305), .ZN(n4310) );
  INV_X1 U5402 ( .A(n4319), .ZN(n4307) );
  NAND3_X1 U5403 ( .A1(n4269), .A2(n4306), .A3(n4307), .ZN(n4308) );
  NOR2_X1 U5404 ( .A1(n4482), .A2(n4308), .ZN(n4309) );
  AND2_X1 U5405 ( .A1(n4310), .A2(n4309), .ZN(n4462) );
  INV_X1 U5406 ( .A(n4462), .ZN(n4946) );
  AOI22_X1 U5407 ( .A1(n4946), .A2(n3466), .B1(n4948), .B2(n3018), .ZN(n4944)
         );
  INV_X1 U5408 ( .A(n5260), .ZN(n6133) );
  OAI22_X1 U5409 ( .A1(n4944), .A2(n6133), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6747), .ZN(n4311) );
  OAI22_X1 U5410 ( .A1(n5188), .A2(n4311), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6135), .ZN(n4313) );
  NAND3_X1 U5411 ( .A1(n4950), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n5260), .ZN(n4312) );
  NAND2_X1 U5412 ( .A1(n4313), .A2(n4312), .ZN(U3461) );
  INV_X1 U5413 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4314) );
  OAI222_X1 U5414 ( .A1(n4314), .A2(n6369), .B1(n6791), .B2(n5769), .C1(n5551), 
        .C2(n6392), .ZN(U2910) );
  OAI21_X1 U5415 ( .B1(n4317), .B2(n4316), .A(n4315), .ZN(n5463) );
  AND3_X1 U5416 ( .A1(n5251), .A2(n3398), .A3(n3289), .ZN(n4318) );
  NAND2_X1 U5417 ( .A1(n4319), .A2(n4318), .ZN(n4505) );
  OAI22_X1 U5418 ( .A1(n4448), .A2(n4386), .B1(n4395), .B2(n4505), .ZN(n4320)
         );
  AND2_X1 U5419 ( .A1(n6335), .A2(n3385), .ZN(n6332) );
  NAND2_X1 U5420 ( .A1(n6335), .A2(n5251), .ZN(n5519) );
  XNOR2_X1 U5421 ( .A(n4321), .B(n4395), .ZN(n5459) );
  AOI22_X1 U5422 ( .A1(n6331), .A2(n5459), .B1(n5504), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4322) );
  OAI21_X1 U5423 ( .B1(n5463), .B2(n5521), .A(n4322), .ZN(U2858) );
  AOI22_X1 U5424 ( .A1(n6420), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6419), .ZN(n4323) );
  NAND2_X1 U5425 ( .A1(n6409), .A2(DATAI_6_), .ZN(n4324) );
  NAND2_X1 U5426 ( .A1(n4323), .A2(n4324), .ZN(U2945) );
  AOI22_X1 U5427 ( .A1(n6420), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6419), .ZN(n4325) );
  NAND2_X1 U5428 ( .A1(n4325), .A2(n4324), .ZN(U2930) );
  AOI22_X1 U5429 ( .A1(n6420), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6419), .ZN(n4326) );
  NAND2_X1 U5430 ( .A1(n6409), .A2(DATAI_7_), .ZN(n4352) );
  NAND2_X1 U5431 ( .A1(n4326), .A2(n4352), .ZN(U2946) );
  AOI22_X1 U5432 ( .A1(n6420), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6419), .ZN(n4327) );
  NAND2_X1 U5433 ( .A1(n6409), .A2(DATAI_4_), .ZN(n4360) );
  NAND2_X1 U5434 ( .A1(n4327), .A2(n4360), .ZN(U2943) );
  AOI22_X1 U5435 ( .A1(n6420), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6419), .ZN(n4328) );
  NAND2_X1 U5436 ( .A1(n6409), .A2(DATAI_5_), .ZN(n4356) );
  NAND2_X1 U5437 ( .A1(n4328), .A2(n4356), .ZN(U2944) );
  AOI22_X1 U5438 ( .A1(n6420), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n6419), .ZN(n4329) );
  INV_X1 U5439 ( .A(DATAI_9_), .ZN(n5124) );
  OR2_X1 U5440 ( .A1(n6406), .A2(n5124), .ZN(n4331) );
  NAND2_X1 U5441 ( .A1(n4329), .A2(n4331), .ZN(U2933) );
  AOI22_X1 U5442 ( .A1(n6420), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6419), .ZN(n4330) );
  NAND2_X1 U5443 ( .A1(n6409), .A2(DATAI_3_), .ZN(n4354) );
  NAND2_X1 U5444 ( .A1(n4330), .A2(n4354), .ZN(U2942) );
  AOI22_X1 U5445 ( .A1(n6420), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6419), .ZN(n4332) );
  NAND2_X1 U5446 ( .A1(n4332), .A2(n4331), .ZN(U2948) );
  INV_X1 U5447 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4334) );
  INV_X1 U5448 ( .A(n6359), .ZN(n4362) );
  INV_X1 U5449 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n4333) );
  OAI222_X1 U5450 ( .A1(n4334), .A2(n6369), .B1(n4362), .B2(n3876), .C1(n6791), 
        .C2(n4333), .ZN(U2898) );
  INV_X1 U5451 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4337) );
  INV_X1 U5452 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4336) );
  INV_X1 U5453 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4335) );
  OAI222_X1 U5454 ( .A1(n4337), .A2(n6369), .B1(n4362), .B2(n4336), .C1(n6791), 
        .C2(n4335), .ZN(U2900) );
  INV_X1 U5455 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4339) );
  INV_X1 U5456 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n4338) );
  OAI222_X1 U5457 ( .A1(n4339), .A2(n6369), .B1(n4362), .B2(n3832), .C1(n6791), 
        .C2(n4338), .ZN(U2902) );
  INV_X1 U5458 ( .A(n4340), .ZN(n4341) );
  OAI21_X1 U5459 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n4342), .A(n4341), 
        .ZN(n5464) );
  OAI21_X1 U5460 ( .B1(n4345), .B2(n4344), .A(n4343), .ZN(n5470) );
  OAI222_X1 U5461 ( .A1(n5464), .A2(n5519), .B1(n6335), .B2(n5465), .C1(n5470), 
        .C2(n5521), .ZN(U2859) );
  INV_X1 U5462 ( .A(DATAI_0_), .ZN(n4519) );
  AOI22_X1 U5463 ( .A1(n6420), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6419), .ZN(n4346) );
  OAI21_X1 U5464 ( .B1(n4519), .B2(n6406), .A(n4346), .ZN(U2939) );
  INV_X1 U5465 ( .A(DATAI_15_), .ZN(n6348) );
  AOI22_X1 U5466 ( .A1(n6420), .A2(LWORD_REG_15__SCAN_IN), .B1(
        EAX_REG_15__SCAN_IN), .B2(n6419), .ZN(n4347) );
  OAI21_X1 U5467 ( .B1(n6348), .B2(n6406), .A(n4347), .ZN(U2954) );
  INV_X1 U5468 ( .A(DATAI_2_), .ZN(n4514) );
  AOI22_X1 U5469 ( .A1(n6420), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6419), .ZN(n4348) );
  OAI21_X1 U5470 ( .B1(n4514), .B2(n6406), .A(n4348), .ZN(U2941) );
  INV_X1 U5471 ( .A(DATAI_1_), .ZN(n4515) );
  AOI22_X1 U5472 ( .A1(n6420), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6419), .ZN(n4349) );
  OAI21_X1 U5473 ( .B1(n4515), .B2(n6406), .A(n4349), .ZN(U2940) );
  AOI22_X1 U5474 ( .A1(n6416), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6419), .ZN(n4351) );
  INV_X1 U5475 ( .A(DATAI_10_), .ZN(n5178) );
  OR2_X1 U5476 ( .A1(n6406), .A2(n5178), .ZN(n4358) );
  NAND2_X1 U5477 ( .A1(n4351), .A2(n4358), .ZN(U2949) );
  AOI22_X1 U5478 ( .A1(n6416), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6419), .ZN(n4353) );
  NAND2_X1 U5479 ( .A1(n4353), .A2(n4352), .ZN(U2931) );
  AOI22_X1 U5480 ( .A1(n6416), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6419), .ZN(n4355) );
  NAND2_X1 U5481 ( .A1(n4355), .A2(n4354), .ZN(U2927) );
  AOI22_X1 U5482 ( .A1(n6416), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6419), .ZN(n4357) );
  NAND2_X1 U5483 ( .A1(n4357), .A2(n4356), .ZN(U2929) );
  AOI22_X1 U5484 ( .A1(n6416), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n6419), .ZN(n4359) );
  NAND2_X1 U5485 ( .A1(n4359), .A2(n4358), .ZN(U2934) );
  AOI22_X1 U5486 ( .A1(n6416), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6419), .ZN(n4361) );
  NAND2_X1 U5487 ( .A1(n4361), .A2(n4360), .ZN(U2928) );
  INV_X1 U5488 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4364) );
  OAI222_X1 U5489 ( .A1(n4364), .A2(n6369), .B1(n6791), .B2(n5801), .C1(n4363), 
        .C2(n4362), .ZN(U2894) );
  NAND2_X1 U5490 ( .A1(n4492), .A2(n3920), .ZN(n4368) );
  INV_X1 U5491 ( .A(n4254), .ZN(n4365) );
  OAI21_X1 U5492 ( .B1(n6796), .B2(n4619), .A(n4365), .ZN(n4366) );
  INV_X1 U5493 ( .A(n4366), .ZN(n4367) );
  NAND2_X1 U5494 ( .A1(n4368), .A2(n4367), .ZN(n4437) );
  XNOR2_X1 U5495 ( .A(n4437), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4413)
         );
  INV_X1 U5496 ( .A(n5470), .ZN(n4377) );
  INV_X1 U5497 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6788) );
  NOR2_X1 U5498 ( .A1(n6120), .A2(n6788), .ZN(n4405) );
  NAND2_X1 U5499 ( .A1(n4370), .A2(n6678), .ZN(n6792) );
  NAND2_X1 U5500 ( .A1(n6792), .A2(n4488), .ZN(n4371) );
  NAND2_X1 U5501 ( .A1(n4488), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U5502 ( .A1(n6160), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4372) );
  NAND2_X1 U5503 ( .A1(n4373), .A2(n4372), .ZN(n4656) );
  INV_X1 U5504 ( .A(n4656), .ZN(n4375) );
  INV_X1 U5505 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4374) );
  AOI21_X1 U5506 ( .B1(n5879), .B2(n4375), .A(n4374), .ZN(n4376) );
  AOI211_X1 U5507 ( .C1(n4377), .C2(n6456), .A(n4405), .B(n4376), .ZN(n4378)
         );
  OAI21_X1 U5508 ( .B1(n4413), .B2(n6161), .A(n4378), .ZN(U2986) );
  INV_X1 U5509 ( .A(n4379), .ZN(n4385) );
  NAND3_X1 U5510 ( .A1(n4382), .A2(n4381), .A3(n3384), .ZN(n4383) );
  OAI211_X1 U5511 ( .C1(n4386), .C2(n4385), .A(n4384), .B(n4383), .ZN(n4387)
         );
  NAND2_X1 U5512 ( .A1(n4387), .A2(n6750), .ZN(n4394) );
  NAND2_X1 U5513 ( .A1(n4388), .A2(n4179), .ZN(n4389) );
  INV_X1 U5514 ( .A(n4512), .ZN(n4510) );
  OAI211_X1 U5515 ( .C1(n4269), .C2(n4389), .A(n2976), .B(n4510), .ZN(n4390)
         );
  INV_X1 U5516 ( .A(n4390), .ZN(n4391) );
  NAND2_X2 U5517 ( .A1(n4394), .A2(n4393), .ZN(n4410) );
  INV_X1 U5518 ( .A(n4482), .ZN(n4398) );
  OAI22_X1 U5519 ( .A1(n4395), .A2(n4269), .B1(n4401), .B2(n3398), .ZN(n4396)
         );
  INV_X1 U5520 ( .A(n4396), .ZN(n4397) );
  NAND4_X1 U5521 ( .A1(n4398), .A2(n4397), .A3(n4964), .A4(n4447), .ZN(n4399)
         );
  INV_X1 U5522 ( .A(n5464), .ZN(n4406) );
  OAI21_X1 U5523 ( .B1(n4401), .B2(n4400), .A(n4973), .ZN(n4402) );
  INV_X1 U5524 ( .A(n4410), .ZN(n4403) );
  NAND2_X1 U5525 ( .A1(n4403), .A2(n6120), .ZN(n4440) );
  NAND2_X1 U5526 ( .A1(n4410), .A2(n4950), .ZN(n6096) );
  AOI21_X1 U5527 ( .B1(n4440), .B2(n6096), .A(n6074), .ZN(n4404) );
  AOI211_X1 U5528 ( .C1(n4406), .C2(n6534), .A(n4405), .B(n4404), .ZN(n4412)
         );
  INV_X1 U5529 ( .A(n4407), .ZN(n4408) );
  NAND2_X1 U5530 ( .A1(n4410), .A2(n4408), .ZN(n6075) );
  INV_X1 U5531 ( .A(n6075), .ZN(n4411) );
  NAND2_X1 U5532 ( .A1(n4443), .A2(n6074), .ZN(n4439) );
  OAI211_X1 U5533 ( .C1(n4413), .C2(n6483), .A(n4412), .B(n4439), .ZN(U3018)
         );
  AOI222_X1 U5534 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6359), .B1(n6385), .B2(
        DATAO_REG_17__SCAN_IN), .C1(n6390), .C2(UWORD_REG_1__SCAN_IN), .ZN(
        n4414) );
  INV_X1 U5535 ( .A(n4414), .ZN(U2906) );
  AOI222_X1 U5536 ( .A1(EAX_REG_16__SCAN_IN), .A2(n6359), .B1(n6385), .B2(
        DATAO_REG_16__SCAN_IN), .C1(n6390), .C2(UWORD_REG_0__SCAN_IN), .ZN(
        n4415) );
  INV_X1 U5537 ( .A(n4415), .ZN(U2907) );
  AOI222_X1 U5538 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6359), .B1(n6385), .B2(
        DATAO_REG_27__SCAN_IN), .C1(n6390), .C2(UWORD_REG_11__SCAN_IN), .ZN(
        n4416) );
  INV_X1 U5539 ( .A(n4416), .ZN(U2896) );
  AOI222_X1 U5540 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6359), .B1(n6385), .B2(
        DATAO_REG_24__SCAN_IN), .C1(n6390), .C2(UWORD_REG_8__SCAN_IN), .ZN(
        n4417) );
  INV_X1 U5541 ( .A(n4417), .ZN(U2899) );
  AOI222_X1 U5542 ( .A1(EAX_REG_18__SCAN_IN), .A2(n6359), .B1(n6385), .B2(
        DATAO_REG_18__SCAN_IN), .C1(n6390), .C2(UWORD_REG_2__SCAN_IN), .ZN(
        n4418) );
  INV_X1 U5543 ( .A(n4418), .ZN(U2905) );
  AOI222_X1 U5544 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6359), .B1(n6385), .B2(
        DATAO_REG_28__SCAN_IN), .C1(n6390), .C2(UWORD_REG_12__SCAN_IN), .ZN(
        n4419) );
  INV_X1 U5545 ( .A(n4419), .ZN(U2895) );
  AOI222_X1 U5546 ( .A1(EAX_REG_22__SCAN_IN), .A2(n6359), .B1(n6385), .B2(
        DATAO_REG_22__SCAN_IN), .C1(n6390), .C2(UWORD_REG_6__SCAN_IN), .ZN(
        n4420) );
  INV_X1 U5547 ( .A(n4420), .ZN(U2901) );
  AOI222_X1 U5548 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6359), .B1(n6390), .B2(
        UWORD_REG_4__SCAN_IN), .C1(DATAO_REG_20__SCAN_IN), .C2(n6385), .ZN(
        n4421) );
  INV_X1 U5549 ( .A(n4421), .ZN(U2903) );
  OR2_X1 U5550 ( .A1(n4423), .A2(n4422), .ZN(n4425) );
  NAND2_X1 U5551 ( .A1(n4425), .A2(n4424), .ZN(n6529) );
  INV_X1 U5552 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4430) );
  INV_X1 U5553 ( .A(n4426), .ZN(n4427) );
  OAI21_X1 U5554 ( .B1(n4429), .B2(n4428), .A(n4427), .ZN(n6451) );
  OAI222_X1 U5555 ( .A1(n6529), .A2(n5519), .B1(n6335), .B2(n4430), .C1(n6451), 
        .C2(n5521), .ZN(U2857) );
  INV_X2 U5556 ( .A(n4495), .ZN(n4849) );
  XNOR2_X1 U5557 ( .A(n4619), .B(n4618), .ZN(n4433) );
  OAI211_X1 U5558 ( .C1(n6796), .C2(n4433), .A(n4431), .B(n4432), .ZN(n4434)
         );
  AOI21_X1 U5559 ( .B1(n4849), .B2(n3920), .A(n4434), .ZN(n4624) );
  NAND2_X1 U5560 ( .A1(n4437), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4435)
         );
  INV_X1 U5561 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U5562 ( .A1(n4435), .A2(n5189), .ZN(n4438) );
  AND2_X1 U5563 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5564 ( .A1(n4437), .A2(n4436), .ZN(n4625) );
  NAND2_X1 U5565 ( .A1(n4438), .A2(n4625), .ZN(n4623) );
  XNOR2_X1 U5566 ( .A(n4624), .B(n4623), .ZN(n4680) );
  NAND2_X1 U5567 ( .A1(n4440), .A2(n4439), .ZN(n4668) );
  INV_X1 U5568 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6782) );
  NOR2_X1 U5569 ( .A1(n6120), .A2(n6782), .ZN(n4677) );
  INV_X1 U5570 ( .A(n5459), .ZN(n4441) );
  NOR2_X1 U5571 ( .A1(n6121), .A2(n4441), .ZN(n4442) );
  AOI211_X1 U5572 ( .C1(INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n4668), .A(n4677), 
        .B(n4442), .ZN(n4445) );
  NAND2_X1 U5573 ( .A1(n6081), .A2(n6096), .ZN(n6496) );
  INV_X1 U5574 ( .A(n6496), .ZN(n6119) );
  AND2_X1 U5575 ( .A1(n6096), .A2(n6074), .ZN(n4667) );
  OR3_X1 U5576 ( .A1(n6119), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4667), 
        .ZN(n4444) );
  OAI211_X1 U5577 ( .C1(n4680), .C2(n6483), .A(n4445), .B(n4444), .ZN(U3017)
         );
  NAND2_X1 U5578 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6162), .ZN(n4479) );
  NAND2_X1 U5579 ( .A1(n4448), .A2(n4447), .ZN(n4470) );
  INV_X1 U5580 ( .A(n4470), .ZN(n4457) );
  INV_X1 U5581 ( .A(n4449), .ZN(n5257) );
  NAND2_X1 U5582 ( .A1(n5257), .A2(n5264), .ZN(n4464) );
  XNOR2_X1 U5583 ( .A(n4464), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4456)
         );
  NAND2_X1 U5584 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4450) );
  XNOR2_X1 U5585 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n4450), .ZN(n4454)
         );
  INV_X1 U5586 ( .A(n4467), .ZN(n4453) );
  AOI211_X1 U5587 ( .C1(n4452), .C2(n5257), .A(n4451), .B(n3824), .ZN(n6130)
         );
  AOI22_X1 U5588 ( .A1(n4950), .A2(n4454), .B1(n4453), .B2(n6130), .ZN(n4455)
         );
  OAI21_X1 U5589 ( .B1(n4457), .B2(n4456), .A(n4455), .ZN(n4458) );
  AOI21_X1 U5590 ( .B1(n2977), .B2(n4946), .A(n4458), .ZN(n6134) );
  NAND2_X1 U5591 ( .A1(n4954), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4459) );
  OAI21_X1 U5592 ( .B1(n4954), .B2(n6134), .A(n4459), .ZN(n4961) );
  INV_X1 U5593 ( .A(n4954), .ZN(n4473) );
  OR2_X1 U5594 ( .A1(n4461), .A2(n4462), .ZN(n4472) );
  NAND2_X1 U5595 ( .A1(n4449), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U5596 ( .A1(n4464), .A2(n4463), .ZN(n4469) );
  XNOR2_X1 U5597 ( .A(n5264), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4465)
         );
  NAND2_X1 U5598 ( .A1(n4950), .A2(n4465), .ZN(n4466) );
  OAI21_X1 U5599 ( .B1(n4469), .B2(n4467), .A(n4466), .ZN(n4468) );
  AOI21_X1 U5600 ( .B1(n4470), .B2(n4469), .A(n4468), .ZN(n4471) );
  NAND2_X1 U5601 ( .A1(n4472), .A2(n4471), .ZN(n5261) );
  NAND2_X1 U5602 ( .A1(n4473), .A2(n5261), .ZN(n4475) );
  NAND2_X1 U5603 ( .A1(n4954), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4474) );
  INV_X1 U5604 ( .A(n4959), .ZN(n4476) );
  NAND3_X1 U5605 ( .A1(n4961), .A2(n6747), .A3(n4476), .ZN(n4477) );
  OAI21_X1 U5606 ( .B1(n4479), .B2(n4478), .A(n4477), .ZN(n4968) );
  INV_X1 U5607 ( .A(n4480), .ZN(n4481) );
  NAND2_X1 U5608 ( .A1(n4968), .A2(n4481), .ZN(n4491) );
  MUX2_X1 U5609 ( .A(n4954), .B(n6162), .S(STATE2_REG_1__SCAN_IN), .Z(n4484)
         );
  AND2_X1 U5610 ( .A1(n4482), .A2(n6747), .ZN(n4483) );
  AOI22_X1 U5611 ( .A1(n4484), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(n6301), .B2(n4483), .ZN(n4966) );
  AND2_X1 U5612 ( .A1(n4966), .A2(n6162), .ZN(n4485) );
  AOI21_X1 U5613 ( .B1(n4491), .B2(n4485), .A(n6767), .ZN(n4489) );
  INV_X1 U5614 ( .A(n6797), .ZN(n4975) );
  INV_X1 U5615 ( .A(n4490), .ZN(n4486) );
  NAND2_X1 U5616 ( .A1(n4975), .A2(n4486), .ZN(n4487) );
  AND3_X1 U5617 ( .A1(n4491), .A2(n4490), .A3(n4966), .ZN(n4976) );
  NOR2_X1 U5618 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6747), .ZN(n4497) );
  OAI22_X1 U5619 ( .A1(n4858), .A2(n6678), .B1(n4497), .B2(n4866), .ZN(n4493)
         );
  OAI21_X1 U5620 ( .B1(n4976), .B2(n4493), .A(n6778), .ZN(n4494) );
  OAI21_X1 U5621 ( .B1(n6778), .B2(n6626), .A(n4494), .ZN(U3465) );
  NOR2_X1 U5622 ( .A1(n4764), .A2(n6160), .ZN(n6679) );
  XNOR2_X1 U5623 ( .A(n6679), .B(n6551), .ZN(n4498) );
  INV_X1 U5624 ( .A(n4461), .ZN(n5446) );
  INV_X1 U5625 ( .A(n4497), .ZN(n6777) );
  AOI22_X1 U5626 ( .A1(n4498), .A2(n6774), .B1(n5446), .B2(n6777), .ZN(n4500)
         );
  NAND2_X1 U5627 ( .A1(n6781), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4499) );
  OAI21_X1 U5628 ( .B1(n6781), .B2(n4500), .A(n4499), .ZN(U3463) );
  AOI211_X1 U5629 ( .C1(n6160), .C2(n4764), .A(n6678), .B(n6679), .ZN(n4502)
         );
  AOI21_X1 U5630 ( .B1(n5452), .B2(n6777), .A(n4502), .ZN(n4504) );
  NAND2_X1 U5631 ( .A1(n6781), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4503) );
  OAI21_X1 U5632 ( .B1(n6781), .B2(n4504), .A(n4503), .ZN(U3464) );
  NOR2_X1 U5633 ( .A1(n4505), .A2(n3910), .ZN(n4506) );
  AND2_X1 U5634 ( .A1(n4510), .A2(n4509), .ZN(n4511) );
  INV_X1 U5635 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6389) );
  OAI222_X1 U5636 ( .A1(n6451), .A2(n6148), .B1(n6349), .B2(n4514), .C1(n6354), 
        .C2(n6389), .ZN(U2889) );
  INV_X1 U5637 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6393) );
  OAI222_X1 U5638 ( .A1(n5463), .A2(n6148), .B1(n6349), .B2(n4515), .C1(n6354), 
        .C2(n6393), .ZN(U2890) );
  XNOR2_X1 U5639 ( .A(n4426), .B(n4516), .ZN(n6330) );
  INV_X1 U5640 ( .A(DATAI_3_), .ZN(n4517) );
  INV_X1 U5641 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6387) );
  OAI222_X1 U5642 ( .A1(n6330), .A2(n6148), .B1(n6349), .B2(n4517), .C1(n6354), 
        .C2(n6387), .ZN(U2888) );
  INV_X1 U5643 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4518) );
  OAI222_X1 U5644 ( .A1(n5470), .A2(n6148), .B1(n6349), .B2(n4519), .C1(n6354), 
        .C2(n4518), .ZN(U2891) );
  NAND2_X1 U5645 ( .A1(n4849), .A2(n4520), .ZN(n4521) );
  INV_X1 U5646 ( .A(n4531), .ZN(n4522) );
  OAI21_X1 U5647 ( .B1(n4522), .B2(n5886), .A(n4982), .ZN(n4526) );
  AND2_X1 U5648 ( .A1(n3466), .A2(n2977), .ZN(n4725) );
  INV_X1 U5649 ( .A(n4523), .ZN(n4567) );
  AOI21_X1 U5650 ( .B1(n4725), .B2(n4765), .A(n4567), .ZN(n4528) );
  NAND2_X1 U5651 ( .A1(n6626), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4524) );
  OAI21_X1 U5652 ( .B1(n6774), .B2(n4684), .A(n6687), .ZN(n4525) );
  INV_X1 U5653 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5807) );
  INV_X1 U5654 ( .A(n4684), .ZN(n4527) );
  OAI22_X1 U5655 ( .A1(n4528), .A2(n6678), .B1(n4686), .B2(n4527), .ZN(n4568)
         );
  INV_X1 U5656 ( .A(n6705), .ZN(n6642) );
  INV_X1 U5657 ( .A(n5137), .ZN(n6700) );
  AOI22_X1 U5658 ( .A1(n4568), .A2(n6642), .B1(n4567), .B2(n6700), .ZN(n4534)
         );
  INV_X1 U5659 ( .A(DATAI_26_), .ZN(n4530) );
  OR2_X1 U5660 ( .A1(n5886), .A2(n4530), .ZN(n6603) );
  INV_X1 U5661 ( .A(n6603), .ZN(n6702) );
  INV_X1 U5662 ( .A(DATAI_18_), .ZN(n4532) );
  OR2_X1 U5663 ( .A1(n5886), .A2(n4532), .ZN(n6645) );
  INV_X1 U5664 ( .A(n6645), .ZN(n6701) );
  AOI22_X1 U5665 ( .A1(n6702), .A2(n4688), .B1(n4938), .B2(n6701), .ZN(n4533)
         );
  OAI211_X1 U5666 ( .C1(n4574), .C2(n5807), .A(n4534), .B(n4533), .ZN(U3142)
         );
  INV_X1 U5667 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4540) );
  INV_X1 U5668 ( .A(n6711), .ZN(n6646) );
  INV_X1 U5669 ( .A(n5141), .ZN(n6706) );
  AOI22_X1 U5670 ( .A1(n4568), .A2(n6646), .B1(n4567), .B2(n6706), .ZN(n4539)
         );
  INV_X1 U5671 ( .A(DATAI_27_), .ZN(n4536) );
  INV_X1 U5672 ( .A(n6606), .ZN(n6708) );
  INV_X1 U5673 ( .A(DATAI_19_), .ZN(n4537) );
  OR2_X1 U5674 ( .A1(n5886), .A2(n4537), .ZN(n6649) );
  INV_X1 U5675 ( .A(n6649), .ZN(n6707) );
  AOI22_X1 U5676 ( .A1(n6708), .A2(n4688), .B1(n4938), .B2(n6707), .ZN(n4538)
         );
  OAI211_X1 U5677 ( .C1(n4574), .C2(n4540), .A(n4539), .B(n4538), .ZN(U3143)
         );
  INV_X1 U5678 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4546) );
  INV_X1 U5679 ( .A(n6733), .ZN(n6662) );
  INV_X1 U5680 ( .A(n5145), .ZN(n6727) );
  AOI22_X1 U5681 ( .A1(n4568), .A2(n6662), .B1(n4567), .B2(n6727), .ZN(n4545)
         );
  INV_X1 U5682 ( .A(DATAI_30_), .ZN(n4542) );
  OR2_X1 U5683 ( .A1(n5886), .A2(n4542), .ZN(n6613) );
  INV_X1 U5684 ( .A(n6613), .ZN(n6730) );
  INV_X1 U5685 ( .A(DATAI_22_), .ZN(n4543) );
  INV_X1 U5686 ( .A(n6665), .ZN(n6728) );
  AOI22_X1 U5687 ( .A1(n6730), .A2(n4688), .B1(n4938), .B2(n6728), .ZN(n4544)
         );
  OAI211_X1 U5688 ( .C1(n4574), .C2(n4546), .A(n4545), .B(n4544), .ZN(U3146)
         );
  INV_X1 U5689 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4550) );
  INV_X1 U5690 ( .A(n6725), .ZN(n6657) );
  INV_X1 U5691 ( .A(n6719), .ZN(n6656) );
  AOI22_X1 U5692 ( .A1(n4568), .A2(n6657), .B1(n4567), .B2(n6656), .ZN(n4549)
         );
  INV_X1 U5693 ( .A(DATAI_29_), .ZN(n4547) );
  OR2_X1 U5694 ( .A1(n5886), .A2(n4547), .ZN(n6720) );
  INV_X1 U5695 ( .A(n6720), .ZN(n6658) );
  INV_X1 U5696 ( .A(DATAI_21_), .ZN(n5719) );
  OR2_X1 U5697 ( .A1(n5886), .A2(n5719), .ZN(n6661) );
  INV_X1 U5698 ( .A(n6661), .ZN(n6722) );
  AOI22_X1 U5699 ( .A1(n6658), .A2(n4688), .B1(n4938), .B2(n6722), .ZN(n4548)
         );
  OAI211_X1 U5700 ( .C1(n4574), .C2(n4550), .A(n4549), .B(n4548), .ZN(U3145)
         );
  INV_X1 U5701 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4555) );
  INV_X1 U5702 ( .A(n6718), .ZN(n6651) );
  INV_X1 U5703 ( .A(n6712), .ZN(n6650) );
  AOI22_X1 U5704 ( .A1(n4568), .A2(n6651), .B1(n4567), .B2(n6650), .ZN(n4554)
         );
  INV_X1 U5705 ( .A(DATAI_28_), .ZN(n4551) );
  OR2_X1 U5706 ( .A1(n5886), .A2(n4551), .ZN(n6713) );
  INV_X1 U5707 ( .A(n6713), .ZN(n6652) );
  INV_X1 U5708 ( .A(DATAI_20_), .ZN(n4552) );
  OR2_X1 U5709 ( .A1(n5886), .A2(n4552), .ZN(n6655) );
  AOI22_X1 U5710 ( .A1(n6652), .A2(n4688), .B1(n4938), .B2(n6715), .ZN(n4553)
         );
  OAI211_X1 U5711 ( .C1(n4574), .C2(n4555), .A(n4554), .B(n4553), .ZN(U3144)
         );
  INV_X1 U5712 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4560) );
  INV_X1 U5713 ( .A(n6744), .ZN(n6668) );
  INV_X1 U5714 ( .A(n6735), .ZN(n6667) );
  AOI22_X1 U5715 ( .A1(n4568), .A2(n6668), .B1(n4567), .B2(n6667), .ZN(n4559)
         );
  INV_X1 U5716 ( .A(DATAI_31_), .ZN(n4556) );
  OR2_X1 U5717 ( .A1(n5886), .A2(n4556), .ZN(n6736) );
  INV_X1 U5718 ( .A(n6736), .ZN(n6671) );
  INV_X1 U5719 ( .A(DATAI_23_), .ZN(n4557) );
  OR2_X1 U5720 ( .A1(n5886), .A2(n4557), .ZN(n6676) );
  AOI22_X1 U5721 ( .A1(n6671), .A2(n4688), .B1(n4938), .B2(n6740), .ZN(n4558)
         );
  OAI211_X1 U5722 ( .C1(n4574), .C2(n4560), .A(n4559), .B(n4558), .ZN(U3147)
         );
  INV_X1 U5723 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4565) );
  INV_X1 U5724 ( .A(n6693), .ZN(n6628) );
  OR2_X1 U5725 ( .A1(n4566), .A2(n4561), .ZN(n5158) );
  AOI22_X1 U5726 ( .A1(n4568), .A2(n6628), .B1(n4567), .B2(n6683), .ZN(n4564)
         );
  INV_X1 U5727 ( .A(DATAI_24_), .ZN(n4562) );
  OR2_X1 U5728 ( .A1(n5886), .A2(n4562), .ZN(n6597) );
  INV_X1 U5729 ( .A(n6597), .ZN(n6690) );
  OR2_X1 U5730 ( .A1(n5886), .A2(n5812), .ZN(n6637) );
  INV_X1 U5731 ( .A(n6637), .ZN(n6684) );
  AOI22_X1 U5732 ( .A1(n6690), .A2(n4688), .B1(n4938), .B2(n6684), .ZN(n4563)
         );
  OAI211_X1 U5733 ( .C1(n4574), .C2(n4565), .A(n4564), .B(n4563), .ZN(U3140)
         );
  INV_X1 U5734 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4573) );
  INV_X1 U5735 ( .A(n6699), .ZN(n6638) );
  INV_X1 U5736 ( .A(n5164), .ZN(n6694) );
  AOI22_X1 U5737 ( .A1(n4568), .A2(n6638), .B1(n4567), .B2(n6694), .ZN(n4572)
         );
  INV_X1 U5738 ( .A(DATAI_25_), .ZN(n4569) );
  OR2_X1 U5739 ( .A1(n5886), .A2(n4569), .ZN(n6600) );
  INV_X1 U5740 ( .A(n6600), .ZN(n6696) );
  INV_X1 U5741 ( .A(DATAI_17_), .ZN(n4570) );
  AOI22_X1 U5742 ( .A1(n6696), .A2(n4688), .B1(n4938), .B2(n6695), .ZN(n4571)
         );
  OAI211_X1 U5743 ( .C1(n4574), .C2(n4573), .A(n4572), .B(n4571), .ZN(U3141)
         );
  INV_X1 U5744 ( .A(n4575), .ZN(n4759) );
  AOI21_X1 U5745 ( .B1(n4577), .B2(n4576), .A(n4759), .ZN(n6313) );
  INV_X1 U5746 ( .A(n6313), .ZN(n4617) );
  INV_X1 U5747 ( .A(DATAI_4_), .ZN(n4578) );
  INV_X1 U5748 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6384) );
  OAI222_X1 U5749 ( .A1(n4617), .A2(n6148), .B1(n6349), .B2(n4578), .C1(n6354), 
        .C2(n6384), .ZN(U2887) );
  NAND2_X1 U5750 ( .A1(n4520), .A2(n4764), .ZN(n4579) );
  NAND2_X1 U5751 ( .A1(n4584), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6550) );
  AND2_X1 U5752 ( .A1(n4581), .A2(n4580), .ZN(n5091) );
  AND2_X1 U5753 ( .A1(n5091), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4585)
         );
  AOI21_X1 U5754 ( .B1(n4725), .B2(n5094), .A(n4585), .ZN(n4587) );
  INV_X1 U5755 ( .A(n4587), .ZN(n4582) );
  INV_X1 U5756 ( .A(n4584), .ZN(n4583) );
  INV_X1 U5757 ( .A(n4585), .ZN(n4610) );
  OAI22_X1 U5758 ( .A1(n4690), .A2(n6661), .B1(n6719), .B2(n4610), .ZN(n4586)
         );
  AOI21_X1 U5759 ( .B1(n6658), .B2(n5120), .A(n4586), .ZN(n4591) );
  NAND2_X1 U5760 ( .A1(n4588), .A2(n4587), .ZN(n4589) );
  NAND2_X1 U5761 ( .A1(n4612), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4590)
         );
  OAI211_X1 U5762 ( .C1(n4615), .C2(n6725), .A(n4591), .B(n4590), .ZN(U3129)
         );
  OAI22_X1 U5763 ( .A1(n4690), .A2(n6641), .B1(n5164), .B2(n4610), .ZN(n4592)
         );
  AOI21_X1 U5764 ( .B1(n6696), .B2(n5120), .A(n4592), .ZN(n4594) );
  NAND2_X1 U5765 ( .A1(n4612), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4593)
         );
  OAI211_X1 U5766 ( .C1(n4615), .C2(n6699), .A(n4594), .B(n4593), .ZN(U3125)
         );
  OAI22_X1 U5767 ( .A1(n4690), .A2(n6649), .B1(n5141), .B2(n4610), .ZN(n4595)
         );
  AOI21_X1 U5768 ( .B1(n6708), .B2(n5120), .A(n4595), .ZN(n4597) );
  NAND2_X1 U5769 ( .A1(n4612), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4596)
         );
  OAI211_X1 U5770 ( .C1(n4615), .C2(n6711), .A(n4597), .B(n4596), .ZN(U3127)
         );
  OAI22_X1 U5771 ( .A1(n4690), .A2(n6676), .B1(n6735), .B2(n4610), .ZN(n4598)
         );
  AOI21_X1 U5772 ( .B1(n6671), .B2(n5120), .A(n4598), .ZN(n4600) );
  NAND2_X1 U5773 ( .A1(n4612), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4599)
         );
  OAI211_X1 U5774 ( .C1(n4615), .C2(n6744), .A(n4600), .B(n4599), .ZN(U3131)
         );
  OAI22_X1 U5775 ( .A1(n4690), .A2(n6655), .B1(n6712), .B2(n4610), .ZN(n4601)
         );
  AOI21_X1 U5776 ( .B1(n6652), .B2(n5120), .A(n4601), .ZN(n4603) );
  NAND2_X1 U5777 ( .A1(n4612), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4602)
         );
  OAI211_X1 U5778 ( .C1(n4615), .C2(n6718), .A(n4603), .B(n4602), .ZN(U3128)
         );
  OAI22_X1 U5779 ( .A1(n4690), .A2(n6645), .B1(n5137), .B2(n4610), .ZN(n4604)
         );
  AOI21_X1 U5780 ( .B1(n6702), .B2(n5120), .A(n4604), .ZN(n4606) );
  NAND2_X1 U5781 ( .A1(n4612), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4605)
         );
  OAI211_X1 U5782 ( .C1(n4615), .C2(n6705), .A(n4606), .B(n4605), .ZN(U3126)
         );
  OAI22_X1 U5783 ( .A1(n4690), .A2(n6665), .B1(n5145), .B2(n4610), .ZN(n4607)
         );
  AOI21_X1 U5784 ( .B1(n6730), .B2(n5120), .A(n4607), .ZN(n4609) );
  NAND2_X1 U5785 ( .A1(n4612), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4608)
         );
  OAI211_X1 U5786 ( .C1(n4615), .C2(n6733), .A(n4609), .B(n4608), .ZN(U3130)
         );
  OAI22_X1 U5787 ( .A1(n4690), .A2(n6637), .B1(n5158), .B2(n4610), .ZN(n4611)
         );
  AOI21_X1 U5788 ( .B1(n6690), .B2(n5120), .A(n4611), .ZN(n4614) );
  NAND2_X1 U5789 ( .A1(n4612), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4613)
         );
  OAI211_X1 U5790 ( .C1(n4615), .C2(n6693), .A(n4614), .B(n4613), .ZN(U3124)
         );
  OAI21_X1 U5791 ( .B1(n4616), .B2(n5432), .A(n4663), .ZN(n4666) );
  INV_X1 U5792 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5746) );
  OAI222_X1 U5793 ( .A1(n4666), .A2(n5519), .B1(n6335), .B2(n5746), .C1(n4617), 
        .C2(n5521), .ZN(U2855) );
  NAND2_X1 U5794 ( .A1(n4619), .A2(n4618), .ZN(n4628) );
  INV_X1 U5795 ( .A(n4620), .ZN(n4627) );
  XNOR2_X1 U5796 ( .A(n4628), .B(n4627), .ZN(n4621) );
  AOI21_X1 U5797 ( .B1(n4621), .B2(n5216), .A(n4254), .ZN(n4622) );
  OR2_X1 U5798 ( .A1(n4624), .A2(n4623), .ZN(n4626) );
  NAND2_X1 U5799 ( .A1(n4628), .A2(n4627), .ZN(n4650) );
  INV_X1 U5800 ( .A(n4649), .ZN(n4629) );
  XNOR2_X1 U5801 ( .A(n4650), .B(n4629), .ZN(n4630) );
  NAND2_X1 U5802 ( .A1(n4630), .A2(n5216), .ZN(n4644) );
  NAND2_X1 U5803 ( .A1(n4644), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4634)
         );
  AND2_X1 U5804 ( .A1(n3920), .A2(n6527), .ZN(n4633) );
  NAND2_X1 U5805 ( .A1(n3535), .A2(n4633), .ZN(n4631) );
  OAI21_X1 U5806 ( .B1(n3535), .B2(n4634), .A(n4631), .ZN(n4632) );
  INV_X1 U5807 ( .A(n4633), .ZN(n4637) );
  INV_X1 U5808 ( .A(n4634), .ZN(n4635) );
  NAND2_X1 U5809 ( .A1(n3535), .A2(n4635), .ZN(n4636) );
  OAI21_X1 U5810 ( .B1(n3535), .B2(n4637), .A(n4636), .ZN(n4639) );
  INV_X1 U5811 ( .A(n4520), .ZN(n4638) );
  NAND2_X1 U5812 ( .A1(n3919), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4640)
         );
  MUX2_X1 U5813 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .B(n4640), .S(n4644), 
        .Z(n4641) );
  NAND2_X1 U5814 ( .A1(n4642), .A2(n3920), .ZN(n4645) );
  NAND2_X1 U5815 ( .A1(n4645), .A2(n4644), .ZN(n4646) );
  NAND2_X1 U5816 ( .A1(n4646), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4647)
         );
  NAND2_X1 U5817 ( .A1(n4648), .A2(n3920), .ZN(n4653) );
  NAND2_X1 U5818 ( .A1(n4650), .A2(n4649), .ZN(n5023) );
  XNOR2_X1 U5819 ( .A(n5023), .B(n5021), .ZN(n4651) );
  NAND2_X1 U5820 ( .A1(n4651), .A2(n5216), .ZN(n4652) );
  NAND2_X1 U5821 ( .A1(n4653), .A2(n4652), .ZN(n5017) );
  INV_X1 U5822 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4670) );
  XNOR2_X1 U5823 ( .A(n5017), .B(n4670), .ZN(n4654) );
  NAND2_X1 U5824 ( .A1(n4655), .A2(n4654), .ZN(n5019) );
  OAI21_X1 U5825 ( .B1(n4655), .B2(n4654), .A(n5019), .ZN(n4675) );
  NAND2_X1 U5826 ( .A1(n6313), .A2(n6456), .ZN(n4660) );
  AND2_X1 U5827 ( .A1(n6490), .A2(REIP_REG_4__SCAN_IN), .ZN(n4673) );
  NOR2_X1 U5828 ( .A1(n5879), .A2(n4657), .ZN(n4658) );
  AOI211_X1 U5829 ( .C1(n5882), .C2(n6312), .A(n4673), .B(n4658), .ZN(n4659)
         );
  OAI211_X1 U5830 ( .C1(n4675), .C2(n6161), .A(n4660), .B(n4659), .ZN(U2982)
         );
  XNOR2_X1 U5831 ( .A(n4575), .B(n4661), .ZN(n6437) );
  INV_X1 U5832 ( .A(n6437), .ZN(n4682) );
  AOI21_X1 U5833 ( .B1(n4664), .B2(n4663), .A(n4662), .ZN(n6510) );
  AOI22_X1 U5834 ( .A1(n6331), .A2(n6510), .B1(EBX_REG_5__SCAN_IN), .B2(n5504), 
        .ZN(n4665) );
  OAI21_X1 U5835 ( .B1(n4682), .B2(n5521), .A(n4665), .ZN(U2854) );
  INV_X1 U5836 ( .A(n4666), .ZN(n6304) );
  NAND2_X1 U5837 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6511) );
  INV_X1 U5838 ( .A(n6511), .ZN(n5891) );
  OR2_X2 U5839 ( .A1(n6116), .A2(n4667), .ZN(n6539) );
  NAND2_X1 U5840 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6512) );
  OAI21_X1 U5841 ( .B1(n6539), .B2(n6512), .A(n6531), .ZN(n6521) );
  NAND2_X1 U5842 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U5843 ( .A1(n6540), .A2(n6530), .ZN(n6522) );
  OAI211_X1 U5844 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6521), .B(n6522), .ZN(n4671) );
  NOR2_X1 U5845 ( .A1(n6531), .A2(n6522), .ZN(n6533) );
  INV_X1 U5846 ( .A(n6512), .ZN(n4669) );
  NAND2_X1 U5847 ( .A1(n6531), .A2(n4668), .ZN(n6114) );
  OAI21_X1 U5848 ( .B1(n6116), .B2(n4669), .A(n6114), .ZN(n6538) );
  NOR2_X1 U5849 ( .A1(n6533), .A2(n6538), .ZN(n6528) );
  OAI22_X1 U5850 ( .A1(n5891), .A2(n4671), .B1(n6528), .B2(n4670), .ZN(n4672)
         );
  AOI211_X1 U5851 ( .C1(n6534), .C2(n6304), .A(n4673), .B(n4672), .ZN(n4674)
         );
  OAI21_X1 U5852 ( .B1(n6483), .B2(n4675), .A(n4674), .ZN(U3014) );
  INV_X1 U5853 ( .A(n5463), .ZN(n4678) );
  MUX2_X1 U5854 ( .A(n5882), .B(n6450), .S(PHYADDRPOINTER_REG_1__SCAN_IN), .Z(
        n4676) );
  AOI211_X1 U5855 ( .C1(n4678), .C2(n6456), .A(n4677), .B(n4676), .ZN(n4679)
         );
  OAI21_X1 U5856 ( .B1(n4680), .B2(n6161), .A(n4679), .ZN(U2985) );
  INV_X1 U5857 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6382) );
  INV_X1 U5858 ( .A(DATAI_5_), .ZN(n4681) );
  OAI222_X1 U5859 ( .A1(n6148), .A2(n4682), .B1(n6354), .B2(n6382), .C1(n4681), 
        .C2(n6349), .ZN(U2886) );
  OR2_X1 U5860 ( .A1(n2977), .A2(n6678), .ZN(n6625) );
  INV_X1 U5861 ( .A(n6625), .ZN(n4683) );
  AND2_X1 U5862 ( .A1(n6624), .A2(n6774), .ZN(n6629) );
  OAI21_X1 U5863 ( .B1(n4683), .B2(n6629), .A(n4690), .ZN(n4689) );
  NAND2_X1 U5864 ( .A1(n4684), .A2(n6626), .ZN(n4715) );
  NAND2_X1 U5865 ( .A1(n6780), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6555) );
  INV_X1 U5866 ( .A(n6555), .ZN(n5054) );
  NAND2_X1 U5867 ( .A1(n5051), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4685) );
  OR2_X1 U5868 ( .A1(n4691), .A2(n4686), .ZN(n6592) );
  OAI211_X1 U5869 ( .C1(n4765), .C2(n4982), .A(n5056), .B(n6592), .ZN(n6630)
         );
  AOI211_X1 U5870 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4715), .A(n5054), .B(
        n6630), .ZN(n4687) );
  NAND2_X1 U5871 ( .A1(n4714), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4695)
         );
  INV_X1 U5872 ( .A(n2977), .ZN(n5128) );
  NOR2_X1 U5873 ( .A1(n5128), .A2(n6678), .ZN(n5136) );
  NAND2_X1 U5874 ( .A1(n4691), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5131) );
  NOR3_X1 U5875 ( .A1(n5131), .A2(n5051), .A3(n6780), .ZN(n4692) );
  AOI21_X1 U5876 ( .B1(n5136), .B2(n4765), .A(n4692), .ZN(n4716) );
  OAI22_X1 U5877 ( .A1(n4716), .A2(n6711), .B1(n5141), .B2(n4715), .ZN(n4693)
         );
  AOI21_X1 U5878 ( .B1(n6708), .B2(n4718), .A(n4693), .ZN(n4694) );
  OAI211_X1 U5879 ( .C1(n4721), .C2(n6649), .A(n4695), .B(n4694), .ZN(U3135)
         );
  NAND2_X1 U5880 ( .A1(n4714), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4698)
         );
  OAI22_X1 U5881 ( .A1(n4716), .A2(n6705), .B1(n5137), .B2(n4715), .ZN(n4696)
         );
  AOI21_X1 U5882 ( .B1(n6702), .B2(n4718), .A(n4696), .ZN(n4697) );
  OAI211_X1 U5883 ( .C1(n4721), .C2(n6645), .A(n4698), .B(n4697), .ZN(U3134)
         );
  NAND2_X1 U5884 ( .A1(n4714), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4701)
         );
  OAI22_X1 U5885 ( .A1(n4716), .A2(n6693), .B1(n5158), .B2(n4715), .ZN(n4699)
         );
  AOI21_X1 U5886 ( .B1(n6690), .B2(n4718), .A(n4699), .ZN(n4700) );
  OAI211_X1 U5887 ( .C1(n4721), .C2(n6637), .A(n4701), .B(n4700), .ZN(U3132)
         );
  NAND2_X1 U5888 ( .A1(n4714), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4704)
         );
  OAI22_X1 U5889 ( .A1(n4716), .A2(n6725), .B1(n6719), .B2(n4715), .ZN(n4702)
         );
  AOI21_X1 U5890 ( .B1(n6658), .B2(n4718), .A(n4702), .ZN(n4703) );
  OAI211_X1 U5891 ( .C1(n4721), .C2(n6661), .A(n4704), .B(n4703), .ZN(U3137)
         );
  NAND2_X1 U5892 ( .A1(n4714), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4707)
         );
  OAI22_X1 U5893 ( .A1(n4716), .A2(n6699), .B1(n5164), .B2(n4715), .ZN(n4705)
         );
  AOI21_X1 U5894 ( .B1(n6696), .B2(n4718), .A(n4705), .ZN(n4706) );
  OAI211_X1 U5895 ( .C1(n4721), .C2(n6641), .A(n4707), .B(n4706), .ZN(U3133)
         );
  NAND2_X1 U5896 ( .A1(n4714), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4710)
         );
  OAI22_X1 U5897 ( .A1(n4716), .A2(n6744), .B1(n6735), .B2(n4715), .ZN(n4708)
         );
  AOI21_X1 U5898 ( .B1(n6671), .B2(n4718), .A(n4708), .ZN(n4709) );
  OAI211_X1 U5899 ( .C1(n4721), .C2(n6676), .A(n4710), .B(n4709), .ZN(U3139)
         );
  NAND2_X1 U5900 ( .A1(n4714), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4713)
         );
  OAI22_X1 U5901 ( .A1(n4716), .A2(n6718), .B1(n6712), .B2(n4715), .ZN(n4711)
         );
  AOI21_X1 U5902 ( .B1(n6652), .B2(n4718), .A(n4711), .ZN(n4712) );
  OAI211_X1 U5903 ( .C1(n4721), .C2(n6655), .A(n4713), .B(n4712), .ZN(U3136)
         );
  NAND2_X1 U5904 ( .A1(n4714), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4720)
         );
  OAI22_X1 U5905 ( .A1(n4716), .A2(n6733), .B1(n5145), .B2(n4715), .ZN(n4717)
         );
  AOI21_X1 U5906 ( .B1(n6730), .B2(n4718), .A(n4717), .ZN(n4719) );
  OAI211_X1 U5907 ( .C1(n4721), .C2(n6665), .A(n4720), .B(n4719), .ZN(U3138)
         );
  AOI21_X1 U5908 ( .B1(n4727), .B2(STATEBS16_REG_SCAN_IN), .A(n6678), .ZN(
        n4730) );
  NAND2_X1 U5909 ( .A1(n4461), .A2(n4722), .ZN(n5127) );
  INV_X1 U5910 ( .A(n5127), .ZN(n5135) );
  NOR2_X1 U5911 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4723) );
  AND2_X1 U5912 ( .A1(n4723), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5129)
         );
  NAND2_X1 U5913 ( .A1(n5129), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4752) );
  INV_X1 U5914 ( .A(n4752), .ZN(n4724) );
  AOI21_X1 U5915 ( .B1(n4725), .B2(n5135), .A(n4724), .ZN(n4729) );
  INV_X1 U5916 ( .A(n4729), .ZN(n4726) );
  OAI22_X1 U5917 ( .A1(n5058), .A2(n6649), .B1(n5141), .B2(n4752), .ZN(n4728)
         );
  AOI21_X1 U5918 ( .B1(n6708), .B2(n5125), .A(n4728), .ZN(n4733) );
  NAND2_X1 U5919 ( .A1(n4730), .A2(n4729), .ZN(n4731) );
  NAND2_X1 U5920 ( .A1(n4754), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4732) );
  OAI211_X1 U5921 ( .C1(n4757), .C2(n6711), .A(n4733), .B(n4732), .ZN(U3095)
         );
  OAI22_X1 U5922 ( .A1(n5058), .A2(n6661), .B1(n6719), .B2(n4752), .ZN(n4734)
         );
  AOI21_X1 U5923 ( .B1(n6658), .B2(n5125), .A(n4734), .ZN(n4736) );
  NAND2_X1 U5924 ( .A1(n4754), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4735) );
  OAI211_X1 U5925 ( .C1(n4757), .C2(n6725), .A(n4736), .B(n4735), .ZN(U3097)
         );
  OAI22_X1 U5926 ( .A1(n5058), .A2(n6655), .B1(n6712), .B2(n4752), .ZN(n4737)
         );
  AOI21_X1 U5927 ( .B1(n6652), .B2(n5125), .A(n4737), .ZN(n4739) );
  NAND2_X1 U5928 ( .A1(n4754), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4738) );
  OAI211_X1 U5929 ( .C1(n4757), .C2(n6718), .A(n4739), .B(n4738), .ZN(U3096)
         );
  OAI22_X1 U5930 ( .A1(n5058), .A2(n6665), .B1(n5145), .B2(n4752), .ZN(n4740)
         );
  AOI21_X1 U5931 ( .B1(n6730), .B2(n5125), .A(n4740), .ZN(n4742) );
  NAND2_X1 U5932 ( .A1(n4754), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4741) );
  OAI211_X1 U5933 ( .C1(n4757), .C2(n6733), .A(n4742), .B(n4741), .ZN(U3098)
         );
  OAI22_X1 U5934 ( .A1(n5058), .A2(n6676), .B1(n6735), .B2(n4752), .ZN(n4743)
         );
  AOI21_X1 U5935 ( .B1(n6671), .B2(n5125), .A(n4743), .ZN(n4745) );
  NAND2_X1 U5936 ( .A1(n4754), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4744) );
  OAI211_X1 U5937 ( .C1(n4757), .C2(n6744), .A(n4745), .B(n4744), .ZN(U3099)
         );
  OAI22_X1 U5938 ( .A1(n5058), .A2(n6645), .B1(n5137), .B2(n4752), .ZN(n4746)
         );
  AOI21_X1 U5939 ( .B1(n6702), .B2(n5125), .A(n4746), .ZN(n4748) );
  NAND2_X1 U5940 ( .A1(n4754), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4747) );
  OAI211_X1 U5941 ( .C1(n4757), .C2(n6705), .A(n4748), .B(n4747), .ZN(U3094)
         );
  OAI22_X1 U5942 ( .A1(n5058), .A2(n6637), .B1(n5158), .B2(n4752), .ZN(n4749)
         );
  AOI21_X1 U5943 ( .B1(n6690), .B2(n5125), .A(n4749), .ZN(n4751) );
  NAND2_X1 U5944 ( .A1(n4754), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4750) );
  OAI211_X1 U5945 ( .C1(n4757), .C2(n6693), .A(n4751), .B(n4750), .ZN(U3092)
         );
  OAI22_X1 U5946 ( .A1(n5058), .A2(n6641), .B1(n5164), .B2(n4752), .ZN(n4753)
         );
  AOI21_X1 U5947 ( .B1(n6696), .B2(n5125), .A(n4753), .ZN(n4756) );
  NAND2_X1 U5948 ( .A1(n4754), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4755) );
  OAI211_X1 U5949 ( .C1(n4757), .C2(n6699), .A(n4756), .B(n4755), .ZN(U3093)
         );
  AOI21_X1 U5950 ( .B1(n4759), .B2(n4661), .A(n4758), .ZN(n4761) );
  NOR2_X1 U5951 ( .A1(n4761), .A2(n4760), .ZN(n5426) );
  INV_X1 U5952 ( .A(n5426), .ZN(n4797) );
  XOR2_X1 U5953 ( .A(n4662), .B(n4762), .Z(n6499) );
  AOI22_X1 U5954 ( .A1(n6331), .A2(n6499), .B1(n5504), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4763) );
  OAI21_X1 U5955 ( .B1(n4797), .B2(n5521), .A(n4763), .ZN(U2853) );
  NAND3_X1 U5956 ( .A1(n4765), .A2(n5087), .A3(n3466), .ZN(n4766) );
  AOI21_X1 U5957 ( .B1(n4766), .B2(n4791), .A(n6678), .ZN(n4767) );
  AOI21_X1 U5958 ( .B1(n6627), .B2(STATE2_REG_2__SCAN_IN), .A(n4767), .ZN(
        n4792) );
  OAI22_X1 U5959 ( .A1(n4792), .A2(n6693), .B1(n4791), .B2(n5158), .ZN(n4768)
         );
  AOI21_X1 U5960 ( .B1(n6684), .B2(n5167), .A(n4768), .ZN(n4772) );
  INV_X1 U5961 ( .A(n4803), .ZN(n4769) );
  NAND2_X1 U5962 ( .A1(n4769), .A2(n6679), .ZN(n6772) );
  NOR2_X1 U5963 ( .A1(n6772), .A2(n6678), .ZN(n4770) );
  NAND2_X1 U5964 ( .A1(n4794), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4771) );
  OAI211_X1 U5965 ( .C1(n6675), .C2(n6597), .A(n4772), .B(n4771), .ZN(U3076)
         );
  OAI22_X1 U5966 ( .A1(n4792), .A2(n6725), .B1(n4791), .B2(n6719), .ZN(n4773)
         );
  AOI21_X1 U5967 ( .B1(n6722), .B2(n5167), .A(n4773), .ZN(n4775) );
  NAND2_X1 U5968 ( .A1(n4794), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4774) );
  OAI211_X1 U5969 ( .C1(n6675), .C2(n6720), .A(n4775), .B(n4774), .ZN(U3081)
         );
  OAI22_X1 U5970 ( .A1(n4792), .A2(n6699), .B1(n4791), .B2(n5164), .ZN(n4776)
         );
  AOI21_X1 U5971 ( .B1(n6695), .B2(n5167), .A(n4776), .ZN(n4778) );
  NAND2_X1 U5972 ( .A1(n4794), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4777) );
  OAI211_X1 U5973 ( .C1(n6675), .C2(n6600), .A(n4778), .B(n4777), .ZN(U3077)
         );
  OAI22_X1 U5974 ( .A1(n4792), .A2(n6705), .B1(n4791), .B2(n5137), .ZN(n4779)
         );
  AOI21_X1 U5975 ( .B1(n6701), .B2(n5167), .A(n4779), .ZN(n4781) );
  NAND2_X1 U5976 ( .A1(n4794), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4780) );
  OAI211_X1 U5977 ( .C1(n6675), .C2(n6603), .A(n4781), .B(n4780), .ZN(U3078)
         );
  OAI22_X1 U5978 ( .A1(n4792), .A2(n6733), .B1(n4791), .B2(n5145), .ZN(n4782)
         );
  AOI21_X1 U5979 ( .B1(n6728), .B2(n5167), .A(n4782), .ZN(n4784) );
  NAND2_X1 U5980 ( .A1(n4794), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4783) );
  OAI211_X1 U5981 ( .C1(n6675), .C2(n6613), .A(n4784), .B(n4783), .ZN(U3082)
         );
  OAI22_X1 U5982 ( .A1(n4792), .A2(n6718), .B1(n4791), .B2(n6712), .ZN(n4785)
         );
  AOI21_X1 U5983 ( .B1(n6715), .B2(n5167), .A(n4785), .ZN(n4787) );
  NAND2_X1 U5984 ( .A1(n4794), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4786) );
  OAI211_X1 U5985 ( .C1(n6675), .C2(n6713), .A(n4787), .B(n4786), .ZN(U3080)
         );
  OAI22_X1 U5986 ( .A1(n4792), .A2(n6711), .B1(n4791), .B2(n5141), .ZN(n4788)
         );
  AOI21_X1 U5987 ( .B1(n6707), .B2(n5167), .A(n4788), .ZN(n4790) );
  NAND2_X1 U5988 ( .A1(n4794), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4789) );
  OAI211_X1 U5989 ( .C1(n6675), .C2(n6606), .A(n4790), .B(n4789), .ZN(U3079)
         );
  OAI22_X1 U5990 ( .A1(n4792), .A2(n6744), .B1(n4791), .B2(n6735), .ZN(n4793)
         );
  AOI21_X1 U5991 ( .B1(n6740), .B2(n5167), .A(n4793), .ZN(n4796) );
  NAND2_X1 U5992 ( .A1(n4794), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4795) );
  OAI211_X1 U5993 ( .C1(n6675), .C2(n6736), .A(n4796), .B(n4795), .ZN(U3083)
         );
  INV_X1 U5994 ( .A(DATAI_6_), .ZN(n5809) );
  INV_X1 U5995 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6380) );
  OAI222_X1 U5996 ( .A1(n4797), .A2(n6148), .B1(n6349), .B2(n5809), .C1(n6354), 
        .C2(n6380), .ZN(U2885) );
  XNOR2_X1 U5997 ( .A(n4798), .B(n4760), .ZN(n6429) );
  INV_X1 U5998 ( .A(n4799), .ZN(n4800) );
  XNOR2_X1 U5999 ( .A(n4801), .B(n4800), .ZN(n6488) );
  AOI22_X1 U6000 ( .A1(n6331), .A2(n6488), .B1(n5504), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4802) );
  OAI21_X1 U6001 ( .B1(n6429), .B2(n5521), .A(n4802), .ZN(U2852) );
  AOI21_X1 U6002 ( .B1(n4807), .B2(STATEBS16_REG_SCAN_IN), .A(n6678), .ZN(
        n6589) );
  NAND2_X1 U6003 ( .A1(n5094), .A2(n5087), .ZN(n6588) );
  NOR2_X1 U6004 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4853) );
  AND2_X1 U6005 ( .A1(n4853), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6587)
         );
  NAND2_X1 U6006 ( .A1(n6587), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4831) );
  INV_X1 U6007 ( .A(n4809), .ZN(n4805) );
  INV_X1 U6008 ( .A(n4807), .ZN(n4806) );
  OAI22_X1 U6009 ( .A1(n6634), .A2(n6665), .B1(n5145), .B2(n4831), .ZN(n4808)
         );
  AOI21_X1 U6010 ( .B1(n6730), .B2(n6616), .A(n4808), .ZN(n4812) );
  NAND2_X1 U6011 ( .A1(n6589), .A2(n4809), .ZN(n4810) );
  NAND2_X1 U6012 ( .A1(n4833), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4811) );
  OAI211_X1 U6013 ( .C1(n4836), .C2(n6733), .A(n4812), .B(n4811), .ZN(U3066)
         );
  OAI22_X1 U6014 ( .A1(n6634), .A2(n6661), .B1(n6719), .B2(n4831), .ZN(n4813)
         );
  AOI21_X1 U6015 ( .B1(n6658), .B2(n6616), .A(n4813), .ZN(n4815) );
  NAND2_X1 U6016 ( .A1(n4833), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4814) );
  OAI211_X1 U6017 ( .C1(n4836), .C2(n6725), .A(n4815), .B(n4814), .ZN(U3065)
         );
  OAI22_X1 U6018 ( .A1(n6634), .A2(n6655), .B1(n6712), .B2(n4831), .ZN(n4816)
         );
  AOI21_X1 U6019 ( .B1(n6652), .B2(n6616), .A(n4816), .ZN(n4818) );
  NAND2_X1 U6020 ( .A1(n4833), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4817) );
  OAI211_X1 U6021 ( .C1(n4836), .C2(n6718), .A(n4818), .B(n4817), .ZN(U3064)
         );
  OAI22_X1 U6022 ( .A1(n6634), .A2(n6649), .B1(n5141), .B2(n4831), .ZN(n4819)
         );
  AOI21_X1 U6023 ( .B1(n6708), .B2(n6616), .A(n4819), .ZN(n4821) );
  NAND2_X1 U6024 ( .A1(n4833), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4820) );
  OAI211_X1 U6025 ( .C1(n4836), .C2(n6711), .A(n4821), .B(n4820), .ZN(U3063)
         );
  OAI22_X1 U6026 ( .A1(n6634), .A2(n6645), .B1(n5137), .B2(n4831), .ZN(n4822)
         );
  AOI21_X1 U6027 ( .B1(n6702), .B2(n6616), .A(n4822), .ZN(n4824) );
  NAND2_X1 U6028 ( .A1(n4833), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4823) );
  OAI211_X1 U6029 ( .C1(n4836), .C2(n6705), .A(n4824), .B(n4823), .ZN(U3062)
         );
  OAI22_X1 U6030 ( .A1(n6634), .A2(n6637), .B1(n5158), .B2(n4831), .ZN(n4825)
         );
  AOI21_X1 U6031 ( .B1(n6690), .B2(n6616), .A(n4825), .ZN(n4827) );
  NAND2_X1 U6032 ( .A1(n4833), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4826) );
  OAI211_X1 U6033 ( .C1(n4836), .C2(n6693), .A(n4827), .B(n4826), .ZN(U3060)
         );
  OAI22_X1 U6034 ( .A1(n6634), .A2(n6641), .B1(n5164), .B2(n4831), .ZN(n4828)
         );
  AOI21_X1 U6035 ( .B1(n6696), .B2(n6616), .A(n4828), .ZN(n4830) );
  NAND2_X1 U6036 ( .A1(n4833), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4829) );
  OAI211_X1 U6037 ( .C1(n4836), .C2(n6699), .A(n4830), .B(n4829), .ZN(U3061)
         );
  OAI22_X1 U6038 ( .A1(n6634), .A2(n6676), .B1(n6735), .B2(n4831), .ZN(n4832)
         );
  AOI21_X1 U6039 ( .B1(n6671), .B2(n6616), .A(n4832), .ZN(n4835) );
  NAND2_X1 U6040 ( .A1(n4833), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4834) );
  OAI211_X1 U6041 ( .C1(n4836), .C2(n6744), .A(n4835), .B(n4834), .ZN(U3067)
         );
  INV_X1 U6042 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6378) );
  INV_X1 U6043 ( .A(DATAI_7_), .ZN(n4837) );
  OAI222_X1 U6044 ( .A1(n6148), .A2(n6429), .B1(n6354), .B2(n6378), .C1(n4837), 
        .C2(n6349), .ZN(U2884) );
  NAND2_X1 U6045 ( .A1(n4839), .A2(n4840), .ZN(n4841) );
  NAND2_X1 U6046 ( .A1(n4838), .A2(n4841), .ZN(n5885) );
  AOI22_X1 U6047 ( .A1(n6350), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6345), .ZN(n4842) );
  OAI21_X1 U6048 ( .B1(n5885), .B2(n6148), .A(n4842), .ZN(U2883) );
  OR2_X1 U6049 ( .A1(n4844), .A2(n4843), .ZN(n4846) );
  NAND2_X1 U6050 ( .A1(n4846), .A2(n4845), .ZN(n5411) );
  INV_X1 U6051 ( .A(n5411), .ZN(n6478) );
  AOI22_X1 U6052 ( .A1(n6331), .A2(n6478), .B1(n5504), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4847) );
  OAI21_X1 U6053 ( .B1(n5885), .B2(n5521), .A(n4847), .ZN(U2851) );
  OR2_X1 U6054 ( .A1(n2977), .A2(n5127), .ZN(n4867) );
  INV_X1 U6055 ( .A(n4867), .ZN(n4851) );
  INV_X1 U6056 ( .A(n4871), .ZN(n4850) );
  AOI211_X1 U6057 ( .C1(n4938), .C2(n4982), .A(n4851), .B(n4876), .ZN(n4857)
         );
  NAND2_X1 U6058 ( .A1(n4853), .A2(n4852), .ZN(n4873) );
  NOR2_X1 U6059 ( .A1(n4873), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4903)
         );
  INV_X1 U6060 ( .A(n5051), .ZN(n6621) );
  NAND2_X1 U6061 ( .A1(n6621), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4854) );
  NAND2_X1 U6062 ( .A1(n4855), .A2(n4854), .ZN(n5090) );
  AOI21_X1 U6063 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6585), .A(n5090), .ZN(
        n6593) );
  OAI211_X1 U6064 ( .C1(n4903), .C2(n6769), .A(n6593), .B(n5131), .ZN(n4856)
         );
  INV_X1 U6065 ( .A(n4938), .ZN(n4862) );
  NOR2_X1 U6066 ( .A1(n6592), .A2(n6621), .ZN(n5134) );
  INV_X1 U6067 ( .A(n6585), .ZN(n4859) );
  NAND2_X1 U6068 ( .A1(n5134), .A2(n4859), .ZN(n4860) );
  OAI21_X1 U6069 ( .B1(n6625), .B2(n5127), .A(n4860), .ZN(n4934) );
  AOI22_X1 U6070 ( .A1(n4934), .A2(n6628), .B1(n6683), .B2(n4903), .ZN(n4861)
         );
  OAI21_X1 U6071 ( .B1(n4862), .B2(n6597), .A(n4861), .ZN(n4863) );
  AOI21_X1 U6072 ( .B1(n4939), .B2(n6684), .A(n4863), .ZN(n4864) );
  OAI21_X1 U6073 ( .B1(n4943), .B2(n4865), .A(n4864), .ZN(U3020) );
  INV_X1 U6074 ( .A(n4876), .ZN(n4869) );
  OR2_X1 U6075 ( .A1(n4873), .A2(n6626), .ZN(n4897) );
  OAI21_X1 U6076 ( .B1(n4867), .B2(n4866), .A(n4897), .ZN(n4875) );
  INV_X1 U6077 ( .A(n4873), .ZN(n4868) );
  OAI22_X1 U6078 ( .A1(n5016), .A2(n6641), .B1(n5164), .B2(n4897), .ZN(n4872)
         );
  AOI21_X1 U6079 ( .B1(n6696), .B2(n4939), .A(n4872), .ZN(n4878) );
  AOI21_X1 U6080 ( .B1(n6678), .B2(n4873), .A(n6558), .ZN(n4874) );
  NAND2_X1 U6081 ( .A1(n4899), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4877) );
  OAI211_X1 U6082 ( .C1(n4902), .C2(n6699), .A(n4878), .B(n4877), .ZN(U3029)
         );
  OAI22_X1 U6083 ( .A1(n5016), .A2(n6637), .B1(n5158), .B2(n4897), .ZN(n4879)
         );
  AOI21_X1 U6084 ( .B1(n6690), .B2(n4939), .A(n4879), .ZN(n4881) );
  NAND2_X1 U6085 ( .A1(n4899), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4880) );
  OAI211_X1 U6086 ( .C1(n4902), .C2(n6693), .A(n4881), .B(n4880), .ZN(U3028)
         );
  OAI22_X1 U6087 ( .A1(n5016), .A2(n6665), .B1(n5145), .B2(n4897), .ZN(n4882)
         );
  AOI21_X1 U6088 ( .B1(n6730), .B2(n4939), .A(n4882), .ZN(n4884) );
  NAND2_X1 U6089 ( .A1(n4899), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4883) );
  OAI211_X1 U6090 ( .C1(n4902), .C2(n6733), .A(n4884), .B(n4883), .ZN(U3034)
         );
  OAI22_X1 U6091 ( .A1(n5016), .A2(n6645), .B1(n5137), .B2(n4897), .ZN(n4885)
         );
  AOI21_X1 U6092 ( .B1(n6702), .B2(n4939), .A(n4885), .ZN(n4887) );
  NAND2_X1 U6093 ( .A1(n4899), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4886) );
  OAI211_X1 U6094 ( .C1(n4902), .C2(n6705), .A(n4887), .B(n4886), .ZN(U3030)
         );
  OAI22_X1 U6095 ( .A1(n5016), .A2(n6661), .B1(n6719), .B2(n4897), .ZN(n4888)
         );
  AOI21_X1 U6096 ( .B1(n6658), .B2(n4939), .A(n4888), .ZN(n4890) );
  NAND2_X1 U6097 ( .A1(n4899), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4889) );
  OAI211_X1 U6098 ( .C1(n4902), .C2(n6725), .A(n4890), .B(n4889), .ZN(U3033)
         );
  OAI22_X1 U6099 ( .A1(n5016), .A2(n6655), .B1(n6712), .B2(n4897), .ZN(n4891)
         );
  AOI21_X1 U6100 ( .B1(n6652), .B2(n4939), .A(n4891), .ZN(n4893) );
  NAND2_X1 U6101 ( .A1(n4899), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4892) );
  OAI211_X1 U6102 ( .C1(n4902), .C2(n6718), .A(n4893), .B(n4892), .ZN(U3032)
         );
  OAI22_X1 U6103 ( .A1(n5016), .A2(n6649), .B1(n5141), .B2(n4897), .ZN(n4894)
         );
  AOI21_X1 U6104 ( .B1(n6708), .B2(n4939), .A(n4894), .ZN(n4896) );
  NAND2_X1 U6105 ( .A1(n4899), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4895) );
  OAI211_X1 U6106 ( .C1(n4902), .C2(n6711), .A(n4896), .B(n4895), .ZN(U3031)
         );
  OAI22_X1 U6107 ( .A1(n5016), .A2(n6676), .B1(n6735), .B2(n4897), .ZN(n4898)
         );
  AOI21_X1 U6108 ( .B1(n6671), .B2(n4939), .A(n4898), .ZN(n4901) );
  NAND2_X1 U6109 ( .A1(n4899), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4900) );
  OAI211_X1 U6110 ( .C1(n4902), .C2(n6744), .A(n4901), .B(n4900), .ZN(U3035)
         );
  INV_X1 U6111 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4908) );
  INV_X1 U6112 ( .A(n4903), .ZN(n4936) );
  NAND2_X1 U6113 ( .A1(n4934), .A2(n6651), .ZN(n4904) );
  OAI21_X1 U6114 ( .B1(n4936), .B2(n6712), .A(n4904), .ZN(n4905) );
  AOI21_X1 U6115 ( .B1(n4938), .B2(n6652), .A(n4905), .ZN(n4907) );
  NAND2_X1 U6116 ( .A1(n4939), .A2(n6715), .ZN(n4906) );
  OAI211_X1 U6117 ( .C1(n4943), .C2(n4908), .A(n4907), .B(n4906), .ZN(U3024)
         );
  INV_X1 U6118 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4913) );
  NAND2_X1 U6119 ( .A1(n4934), .A2(n6657), .ZN(n4909) );
  OAI21_X1 U6120 ( .B1(n4936), .B2(n6719), .A(n4909), .ZN(n4910) );
  AOI21_X1 U6121 ( .B1(n4938), .B2(n6658), .A(n4910), .ZN(n4912) );
  NAND2_X1 U6122 ( .A1(n4939), .A2(n6722), .ZN(n4911) );
  OAI211_X1 U6123 ( .C1(n4943), .C2(n4913), .A(n4912), .B(n4911), .ZN(U3025)
         );
  NAND2_X1 U6124 ( .A1(n4934), .A2(n6638), .ZN(n4914) );
  OAI21_X1 U6125 ( .B1(n4936), .B2(n5164), .A(n4914), .ZN(n4915) );
  AOI21_X1 U6126 ( .B1(n4938), .B2(n6696), .A(n4915), .ZN(n4917) );
  NAND2_X1 U6127 ( .A1(n4939), .A2(n6695), .ZN(n4916) );
  OAI211_X1 U6128 ( .C1(n4943), .C2(n4918), .A(n4917), .B(n4916), .ZN(U3021)
         );
  INV_X1 U6129 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U6130 ( .A1(n4934), .A2(n6662), .ZN(n4919) );
  OAI21_X1 U6131 ( .B1(n4936), .B2(n5145), .A(n4919), .ZN(n4920) );
  AOI21_X1 U6132 ( .B1(n4938), .B2(n6730), .A(n4920), .ZN(n4922) );
  NAND2_X1 U6133 ( .A1(n4939), .A2(n6728), .ZN(n4921) );
  OAI211_X1 U6134 ( .C1(n4943), .C2(n4923), .A(n4922), .B(n4921), .ZN(U3026)
         );
  INV_X1 U6135 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4928) );
  NAND2_X1 U6136 ( .A1(n4934), .A2(n6642), .ZN(n4924) );
  OAI21_X1 U6137 ( .B1(n4936), .B2(n5137), .A(n4924), .ZN(n4925) );
  AOI21_X1 U6138 ( .B1(n4938), .B2(n6702), .A(n4925), .ZN(n4927) );
  NAND2_X1 U6139 ( .A1(n4939), .A2(n6701), .ZN(n4926) );
  OAI211_X1 U6140 ( .C1(n4943), .C2(n4928), .A(n4927), .B(n4926), .ZN(U3022)
         );
  NAND2_X1 U6141 ( .A1(n4934), .A2(n6668), .ZN(n4929) );
  OAI21_X1 U6142 ( .B1(n4936), .B2(n6735), .A(n4929), .ZN(n4930) );
  AOI21_X1 U6143 ( .B1(n4938), .B2(n6671), .A(n4930), .ZN(n4932) );
  NAND2_X1 U6144 ( .A1(n4939), .A2(n6740), .ZN(n4931) );
  OAI211_X1 U6145 ( .C1(n4943), .C2(n4933), .A(n4932), .B(n4931), .ZN(U3027)
         );
  INV_X1 U6146 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4942) );
  NAND2_X1 U6147 ( .A1(n4934), .A2(n6646), .ZN(n4935) );
  OAI21_X1 U6148 ( .B1(n4936), .B2(n5141), .A(n4935), .ZN(n4937) );
  AOI21_X1 U6149 ( .B1(n4938), .B2(n6708), .A(n4937), .ZN(n4941) );
  NAND2_X1 U6150 ( .A1(n4939), .A2(n6707), .ZN(n4940) );
  OAI211_X1 U6151 ( .C1(n4943), .C2(n4942), .A(n4941), .B(n4940), .ZN(U3023)
         );
  INV_X1 U6152 ( .A(n4944), .ZN(n4945) );
  AOI211_X1 U6153 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n4950), .A(n6626), .B(n4945), .ZN(n4955) );
  NAND2_X1 U6154 ( .A1(n4955), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4957) );
  NAND2_X1 U6155 ( .A1(n5452), .A2(n4946), .ZN(n4952) );
  NOR2_X1 U6156 ( .A1(n4480), .A2(n4449), .ZN(n4949) );
  AOI22_X1 U6157 ( .A1(n4950), .A2(n5194), .B1(n4949), .B2(n4948), .ZN(n4951)
         );
  NAND2_X1 U6158 ( .A1(n4952), .A2(n4951), .ZN(n5192) );
  INV_X1 U6159 ( .A(n5192), .ZN(n4953) );
  OAI22_X1 U6160 ( .A1(n4955), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n4954), .B2(n4953), .ZN(n4956) );
  NAND2_X1 U6161 ( .A1(n4957), .A2(n4956), .ZN(n4958) );
  AOI222_X1 U6162 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n4959), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n4958), .C1(n4959), .C2(n4958), 
        .ZN(n4960) );
  AOI222_X1 U6163 ( .A1(n4961), .A2(n6780), .B1(n4961), .B2(n4960), .C1(n6780), 
        .C2(n4960), .ZN(n4970) );
  OAI21_X1 U6164 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n4962), 
        .ZN(n4963) );
  NAND4_X1 U6165 ( .A1(n4966), .A2(n4965), .A3(n4964), .A4(n4963), .ZN(n4967)
         );
  NOR2_X1 U6166 ( .A1(n4968), .A2(n4967), .ZN(n4969) );
  OAI21_X1 U6167 ( .B1(n4970), .B2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n4969), 
        .ZN(n4971) );
  INV_X1 U6168 ( .A(n4971), .ZN(n4981) );
  OAI22_X1 U6169 ( .A1(n4971), .A2(n6155), .B1(n6791), .B2(n4179), .ZN(n4972)
         );
  OAI21_X1 U6170 ( .B1(n4974), .B2(n4973), .A(n4972), .ZN(n6770) );
  OAI21_X1 U6171 ( .B1(n4975), .B2(n6132), .A(n6770), .ZN(n4978) );
  OAI21_X1 U6172 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4179), .A(n6770), .ZN(
        n6746) );
  NOR2_X1 U6173 ( .A1(n6746), .A2(n4976), .ZN(n4977) );
  MUX2_X1 U6174 ( .A(n4978), .B(n4977), .S(STATE2_REG_0__SCAN_IN), .Z(n4980)
         );
  OAI211_X1 U6175 ( .C1(n4981), .C2(n6155), .A(n4980), .B(n4979), .ZN(U3148)
         );
  OAI21_X1 U6176 ( .B1(n4983), .B2(n6578), .A(n4982), .ZN(n4984) );
  NAND2_X1 U6177 ( .A1(n4461), .A2(n5452), .ZN(n5049) );
  OR2_X1 U6178 ( .A1(n2977), .A2(n5049), .ZN(n4986) );
  AOI21_X1 U6179 ( .B1(n4984), .B2(n4986), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4985) );
  NAND2_X1 U6180 ( .A1(n6554), .A2(n6780), .ZN(n6559) );
  NOR2_X1 U6181 ( .A1(n6559), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4988)
         );
  NAND2_X1 U6182 ( .A1(n5010), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4991) );
  INV_X1 U6183 ( .A(n4986), .ZN(n6553) );
  NOR3_X1 U6184 ( .A1(n6592), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5051), 
        .ZN(n4987) );
  AOI21_X1 U6185 ( .B1(n6553), .B2(n6774), .A(n4987), .ZN(n5012) );
  INV_X1 U6186 ( .A(n4988), .ZN(n5011) );
  OAI22_X1 U6187 ( .A1(n5012), .A2(n6744), .B1(n5011), .B2(n6735), .ZN(n4989)
         );
  AOI21_X1 U6188 ( .B1(n6578), .B2(n6740), .A(n4989), .ZN(n4990) );
  OAI211_X1 U6189 ( .C1(n5016), .C2(n6736), .A(n4991), .B(n4990), .ZN(U3043)
         );
  NAND2_X1 U6190 ( .A1(n5010), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4994) );
  OAI22_X1 U6191 ( .A1(n5012), .A2(n6693), .B1(n5011), .B2(n5158), .ZN(n4992)
         );
  AOI21_X1 U6192 ( .B1(n6578), .B2(n6684), .A(n4992), .ZN(n4993) );
  OAI211_X1 U6193 ( .C1(n5016), .C2(n6597), .A(n4994), .B(n4993), .ZN(U3036)
         );
  NAND2_X1 U6194 ( .A1(n5010), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4997) );
  OAI22_X1 U6195 ( .A1(n5012), .A2(n6705), .B1(n5011), .B2(n5137), .ZN(n4995)
         );
  AOI21_X1 U6196 ( .B1(n6578), .B2(n6701), .A(n4995), .ZN(n4996) );
  OAI211_X1 U6197 ( .C1(n5016), .C2(n6603), .A(n4997), .B(n4996), .ZN(U3038)
         );
  NAND2_X1 U6198 ( .A1(n5010), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5000) );
  OAI22_X1 U6199 ( .A1(n5012), .A2(n6718), .B1(n5011), .B2(n6712), .ZN(n4998)
         );
  AOI21_X1 U6200 ( .B1(n6578), .B2(n6715), .A(n4998), .ZN(n4999) );
  OAI211_X1 U6201 ( .C1(n5016), .C2(n6713), .A(n5000), .B(n4999), .ZN(U3040)
         );
  NAND2_X1 U6202 ( .A1(n5010), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5003) );
  OAI22_X1 U6203 ( .A1(n5012), .A2(n6733), .B1(n5011), .B2(n5145), .ZN(n5001)
         );
  AOI21_X1 U6204 ( .B1(n6578), .B2(n6728), .A(n5001), .ZN(n5002) );
  OAI211_X1 U6205 ( .C1(n5016), .C2(n6613), .A(n5003), .B(n5002), .ZN(U3042)
         );
  NAND2_X1 U6206 ( .A1(n5010), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5006) );
  OAI22_X1 U6207 ( .A1(n5012), .A2(n6711), .B1(n5011), .B2(n5141), .ZN(n5004)
         );
  AOI21_X1 U6208 ( .B1(n6578), .B2(n6707), .A(n5004), .ZN(n5005) );
  OAI211_X1 U6209 ( .C1(n5016), .C2(n6606), .A(n5006), .B(n5005), .ZN(U3039)
         );
  NAND2_X1 U6210 ( .A1(n5010), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5009) );
  OAI22_X1 U6211 ( .A1(n5012), .A2(n6725), .B1(n5011), .B2(n6719), .ZN(n5007)
         );
  AOI21_X1 U6212 ( .B1(n6578), .B2(n6722), .A(n5007), .ZN(n5008) );
  OAI211_X1 U6213 ( .C1(n5016), .C2(n6720), .A(n5009), .B(n5008), .ZN(U3041)
         );
  NAND2_X1 U6214 ( .A1(n5010), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5015) );
  OAI22_X1 U6215 ( .A1(n5012), .A2(n6699), .B1(n5011), .B2(n5164), .ZN(n5013)
         );
  AOI21_X1 U6216 ( .B1(n6578), .B2(n6695), .A(n5013), .ZN(n5014) );
  OAI211_X1 U6217 ( .C1(n5016), .C2(n6600), .A(n5015), .B(n5014), .ZN(U3037)
         );
  NAND2_X1 U6218 ( .A1(n5017), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5018)
         );
  NAND2_X1 U6219 ( .A1(n5020), .A2(n3920), .ZN(n5026) );
  INV_X1 U6220 ( .A(n5021), .ZN(n5022) );
  OR2_X1 U6221 ( .A1(n5023), .A2(n5022), .ZN(n5031) );
  XNOR2_X1 U6222 ( .A(n5031), .B(n5032), .ZN(n5024) );
  NAND2_X1 U6223 ( .A1(n5024), .A2(n5216), .ZN(n5025) );
  NAND2_X1 U6224 ( .A1(n5026), .A2(n5025), .ZN(n5027) );
  INV_X1 U6225 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U6226 ( .A1(n5027), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5028)
         );
  NAND3_X1 U6227 ( .A1(n5029), .A2(n5030), .A3(n3920), .ZN(n5036) );
  INV_X1 U6228 ( .A(n5031), .ZN(n5033) );
  NAND2_X1 U6229 ( .A1(n5033), .A2(n5032), .ZN(n5202) );
  XNOR2_X1 U6230 ( .A(n5202), .B(n5203), .ZN(n5034) );
  NAND2_X1 U6231 ( .A1(n5034), .A2(n5216), .ZN(n5035) );
  NAND2_X1 U6232 ( .A1(n5036), .A2(n5035), .ZN(n5208) );
  XOR2_X1 U6233 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .B(n5208), .Z(n5037) );
  NAND2_X1 U6234 ( .A1(n5212), .A2(n5037), .ZN(n6427) );
  OAI21_X1 U6235 ( .B1(n5212), .B2(n5037), .A(n6427), .ZN(n6500) );
  INV_X1 U6236 ( .A(n5038), .ZN(n5428) );
  NAND2_X1 U6237 ( .A1(n6450), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5039)
         );
  NAND2_X1 U6238 ( .A1(n6490), .A2(REIP_REG_6__SCAN_IN), .ZN(n6497) );
  OAI211_X1 U6239 ( .C1(n6461), .C2(n5428), .A(n5039), .B(n6497), .ZN(n5040)
         );
  AOI21_X1 U6240 ( .B1(n5426), .B2(n6456), .A(n5040), .ZN(n5041) );
  OAI21_X1 U6241 ( .B1(n6500), .B2(n6161), .A(n5041), .ZN(U2980) );
  NAND2_X1 U6242 ( .A1(n4838), .A2(n5043), .ZN(n5044) );
  NAND2_X1 U6243 ( .A1(n5042), .A2(n5044), .ZN(n5873) );
  AOI21_X1 U6244 ( .B1(n5045), .B2(n4845), .A(n5174), .ZN(n6472) );
  AOI22_X1 U6245 ( .A1(n6331), .A2(n6472), .B1(EBX_REG_9__SCAN_IN), .B2(n5504), 
        .ZN(n5046) );
  OAI21_X1 U6246 ( .B1(n5873), .B2(n5521), .A(n5046), .ZN(U2850) );
  NOR2_X1 U6247 ( .A1(n6729), .A2(n6678), .ZN(n5048) );
  AOI21_X1 U6248 ( .B1(n5048), .B2(n5058), .A(n6776), .ZN(n5057) );
  INV_X1 U6249 ( .A(n5057), .ZN(n5053) );
  INV_X1 U6250 ( .A(n5049), .ZN(n5050) );
  NOR3_X1 U6251 ( .A1(n6592), .A2(n5051), .A3(n6780), .ZN(n5052) );
  AND2_X1 U6252 ( .A1(n6554), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6689)
         );
  NAND2_X1 U6253 ( .A1(n6689), .A2(n6626), .ZN(n5081) );
  INV_X1 U6254 ( .A(n5131), .ZN(n6622) );
  AOI211_X1 U6255 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5081), .A(n5054), .B(
        n6622), .ZN(n5055) );
  NAND2_X1 U6256 ( .A1(n5080), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5061)
         );
  OAI22_X1 U6257 ( .A1(n6737), .A2(n6649), .B1(n5141), .B2(n5081), .ZN(n5059)
         );
  AOI21_X1 U6258 ( .B1(n5083), .B2(n6708), .A(n5059), .ZN(n5060) );
  OAI211_X1 U6259 ( .C1(n5086), .C2(n6711), .A(n5061), .B(n5060), .ZN(U3103)
         );
  NAND2_X1 U6260 ( .A1(n5080), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5064)
         );
  OAI22_X1 U6261 ( .A1(n6737), .A2(n6641), .B1(n5164), .B2(n5081), .ZN(n5062)
         );
  AOI21_X1 U6262 ( .B1(n5083), .B2(n6696), .A(n5062), .ZN(n5063) );
  OAI211_X1 U6263 ( .C1(n5086), .C2(n6699), .A(n5064), .B(n5063), .ZN(U3101)
         );
  NAND2_X1 U6264 ( .A1(n5080), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5067)
         );
  OAI22_X1 U6265 ( .A1(n6737), .A2(n6637), .B1(n5158), .B2(n5081), .ZN(n5065)
         );
  AOI21_X1 U6266 ( .B1(n5083), .B2(n6690), .A(n5065), .ZN(n5066) );
  OAI211_X1 U6267 ( .C1(n5086), .C2(n6693), .A(n5067), .B(n5066), .ZN(U3100)
         );
  NAND2_X1 U6268 ( .A1(n5080), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5070)
         );
  OAI22_X1 U6269 ( .A1(n6737), .A2(n6655), .B1(n6712), .B2(n5081), .ZN(n5068)
         );
  AOI21_X1 U6270 ( .B1(n5083), .B2(n6652), .A(n5068), .ZN(n5069) );
  OAI211_X1 U6271 ( .C1(n5086), .C2(n6718), .A(n5070), .B(n5069), .ZN(U3104)
         );
  NAND2_X1 U6272 ( .A1(n5080), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5073)
         );
  OAI22_X1 U6273 ( .A1(n6737), .A2(n6676), .B1(n6735), .B2(n5081), .ZN(n5071)
         );
  AOI21_X1 U6274 ( .B1(n5083), .B2(n6671), .A(n5071), .ZN(n5072) );
  OAI211_X1 U6275 ( .C1(n5086), .C2(n6744), .A(n5073), .B(n5072), .ZN(U3107)
         );
  NAND2_X1 U6276 ( .A1(n5080), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5076)
         );
  OAI22_X1 U6277 ( .A1(n6737), .A2(n6645), .B1(n5137), .B2(n5081), .ZN(n5074)
         );
  AOI21_X1 U6278 ( .B1(n5083), .B2(n6702), .A(n5074), .ZN(n5075) );
  OAI211_X1 U6279 ( .C1(n5086), .C2(n6705), .A(n5076), .B(n5075), .ZN(U3102)
         );
  NAND2_X1 U6280 ( .A1(n5080), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5079)
         );
  OAI22_X1 U6281 ( .A1(n6737), .A2(n6661), .B1(n6719), .B2(n5081), .ZN(n5077)
         );
  AOI21_X1 U6282 ( .B1(n5083), .B2(n6658), .A(n5077), .ZN(n5078) );
  OAI211_X1 U6283 ( .C1(n5086), .C2(n6725), .A(n5079), .B(n5078), .ZN(U3105)
         );
  NAND2_X1 U6284 ( .A1(n5080), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5085)
         );
  OAI22_X1 U6285 ( .A1(n6737), .A2(n6665), .B1(n5145), .B2(n5081), .ZN(n5082)
         );
  AOI21_X1 U6286 ( .B1(n5083), .B2(n6730), .A(n5082), .ZN(n5084) );
  OAI211_X1 U6287 ( .C1(n5086), .C2(n6733), .A(n5085), .B(n5084), .ZN(U3106)
         );
  NOR3_X1 U6288 ( .A1(n5120), .A2(n6739), .A3(n6678), .ZN(n5088) );
  OAI22_X1 U6289 ( .A1(n5088), .A2(n6776), .B1(n5087), .B2(n6586), .ZN(n5093)
         );
  NOR2_X1 U6290 ( .A1(n6585), .A2(n4686), .ZN(n5089) );
  NOR2_X1 U6291 ( .A1(n5090), .A2(n5089), .ZN(n5132) );
  NAND2_X1 U6292 ( .A1(n5091), .A2(n6626), .ZN(n5117) );
  NAND2_X1 U6293 ( .A1(n5117), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5092) );
  NAND4_X1 U6294 ( .A1(n5093), .A2(n5132), .A3(n6592), .A4(n5092), .ZN(n5116)
         );
  NAND2_X1 U6295 ( .A1(n5116), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5097)
         );
  NOR2_X1 U6296 ( .A1(n5131), .A2(n6621), .ZN(n6583) );
  AOI22_X1 U6297 ( .A1(n5136), .A2(n5094), .B1(n6585), .B2(n6583), .ZN(n5118)
         );
  OAI22_X1 U6298 ( .A1(n5118), .A2(n6693), .B1(n5158), .B2(n5117), .ZN(n5095)
         );
  AOI21_X1 U6299 ( .B1(n5120), .B2(n6684), .A(n5095), .ZN(n5096) );
  OAI211_X1 U6300 ( .C1(n5123), .C2(n6597), .A(n5097), .B(n5096), .ZN(U3116)
         );
  NAND2_X1 U6301 ( .A1(n5116), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5100)
         );
  OAI22_X1 U6302 ( .A1(n5118), .A2(n6733), .B1(n5145), .B2(n5117), .ZN(n5098)
         );
  AOI21_X1 U6303 ( .B1(n5120), .B2(n6728), .A(n5098), .ZN(n5099) );
  OAI211_X1 U6304 ( .C1(n5123), .C2(n6613), .A(n5100), .B(n5099), .ZN(U3122)
         );
  NAND2_X1 U6305 ( .A1(n5116), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5103)
         );
  OAI22_X1 U6306 ( .A1(n5118), .A2(n6725), .B1(n6719), .B2(n5117), .ZN(n5101)
         );
  AOI21_X1 U6307 ( .B1(n5120), .B2(n6722), .A(n5101), .ZN(n5102) );
  OAI211_X1 U6308 ( .C1(n5123), .C2(n6720), .A(n5103), .B(n5102), .ZN(U3121)
         );
  NAND2_X1 U6309 ( .A1(n5116), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5106)
         );
  OAI22_X1 U6310 ( .A1(n5118), .A2(n6718), .B1(n6712), .B2(n5117), .ZN(n5104)
         );
  AOI21_X1 U6311 ( .B1(n5120), .B2(n6715), .A(n5104), .ZN(n5105) );
  OAI211_X1 U6312 ( .C1(n5123), .C2(n6713), .A(n5106), .B(n5105), .ZN(U3120)
         );
  NAND2_X1 U6313 ( .A1(n5116), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5109)
         );
  OAI22_X1 U6314 ( .A1(n5118), .A2(n6711), .B1(n5141), .B2(n5117), .ZN(n5107)
         );
  AOI21_X1 U6315 ( .B1(n5120), .B2(n6707), .A(n5107), .ZN(n5108) );
  OAI211_X1 U6316 ( .C1(n5123), .C2(n6606), .A(n5109), .B(n5108), .ZN(U3119)
         );
  NAND2_X1 U6317 ( .A1(n5116), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5112)
         );
  OAI22_X1 U6318 ( .A1(n5118), .A2(n6705), .B1(n5137), .B2(n5117), .ZN(n5110)
         );
  AOI21_X1 U6319 ( .B1(n5120), .B2(n6701), .A(n5110), .ZN(n5111) );
  OAI211_X1 U6320 ( .C1(n5123), .C2(n6603), .A(n5112), .B(n5111), .ZN(U3118)
         );
  NAND2_X1 U6321 ( .A1(n5116), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5115)
         );
  OAI22_X1 U6322 ( .A1(n5118), .A2(n6699), .B1(n5164), .B2(n5117), .ZN(n5113)
         );
  AOI21_X1 U6323 ( .B1(n5120), .B2(n6695), .A(n5113), .ZN(n5114) );
  OAI211_X1 U6324 ( .C1(n5123), .C2(n6600), .A(n5115), .B(n5114), .ZN(U3117)
         );
  NAND2_X1 U6325 ( .A1(n5116), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5122)
         );
  OAI22_X1 U6326 ( .A1(n5118), .A2(n6744), .B1(n6735), .B2(n5117), .ZN(n5119)
         );
  AOI21_X1 U6327 ( .B1(n5120), .B2(n6740), .A(n5119), .ZN(n5121) );
  OAI211_X1 U6328 ( .C1(n5123), .C2(n6736), .A(n5122), .B(n5121), .ZN(U3123)
         );
  INV_X1 U6329 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6374) );
  OAI222_X1 U6330 ( .A1(n5873), .A2(n6148), .B1(n6349), .B2(n5124), .C1(n6354), 
        .C2(n6374), .ZN(U2882) );
  OAI21_X1 U6331 ( .B1(n5125), .B2(n5167), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5126) );
  OAI211_X1 U6332 ( .C1(n5128), .C2(n5127), .A(n5126), .B(n6774), .ZN(n5133)
         );
  NAND2_X1 U6333 ( .A1(n5129), .A2(n6626), .ZN(n5163) );
  NAND2_X1 U6334 ( .A1(n5163), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5130) );
  NAND4_X1 U6335 ( .A1(n5133), .A2(n5132), .A3(n5131), .A4(n5130), .ZN(n5162)
         );
  NAND2_X1 U6336 ( .A1(n5162), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5140) );
  AOI22_X1 U6337 ( .A1(n5136), .A2(n5135), .B1(n6585), .B2(n5134), .ZN(n5165)
         );
  OAI22_X1 U6338 ( .A1(n5165), .A2(n6705), .B1(n5137), .B2(n5163), .ZN(n5138)
         );
  AOI21_X1 U6339 ( .B1(n6702), .B2(n5167), .A(n5138), .ZN(n5139) );
  OAI211_X1 U6340 ( .C1(n5170), .C2(n6645), .A(n5140), .B(n5139), .ZN(U3086)
         );
  NAND2_X1 U6341 ( .A1(n5162), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5144) );
  OAI22_X1 U6342 ( .A1(n5165), .A2(n6711), .B1(n5141), .B2(n5163), .ZN(n5142)
         );
  AOI21_X1 U6343 ( .B1(n6708), .B2(n5167), .A(n5142), .ZN(n5143) );
  OAI211_X1 U6344 ( .C1(n5170), .C2(n6649), .A(n5144), .B(n5143), .ZN(U3087)
         );
  NAND2_X1 U6345 ( .A1(n5162), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5148) );
  OAI22_X1 U6346 ( .A1(n5165), .A2(n6733), .B1(n5145), .B2(n5163), .ZN(n5146)
         );
  AOI21_X1 U6347 ( .B1(n6730), .B2(n5167), .A(n5146), .ZN(n5147) );
  OAI211_X1 U6348 ( .C1(n5170), .C2(n6665), .A(n5148), .B(n5147), .ZN(U3090)
         );
  NAND2_X1 U6349 ( .A1(n5162), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5151) );
  OAI22_X1 U6350 ( .A1(n5165), .A2(n6744), .B1(n6735), .B2(n5163), .ZN(n5149)
         );
  AOI21_X1 U6351 ( .B1(n6671), .B2(n5167), .A(n5149), .ZN(n5150) );
  OAI211_X1 U6352 ( .C1(n5170), .C2(n6676), .A(n5151), .B(n5150), .ZN(U3091)
         );
  NAND2_X1 U6353 ( .A1(n5162), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5154) );
  OAI22_X1 U6354 ( .A1(n5165), .A2(n6725), .B1(n6719), .B2(n5163), .ZN(n5152)
         );
  AOI21_X1 U6355 ( .B1(n6658), .B2(n5167), .A(n5152), .ZN(n5153) );
  OAI211_X1 U6356 ( .C1(n5170), .C2(n6661), .A(n5154), .B(n5153), .ZN(U3089)
         );
  NAND2_X1 U6357 ( .A1(n5162), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5157) );
  OAI22_X1 U6358 ( .A1(n5165), .A2(n6718), .B1(n6712), .B2(n5163), .ZN(n5155)
         );
  AOI21_X1 U6359 ( .B1(n6652), .B2(n5167), .A(n5155), .ZN(n5156) );
  OAI211_X1 U6360 ( .C1(n5170), .C2(n6655), .A(n5157), .B(n5156), .ZN(U3088)
         );
  NAND2_X1 U6361 ( .A1(n5162), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5161) );
  OAI22_X1 U6362 ( .A1(n5165), .A2(n6693), .B1(n5158), .B2(n5163), .ZN(n5159)
         );
  AOI21_X1 U6363 ( .B1(n6690), .B2(n5167), .A(n5159), .ZN(n5160) );
  OAI211_X1 U6364 ( .C1(n5170), .C2(n6637), .A(n5161), .B(n5160), .ZN(U3084)
         );
  NAND2_X1 U6365 ( .A1(n5162), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5169) );
  OAI22_X1 U6366 ( .A1(n5165), .A2(n6699), .B1(n5164), .B2(n5163), .ZN(n5166)
         );
  AOI21_X1 U6367 ( .B1(n6696), .B2(n5167), .A(n5166), .ZN(n5168) );
  OAI211_X1 U6368 ( .C1(n5170), .C2(n6641), .A(n5169), .B(n5168), .ZN(U3085)
         );
  AOI21_X1 U6369 ( .B1(n5173), .B2(n5042), .A(n5172), .ZN(n6265) );
  INV_X1 U6370 ( .A(n6265), .ZN(n5179) );
  OAI21_X1 U6371 ( .B1(n5175), .B2(n5174), .A(n5185), .ZN(n6261) );
  INV_X1 U6372 ( .A(n6261), .ZN(n5176) );
  AOI22_X1 U6373 ( .A1(n6331), .A2(n5176), .B1(EBX_REG_10__SCAN_IN), .B2(n5504), .ZN(n5177) );
  OAI21_X1 U6374 ( .B1(n5179), .B2(n5521), .A(n5177), .ZN(U2849) );
  INV_X1 U6375 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6372) );
  OAI222_X1 U6376 ( .A1(n5179), .A2(n6148), .B1(n6349), .B2(n5178), .C1(n6354), 
        .C2(n6372), .ZN(U2881) );
  OR2_X1 U6377 ( .A1(n5172), .A2(n5181), .ZN(n5182) );
  NAND2_X1 U6378 ( .A1(n5180), .A2(n5182), .ZN(n6251) );
  AOI22_X1 U6379 ( .A1(n6350), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6345), .ZN(n5183) );
  OAI21_X1 U6380 ( .B1(n6251), .B2(n6148), .A(n5183), .ZN(U2880) );
  AOI21_X1 U6381 ( .B1(n5186), .B2(n5185), .A(n5184), .ZN(n6463) );
  AOI22_X1 U6382 ( .A1(n6331), .A2(n6463), .B1(EBX_REG_11__SCAN_IN), .B2(n5504), .ZN(n5187) );
  OAI21_X1 U6383 ( .B1(n6251), .B2(n5521), .A(n5187), .ZN(U2848) );
  INV_X1 U6384 ( .A(n5188), .ZN(n5195) );
  INV_X1 U6385 ( .A(n6135), .ZN(n5263) );
  AOI22_X1 U6386 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5916), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5189), .ZN(n5256) );
  NOR2_X1 U6387 ( .A1(n6747), .A2(n6074), .ZN(n5191) );
  INV_X1 U6388 ( .A(n6132), .ZN(n5255) );
  AOI222_X1 U6389 ( .A1(n5192), .A2(n5260), .B1(n5256), .B2(n5191), .C1(n5190), 
        .C2(n5255), .ZN(n5193) );
  OAI22_X1 U6390 ( .A1(n5195), .A2(n5194), .B1(n5263), .B2(n5193), .ZN(U3460)
         );
  AND2_X1 U6391 ( .A1(n6490), .A2(REIP_REG_30__SCAN_IN), .ZN(n5923) );
  NOR2_X1 U6392 ( .A1(n5196), .A2(n6461), .ZN(n5197) );
  AOI211_X1 U6393 ( .C1(n6450), .C2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5923), 
        .B(n5197), .ZN(n5239) );
  INV_X1 U6394 ( .A(n5198), .ZN(n5199) );
  AND2_X1 U6395 ( .A1(n5208), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6423)
         );
  NAND2_X1 U6396 ( .A1(n5201), .A2(n3920), .ZN(n5207) );
  INV_X1 U6397 ( .A(n5202), .ZN(n5204) );
  NAND2_X1 U6398 ( .A1(n5204), .A2(n5203), .ZN(n5218) );
  XNOR2_X1 U6399 ( .A(n5218), .B(n5215), .ZN(n5205) );
  NAND2_X1 U6400 ( .A1(n5205), .A2(n5216), .ZN(n5206) );
  NAND2_X1 U6401 ( .A1(n5207), .A2(n5206), .ZN(n5213) );
  XNOR2_X1 U6402 ( .A(n5213), .B(n6493), .ZN(n6424) );
  NAND2_X1 U6403 ( .A1(n5213), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5865)
         );
  NAND2_X1 U6404 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  OR2_X1 U6405 ( .A1(n5218), .A2(n5217), .ZN(n5219) );
  NAND2_X1 U6406 ( .A1(n5214), .A2(n5219), .ZN(n5866) );
  NAND2_X1 U6407 ( .A1(n5866), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5862)
         );
  NAND3_X1 U6408 ( .A1(n6425), .A2(n5865), .A3(n5862), .ZN(n5222) );
  XNOR2_X1 U6409 ( .A(n5214), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5863)
         );
  OR2_X1 U6410 ( .A1(n5866), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5220)
         );
  AND2_X1 U6411 ( .A1(n5863), .A2(n5220), .ZN(n5221) );
  INV_X1 U6412 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5223) );
  AND3_X1 U6413 ( .A1(n5223), .A2(n5837), .A3(n6468), .ZN(n5224) );
  OR2_X1 U6414 ( .A1(n5214), .A2(n5224), .ZN(n5225) );
  INV_X1 U6415 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U6416 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5226) );
  OAI21_X1 U6417 ( .B1(n6104), .B2(n5226), .A(n5214), .ZN(n5227) );
  INV_X1 U6418 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6077) );
  XNOR2_X1 U6419 ( .A(n3093), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5824)
         );
  NAND2_X1 U6420 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6421 ( .A1(n3093), .A2(n5228), .ZN(n5229) );
  INV_X1 U6422 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6040) );
  NAND4_X1 U6423 ( .A1(n6049), .A2(n6040), .A3(n6063), .A4(n6068), .ZN(n5230)
         );
  NAND2_X1 U6424 ( .A1(n5610), .A2(n5230), .ZN(n5231) );
  NAND2_X1 U6425 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5896) );
  OAI21_X1 U6426 ( .B1(n6063), .B2(n5896), .A(n5214), .ZN(n5233) );
  AND2_X1 U6427 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6021) );
  AND2_X1 U6428 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U6429 ( .A1(n6021), .A2(n5899), .ZN(n5620) );
  NAND2_X1 U6430 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5910) );
  NOR2_X1 U6431 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6022) );
  NOR2_X1 U6432 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5978) );
  INV_X1 U6433 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5997) );
  XNOR2_X1 U6434 ( .A(n3093), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5601)
         );
  AOI21_X1 U6435 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5610), .ZN(n5234) );
  NOR2_X1 U6436 ( .A1(n3093), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5589)
         );
  NOR2_X1 U6437 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6438 ( .A1(n5589), .A2(n5235), .ZN(n5244) );
  INV_X1 U6439 ( .A(n5244), .ZN(n5236) );
  XNOR2_X1 U6440 ( .A(n5237), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5921)
         );
  NAND2_X1 U6441 ( .A1(n5921), .A2(n6455), .ZN(n5238) );
  OAI211_X1 U6442 ( .C1(n5243), .C2(n5886), .A(n5239), .B(n5238), .ZN(U2956)
         );
  AOI22_X1 U6443 ( .A1(n6340), .A2(DATAI_30_), .B1(n6345), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6444 ( .A1(n6342), .A2(DATAI_14_), .ZN(n5240) );
  OAI211_X1 U6445 ( .C1(n5243), .C2(n6148), .A(n5241), .B(n5240), .ZN(U2861)
         );
  INV_X1 U6446 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5242) );
  OAI222_X1 U6447 ( .A1(n5521), .A2(n5243), .B1(n5242), .B2(n6335), .C1(n5922), 
        .C2(n5519), .ZN(U2829) );
  AND2_X1 U6448 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5913) );
  NOR4_X1 U6449 ( .A1(n5600), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n5244), .ZN(n5245) );
  AOI21_X1 U6450 ( .B1(n5553), .B2(n5913), .A(n5245), .ZN(n5246) );
  XNOR2_X1 U6451 ( .A(n5246), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5887)
         );
  NAND2_X1 U6452 ( .A1(n6490), .A2(REIP_REG_31__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U6453 ( .A1(n6450), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5247)
         );
  OAI211_X1 U6454 ( .C1(n5248), .C2(n6461), .A(n5915), .B(n5247), .ZN(n5249)
         );
  AOI21_X1 U6455 ( .B1(n5887), .B2(n6455), .A(n5249), .ZN(n5250) );
  OAI21_X1 U6456 ( .B1(n5254), .B2(n5886), .A(n5250), .ZN(U2955) );
  NAND2_X1 U6457 ( .A1(n6354), .A2(n5251), .ZN(n5253) );
  AOI22_X1 U6458 ( .A1(n6340), .A2(DATAI_31_), .B1(n6345), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5252) );
  OAI21_X1 U6459 ( .B1(n5254), .B2(n5253), .A(n5252), .ZN(U2860) );
  AOI21_X1 U6460 ( .B1(n5255), .B2(n5257), .A(n5263), .ZN(n5265) );
  NOR3_X1 U6461 ( .A1(n6747), .A2(n6074), .A3(n5256), .ZN(n5259) );
  NOR3_X1 U6462 ( .A1(n6132), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5257), 
        .ZN(n5258) );
  AOI211_X1 U6463 ( .C1(n5261), .C2(n5260), .A(n5259), .B(n5258), .ZN(n5262)
         );
  OAI22_X1 U6464 ( .A1(n5265), .A2(n5264), .B1(n5263), .B2(n5262), .ZN(U3459)
         );
  OR2_X1 U6465 ( .A1(n5392), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5268) );
  INV_X1 U6466 ( .A(n5266), .ZN(n5267) );
  MUX2_X1 U6467 ( .A(n5268), .B(n5267), .S(n6794), .Z(U3474) );
  MUX2_X1 U6468 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6137), .Z(U3473) );
  INV_X1 U6469 ( .A(n5272), .ZN(n5277) );
  OAI21_X1 U6470 ( .B1(n5286), .B2(n5273), .A(n2983), .ZN(n5941) );
  AOI22_X1 U6471 ( .A1(n6303), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6306), .ZN(n5274) );
  OAI21_X1 U6472 ( .B1(n5941), .B2(n6260), .A(n5274), .ZN(n5276) );
  NOR2_X1 U6473 ( .A1(n6299), .A2(n5572), .ZN(n5275) );
  AOI211_X1 U6474 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5277), .A(n5276), .B(n5275), .ZN(n5280) );
  NAND3_X1 U6475 ( .A1(n5278), .A2(REIP_REG_27__SCAN_IN), .A3(n5793), .ZN(
        n5279) );
  OAI211_X1 U6476 ( .C1(n5571), .C2(n6282), .A(n5280), .B(n5279), .ZN(U2799)
         );
  AOI21_X1 U6477 ( .B1(n5282), .B2(n5281), .A(n5269), .ZN(n5585) );
  NAND2_X1 U6478 ( .A1(n5585), .A2(n6266), .ZN(n5292) );
  NOR2_X1 U6479 ( .A1(n5283), .A2(n5284), .ZN(n5285) );
  AOI22_X1 U6480 ( .A1(n6303), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6306), .ZN(n5287) );
  OAI21_X1 U6481 ( .B1(n5948), .B2(n6260), .A(n5287), .ZN(n5290) );
  NOR2_X1 U6482 ( .A1(n5300), .A2(n5288), .ZN(n5289) );
  AOI211_X1 U6483 ( .C1(n6311), .C2(n5581), .A(n5290), .B(n5289), .ZN(n5291)
         );
  OAI211_X1 U6484 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5293), .A(n5292), .B(n5291), .ZN(U2800) );
  OAI21_X1 U6485 ( .B1(n5294), .B2(n5295), .A(n5281), .ZN(n5596) );
  INV_X1 U6486 ( .A(n5587), .ZN(n5305) );
  NOR2_X1 U6487 ( .A1(n5296), .A2(n5297), .ZN(n5298) );
  OR2_X1 U6488 ( .A1(n5283), .A2(n5298), .ZN(n5959) );
  AOI22_X1 U6489 ( .A1(n6303), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6306), .ZN(n5299) );
  OAI21_X1 U6490 ( .B1(n5959), .B2(n6260), .A(n5299), .ZN(n5304) );
  NAND3_X1 U6491 ( .A1(n5330), .A2(REIP_REG_25__SCAN_IN), .A3(
        REIP_REG_24__SCAN_IN), .ZN(n5302) );
  AOI21_X1 U6492 ( .B1(n5302), .B2(n5301), .A(n5300), .ZN(n5303) );
  AOI211_X1 U6493 ( .C1(n6311), .C2(n5305), .A(n5304), .B(n5303), .ZN(n5306)
         );
  OAI21_X1 U6494 ( .B1(n5596), .B2(n6282), .A(n5306), .ZN(U2801) );
  AOI21_X1 U6496 ( .B1(n5309), .B2(n5308), .A(n5294), .ZN(n5310) );
  INV_X1 U6497 ( .A(n5310), .ZN(n5605) );
  INV_X1 U6498 ( .A(n5296), .ZN(n5313) );
  NAND2_X1 U6499 ( .A1(n5323), .A2(n5311), .ZN(n5312) );
  NAND2_X1 U6500 ( .A1(n5313), .A2(n5312), .ZN(n5969) );
  NAND2_X1 U6501 ( .A1(n5342), .A2(REIP_REG_25__SCAN_IN), .ZN(n5315) );
  AOI22_X1 U6502 ( .A1(n6303), .A2(EBX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6306), .ZN(n5314) );
  OAI211_X1 U6503 ( .C1(n5969), .C2(n6260), .A(n5315), .B(n5314), .ZN(n5316)
         );
  AOI21_X1 U6504 ( .B1(n6311), .B2(n5599), .A(n5316), .ZN(n5319) );
  XOR2_X1 U6505 ( .A(REIP_REG_25__SCAN_IN), .B(REIP_REG_24__SCAN_IN), .Z(n5317) );
  NAND2_X1 U6506 ( .A1(n5330), .A2(n5317), .ZN(n5318) );
  OAI211_X1 U6507 ( .C1(n5605), .C2(n6282), .A(n5319), .B(n5318), .ZN(U2802)
         );
  OAI21_X1 U6508 ( .B1(n5320), .B2(n5321), .A(n5308), .ZN(n5613) );
  OAI21_X1 U6509 ( .B1(n5322), .B2(n5324), .A(n5323), .ZN(n5974) );
  OAI22_X1 U6510 ( .A1(n5974), .A2(n6260), .B1(n5615), .B2(n6294), .ZN(n5325)
         );
  AOI21_X1 U6511 ( .B1(EBX_REG_24__SCAN_IN), .B2(n6229), .A(n5325), .ZN(n5327)
         );
  NAND2_X1 U6512 ( .A1(n5342), .A2(REIP_REG_24__SCAN_IN), .ZN(n5326) );
  OAI211_X1 U6513 ( .C1(n6299), .C2(n5614), .A(n5327), .B(n5326), .ZN(n5328)
         );
  AOI21_X1 U6514 ( .B1(n5330), .B2(n5329), .A(n5328), .ZN(n5331) );
  OAI21_X1 U6515 ( .B1(n5613), .B2(n6282), .A(n5331), .ZN(U2803) );
  INV_X1 U6516 ( .A(n5332), .ZN(n5347) );
  AOI21_X1 U6517 ( .B1(n5333), .B2(n5347), .A(n5320), .ZN(n5628) );
  INV_X1 U6518 ( .A(n5628), .ZN(n5538) );
  NAND2_X1 U6519 ( .A1(n5334), .A2(n5335), .ZN(n5336) );
  NAND2_X1 U6520 ( .A1(n5337), .A2(n5336), .ZN(n5985) );
  OAI22_X1 U6521 ( .A1(n5985), .A2(n6260), .B1(n5626), .B2(n6294), .ZN(n5340)
         );
  INV_X1 U6522 ( .A(n5624), .ZN(n5338) );
  NOR2_X1 U6523 ( .A1(n6299), .A2(n5338), .ZN(n5339) );
  AOI211_X1 U6524 ( .C1(EBX_REG_23__SCAN_IN), .C2(n6229), .A(n5340), .B(n5339), 
        .ZN(n5345) );
  INV_X1 U6525 ( .A(n5358), .ZN(n5370) );
  NOR2_X1 U6526 ( .A1(n5370), .A2(n5341), .ZN(n5343) );
  OAI21_X1 U6527 ( .B1(n5343), .B2(REIP_REG_23__SCAN_IN), .A(n5342), .ZN(n5344) );
  OAI211_X1 U6528 ( .C1(n5538), .C2(n6282), .A(n5345), .B(n5344), .ZN(U2804)
         );
  AOI21_X1 U6529 ( .B1(n5348), .B2(n5346), .A(n5332), .ZN(n5636) );
  INV_X1 U6530 ( .A(n5636), .ZN(n5541) );
  XOR2_X1 U6531 ( .A(REIP_REG_21__SCAN_IN), .B(REIP_REG_22__SCAN_IN), .Z(n5357) );
  OAI21_X1 U6532 ( .B1(n5363), .B2(n5350), .A(n5334), .ZN(n5993) );
  OAI22_X1 U6533 ( .A1(n6260), .A2(n5993), .B1(n5351), .B2(n6294), .ZN(n5354)
         );
  NOR2_X1 U6534 ( .A1(n5383), .A2(n5352), .ZN(n5353) );
  AOI211_X1 U6535 ( .C1(EBX_REG_22__SCAN_IN), .C2(n6229), .A(n5354), .B(n5353), 
        .ZN(n5355) );
  OAI21_X1 U6536 ( .B1(n6299), .B2(n5634), .A(n5355), .ZN(n5356) );
  AOI21_X1 U6537 ( .B1(n5358), .B2(n5357), .A(n5356), .ZN(n5359) );
  OAI21_X1 U6538 ( .B1(n5541), .B2(n6282), .A(n5359), .ZN(U2805) );
  XOR2_X1 U6539 ( .A(n5362), .B(n5361), .Z(n5644) );
  INV_X1 U6540 ( .A(n5644), .ZN(n5544) );
  INV_X1 U6541 ( .A(n5363), .ZN(n5364) );
  OAI21_X1 U6542 ( .B1(n5366), .B2(n5365), .A(n5364), .ZN(n6004) );
  OAI22_X1 U6543 ( .A1(n6260), .A2(n6004), .B1(n5642), .B2(n6294), .ZN(n5367)
         );
  AOI21_X1 U6544 ( .B1(EBX_REG_21__SCAN_IN), .B2(n6229), .A(n5367), .ZN(n5368)
         );
  OAI21_X1 U6545 ( .B1(n5383), .B2(n5369), .A(n5368), .ZN(n5372) );
  NOR2_X1 U6546 ( .A1(n5370), .A2(REIP_REG_21__SCAN_IN), .ZN(n5371) );
  AOI211_X1 U6547 ( .C1(n6311), .C2(n5640), .A(n5372), .B(n5371), .ZN(n5373)
         );
  OAI21_X1 U6548 ( .B1(n5544), .B2(n6282), .A(n5373), .ZN(U2806) );
  AND2_X1 U6549 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  NOR2_X1 U6550 ( .A1(n5361), .A2(n5376), .ZN(n6149) );
  INV_X1 U6551 ( .A(n6149), .ZN(n5483) );
  MUX2_X1 U6552 ( .A(n5486), .B(n5377), .S(n2995), .Z(n5378) );
  XOR2_X1 U6553 ( .A(n5379), .B(n5378), .Z(n6020) );
  NOR2_X1 U6554 ( .A1(n6020), .A2(n6260), .ZN(n5381) );
  OAI22_X1 U6555 ( .A1(n6259), .A2(n5482), .B1(n5650), .B2(n6294), .ZN(n5380)
         );
  AOI211_X1 U6556 ( .C1(n6311), .C2(n5648), .A(n5381), .B(n5380), .ZN(n5387)
         );
  NAND2_X1 U6557 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n6140) );
  INV_X1 U6558 ( .A(n5382), .ZN(n6179) );
  OAI21_X1 U6559 ( .B1(n6140), .B2(n6179), .A(n4197), .ZN(n5385) );
  INV_X1 U6560 ( .A(n5383), .ZN(n5384) );
  NAND2_X1 U6561 ( .A1(n5385), .A2(n5384), .ZN(n5386) );
  OAI211_X1 U6562 ( .C1(n5483), .C2(n6282), .A(n5387), .B(n5386), .ZN(U2807)
         );
  OAI21_X1 U6563 ( .B1(n5388), .B2(n5390), .A(n5389), .ZN(n5673) );
  INV_X1 U6564 ( .A(n5391), .ZN(n6183) );
  OAI21_X1 U6565 ( .B1(n6205), .B2(n6199), .A(n4230), .ZN(n5401) );
  NAND2_X1 U6566 ( .A1(n6233), .A2(n5392), .ZN(n6308) );
  INV_X1 U6567 ( .A(n6308), .ZN(n6263) );
  NAND2_X1 U6568 ( .A1(n5393), .A2(n5394), .ZN(n5395) );
  NAND2_X1 U6569 ( .A1(n2985), .A2(n5395), .ZN(n6045) );
  NOR2_X1 U6570 ( .A1(n6260), .A2(n6045), .ZN(n5396) );
  AOI211_X1 U6571 ( .C1(n6306), .C2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n6263), 
        .B(n5396), .ZN(n5397) );
  OAI21_X1 U6572 ( .B1(n5398), .B2(n6259), .A(n5397), .ZN(n5400) );
  NOR2_X1 U6573 ( .A1(n6299), .A2(n5675), .ZN(n5399) );
  AOI211_X1 U6574 ( .C1(n6183), .C2(n5401), .A(n5400), .B(n5399), .ZN(n5402)
         );
  OAI21_X1 U6575 ( .B1(n5673), .B2(n6282), .A(n5402), .ZN(U2810) );
  AOI22_X1 U6576 ( .A1(n6305), .A2(n6472), .B1(n6229), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5403) );
  OAI21_X1 U6577 ( .B1(n6299), .B2(n5869), .A(n5403), .ZN(n5408) );
  INV_X1 U6578 ( .A(n6233), .ZN(n5453) );
  INV_X1 U6579 ( .A(n5404), .ZN(n5405) );
  NOR2_X1 U6580 ( .A1(n6289), .A2(n5405), .ZN(n5415) );
  OR2_X1 U6581 ( .A1(n5453), .A2(n5415), .ZN(n6267) );
  NOR2_X1 U6582 ( .A1(n6289), .A2(REIP_REG_9__SCAN_IN), .ZN(n6268) );
  AOI22_X1 U6583 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6267), .B1(n5405), .B2(n6268), .ZN(n5406) );
  OAI211_X1 U6584 ( .C1(n6294), .C2(n5728), .A(n5406), .B(n6308), .ZN(n5407)
         );
  NOR2_X1 U6585 ( .A1(n5408), .A2(n5407), .ZN(n5409) );
  OAI21_X1 U6586 ( .B1(n6282), .B2(n5873), .A(n5409), .ZN(U2818) );
  NAND2_X1 U6587 ( .A1(n6311), .A2(n5881), .ZN(n5417) );
  AOI22_X1 U6588 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6306), .B1(
        EBX_REG_8__SCAN_IN), .B2(n6303), .ZN(n5410) );
  OAI211_X1 U6589 ( .C1(n6260), .C2(n5411), .A(n5410), .B(n6308), .ZN(n5413)
         );
  AND2_X1 U6590 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6267), .ZN(n5412) );
  AOI211_X1 U6591 ( .C1(n5415), .C2(n5414), .A(n5413), .B(n5412), .ZN(n5416)
         );
  OAI211_X1 U6592 ( .C1(n5885), .C2(n6282), .A(n5417), .B(n5416), .ZN(U2819)
         );
  AOI22_X1 U6593 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6306), .B1(n6305), 
        .B2(n6499), .ZN(n5418) );
  NAND2_X1 U6594 ( .A1(n5418), .A2(n6308), .ZN(n5425) );
  OAI21_X1 U6595 ( .B1(n6289), .B2(n5419), .A(n6233), .ZN(n6291) );
  INV_X1 U6596 ( .A(n6291), .ZN(n5423) );
  NAND2_X1 U6597 ( .A1(n5422), .A2(n5419), .ZN(n5420) );
  NOR2_X1 U6598 ( .A1(n6289), .A2(n5420), .ZN(n6284) );
  AOI21_X1 U6599 ( .B1(EBX_REG_6__SCAN_IN), .B2(n6229), .A(n6284), .ZN(n5421)
         );
  OAI21_X1 U6600 ( .B1(n5423), .B2(n5422), .A(n5421), .ZN(n5424) );
  AOI211_X1 U6601 ( .C1(n6266), .C2(n5426), .A(n5425), .B(n5424), .ZN(n5427)
         );
  OAI21_X1 U6602 ( .B1(n5428), .B2(n6299), .A(n5427), .ZN(U2821) );
  INV_X1 U6603 ( .A(n5435), .ZN(n5429) );
  INV_X1 U6604 ( .A(n6448), .ZN(n5441) );
  NAND2_X1 U6605 ( .A1(n6233), .A2(REIP_REG_2__SCAN_IN), .ZN(n5430) );
  AOI21_X1 U6606 ( .B1(n6319), .B2(n6782), .A(n5430), .ZN(n5443) );
  NAND2_X1 U6607 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .ZN(
        n6315) );
  OAI21_X1 U6608 ( .B1(n6315), .B2(n5430), .A(n6191), .ZN(n5431) );
  INV_X1 U6609 ( .A(n5431), .ZN(n6302) );
  OAI21_X1 U6610 ( .B1(n5443), .B2(REIP_REG_3__SCAN_IN), .A(n6302), .ZN(n5439)
         );
  AOI21_X1 U6611 ( .B1(n5433), .B2(n4424), .A(n5432), .ZN(n6520) );
  AOI22_X1 U6612 ( .A1(n6305), .A2(n6520), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n6306), .ZN(n5438) );
  NOR2_X1 U6613 ( .A1(n5435), .A2(n5434), .ZN(n6300) );
  NAND2_X1 U6614 ( .A1(n6300), .A2(n2977), .ZN(n5437) );
  NAND2_X1 U6615 ( .A1(n6303), .A2(EBX_REG_3__SCAN_IN), .ZN(n5436) );
  NAND4_X1 U6616 ( .A1(n5439), .A2(n5438), .A3(n5437), .A4(n5436), .ZN(n5440)
         );
  AOI21_X1 U6617 ( .B1(n5441), .B2(n6311), .A(n5440), .ZN(n5442) );
  OAI21_X1 U6618 ( .B1(n6292), .B2(n6330), .A(n5442), .ZN(U2824) );
  INV_X1 U6619 ( .A(n6460), .ZN(n5450) );
  INV_X1 U6620 ( .A(n5443), .ZN(n5445) );
  OAI21_X1 U6621 ( .B1(n6289), .B2(n6782), .A(n6316), .ZN(n5444) );
  AOI22_X1 U6622 ( .A1(n5445), .A2(n5444), .B1(EBX_REG_2__SCAN_IN), .B2(n6229), 
        .ZN(n5448) );
  AOI22_X1 U6623 ( .A1(n6300), .A2(n5446), .B1(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6306), .ZN(n5447) );
  OAI211_X1 U6624 ( .C1(n6260), .C2(n6529), .A(n5448), .B(n5447), .ZN(n5449)
         );
  AOI21_X1 U6625 ( .B1(n6311), .B2(n5450), .A(n5449), .ZN(n5451) );
  OAI21_X1 U6626 ( .B1(n6292), .B2(n6451), .A(n5451), .ZN(U2825) );
  NAND2_X1 U6627 ( .A1(n6300), .A2(n5452), .ZN(n5455) );
  NAND2_X1 U6628 ( .A1(n5453), .A2(REIP_REG_1__SCAN_IN), .ZN(n5454) );
  OAI211_X1 U6629 ( .C1(REIP_REG_1__SCAN_IN), .C2(n6289), .A(n5455), .B(n5454), 
        .ZN(n5458) );
  NOR2_X1 U6630 ( .A1(n6259), .A2(n5456), .ZN(n5457) );
  AOI211_X1 U6631 ( .C1(n6305), .C2(n5459), .A(n5458), .B(n5457), .ZN(n5462)
         );
  MUX2_X1 U6632 ( .A(n6311), .B(n6306), .S(PHYADDRPOINTER_REG_1__SCAN_IN), .Z(
        n5460) );
  INV_X1 U6633 ( .A(n5460), .ZN(n5461) );
  OAI211_X1 U6634 ( .C1(n6292), .C2(n5463), .A(n5462), .B(n5461), .ZN(U2826)
         );
  NOR2_X1 U6635 ( .A1(n6260), .A2(n5464), .ZN(n5467) );
  OAI22_X1 U6636 ( .A1(n6259), .A2(n5465), .B1(n6232), .B2(n6788), .ZN(n5466)
         );
  AOI211_X1 U6637 ( .C1(n6300), .C2(n3466), .A(n5467), .B(n5466), .ZN(n5469)
         );
  OAI21_X1 U6638 ( .B1(n6311), .B2(n6306), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5468) );
  OAI211_X1 U6639 ( .C1(n6292), .C2(n5470), .A(n5469), .B(n5468), .ZN(U2827)
         );
  INV_X1 U6640 ( .A(n5918), .ZN(n5471) );
  OAI22_X1 U6641 ( .A1(n5471), .A2(n5519), .B1(n6335), .B2(n5766), .ZN(U2828)
         );
  AOI22_X1 U6642 ( .A1(n5472), .A2(n6331), .B1(EBX_REG_29__SCAN_IN), .B2(n5504), .ZN(n5473) );
  OAI21_X1 U6643 ( .B1(n4100), .B2(n5521), .A(n5473), .ZN(U2830) );
  OAI222_X1 U6644 ( .A1(n5571), .A2(n5521), .B1(n5474), .B2(n6335), .C1(n5941), 
        .C2(n5519), .ZN(U2831) );
  INV_X1 U6645 ( .A(n5585), .ZN(n5529) );
  OAI222_X1 U6646 ( .A1(n5521), .A2(n5529), .B1(n5475), .B2(n6335), .C1(n5948), 
        .C2(n5519), .ZN(U2832) );
  OAI222_X1 U6647 ( .A1(n5596), .A2(n5521), .B1(n5476), .B2(n6335), .C1(n5959), 
        .C2(n5519), .ZN(U2833) );
  INV_X1 U6648 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5477) );
  OAI222_X1 U6649 ( .A1(n5969), .A2(n5519), .B1(n5477), .B2(n6335), .C1(n5605), 
        .C2(n5521), .ZN(U2834) );
  INV_X1 U6650 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5478) );
  OAI222_X1 U6651 ( .A1(n5521), .A2(n5613), .B1(n5478), .B2(n6335), .C1(n5974), 
        .C2(n5519), .ZN(U2835) );
  OAI222_X1 U6652 ( .A1(n5521), .A2(n5538), .B1(n5479), .B2(n6335), .C1(n5985), 
        .C2(n5519), .ZN(U2836) );
  INV_X1 U6653 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5480) );
  OAI222_X1 U6654 ( .A1(n5521), .A2(n5541), .B1(n5480), .B2(n6335), .C1(n5993), 
        .C2(n5519), .ZN(U2837) );
  INV_X1 U6655 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5481) );
  OAI222_X1 U6656 ( .A1(n5544), .A2(n5521), .B1(n5481), .B2(n6335), .C1(n6004), 
        .C2(n5519), .ZN(U2838) );
  OAI222_X1 U6657 ( .A1(n5483), .A2(n5521), .B1(n5482), .B2(n6335), .C1(n5519), 
        .C2(n6020), .ZN(U2839) );
  XNOR2_X1 U6658 ( .A(n2986), .B(n5484), .ZN(n6152) );
  INV_X1 U6659 ( .A(n6152), .ZN(n5489) );
  MUX2_X1 U6660 ( .A(n5486), .B(n5485), .S(n6802), .Z(n5491) );
  XNOR2_X1 U6661 ( .A(n5493), .B(n5487), .ZN(n6143) );
  AOI22_X1 U6662 ( .A1(n6331), .A2(n6143), .B1(EBX_REG_19__SCAN_IN), .B2(n5504), .ZN(n5488) );
  OAI21_X1 U6663 ( .B1(n5489), .B2(n5521), .A(n5488), .ZN(U2840) );
  AOI21_X1 U6664 ( .B1(n5490), .B2(n5389), .A(n2986), .ZN(n6336) );
  INV_X1 U6665 ( .A(n6336), .ZN(n5495) );
  NAND2_X1 U6666 ( .A1(n2985), .A2(n5491), .ZN(n5492) );
  NAND2_X1 U6667 ( .A1(n5493), .A2(n5492), .ZN(n6189) );
  OAI222_X1 U6668 ( .A1(n5495), .A2(n5521), .B1(n5494), .B2(n6335), .C1(n6189), 
        .C2(n5519), .ZN(U2841) );
  INV_X1 U6669 ( .A(n6045), .ZN(n5496) );
  AOI22_X1 U6670 ( .A1(n6331), .A2(n5496), .B1(EBX_REG_17__SCAN_IN), .B2(n5504), .ZN(n5497) );
  OAI21_X1 U6671 ( .B1(n5673), .B2(n5521), .A(n5497), .ZN(U2842) );
  AND2_X1 U6672 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  OR2_X1 U6673 ( .A1(n5500), .A2(n5388), .ZN(n6339) );
  OR2_X1 U6674 ( .A1(n5501), .A2(n5502), .ZN(n5503) );
  AND2_X1 U6675 ( .A1(n5393), .A2(n5503), .ZN(n6196) );
  AOI22_X1 U6676 ( .A1(n6331), .A2(n6196), .B1(EBX_REG_16__SCAN_IN), .B2(n5504), .ZN(n5505) );
  OAI21_X1 U6677 ( .B1(n6339), .B2(n5521), .A(n5505), .ZN(U2843) );
  OR2_X1 U6678 ( .A1(n5507), .A2(n5508), .ZN(n5509) );
  NAND2_X1 U6679 ( .A1(n5506), .A2(n5509), .ZN(n6219) );
  INV_X1 U6680 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5515) );
  OR2_X1 U6681 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  NAND2_X1 U6682 ( .A1(n5511), .A2(n5514), .ZN(n6222) );
  OAI222_X1 U6683 ( .A1(n6219), .A2(n5519), .B1(n5515), .B2(n6335), .C1(n6222), 
        .C2(n5521), .ZN(U2845) );
  AOI21_X1 U6684 ( .B1(n5516), .B2(n5180), .A(n2978), .ZN(n6352) );
  INV_X1 U6685 ( .A(n6352), .ZN(n5522) );
  INV_X1 U6686 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5520) );
  AND2_X1 U6687 ( .A1(n3112), .A2(n5517), .ZN(n5518) );
  OR2_X1 U6688 ( .A1(n5518), .A2(n6091), .ZN(n6238) );
  OAI222_X1 U6689 ( .A1(n5522), .A2(n5521), .B1(n5520), .B2(n6335), .C1(n6238), 
        .C2(n5519), .ZN(U2847) );
  AOI22_X1 U6690 ( .A1(n6340), .A2(DATAI_29_), .B1(n6345), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6691 ( .A1(n6342), .A2(DATAI_13_), .ZN(n5523) );
  OAI211_X1 U6692 ( .C1(n4100), .C2(n6148), .A(n5524), .B(n5523), .ZN(U2862)
         );
  AOI22_X1 U6693 ( .A1(n6340), .A2(DATAI_28_), .B1(n6345), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6694 ( .A1(n6342), .A2(DATAI_12_), .ZN(n5525) );
  OAI211_X1 U6695 ( .C1(n5571), .C2(n6148), .A(n5526), .B(n5525), .ZN(U2863)
         );
  AOI22_X1 U6696 ( .A1(n6340), .A2(DATAI_27_), .B1(n6345), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U6697 ( .A1(n6342), .A2(DATAI_11_), .ZN(n5527) );
  OAI211_X1 U6698 ( .C1(n5529), .C2(n6148), .A(n5528), .B(n5527), .ZN(U2864)
         );
  AOI22_X1 U6699 ( .A1(n6340), .A2(DATAI_26_), .B1(n6345), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U6700 ( .A1(n6342), .A2(DATAI_10_), .ZN(n5530) );
  OAI211_X1 U6701 ( .C1(n5596), .C2(n6148), .A(n5531), .B(n5530), .ZN(U2865)
         );
  AOI22_X1 U6702 ( .A1(n6340), .A2(DATAI_25_), .B1(n6345), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U6703 ( .A1(n6342), .A2(DATAI_9_), .ZN(n5532) );
  OAI211_X1 U6704 ( .C1(n5605), .C2(n6148), .A(n5533), .B(n5532), .ZN(U2866)
         );
  AOI22_X1 U6705 ( .A1(n6340), .A2(DATAI_24_), .B1(n6345), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6706 ( .A1(n6342), .A2(DATAI_8_), .ZN(n5534) );
  OAI211_X1 U6707 ( .C1(n5613), .C2(n6148), .A(n5535), .B(n5534), .ZN(U2867)
         );
  AOI22_X1 U6708 ( .A1(n6340), .A2(DATAI_23_), .B1(n6345), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U6709 ( .A1(n6342), .A2(DATAI_7_), .ZN(n5536) );
  OAI211_X1 U6710 ( .C1(n5538), .C2(n6148), .A(n5537), .B(n5536), .ZN(U2868)
         );
  AOI22_X1 U6711 ( .A1(n6340), .A2(DATAI_22_), .B1(n6345), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U6712 ( .A1(n6342), .A2(DATAI_6_), .ZN(n5539) );
  OAI211_X1 U6713 ( .C1(n5541), .C2(n6148), .A(n5540), .B(n5539), .ZN(U2869)
         );
  AOI22_X1 U6714 ( .A1(n6340), .A2(DATAI_21_), .B1(n6345), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U6715 ( .A1(n6342), .A2(DATAI_5_), .ZN(n5542) );
  OAI211_X1 U6716 ( .C1(n5544), .C2(n6148), .A(n5543), .B(n5542), .ZN(U2870)
         );
  AOI22_X1 U6717 ( .A1(n6340), .A2(DATAI_17_), .B1(n6345), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U6718 ( .A1(n6342), .A2(DATAI_1_), .ZN(n5545) );
  OAI211_X1 U6719 ( .C1(n5673), .C2(n6148), .A(n5546), .B(n5545), .ZN(U2874)
         );
  AOI22_X1 U6720 ( .A1(n6350), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6345), .ZN(n5547) );
  OAI21_X1 U6721 ( .B1(n6222), .B2(n6148), .A(n5547), .ZN(U2877) );
  INV_X1 U6722 ( .A(DATAI_13_), .ZN(n5550) );
  XNOR2_X1 U6723 ( .A(n2978), .B(n5548), .ZN(n6327) );
  INV_X1 U6724 ( .A(n6327), .ZN(n5549) );
  OAI222_X1 U6725 ( .A1(n6354), .A2(n5551), .B1(n5550), .B2(n6349), .C1(n6148), 
        .C2(n5549), .ZN(U2878) );
  INV_X1 U6726 ( .A(n5553), .ZN(n5557) );
  INV_X1 U6727 ( .A(n5552), .ZN(n5556) );
  INV_X1 U6728 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5934) );
  INV_X1 U6731 ( .A(n5558), .ZN(n5937) );
  NAND2_X1 U6732 ( .A1(n5559), .A2(n5882), .ZN(n5560) );
  NAND2_X1 U6733 ( .A1(n6490), .A2(REIP_REG_29__SCAN_IN), .ZN(n5931) );
  OAI211_X1 U6734 ( .C1(n5879), .C2(n5561), .A(n5560), .B(n5931), .ZN(n5562)
         );
  AOI21_X1 U6735 ( .B1(n5563), .B2(n6456), .A(n5562), .ZN(n5564) );
  OAI21_X1 U6736 ( .B1(n5937), .B2(n6161), .A(n5564), .ZN(U2957) );
  NAND2_X1 U6737 ( .A1(n5565), .A2(n5589), .ZN(n5567) );
  NAND2_X1 U6738 ( .A1(n3093), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U6739 ( .A1(n5579), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5566) );
  OAI21_X1 U6740 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5567), .A(n5566), 
        .ZN(n5570) );
  INV_X1 U6741 ( .A(n5567), .ZN(n5578) );
  NOR3_X1 U6742 ( .A1(n5578), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5939), 
        .ZN(n5569) );
  NAND2_X1 U6743 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5912) );
  NOR2_X1 U6744 ( .A1(n5579), .A2(n5912), .ZN(n5568) );
  INV_X1 U6745 ( .A(n5571), .ZN(n5576) );
  NOR2_X1 U6746 ( .A1(n5572), .A2(n6461), .ZN(n5575) );
  NAND2_X1 U6747 ( .A1(n6490), .A2(REIP_REG_28__SCAN_IN), .ZN(n5940) );
  OAI21_X1 U6748 ( .B1(n5879), .B2(n5573), .A(n5940), .ZN(n5574) );
  OAI21_X1 U6749 ( .B1(n5946), .B2(n6161), .A(n5577), .ZN(U2958) );
  NOR2_X1 U6750 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  XOR2_X1 U6751 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(n5580), .Z(n5955) );
  NAND2_X1 U6752 ( .A1(n5581), .A2(n5882), .ZN(n5582) );
  NAND2_X1 U6753 ( .A1(n6490), .A2(REIP_REG_27__SCAN_IN), .ZN(n5947) );
  OAI211_X1 U6754 ( .C1(n5879), .C2(n5583), .A(n5582), .B(n5947), .ZN(n5584)
         );
  AOI21_X1 U6755 ( .B1(n5585), .B2(n6456), .A(n5584), .ZN(n5586) );
  OAI21_X1 U6756 ( .B1(n5955), .B2(n6161), .A(n5586), .ZN(U2959) );
  AND2_X1 U6757 ( .A1(n6490), .A2(REIP_REG_26__SCAN_IN), .ZN(n5957) );
  NOR2_X1 U6758 ( .A1(n5587), .A2(n6461), .ZN(n5588) );
  AOI211_X1 U6759 ( .C1(n6450), .C2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5957), 
        .B(n5588), .ZN(n5595) );
  INV_X1 U6760 ( .A(n5589), .ZN(n5591) );
  NAND2_X1 U6761 ( .A1(n5591), .A2(n5590), .ZN(n5592) );
  XNOR2_X1 U6762 ( .A(n5593), .B(n5592), .ZN(n5956) );
  NAND2_X1 U6763 ( .A1(n5956), .A2(n6455), .ZN(n5594) );
  OAI211_X1 U6764 ( .C1(n5596), .C2(n5886), .A(n5595), .B(n5594), .ZN(U2960)
         );
  NAND2_X1 U6765 ( .A1(n6490), .A2(REIP_REG_25__SCAN_IN), .ZN(n5968) );
  OAI21_X1 U6766 ( .B1(n5879), .B2(n5597), .A(n5968), .ZN(n5598) );
  AOI21_X1 U6767 ( .B1(n5599), .B2(n5882), .A(n5598), .ZN(n5604) );
  OAI21_X1 U6768 ( .B1(n5602), .B2(n5601), .A(n5600), .ZN(n5967) );
  NAND2_X1 U6769 ( .A1(n5967), .A2(n6455), .ZN(n5603) );
  OAI211_X1 U6770 ( .C1(n5605), .C2(n5886), .A(n5604), .B(n5603), .ZN(U2961)
         );
  INV_X1 U6771 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6032) );
  AND2_X1 U6772 ( .A1(n3093), .A2(n6032), .ZN(n5655) );
  INV_X1 U6773 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U6774 ( .A1(n3093), .A2(n5607), .ZN(n5606) );
  OR2_X1 U6775 ( .A1(n3093), .A2(n5607), .ZN(n5608) );
  XNOR2_X1 U6776 ( .A(n3093), .B(n6007), .ZN(n5639) );
  OR2_X1 U6777 ( .A1(n3093), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5630)
         );
  NAND2_X1 U6778 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5609) );
  OR3_X1 U6779 ( .A1(n5631), .A2(n5610), .A3(n5609), .ZN(n5611) );
  XNOR2_X1 U6780 ( .A(n5612), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5983)
         );
  INV_X1 U6781 ( .A(n5613), .ZN(n5618) );
  NOR2_X1 U6782 ( .A1(n5614), .A2(n6461), .ZN(n5617) );
  NAND2_X1 U6783 ( .A1(n6490), .A2(REIP_REG_24__SCAN_IN), .ZN(n5975) );
  OAI21_X1 U6784 ( .B1(n5879), .B2(n5615), .A(n5975), .ZN(n5616) );
  AOI211_X1 U6785 ( .C1(n5618), .C2(n6456), .A(n5617), .B(n5616), .ZN(n5619)
         );
  OAI21_X1 U6786 ( .B1(n5983), .B2(n6161), .A(n5619), .ZN(U2962) );
  INV_X1 U6787 ( .A(n5620), .ZN(n5909) );
  NAND2_X1 U6788 ( .A1(n5653), .A2(n5909), .ZN(n5622) );
  OAI21_X1 U6789 ( .B1(n5657), .B2(n5622), .A(n5621), .ZN(n5623) );
  XNOR2_X1 U6790 ( .A(n5623), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5992)
         );
  NAND2_X1 U6791 ( .A1(n5624), .A2(n5882), .ZN(n5625) );
  NAND2_X1 U6792 ( .A1(n6490), .A2(REIP_REG_23__SCAN_IN), .ZN(n5984) );
  OAI211_X1 U6793 ( .C1(n5879), .C2(n5626), .A(n5625), .B(n5984), .ZN(n5627)
         );
  AOI21_X1 U6794 ( .B1(n5628), .B2(n6456), .A(n5627), .ZN(n5629) );
  OAI21_X1 U6795 ( .B1(n5992), .B2(n6161), .A(n5629), .ZN(U2963) );
  OAI21_X1 U6796 ( .B1(n5610), .B2(n5997), .A(n5630), .ZN(n5632) );
  XOR2_X1 U6797 ( .A(n5632), .B(n5631), .Z(n6001) );
  AND2_X1 U6798 ( .A1(n6490), .A2(REIP_REG_22__SCAN_IN), .ZN(n5994) );
  AOI21_X1 U6799 ( .B1(n6450), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5994), 
        .ZN(n5633) );
  OAI21_X1 U6800 ( .B1(n5634), .B2(n6461), .A(n5633), .ZN(n5635) );
  AOI21_X1 U6801 ( .B1(n5636), .B2(n6456), .A(n5635), .ZN(n5637) );
  OAI21_X1 U6802 ( .B1(n6001), .B2(n6161), .A(n5637), .ZN(U2964) );
  AOI21_X1 U6803 ( .B1(n5639), .B2(n5638), .A(n2993), .ZN(n6010) );
  NAND2_X1 U6804 ( .A1(n5640), .A2(n5882), .ZN(n5641) );
  NAND2_X1 U6805 ( .A1(n6490), .A2(REIP_REG_21__SCAN_IN), .ZN(n6003) );
  OAI211_X1 U6806 ( .C1(n5879), .C2(n5642), .A(n5641), .B(n6003), .ZN(n5643)
         );
  AOI21_X1 U6807 ( .B1(n5644), .B2(n6456), .A(n5643), .ZN(n5645) );
  OAI21_X1 U6808 ( .B1(n6010), .B2(n6161), .A(n5645), .ZN(U2965) );
  XNOR2_X1 U6809 ( .A(n3093), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5646)
         );
  XNOR2_X1 U6810 ( .A(n5647), .B(n5646), .ZN(n6027) );
  NAND2_X1 U6811 ( .A1(n5648), .A2(n5882), .ZN(n5649) );
  NAND2_X1 U6812 ( .A1(n6490), .A2(REIP_REG_20__SCAN_IN), .ZN(n6019) );
  OAI211_X1 U6813 ( .C1(n5879), .C2(n5650), .A(n5649), .B(n6019), .ZN(n5651)
         );
  AOI21_X1 U6814 ( .B1(n6149), .B2(n6456), .A(n5651), .ZN(n5652) );
  OAI21_X1 U6815 ( .B1(n6027), .B2(n6161), .A(n5652), .ZN(U2966) );
  OAI21_X1 U6816 ( .B1(n3036), .B2(n5655), .A(n5654), .ZN(n5656) );
  OAI21_X1 U6817 ( .B1(n5657), .B2(n3036), .A(n5656), .ZN(n6036) );
  NAND2_X1 U6818 ( .A1(n6142), .A2(n5882), .ZN(n5658) );
  NAND2_X1 U6819 ( .A1(n6490), .A2(REIP_REG_19__SCAN_IN), .ZN(n6028) );
  OAI211_X1 U6820 ( .C1(n5879), .C2(n5659), .A(n5658), .B(n6028), .ZN(n5660)
         );
  AOI21_X1 U6821 ( .B1(n6152), .B2(n6456), .A(n5660), .ZN(n5661) );
  OAI21_X1 U6822 ( .B1(n6161), .B2(n6036), .A(n5661), .ZN(U2967) );
  OAI21_X1 U6823 ( .B1(n5610), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5823), 
        .ZN(n5687) );
  XNOR2_X1 U6824 ( .A(n3093), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5686)
         );
  NAND2_X1 U6825 ( .A1(n5687), .A2(n5686), .ZN(n5685) );
  OAI21_X1 U6826 ( .B1(n5610), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5685), 
        .ZN(n5680) );
  AOI21_X1 U6827 ( .B1(n3093), .B2(n6063), .A(n5680), .ZN(n5667) );
  NAND3_X1 U6828 ( .A1(n5667), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n3093), .ZN(n5672) );
  INV_X1 U6829 ( .A(n5685), .ZN(n5662) );
  NOR2_X1 U6830 ( .A1(n3093), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5679)
         );
  NAND3_X1 U6831 ( .A1(n5662), .A2(n5679), .A3(n6049), .ZN(n5669) );
  NAND2_X1 U6832 ( .A1(n5672), .A2(n5669), .ZN(n5663) );
  XNOR2_X1 U6833 ( .A(n5663), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6043)
         );
  NAND2_X1 U6834 ( .A1(n6490), .A2(REIP_REG_18__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U6835 ( .A1(n6450), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5664)
         );
  OAI211_X1 U6836 ( .C1(n6186), .C2(n6461), .A(n6037), .B(n5664), .ZN(n5665)
         );
  AOI21_X1 U6837 ( .B1(n6336), .B2(n6456), .A(n5665), .ZN(n5666) );
  OAI21_X1 U6838 ( .B1(n6043), .B2(n6161), .A(n5666), .ZN(U2968) );
  OAI21_X1 U6839 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n3093), .A(n5667), 
        .ZN(n5668) );
  OAI21_X1 U6840 ( .B1(n5679), .B2(n6049), .A(n5668), .ZN(n5671) );
  INV_X1 U6841 ( .A(n5669), .ZN(n5670) );
  AOI21_X1 U6842 ( .B1(n5672), .B2(n5671), .A(n5670), .ZN(n6052) );
  INV_X1 U6843 ( .A(n5673), .ZN(n5677) );
  NAND2_X1 U6844 ( .A1(n6490), .A2(REIP_REG_17__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U6845 ( .A1(n6450), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5674)
         );
  OAI211_X1 U6846 ( .C1(n5675), .C2(n6461), .A(n6044), .B(n5674), .ZN(n5676)
         );
  AOI21_X1 U6847 ( .B1(n5677), .B2(n6456), .A(n5676), .ZN(n5678) );
  OAI21_X1 U6848 ( .B1(n6052), .B2(n6161), .A(n5678), .ZN(U2969) );
  AOI21_X1 U6849 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n3093), .A(n5679), 
        .ZN(n5681) );
  XOR2_X1 U6850 ( .A(n5681), .B(n5680), .Z(n6058) );
  NAND2_X1 U6851 ( .A1(n6058), .A2(n6455), .ZN(n5684) );
  AND2_X1 U6852 ( .A1(n6490), .A2(REIP_REG_16__SCAN_IN), .ZN(n6060) );
  NOR2_X1 U6853 ( .A1(n6461), .A2(n6193), .ZN(n5682) );
  AOI211_X1 U6854 ( .C1(n6450), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6060), 
        .B(n5682), .ZN(n5683) );
  OAI211_X1 U6855 ( .C1(n5886), .C2(n6339), .A(n5684), .B(n5683), .ZN(U2970)
         );
  OAI21_X1 U6856 ( .B1(n5687), .B2(n5686), .A(n5685), .ZN(n5688) );
  INV_X1 U6857 ( .A(n5688), .ZN(n6072) );
  XOR2_X1 U6858 ( .A(n5689), .B(n5511), .Z(n6346) );
  NOR2_X1 U6859 ( .A1(n6120), .A2(n6206), .ZN(n6070) );
  AOI21_X1 U6860 ( .B1(n6450), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6070), 
        .ZN(n5690) );
  OAI21_X1 U6861 ( .B1(n6211), .B2(n6461), .A(n5690), .ZN(n5691) );
  AOI21_X1 U6862 ( .B1(n6346), .B2(n6456), .A(n5691), .ZN(n5692) );
  OAI21_X1 U6863 ( .B1(n6072), .B2(n6161), .A(n5692), .ZN(U2971) );
  INV_X1 U6864 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5799) );
  NOR4_X1 U6865 ( .A1(EBX_REG_7__SCAN_IN), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), 
        .A3(ADDRESS_REG_21__SCAN_IN), .A4(n5799), .ZN(n5780) );
  NOR4_X1 U6866 ( .A1(EAX_REG_9__SCAN_IN), .A2(DATAI_25_), .A3(
        BYTEENABLE_REG_3__SCAN_IN), .A4(n5877), .ZN(n5702) );
  NAND3_X1 U6867 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(EBX_REG_24__SCAN_IN), 
        .A3(EAX_REG_12__SCAN_IN), .ZN(n5695) );
  NAND4_X1 U6868 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(
        INSTQUEUE_REG_15__2__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAO_REG_26__SCAN_IN), .ZN(n5694) );
  NAND4_X1 U6869 ( .A1(DATAI_6_), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .A3(
        DATAO_REG_30__SCAN_IN), .A4(n5812), .ZN(n5693) );
  NOR4_X1 U6870 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n5695), .A3(n5694), .A4(
        n5693), .ZN(n5701) );
  NOR4_X1 U6871 ( .A1(DATAI_26_), .A2(EBX_REG_4__SCAN_IN), .A3(
        BE_N_REG_0__SCAN_IN), .A4(n5997), .ZN(n5700) );
  INV_X1 U6872 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5736) );
  NAND3_X1 U6873 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(EAX_REG_20__SCAN_IN), 
        .A3(n5736), .ZN(n5698) );
  INV_X1 U6874 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5768) );
  NAND4_X1 U6875 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        DATAO_REG_19__SCAN_IN), .A3(n5768), .A4(n5769), .ZN(n5697) );
  NAND4_X1 U6876 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(
        INSTQUEUE_REG_9__5__SCAN_IN), .A3(EBX_REG_31__SCAN_IN), .A4(
        DATAWIDTH_REG_7__SCAN_IN), .ZN(n5696) );
  NOR4_X1 U6877 ( .A1(ADDRESS_REG_12__SCAN_IN), .A2(n5698), .A3(n5697), .A4(
        n5696), .ZN(n5699) );
  NAND4_X1 U6878 ( .A1(n5702), .A2(n5701), .A3(n5700), .A4(n5699), .ZN(n5713)
         );
  INV_X1 U6879 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6757) );
  NAND4_X1 U6880 ( .A1(EAX_REG_5__SCAN_IN), .A2(INSTQUEUE_REG_8__3__SCAN_IN), 
        .A3(REIP_REG_28__SCAN_IN), .A4(n6757), .ZN(n5712) );
  NAND4_X1 U6881 ( .A1(EAX_REG_10__SCAN_IN), .A2(INSTQUEUE_REG_5__7__SCAN_IN), 
        .A3(FLUSH_REG_SCAN_IN), .A4(n4542), .ZN(n5711) );
  INV_X1 U6882 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n5705) );
  INV_X1 U6883 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5755) );
  NAND4_X1 U6884 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(
        BYTEENABLE_REG_2__SCAN_IN), .A3(n5755), .A4(n6348), .ZN(n5704) );
  INV_X1 U6885 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n5748) );
  NAND4_X1 U6886 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTQUEUE_REG_9__3__SCAN_IN), .A3(EAX_REG_3__SCAN_IN), .A4(n5748), 
        .ZN(n5703) );
  OR4_X1 U6887 ( .A1(n5705), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .A3(n5704), 
        .A4(n5703), .ZN(n5709) );
  NAND4_X1 U6888 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        REIP_REG_13__SCAN_IN), .A3(ADDRESS_REG_27__SCAN_IN), .A4(n5939), .ZN(
        n5708) );
  INV_X1 U6889 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6370) );
  NAND4_X1 U6890 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(DATAI_21_), .A3(n5650), .A4(n6370), .ZN(n5707) );
  OR4_X1 U6891 ( .A1(n5709), .A2(n5708), .A3(n5707), .A4(n5706), .ZN(n5710) );
  NOR4_X1 U6892 ( .A1(n5713), .A2(n5712), .A3(n5711), .A4(n5710), .ZN(n5779)
         );
  INV_X1 U6893 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5715) );
  AOI22_X1 U6894 ( .A1(n5715), .A2(keyinput43), .B1(keyinput36), .B2(n6387), 
        .ZN(n5714) );
  OAI221_X1 U6895 ( .B1(n5715), .B2(keyinput43), .C1(n6387), .C2(keyinput36), 
        .A(n5714), .ZN(n5724) );
  AOI22_X1 U6896 ( .A1(n3881), .A2(keyinput25), .B1(keyinput21), .B2(n5650), 
        .ZN(n5716) );
  OAI221_X1 U6897 ( .B1(n3881), .B2(keyinput25), .C1(n5650), .C2(keyinput21), 
        .A(n5716), .ZN(n5723) );
  INV_X1 U6898 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6784) );
  AOI22_X1 U6899 ( .A1(n6784), .A2(keyinput2), .B1(keyinput62), .B2(n6348), 
        .ZN(n5717) );
  OAI221_X1 U6900 ( .B1(n6784), .B2(keyinput2), .C1(n6348), .C2(keyinput62), 
        .A(n5717), .ZN(n5722) );
  INV_X1 U6901 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5720) );
  AOI22_X1 U6902 ( .A1(n5720), .A2(keyinput54), .B1(keyinput22), .B2(n5719), 
        .ZN(n5718) );
  OAI221_X1 U6903 ( .B1(n5720), .B2(keyinput54), .C1(n5719), .C2(keyinput22), 
        .A(n5718), .ZN(n5721) );
  NOR4_X1 U6904 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n5777)
         );
  INV_X1 U6905 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n6361) );
  AOI22_X1 U6906 ( .A1(n3025), .A2(keyinput45), .B1(keyinput42), .B2(n6361), 
        .ZN(n5725) );
  OAI221_X1 U6907 ( .B1(n3025), .B2(keyinput45), .C1(n6361), .C2(keyinput42), 
        .A(n5725), .ZN(n5733) );
  INV_X1 U6908 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6177) );
  AOI22_X1 U6909 ( .A1(n5877), .A2(keyinput16), .B1(keyinput33), .B2(n6177), 
        .ZN(n5726) );
  OAI221_X1 U6910 ( .B1(n5877), .B2(keyinput16), .C1(n6177), .C2(keyinput33), 
        .A(n5726), .ZN(n5732) );
  AOI22_X1 U6911 ( .A1(n5728), .A2(keyinput27), .B1(keyinput60), .B2(n5705), 
        .ZN(n5727) );
  OAI221_X1 U6912 ( .B1(n5728), .B2(keyinput27), .C1(n5705), .C2(keyinput60), 
        .A(n5727), .ZN(n5731) );
  AOI22_X1 U6913 ( .A1(n6757), .A2(keyinput18), .B1(n6382), .B2(keyinput5), 
        .ZN(n5729) );
  OAI221_X1 U6914 ( .B1(n6757), .B2(keyinput18), .C1(n6382), .C2(keyinput5), 
        .A(n5729), .ZN(n5730) );
  NOR4_X1 U6915 ( .A1(n5733), .A2(n5732), .A3(n5731), .A4(n5730), .ZN(n5776)
         );
  AOI22_X1 U6916 ( .A1(n6370), .A2(keyinput4), .B1(n4542), .B2(keyinput23), 
        .ZN(n5734) );
  OAI221_X1 U6917 ( .B1(n6370), .B2(keyinput4), .C1(n4542), .C2(keyinput23), 
        .A(n5734), .ZN(n5744) );
  AOI22_X1 U6918 ( .A1(n5737), .A2(keyinput44), .B1(n5736), .B2(keyinput50), 
        .ZN(n5735) );
  OAI221_X1 U6919 ( .B1(n5737), .B2(keyinput44), .C1(n5736), .C2(keyinput50), 
        .A(n5735), .ZN(n5743) );
  AOI22_X1 U6920 ( .A1(n4569), .A2(keyinput19), .B1(n6374), .B2(keyinput24), 
        .ZN(n5738) );
  OAI221_X1 U6921 ( .B1(n4569), .B2(keyinput19), .C1(n6374), .C2(keyinput24), 
        .A(n5738), .ZN(n5742) );
  INV_X1 U6922 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6758) );
  INV_X1 U6923 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5740) );
  AOI22_X1 U6924 ( .A1(n6758), .A2(keyinput8), .B1(n5740), .B2(keyinput51), 
        .ZN(n5739) );
  OAI221_X1 U6925 ( .B1(n6758), .B2(keyinput8), .C1(n5740), .C2(keyinput51), 
        .A(n5739), .ZN(n5741) );
  NOR4_X1 U6926 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n5741), .ZN(n5775)
         );
  AOI22_X1 U6927 ( .A1(n5746), .A2(keyinput47), .B1(n5997), .B2(keyinput6), 
        .ZN(n5745) );
  OAI221_X1 U6928 ( .B1(n5746), .B2(keyinput47), .C1(n5997), .C2(keyinput6), 
        .A(n5745), .ZN(n5747) );
  INV_X1 U6929 ( .A(n5747), .ZN(n5763) );
  XNOR2_X1 U6930 ( .A(keyinput56), .B(n5748), .ZN(n5750) );
  XNOR2_X1 U6931 ( .A(keyinput26), .B(n3813), .ZN(n5749) );
  NOR2_X1 U6932 ( .A1(n5750), .A2(n5749), .ZN(n5762) );
  XNOR2_X1 U6933 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .B(keyinput30), .ZN(n5754) );
  XNOR2_X1 U6934 ( .A(EBX_REG_24__SCAN_IN), .B(keyinput20), .ZN(n5753) );
  XNOR2_X1 U6935 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput17), .ZN(
        n5752) );
  XNOR2_X1 U6936 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .B(keyinput48), .ZN(n5751)
         );
  NAND4_X1 U6937 ( .A1(n5754), .A2(n5753), .A3(n5752), .A4(n5751), .ZN(n5760)
         );
  XNOR2_X1 U6938 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .B(keyinput32), .ZN(n5758) );
  XNOR2_X1 U6939 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .B(keyinput40), .ZN(n5757) );
  XNOR2_X1 U6940 ( .A(keyinput7), .B(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5756)
         );
  NAND3_X1 U6941 ( .A1(n5758), .A2(n5757), .A3(n5756), .ZN(n5759) );
  NOR2_X1 U6942 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  NAND3_X1 U6943 ( .A1(n5763), .A2(n5762), .A3(n5761), .ZN(n5773) );
  INV_X1 U6944 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5765) );
  AOI22_X1 U6945 ( .A1(n5766), .A2(keyinput37), .B1(n5765), .B2(keyinput28), 
        .ZN(n5764) );
  OAI221_X1 U6946 ( .B1(n5766), .B2(keyinput37), .C1(n5765), .C2(keyinput28), 
        .A(n5764), .ZN(n5772) );
  AOI22_X1 U6947 ( .A1(n5769), .A2(keyinput57), .B1(n5768), .B2(keyinput46), 
        .ZN(n5767) );
  OAI221_X1 U6948 ( .B1(n5769), .B2(keyinput57), .C1(n5768), .C2(keyinput46), 
        .A(n5767), .ZN(n5771) );
  INV_X1 U6949 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6759) );
  XNOR2_X1 U6950 ( .A(n6759), .B(keyinput14), .ZN(n5770) );
  NOR4_X1 U6951 ( .A1(n5773), .A2(n5772), .A3(n5771), .A4(n5770), .ZN(n5774)
         );
  NAND4_X1 U6952 ( .A1(n5777), .A2(n5776), .A3(n5775), .A4(n5774), .ZN(n5778)
         );
  AOI21_X1 U6953 ( .B1(n5780), .B2(n5779), .A(n5778), .ZN(n5822) );
  AOI22_X1 U6954 ( .A1(n6372), .A2(keyinput29), .B1(keyinput9), .B2(n5782), 
        .ZN(n5781) );
  OAI221_X1 U6955 ( .B1(n6372), .B2(keyinput29), .C1(n5782), .C2(keyinput9), 
        .A(n5781), .ZN(n5791) );
  INV_X1 U6956 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5784) );
  AOI22_X1 U6957 ( .A1(n6162), .A2(keyinput38), .B1(n5784), .B2(keyinput12), 
        .ZN(n5783) );
  OAI221_X1 U6958 ( .B1(n6162), .B2(keyinput38), .C1(n5784), .C2(keyinput12), 
        .A(n5783), .ZN(n5790) );
  AOI22_X1 U6959 ( .A1(n5939), .A2(keyinput53), .B1(keyinput52), .B2(n6104), 
        .ZN(n5785) );
  OAI221_X1 U6960 ( .B1(n5939), .B2(keyinput53), .C1(n6104), .C2(keyinput52), 
        .A(n5785), .ZN(n5789) );
  AOI22_X1 U6961 ( .A1(n5787), .A2(keyinput39), .B1(n6780), .B2(keyinput61), 
        .ZN(n5786) );
  OAI221_X1 U6962 ( .B1(n5787), .B2(keyinput39), .C1(n6780), .C2(keyinput61), 
        .A(n5786), .ZN(n5788) );
  NOR4_X1 U6963 ( .A1(n5791), .A2(n5790), .A3(n5789), .A4(n5788), .ZN(n5821)
         );
  INV_X1 U6964 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5794) );
  AOI22_X1 U6965 ( .A1(n5794), .A2(keyinput13), .B1(keyinput59), .B2(n5793), 
        .ZN(n5792) );
  OAI221_X1 U6966 ( .B1(n5794), .B2(keyinput13), .C1(n5793), .C2(keyinput59), 
        .A(n5792), .ZN(n5805) );
  INV_X1 U6967 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6295) );
  AOI22_X1 U6968 ( .A1(n6295), .A2(keyinput15), .B1(n5796), .B2(keyinput31), 
        .ZN(n5795) );
  OAI221_X1 U6969 ( .B1(n6295), .B2(keyinput15), .C1(n5796), .C2(keyinput31), 
        .A(n5795), .ZN(n5804) );
  AOI22_X1 U6970 ( .A1(n5799), .A2(keyinput11), .B1(keyinput41), .B2(n5798), 
        .ZN(n5797) );
  OAI221_X1 U6971 ( .B1(n5799), .B2(keyinput11), .C1(n5798), .C2(keyinput41), 
        .A(n5797), .ZN(n5803) );
  AOI22_X1 U6972 ( .A1(n5801), .A2(keyinput63), .B1(n3677), .B2(keyinput58), 
        .ZN(n5800) );
  OAI221_X1 U6973 ( .B1(n5801), .B2(keyinput63), .C1(n3677), .C2(keyinput58), 
        .A(n5800), .ZN(n5802) );
  NOR4_X1 U6974 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n5820)
         );
  INV_X1 U6975 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6358) );
  AOI22_X1 U6976 ( .A1(n5807), .A2(keyinput3), .B1(keyinput34), .B2(n6358), 
        .ZN(n5806) );
  OAI221_X1 U6977 ( .B1(n5807), .B2(keyinput3), .C1(n6358), .C2(keyinput34), 
        .A(n5806), .ZN(n5818) );
  AOI22_X1 U6978 ( .A1(n5810), .A2(keyinput0), .B1(keyinput35), .B2(n5809), 
        .ZN(n5808) );
  OAI221_X1 U6979 ( .B1(n5810), .B2(keyinput0), .C1(n5809), .C2(keyinput35), 
        .A(n5808), .ZN(n5817) );
  INV_X1 U6980 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n6356) );
  AOI22_X1 U6981 ( .A1(n6356), .A2(keyinput55), .B1(keyinput49), .B2(n5812), 
        .ZN(n5811) );
  OAI221_X1 U6982 ( .B1(n6356), .B2(keyinput55), .C1(n5812), .C2(keyinput49), 
        .A(n5811), .ZN(n5816) );
  INV_X1 U6983 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n5814) );
  AOI22_X1 U6984 ( .A1(n4530), .A2(keyinput10), .B1(keyinput1), .B2(n5814), 
        .ZN(n5813) );
  OAI221_X1 U6985 ( .B1(n4530), .B2(keyinput10), .C1(n5814), .C2(keyinput1), 
        .A(n5813), .ZN(n5815) );
  NOR4_X1 U6986 ( .A1(n5818), .A2(n5817), .A3(n5816), .A4(n5815), .ZN(n5819)
         );
  NAND4_X1 U6987 ( .A1(n5822), .A2(n5821), .A3(n5820), .A4(n5819), .ZN(n5830)
         );
  OAI21_X1 U6988 ( .B1(n5825), .B2(n5824), .A(n5823), .ZN(n6073) );
  NAND2_X1 U6989 ( .A1(n6490), .A2(REIP_REG_14__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U6990 ( .A1(n6450), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5826)
         );
  OAI211_X1 U6991 ( .C1(n6461), .C2(n6221), .A(n6085), .B(n5826), .ZN(n5828)
         );
  NOR2_X1 U6992 ( .A1(n6222), .A2(n5886), .ZN(n5827) );
  AOI211_X1 U6993 ( .C1(n6455), .C2(n6073), .A(n5828), .B(n5827), .ZN(n5829)
         );
  XOR2_X1 U6994 ( .A(n5830), .B(n5829), .Z(U2972) );
  XOR2_X1 U6995 ( .A(n5832), .B(n5831), .Z(n6103) );
  NOR2_X1 U6996 ( .A1(n6120), .A2(n5787), .ZN(n6098) );
  AOI21_X1 U6997 ( .B1(n6450), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6098), 
        .ZN(n5833) );
  OAI21_X1 U6998 ( .B1(n6230), .B2(n6461), .A(n5833), .ZN(n5834) );
  AOI21_X1 U6999 ( .B1(n6327), .B2(n6456), .A(n5834), .ZN(n5835) );
  OAI21_X1 U7000 ( .B1(n6103), .B2(n6161), .A(n5835), .ZN(U2973) );
  INV_X1 U7001 ( .A(n5836), .ZN(n5867) );
  AOI21_X1 U7002 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5610), .A(n5867), 
        .ZN(n5853) );
  NOR2_X1 U7003 ( .A1(n5610), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5854)
         );
  NOR2_X1 U7004 ( .A1(n5853), .A2(n5854), .ZN(n5852) );
  NOR2_X1 U7005 ( .A1(n3093), .A2(n5837), .ZN(n5856) );
  NOR2_X1 U7006 ( .A1(n5852), .A2(n5856), .ZN(n5848) );
  NOR2_X1 U7007 ( .A1(n5610), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5846)
         );
  NAND2_X1 U7008 ( .A1(n5610), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5844) );
  OAI21_X1 U7009 ( .B1(n5848), .B2(n5846), .A(n5844), .ZN(n5839) );
  XNOR2_X1 U7010 ( .A(n3093), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5838)
         );
  XNOR2_X1 U7011 ( .A(n5839), .B(n5838), .ZN(n6113) );
  INV_X1 U7012 ( .A(n6242), .ZN(n5841) );
  NAND2_X1 U7013 ( .A1(n6490), .A2(REIP_REG_12__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7014 ( .A1(n6450), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5840)
         );
  OAI211_X1 U7015 ( .C1(n6461), .C2(n5841), .A(n6105), .B(n5840), .ZN(n5842)
         );
  AOI21_X1 U7016 ( .B1(n6352), .B2(n6456), .A(n5842), .ZN(n5843) );
  OAI21_X1 U7017 ( .B1(n6113), .B2(n6161), .A(n5843), .ZN(U2974) );
  INV_X1 U7018 ( .A(n5844), .ZN(n5845) );
  NOR2_X1 U7019 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  XNOR2_X1 U7020 ( .A(n5848), .B(n5847), .ZN(n6465) );
  NAND2_X1 U7021 ( .A1(n6465), .A2(n6455), .ZN(n5851) );
  AND2_X1 U7022 ( .A1(n6490), .A2(REIP_REG_11__SCAN_IN), .ZN(n6462) );
  NOR2_X1 U7023 ( .A1(n6461), .A2(n6252), .ZN(n5849) );
  AOI211_X1 U7024 ( .C1(n6450), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6462), 
        .B(n5849), .ZN(n5850) );
  OAI211_X1 U7025 ( .C1(n5886), .C2(n6251), .A(n5851), .B(n5850), .ZN(U2975)
         );
  INV_X1 U7026 ( .A(n5852), .ZN(n5857) );
  OAI21_X1 U7027 ( .B1(n5856), .B2(n5854), .A(n5853), .ZN(n5855) );
  OAI21_X1 U7028 ( .B1(n5857), .B2(n5856), .A(n5855), .ZN(n6129) );
  AOI22_X1 U7029 ( .A1(n6450), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6490), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5858) );
  OAI21_X1 U7030 ( .B1(n6461), .B2(n5859), .A(n5858), .ZN(n5860) );
  AOI21_X1 U7031 ( .B1(n6265), .B2(n6456), .A(n5860), .ZN(n5861) );
  OAI21_X1 U7032 ( .B1(n6129), .B2(n6161), .A(n5861), .ZN(U2976) );
  INV_X1 U7033 ( .A(n5862), .ZN(n5864) );
  NOR2_X1 U7034 ( .A1(n5864), .A2(n5863), .ZN(n5868) );
  NAND2_X1 U7035 ( .A1(n6425), .A2(n5865), .ZN(n5876) );
  XNOR2_X1 U7036 ( .A(n5866), .B(n6487), .ZN(n5875) );
  NAND2_X1 U7037 ( .A1(n5876), .A2(n5875), .ZN(n5874) );
  AOI21_X1 U7038 ( .B1(n5868), .B2(n5874), .A(n5867), .ZN(n6474) );
  NAND2_X1 U7039 ( .A1(n6474), .A2(n6455), .ZN(n5872) );
  AND2_X1 U7040 ( .A1(n6490), .A2(REIP_REG_9__SCAN_IN), .ZN(n6471) );
  NOR2_X1 U7041 ( .A1(n6461), .A2(n5869), .ZN(n5870) );
  AOI211_X1 U7042 ( .C1(n6450), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6471), 
        .B(n5870), .ZN(n5871) );
  OAI211_X1 U7043 ( .C1(n5886), .C2(n5873), .A(n5872), .B(n5871), .ZN(U2977)
         );
  OAI21_X1 U7044 ( .B1(n5876), .B2(n5875), .A(n5874), .ZN(n6484) );
  OR2_X1 U7045 ( .A1(n6484), .A2(n6161), .ZN(n5884) );
  INV_X1 U7046 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5878) );
  OAI22_X1 U7047 ( .A1(n5879), .A2(n5878), .B1(n6120), .B2(n5877), .ZN(n5880)
         );
  AOI21_X1 U7048 ( .B1(n5882), .B2(n5881), .A(n5880), .ZN(n5883) );
  OAI211_X1 U7049 ( .C1(n5886), .C2(n5885), .A(n5884), .B(n5883), .ZN(U2978)
         );
  INV_X1 U7050 ( .A(n5887), .ZN(n5920) );
  INV_X1 U7051 ( .A(n5913), .ZN(n5905) );
  INV_X1 U7052 ( .A(n5912), .ZN(n5904) );
  NAND2_X1 U7053 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7054 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5892) );
  NOR3_X1 U7055 ( .A1(n6512), .A2(n6511), .A3(n5892), .ZN(n6115) );
  NAND2_X1 U7056 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7057 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6124) );
  NOR2_X1 U7058 ( .A1(n6123), .A2(n6124), .ZN(n5893) );
  NAND2_X1 U7059 ( .A1(n6115), .A2(n5893), .ZN(n6095) );
  INV_X1 U7060 ( .A(n6095), .ZN(n5888) );
  OR2_X1 U7061 ( .A1(n6116), .A2(n5888), .ZN(n5889) );
  NAND2_X1 U7062 ( .A1(n5889), .A2(n6114), .ZN(n6053) );
  NAND2_X1 U7063 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6076) );
  NOR2_X1 U7064 ( .A1(n6076), .A2(n6077), .ZN(n6084) );
  NAND2_X1 U7065 ( .A1(n6084), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5907) );
  NOR3_X1 U7066 ( .A1(n6068), .A2(n6063), .A3(n5907), .ZN(n5894) );
  NOR2_X1 U7067 ( .A1(n6116), .A2(n5894), .ZN(n5890) );
  NOR2_X1 U7068 ( .A1(n6053), .A2(n5890), .ZN(n6014) );
  NAND2_X1 U7069 ( .A1(n5891), .A2(n6522), .ZN(n6501) );
  NOR2_X1 U7070 ( .A1(n5892), .A2(n6501), .ZN(n6122) );
  NAND2_X1 U7071 ( .A1(n5893), .A2(n6122), .ZN(n6054) );
  INV_X1 U7072 ( .A(n5894), .ZN(n5895) );
  NOR2_X1 U7073 ( .A1(n6054), .A2(n5895), .ZN(n6011) );
  INV_X1 U7074 ( .A(n5896), .ZN(n6016) );
  NAND3_X1 U7075 ( .A1(n6011), .A2(n6016), .A3(n6021), .ZN(n5897) );
  NAND2_X1 U7076 ( .A1(n6496), .A2(n5897), .ZN(n5898) );
  AND2_X1 U7077 ( .A1(n6014), .A2(n5898), .ZN(n6002) );
  INV_X1 U7078 ( .A(n5899), .ZN(n5900) );
  NAND2_X1 U7079 ( .A1(n6496), .A2(n5900), .ZN(n5901) );
  AND2_X1 U7080 ( .A1(n6002), .A2(n5901), .ZN(n5986) );
  NAND2_X1 U7081 ( .A1(n6539), .A2(n6531), .ZN(n5902) );
  NAND2_X1 U7082 ( .A1(n5902), .A2(n5910), .ZN(n5903) );
  NAND2_X1 U7083 ( .A1(n5986), .A2(n5903), .ZN(n5980) );
  AOI21_X1 U7084 ( .B1(n5960), .B2(n6496), .A(n5980), .ZN(n5949) );
  OAI21_X1 U7085 ( .B1(n5904), .B2(n6119), .A(n5949), .ZN(n5929) );
  AOI21_X1 U7086 ( .B1(n5905), .B2(n6496), .A(n5929), .ZN(n5927) );
  INV_X1 U7087 ( .A(n6054), .ZN(n5906) );
  NAND2_X1 U7088 ( .A1(n6508), .A2(n5906), .ZN(n6079) );
  INV_X1 U7089 ( .A(n5907), .ZN(n6055) );
  NAND2_X1 U7090 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5908) );
  INV_X1 U7091 ( .A(n5910), .ZN(n5911) );
  NAND2_X1 U7092 ( .A1(n5990), .A2(n5911), .ZN(n5973) );
  NAND3_X1 U7093 ( .A1(n5935), .A2(n5913), .A3(n5916), .ZN(n5914) );
  OAI211_X1 U7094 ( .C1(n5927), .C2(n5916), .A(n5915), .B(n5914), .ZN(n5917)
         );
  AOI21_X1 U7095 ( .B1(n6534), .B2(n5918), .A(n5917), .ZN(n5919) );
  OAI21_X1 U7096 ( .B1(n5920), .B2(n6483), .A(n5919), .ZN(U2987) );
  AOI21_X1 U7097 ( .B1(n5935), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7098 ( .A1(n5921), .A2(n6537), .ZN(n5926) );
  INV_X1 U7099 ( .A(n5922), .ZN(n5924) );
  AOI21_X1 U7100 ( .B1(n5924), .B2(n6534), .A(n5923), .ZN(n5925) );
  OAI211_X1 U7101 ( .C1(n5928), .C2(n5927), .A(n5926), .B(n5925), .ZN(U2988)
         );
  INV_X1 U7102 ( .A(n5472), .ZN(n5932) );
  NAND2_X1 U7103 ( .A1(n5929), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5930) );
  OAI211_X1 U7104 ( .C1(n5932), .C2(n6121), .A(n5931), .B(n5930), .ZN(n5933)
         );
  AOI21_X1 U7105 ( .B1(n5935), .B2(n5934), .A(n5933), .ZN(n5936) );
  OAI21_X1 U7106 ( .B1(n5937), .B2(n6483), .A(n5936), .ZN(U2989) );
  XNOR2_X1 U7107 ( .A(n5939), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5944)
         );
  INV_X1 U7108 ( .A(n5938), .ZN(n5953) );
  NOR2_X1 U7109 ( .A1(n5949), .A2(n5939), .ZN(n5943) );
  OAI21_X1 U7110 ( .B1(n5941), .B2(n6121), .A(n5940), .ZN(n5942) );
  AOI211_X1 U7111 ( .C1(n5944), .C2(n5953), .A(n5943), .B(n5942), .ZN(n5945)
         );
  OAI21_X1 U7112 ( .B1(n5946), .B2(n6483), .A(n5945), .ZN(U2990) );
  OAI21_X1 U7113 ( .B1(n5948), .B2(n6121), .A(n5947), .ZN(n5951) );
  NOR2_X1 U7114 ( .A1(n5949), .A2(n5952), .ZN(n5950) );
  AOI211_X1 U7115 ( .C1(n5953), .C2(n5952), .A(n5951), .B(n5950), .ZN(n5954)
         );
  OAI21_X1 U7116 ( .B1(n5955), .B2(n6483), .A(n5954), .ZN(U2991) );
  INV_X1 U7117 ( .A(n5956), .ZN(n5966) );
  INV_X1 U7118 ( .A(n5957), .ZN(n5958) );
  OAI21_X1 U7119 ( .B1(n5959), .B2(n6121), .A(n5958), .ZN(n5964) );
  INV_X1 U7120 ( .A(n5960), .ZN(n5961) );
  AOI211_X1 U7121 ( .C1(n3080), .C2(n5962), .A(n5961), .B(n5973), .ZN(n5963)
         );
  AOI211_X1 U7122 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5980), .A(n5964), .B(n5963), .ZN(n5965) );
  OAI21_X1 U7123 ( .B1(n5966), .B2(n6483), .A(n5965), .ZN(U2992) );
  NAND2_X1 U7124 ( .A1(n5967), .A2(n6537), .ZN(n5972) );
  OAI21_X1 U7125 ( .B1(n5969), .B2(n6121), .A(n5968), .ZN(n5970) );
  AOI21_X1 U7126 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5980), .A(n5970), 
        .ZN(n5971) );
  OAI211_X1 U7127 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5973), .A(n5972), .B(n5971), .ZN(U2993) );
  INV_X1 U7128 ( .A(n5974), .ZN(n5977) );
  INV_X1 U7129 ( .A(n5975), .ZN(n5976) );
  AOI21_X1 U7130 ( .B1(n5977), .B2(n6534), .A(n5976), .ZN(n5982) );
  INV_X1 U7131 ( .A(n5978), .ZN(n5979) );
  OAI211_X1 U7132 ( .C1(n5990), .C2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n5980), .B(n5979), .ZN(n5981) );
  OAI211_X1 U7133 ( .C1(n5983), .C2(n6483), .A(n5982), .B(n5981), .ZN(U2994)
         );
  INV_X1 U7134 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5989) );
  OAI21_X1 U7135 ( .B1(n5985), .B2(n6121), .A(n5984), .ZN(n5988) );
  NOR2_X1 U7136 ( .A1(n5986), .A2(n5989), .ZN(n5987) );
  AOI211_X1 U7137 ( .C1(n5990), .C2(n5989), .A(n5988), .B(n5987), .ZN(n5991)
         );
  OAI21_X1 U7138 ( .B1(n5992), .B2(n6483), .A(n5991), .ZN(U2995) );
  AND2_X1 U7139 ( .A1(n6033), .A2(n6021), .ZN(n6008) );
  XNOR2_X1 U7140 ( .A(n6007), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5999)
         );
  INV_X1 U7141 ( .A(n5993), .ZN(n5995) );
  AOI21_X1 U7142 ( .B1(n5995), .B2(n6534), .A(n5994), .ZN(n5996) );
  OAI21_X1 U7143 ( .B1(n6002), .B2(n5997), .A(n5996), .ZN(n5998) );
  AOI21_X1 U7144 ( .B1(n6008), .B2(n5999), .A(n5998), .ZN(n6000) );
  OAI21_X1 U7145 ( .B1(n6001), .B2(n6483), .A(n6000), .ZN(U2996) );
  NOR2_X1 U7146 ( .A1(n6002), .A2(n6007), .ZN(n6006) );
  OAI21_X1 U7147 ( .B1(n6004), .B2(n6121), .A(n6003), .ZN(n6005) );
  AOI211_X1 U7148 ( .C1(n6008), .C2(n6007), .A(n6006), .B(n6005), .ZN(n6009)
         );
  OAI21_X1 U7149 ( .B1(n6010), .B2(n6483), .A(n6009), .ZN(U2997) );
  AOI21_X1 U7150 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6011), .A(n6531), 
        .ZN(n6012) );
  INV_X1 U7151 ( .A(n6012), .ZN(n6013) );
  AND2_X1 U7152 ( .A1(n6014), .A2(n6013), .ZN(n6046) );
  NAND2_X1 U7153 ( .A1(n6508), .A2(n6040), .ZN(n6015) );
  OAI21_X1 U7154 ( .B1(n6116), .B2(n6016), .A(n6015), .ZN(n6017) );
  INV_X1 U7155 ( .A(n6017), .ZN(n6018) );
  NAND2_X1 U7156 ( .A1(n6046), .A2(n6018), .ZN(n6031) );
  OAI21_X1 U7157 ( .B1(n6020), .B2(n6121), .A(n6019), .ZN(n6025) );
  INV_X1 U7158 ( .A(n6033), .ZN(n6023) );
  NOR3_X1 U7159 ( .A1(n6023), .A2(n6022), .A3(n6021), .ZN(n6024) );
  AOI211_X1 U7160 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n6031), .A(n6025), .B(n6024), .ZN(n6026) );
  OAI21_X1 U7161 ( .B1(n6027), .B2(n6483), .A(n6026), .ZN(U2998) );
  NAND2_X1 U7162 ( .A1(n6143), .A2(n6534), .ZN(n6029) );
  NAND2_X1 U7163 ( .A1(n6029), .A2(n6028), .ZN(n6030) );
  AOI21_X1 U7164 ( .B1(n6031), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6030), 
        .ZN(n6035) );
  NAND2_X1 U7165 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  OAI211_X1 U7166 ( .C1(n6036), .C2(n6483), .A(n6035), .B(n6034), .ZN(U2999)
         );
  OAI21_X1 U7167 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6539), .A(n6046), 
        .ZN(n6039) );
  OAI21_X1 U7168 ( .B1(n6121), .B2(n6189), .A(n6037), .ZN(n6038) );
  AOI21_X1 U7169 ( .B1(n6039), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n6038), 
        .ZN(n6042) );
  NAND3_X1 U7170 ( .A1(n6050), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n6040), .ZN(n6041) );
  OAI211_X1 U7171 ( .C1(n6043), .C2(n6483), .A(n6042), .B(n6041), .ZN(U3000)
         );
  OAI21_X1 U7172 ( .B1(n6121), .B2(n6045), .A(n6044), .ZN(n6048) );
  NOR2_X1 U7173 ( .A1(n6046), .A2(n6049), .ZN(n6047) );
  AOI211_X1 U7174 ( .C1(n6050), .C2(n6049), .A(n6048), .B(n6047), .ZN(n6051)
         );
  OAI21_X1 U7175 ( .B1(n6052), .B2(n6483), .A(n6051), .ZN(U3001) );
  INV_X1 U7176 ( .A(n6067), .ZN(n6057) );
  AOI21_X1 U7177 ( .B1(n6054), .B2(n6508), .A(n6053), .ZN(n6469) );
  OAI21_X1 U7178 ( .B1(n6055), .B2(n6119), .A(n6469), .ZN(n6056) );
  AOI21_X1 U7179 ( .B1(n6057), .B2(n6068), .A(n6056), .ZN(n6066) );
  NAND2_X1 U7180 ( .A1(n6058), .A2(n6537), .ZN(n6062) );
  NOR3_X1 U7181 ( .A1(n6067), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6068), 
        .ZN(n6059) );
  AOI211_X1 U7182 ( .C1(n6534), .C2(n6196), .A(n6060), .B(n6059), .ZN(n6061)
         );
  OAI211_X1 U7183 ( .C1(n6066), .C2(n6063), .A(n6062), .B(n6061), .ZN(U3002)
         );
  AND2_X1 U7184 ( .A1(n5506), .A2(n6064), .ZN(n6065) );
  AOI21_X1 U7185 ( .B1(n6068), .B2(n6067), .A(n6066), .ZN(n6069) );
  AOI211_X1 U7186 ( .C1(n6534), .C2(n3135), .A(n6070), .B(n6069), .ZN(n6071)
         );
  OAI21_X1 U7187 ( .B1(n6072), .B2(n6483), .A(n6071), .ZN(U3003) );
  INV_X1 U7188 ( .A(n6073), .ZN(n6089) );
  INV_X1 U7189 ( .A(n6469), .ZN(n6110) );
  OR3_X1 U7190 ( .A1(n6075), .A2(n6074), .A3(n6095), .ZN(n6078) );
  INV_X1 U7191 ( .A(n6076), .ZN(n6080) );
  NAND2_X1 U7192 ( .A1(n6080), .A2(n6077), .ZN(n6094) );
  AOI21_X1 U7193 ( .B1(n6079), .B2(n6078), .A(n6094), .ZN(n6100) );
  OAI22_X1 U7194 ( .A1(n6081), .A2(n6080), .B1(n6084), .B2(n6096), .ZN(n6082)
         );
  INV_X1 U7195 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6083) );
  NAND3_X1 U7196 ( .A1(n6464), .A2(n6084), .A3(n6083), .ZN(n6086) );
  OAI211_X1 U7197 ( .C1(n6121), .C2(n6219), .A(n6086), .B(n6085), .ZN(n6087)
         );
  AOI21_X1 U7198 ( .B1(n6099), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n6087), 
        .ZN(n6088) );
  OAI21_X1 U7199 ( .B1(n6089), .B2(n6483), .A(n6088), .ZN(U3004) );
  INV_X1 U7200 ( .A(n6090), .ZN(n6093) );
  INV_X1 U7201 ( .A(n6091), .ZN(n6092) );
  AOI21_X1 U7202 ( .B1(n6093), .B2(n6092), .A(n5507), .ZN(n6326) );
  NOR3_X1 U7203 ( .A1(n6096), .A2(n6095), .A3(n6094), .ZN(n6097) );
  AOI211_X1 U7204 ( .C1(n6534), .C2(n6326), .A(n6098), .B(n6097), .ZN(n6102)
         );
  OAI21_X1 U7205 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6100), .A(n6099), 
        .ZN(n6101) );
  OAI211_X1 U7206 ( .C1(n6103), .C2(n6483), .A(n6102), .B(n6101), .ZN(U3005)
         );
  NAND3_X1 U7207 ( .A1(n6464), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n6104), .ZN(n6106) );
  OAI211_X1 U7208 ( .C1(n6121), .C2(n6238), .A(n6106), .B(n6105), .ZN(n6107)
         );
  INV_X1 U7209 ( .A(n6107), .ZN(n6112) );
  AOI21_X1 U7210 ( .B1(n6108), .B2(n6531), .A(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n6109) );
  OAI21_X1 U7211 ( .B1(n6110), .B2(n6109), .A(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n6111) );
  OAI211_X1 U7212 ( .C1(n6113), .C2(n6483), .A(n6112), .B(n6111), .ZN(U3006)
         );
  INV_X1 U7213 ( .A(n6123), .ZN(n6479) );
  INV_X1 U7214 ( .A(n6114), .ZN(n6118) );
  OAI22_X1 U7215 ( .A1(n6116), .A2(n6115), .B1(n6122), .B2(n6531), .ZN(n6117)
         );
  NOR2_X1 U7216 ( .A1(n6118), .A2(n6117), .ZN(n6492) );
  OAI21_X1 U7217 ( .B1(n6479), .B2(n6119), .A(n6492), .ZN(n6470) );
  OAI22_X1 U7218 ( .A1(n6121), .A2(n6261), .B1(n6270), .B2(n6120), .ZN(n6127)
         );
  NAND2_X1 U7219 ( .A1(n6122), .A2(n6521), .ZN(n6494) );
  NOR2_X1 U7220 ( .A1(n6123), .A2(n6494), .ZN(n6473) );
  OAI211_X1 U7221 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6473), .B(n6124), .ZN(n6125) );
  INV_X1 U7222 ( .A(n6125), .ZN(n6126) );
  AOI211_X1 U7223 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6470), .A(n6127), .B(n6126), .ZN(n6128) );
  OAI21_X1 U7224 ( .B1(n6129), .B2(n6483), .A(n6128), .ZN(U3008) );
  INV_X1 U7225 ( .A(n6130), .ZN(n6131) );
  OAI22_X1 U7226 ( .A1(n6134), .A2(n6133), .B1(n6132), .B2(n6131), .ZN(n6136)
         );
  MUX2_X1 U7227 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6136), .S(n6135), 
        .Z(U3456) );
  MUX2_X1 U7228 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6137), .Z(U3447) );
  MUX2_X1 U7229 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6137), .Z(U3446) );
  MUX2_X1 U7230 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6137), .Z(U3445) );
  AND2_X1 U7231 ( .A1(n6385), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U7232 ( .B1(n6139), .B2(n6138), .A(n6179), .ZN(n6141) );
  AOI22_X1 U7233 ( .A1(n6142), .A2(n6311), .B1(n6141), .B2(n6140), .ZN(n6147)
         );
  AOI22_X1 U7234 ( .A1(n6303), .A2(EBX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6306), .ZN(n6146) );
  AOI21_X1 U7235 ( .B1(REIP_REG_19__SCAN_IN), .B2(n6183), .A(n6263), .ZN(n6145) );
  AOI22_X1 U7236 ( .A1(n6152), .A2(n6266), .B1(n6305), .B2(n6143), .ZN(n6144)
         );
  NAND4_X1 U7237 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(U2808)
         );
  AOI22_X1 U7238 ( .A1(n6149), .A2(n6351), .B1(n6340), .B2(DATAI_20_), .ZN(
        n6151) );
  AOI22_X1 U7239 ( .A1(n6342), .A2(DATAI_4_), .B1(n6345), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7240 ( .A1(n6151), .A2(n6150), .ZN(U2871) );
  AOI22_X1 U7241 ( .A1(n6152), .A2(n6351), .B1(n6340), .B2(DATAI_19_), .ZN(
        n6154) );
  AOI22_X1 U7242 ( .A1(n6342), .A2(DATAI_3_), .B1(n6345), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7243 ( .A1(n6154), .A2(n6153), .ZN(U2872) );
  OAI21_X1 U7244 ( .B1(n6156), .B2(n6155), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6157) );
  OAI21_X1 U7245 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6158), .A(n6157), .ZN(
        U2790) );
  OAI21_X1 U7246 ( .B1(BS16_N), .B2(n6159), .A(n6765), .ZN(n6763) );
  OAI21_X1 U7247 ( .B1(n6765), .B2(n6160), .A(n6763), .ZN(U2792) );
  OAI21_X1 U7248 ( .B1(n6163), .B2(n6162), .A(n6161), .ZN(U2793) );
  NOR4_X1 U7249 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6167) );
  NOR4_X1 U7250 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n6166) );
  NOR4_X1 U7251 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6165) );
  NOR4_X1 U7252 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6164) );
  NAND4_X1 U7253 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n6173)
         );
  NOR4_X1 U7254 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6171) );
  AOI211_X1 U7255 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_15__SCAN_IN), .B(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6170) );
  NOR4_X1 U7256 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6169)
         );
  NOR4_X1 U7257 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6168) );
  NAND4_X1 U7258 ( .A1(n6171), .A2(n6170), .A3(n6169), .A4(n6168), .ZN(n6172)
         );
  NOR2_X1 U7259 ( .A1(n6173), .A2(n6172), .ZN(n6786) );
  INV_X1 U7260 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6175) );
  NOR3_X1 U7261 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6176) );
  OAI21_X1 U7262 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6176), .A(n6786), .ZN(n6174)
         );
  OAI21_X1 U7263 ( .B1(n6786), .B2(n6175), .A(n6174), .ZN(U2794) );
  INV_X1 U7264 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6764) );
  AOI21_X1 U7265 ( .B1(n6782), .B2(n6764), .A(n6176), .ZN(n6178) );
  INV_X1 U7266 ( .A(n6786), .ZN(n6789) );
  AOI22_X1 U7267 ( .A1(n6786), .A2(n6178), .B1(n6177), .B2(n6789), .ZN(U2795)
         );
  OAI21_X1 U7268 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6179), .A(n6308), .ZN(n6182) );
  INV_X1 U7269 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6180) );
  NOR2_X1 U7270 ( .A1(n6294), .A2(n6180), .ZN(n6181) );
  AOI211_X1 U7271 ( .C1(EBX_REG_18__SCAN_IN), .C2(n6303), .A(n6182), .B(n6181), 
        .ZN(n6185) );
  NAND2_X1 U7272 ( .A1(n6183), .A2(REIP_REG_18__SCAN_IN), .ZN(n6184) );
  OAI211_X1 U7273 ( .C1(n6299), .C2(n6186), .A(n6185), .B(n6184), .ZN(n6187)
         );
  AOI21_X1 U7274 ( .B1(n6336), .B2(n6266), .A(n6187), .ZN(n6188) );
  OAI21_X1 U7275 ( .B1(n6260), .B2(n6189), .A(n6188), .ZN(U2809) );
  NAND2_X1 U7276 ( .A1(n6191), .A2(n6190), .ZN(n6215) );
  NAND2_X1 U7277 ( .A1(n6192), .A2(n6206), .ZN(n6207) );
  INV_X1 U7278 ( .A(n6193), .ZN(n6201) );
  NAND2_X1 U7279 ( .A1(n6306), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6194)
         );
  NAND2_X1 U7280 ( .A1(n6194), .A2(n6308), .ZN(n6195) );
  AOI21_X1 U7281 ( .B1(n6305), .B2(n6196), .A(n6195), .ZN(n6198) );
  NAND2_X1 U7282 ( .A1(n6229), .A2(EBX_REG_16__SCAN_IN), .ZN(n6197) );
  OAI211_X1 U7283 ( .C1(n6199), .C2(REIP_REG_16__SCAN_IN), .A(n6198), .B(n6197), .ZN(n6200) );
  AOI21_X1 U7284 ( .B1(n6311), .B2(n6201), .A(n6200), .ZN(n6202) );
  OAI21_X1 U7285 ( .B1(n6339), .B2(n6282), .A(n6202), .ZN(n6203) );
  INV_X1 U7286 ( .A(n6203), .ZN(n6204) );
  OAI221_X1 U7287 ( .B1(n6205), .B2(n6215), .C1(n6205), .C2(n6207), .A(n6204), 
        .ZN(U2811) );
  OAI22_X1 U7288 ( .A1(n6259), .A2(n6325), .B1(n6206), .B2(n6215), .ZN(n6210)
         );
  OAI211_X1 U7289 ( .C1(n6294), .C2(n6208), .A(n6308), .B(n6207), .ZN(n6209)
         );
  AOI211_X1 U7290 ( .C1(n6305), .C2(n3135), .A(n6210), .B(n6209), .ZN(n6214)
         );
  INV_X1 U7291 ( .A(n6211), .ZN(n6212) );
  AOI22_X1 U7292 ( .A1(n6346), .A2(n6266), .B1(n6311), .B2(n6212), .ZN(n6213)
         );
  NAND2_X1 U7293 ( .A1(n6214), .A2(n6213), .ZN(U2812) );
  AOI21_X1 U7294 ( .B1(n6217), .B2(n6216), .A(n6215), .ZN(n6218) );
  AOI21_X1 U7295 ( .B1(EBX_REG_14__SCAN_IN), .B2(n6303), .A(n6218), .ZN(n6226)
         );
  INV_X1 U7296 ( .A(n6219), .ZN(n6220) );
  AOI22_X1 U7297 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n6306), .B1(n6305), 
        .B2(n6220), .ZN(n6225) );
  OAI22_X1 U7298 ( .A1(n6222), .A2(n6282), .B1(n6221), .B2(n6299), .ZN(n6223)
         );
  INV_X1 U7299 ( .A(n6223), .ZN(n6224) );
  NAND4_X1 U7300 ( .A1(n6226), .A2(n6225), .A3(n6224), .A4(n6308), .ZN(U2813)
         );
  NOR3_X1 U7301 ( .A1(n6289), .A2(REIP_REG_13__SCAN_IN), .A3(n6227), .ZN(n6228) );
  AOI211_X1 U7302 ( .C1(n6306), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6263), 
        .B(n6228), .ZN(n6237) );
  AOI22_X1 U7303 ( .A1(n6305), .A2(n6326), .B1(n6229), .B2(EBX_REG_13__SCAN_IN), .ZN(n6236) );
  INV_X1 U7304 ( .A(n6230), .ZN(n6231) );
  AOI22_X1 U7305 ( .A1(n6327), .A2(n6266), .B1(n6231), .B2(n6311), .ZN(n6235)
         );
  AOI21_X1 U7306 ( .B1(n6241), .B2(n6233), .A(n6232), .ZN(n6250) );
  NOR2_X1 U7307 ( .A1(n6289), .A2(REIP_REG_12__SCAN_IN), .ZN(n6240) );
  OAI21_X1 U7308 ( .B1(n6250), .B2(n6240), .A(REIP_REG_13__SCAN_IN), .ZN(n6234) );
  NAND4_X1 U7309 ( .A1(n6237), .A2(n6236), .A3(n6235), .A4(n6234), .ZN(U2814)
         );
  INV_X1 U7310 ( .A(n6238), .ZN(n6239) );
  AOI22_X1 U7311 ( .A1(n6305), .A2(n6239), .B1(REIP_REG_12__SCAN_IN), .B2(
        n6250), .ZN(n6246) );
  AOI22_X1 U7312 ( .A1(n6303), .A2(EBX_REG_12__SCAN_IN), .B1(n6306), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6245) );
  AOI21_X1 U7313 ( .B1(n6241), .B2(n6240), .A(n6263), .ZN(n6244) );
  AOI22_X1 U7314 ( .A1(n6352), .A2(n6266), .B1(n6242), .B2(n6311), .ZN(n6243)
         );
  NAND4_X1 U7315 ( .A1(n6246), .A2(n6245), .A3(n6244), .A4(n6243), .ZN(U2815)
         );
  OAI21_X1 U7316 ( .B1(n6289), .B2(n6248), .A(n6247), .ZN(n6249) );
  AOI22_X1 U7317 ( .A1(n6250), .A2(n6249), .B1(EBX_REG_11__SCAN_IN), .B2(n6303), .ZN(n6257) );
  AOI22_X1 U7318 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6306), .B1(n6305), 
        .B2(n6463), .ZN(n6256) );
  INV_X1 U7319 ( .A(n6251), .ZN(n6254) );
  INV_X1 U7320 ( .A(n6252), .ZN(n6253) );
  AOI22_X1 U7321 ( .A1(n6266), .A2(n6254), .B1(n6311), .B2(n6253), .ZN(n6255)
         );
  NAND4_X1 U7322 ( .A1(n6257), .A2(n6256), .A3(n6255), .A4(n6308), .ZN(U2816)
         );
  OAI22_X1 U7323 ( .A1(n6261), .A2(n6260), .B1(n6259), .B2(n6258), .ZN(n6262)
         );
  AOI211_X1 U7324 ( .C1(n6306), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6263), 
        .B(n6262), .ZN(n6274) );
  AOI22_X1 U7325 ( .A1(n6266), .A2(n6265), .B1(n6311), .B2(n6264), .ZN(n6273)
         );
  OAI21_X1 U7326 ( .B1(n6268), .B2(n6267), .A(REIP_REG_10__SCAN_IN), .ZN(n6272) );
  NAND3_X1 U7327 ( .A1(n6319), .A2(n6270), .A3(n6269), .ZN(n6271) );
  NAND4_X1 U7328 ( .A1(n6274), .A2(n6273), .A3(n6272), .A4(n6271), .ZN(U2817)
         );
  INV_X1 U7329 ( .A(n6275), .ZN(n6276) );
  NAND2_X1 U7330 ( .A1(n4209), .A2(n6276), .ZN(n6278) );
  NAND2_X1 U7331 ( .A1(n6306), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6277)
         );
  OAI211_X1 U7332 ( .C1(n6289), .C2(n6278), .A(n6308), .B(n6277), .ZN(n6279)
         );
  AOI21_X1 U7333 ( .B1(n6305), .B2(n6488), .A(n6279), .ZN(n6281) );
  NAND2_X1 U7334 ( .A1(n6229), .A2(EBX_REG_7__SCAN_IN), .ZN(n6280) );
  OAI211_X1 U7335 ( .C1(n6282), .C2(n6429), .A(n6281), .B(n6280), .ZN(n6283)
         );
  INV_X1 U7336 ( .A(n6283), .ZN(n6286) );
  OAI21_X1 U7337 ( .B1(n6291), .B2(n6284), .A(REIP_REG_7__SCAN_IN), .ZN(n6285)
         );
  OAI211_X1 U7338 ( .C1(n6299), .C2(n6433), .A(n6286), .B(n6285), .ZN(U2820)
         );
  OAI21_X1 U7339 ( .B1(n6289), .B2(n6288), .A(n6287), .ZN(n6290) );
  AOI22_X1 U7340 ( .A1(n6291), .A2(n6290), .B1(n6303), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n6298) );
  INV_X1 U7341 ( .A(n6292), .ZN(n6314) );
  NAND2_X1 U7342 ( .A1(n6305), .A2(n6510), .ZN(n6293) );
  OAI211_X1 U7343 ( .C1(n6295), .C2(n6294), .A(n6293), .B(n6308), .ZN(n6296)
         );
  AOI21_X1 U7344 ( .B1(n6314), .B2(n6437), .A(n6296), .ZN(n6297) );
  OAI211_X1 U7345 ( .C1(n6440), .C2(n6299), .A(n6298), .B(n6297), .ZN(U2822)
         );
  AOI22_X1 U7346 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6302), .B1(n6301), .B2(n6300), .ZN(n6323) );
  NAND2_X1 U7347 ( .A1(n6303), .A2(EBX_REG_4__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7348 ( .A1(n6305), .A2(n6304), .ZN(n6309) );
  NAND2_X1 U7349 ( .A1(n6306), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6307)
         );
  AND4_X1 U7350 ( .A1(n6310), .A2(n6309), .A3(n6308), .A4(n6307), .ZN(n6322)
         );
  AOI22_X1 U7351 ( .A1(n6314), .A2(n6313), .B1(n6312), .B2(n6311), .ZN(n6321)
         );
  NOR2_X1 U7352 ( .A1(n6316), .A2(n6315), .ZN(n6317) );
  NAND3_X1 U7353 ( .A1(n6319), .A2(n6318), .A3(n6317), .ZN(n6320) );
  NAND4_X1 U7354 ( .A1(n6323), .A2(n6322), .A3(n6321), .A4(n6320), .ZN(U2823)
         );
  AOI22_X1 U7355 ( .A1(n6346), .A2(n6332), .B1(n6331), .B2(n3135), .ZN(n6324)
         );
  OAI21_X1 U7356 ( .B1(n6335), .B2(n6325), .A(n6324), .ZN(U2844) );
  AOI22_X1 U7357 ( .A1(n6327), .A2(n6332), .B1(n6331), .B2(n6326), .ZN(n6328)
         );
  OAI21_X1 U7358 ( .B1(n6335), .B2(n6329), .A(n6328), .ZN(U2846) );
  INV_X1 U7359 ( .A(n6330), .ZN(n6445) );
  AOI22_X1 U7360 ( .A1(n6445), .A2(n6332), .B1(n6331), .B2(n6520), .ZN(n6333)
         );
  OAI21_X1 U7361 ( .B1(n6335), .B2(n6334), .A(n6333), .ZN(U2856) );
  AOI22_X1 U7362 ( .A1(n6336), .A2(n6351), .B1(n6340), .B2(DATAI_18_), .ZN(
        n6338) );
  AOI22_X1 U7363 ( .A1(n6342), .A2(DATAI_2_), .B1(n6345), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7364 ( .A1(n6338), .A2(n6337), .ZN(U2873) );
  INV_X1 U7365 ( .A(n6339), .ZN(n6341) );
  AOI22_X1 U7366 ( .A1(n6341), .A2(n6351), .B1(n6340), .B2(DATAI_16_), .ZN(
        n6344) );
  AOI22_X1 U7367 ( .A1(n6342), .A2(DATAI_0_), .B1(n6345), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U7368 ( .A1(n6344), .A2(n6343), .ZN(U2875) );
  AOI22_X1 U7369 ( .A1(n6346), .A2(n6351), .B1(EAX_REG_15__SCAN_IN), .B2(n6345), .ZN(n6347) );
  OAI21_X1 U7370 ( .B1(n6349), .B2(n6348), .A(n6347), .ZN(U2876) );
  AOI22_X1 U7371 ( .A1(n6352), .A2(n6351), .B1(DATAI_12_), .B2(n6350), .ZN(
        n6353) );
  OAI21_X1 U7372 ( .B1(n3677), .B2(n6354), .A(n6353), .ZN(U2879) );
  AOI22_X1 U7373 ( .A1(n6359), .A2(EAX_REG_30__SCAN_IN), .B1(n6390), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6355) );
  OAI21_X1 U7374 ( .B1(n6356), .B2(n6369), .A(n6355), .ZN(U2893) );
  AOI22_X1 U7375 ( .A1(n6359), .A2(EAX_REG_26__SCAN_IN), .B1(n6390), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6357) );
  OAI21_X1 U7376 ( .B1(n6358), .B2(n6369), .A(n6357), .ZN(U2897) );
  AOI22_X1 U7377 ( .A1(n6359), .A2(EAX_REG_19__SCAN_IN), .B1(n6390), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n6360) );
  OAI21_X1 U7378 ( .B1(n6361), .B2(n6369), .A(n6360), .ZN(U2904) );
  INV_X1 U7379 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6363) );
  AOI22_X1 U7380 ( .A1(n6385), .A2(DATAO_REG_15__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6362) );
  OAI21_X1 U7381 ( .B1(n6363), .B2(n6392), .A(n6362), .ZN(U2908) );
  INV_X1 U7382 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6365) );
  AOI22_X1 U7383 ( .A1(n6385), .A2(DATAO_REG_14__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6364) );
  OAI21_X1 U7384 ( .B1(n6365), .B2(n6392), .A(n6364), .ZN(U2909) );
  AOI22_X1 U7385 ( .A1(n6385), .A2(DATAO_REG_12__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6366) );
  OAI21_X1 U7386 ( .B1(n3677), .B2(n6392), .A(n6366), .ZN(U2911) );
  AOI22_X1 U7387 ( .A1(n6367), .A2(EAX_REG_11__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6368) );
  OAI21_X1 U7388 ( .B1(n6370), .B2(n6369), .A(n6368), .ZN(U2912) );
  AOI22_X1 U7389 ( .A1(n6385), .A2(DATAO_REG_10__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6371) );
  OAI21_X1 U7390 ( .B1(n6372), .B2(n6392), .A(n6371), .ZN(U2913) );
  AOI22_X1 U7391 ( .A1(n6385), .A2(DATAO_REG_9__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6373) );
  OAI21_X1 U7392 ( .B1(n6374), .B2(n6392), .A(n6373), .ZN(U2914) );
  INV_X1 U7393 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6376) );
  AOI22_X1 U7394 ( .A1(n6385), .A2(DATAO_REG_8__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6375) );
  OAI21_X1 U7395 ( .B1(n6376), .B2(n6392), .A(n6375), .ZN(U2915) );
  AOI22_X1 U7396 ( .A1(n6385), .A2(DATAO_REG_7__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n6377) );
  OAI21_X1 U7397 ( .B1(n6378), .B2(n6392), .A(n6377), .ZN(U2916) );
  AOI22_X1 U7398 ( .A1(n6385), .A2(DATAO_REG_6__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n6379) );
  OAI21_X1 U7399 ( .B1(n6380), .B2(n6392), .A(n6379), .ZN(U2917) );
  AOI22_X1 U7400 ( .A1(n6385), .A2(DATAO_REG_5__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n6381) );
  OAI21_X1 U7401 ( .B1(n6382), .B2(n6392), .A(n6381), .ZN(U2918) );
  AOI22_X1 U7402 ( .A1(n6385), .A2(DATAO_REG_4__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n6383) );
  OAI21_X1 U7403 ( .B1(n6384), .B2(n6392), .A(n6383), .ZN(U2919) );
  AOI22_X1 U7404 ( .A1(n6385), .A2(DATAO_REG_3__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n6386) );
  OAI21_X1 U7405 ( .B1(n6387), .B2(n6392), .A(n6386), .ZN(U2920) );
  AOI22_X1 U7406 ( .A1(n6385), .A2(DATAO_REG_2__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n6388) );
  OAI21_X1 U7407 ( .B1(n6389), .B2(n6392), .A(n6388), .ZN(U2921) );
  AOI22_X1 U7408 ( .A1(n6385), .A2(DATAO_REG_1__SCAN_IN), .B1(n6390), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n6391) );
  OAI21_X1 U7409 ( .B1(n6393), .B2(n6392), .A(n6391), .ZN(U2922) );
  INV_X1 U7410 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6395) );
  AOI22_X1 U7411 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6416), .B1(n6409), .B2(
        DATAI_0_), .ZN(n6394) );
  OAI21_X1 U7412 ( .B1(n6395), .B2(n6418), .A(n6394), .ZN(U2924) );
  INV_X1 U7413 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6397) );
  AOI22_X1 U7414 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6416), .B1(n6409), .B2(
        DATAI_1_), .ZN(n6396) );
  OAI21_X1 U7415 ( .B1(n6397), .B2(n6418), .A(n6396), .ZN(U2925) );
  INV_X1 U7416 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6399) );
  AOI22_X1 U7417 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6416), .B1(n6409), .B2(
        DATAI_2_), .ZN(n6398) );
  OAI21_X1 U7418 ( .B1(n6399), .B2(n6418), .A(n6398), .ZN(U2926) );
  INV_X1 U7419 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U7420 ( .A1(n6409), .A2(DATAI_8_), .ZN(n6411) );
  INV_X1 U7421 ( .A(n6411), .ZN(n6400) );
  AOI21_X1 U7422 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6416), .A(n6400), .ZN(n6401) );
  OAI21_X1 U7423 ( .B1(n6402), .B2(n6418), .A(n6401), .ZN(U2932) );
  NAND2_X1 U7424 ( .A1(n6409), .A2(DATAI_11_), .ZN(n6413) );
  INV_X1 U7425 ( .A(n6413), .ZN(n6403) );
  AOI21_X1 U7426 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6416), .A(n6403), .ZN(
        n6404) );
  OAI21_X1 U7427 ( .B1(n3891), .B2(n6418), .A(n6404), .ZN(U2935) );
  INV_X1 U7428 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6408) );
  INV_X1 U7429 ( .A(DATAI_12_), .ZN(n6405) );
  NOR2_X1 U7430 ( .A1(n6406), .A2(n6405), .ZN(n6415) );
  AOI21_X1 U7431 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6416), .A(n6415), .ZN(
        n6407) );
  OAI21_X1 U7432 ( .B1(n6408), .B2(n6418), .A(n6407), .ZN(U2936) );
  AOI22_X1 U7433 ( .A1(n6416), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n6419), .ZN(n6410) );
  NAND2_X1 U7434 ( .A1(n6409), .A2(DATAI_14_), .ZN(n6421) );
  NAND2_X1 U7435 ( .A1(n6410), .A2(n6421), .ZN(U2938) );
  AOI22_X1 U7436 ( .A1(n6420), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6419), .ZN(n6412) );
  NAND2_X1 U7437 ( .A1(n6412), .A2(n6411), .ZN(U2947) );
  AOI22_X1 U7438 ( .A1(n6420), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n6419), .ZN(n6414) );
  NAND2_X1 U7439 ( .A1(n6414), .A2(n6413), .ZN(U2950) );
  AOI21_X1 U7440 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6416), .A(n6415), .ZN(
        n6417) );
  OAI21_X1 U7441 ( .B1(n3677), .B2(n6418), .A(n6417), .ZN(U2951) );
  AOI22_X1 U7442 ( .A1(n6420), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6419), .ZN(n6422) );
  NAND2_X1 U7443 ( .A1(n6422), .A2(n6421), .ZN(U2953) );
  AOI22_X1 U7444 ( .A1(n6450), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .B1(n6490), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6432) );
  NOR2_X1 U7445 ( .A1(n6424), .A2(n6423), .ZN(n6428) );
  INV_X1 U7446 ( .A(n6425), .ZN(n6426) );
  AOI21_X1 U7447 ( .B1(n6428), .B2(n6427), .A(n6426), .ZN(n6489) );
  INV_X1 U7448 ( .A(n6429), .ZN(n6430) );
  AOI22_X1 U7449 ( .A1(n6489), .A2(n6455), .B1(n6456), .B2(n6430), .ZN(n6431)
         );
  OAI211_X1 U7450 ( .C1(n6461), .C2(n6433), .A(n6432), .B(n6431), .ZN(U2979)
         );
  AND2_X1 U7451 ( .A1(n6490), .A2(REIP_REG_5__SCAN_IN), .ZN(n6509) );
  AOI21_X1 U7452 ( .B1(n6450), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6509), 
        .ZN(n6439) );
  INV_X1 U7453 ( .A(n6436), .ZN(n6514) );
  AOI22_X1 U7454 ( .A1(n6514), .A2(n6455), .B1(n6456), .B2(n6437), .ZN(n6438)
         );
  OAI211_X1 U7455 ( .C1(n6461), .C2(n6440), .A(n6439), .B(n6438), .ZN(U2981)
         );
  AND2_X1 U7456 ( .A1(n6490), .A2(REIP_REG_3__SCAN_IN), .ZN(n6519) );
  AOI21_X1 U7457 ( .B1(n6450), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6519), 
        .ZN(n6447) );
  INV_X1 U7458 ( .A(n6441), .ZN(n6442) );
  AOI21_X1 U7459 ( .B1(n6444), .B2(n6443), .A(n6442), .ZN(n6523) );
  AOI22_X1 U7460 ( .A1(n6523), .A2(n6455), .B1(n6456), .B2(n6445), .ZN(n6446)
         );
  OAI211_X1 U7461 ( .C1(n6461), .C2(n6448), .A(n6447), .B(n6446), .ZN(U2983)
         );
  NAND2_X1 U7462 ( .A1(n6490), .A2(REIP_REG_2__SCAN_IN), .ZN(n6543) );
  INV_X1 U7463 ( .A(n6543), .ZN(n6449) );
  AOI21_X1 U7464 ( .B1(n6450), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n6449), 
        .ZN(n6459) );
  INV_X1 U7465 ( .A(n6451), .ZN(n6457) );
  XNOR2_X1 U7466 ( .A(n6452), .B(n6540), .ZN(n6454) );
  XNOR2_X1 U7467 ( .A(n6454), .B(n6453), .ZN(n6536) );
  AOI22_X1 U7468 ( .A1(n6457), .A2(n6456), .B1(n6455), .B2(n6536), .ZN(n6458)
         );
  OAI211_X1 U7469 ( .C1(n6461), .C2(n6460), .A(n6459), .B(n6458), .ZN(U2984)
         );
  AOI21_X1 U7470 ( .B1(n6534), .B2(n6463), .A(n6462), .ZN(n6467) );
  AOI22_X1 U7471 ( .A1(n6465), .A2(n6537), .B1(n6468), .B2(n6464), .ZN(n6466)
         );
  OAI211_X1 U7472 ( .C1(n6469), .C2(n6468), .A(n6467), .B(n6466), .ZN(U3007)
         );
  INV_X1 U7473 ( .A(n6470), .ZN(n6477) );
  AOI21_X1 U7474 ( .B1(n6534), .B2(n6472), .A(n6471), .ZN(n6476) );
  AOI22_X1 U7475 ( .A1(n6474), .A2(n6537), .B1(n5223), .B2(n6473), .ZN(n6475)
         );
  OAI211_X1 U7476 ( .C1(n6477), .C2(n5223), .A(n6476), .B(n6475), .ZN(U3009)
         );
  AOI22_X1 U7477 ( .A1(n6534), .A2(n6478), .B1(n6490), .B2(REIP_REG_8__SCAN_IN), .ZN(n6482) );
  AOI211_X1 U7478 ( .C1(n6493), .C2(n6487), .A(n6479), .B(n6494), .ZN(n6480)
         );
  INV_X1 U7479 ( .A(n6480), .ZN(n6481) );
  OAI211_X1 U7480 ( .C1(n6484), .C2(n6483), .A(n6482), .B(n6481), .ZN(n6485)
         );
  INV_X1 U7481 ( .A(n6485), .ZN(n6486) );
  OAI21_X1 U7482 ( .B1(n6492), .B2(n6487), .A(n6486), .ZN(U3010) );
  AOI222_X1 U7483 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6490), .B1(n6537), .B2(
        n6489), .C1(n6488), .C2(n6534), .ZN(n6491) );
  OAI221_X1 U7484 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n6494), .C1(n6493), .C2(n6492), .A(n6491), .ZN(U3011) );
  INV_X1 U7485 ( .A(n6501), .ZN(n6507) );
  NAND2_X1 U7486 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6507), .ZN(n6495)
         );
  AOI21_X1 U7487 ( .B1(n6496), .B2(n6495), .A(n6538), .ZN(n6518) );
  INV_X1 U7488 ( .A(n6497), .ZN(n6498) );
  AOI21_X1 U7489 ( .B1(n6534), .B2(n6499), .A(n6498), .ZN(n6506) );
  INV_X1 U7490 ( .A(n6500), .ZN(n6504) );
  NOR3_X1 U7491 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6502), .A3(n6501), 
        .ZN(n6503) );
  AOI22_X1 U7492 ( .A1(n6504), .A2(n6537), .B1(n6503), .B2(n6521), .ZN(n6505)
         );
  OAI211_X1 U7493 ( .C1(n6518), .C2(n5209), .A(n6506), .B(n6505), .ZN(U3012)
         );
  AOI21_X1 U7494 ( .B1(n6508), .B2(n6507), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6517) );
  AOI21_X1 U7495 ( .B1(n6534), .B2(n6510), .A(n6509), .ZN(n6516) );
  NOR4_X1 U7496 ( .A1(n6539), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6512), 
        .A4(n6511), .ZN(n6513) );
  AOI21_X1 U7497 ( .B1(n6514), .B2(n6537), .A(n6513), .ZN(n6515) );
  OAI211_X1 U7498 ( .C1(n6518), .C2(n6517), .A(n6516), .B(n6515), .ZN(U3013)
         );
  AOI21_X1 U7499 ( .B1(n6534), .B2(n6520), .A(n6519), .ZN(n6526) );
  AND2_X1 U7500 ( .A1(n6522), .A2(n6521), .ZN(n6524) );
  AOI22_X1 U7501 ( .A1(n6524), .A2(n6527), .B1(n6523), .B2(n6537), .ZN(n6525)
         );
  OAI211_X1 U7502 ( .C1(n6528), .C2(n6527), .A(n6526), .B(n6525), .ZN(U3015)
         );
  INV_X1 U7503 ( .A(n6529), .ZN(n6535) );
  NOR3_X1 U7504 ( .A1(n6540), .A2(n6531), .A3(n6530), .ZN(n6532) );
  AOI211_X1 U7505 ( .C1(n6535), .C2(n6534), .A(n6533), .B(n6532), .ZN(n6545)
         );
  AOI22_X1 U7506 ( .A1(n6538), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6537), 
        .B2(n6536), .ZN(n6544) );
  INV_X1 U7507 ( .A(n6539), .ZN(n6541) );
  NAND3_X1 U7508 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6541), .A3(n6540), 
        .ZN(n6542) );
  NAND4_X1 U7509 ( .A1(n6545), .A2(n6544), .A3(n6543), .A4(n6542), .ZN(U3016)
         );
  NOR2_X1 U7510 ( .A1(n6546), .A2(n6778), .ZN(U3019) );
  AND2_X1 U7511 ( .A1(n6780), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6549)
         );
  AND2_X1 U7512 ( .A1(n6554), .A2(n6549), .ZN(n6577) );
  AOI22_X1 U7513 ( .A1(n6578), .A2(n6690), .B1(n6683), .B2(n6577), .ZN(n6564)
         );
  NAND2_X1 U7514 ( .A1(n6550), .A2(n6677), .ZN(n6771) );
  NAND2_X1 U7515 ( .A1(n6679), .A2(n6551), .ZN(n6552) );
  OAI21_X1 U7516 ( .B1(n6771), .B2(n6552), .A(n6774), .ZN(n6562) );
  AOI21_X1 U7517 ( .B1(n6553), .B2(n3466), .A(n6577), .ZN(n6557) );
  INV_X1 U7518 ( .A(n6554), .ZN(n6556) );
  OAI22_X1 U7519 ( .A1(n6562), .A2(n6557), .B1(n6556), .B2(n6555), .ZN(n6580)
         );
  INV_X1 U7520 ( .A(n6557), .ZN(n6561) );
  AOI21_X1 U7521 ( .B1(n6678), .B2(n6559), .A(n6558), .ZN(n6560) );
  AOI22_X1 U7522 ( .A1(n6628), .A2(n6580), .B1(n6579), .B2(
        INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6563) );
  OAI211_X1 U7523 ( .C1(n6637), .C2(n6620), .A(n6564), .B(n6563), .ZN(U3044)
         );
  AOI22_X1 U7524 ( .A1(n6578), .A2(n6696), .B1(n6694), .B2(n6577), .ZN(n6566)
         );
  AOI22_X1 U7525 ( .A1(n6638), .A2(n6580), .B1(n6579), .B2(
        INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6565) );
  OAI211_X1 U7526 ( .C1(n6641), .C2(n6620), .A(n6566), .B(n6565), .ZN(U3045)
         );
  AOI22_X1 U7527 ( .A1(n6578), .A2(n6702), .B1(n6700), .B2(n6577), .ZN(n6568)
         );
  AOI22_X1 U7528 ( .A1(n6642), .A2(n6580), .B1(n6579), .B2(
        INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6567) );
  OAI211_X1 U7529 ( .C1(n6645), .C2(n6620), .A(n6568), .B(n6567), .ZN(U3046)
         );
  AOI22_X1 U7530 ( .A1(n6578), .A2(n6708), .B1(n6706), .B2(n6577), .ZN(n6570)
         );
  AOI22_X1 U7531 ( .A1(n6646), .A2(n6580), .B1(n6579), .B2(
        INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6569) );
  OAI211_X1 U7532 ( .C1(n6649), .C2(n6620), .A(n6570), .B(n6569), .ZN(U3047)
         );
  AOI22_X1 U7533 ( .A1(n6578), .A2(n6652), .B1(n6650), .B2(n6577), .ZN(n6572)
         );
  AOI22_X1 U7534 ( .A1(n6651), .A2(n6580), .B1(n6579), .B2(
        INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6571) );
  OAI211_X1 U7535 ( .C1(n6655), .C2(n6620), .A(n6572), .B(n6571), .ZN(U3048)
         );
  AOI22_X1 U7536 ( .A1(n6578), .A2(n6658), .B1(n6656), .B2(n6577), .ZN(n6574)
         );
  AOI22_X1 U7537 ( .A1(n6657), .A2(n6580), .B1(n6579), .B2(
        INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6573) );
  OAI211_X1 U7538 ( .C1(n6661), .C2(n6620), .A(n6574), .B(n6573), .ZN(U3049)
         );
  AOI22_X1 U7539 ( .A1(n6578), .A2(n6730), .B1(n6727), .B2(n6577), .ZN(n6576)
         );
  AOI22_X1 U7540 ( .A1(n6662), .A2(n6580), .B1(n6579), .B2(
        INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6575) );
  OAI211_X1 U7541 ( .C1(n6665), .C2(n6620), .A(n6576), .B(n6575), .ZN(U3050)
         );
  AOI22_X1 U7542 ( .A1(n6578), .A2(n6671), .B1(n6667), .B2(n6577), .ZN(n6582)
         );
  AOI22_X1 U7543 ( .A1(n6668), .A2(n6580), .B1(n6579), .B2(
        INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6581) );
  OAI211_X1 U7544 ( .C1(n6676), .C2(n6620), .A(n6582), .B(n6581), .ZN(U3051)
         );
  INV_X1 U7545 ( .A(n6583), .ZN(n6584) );
  OAI22_X1 U7546 ( .A1(n6625), .A2(n6586), .B1(n6585), .B2(n6584), .ZN(n6615)
         );
  NAND2_X1 U7547 ( .A1(n6587), .A2(n6626), .ZN(n6590) );
  AOI22_X1 U7548 ( .A1(n6615), .A2(n6628), .B1(n6683), .B2(n6614), .ZN(n6596)
         );
  OAI211_X1 U7549 ( .C1(n6776), .C2(n6620), .A(n6589), .B(n6588), .ZN(n6594)
         );
  NAND2_X1 U7550 ( .A1(n6590), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6591) );
  NAND4_X1 U7551 ( .A1(n6594), .A2(n6593), .A3(n6592), .A4(n6591), .ZN(n6617)
         );
  AOI22_X1 U7552 ( .A1(n6617), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6684), 
        .B2(n6616), .ZN(n6595) );
  OAI211_X1 U7553 ( .C1(n6597), .C2(n6620), .A(n6596), .B(n6595), .ZN(U3052)
         );
  AOI22_X1 U7554 ( .A1(n6615), .A2(n6638), .B1(n6694), .B2(n6614), .ZN(n6599)
         );
  AOI22_X1 U7555 ( .A1(n6617), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6695), 
        .B2(n6616), .ZN(n6598) );
  OAI211_X1 U7556 ( .C1(n6600), .C2(n6620), .A(n6599), .B(n6598), .ZN(U3053)
         );
  AOI22_X1 U7557 ( .A1(n6615), .A2(n6642), .B1(n6700), .B2(n6614), .ZN(n6602)
         );
  AOI22_X1 U7558 ( .A1(n6617), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6701), 
        .B2(n6616), .ZN(n6601) );
  OAI211_X1 U7559 ( .C1(n6603), .C2(n6620), .A(n6602), .B(n6601), .ZN(U3054)
         );
  AOI22_X1 U7560 ( .A1(n6615), .A2(n6646), .B1(n6706), .B2(n6614), .ZN(n6605)
         );
  AOI22_X1 U7561 ( .A1(n6617), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6707), 
        .B2(n6616), .ZN(n6604) );
  OAI211_X1 U7562 ( .C1(n6606), .C2(n6620), .A(n6605), .B(n6604), .ZN(U3055)
         );
  AOI22_X1 U7563 ( .A1(n6615), .A2(n6651), .B1(n6650), .B2(n6614), .ZN(n6608)
         );
  AOI22_X1 U7564 ( .A1(n6617), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6715), 
        .B2(n6616), .ZN(n6607) );
  OAI211_X1 U7565 ( .C1(n6713), .C2(n6620), .A(n6608), .B(n6607), .ZN(U3056)
         );
  AOI22_X1 U7566 ( .A1(n6615), .A2(n6657), .B1(n6656), .B2(n6614), .ZN(n6610)
         );
  AOI22_X1 U7567 ( .A1(n6617), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6722), 
        .B2(n6616), .ZN(n6609) );
  OAI211_X1 U7568 ( .C1(n6720), .C2(n6620), .A(n6610), .B(n6609), .ZN(U3057)
         );
  AOI22_X1 U7569 ( .A1(n6615), .A2(n6662), .B1(n6727), .B2(n6614), .ZN(n6612)
         );
  AOI22_X1 U7570 ( .A1(n6617), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6728), 
        .B2(n6616), .ZN(n6611) );
  OAI211_X1 U7571 ( .C1(n6613), .C2(n6620), .A(n6612), .B(n6611), .ZN(U3058)
         );
  AOI22_X1 U7572 ( .A1(n6615), .A2(n6668), .B1(n6667), .B2(n6614), .ZN(n6619)
         );
  AOI22_X1 U7573 ( .A1(n6617), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6740), 
        .B2(n6616), .ZN(n6618) );
  OAI211_X1 U7574 ( .C1(n6736), .C2(n6620), .A(n6619), .B(n6618), .ZN(U3059)
         );
  NAND3_X1 U7575 ( .A1(n6622), .A2(n6621), .A3(n6780), .ZN(n6623) );
  OAI21_X1 U7576 ( .B1(n6625), .B2(n6624), .A(n6623), .ZN(n6669) );
  NAND2_X1 U7577 ( .A1(n6627), .A2(n6626), .ZN(n6631) );
  INV_X1 U7578 ( .A(n6631), .ZN(n6666) );
  AOI22_X1 U7579 ( .A1(n6669), .A2(n6628), .B1(n6683), .B2(n6666), .ZN(n6636)
         );
  NAND3_X1 U7580 ( .A1(n6634), .A2(n6629), .A3(n6675), .ZN(n6633) );
  AOI211_X1 U7581 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6631), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6630), .ZN(n6632) );
  AOI22_X1 U7582 ( .A1(n6672), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6690), 
        .B2(n6670), .ZN(n6635) );
  OAI211_X1 U7583 ( .C1(n6637), .C2(n6675), .A(n6636), .B(n6635), .ZN(U3068)
         );
  AOI22_X1 U7584 ( .A1(n6669), .A2(n6638), .B1(n6694), .B2(n6666), .ZN(n6640)
         );
  AOI22_X1 U7585 ( .A1(n6672), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6696), 
        .B2(n6670), .ZN(n6639) );
  OAI211_X1 U7586 ( .C1(n6641), .C2(n6675), .A(n6640), .B(n6639), .ZN(U3069)
         );
  AOI22_X1 U7587 ( .A1(n6669), .A2(n6642), .B1(n6700), .B2(n6666), .ZN(n6644)
         );
  AOI22_X1 U7588 ( .A1(n6672), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6702), 
        .B2(n6670), .ZN(n6643) );
  OAI211_X1 U7589 ( .C1(n6645), .C2(n6675), .A(n6644), .B(n6643), .ZN(U3070)
         );
  AOI22_X1 U7590 ( .A1(n6669), .A2(n6646), .B1(n6706), .B2(n6666), .ZN(n6648)
         );
  AOI22_X1 U7591 ( .A1(n6672), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6708), 
        .B2(n6670), .ZN(n6647) );
  OAI211_X1 U7592 ( .C1(n6649), .C2(n6675), .A(n6648), .B(n6647), .ZN(U3071)
         );
  AOI22_X1 U7593 ( .A1(n6669), .A2(n6651), .B1(n6650), .B2(n6666), .ZN(n6654)
         );
  AOI22_X1 U7594 ( .A1(n6672), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6652), 
        .B2(n6670), .ZN(n6653) );
  OAI211_X1 U7595 ( .C1(n6655), .C2(n6675), .A(n6654), .B(n6653), .ZN(U3072)
         );
  AOI22_X1 U7596 ( .A1(n6669), .A2(n6657), .B1(n6656), .B2(n6666), .ZN(n6660)
         );
  AOI22_X1 U7597 ( .A1(n6672), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6658), 
        .B2(n6670), .ZN(n6659) );
  OAI211_X1 U7598 ( .C1(n6661), .C2(n6675), .A(n6660), .B(n6659), .ZN(U3073)
         );
  AOI22_X1 U7599 ( .A1(n6669), .A2(n6662), .B1(n6727), .B2(n6666), .ZN(n6664)
         );
  AOI22_X1 U7600 ( .A1(n6672), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6730), 
        .B2(n6670), .ZN(n6663) );
  OAI211_X1 U7601 ( .C1(n6665), .C2(n6675), .A(n6664), .B(n6663), .ZN(U3074)
         );
  AOI22_X1 U7602 ( .A1(n6669), .A2(n6668), .B1(n6667), .B2(n6666), .ZN(n6674)
         );
  AOI22_X1 U7603 ( .A1(n6672), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6671), 
        .B2(n6670), .ZN(n6673) );
  OAI211_X1 U7604 ( .C1(n6676), .C2(n6675), .A(n6674), .B(n6673), .ZN(U3075)
         );
  INV_X1 U7605 ( .A(n6677), .ZN(n6680) );
  AOI21_X1 U7606 ( .B1(n6680), .B2(n6679), .A(n6678), .ZN(n6686) );
  AND2_X1 U7607 ( .A1(n6689), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6726)
         );
  AOI21_X1 U7608 ( .B1(n6681), .B2(n3466), .A(n6726), .ZN(n6685) );
  INV_X1 U7609 ( .A(n6685), .ZN(n6682) );
  AOI22_X1 U7610 ( .A1(n6739), .A2(n6684), .B1(n6683), .B2(n6726), .ZN(n6692)
         );
  NAND2_X1 U7611 ( .A1(n6686), .A2(n6685), .ZN(n6688) );
  OAI211_X1 U7612 ( .C1(n6774), .C2(n6689), .A(n6688), .B(n6687), .ZN(n6741)
         );
  AOI22_X1 U7613 ( .A1(n6741), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n6690), 
        .B2(n6729), .ZN(n6691) );
  OAI211_X1 U7614 ( .C1(n6745), .C2(n6693), .A(n6692), .B(n6691), .ZN(U3108)
         );
  AOI22_X1 U7615 ( .A1(n6739), .A2(n6695), .B1(n6694), .B2(n6726), .ZN(n6698)
         );
  AOI22_X1 U7616 ( .A1(n6741), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n6696), 
        .B2(n6729), .ZN(n6697) );
  OAI211_X1 U7617 ( .C1(n6745), .C2(n6699), .A(n6698), .B(n6697), .ZN(U3109)
         );
  AOI22_X1 U7618 ( .A1(n6739), .A2(n6701), .B1(n6700), .B2(n6726), .ZN(n6704)
         );
  AOI22_X1 U7619 ( .A1(n6741), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n6702), 
        .B2(n6729), .ZN(n6703) );
  OAI211_X1 U7620 ( .C1(n6745), .C2(n6705), .A(n6704), .B(n6703), .ZN(U3110)
         );
  AOI22_X1 U7621 ( .A1(n6739), .A2(n6707), .B1(n6706), .B2(n6726), .ZN(n6710)
         );
  AOI22_X1 U7622 ( .A1(n6741), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n6708), 
        .B2(n6729), .ZN(n6709) );
  OAI211_X1 U7623 ( .C1(n6745), .C2(n6711), .A(n6710), .B(n6709), .ZN(U3111)
         );
  INV_X1 U7624 ( .A(n6726), .ZN(n6734) );
  OAI22_X1 U7625 ( .A1(n6737), .A2(n6713), .B1(n6712), .B2(n6734), .ZN(n6714)
         );
  INV_X1 U7626 ( .A(n6714), .ZN(n6717) );
  AOI22_X1 U7627 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6741), .B1(n6715), 
        .B2(n6739), .ZN(n6716) );
  OAI211_X1 U7628 ( .C1(n6745), .C2(n6718), .A(n6717), .B(n6716), .ZN(U3112)
         );
  OAI22_X1 U7629 ( .A1(n6737), .A2(n6720), .B1(n6719), .B2(n6734), .ZN(n6721)
         );
  INV_X1 U7630 ( .A(n6721), .ZN(n6724) );
  AOI22_X1 U7631 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6741), .B1(n6722), 
        .B2(n6739), .ZN(n6723) );
  OAI211_X1 U7632 ( .C1(n6745), .C2(n6725), .A(n6724), .B(n6723), .ZN(U3113)
         );
  AOI22_X1 U7633 ( .A1(n6739), .A2(n6728), .B1(n6727), .B2(n6726), .ZN(n6732)
         );
  AOI22_X1 U7634 ( .A1(n6741), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n6730), 
        .B2(n6729), .ZN(n6731) );
  OAI211_X1 U7635 ( .C1(n6745), .C2(n6733), .A(n6732), .B(n6731), .ZN(U3114)
         );
  OAI22_X1 U7636 ( .A1(n6737), .A2(n6736), .B1(n6735), .B2(n6734), .ZN(n6738)
         );
  INV_X1 U7637 ( .A(n6738), .ZN(n6743) );
  AOI22_X1 U7638 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6741), .B1(n6740), 
        .B2(n6739), .ZN(n6742) );
  OAI211_X1 U7639 ( .C1(n6745), .C2(n6744), .A(n6743), .B(n6742), .ZN(U3115)
         );
  INV_X1 U7640 ( .A(n6746), .ZN(n6749) );
  NOR3_X1 U7641 ( .A1(n6749), .A2(n6748), .A3(n6747), .ZN(n6755) );
  INV_X1 U7642 ( .A(n6770), .ZN(n6753) );
  AOI21_X1 U7643 ( .B1(n6751), .B2(n4179), .A(n6750), .ZN(n6752) );
  NOR2_X1 U7644 ( .A1(n6753), .A2(n6752), .ZN(n6754) );
  OR3_X1 U7645 ( .A1(n6756), .A2(n6755), .A3(n6754), .ZN(U3149) );
  AND2_X1 U7646 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6761), .ZN(U3151) );
  NOR2_X1 U7647 ( .A1(n6765), .A2(n6757), .ZN(U3152) );
  AND2_X1 U7648 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6761), .ZN(U3153) );
  AND2_X1 U7649 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6761), .ZN(U3154) );
  AND2_X1 U7650 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6761), .ZN(U3155) );
  AND2_X1 U7651 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6761), .ZN(U3156) );
  AND2_X1 U7652 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6761), .ZN(U3157) );
  AND2_X1 U7653 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6761), .ZN(U3158) );
  AND2_X1 U7654 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6761), .ZN(U3159) );
  AND2_X1 U7655 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6761), .ZN(U3160) );
  NOR2_X1 U7656 ( .A1(n6765), .A2(n6758), .ZN(U3161) );
  AND2_X1 U7657 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6761), .ZN(U3162) );
  AND2_X1 U7658 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6761), .ZN(U3163) );
  AND2_X1 U7659 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6761), .ZN(U3164) );
  AND2_X1 U7660 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6761), .ZN(U3165) );
  AND2_X1 U7661 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6761), .ZN(U3166) );
  NOR2_X1 U7662 ( .A1(n6765), .A2(n5705), .ZN(U3167) );
  AND2_X1 U7663 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6761), .ZN(U3168) );
  AND2_X1 U7664 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6761), .ZN(U3169) );
  AND2_X1 U7665 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6761), .ZN(U3170) );
  AND2_X1 U7666 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6761), .ZN(U3171) );
  AND2_X1 U7667 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6761), .ZN(U3172) );
  AND2_X1 U7668 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6761), .ZN(U3173) );
  AND2_X1 U7669 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6761), .ZN(U3174) );
  NOR2_X1 U7670 ( .A1(n6765), .A2(n6759), .ZN(U3175) );
  AND2_X1 U7671 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6761), .ZN(U3176) );
  AND2_X1 U7672 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6761), .ZN(U3177) );
  AND2_X1 U7673 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6761), .ZN(U3178) );
  AND2_X1 U7674 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6761), .ZN(U3179) );
  AND2_X1 U7675 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6761), .ZN(U3180) );
  INV_X1 U7676 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6762) );
  INV_X1 U7677 ( .A(n6763), .ZN(n6760) );
  AOI21_X1 U7678 ( .B1(n6762), .B2(n6761), .A(n6760), .ZN(U3451) );
  OAI21_X1 U7679 ( .B1(n6765), .B2(n6764), .A(n6763), .ZN(U3452) );
  INV_X1 U7680 ( .A(n6766), .ZN(n6768) );
  OAI211_X1 U7681 ( .C1(n6770), .C2(n6769), .A(n6768), .B(n6767), .ZN(U3453)
         );
  INV_X1 U7682 ( .A(n6771), .ZN(n6773) );
  NAND2_X1 U7683 ( .A1(n6773), .A2(n6772), .ZN(n6775) );
  AOI222_X1 U7684 ( .A1(n6777), .A2(n2977), .B1(n4642), .B2(n6776), .C1(n6775), 
        .C2(n6774), .ZN(n6779) );
  AOI22_X1 U7685 ( .A1(n6781), .A2(n6780), .B1(n6779), .B2(n6778), .ZN(U3462)
         );
  AOI21_X1 U7686 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6783) );
  AOI22_X1 U7687 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6783), .B2(n6782), .ZN(n6785) );
  AOI22_X1 U7688 ( .A1(n6786), .A2(n6785), .B1(n6784), .B2(n6789), .ZN(U3468)
         );
  NOR2_X1 U7689 ( .A1(n6789), .A2(REIP_REG_1__SCAN_IN), .ZN(n6787) );
  AOI22_X1 U7690 ( .A1(n6790), .A2(n6789), .B1(n6788), .B2(n6787), .ZN(U3469)
         );
  NOR2_X1 U7691 ( .A1(n6791), .A2(READY_N), .ZN(n6793) );
  NOR3_X1 U7692 ( .A1(n6794), .A2(n6793), .A3(n6792), .ZN(n6801) );
  OAI211_X1 U7693 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6796), .A(n6795), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6798) );
  AOI21_X1 U7694 ( .B1(n6798), .B2(STATE2_REG_0__SCAN_IN), .A(n6797), .ZN(
        n6800) );
  NAND2_X1 U7695 ( .A1(n6801), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6799) );
  OAI21_X1 U7696 ( .B1(n6801), .B2(n6800), .A(n6799), .ZN(U3472) );
  AND2_X1 U4018 ( .A1(n3143), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3148)
         );
  AND2_X1 U3431 ( .A1(n4449), .A2(n3011), .ZN(n3310) );
  BUF_X1 U34640 ( .A(n3301), .Z(n4400) );
  OR2_X1 U4092 ( .A1(n3260), .A2(n3259), .ZN(n3385) );
  OR2_X1 U3425 ( .A1(n3246), .A2(n3245), .ZN(n3289) );
  CLKBUF_X1 U3437 ( .A(n3248), .Z(n4432) );
  CLKBUF_X2 U34600 ( .A(n3310), .Z(n3824) );
  CLKBUF_X1 U3504 ( .A(n4495), .Z(n4764) );
  CLKBUF_X1 U3816 ( .A(n5307), .Z(n5308) );
  CLKBUF_X1 U3884 ( .A(n4501), .Z(n5452) );
  CLKBUF_X1 U3887 ( .A(n4446), .Z(n2977) );
  AOI211_X1 U4051 ( .C1(n5576), .C2(n6456), .A(n5575), .B(n5574), .ZN(n5577)
         );
  AND2_X2 U4052 ( .A1(n3383), .A2(n3031), .ZN(n6802) );
  OR3_X1 U4078 ( .A1(n5553), .A2(n2991), .A3(n5934), .ZN(n6803) );
  CLKBUF_X1 U4326 ( .A(n3436), .Z(n3437) );
endmodule

