

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566;

  OR2_X1 U4878 ( .A1(n6394), .A2(n6393), .ZN(n4471) );
  NAND2_X2 U4879 ( .A1(n5246), .A2(n5245), .ZN(n8677) );
  CLKBUF_X2 U4880 ( .A(n6934), .Z(n7043) );
  INV_X1 U4881 ( .A(n9431), .ZN(n6518) );
  INV_X1 U4882 ( .A(n5336), .ZN(n5799) );
  CLKBUF_X1 U4883 ( .A(n5298), .Z(n5800) );
  INV_X1 U4884 ( .A(n5298), .ZN(n5776) );
  CLKBUF_X1 U4885 ( .A(n5300), .Z(n5733) );
  CLKBUF_X2 U4886 ( .A(n6074), .Z(n4384) );
  MUX2_X1 U4887 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6089), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n6090) );
  AND2_X1 U4888 ( .A1(n4372), .A2(n5171), .ZN(n5183) );
  AOI21_X1 U4889 ( .B1(n8406), .B2(n8398), .A(n8400), .ZN(n6707) );
  INV_X1 U4890 ( .A(n6905), .ZN(n6897) );
  NOR2_X1 U4891 ( .A1(n8115), .A2(n8114), .ZN(n8197) );
  INV_X1 U4892 ( .A(n4383), .ZN(n6203) );
  INV_X1 U4893 ( .A(n4384), .ZN(n6047) );
  NAND2_X1 U4894 ( .A1(n10350), .A2(n10079), .ZN(n9492) );
  AND2_X1 U4895 ( .A1(n5328), .A2(n5847), .ZN(n8687) );
  INV_X2 U4896 ( .A(n5325), .ZN(n5569) );
  XNOR2_X1 U4897 ( .A(n5231), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U4898 ( .A1(n9188), .A2(n9189), .ZN(n9187) );
  INV_X1 U4899 ( .A(n4380), .ZN(n9546) );
  BUF_X1 U4900 ( .A(n6403), .Z(n4386) );
  NAND2_X1 U4901 ( .A1(n9507), .A2(n9944), .ZN(n9965) );
  NAND2_X1 U4902 ( .A1(n6090), .A2(n10279), .ZN(n6091) );
  INV_X1 U4903 ( .A(n8041), .ZN(n8216) );
  NAND2_X1 U4904 ( .A1(n5588), .A2(n5587), .ZN(n8499) );
  INV_X1 U4905 ( .A(n8092), .ZN(n8711) );
  INV_X1 U4906 ( .A(n9551), .ZN(n9540) );
  OAI211_X1 U4907 ( .C1(n7173), .C2(n9614), .A(n5968), .B(n5967), .ZN(n10360)
         );
  NAND4_X1 U4908 ( .A1(n6080), .A2(n5026), .A3(n4696), .A4(n5932), .ZN(n6088)
         );
  OAI21_X1 U4909 ( .B1(n6103), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U4910 ( .A1(n5931), .A2(n6088), .ZN(n6095) );
  XNOR2_X1 U4911 ( .A(n6082), .B(n6104), .ZN(n9431) );
  AND4_X1 U4912 ( .A1(n5168), .A2(n5217), .A3(n5220), .A4(n5241), .ZN(n4372)
         );
  NAND2_X2 U4913 ( .A1(n7446), .A2(n6603), .ZN(n6604) );
  INV_X4 U4914 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8078) );
  NAND3_X1 U4915 ( .A1(n6883), .A2(n9950), .A3(n6886), .ZN(n4373) );
  NAND3_X2 U4916 ( .A1(n6883), .A2(n9950), .A3(n6886), .ZN(n7076) );
  NAND3_X2 U4917 ( .A1(n4854), .A2(n5308), .A3(n4855), .ZN(n5419) );
  NAND2_X2 U4918 ( .A1(n9214), .A2(n10104), .ZN(n9322) );
  NAND2_X2 U4919 ( .A1(n8030), .A2(n6187), .ZN(n6189) );
  AOI22_X2 U4920 ( .A1(n8317), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n6612), .B2(
        n4647), .ZN(n8322) );
  NAND2_X1 U4921 ( .A1(n6096), .A2(n6095), .ZN(n4374) );
  NAND2_X1 U4922 ( .A1(n6096), .A2(n6095), .ZN(n4375) );
  NAND2_X2 U4923 ( .A1(n6096), .A2(n6095), .ZN(n7173) );
  NAND2_X2 U4924 ( .A1(n8798), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5193) );
  OAI21_X1 U4925 ( .B1(n6759), .B2(n6758), .A(n6757), .ZN(n4376) );
  INV_X1 U4926 ( .A(n9571), .ZN(n10108) );
  OAI21_X2 U4927 ( .B1(n8456), .B2(n6193), .A(n6192), .ZN(n8446) );
  NAND2_X2 U4928 ( .A1(n4977), .A2(n4974), .ZN(n8456) );
  OAI21_X2 U4929 ( .B1(n5401), .B2(n4803), .A(n5074), .ZN(n5439) );
  NAND2_X2 U4930 ( .A1(n5116), .A2(n5115), .ZN(n5401) );
  NOR2_X2 U4931 ( .A1(n9211), .A2(n5090), .ZN(n7824) );
  NAND2_X2 U4932 ( .A1(n4527), .A2(n6052), .ZN(n10256) );
  NAND2_X2 U4933 ( .A1(n5256), .A2(n5255), .ZN(n8579) );
  OAI222_X1 U4934 ( .A1(n8105), .A2(n7793), .B1(P1_U3086), .B2(n9431), .C1(
        n10283), .C2(n7792), .ZN(P1_U3334) );
  NAND2_X2 U4935 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  NOR3_X1 U4936 ( .A1(n9421), .A2(n9707), .A3(n9447), .ZN(n9424) );
  NAND2_X1 U4937 ( .A1(n6062), .A2(n6061), .ZN(n9735) );
  NAND2_X1 U4938 ( .A1(n8893), .A2(n6987), .ZN(n9188) );
  AND2_X1 U4939 ( .A1(n6505), .A2(n9820), .ZN(n9523) );
  NOR2_X1 U4940 ( .A1(n9965), .A2(n5021), .ZN(n5024) );
  OR2_X1 U4941 ( .A1(n9955), .A2(n9967), .ZN(n9508) );
  INV_X2 U4942 ( .A(n10112), .ZN(n4377) );
  NAND2_X1 U4943 ( .A1(n9492), .A2(n10031), .ZN(n10074) );
  NAND2_X2 U4944 ( .A1(n9490), .A2(n6472), .ZN(n10366) );
  INV_X2 U4945 ( .A(n9568), .ZN(n10350) );
  INV_X1 U4946 ( .A(n10343), .ZN(n10403) );
  INV_X1 U4947 ( .A(n10364), .ZN(n10361) );
  AND4_X1 U4948 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(n10058)
         );
  INV_X2 U4949 ( .A(n10360), .ZN(n10392) );
  NAND2_X1 U4950 ( .A1(n4373), .A2(n6934), .ZN(n6905) );
  NAND2_X2 U4951 ( .A1(n6886), .A2(n6885), .ZN(n7070) );
  INV_X1 U4952 ( .A(n5305), .ZN(n4379) );
  INV_X2 U4953 ( .A(n6436), .ZN(n6533) );
  INV_X1 U4954 ( .A(n6263), .ZN(n6303) );
  CLKBUF_X2 U4955 ( .A(n6265), .Z(n6436) );
  INV_X4 U4956 ( .A(n6067), .ZN(n5983) );
  INV_X1 U4957 ( .A(n6259), .ZN(n4378) );
  INV_X1 U4958 ( .A(n6091), .ZN(n6246) );
  OR2_X1 U4959 ( .A1(n6297), .A2(n6296), .ZN(n6312) );
  AOI21_X1 U4960 ( .B1(n4547), .B2(n8696), .A(n4544), .ZN(n8721) );
  XNOR2_X1 U4961 ( .A(n8439), .B(n8438), .ZN(n4547) );
  OR3_X1 U4962 ( .A1(n8816), .A2(n7086), .A3(n7084), .ZN(n7112) );
  INV_X1 U4963 ( .A(n8446), .ZN(n4998) );
  OR2_X1 U4964 ( .A1(n4683), .A2(n5897), .ZN(n4680) );
  OAI211_X1 U4965 ( .C1(n5748), .C2(n4698), .A(n4453), .B(n4697), .ZN(n4812)
         );
  CLKBUF_X1 U4966 ( .A(n9200), .Z(n9201) );
  OAI21_X1 U4967 ( .B1(n9200), .B2(n5042), .A(n4412), .ZN(n9286) );
  XNOR2_X1 U4968 ( .A(n5796), .B(n5795), .ZN(n8797) );
  NAND2_X1 U4969 ( .A1(n6185), .A2(n4396), .ZN(n4967) );
  OR2_X1 U4970 ( .A1(n6522), .A2(n7106), .ZN(n5086) );
  INV_X1 U4971 ( .A(n9444), .ZN(n4958) );
  NAND2_X1 U4972 ( .A1(n4626), .A2(n6511), .ZN(n9758) );
  AND2_X1 U4973 ( .A1(n9407), .A2(n9411), .ZN(n9444) );
  NAND2_X1 U4974 ( .A1(n9799), .A2(n9386), .ZN(n9800) );
  NOR2_X1 U4975 ( .A1(n8376), .A2(n8540), .ZN(n8395) );
  OR2_X1 U4976 ( .A1(n8136), .A2(n6816), .ZN(n6819) );
  NAND2_X1 U4977 ( .A1(n4462), .A2(n8520), .ZN(n4667) );
  NAND2_X2 U4978 ( .A1(n9276), .A2(n9271), .ZN(n8857) );
  XNOR2_X1 U4979 ( .A(n5723), .B(n5722), .ZN(n7976) );
  NAND2_X1 U4980 ( .A1(n4824), .A2(n5691), .ZN(n5723) );
  INV_X1 U4981 ( .A(n4981), .ZN(n4980) );
  AOI21_X1 U4982 ( .B1(n4865), .B2(n8282), .A(n4503), .ZN(n4864) );
  NAND2_X1 U4983 ( .A1(n5686), .A2(n5685), .ZN(n5713) );
  NAND2_X1 U4984 ( .A1(n6058), .A2(n6057), .ZN(n9767) );
  NAND2_X1 U4985 ( .A1(n4929), .A2(n4928), .ZN(n9922) );
  OAI21_X1 U4986 ( .B1(n9241), .B2(n4463), .A(n5052), .ZN(n6985) );
  NAND2_X1 U4987 ( .A1(n6056), .A2(n6055), .ZN(n9787) );
  OR2_X1 U4988 ( .A1(n9368), .A2(n9367), .ZN(n4772) );
  AND2_X1 U4989 ( .A1(n4775), .A2(n4774), .ZN(n4773) );
  NAND2_X1 U4990 ( .A1(n9242), .A2(n9243), .ZN(n9241) );
  NAND2_X1 U4991 ( .A1(n7979), .A2(n6971), .ZN(n9242) );
  NOR2_X1 U4992 ( .A1(n9373), .A2(n9372), .ZN(n4775) );
  NAND2_X1 U4993 ( .A1(n4862), .A2(n4441), .ZN(n7492) );
  INV_X1 U4994 ( .A(n9853), .ZN(n10180) );
  NAND2_X1 U4995 ( .A1(n7372), .A2(n6780), .ZN(n7435) );
  AND2_X1 U4996 ( .A1(n6051), .A2(n6050), .ZN(n9853) );
  NAND2_X1 U4997 ( .A1(n6054), .A2(n6053), .ZN(n9808) );
  NAND2_X1 U4998 ( .A1(n6036), .A2(n6035), .ZN(n9881) );
  NAND2_X1 U4999 ( .A1(n5553), .A2(n5552), .ZN(n8755) );
  AND2_X1 U5000 ( .A1(n5571), .A2(n5570), .ZN(n8041) );
  NAND2_X1 U5001 ( .A1(n6777), .A2(n4493), .ZN(n7372) );
  NAND2_X1 U5002 ( .A1(n5224), .A2(n5223), .ZN(n8767) );
  NAND2_X1 U5003 ( .A1(n4844), .A2(n5167), .ZN(n5544) );
  NAND2_X1 U5004 ( .A1(n9508), .A2(n9354), .ZN(n9947) );
  NAND2_X1 U5005 ( .A1(n6028), .A2(n6027), .ZN(n10271) );
  NAND2_X1 U5006 ( .A1(n5500), .A2(n5499), .ZN(n8785) );
  NAND2_X1 U5007 ( .A1(n5162), .A2(n5161), .ZN(n5211) );
  NAND2_X1 U5008 ( .A1(n6022), .A2(n6021), .ZN(n10208) );
  OR2_X1 U5009 ( .A1(n7445), .A2(n7444), .ZN(n7642) );
  NAND2_X1 U5010 ( .A1(n6007), .A2(n6006), .ZN(n7994) );
  XNOR2_X1 U5011 ( .A(n5496), .B(n5495), .ZN(n7204) );
  NOR2_X1 U5012 ( .A1(n6904), .A2(n6901), .ZN(n7358) );
  NAND2_X1 U5013 ( .A1(n5494), .A2(n5493), .ZN(n5496) );
  NAND2_X1 U5014 ( .A1(n5996), .A2(n5995), .ZN(n10227) );
  NAND2_X1 U5015 ( .A1(n10058), .A2(n10050), .ZN(n9496) );
  INV_X2 U5016 ( .A(n6897), .ZN(n7045) );
  NAND2_X1 U5017 ( .A1(n5406), .A2(n5405), .ZN(n7780) );
  OR2_X1 U5018 ( .A1(n10064), .A2(n10334), .ZN(n10033) );
  AND2_X1 U5019 ( .A1(n5422), .A2(n5421), .ZN(n7814) );
  INV_X1 U5020 ( .A(n10058), .ZN(n10018) );
  XNOR2_X1 U5021 ( .A(n5390), .B(n5389), .ZN(n7144) );
  INV_X1 U5022 ( .A(n10073), .ZN(n9569) );
  INV_X1 U5023 ( .A(n7329), .ZN(n6771) );
  INV_X1 U5024 ( .A(n7348), .ZN(n8303) );
  NAND2_X1 U5025 ( .A1(n6378), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U5026 ( .A1(n5279), .A2(n5280), .ZN(n7475) );
  AND4_X1 U5027 ( .A1(n6327), .A2(n6326), .A3(n6325), .A4(n6324), .ZN(n10043)
         );
  NAND4_X1 U5028 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), .ZN(n8302)
         );
  NOR2_X1 U5029 ( .A1(n5286), .A2(n4444), .ZN(n7337) );
  AND4_X1 U5030 ( .A1(n5319), .A2(n5318), .A3(n5317), .A4(n5316), .ZN(n7329)
         );
  INV_X4 U5031 ( .A(n7070), .ZN(n7002) );
  NAND4_X2 U5032 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(n10364)
         );
  INV_X2 U5033 ( .A(n6207), .ZN(n6564) );
  NAND2_X2 U5034 ( .A1(n6200), .A2(n6201), .ZN(n6846) );
  CLKBUF_X1 U5035 ( .A(n6886), .Z(n7175) );
  NAND2_X1 U5036 ( .A1(n6574), .A2(n7152), .ZN(n7450) );
  MUX2_X1 U5037 ( .A(n10448), .B(n8813), .S(n6207), .Z(n10472) );
  NAND2_X2 U5038 ( .A1(n6121), .A2(n6120), .ZN(n6886) );
  AND2_X1 U5039 ( .A1(n7690), .A2(n7503), .ZN(n6225) );
  INV_X4 U5040 ( .A(n5315), .ZN(n5752) );
  NAND3_X2 U5041 ( .A1(n5947), .A2(n5946), .A3(n5945), .ZN(n7518) );
  INV_X2 U5042 ( .A(n9315), .ZN(n4380) );
  BUF_X2 U5044 ( .A(n5288), .Z(n6207) );
  INV_X2 U5045 ( .A(n6303), .ZN(n6413) );
  NAND2_X1 U5046 ( .A1(n6708), .A2(n4382), .ZN(n5288) );
  INV_X2 U5047 ( .A(n6436), .ZN(n4381) );
  XNOR2_X1 U5048 ( .A(n5916), .B(n5915), .ZN(n6216) );
  NOR2_X1 U5049 ( .A1(n6122), .A2(n7975), .ZN(n6120) );
  NAND2_X1 U5050 ( .A1(n4845), .A2(n5918), .ZN(n6214) );
  NAND2_X1 U5051 ( .A1(n5809), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5231) );
  XNOR2_X1 U5052 ( .A(n6110), .B(n6109), .ZN(n6125) );
  NAND2_X1 U5053 ( .A1(n8007), .A2(n6246), .ZN(n6265) );
  AND2_X1 U5054 ( .A1(n6245), .A2(n6091), .ZN(n6374) );
  NAND2_X1 U5055 ( .A1(n6113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6110) );
  MUX2_X1 U5056 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6112), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6114) );
  OAI21_X1 U5057 ( .B1(n5923), .B2(n5180), .A(n4403), .ZN(n4780) );
  INV_X1 U5058 ( .A(n6123), .ZN(n7975) );
  XNOR2_X1 U5059 ( .A(n6100), .B(n6105), .ZN(n7732) );
  XNOR2_X1 U5060 ( .A(n6087), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U5061 ( .A1(n5187), .A2(n5186), .ZN(n5549) );
  XNOR2_X1 U5062 ( .A(n6083), .B(n9087), .ZN(n9539) );
  NAND2_X1 U5063 ( .A1(n5034), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6030) );
  XNOR2_X1 U5064 ( .A(n5350), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6631) );
  XNOR2_X1 U5065 ( .A(n4604), .B(n5932), .ZN(n6096) );
  MUX2_X1 U5066 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5930), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5931) );
  NAND2_X1 U5067 ( .A1(n6106), .A2(n5078), .ZN(n6111) );
  NAND2_X1 U5068 ( .A1(n10279), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6087) );
  OR2_X1 U5069 ( .A1(n6117), .A2(n10278), .ZN(n4604) );
  NAND2_X1 U5070 ( .A1(n6117), .A2(n4777), .ZN(n10279) );
  NAND2_X1 U5071 ( .A1(n6285), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6305) );
  NAND3_X1 U5072 ( .A1(n5092), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4804) );
  AND2_X1 U5073 ( .A1(n4654), .A2(n4653), .ZN(n4854) );
  NAND2_X1 U5074 ( .A1(n4650), .A2(n4651), .ZN(n4652) );
  AND4_X1 U5075 ( .A1(n5215), .A2(n5213), .A3(n5170), .A4(n5169), .ZN(n5171)
         );
  NOR2_X1 U5076 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4890) );
  INV_X1 U5077 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6031) );
  INV_X1 U5078 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5035) );
  NOR2_X1 U5079 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4889) );
  INV_X2 U5080 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8934) );
  NOR2_X1 U5081 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4689) );
  NOR2_X1 U5082 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4690) );
  NOR2_X1 U5083 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4748) );
  BUF_X1 U5084 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n10448) );
  INV_X1 U5085 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9055) );
  INV_X1 U5086 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6040) );
  INV_X4 U5087 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X4 U5088 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5089 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4651) );
  NOR2_X1 U5090 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4653) );
  NOR2_X1 U5091 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4654) );
  NOR2_X1 U5092 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5174) );
  INV_X1 U5093 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5182) );
  INV_X1 U5094 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5915) );
  INV_X1 U5095 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5241) );
  INV_X1 U5096 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5213) );
  INV_X1 U5097 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5215) );
  NOR2_X1 U5098 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5172) );
  INV_X1 U5099 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5217) );
  INV_X1 U5100 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5220) );
  INV_X1 U5101 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5186) );
  NOR2_X1 U5102 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5168) );
  NOR2_X1 U5103 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4888) );
  AOI21_X2 U5104 ( .B1(n8125), .B2(n4850), .A(n4847), .ZN(n4846) );
  NAND2_X2 U5105 ( .A1(n6792), .A2(n6791), .ZN(n8125) );
  BUF_X1 U5106 ( .A(n10445), .Z(n4382) );
  BUF_X8 U5107 ( .A(n10445), .Z(n4383) );
  NAND2_X2 U5108 ( .A1(n4780), .A2(n5181), .ZN(n10445) );
  INV_X1 U5109 ( .A(n9729), .ZN(n6450) );
  NAND2_X1 U5110 ( .A1(n5288), .A2(n5936), .ZN(n5325) );
  OR2_X2 U5111 ( .A1(n8801), .A2(n5207), .ZN(n5298) );
  NAND2_X2 U5112 ( .A1(n9926), .A2(n9370), .ZN(n9911) );
  AND2_X1 U5113 ( .A1(n6246), .A2(n6245), .ZN(n6263) );
  INV_X2 U5114 ( .A(n6380), .ZN(n6404) );
  INV_X2 U5115 ( .A(n6380), .ZN(n6541) );
  INV_X2 U5116 ( .A(n6374), .ZN(n6380) );
  OR2_X1 U5117 ( .A1(n6074), .A2(n7131), .ZN(n5947) );
  OR2_X1 U5118 ( .A1(n6067), .A2(n7155), .ZN(n5945) );
  INV_X2 U5119 ( .A(n6390), .ZN(n6403) );
  NAND2_X1 U5120 ( .A1(n6091), .A2(n8007), .ZN(n6259) );
  INV_X1 U5121 ( .A(n6265), .ZN(n6274) );
  AOI21_X2 U5122 ( .B1(n8857), .B2(n4442), .A(n5044), .ZN(n5043) );
  XNOR2_X2 U5123 ( .A(n5193), .B(n5192), .ZN(n8801) );
  INV_X2 U5124 ( .A(n9480), .ZN(n9572) );
  BUF_X2 U5125 ( .A(n6074), .Z(n4385) );
  NAND2_X1 U5126 ( .A1(n4374), .A2(n7132), .ZN(n6074) );
  NAND2_X2 U5127 ( .A1(n5989), .A2(n5988), .ZN(n10050) );
  NOR2_X2 U5128 ( .A1(n5086), .A2(n6556), .ZN(n9712) );
  NAND2_X1 U5129 ( .A1(n4374), .A2(n5936), .ZN(n4387) );
  INV_X1 U5130 ( .A(n6303), .ZN(n4388) );
  INV_X2 U5131 ( .A(n6303), .ZN(n4389) );
  NAND2_X1 U5132 ( .A1(n4375), .A2(n7132), .ZN(n4390) );
  INV_X4 U5133 ( .A(n4391), .ZN(n10122) );
  OAI222_X1 U5134 ( .A1(P1_U3086), .A2(n7228), .B1(n8004), .B2(n7172), .C1(
        n7171), .C2(n8105), .ZN(P1_U3354) );
  OAI222_X1 U5135 ( .A1(P1_U3086), .A2(n6125), .B1(n8004), .B2(n8010), .C1(
        n9063), .C2(n8105), .ZN(P1_U3330) );
  INV_X2 U5136 ( .A(n10281), .ZN(n8105) );
  INV_X1 U5137 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U5138 ( .A1(n4498), .A2(n4380), .ZN(n4760) );
  NAND2_X1 U5139 ( .A1(n4537), .A2(n4536), .ZN(n9417) );
  AND2_X1 U5140 ( .A1(n9469), .A2(n4469), .ZN(n4536) );
  AOI21_X1 U5141 ( .B1(n4680), .B2(n4681), .A(n4678), .ZN(n4677) );
  INV_X1 U5142 ( .A(n6146), .ZN(n4678) );
  AND2_X1 U5143 ( .A1(n8801), .A2(n5207), .ZN(n5264) );
  OR2_X1 U5144 ( .A1(n5785), .A2(n8422), .ZN(n6146) );
  OR2_X1 U5145 ( .A1(n8772), .A2(n8557), .ZN(n5876) );
  NAND2_X1 U5146 ( .A1(n6514), .A2(n6513), .ZN(n4949) );
  AOI21_X1 U5147 ( .B1(n4956), .B2(n4959), .A(n4955), .ZN(n4954) );
  NOR2_X1 U5148 ( .A1(n8821), .A2(n9732), .ZN(n4955) );
  INV_X1 U5149 ( .A(n5048), .ZN(n5047) );
  OAI21_X1 U5150 ( .B1(n5049), .B2(n5051), .A(n7020), .ZN(n5048) );
  NAND2_X1 U5151 ( .A1(n4375), .A2(n5936), .ZN(n6067) );
  AND2_X1 U5152 ( .A1(n4472), .A2(n5580), .ZN(n4784) );
  AND2_X1 U5153 ( .A1(n4841), .A2(n4840), .ZN(n4839) );
  INV_X1 U5154 ( .A(n5607), .ZN(n4840) );
  INV_X1 U5155 ( .A(n4418), .ZN(n5056) );
  INV_X1 U5156 ( .A(n4826), .ZN(n4825) );
  OAI21_X1 U5157 ( .B1(n5714), .B2(n4827), .A(n5722), .ZN(n4826) );
  AND2_X1 U5158 ( .A1(n5154), .A2(n5513), .ZN(n4596) );
  INV_X1 U5159 ( .A(n5400), .ZN(n5386) );
  NAND2_X1 U5160 ( .A1(n5121), .A2(n7170), .ZN(n4550) );
  OAI21_X1 U5161 ( .B1(n5121), .B2(n4569), .A(n4568), .ZN(n5108) );
  NAND2_X1 U5162 ( .A1(n5121), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4568) );
  OAI211_X1 U5163 ( .C1(n4812), .C2(n4459), .A(n4808), .B(n5781), .ZN(n5784)
         );
  NAND2_X1 U5164 ( .A1(n4809), .A2(n8092), .ZN(n4808) );
  NAND2_X1 U5165 ( .A1(n4711), .A2(n6594), .ZN(n6595) );
  NAND2_X1 U5166 ( .A1(n4549), .A2(n7400), .ZN(n4901) );
  INV_X1 U5167 ( .A(n6574), .ZN(n4549) );
  OR2_X1 U5168 ( .A1(n5298), .A2(n7473), .ZN(n5267) );
  INV_X1 U5169 ( .A(n6194), .ZN(n4996) );
  INV_X1 U5170 ( .A(n5886), .ZN(n4738) );
  OR2_X1 U5171 ( .A1(n8499), .A2(n8483), .ZN(n5884) );
  OR2_X1 U5172 ( .A1(n8755), .A2(n8214), .ZN(n5881) );
  OR2_X1 U5173 ( .A1(n7700), .A2(n7512), .ZN(n5854) );
  INV_X1 U5174 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4855) );
  INV_X2 U5175 ( .A(n4652), .ZN(n5308) );
  NAND2_X1 U5176 ( .A1(n6936), .A2(n5068), .ZN(n5067) );
  INV_X1 U5177 ( .A(n6937), .ZN(n5068) );
  NAND2_X1 U5178 ( .A1(n9743), .A2(n9457), .ZN(n9729) );
  AOI21_X1 U5179 ( .B1(n9910), .B2(n6497), .A(n4937), .ZN(n4936) );
  INV_X1 U5180 ( .A(n6498), .ZN(n4937) );
  NAND2_X1 U5181 ( .A1(n6480), .A2(n4609), .ZN(n4608) );
  NOR2_X1 U5182 ( .A1(n9749), .A2(n9735), .ZN(n6521) );
  AND2_X1 U5183 ( .A1(n5685), .A2(n5672), .ZN(n5683) );
  NAND2_X1 U5184 ( .A1(n4843), .A2(n4833), .ZN(n4834) );
  INV_X1 U5185 ( .A(n5525), .ZN(n5159) );
  OR2_X1 U5186 ( .A1(n6000), .A2(n5999), .ZN(n6003) );
  INV_X1 U5187 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5998) );
  NOR4_X1 U5188 ( .A1(n5898), .A2(n5839), .A3(n5838), .A4(n5837), .ZN(n5906)
         );
  OR2_X1 U5189 ( .A1(n6237), .A2(n5733), .ZN(n5805) );
  INV_X1 U5190 ( .A(n5733), .ZN(n5751) );
  OAI211_X1 U5191 ( .C1(n5336), .C2(n5282), .A(n5284), .B(n5285), .ZN(n5286)
         );
  NAND2_X1 U5192 ( .A1(n4634), .A2(n8393), .ZN(n8392) );
  OR2_X1 U5193 ( .A1(n5707), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5749) );
  INV_X1 U5194 ( .A(n8296), .ZN(n8556) );
  AND2_X1 U5195 ( .A1(n5288), .A2(n7132), .ZN(n5305) );
  OR2_X1 U5196 ( .A1(n7122), .A2(n6235), .ZN(n6238) );
  NAND2_X1 U5197 ( .A1(n4915), .A2(n5895), .ZN(n8428) );
  AND2_X1 U5198 ( .A1(n4741), .A2(n4482), .ZN(n4736) );
  AOI21_X1 U5199 ( .B1(n4980), .B2(n4976), .A(n4975), .ZN(n4974) );
  NOR2_X1 U5200 ( .A1(n8123), .A2(n8484), .ZN(n4975) );
  NAND2_X1 U5201 ( .A1(n4424), .A2(n4737), .ZN(n4741) );
  NOR2_X1 U5202 ( .A1(n8485), .A2(n4738), .ZN(n4737) );
  OR2_X1 U5203 ( .A1(n6846), .A2(n6871), .ZN(n8694) );
  AOI21_X1 U5204 ( .B1(n4985), .B2(n4983), .A(n4456), .ZN(n4982) );
  INV_X1 U5205 ( .A(n4985), .ZN(n4984) );
  AOI21_X1 U5206 ( .B1(n4430), .B2(n4663), .A(n4659), .ZN(n4658) );
  INV_X1 U5207 ( .A(n5874), .ZN(n4663) );
  NAND2_X1 U5208 ( .A1(n6202), .A2(n6742), .ZN(n8696) );
  XNOR2_X1 U5209 ( .A(n6214), .B(P2_B_REG_SCAN_IN), .ZN(n6215) );
  NAND2_X1 U5210 ( .A1(n5178), .A2(n5180), .ZN(n4939) );
  NAND2_X1 U5211 ( .A1(n5913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U5212 ( .A1(n4858), .A2(n4856), .ZN(n5913) );
  INV_X1 U5213 ( .A(n4857), .ZN(n4856) );
  INV_X1 U5214 ( .A(n6441), .ZN(n6431) );
  NAND2_X1 U5215 ( .A1(n5047), .A2(n4433), .ZN(n5045) );
  NAND2_X1 U5216 ( .A1(n8883), .A2(n5041), .ZN(n5040) );
  INV_X1 U5217 ( .A(n7040), .ZN(n5041) );
  INV_X1 U5218 ( .A(n4948), .ZN(n4947) );
  NOR2_X1 U5219 ( .A1(n4957), .A2(n4952), .ZN(n4951) );
  NAND2_X1 U5220 ( .A1(n9870), .A2(n6501), .ZN(n4935) );
  OR2_X1 U5221 ( .A1(n7994), .A2(n9968), .ZN(n9360) );
  NAND2_X1 U5222 ( .A1(n6070), .A2(n6069), .ZN(n6556) );
  NAND2_X1 U5223 ( .A1(n6068), .A2(n5983), .ZN(n6070) );
  NAND3_X1 U5224 ( .A1(n9548), .A2(n7175), .A3(P1_STATE_REG_SCAN_IN), .ZN(
        n7190) );
  INV_X1 U5225 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4887) );
  INV_X1 U5226 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5027) );
  XNOR2_X1 U5227 ( .A(n6147), .B(n6197), .ZN(n6737) );
  OAI21_X1 U5228 ( .B1(n8428), .B2(n4681), .A(n4680), .ZN(n6147) );
  XNOR2_X1 U5229 ( .A(n6548), .B(n4958), .ZN(n9725) );
  NAND2_X1 U5230 ( .A1(n4953), .A2(n4959), .ZN(n6548) );
  NAND2_X1 U5231 ( .A1(n9742), .A2(n4962), .ZN(n4953) );
  OAI22_X1 U5232 ( .A1(n8818), .A2(n6461), .B1(n9402), .B2(n6460), .ZN(n6462)
         );
  NAND2_X1 U5233 ( .A1(n9345), .A2(n4380), .ZN(n4757) );
  NAND3_X1 U5234 ( .A1(n6318), .A2(n9315), .A3(n10034), .ZN(n4754) );
  NAND3_X1 U5235 ( .A1(n4756), .A2(n4458), .A3(n4380), .ZN(n4753) );
  INV_X1 U5236 ( .A(n9345), .ZN(n4756) );
  NAND2_X1 U5237 ( .A1(n4776), .A2(n9513), .ZN(n4771) );
  INV_X1 U5238 ( .A(n5486), .ZN(n4507) );
  NAND2_X1 U5239 ( .A1(n4776), .A2(n4432), .ZN(n4774) );
  NOR2_X1 U5240 ( .A1(n4447), .A2(n4771), .ZN(n4770) );
  NOR2_X1 U5241 ( .A1(n4773), .A2(n4447), .ZN(n4769) );
  AND2_X1 U5242 ( .A1(n5881), .A2(n8521), .ZN(n4788) );
  NAND2_X1 U5243 ( .A1(n4781), .A2(n4450), .ZN(n4783) );
  NAND2_X1 U5244 ( .A1(n5563), .A2(n4786), .ZN(n4781) );
  NAND2_X1 U5245 ( .A1(n4786), .A2(n6846), .ZN(n4598) );
  INV_X1 U5246 ( .A(n8447), .ZN(n4791) );
  NOR2_X1 U5247 ( .A1(n4593), .A2(n4454), .ZN(n4592) );
  NAND2_X1 U5248 ( .A1(n6318), .A2(n4401), .ZN(n9497) );
  NOR2_X1 U5249 ( .A1(n4893), .A2(n9767), .ZN(n4892) );
  NAND2_X1 U5250 ( .A1(n10249), .A2(n10253), .ZN(n4893) );
  AOI21_X1 U5251 ( .B1(n4839), .B2(n4837), .A(n4836), .ZN(n4835) );
  INV_X1 U5252 ( .A(n5606), .ZN(n4836) );
  INV_X1 U5253 ( .A(n4839), .ZN(n4838) );
  NAND2_X1 U5254 ( .A1(n5210), .A2(n5167), .ZN(n4830) );
  NOR2_X1 U5255 ( .A1(n4838), .A2(n4833), .ZN(n4832) );
  NAND2_X1 U5256 ( .A1(n5546), .A2(n5545), .ZN(n5564) );
  INV_X1 U5257 ( .A(n5540), .ZN(n5543) );
  NAND2_X1 U5258 ( .A1(n5145), .A2(n5144), .ZN(n5152) );
  NAND2_X1 U5259 ( .A1(n5150), .A2(n5471), .ZN(n5487) );
  NOR2_X1 U5260 ( .A1(n5252), .A2(n4817), .ZN(n4816) );
  INV_X1 U5261 ( .A(n5134), .ZN(n4817) );
  NAND2_X1 U5262 ( .A1(n7561), .A2(n4438), .ZN(n6572) );
  NAND2_X1 U5263 ( .A1(n7621), .A2(n6573), .ZN(n6574) );
  AOI21_X1 U5264 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7737), .A(n7738), .ZN(
        n6578) );
  INV_X1 U5265 ( .A(n7736), .ZN(n4734) );
  NAND2_X1 U5266 ( .A1(n4407), .A2(n4649), .ZN(n4645) );
  NAND2_X1 U5267 ( .A1(n4647), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U5268 ( .A1(n8324), .A2(n6579), .ZN(n6580) );
  AND2_X1 U5269 ( .A1(n5654), .A2(n4700), .ZN(n4699) );
  INV_X1 U5270 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n4700) );
  INV_X1 U5271 ( .A(n5656), .ZN(n5655) );
  AND2_X1 U5272 ( .A1(n5203), .A2(n4707), .ZN(n4706) );
  INV_X1 U5273 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n4707) );
  INV_X1 U5274 ( .A(n5518), .ZN(n5204) );
  AND2_X1 U5275 ( .A1(n7668), .A2(n5450), .ZN(n7696) );
  INV_X1 U5276 ( .A(n5853), .ZN(n4927) );
  NAND2_X1 U5277 ( .A1(n7495), .A2(n7440), .ZN(n5852) );
  NAND2_X1 U5278 ( .A1(n6761), .A2(n6150), .ZN(n5846) );
  OAI211_X1 U5279 ( .C1(n6567), .C2(n6207), .A(n4528), .B(n4664), .ZN(n5311)
         );
  NAND2_X1 U5280 ( .A1(n4529), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4528) );
  NAND2_X1 U5281 ( .A1(n8306), .A2(n10472), .ZN(n7412) );
  NAND2_X1 U5282 ( .A1(n4993), .A2(n6196), .ZN(n4992) );
  INV_X1 U5283 ( .A(n4999), .ZN(n4993) );
  OR2_X1 U5284 ( .A1(n8728), .A2(n8275), .ZN(n5892) );
  AND2_X1 U5285 ( .A1(n4980), .A2(n4979), .ZN(n4978) );
  INV_X1 U5286 ( .A(n6191), .ZN(n4979) );
  OR2_X1 U5287 ( .A1(n8734), .A2(n8119), .ZN(n5889) );
  OR2_X1 U5288 ( .A1(n8740), .A2(n8484), .ZN(n5887) );
  CLKBUF_X1 U5289 ( .A(n8030), .Z(n8031) );
  NAND2_X1 U5290 ( .A1(n7507), .A2(n7506), .ZN(n4969) );
  OR2_X1 U5291 ( .A1(n8299), .A2(n7780), .ZN(n6164) );
  INV_X1 U5292 ( .A(n7431), .ZN(n7344) );
  INV_X1 U5293 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U5294 ( .A1(n6933), .A2(n5069), .ZN(n5065) );
  INV_X1 U5295 ( .A(n5053), .ZN(n5052) );
  OAI21_X1 U5296 ( .B1(n5057), .B2(n4452), .A(n5054), .ZN(n5053) );
  NOR2_X1 U5297 ( .A1(n4418), .A2(n5058), .ZN(n5057) );
  INV_X1 U5298 ( .A(n6947), .ZN(n5066) );
  INV_X1 U5299 ( .A(n6948), .ZN(n5064) );
  NOR2_X1 U5300 ( .A1(n9924), .A2(n4520), .ZN(n4519) );
  AND2_X1 U5301 ( .A1(n9551), .A2(n9539), .ZN(n6881) );
  INV_X1 U5302 ( .A(n9422), .ZN(n4765) );
  NAND2_X1 U5303 ( .A1(n4958), .A2(n9524), .ZN(n5008) );
  INV_X1 U5304 ( .A(n5010), .ZN(n5009) );
  OAI21_X1 U5305 ( .B1(n6449), .B2(n5011), .A(n9444), .ZN(n5010) );
  OR2_X1 U5306 ( .A1(n9787), .A2(n9803), .ZN(n6511) );
  NOR2_X1 U5307 ( .A1(n6512), .A2(n4628), .ZN(n4627) );
  INV_X1 U5308 ( .A(n6509), .ZN(n4628) );
  OR2_X1 U5309 ( .A1(n9767), .A2(n6429), .ZN(n9454) );
  NAND2_X1 U5310 ( .A1(n9800), .A2(n9310), .ZN(n9777) );
  OR2_X1 U5311 ( .A1(n10271), .A2(n9894), .ZN(n9514) );
  INV_X1 U5312 ( .A(n4931), .ZN(n4930) );
  OAI21_X1 U5313 ( .B1(n9965), .B2(n4932), .A(n6494), .ZN(n4931) );
  INV_X1 U5314 ( .A(n6493), .ZN(n4932) );
  INV_X1 U5315 ( .A(n9360), .ZN(n5021) );
  NAND2_X1 U5316 ( .A1(n9557), .A2(n9551), .ZN(n6884) );
  NAND2_X1 U5317 ( .A1(n6127), .A2(n6126), .ZN(n6129) );
  NAND2_X1 U5318 ( .A1(n5768), .A2(n5767), .ZN(n5793) );
  NAND2_X1 U5319 ( .A1(n4820), .A2(SI_29_), .ZN(n5768) );
  AOI21_X1 U5320 ( .B1(n4825), .B2(n4827), .A(n4823), .ZN(n4822) );
  INV_X1 U5321 ( .A(n5724), .ZN(n4823) );
  AND2_X1 U5322 ( .A1(n5667), .A2(n5651), .ZN(n5665) );
  NAND2_X1 U5323 ( .A1(n6080), .A2(n5035), .ZN(n5034) );
  XNOR2_X1 U5324 ( .A(n5160), .B(SI_16_), .ZN(n5525) );
  NAND2_X1 U5325 ( .A1(n4595), .A2(n5158), .ZN(n5526) );
  XNOR2_X1 U5326 ( .A(n5151), .B(SI_13_), .ZN(n5471) );
  OR2_X1 U5327 ( .A1(n5127), .A2(n5387), .ZN(n5129) );
  OR2_X1 U5328 ( .A1(n5378), .A2(n5110), .ZN(n5111) );
  INV_X1 U5329 ( .A(n4851), .ZN(n4850) );
  OAI21_X1 U5330 ( .B1(n4852), .B2(n6796), .A(n8219), .ZN(n4851) );
  INV_X1 U5331 ( .A(n6808), .ZN(n4866) );
  NAND2_X1 U5332 ( .A1(n5200), .A2(n4428), .ZN(n5257) );
  NAND2_X1 U5333 ( .A1(n8187), .A2(n4494), .ZN(n8190) );
  NAND2_X1 U5334 ( .A1(n4464), .A2(n6788), .ZN(n4874) );
  AOI21_X1 U5335 ( .B1(n4873), .B2(n7714), .A(n4872), .ZN(n4871) );
  NOR2_X1 U5336 ( .A1(n7771), .A2(n7770), .ZN(n4872) );
  INV_X1 U5337 ( .A(n4874), .ZN(n4873) );
  NAND2_X1 U5338 ( .A1(n7435), .A2(n7434), .ZN(n4862) );
  AND2_X1 U5339 ( .A1(n4504), .A2(n5790), .ZN(n5806) );
  OR2_X1 U5340 ( .A1(n5297), .A2(n5296), .ZN(n5303) );
  OAI21_X1 U5341 ( .B1(n7385), .B2(n10451), .A(n6626), .ZN(n7570) );
  XNOR2_X1 U5342 ( .A(n6567), .B(n6588), .ZN(n7564) );
  AOI21_X1 U5343 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n7149), .A(n7449), .ZN(
        n6575) );
  NAND2_X1 U5344 ( .A1(n7909), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U5345 ( .A1(n6580), .A2(n8348), .ZN(n6581) );
  OR2_X1 U5346 ( .A1(n6619), .A2(n6620), .ZN(n6616) );
  INV_X1 U5347 ( .A(n4725), .ZN(n4724) );
  NAND2_X1 U5348 ( .A1(n8406), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U5349 ( .A1(n5732), .A2(n5731), .ZN(n6237) );
  NAND2_X1 U5350 ( .A1(n5655), .A2(n5654), .ZN(n5675) );
  NOR2_X1 U5351 ( .A1(n4738), .A2(n5882), .ZN(n4942) );
  INV_X1 U5352 ( .A(n5885), .ZN(n4521) );
  NOR2_X1 U5353 ( .A1(n8500), .A2(n4743), .ZN(n4742) );
  INV_X1 U5354 ( .A(n5881), .ZN(n4743) );
  OR2_X1 U5355 ( .A1(n5226), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5554) );
  OR2_X1 U5356 ( .A1(n7868), .A2(n7776), .ZN(n8597) );
  OR2_X1 U5357 ( .A1(n5425), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U5358 ( .A1(n5200), .A2(n5199), .ZN(n5444) );
  INV_X1 U5359 ( .A(n4672), .ZN(n4671) );
  NOR2_X1 U5360 ( .A1(n4675), .A2(n4676), .ZN(n4674) );
  INV_X1 U5361 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5196) );
  INV_X1 U5362 ( .A(n5311), .ZN(n7328) );
  XNOR2_X1 U5363 ( .A(n8711), .B(n8432), .ZN(n8420) );
  NAND2_X1 U5364 ( .A1(n5896), .A2(n5719), .ZN(n8430) );
  NAND2_X1 U5365 ( .A1(n4997), .A2(n6194), .ZN(n8439) );
  NAND2_X1 U5366 ( .A1(n8440), .A2(n8692), .ZN(n4546) );
  AND2_X1 U5367 ( .A1(n8493), .A2(n5079), .ZN(n6187) );
  NAND2_X1 U5368 ( .A1(n5879), .A2(n4670), .ZN(n4740) );
  INV_X1 U5369 ( .A(n4667), .ZN(n4670) );
  NAND2_X1 U5370 ( .A1(n5613), .A2(n5612), .ZN(n8230) );
  AND2_X1 U5371 ( .A1(n5881), .A2(n5880), .ZN(n8512) );
  INV_X1 U5372 ( .A(n6178), .ZN(n4988) );
  AND2_X1 U5373 ( .A1(n5876), .A2(n5875), .ZN(n8545) );
  NAND2_X1 U5374 ( .A1(n5872), .A2(n5871), .ZN(n8561) );
  NOR2_X1 U5375 ( .A1(n5870), .A2(n5507), .ZN(n4945) );
  OR2_X1 U5376 ( .A1(n5509), .A2(n5870), .ZN(n8575) );
  INV_X1 U5377 ( .A(n8694), .ZN(n8609) );
  NAND2_X1 U5378 ( .A1(n7787), .A2(n7730), .ZN(n10488) );
  NOR2_X1 U5379 ( .A1(n7119), .A2(n6741), .ZN(n6865) );
  OR2_X1 U5380 ( .A1(n6743), .A2(n6200), .ZN(n6848) );
  INV_X1 U5381 ( .A(n8696), .ZN(n10469) );
  AND2_X1 U5382 ( .A1(n6861), .A2(n7195), .ZN(n7160) );
  INV_X1 U5383 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U5384 ( .A1(n5917), .A2(n5914), .ZN(n5918) );
  NAND3_X1 U5385 ( .A1(n5235), .A2(n5234), .A3(n5233), .ZN(n5237) );
  NAND2_X1 U5386 ( .A1(n4860), .A2(n5238), .ZN(n5840) );
  INV_X1 U5387 ( .A(n5237), .ZN(n4860) );
  BUF_X1 U5388 ( .A(n6754), .Z(n6200) );
  NAND2_X1 U5389 ( .A1(n4652), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U5390 ( .A1(n9241), .A2(n4426), .ZN(n8825) );
  INV_X1 U5391 ( .A(n6934), .ZN(n7073) );
  AND2_X1 U5392 ( .A1(n7060), .A2(n7059), .ZN(n7085) );
  NAND2_X1 U5393 ( .A1(n6411), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6421) );
  INV_X1 U5394 ( .A(n4576), .ZN(n6430) );
  NAND2_X1 U5395 ( .A1(n6356), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6363) );
  INV_X1 U5396 ( .A(n9471), .ZN(n4579) );
  AND2_X1 U5397 ( .A1(n9557), .A2(n6518), .ZN(n9472) );
  NOR2_X1 U5398 ( .A1(n9535), .A2(n4581), .ZN(n4580) );
  NOR2_X1 U5399 ( .A1(n10236), .A2(n9562), .ZN(n4581) );
  OAI21_X1 U5400 ( .B1(n9531), .B2(n4584), .A(n4583), .ZN(n4582) );
  INV_X1 U5401 ( .A(n9533), .ZN(n4583) );
  INV_X1 U5402 ( .A(n6881), .ZN(n5033) );
  AND4_X1 U5403 ( .A1(n6252), .A2(n6251), .A3(n6250), .A4(n6249), .ZN(n7104)
         );
  AOI21_X1 U5404 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n10293), .A(n10296), .ZN(
        n8048) );
  OR2_X1 U5405 ( .A1(n7106), .A2(n8818), .ZN(n9449) );
  AND2_X1 U5406 ( .A1(n9449), .A2(n9412), .ZN(n6722) );
  INV_X1 U5407 ( .A(n4960), .ZN(n4959) );
  OAI21_X1 U5408 ( .B1(n6517), .B2(n4961), .A(n6516), .ZN(n4960) );
  NAND2_X1 U5409 ( .A1(n6515), .A2(n4964), .ZN(n4961) );
  AND2_X1 U5410 ( .A1(n6444), .A2(n6443), .ZN(n9736) );
  NAND2_X1 U5411 ( .A1(n6441), .A2(n6442), .ZN(n6444) );
  NAND2_X1 U5412 ( .A1(n4622), .A2(n4620), .ZN(n9742) );
  AOI21_X1 U5413 ( .B1(n4623), .B2(n4621), .A(n4952), .ZN(n4620) );
  OR2_X1 U5414 ( .A1(n6510), .A2(n4624), .ZN(n4622) );
  INV_X1 U5415 ( .A(n4627), .ZN(n4621) );
  NAND2_X1 U5416 ( .A1(n9779), .A2(n9451), .ZN(n9760) );
  NAND2_X1 U5417 ( .A1(n9819), .A2(n9523), .ZN(n9799) );
  AND2_X1 U5418 ( .A1(n9380), .A2(n9520), .ZN(n9857) );
  NAND2_X1 U5419 ( .A1(n4615), .A2(n4613), .ZN(n6500) );
  AND2_X1 U5420 ( .A1(n4936), .A2(n4614), .ZN(n4613) );
  OR2_X2 U5421 ( .A1(n10197), .A2(n9877), .ZN(n9871) );
  NAND2_X1 U5422 ( .A1(n4616), .A2(n6495), .ZN(n9903) );
  NAND2_X1 U5423 ( .A1(n9922), .A2(n9924), .ZN(n4616) );
  OR2_X1 U5424 ( .A1(n9903), .A2(n9910), .ZN(n9905) );
  NAND2_X1 U5425 ( .A1(n4577), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U5426 ( .A1(n7997), .A2(n9439), .ZN(n5025) );
  CLKBUF_X1 U5427 ( .A(n7996), .Z(n7997) );
  NAND2_X1 U5428 ( .A1(n4608), .A2(n4607), .ZN(n6482) );
  INV_X1 U5429 ( .A(n4606), .ZN(n4607) );
  AOI21_X1 U5430 ( .B1(n10366), .B2(n9320), .A(n6476), .ZN(n6477) );
  NAND2_X1 U5431 ( .A1(n6060), .A2(n6059), .ZN(n10153) );
  NAND2_X1 U5432 ( .A1(n6049), .A2(n6048), .ZN(n9864) );
  OAI211_X1 U5433 ( .C1(n7173), .C2(n7228), .A(n5938), .B(n5937), .ZN(n6467)
         );
  OR2_X1 U5434 ( .A1(n4387), .A2(n7172), .ZN(n5937) );
  OR2_X1 U5435 ( .A1(n4390), .A2(n7171), .ZN(n5938) );
  AND2_X1 U5436 ( .A1(n10133), .A2(n5033), .ZN(n10228) );
  AND2_X1 U5437 ( .A1(n7732), .A2(n9431), .ZN(n10133) );
  AND2_X1 U5438 ( .A1(n5646), .A2(n5634), .ZN(n5644) );
  XNOR2_X1 U5439 ( .A(n5586), .B(n5585), .ZN(n7786) );
  INV_X1 U5440 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6011) );
  NOR2_X1 U5441 ( .A1(n6003), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6012) );
  OR2_X1 U5442 ( .A1(n5121), .A2(n4437), .ZN(n4559) );
  NOR2_X2 U5443 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5943) );
  AND2_X1 U5444 ( .A1(n8093), .A2(n8271), .ZN(n4523) );
  AND2_X1 U5445 ( .A1(n5620), .A2(n5619), .ZN(n8496) );
  AND4_X1 U5446 ( .A1(n5373), .A2(n5372), .A3(n5371), .A4(n5370), .ZN(n7700)
         );
  INV_X1 U5447 ( .A(n8302), .ZN(n7495) );
  AND3_X1 U5448 ( .A1(n5229), .A2(n5228), .A3(n5227), .ZN(n8261) );
  AND2_X1 U5449 ( .A1(n7489), .A2(n10473), .ZN(n8263) );
  AND2_X1 U5450 ( .A1(n5704), .A2(n5703), .ZN(n8421) );
  INV_X1 U5451 ( .A(n7730), .ZN(n6201) );
  INV_X1 U5452 ( .A(n8090), .ZN(n8432) );
  INV_X1 U5453 ( .A(n8421), .ZN(n8440) );
  NAND2_X1 U5454 ( .A1(n5712), .A2(n5711), .ZN(n8448) );
  NAND2_X1 U5455 ( .A1(n5681), .A2(n5680), .ZN(n8458) );
  NAND2_X1 U5456 ( .A1(n5643), .A2(n5642), .ZN(n8457) );
  NAND2_X1 U5457 ( .A1(n5578), .A2(n5577), .ZN(n8515) );
  INV_X1 U5458 ( .A(P2_U3893), .ZN(n8402) );
  INV_X1 U5459 ( .A(n8261), .ZN(n8547) );
  AND3_X1 U5460 ( .A1(n5535), .A2(n5534), .A3(n5533), .ZN(n8557) );
  INV_X1 U5461 ( .A(n10444), .ZN(n8401) );
  NAND2_X1 U5462 ( .A1(n7634), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4712) );
  OAI21_X1 U5463 ( .B1(n4724), .B2(n6702), .A(n4720), .ZN(n4719) );
  NAND2_X1 U5464 ( .A1(n4724), .A2(n4721), .ZN(n4720) );
  NAND2_X1 U5465 ( .A1(n4728), .A2(n6705), .ZN(n4721) );
  AND2_X1 U5466 ( .A1(n4548), .A2(n4902), .ZN(n4562) );
  NAND2_X1 U5467 ( .A1(n4563), .A2(n4492), .ZN(n4548) );
  NOR2_X1 U5468 ( .A1(n8389), .A2(n4904), .ZN(n4903) );
  INV_X1 U5469 ( .A(n10464), .ZN(n10466) );
  NAND2_X1 U5470 ( .A1(n4916), .A2(n7415), .ZN(n7416) );
  OAI21_X1 U5471 ( .B1(n6737), .B2(n7878), .A(n6211), .ZN(n6739) );
  OAI21_X1 U5472 ( .B1(n8806), .B2(n4379), .A(n5730), .ZN(n5785) );
  AND2_X1 U5473 ( .A1(n6221), .A2(n6220), .ZN(n8796) );
  OR2_X1 U5474 ( .A1(n6219), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6221) );
  XNOR2_X1 U5475 ( .A(n6102), .B(n8934), .ZN(n9548) );
  NAND2_X1 U5476 ( .A1(n5045), .A2(n7029), .ZN(n5044) );
  OR2_X1 U5477 ( .A1(n7085), .A2(n9307), .ZN(n7084) );
  NAND2_X1 U5478 ( .A1(n7069), .A2(n5039), .ZN(n5038) );
  NAND2_X1 U5479 ( .A1(n4412), .A2(n5042), .ZN(n5039) );
  AND4_X1 U5480 ( .A1(n6340), .A2(n6339), .A3(n6338), .A4(n6337), .ZN(n9968)
         );
  INV_X1 U5481 ( .A(n9307), .ZN(n9287) );
  NAND2_X1 U5482 ( .A1(n6439), .A2(n6438), .ZN(n9762) );
  OR2_X1 U5483 ( .A1(n9751), .A2(n6433), .ZN(n6439) );
  AOI21_X1 U5484 ( .B1(n9724), .B2(n10372), .A(n9723), .ZN(n5030) );
  OR2_X1 U5485 ( .A1(n7088), .A2(n7190), .ZN(n10097) );
  NAND2_X1 U5486 ( .A1(n6727), .A2(n4574), .ZN(n6732) );
  INV_X1 U5487 ( .A(n4575), .ZN(n4574) );
  OAI21_X1 U5488 ( .B1(n8088), .B2(n10225), .A(n6726), .ZN(n4575) );
  NAND2_X1 U5489 ( .A1(n4612), .A2(n10424), .ZN(n4611) );
  INV_X1 U5490 ( .A(n9725), .ZN(n4612) );
  AND2_X1 U5491 ( .A1(n9710), .A2(n10142), .ZN(n6561) );
  AND2_X1 U5492 ( .A1(n4877), .A2(n4695), .ZN(n4694) );
  INV_X1 U5493 ( .A(n8025), .ZN(n4695) );
  NOR2_X1 U5494 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(n6085), .ZN(n4777) );
  OR2_X1 U5495 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6085) );
  CLKBUF_X1 U5496 ( .A(n5846), .Z(n5294) );
  OAI21_X1 U5497 ( .B1(n4916), .B2(n5820), .A(n5294), .ZN(n5289) );
  NAND2_X1 U5498 ( .A1(n5412), .A2(n6846), .ZN(n4510) );
  INV_X1 U5499 ( .A(n4509), .ZN(n4508) );
  AND3_X1 U5500 ( .A1(n4754), .A2(n4753), .A3(n9347), .ZN(n4752) );
  NAND2_X1 U5501 ( .A1(n4752), .A2(n4750), .ZN(n4749) );
  INV_X1 U5502 ( .A(n4416), .ZN(n4750) );
  NAND2_X1 U5503 ( .A1(n9342), .A2(n4416), .ZN(n4755) );
  OR2_X1 U5504 ( .A1(n4799), .A2(n8560), .ZN(n4798) );
  INV_X1 U5505 ( .A(n4771), .ZN(n4768) );
  AND2_X1 U5506 ( .A1(n5484), .A2(n4506), .ZN(n4505) );
  NAND2_X1 U5507 ( .A1(n4507), .A2(n6846), .ZN(n4506) );
  AND2_X1 U5508 ( .A1(n5511), .A2(n4475), .ZN(n4796) );
  NOR2_X1 U5509 ( .A1(n4794), .A2(n6182), .ZN(n4793) );
  NOR2_X1 U5510 ( .A1(n4797), .A2(n4795), .ZN(n4794) );
  INV_X1 U5511 ( .A(n5537), .ZN(n4795) );
  AND2_X1 U5512 ( .A1(n4798), .A2(n4480), .ZN(n4797) );
  NAND2_X1 U5513 ( .A1(n4540), .A2(n4539), .ZN(n9379) );
  INV_X1 U5514 ( .A(n4769), .ZN(n4539) );
  AOI21_X1 U5515 ( .B1(n4772), .B2(n4770), .A(n4461), .ZN(n4540) );
  AND2_X1 U5516 ( .A1(n4599), .A2(n4484), .ZN(n4786) );
  OR2_X1 U5517 ( .A1(n4788), .A2(n6846), .ZN(n4599) );
  AND2_X1 U5518 ( .A1(n5884), .A2(n5883), .ZN(n4787) );
  INV_X1 U5519 ( .A(n5664), .ZN(n4593) );
  INV_X1 U5520 ( .A(n8604), .ZN(n4564) );
  NOR2_X1 U5521 ( .A1(n10467), .A2(n4916), .ZN(n5822) );
  AND2_X1 U5522 ( .A1(n9407), .A2(n9315), .ZN(n4538) );
  NOR2_X1 U5523 ( .A1(n4566), .A2(n8575), .ZN(n4565) );
  NAND2_X1 U5524 ( .A1(n5830), .A2(n8545), .ZN(n4566) );
  INV_X1 U5525 ( .A(n5763), .ZN(n4811) );
  NAND2_X1 U5526 ( .A1(n4790), .A2(n5682), .ZN(n4698) );
  AOI21_X1 U5527 ( .B1(n8379), .B2(n8380), .A(n6697), .ZN(n6701) );
  INV_X1 U5528 ( .A(n5855), .ZN(n4922) );
  INV_X1 U5529 ( .A(n5854), .ZN(n4923) );
  INV_X1 U5530 ( .A(n7155), .ZN(n4665) );
  NAND2_X1 U5531 ( .A1(n4927), .A2(n5854), .ZN(n4926) );
  INV_X1 U5532 ( .A(n6978), .ZN(n5058) );
  OR2_X1 U5533 ( .A1(n4426), .A2(n5055), .ZN(n5054) );
  INV_X1 U5534 ( .A(n8826), .ZN(n5055) );
  NAND2_X1 U5535 ( .A1(n9418), .A2(n4380), .ZN(n9419) );
  INV_X1 U5536 ( .A(n6495), .ZN(n4619) );
  INV_X1 U5537 ( .A(n4618), .ZN(n4617) );
  OAI21_X1 U5538 ( .B1(n9924), .B2(n4619), .A(n6497), .ZN(n4618) );
  NAND2_X1 U5539 ( .A1(n10013), .A2(n9356), .ZN(n5003) );
  NAND2_X1 U5540 ( .A1(n4425), .A2(n4885), .ZN(n4884) );
  INV_X1 U5541 ( .A(n4886), .ZN(n4885) );
  XNOR2_X1 U5542 ( .A(n5766), .B(n5764), .ZN(n4820) );
  INV_X1 U5543 ( .A(n5691), .ZN(n4827) );
  AOI21_X1 U5544 ( .B1(n4843), .B2(n5543), .A(n4842), .ZN(n4841) );
  INV_X1 U5545 ( .A(n5564), .ZN(n4842) );
  INV_X1 U5546 ( .A(n5240), .ZN(n5488) );
  INV_X1 U5547 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4807) );
  INV_X1 U5548 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4806) );
  AOI21_X1 U5549 ( .B1(n4871), .B2(n4874), .A(n4870), .ZN(n4869) );
  INV_X1 U5550 ( .A(n7804), .ZN(n4870) );
  INV_X1 U5551 ( .A(n4871), .ZN(n4867) );
  OR2_X1 U5552 ( .A1(n5336), .A2(n5313), .ZN(n5319) );
  AOI21_X1 U5553 ( .B1(n6605), .B2(n7768), .A(n4714), .ZN(n4713) );
  INV_X1 U5554 ( .A(n7576), .ZN(n4714) );
  OAI21_X1 U5555 ( .B1(n8322), .B2(n8323), .A(n4716), .ZN(n6613) );
  OR2_X1 U5556 ( .A1(n6680), .A2(n8672), .ZN(n4716) );
  INV_X1 U5557 ( .A(n8391), .ZN(n4727) );
  INV_X1 U5558 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n4704) );
  NOR2_X1 U5559 ( .A1(n5572), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5589) );
  INV_X1 U5560 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8931) );
  INV_X1 U5561 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5199) );
  INV_X1 U5562 ( .A(n5408), .ZN(n5200) );
  INV_X1 U5563 ( .A(n7675), .ZN(n4675) );
  INV_X1 U5564 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4701) );
  OR2_X1 U5565 ( .A1(n8722), .A2(n8448), .ZN(n5000) );
  NAND2_X1 U5566 ( .A1(n4997), .A2(n4994), .ZN(n5001) );
  NOR2_X1 U5567 ( .A1(n6191), .A2(n8485), .ZN(n4976) );
  NOR2_X1 U5568 ( .A1(n8545), .A2(n4986), .ZN(n4985) );
  INV_X1 U5569 ( .A(n6181), .ZN(n4986) );
  INV_X1 U5570 ( .A(n4417), .ZN(n4983) );
  NAND2_X1 U5571 ( .A1(n4662), .A2(n5874), .ZN(n4661) );
  INV_X1 U5572 ( .A(n5873), .ZN(n4662) );
  INV_X1 U5573 ( .A(n5876), .ZN(n4659) );
  NOR2_X1 U5574 ( .A1(n6174), .A2(n4973), .ZN(n4971) );
  OR2_X1 U5575 ( .A1(n8677), .A2(n8246), .ZN(n5867) );
  OR2_X1 U5576 ( .A1(n6219), .A2(n6234), .ZN(n6745) );
  OAI21_X1 U5577 ( .B1(n5238), .B2(n4859), .A(n9055), .ZN(n4857) );
  OR2_X1 U5578 ( .A1(n5391), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5440) );
  OR2_X1 U5579 ( .A1(n5349), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5363) );
  NOR2_X1 U5580 ( .A1(n6421), .A2(n9204), .ZN(n4576) );
  NAND2_X1 U5581 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n4588) );
  AND2_X1 U5582 ( .A1(n6905), .A2(n10137), .ZN(n6902) );
  OR2_X1 U5583 ( .A1(n6556), .A2(n6539), .ZN(n9450) );
  NAND2_X1 U5584 ( .A1(n6556), .A2(n6539), .ZN(n9469) );
  NAND2_X1 U5585 ( .A1(n4958), .A2(n4959), .ZN(n4957) );
  OR2_X1 U5586 ( .A1(n10153), .A2(n6440), .ZN(n9457) );
  INV_X1 U5587 ( .A(n6511), .ZN(n4625) );
  NAND2_X1 U5588 ( .A1(n4617), .A2(n4619), .ZN(n4614) );
  NOR2_X1 U5589 ( .A1(n10039), .A2(n4881), .ZN(n9951) );
  NAND2_X1 U5590 ( .A1(n4883), .A2(n4882), .ZN(n4881) );
  INV_X1 U5591 ( .A(n4884), .ZN(n4883) );
  NOR2_X1 U5592 ( .A1(n6335), .A2(n7310), .ZN(n4577) );
  NAND2_X1 U5593 ( .A1(n10423), .A2(n10416), .ZN(n4886) );
  NAND2_X1 U5594 ( .A1(n10029), .A2(n6311), .ZN(n6321) );
  INV_X1 U5595 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7225) );
  OAI21_X1 U5596 ( .B1(n10336), .B2(n4422), .A(n10061), .ZN(n4606) );
  INV_X1 U5597 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6304) );
  INV_X1 U5598 ( .A(n9490), .ZN(n5020) );
  NAND2_X1 U5599 ( .A1(n10108), .A2(n4880), .ZN(n7754) );
  NAND2_X1 U5600 ( .A1(n4880), .A2(n9571), .ZN(n9482) );
  AND2_X1 U5601 ( .A1(n4880), .A2(n7277), .ZN(n4879) );
  NAND2_X1 U5602 ( .A1(n9832), .A2(n4402), .ZN(n9749) );
  NAND2_X1 U5603 ( .A1(n9832), .A2(n4892), .ZN(n9765) );
  NAND2_X1 U5604 ( .A1(n9832), .A2(n4894), .ZN(n9784) );
  INV_X1 U5605 ( .A(n4893), .ZN(n4894) );
  AND2_X1 U5606 ( .A1(n9832), .A2(n10253), .ZN(n9806) );
  AND2_X1 U5607 ( .A1(n9829), .A2(n9837), .ZN(n9832) );
  NOR2_X1 U5608 ( .A1(n9862), .A2(n10180), .ZN(n9829) );
  AND2_X1 U5609 ( .A1(n5724), .A2(n5696), .ZN(n5722) );
  AND2_X1 U5610 ( .A1(n5691), .A2(n5690), .ZN(n5714) );
  INV_X1 U5611 ( .A(n4829), .ZN(n4828) );
  OAI21_X1 U5612 ( .B1(n4838), .B2(n4830), .A(n4835), .ZN(n4829) );
  NOR2_X1 U5613 ( .A1(n5487), .A2(n5495), .ZN(n5081) );
  AND2_X1 U5614 ( .A1(n5491), .A2(n5148), .ZN(n5149) );
  NAND2_X1 U5615 ( .A1(n4815), .A2(n4813), .ZN(n5470) );
  NOR2_X1 U5616 ( .A1(n5488), .A2(n4814), .ZN(n4813) );
  INV_X1 U5617 ( .A(n5141), .ZN(n4814) );
  XNOR2_X1 U5618 ( .A(n5142), .B(SI_12_), .ZN(n5240) );
  NAND2_X1 U5619 ( .A1(n5118), .A2(n5117), .ZN(n5387) );
  NAND2_X1 U5620 ( .A1(n5121), .A2(n7130), .ZN(n4541) );
  OAI21_X1 U5621 ( .B1(n5121), .B2(n4531), .A(n4530), .ZN(n5107) );
  NAND2_X1 U5622 ( .A1(n5121), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4530) );
  NAND2_X1 U5623 ( .A1(n6773), .A2(n6772), .ZN(n7349) );
  NAND2_X1 U5624 ( .A1(n4876), .A2(n4875), .ZN(n7711) );
  XNOR2_X1 U5625 ( .A(n6810), .B(n8547), .ZN(n8187) );
  NAND2_X1 U5626 ( .A1(n4853), .A2(n6800), .ZN(n4852) );
  INV_X1 U5627 ( .A(n8297), .ZN(n8246) );
  INV_X1 U5628 ( .A(n8458), .ZN(n8275) );
  NAND2_X1 U5629 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n4859), .ZN(n4779) );
  AND2_X1 U5630 ( .A1(n5805), .A2(n5804), .ZN(n8413) );
  AND4_X1 U5631 ( .A1(n5262), .A2(n5261), .A3(n5260), .A4(n5259), .ZN(n8157)
         );
  OAI21_X1 U5632 ( .B1(n4383), .B2(n7473), .A(n4551), .ZN(n6625) );
  NAND2_X1 U5633 ( .A1(n4383), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4551) );
  OR2_X1 U5634 ( .A1(n7389), .A2(n7473), .ZN(n7387) );
  NAND2_X1 U5635 ( .A1(n7387), .A2(n6569), .ZN(n7562) );
  NAND2_X1 U5636 ( .A1(n6572), .A2(n7617), .ZN(n7549) );
  XNOR2_X1 U5637 ( .A(n4642), .B(n6595), .ZN(n7551) );
  NAND2_X1 U5638 ( .A1(n4913), .A2(n7616), .ZN(n7621) );
  NAND2_X1 U5639 ( .A1(n6572), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4641) );
  NAND2_X1 U5640 ( .A1(n4914), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7619) );
  INV_X1 U5641 ( .A(n7549), .ZN(n4914) );
  NAND2_X1 U5642 ( .A1(n4901), .A2(n7450), .ZN(n7402) );
  NAND3_X1 U5643 ( .A1(n4901), .A2(P2_REG2_REG_5__SCAN_IN), .A3(n7450), .ZN(
        n7452) );
  AOI21_X1 U5644 ( .B1(n7452), .B2(n7450), .A(n7451), .ZN(n7449) );
  NAND2_X1 U5645 ( .A1(n6647), .A2(n6646), .ZN(n7644) );
  OR2_X1 U5646 ( .A1(n4393), .A2(n7578), .ZN(n4629) );
  NAND2_X1 U5647 ( .A1(n7636), .A2(n4449), .ZN(n4630) );
  AND2_X1 U5648 ( .A1(n4631), .A2(n7146), .ZN(n6577) );
  XNOR2_X1 U5649 ( .A(n6578), .B(n4895), .ZN(n7909) );
  NAND2_X1 U5650 ( .A1(n6665), .A2(n6664), .ZN(n7912) );
  AOI21_X1 U5651 ( .B1(n7650), .B2(n4735), .A(n4732), .ZN(n6610) );
  AND2_X1 U5652 ( .A1(n7736), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4735) );
  OR2_X1 U5653 ( .A1(n4648), .A2(n4647), .ZN(n4911) );
  NAND2_X1 U5654 ( .A1(n4648), .A2(n4647), .ZN(n4912) );
  AND2_X1 U5655 ( .A1(n4646), .A2(n4645), .ZN(n4644) );
  NAND2_X1 U5656 ( .A1(n6677), .A2(n8310), .ZN(n8334) );
  NAND2_X1 U5657 ( .A1(n8351), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8369) );
  AND2_X1 U5658 ( .A1(n8356), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4897) );
  NAND2_X1 U5659 ( .A1(n8391), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4728) );
  NOR2_X1 U5660 ( .A1(n4905), .A2(n4907), .ZN(n4904) );
  INV_X1 U5661 ( .A(n4908), .ZN(n4905) );
  INV_X1 U5662 ( .A(n8392), .ZN(n4563) );
  NAND2_X1 U5663 ( .A1(n4908), .A2(n6704), .ZN(n4906) );
  INV_X1 U5664 ( .A(n4684), .ZN(n4683) );
  OAI21_X1 U5665 ( .B1(n8429), .B2(n4685), .A(n8420), .ZN(n4684) );
  NAND2_X1 U5666 ( .A1(n4686), .A2(n5896), .ZN(n4681) );
  NAND2_X1 U5667 ( .A1(n5655), .A2(n4496), .ZN(n5707) );
  NAND2_X1 U5668 ( .A1(n5655), .A2(n4699), .ZN(n5705) );
  NAND2_X1 U5669 ( .A1(n5589), .A2(n4409), .ZN(n5637) );
  NAND2_X1 U5670 ( .A1(n5589), .A2(n4702), .ZN(n5656) );
  AND2_X1 U5671 ( .A1(n4409), .A2(n4703), .ZN(n4702) );
  INV_X1 U5672 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n4703) );
  NAND2_X1 U5673 ( .A1(n5589), .A2(n8916), .ZN(n5614) );
  OR2_X1 U5674 ( .A1(n5554), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5572) );
  INV_X1 U5675 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U5676 ( .A1(n5204), .A2(n4706), .ZN(n5532) );
  NAND2_X1 U5677 ( .A1(n5204), .A2(n5203), .ZN(n5530) );
  OR2_X1 U5678 ( .A1(n5501), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U5679 ( .A1(n5200), .A2(n4708), .ZN(n5478) );
  AND2_X1 U5680 ( .A1(n4428), .A2(n5201), .ZN(n4708) );
  INV_X1 U5681 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U5682 ( .A1(n5202), .A2(n8931), .ZN(n5501) );
  INV_X1 U5683 ( .A(n5478), .ZN(n5202) );
  OR2_X1 U5684 ( .A1(n7869), .A2(n7873), .ZN(n8598) );
  NAND2_X1 U5685 ( .A1(n6168), .A2(n6167), .ZN(n8605) );
  NAND2_X1 U5686 ( .A1(n5198), .A2(n5197), .ZN(n5425) );
  INV_X1 U5687 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5197) );
  INV_X1 U5688 ( .A(n5423), .ZN(n5198) );
  NAND2_X1 U5689 ( .A1(n4969), .A2(n6161), .ZN(n7697) );
  OAI21_X1 U5690 ( .B1(n7505), .B2(n4927), .A(n5854), .ZN(n7693) );
  OR2_X1 U5691 ( .A1(n5368), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U5692 ( .A1(n7355), .A2(n4701), .ZN(n5354) );
  NAND2_X1 U5693 ( .A1(n5850), .A2(n5849), .ZN(n7537) );
  NAND2_X1 U5694 ( .A1(n8688), .A2(n8687), .ZN(n4656) );
  NAND2_X1 U5695 ( .A1(n5849), .A2(n5819), .ZN(n7429) );
  INV_X1 U5696 ( .A(n8687), .ZN(n8691) );
  NAND2_X1 U5697 ( .A1(n5264), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5268) );
  OR2_X1 U5698 ( .A1(n5300), .A2(n7468), .ZN(n5269) );
  OR2_X1 U5699 ( .A1(n6846), .A2(n6755), .ZN(n7462) );
  OR2_X1 U5700 ( .A1(n10488), .A2(n6236), .ZN(n7118) );
  NOR2_X1 U5701 ( .A1(n8413), .A2(n8412), .ZN(n8704) );
  AOI21_X1 U5702 ( .B1(n4998), .B2(n4445), .A(n4989), .ZN(n6198) );
  NAND2_X1 U5703 ( .A1(n4404), .A2(n4990), .ZN(n4989) );
  NAND2_X1 U5704 ( .A1(n4400), .A2(n4995), .ZN(n4990) );
  AND2_X1 U5705 ( .A1(n5757), .A2(n5756), .ZN(n8090) );
  AND2_X1 U5706 ( .A1(n5761), .A2(n5760), .ZN(n8092) );
  NAND2_X1 U5707 ( .A1(n5001), .A2(n4420), .ZN(n4991) );
  NAND2_X1 U5708 ( .A1(n8429), .A2(n4399), .ZN(n4999) );
  NAND2_X1 U5709 ( .A1(n5001), .A2(n5000), .ZN(n8431) );
  NAND2_X1 U5710 ( .A1(n8432), .A2(n8692), .ZN(n4557) );
  OAI21_X1 U5711 ( .B1(n6188), .B2(n8481), .A(n6190), .ZN(n4981) );
  NAND2_X1 U5712 ( .A1(n4943), .A2(n5881), .ZN(n8501) );
  NAND2_X1 U5713 ( .A1(n4944), .A2(n5880), .ZN(n4943) );
  INV_X1 U5714 ( .A(n7503), .ZN(n6587) );
  OR2_X1 U5715 ( .A1(n8767), .A2(n8261), .ZN(n8522) );
  AND2_X1 U5716 ( .A1(n6162), .A2(n6161), .ZN(n4968) );
  NAND2_X1 U5717 ( .A1(n4920), .A2(n4924), .ZN(n7695) );
  NAND2_X1 U5718 ( .A1(n7505), .A2(n5854), .ZN(n4920) );
  OR2_X1 U5719 ( .A1(n7462), .A2(n8795), .ZN(n6872) );
  INV_X1 U5720 ( .A(n10488), .ZN(n10473) );
  CLKBUF_X1 U5721 ( .A(n5919), .Z(n5920) );
  AND2_X1 U5722 ( .A1(n5382), .A2(n5419), .ZN(n7455) );
  INV_X1 U5723 ( .A(n4421), .ZN(n5051) );
  OAI21_X1 U5724 ( .B1(n4421), .B2(n5050), .A(n8872), .ZN(n5049) );
  INV_X1 U5725 ( .A(n7012), .ZN(n5050) );
  NAND2_X1 U5726 ( .A1(n4467), .A2(n4512), .ZN(n4511) );
  INV_X1 U5727 ( .A(n6965), .ZN(n4512) );
  INV_X1 U5728 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7310) );
  NAND2_X1 U5729 ( .A1(n4576), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6441) );
  OR2_X1 U5730 ( .A1(n8889), .A2(n6984), .ZN(n5076) );
  AND2_X1 U5731 ( .A1(n7040), .A2(n7038), .ZN(n9198) );
  AND2_X1 U5732 ( .A1(n6378), .A2(n4585), .ZN(n6411) );
  NOR2_X1 U5733 ( .A1(n4589), .A2(n4586), .ZN(n4585) );
  OR2_X1 U5734 ( .A1(n4588), .A2(n4587), .ZN(n4586) );
  INV_X1 U5735 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n4587) );
  NOR2_X1 U5736 ( .A1(n6394), .A2(n4588), .ZN(n6401) );
  INV_X1 U5737 ( .A(n5063), .ZN(n9260) );
  AOI21_X1 U5738 ( .B1(n5062), .B2(n4419), .A(n4398), .ZN(n5063) );
  NAND2_X1 U5739 ( .A1(n8882), .A2(n8883), .ZN(n8881) );
  INV_X1 U5740 ( .A(n8883), .ZN(n5042) );
  NAND2_X1 U5741 ( .A1(n8825), .A2(n8826), .ZN(n5060) );
  INV_X1 U5742 ( .A(n9947), .ZN(n4518) );
  NAND2_X1 U5743 ( .A1(n9444), .A2(n4515), .ZN(n4514) );
  AND2_X1 U5744 ( .A1(n9744), .A2(n4516), .ZN(n4515) );
  AND2_X1 U5745 ( .A1(n9823), .A2(n4517), .ZN(n4516) );
  NOR2_X1 U5746 ( .A1(n9757), .A2(n9776), .ZN(n4517) );
  NOR2_X1 U5747 ( .A1(n9424), .A2(n4761), .ZN(n9544) );
  OR2_X1 U5748 ( .A1(n7244), .A2(n7243), .ZN(n7255) );
  OR2_X1 U5749 ( .A1(n7263), .A2(n7264), .ZN(n7304) );
  OR2_X1 U5750 ( .A1(n7257), .A2(n7258), .ZN(n7315) );
  OR2_X1 U5751 ( .A1(n7601), .A2(n7602), .ZN(n8047) );
  OR2_X1 U5752 ( .A1(n7319), .A2(n7318), .ZN(n7592) );
  OR2_X1 U5753 ( .A1(n7594), .A2(n7595), .ZN(n8059) );
  NOR2_X1 U5754 ( .A1(n8049), .A2(n10306), .ZN(n9690) );
  INV_X1 U5755 ( .A(n8016), .ZN(n9446) );
  AND2_X1 U5756 ( .A1(n9450), .A2(n9469), .ZN(n8016) );
  NOR2_X1 U5757 ( .A1(n6517), .A2(n4963), .ZN(n4962) );
  INV_X1 U5758 ( .A(n4964), .ZN(n4963) );
  AND4_X1 U5759 ( .A1(n6459), .A2(n6458), .A3(n6457), .A4(n6456), .ZN(n8818)
         );
  AOI21_X1 U5760 ( .B1(n5009), .B2(n5011), .A(n5007), .ZN(n5006) );
  NOR2_X1 U5761 ( .A1(n5008), .A2(n6449), .ZN(n5007) );
  AOI21_X1 U5762 ( .B1(n5015), .B2(n9776), .A(n5014), .ZN(n5013) );
  INV_X1 U5763 ( .A(n9454), .ZN(n5014) );
  NAND2_X1 U5764 ( .A1(n9745), .A2(n9744), .ZN(n9743) );
  AND2_X1 U5765 ( .A1(n9457), .A2(n9460), .ZN(n9744) );
  NAND2_X1 U5766 ( .A1(n6420), .A2(n6419), .ZN(n9779) );
  INV_X1 U5767 ( .A(n9777), .ZN(n6420) );
  AND2_X1 U5768 ( .A1(n9310), .A2(n9377), .ZN(n9801) );
  NAND2_X1 U5769 ( .A1(n6386), .A2(n9520), .ZN(n9819) );
  NOR2_X1 U5770 ( .A1(n4934), .A2(n4460), .ZN(n4933) );
  INV_X1 U5771 ( .A(n6502), .ZN(n4934) );
  AND2_X1 U5772 ( .A1(n9878), .A2(n10267), .ZN(n9879) );
  NAND2_X1 U5773 ( .A1(n9879), .A2(n10262), .ZN(n9862) );
  AND2_X1 U5774 ( .A1(n6366), .A2(n6365), .ZN(n9894) );
  AOI21_X1 U5775 ( .B1(n4930), .B2(n4932), .A(n4451), .ZN(n4928) );
  INV_X1 U5776 ( .A(n4577), .ZN(n6341) );
  NAND2_X1 U5777 ( .A1(n9961), .A2(n9965), .ZN(n9960) );
  AND4_X1 U5778 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .ZN(n9941)
         );
  NAND2_X1 U5779 ( .A1(n6328), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6335) );
  NOR2_X1 U5780 ( .A1(n10039), .A2(n4886), .ZN(n10021) );
  NAND2_X1 U5781 ( .A1(n5004), .A2(n9496), .ZN(n10012) );
  NAND2_X1 U5782 ( .A1(n6321), .A2(n6320), .ZN(n5004) );
  NAND2_X1 U5783 ( .A1(n10012), .A2(n10013), .ZN(n10011) );
  NOR2_X1 U5784 ( .A1(n10039), .A2(n10050), .ZN(n10041) );
  INV_X1 U5785 ( .A(n6479), .ZN(n4610) );
  AND3_X1 U5786 ( .A1(n5958), .A2(n4395), .A3(n10397), .ZN(n10345) );
  AND4_X1 U5787 ( .A1(n6295), .A2(n6294), .A3(n6293), .A4(n6292), .ZN(n10072)
         );
  NAND2_X1 U5788 ( .A1(n5958), .A2(n4395), .ZN(n10368) );
  NAND2_X1 U5789 ( .A1(n6884), .A2(n5033), .ZN(n6519) );
  XNOR2_X1 U5790 ( .A(n10108), .B(n7518), .ZN(n7520) );
  AND2_X1 U5791 ( .A1(n10122), .A2(n4879), .ZN(n10100) );
  NAND2_X1 U5792 ( .A1(n10122), .A2(n7277), .ZN(n7517) );
  INV_X1 U5793 ( .A(n8080), .ZN(n6726) );
  NAND2_X1 U5794 ( .A1(n6025), .A2(n6024), .ZN(n10197) );
  INV_X1 U5795 ( .A(n7173), .ZN(n6046) );
  INV_X1 U5796 ( .A(n10369), .ZN(n10214) );
  AND2_X1 U5797 ( .A1(n10133), .A2(n9539), .ZN(n10369) );
  OR2_X1 U5798 ( .A1(n9315), .A2(n7087), .ZN(n10401) );
  AND2_X1 U5799 ( .A1(n6128), .A2(n7082), .ZN(n8012) );
  AND3_X1 U5800 ( .A1(n7080), .A2(n7088), .A3(n7079), .ZN(n6525) );
  OAI21_X1 U5801 ( .B1(n5793), .B2(n5792), .A(n5791), .ZN(n5796) );
  XNOR2_X1 U5802 ( .A(n5793), .B(n5792), .ZN(n8006) );
  INV_X1 U5803 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4696) );
  XNOR2_X1 U5804 ( .A(n5758), .B(n5759), .ZN(n8103) );
  NAND2_X1 U5805 ( .A1(n6108), .A2(n6107), .ZN(n6113) );
  INV_X1 U5806 ( .A(n6111), .ZN(n6108) );
  NAND2_X1 U5807 ( .A1(n6081), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6100) );
  INV_X1 U5808 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6104) );
  INV_X1 U5809 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9087) );
  XNOR2_X1 U5810 ( .A(n5582), .B(n5567), .ZN(n7689) );
  NOR2_X1 U5811 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6078) );
  NAND2_X1 U5812 ( .A1(n4600), .A2(n4601), .ZN(n5566) );
  AOI21_X1 U5813 ( .B1(n5210), .B2(n4602), .A(n4405), .ZN(n4601) );
  AND2_X1 U5814 ( .A1(n6034), .A2(n6033), .ZN(n8068) );
  XNOR2_X1 U5815 ( .A(n5211), .B(n5210), .ZN(n7299) );
  OR2_X1 U5816 ( .A1(n6080), .A2(n10278), .ZN(n6026) );
  XNOR2_X1 U5817 ( .A(n5490), .B(n5240), .ZN(n7185) );
  INV_X1 U5818 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U5819 ( .A1(n5414), .A2(n4802), .ZN(n5416) );
  XNOR2_X1 U5820 ( .A(n5107), .B(SI_4_), .ZN(n5346) );
  INV_X1 U5821 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5960) );
  INV_X1 U5822 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4745) );
  INV_X1 U5823 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9088) );
  NOR2_X1 U5824 ( .A1(n6671), .A2(n8585), .ZN(n4649) );
  AND4_X1 U5825 ( .A1(n5409), .A2(n5410), .A3(n5411), .A4(n4801), .ZN(n7770)
         );
  NAND2_X1 U5826 ( .A1(n5265), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n4801) );
  OAI21_X1 U5827 ( .B1(n6814), .B2(n8254), .A(n4457), .ZN(n4503) );
  AND4_X1 U5828 ( .A1(n5399), .A2(n5398), .A3(n5397), .A4(n5396), .ZN(n7776)
         );
  NAND2_X1 U5829 ( .A1(n7711), .A2(n6788), .ZN(n7773) );
  NAND2_X1 U5830 ( .A1(n8284), .A2(n6808), .ZN(n8189) );
  OR2_X1 U5831 ( .A1(n6777), .A2(n4493), .ZN(n7371) );
  INV_X1 U5832 ( .A(n8298), .ZN(n8156) );
  NAND2_X1 U5833 ( .A1(n4868), .A2(n4871), .ZN(n7805) );
  OR2_X1 U5834 ( .A1(n4876), .A2(n4874), .ZN(n4868) );
  INV_X1 U5835 ( .A(n4849), .ZN(n8221) );
  AOI21_X1 U5836 ( .B1(n8125), .B2(n6796), .A(n4852), .ZN(n4849) );
  INV_X1 U5837 ( .A(n8286), .ZN(n8274) );
  INV_X1 U5838 ( .A(n6783), .ZN(n4861) );
  NAND2_X1 U5839 ( .A1(n4862), .A2(n6783), .ZN(n7491) );
  AND2_X1 U5840 ( .A1(n6855), .A2(n7160), .ZN(n7489) );
  AND2_X1 U5841 ( .A1(n6851), .A2(n6850), .ZN(n8271) );
  OR2_X1 U5842 ( .A1(n8283), .A2(n8282), .ZN(n8284) );
  AND2_X1 U5843 ( .A1(n5805), .A2(n5737), .ZN(n8422) );
  NAND2_X1 U5844 ( .A1(n5662), .A2(n5661), .ZN(n8474) );
  INV_X1 U5845 ( .A(n8214), .ZN(n8527) );
  INV_X1 U5846 ( .A(n8157), .ZN(n8607) );
  INV_X1 U5847 ( .A(n7776), .ZN(n8608) );
  INV_X1 U5848 ( .A(n7770), .ZN(n8299) );
  CLKBUF_X1 U5849 ( .A(n6762), .Z(n8304) );
  NAND2_X1 U5850 ( .A1(n4383), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4542) );
  XNOR2_X1 U5851 ( .A(n6575), .B(n7136), .ZN(n7636) );
  NAND2_X1 U5852 ( .A1(n7636), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7635) );
  XNOR2_X1 U5853 ( .A(n6608), .B(n7656), .ZN(n7650) );
  NAND2_X1 U5854 ( .A1(n4733), .A2(n6609), .ZN(n7735) );
  NAND2_X1 U5855 ( .A1(n7650), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4733) );
  AOI21_X1 U5856 ( .B1(n7925), .B2(n4411), .A(n7924), .ZN(n7927) );
  NAND2_X1 U5857 ( .A1(n4912), .A2(n4911), .ZN(n8307) );
  NAND2_X1 U5858 ( .A1(n4502), .A2(n4501), .ZN(n8408) );
  OR2_X1 U5859 ( .A1(n8405), .A2(n4408), .ZN(n4501) );
  NAND2_X1 U5860 ( .A1(n8407), .A2(n6615), .ZN(n4502) );
  NAND2_X1 U5861 ( .A1(n4635), .A2(n6584), .ZN(n4634) );
  NOR2_X1 U5862 ( .A1(n8389), .A2(n6585), .ZN(n4633) );
  NAND2_X1 U5863 ( .A1(n4639), .A2(n8385), .ZN(n4638) );
  NAND2_X1 U5864 ( .A1(n4723), .A2(n8378), .ZN(n4722) );
  NAND2_X1 U5865 ( .A1(n6189), .A2(n6188), .ZN(n8480) );
  NAND2_X1 U5866 ( .A1(n4424), .A2(n5886), .ZN(n4941) );
  NAND2_X1 U5867 ( .A1(n4942), .A2(n4944), .ZN(n4940) );
  NAND2_X1 U5868 ( .A1(n6179), .A2(n6178), .ZN(n8554) );
  NAND2_X1 U5869 ( .A1(n6239), .A2(n8461), .ZN(n8618) );
  OR2_X1 U5870 ( .A1(n7118), .A2(n8795), .ZN(n10458) );
  XNOR2_X1 U5871 ( .A(n7413), .B(n4916), .ZN(n7419) );
  INV_X1 U5872 ( .A(n8618), .ZN(n8589) );
  INV_X1 U5873 ( .A(n10458), .ZN(n8588) );
  NAND2_X2 U5874 ( .A1(n6238), .A2(n10458), .ZN(n10464) );
  NAND2_X1 U5875 ( .A1(n8428), .A2(n8429), .ZN(n4682) );
  AOI21_X1 U5876 ( .B1(n4558), .B2(n8696), .A(n4555), .ZN(n8715) );
  NAND2_X1 U5877 ( .A1(n4557), .A2(n4556), .ZN(n4555) );
  XNOR2_X1 U5878 ( .A(n8431), .B(n8430), .ZN(n4558) );
  NAND2_X1 U5879 ( .A1(n8448), .A2(n8609), .ZN(n4556) );
  NAND2_X1 U5880 ( .A1(n4546), .A2(n4545), .ZN(n4544) );
  NAND2_X1 U5881 ( .A1(n8458), .A2(n8609), .ZN(n4545) );
  NAND2_X1 U5882 ( .A1(n5674), .A2(n5673), .ZN(n8728) );
  NAND2_X1 U5883 ( .A1(n5653), .A2(n5652), .ZN(n8734) );
  NAND2_X1 U5884 ( .A1(n4740), .A2(n4736), .ZN(n8464) );
  NAND2_X1 U5885 ( .A1(n5636), .A2(n5635), .ZN(n8740) );
  AND2_X1 U5886 ( .A1(n4741), .A2(n4427), .ZN(n4739) );
  NAND2_X1 U5887 ( .A1(n4967), .A2(n6186), .ZN(n8511) );
  NAND2_X1 U5888 ( .A1(n5529), .A2(n5528), .ZN(n8772) );
  NAND2_X1 U5889 ( .A1(n4987), .A2(n6181), .ZN(n8546) );
  NAND2_X1 U5890 ( .A1(n6179), .A2(n4417), .ZN(n4987) );
  NAND2_X1 U5891 ( .A1(n8561), .A2(n5873), .ZN(n4660) );
  NAND2_X1 U5892 ( .A1(n5517), .A2(n5516), .ZN(n8779) );
  NAND2_X1 U5893 ( .A1(n4946), .A2(n5869), .ZN(n8576) );
  NAND2_X1 U5894 ( .A1(n5477), .A2(n5476), .ZN(n8227) );
  NAND2_X1 U5895 ( .A1(n5568), .A2(n7139), .ZN(n5406) );
  AND2_X1 U5896 ( .A1(n6860), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7195) );
  INV_X1 U5897 ( .A(n7193), .ZN(n7198) );
  NOR2_X1 U5898 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4800) );
  INV_X1 U5899 ( .A(n6217), .ZN(n7971) );
  NAND2_X1 U5900 ( .A1(n5918), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5916) );
  OR2_X1 U5901 ( .A1(n5917), .A2(n5914), .ZN(n4845) );
  NAND2_X1 U5902 ( .A1(n5239), .A2(n5840), .ZN(n7730) );
  INV_X1 U5903 ( .A(n6200), .ZN(n7787) );
  INV_X1 U5904 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9061) );
  INV_X1 U5905 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9074) );
  INV_X1 U5906 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9107) );
  INV_X1 U5907 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U5908 ( .A1(n4525), .A2(n4524), .ZN(n5310) );
  NAND2_X1 U5909 ( .A1(n5309), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U5910 ( .A1(n4526), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n4525) );
  AND2_X1 U5911 ( .A1(n6454), .A2(n6248), .ZN(n9719) );
  NOR3_X1 U5912 ( .A1(n9250), .A2(n8839), .A3(n8838), .ZN(n8841) );
  AND4_X1 U5913 ( .A1(n6361), .A2(n6360), .A3(n6359), .A4(n6358), .ZN(n9942)
         );
  OR2_X1 U5914 ( .A1(n7091), .A2(n7280), .ZN(n9301) );
  NAND2_X1 U5915 ( .A1(n7089), .A2(n10097), .ZN(n9256) );
  OR2_X1 U5916 ( .A1(n7091), .A2(n6095), .ZN(n9277) );
  NOR2_X1 U5917 ( .A1(n9273), .A2(n5037), .ZN(n5036) );
  INV_X1 U5918 ( .A(n6994), .ZN(n5037) );
  NAND2_X1 U5919 ( .A1(n9187), .A2(n6994), .ZN(n9272) );
  INV_X1 U5920 ( .A(n9301), .ZN(n9289) );
  OR3_X1 U5921 ( .A1(n7099), .A2(n7190), .A3(n7092), .ZN(n9307) );
  OR2_X1 U5922 ( .A1(n7101), .A2(n7100), .ZN(n9305) );
  AOI21_X1 U5923 ( .B1(n9477), .B2(n9475), .A(n9540), .ZN(n9476) );
  NOR2_X1 U5924 ( .A1(n9715), .A2(n4579), .ZN(n4578) );
  OR2_X1 U5925 ( .A1(n9543), .A2(n5033), .ZN(n5032) );
  NAND4_X1 U5926 ( .A1(n6448), .A2(n6447), .A3(n6446), .A4(n6445), .ZN(n9746)
         );
  NAND2_X1 U5927 ( .A1(n6428), .A2(n6427), .ZN(n9781) );
  OR2_X1 U5928 ( .A1(n9768), .A2(n6433), .ZN(n6428) );
  NAND2_X1 U5929 ( .A1(n6418), .A2(n6417), .ZN(n9803) );
  INV_X1 U5930 ( .A(n10334), .ZN(n9566) );
  NAND2_X1 U5931 ( .A1(n6274), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6284) );
  AND2_X1 U5932 ( .A1(n7181), .A2(n7180), .ZN(n7245) );
  OR2_X1 U5933 ( .A1(n7223), .A2(n7224), .ZN(n7261) );
  OR2_X1 U5934 ( .A1(n7308), .A2(n7309), .ZN(n7599) );
  AND2_X1 U5935 ( .A1(n10288), .A2(n10287), .ZN(n10296) );
  INV_X1 U5936 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6017) );
  AOI21_X1 U5937 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n8064), .A(n9688), .ZN(
        n9695) );
  OR2_X1 U5938 ( .A1(n10318), .A2(n10317), .ZN(n10327) );
  NAND2_X1 U5939 ( .A1(n8015), .A2(n6724), .ZN(n8088) );
  AND2_X1 U5940 ( .A1(n6534), .A2(n6455), .ZN(n8081) );
  OAI21_X1 U5941 ( .B1(n9742), .B2(n6515), .A(n4964), .ZN(n9726) );
  NAND2_X1 U5942 ( .A1(n9734), .A2(n9733), .ZN(n10146) );
  NAND2_X1 U5943 ( .A1(n6510), .A2(n6509), .ZN(n9775) );
  NAND2_X1 U5944 ( .A1(n4935), .A2(n6502), .ZN(n9856) );
  NAND2_X1 U5945 ( .A1(n9905), .A2(n6497), .ZN(n9889) );
  NAND2_X1 U5946 ( .A1(n5025), .A2(n9360), .ZN(n9964) );
  OAI21_X1 U5947 ( .B1(n10123), .B2(n4880), .A(n10114), .ZN(n10115) );
  INV_X1 U5948 ( .A(n10123), .ZN(n10359) );
  NOR2_X1 U5949 ( .A1(n10146), .A2(n4570), .ZN(n10237) );
  NAND2_X1 U5950 ( .A1(n4572), .A2(n4571), .ZN(n4570) );
  INV_X1 U5951 ( .A(n10147), .ZN(n4571) );
  NAND2_X1 U5952 ( .A1(n10148), .A2(n10424), .ZN(n4572) );
  INV_X1 U5953 ( .A(n9735), .ZN(n10240) );
  INV_X1 U5954 ( .A(n9787), .ZN(n10249) );
  INV_X1 U5955 ( .A(n9808), .ZN(n10253) );
  NAND2_X1 U5956 ( .A1(n7786), .A2(n5983), .ZN(n4527) );
  INV_X1 U5957 ( .A(n9881), .ZN(n10267) );
  INV_X1 U5958 ( .A(n7994), .ZN(n9981) );
  CLKBUF_X1 U5959 ( .A(n6096), .Z(n7989) );
  INV_X1 U5960 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9063) );
  INV_X1 U5961 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9037) );
  INV_X1 U5962 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9062) );
  INV_X1 U5963 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7734) );
  INV_X1 U5964 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7707) );
  INV_X1 U5965 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7502) );
  INV_X1 U5966 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8948) );
  INV_X1 U5967 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n8944) );
  INV_X1 U5968 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9171) );
  INV_X1 U5969 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6001) );
  INV_X1 U5970 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5969) );
  OAI21_X1 U5971 ( .B1(n5936), .B2(n7133), .A(n4513), .ZN(n5277) );
  NAND2_X1 U5972 ( .A1(n5936), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U5973 ( .A1(n5935), .A2(n5934), .ZN(n7228) );
  OR2_X1 U5974 ( .A1(n7927), .A2(n4649), .ZN(n4648) );
  NAND2_X1 U5975 ( .A1(n4712), .A2(n6605), .ZN(n7577) );
  NAND2_X1 U5976 ( .A1(n4730), .A2(n8385), .ZN(n4729) );
  NAND2_X1 U5977 ( .A1(n6739), .A2(n10464), .ZN(n6244) );
  OAI21_X1 U5978 ( .B1(n6738), .B2(n7125), .A(n7126), .ZN(n4966) );
  AND2_X1 U5979 ( .A1(n7086), .A2(n9287), .ZN(n7110) );
  AOI21_X1 U5980 ( .B1(n8076), .B2(n9551), .A(n4553), .ZN(n4552) );
  INV_X1 U5981 ( .A(n5029), .ZN(n5028) );
  OAI21_X1 U5982 ( .B1(n9725), .B2(n10124), .A(n5030), .ZN(n5029) );
  OAI21_X1 U5983 ( .B1(n6732), .B2(n10440), .A(n6733), .ZN(n6735) );
  NAND2_X1 U5984 ( .A1(n6530), .A2(n6529), .ZN(P1_U3549) );
  NOR2_X1 U5985 ( .A1(n5075), .A2(n6528), .ZN(n6529) );
  OAI22_X1 U5986 ( .A1(n10194), .A2(n4880), .B1(n10442), .B2(n6253), .ZN(n7526) );
  AND2_X1 U5987 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  INV_X1 U5988 ( .A(n6714), .ZN(n6715) );
  OAI21_X1 U5989 ( .B1(n8023), .B2(n10266), .A(n6713), .ZN(n6714) );
  OAI21_X1 U5990 ( .B1(n10266), .B2(n4880), .A(n4605), .ZN(n7524) );
  OR2_X1 U5991 ( .A1(n10430), .A2(n7523), .ZN(n4605) );
  OAI21_X1 U5992 ( .B1(n8806), .B2(n8004), .A(n4692), .ZN(P1_U3326) );
  INV_X1 U5993 ( .A(n4693), .ZN(n4692) );
  NAND2_X1 U5994 ( .A1(n5167), .A2(n5166), .ZN(n5210) );
  INV_X1 U5995 ( .A(n8485), .ZN(n8481) );
  INV_X1 U5996 ( .A(n4378), .ZN(n6390) );
  NOR2_X1 U5997 ( .A1(n6328), .A2(n6323), .ZN(n4392) );
  OR2_X1 U5998 ( .A1(n6575), .A2(n7637), .ZN(n4393) );
  AND3_X1 U5999 ( .A1(n4899), .A2(n6581), .A3(P2_REG2_REG_15__SCAN_IN), .ZN(
        n4394) );
  NAND2_X1 U6000 ( .A1(n6168), .A2(n4972), .ZN(n7886) );
  AND2_X1 U6001 ( .A1(n5957), .A2(n10392), .ZN(n4395) );
  NAND2_X1 U6002 ( .A1(n8761), .A2(n8536), .ZN(n4396) );
  AND2_X1 U6003 ( .A1(n4841), .A2(n4834), .ZN(n4397) );
  INV_X1 U6004 ( .A(n7337), .ZN(n8306) );
  OR2_X1 U6005 ( .A1(n5066), .A2(n4431), .ZN(n4398) );
  OR2_X1 U6006 ( .A1(n8717), .A2(n8440), .ZN(n4399) );
  AND2_X1 U6007 ( .A1(n4420), .A2(n6196), .ZN(n4400) );
  AOI21_X1 U6008 ( .B1(n9241), .B2(n6978), .A(n4410), .ZN(n5061) );
  AND2_X1 U6009 ( .A1(n10031), .A2(n9343), .ZN(n4401) );
  AND2_X1 U6010 ( .A1(n4892), .A2(n4891), .ZN(n4402) );
  NAND2_X1 U6011 ( .A1(n4521), .A2(n5884), .ZN(n5886) );
  INV_X1 U6012 ( .A(n5325), .ZN(n4529) );
  AND2_X1 U6013 ( .A1(n4465), .A2(n4779), .ZN(n4403) );
  AND2_X1 U6014 ( .A1(n4468), .A2(n4992), .ZN(n4404) );
  AND2_X1 U6015 ( .A1(n5542), .A2(SI_18_), .ZN(n4405) );
  INV_X1 U6016 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10278) );
  AND2_X1 U6017 ( .A1(n4911), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4406) );
  AOI21_X1 U6018 ( .B1(n10336), .B2(n4610), .A(n4422), .ZN(n4609) );
  OAI21_X1 U6019 ( .B1(n6480), .B2(n9341), .A(n4609), .ZN(n10060) );
  INV_X1 U6020 ( .A(n6674), .ZN(n4647) );
  OR2_X1 U6021 ( .A1(n4647), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4407) );
  OR2_X1 U6022 ( .A1(n8404), .A2(n6615), .ZN(n4408) );
  NOR2_X1 U6023 ( .A1(n6616), .A2(n4383), .ZN(n8396) );
  AND2_X1 U6024 ( .A1(n8916), .A2(n4704), .ZN(n4409) );
  XOR2_X1 U6025 ( .A(n6979), .B(n7043), .Z(n4410) );
  OR2_X1 U6026 ( .A1(n6578), .A2(n7914), .ZN(n4411) );
  AND2_X1 U6027 ( .A1(n7054), .A2(n5040), .ZN(n4412) );
  NAND2_X1 U6028 ( .A1(n5978), .A2(n5979), .ZN(n5981) );
  NAND2_X1 U6029 ( .A1(n5062), .A2(n5067), .ZN(n7962) );
  NAND2_X1 U6030 ( .A1(n5025), .A2(n5024), .ZN(n9943) );
  NOR2_X1 U6031 ( .A1(n8189), .A2(n8180), .ZN(n4413) );
  AND2_X1 U6032 ( .A1(n4406), .A2(n4912), .ZN(n4414) );
  OR2_X1 U6033 ( .A1(n8834), .A2(n9252), .ZN(n4415) );
  AND3_X1 U6034 ( .A1(n4758), .A2(n9341), .A3(n4757), .ZN(n4416) );
  NOR2_X1 U6035 ( .A1(n6180), .A2(n4988), .ZN(n4417) );
  NOR2_X1 U6036 ( .A1(n6983), .A2(n9298), .ZN(n4418) );
  AND2_X1 U6037 ( .A1(n5067), .A2(n5064), .ZN(n4419) );
  AND2_X1 U6038 ( .A1(n4399), .A2(n5000), .ZN(n4420) );
  NAND2_X1 U6039 ( .A1(n7011), .A2(n8871), .ZN(n4421) );
  AND2_X1 U6040 ( .A1(n10072), .A2(n10403), .ZN(n4422) );
  NOR2_X1 U6041 ( .A1(n6826), .A2(n8231), .ZN(n4423) );
  NAND2_X1 U6042 ( .A1(n5884), .A2(n4742), .ZN(n4424) );
  NOR2_X1 U6043 ( .A1(n10227), .A2(n7994), .ZN(n4425) );
  NOR2_X1 U6044 ( .A1(n5565), .A2(n4405), .ZN(n4843) );
  INV_X1 U6045 ( .A(n4843), .ZN(n4837) );
  AND2_X1 U6046 ( .A1(n6978), .A2(n4410), .ZN(n4426) );
  INV_X1 U6047 ( .A(n7400), .ZN(n7152) );
  OR2_X1 U6048 ( .A1(n8230), .A2(n8496), .ZN(n4427) );
  BUF_X1 U6049 ( .A(n6319), .Z(n10079) );
  AND3_X1 U6050 ( .A1(n5199), .A2(n4710), .A3(n4709), .ZN(n4428) );
  OR2_X1 U6051 ( .A1(n8728), .A2(n8458), .ZN(n4429) );
  OAI21_X1 U6052 ( .B1(n6189), .B2(n8481), .A(n4980), .ZN(n8471) );
  INV_X1 U6053 ( .A(n5849), .ZN(n4676) );
  NAND2_X1 U6054 ( .A1(n9960), .A2(n6493), .ZN(n9940) );
  AND2_X1 U6055 ( .A1(n4740), .A2(n4739), .ZN(n8470) );
  AND2_X1 U6056 ( .A1(n5875), .A2(n4661), .ZN(n4430) );
  AND3_X1 U6057 ( .A1(n6944), .A2(n7963), .A3(n9223), .ZN(n4431) );
  INV_X1 U6058 ( .A(n6513), .ZN(n4952) );
  NAND2_X1 U6059 ( .A1(n5206), .A2(n5207), .ZN(n5300) );
  NAND2_X1 U6060 ( .A1(n5164), .A2(n5163), .ZN(n5167) );
  INV_X1 U6061 ( .A(n5167), .ZN(n4833) );
  AND2_X1 U6062 ( .A1(n9369), .A2(n9546), .ZN(n4432) );
  NAND2_X1 U6063 ( .A1(n10361), .A2(n9216), .ZN(n9489) );
  AND2_X1 U6064 ( .A1(n5049), .A2(n4415), .ZN(n4433) );
  OR3_X1 U6065 ( .A1(n5906), .A2(n6200), .A3(n5905), .ZN(n4434) );
  AND2_X1 U6066 ( .A1(n4419), .A2(n6966), .ZN(n4435) );
  INV_X1 U6067 ( .A(n7714), .ZN(n4875) );
  XNOR2_X1 U6068 ( .A(n5156), .B(SI_15_), .ZN(n5513) );
  AND2_X1 U6069 ( .A1(n4410), .A2(n5055), .ZN(n4436) );
  OR2_X1 U6070 ( .A1(n5094), .A2(n5940), .ZN(n4437) );
  AND2_X1 U6071 ( .A1(n4642), .A2(n6570), .ZN(n4438) );
  INV_X1 U6072 ( .A(n8430), .ZN(n8429) );
  NAND2_X1 U6073 ( .A1(n5060), .A2(n5059), .ZN(n4439) );
  AND2_X1 U6074 ( .A1(n9484), .A2(n9485), .ZN(n4440) );
  NOR2_X1 U6075 ( .A1(n7490), .A2(n4861), .ZN(n4441) );
  AND2_X1 U6076 ( .A1(n5047), .A2(n4415), .ZN(n4442) );
  NAND2_X1 U6077 ( .A1(n10018), .A2(n10416), .ZN(n9347) );
  AND2_X1 U6078 ( .A1(n5524), .A2(n6181), .ZN(n8560) );
  AND2_X1 U6079 ( .A1(n9504), .A2(n5003), .ZN(n4443) );
  NOR2_X1 U6080 ( .A1(n5315), .A2(n10446), .ZN(n4444) );
  INV_X1 U6081 ( .A(n9715), .ZN(n10236) );
  NAND2_X1 U6082 ( .A1(n6072), .A2(n6071), .ZN(n9715) );
  AND2_X1 U6083 ( .A1(n4400), .A2(n4429), .ZN(n4445) );
  NAND2_X1 U6084 ( .A1(n4940), .A2(n4941), .ZN(n4446) );
  NAND2_X1 U6085 ( .A1(n9427), .A2(n9429), .ZN(n4447) );
  NAND2_X1 U6086 ( .A1(n4898), .A2(n4896), .ZN(n4448) );
  INV_X1 U6087 ( .A(n5896), .ZN(n4685) );
  AND2_X1 U6088 ( .A1(n4632), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4449) );
  AND2_X1 U6089 ( .A1(n4598), .A2(n4784), .ZN(n4450) );
  NOR2_X1 U6090 ( .A1(n9955), .A2(n9929), .ZN(n4451) );
  INV_X1 U6091 ( .A(n6182), .ZN(n8534) );
  AND2_X1 U6092 ( .A1(n5056), .A2(n4410), .ZN(n4452) );
  AND2_X1 U6093 ( .A1(n5762), .A2(n5747), .ZN(n4453) );
  INV_X1 U6094 ( .A(n4995), .ZN(n4994) );
  OR2_X1 U6095 ( .A1(n6195), .A2(n4996), .ZN(n4995) );
  AND2_X1 U6096 ( .A1(n8785), .A2(n8556), .ZN(n5870) );
  AND2_X1 U6097 ( .A1(n5834), .A2(n5623), .ZN(n4454) );
  INV_X1 U6098 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5932) );
  AND2_X1 U6099 ( .A1(n6308), .A2(n6310), .ZN(n4455) );
  NOR2_X1 U6100 ( .A1(n8182), .A2(n8557), .ZN(n4456) );
  NAND2_X1 U6101 ( .A1(n6809), .A2(n8139), .ZN(n4457) );
  INV_X1 U6102 ( .A(n4973), .ZN(n4972) );
  NAND2_X1 U6103 ( .A1(n5091), .A2(n6167), .ZN(n4973) );
  NAND2_X1 U6104 ( .A1(n10033), .A2(n9343), .ZN(n4458) );
  AND2_X1 U6105 ( .A1(n5763), .A2(n8711), .ZN(n4459) );
  AND2_X1 U6106 ( .A1(n9864), .A2(n9845), .ZN(n4460) );
  AOI21_X1 U6107 ( .B1(n8857), .B2(n5051), .A(n5049), .ZN(n5046) );
  NAND2_X1 U6108 ( .A1(n9380), .A2(n9428), .ZN(n4461) );
  AND2_X1 U6109 ( .A1(n4942), .A2(n8481), .ZN(n4462) );
  AND2_X1 U6110 ( .A1(n5056), .A2(n4436), .ZN(n4463) );
  OAI21_X1 U6111 ( .B1(n8857), .B2(n5049), .A(n5047), .ZN(n8833) );
  NAND2_X1 U6112 ( .A1(n7771), .A2(n7770), .ZN(n4464) );
  NAND2_X1 U6113 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5180), .ZN(n4465) );
  NOR3_X1 U6114 ( .A1(n7946), .A2(n5829), .A3(n5828), .ZN(n4466) );
  INV_X1 U6115 ( .A(n9371), .ZN(n4776) );
  NAND2_X1 U6116 ( .A1(n4398), .A2(n6966), .ZN(n4467) );
  INV_X1 U6117 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6118 ( .A1(n8711), .A2(n8432), .ZN(n4468) );
  NAND2_X1 U6119 ( .A1(n4682), .A2(n5896), .ZN(n8418) );
  OR2_X1 U6120 ( .A1(n9412), .A2(n4380), .ZN(n4469) );
  INV_X1 U6121 ( .A(n9910), .ZN(n6496) );
  AND3_X1 U6122 ( .A1(n5826), .A2(n7696), .A3(n4564), .ZN(n4470) );
  INV_X1 U6123 ( .A(n9524), .ZN(n5011) );
  INV_X1 U6124 ( .A(n7578), .ZN(n4632) );
  INV_X1 U6125 ( .A(n5897), .ZN(n4686) );
  AND2_X1 U6126 ( .A1(n8502), .A2(n5880), .ZN(n4472) );
  INV_X1 U6127 ( .A(n4669), .ZN(n4944) );
  NAND2_X1 U6128 ( .A1(n5879), .A2(n8520), .ZN(n4669) );
  AND2_X1 U6129 ( .A1(n6076), .A2(n6075), .ZN(n9707) );
  INV_X1 U6130 ( .A(n9707), .ZN(n6141) );
  AND2_X1 U6131 ( .A1(n9360), .A2(n9506), .ZN(n9439) );
  INV_X1 U6132 ( .A(n9439), .ZN(n5023) );
  AND2_X1 U6133 ( .A1(n4665), .A2(n7132), .ZN(n4473) );
  NAND2_X1 U6134 ( .A1(n9347), .A2(n10033), .ZN(n9346) );
  INV_X1 U6135 ( .A(n9346), .ZN(n6318) );
  AND2_X1 U6136 ( .A1(n9993), .A2(n10013), .ZN(n4474) );
  AND2_X1 U6137 ( .A1(n5537), .A2(n5830), .ZN(n4475) );
  AND2_X1 U6138 ( .A1(n8509), .A2(n6186), .ZN(n4476) );
  AND2_X1 U6139 ( .A1(n10403), .A2(n10397), .ZN(n4477) );
  AND2_X1 U6140 ( .A1(n5817), .A2(n6206), .ZN(n4478) );
  AND2_X1 U6141 ( .A1(n4754), .A2(n4753), .ZN(n4479) );
  AND2_X1 U6142 ( .A1(n5536), .A2(n8545), .ZN(n4480) );
  NOR2_X1 U6143 ( .A1(n5543), .A2(n4833), .ZN(n4602) );
  NOR2_X1 U6144 ( .A1(n9757), .A2(n9392), .ZN(n5015) );
  AND2_X1 U6145 ( .A1(n9419), .A2(n9715), .ZN(n4481) );
  AND2_X1 U6146 ( .A1(n5887), .A2(n4427), .ZN(n4482) );
  NAND2_X1 U6147 ( .A1(n6141), .A2(n9423), .ZN(n4483) );
  NAND2_X1 U6148 ( .A1(n5561), .A2(n6846), .ZN(n4484) );
  INV_X1 U6149 ( .A(n9823), .ZN(n9817) );
  AND2_X1 U6150 ( .A1(n6505), .A2(n9376), .ZN(n9823) );
  AND2_X1 U6151 ( .A1(n5834), .A2(n8481), .ZN(n4485) );
  INV_X1 U6152 ( .A(n4925), .ZN(n4924) );
  NAND2_X1 U6153 ( .A1(n4926), .A2(n7696), .ZN(n4925) );
  OR2_X1 U6154 ( .A1(n9443), .A2(n4514), .ZN(n4486) );
  INV_X1 U6155 ( .A(n4624), .ZN(n4623) );
  OR2_X1 U6156 ( .A1(n6514), .A2(n4625), .ZN(n4624) );
  INV_X1 U6157 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5979) );
  INV_X1 U6158 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U6159 ( .A1(n10062), .A2(n5986), .ZN(n10039) );
  INV_X1 U6160 ( .A(n10153), .ZN(n4891) );
  NAND2_X1 U6161 ( .A1(n6066), .A2(n6065), .ZN(n7106) );
  INV_X1 U6162 ( .A(n6671), .ZN(n7928) );
  NAND2_X1 U6163 ( .A1(n10364), .A2(n5957), .ZN(n9484) );
  NAND2_X1 U6164 ( .A1(n6114), .A2(n6113), .ZN(n6122) );
  NAND2_X1 U6165 ( .A1(n6480), .A2(n6479), .ZN(n10333) );
  NAND2_X1 U6166 ( .A1(n4660), .A2(n5874), .ZN(n8544) );
  INV_X1 U6167 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n4709) );
  XNOR2_X1 U6168 ( .A(n5404), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7583) );
  OR2_X1 U6169 ( .A1(n6660), .A2(n8684), .ZN(n4487) );
  AND2_X1 U6170 ( .A1(n9820), .A2(n9821), .ZN(n9843) );
  AND2_X1 U6171 ( .A1(n9472), .A2(n5033), .ZN(n4488) );
  NAND2_X1 U6172 ( .A1(n5840), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5912) );
  AOI21_X1 U6173 ( .B1(n7757), .B2(n9489), .A(n9331), .ZN(n5019) );
  AND2_X1 U6174 ( .A1(n4706), .A2(n4705), .ZN(n4489) );
  OR2_X1 U6175 ( .A1(n7583), .A2(n7724), .ZN(n4490) );
  OR2_X1 U6176 ( .A1(n10039), .A2(n4884), .ZN(n4491) );
  AND2_X2 U6177 ( .A1(n7122), .A2(n7121), .ZN(n10508) );
  NAND2_X1 U6178 ( .A1(n5958), .A2(n5957), .ZN(n7759) );
  INV_X1 U6179 ( .A(n10442), .ZN(n10440) );
  INV_X1 U6180 ( .A(n10222), .ZN(n4882) );
  AND2_X1 U6181 ( .A1(n8396), .A2(n4906), .ZN(n4492) );
  NAND2_X1 U6182 ( .A1(n4656), .A2(n5847), .ZN(n7427) );
  NAND2_X1 U6183 ( .A1(n10453), .A2(n4383), .ZN(n8411) );
  INV_X1 U6184 ( .A(n8411), .ZN(n8385) );
  XOR2_X1 U6185 ( .A(n6778), .B(n8303), .Z(n4493) );
  AND2_X1 U6186 ( .A1(n6811), .A2(n8557), .ZN(n4494) );
  AND2_X1 U6187 ( .A1(n4630), .A2(n4629), .ZN(n4495) );
  AND2_X1 U6188 ( .A1(n4699), .A2(n8970), .ZN(n4496) );
  NAND2_X2 U6189 ( .A1(n8013), .A2(n10097), .ZN(n10112) );
  OR2_X1 U6190 ( .A1(n4728), .A2(n6705), .ZN(n4497) );
  INV_X1 U6191 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n4710) );
  INV_X1 U6192 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n4589) );
  INV_X1 U6193 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7355) );
  INV_X1 U6194 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4569) );
  INV_X1 U6195 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4531) );
  INV_X1 U6196 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n4778) );
  INV_X1 U6197 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4859) );
  XNOR2_X1 U6198 ( .A(n6610), .B(n7914), .ZN(n7908) );
  INV_X1 U6199 ( .A(n7914), .ZN(n4895) );
  OAI22_X1 U6200 ( .A1(n8105), .A2(n8005), .B1(n6091), .B2(P1_U3086), .ZN(
        n4693) );
  INV_X1 U6201 ( .A(n6605), .ZN(n4715) );
  NAND2_X1 U6202 ( .A1(n7610), .A2(n6599), .ZN(n6600) );
  OAI21_X1 U6203 ( .B1(n6609), .B2(n4734), .A(n4487), .ZN(n4732) );
  AOI21_X1 U6204 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8360), .A(n8372), .ZN(
        n6614) );
  XNOR2_X1 U6205 ( .A(n6611), .B(n4647), .ZN(n8317) );
  OAI21_X2 U6206 ( .B1(n6179), .B2(n4984), .A(n4982), .ZN(n8535) );
  NAND2_X1 U6207 ( .A1(n6176), .A2(n6175), .ZN(n8569) );
  INV_X2 U6208 ( .A(n5845), .ZN(n4916) );
  NAND2_X1 U6209 ( .A1(n4991), .A2(n4999), .ZN(n8419) );
  NAND2_X1 U6210 ( .A1(n4916), .A2(n7412), .ZN(n6152) );
  NAND2_X1 U6211 ( .A1(n7872), .A2(n6166), .ZN(n6168) );
  OAI21_X1 U6212 ( .B1(n7634), .B2(n4715), .A(n4713), .ZN(n6607) );
  AOI22_X1 U6213 ( .A1(n7922), .A2(n7923), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n7928), .ZN(n6611) );
  NAND3_X1 U6214 ( .A1(n4759), .A2(n10236), .A3(n4760), .ZN(n4766) );
  NAND2_X1 U6215 ( .A1(n9416), .A2(n9450), .ZN(n4498) );
  NAND2_X1 U6216 ( .A1(n4499), .A2(n9823), .ZN(n9375) );
  NAND3_X1 U6217 ( .A1(n9374), .A2(n9427), .A3(n9520), .ZN(n4499) );
  AOI21_X1 U6218 ( .B1(n9413), .B2(n9468), .A(n9466), .ZN(n9415) );
  OR2_X1 U6219 ( .A1(n5401), .A2(n5400), .ZN(n5388) );
  NAND2_X1 U6220 ( .A1(n5106), .A2(n5105), .ZN(n5413) );
  NAND2_X1 U6221 ( .A1(n6819), .A2(n6818), .ZN(n8209) );
  OAI21_X2 U6222 ( .B1(n7713), .B2(n4867), .A(n4869), .ZN(n6792) );
  NAND2_X2 U6223 ( .A1(n8270), .A2(n6845), .ZN(n6853) );
  OAI21_X2 U6224 ( .B1(n8106), .B2(n8107), .A(n6804), .ZN(n8283) );
  NAND2_X1 U6225 ( .A1(n4848), .A2(n8220), .ZN(n4847) );
  NOR2_X2 U6226 ( .A1(n8161), .A2(n6795), .ZN(n6796) );
  NAND2_X1 U6227 ( .A1(n4818), .A2(n5134), .ZN(n5253) );
  OR2_X2 U6228 ( .A1(n8188), .A2(n6814), .ZN(n6815) );
  NAND2_X1 U6229 ( .A1(n5131), .A2(n5438), .ZN(n4818) );
  INV_X1 U6230 ( .A(n8187), .ZN(n6812) );
  NAND2_X1 U6231 ( .A1(n6842), .A2(n8267), .ZN(n8270) );
  NAND2_X1 U6232 ( .A1(n6716), .A2(n10442), .ZN(n6555) );
  AND2_X2 U6233 ( .A1(n4694), .A2(n8028), .ZN(n6716) );
  NAND2_X1 U6234 ( .A1(n4950), .A2(n4947), .ZN(n6723) );
  NAND2_X1 U6235 ( .A1(n4831), .A2(n4828), .ZN(n5624) );
  NAND2_X1 U6236 ( .A1(n6552), .A2(n6551), .ZN(n4878) );
  NOR2_X1 U6237 ( .A1(n6550), .A2(n4878), .ZN(n4877) );
  OAI21_X1 U6238 ( .B1(n4957), .B2(n4949), .A(n4954), .ZN(n4948) );
  NAND2_X2 U6239 ( .A1(n4500), .A2(n5189), .ZN(n8761) );
  NAND2_X1 U6240 ( .A1(n7366), .A2(n5568), .ZN(n4500) );
  AOI21_X1 U6241 ( .B1(n7570), .B2(n7571), .A(n6630), .ZN(n7557) );
  NOR2_X1 U6242 ( .A1(n8400), .A2(n8399), .ZN(n8405) );
  INV_X1 U6243 ( .A(n4846), .ZN(n8106) );
  OAI21_X1 U6244 ( .B1(n4383), .B2(n10447), .A(n4542), .ZN(n6624) );
  NAND2_X2 U6245 ( .A1(n6273), .A2(n6272), .ZN(n10106) );
  OAI211_X2 U6246 ( .C1(n7173), .C2(n9599), .A(n5956), .B(n5955), .ZN(n9216)
         );
  NAND2_X1 U6247 ( .A1(n5788), .A2(n5789), .ZN(n4504) );
  NAND2_X1 U6248 ( .A1(n4594), .A2(n4592), .ZN(n4790) );
  NAND2_X1 U6249 ( .A1(n5485), .A2(n4505), .ZN(n5512) );
  OAI21_X1 U6250 ( .B1(n5563), .B2(n6846), .A(n4786), .ZN(n4785) );
  NAND2_X1 U6251 ( .A1(n4510), .A2(n4508), .ZN(n5453) );
  AOI21_X1 U6252 ( .B1(n5456), .B2(n8597), .A(n6846), .ZN(n4509) );
  OR2_X1 U6253 ( .A1(n5843), .A2(n6236), .ZN(n4789) );
  NAND3_X1 U6254 ( .A1(n5595), .A2(n6846), .A3(n5884), .ZN(n4590) );
  NAND2_X1 U6255 ( .A1(n4812), .A2(n4810), .ZN(n5786) );
  AOI21_X2 U6256 ( .B1(n5065), .B2(n4435), .A(n4511), .ZN(n7980) );
  NAND3_X1 U6257 ( .A1(n9440), .A2(n4519), .A3(n4518), .ZN(n9441) );
  NAND3_X1 U6258 ( .A1(n9365), .A2(n9439), .A3(n4474), .ZN(n4520) );
  NAND2_X1 U6259 ( .A1(n4818), .A2(n4816), .ZN(n4815) );
  INV_X1 U6260 ( .A(n4736), .ZN(n4668) );
  INV_X1 U6261 ( .A(n5322), .ZN(n5103) );
  OAI211_X1 U6262 ( .C1(n8102), .C2(n8101), .A(n4522), .B(n8100), .ZN(P2_U3160) );
  NAND2_X1 U6263 ( .A1(n8102), .A2(n4523), .ZN(n4522) );
  XNOR2_X1 U6264 ( .A(n4640), .B(n8391), .ZN(n4639) );
  NAND2_X1 U6265 ( .A1(n5120), .A2(n5387), .ZN(n5400) );
  AND2_X1 U6266 ( .A1(n9397), .A2(n9396), .ZN(n4533) );
  OAI21_X1 U6267 ( .B1(n9410), .B2(n9409), .A(n9408), .ZN(n9413) );
  NAND2_X1 U6268 ( .A1(n4767), .A2(n4773), .ZN(n9378) );
  NAND2_X1 U6269 ( .A1(n4755), .A2(n4479), .ZN(n9357) );
  NAND2_X1 U6270 ( .A1(n4850), .A2(n4852), .ZN(n4848) );
  NAND2_X1 U6271 ( .A1(n6796), .A2(n6797), .ZN(n4853) );
  NAND3_X1 U6272 ( .A1(n4532), .A2(n5842), .A3(n4434), .ZN(n4603) );
  NAND2_X1 U6273 ( .A1(n5908), .A2(n5907), .ZN(n4532) );
  OAI21_X4 U6274 ( .B1(n4844), .B2(n4837), .A(n4397), .ZN(n5582) );
  OAI211_X1 U6275 ( .C1(n5879), .C2(n4668), .A(n4666), .B(n5888), .ZN(n5890)
         );
  NAND2_X1 U6276 ( .A1(n4679), .A2(n4677), .ZN(n5900) );
  NAND2_X1 U6277 ( .A1(n9398), .A2(n4533), .ZN(n9400) );
  NAND2_X1 U6278 ( .A1(n4534), .A2(n9420), .ZN(n9421) );
  NAND2_X1 U6279 ( .A1(n4535), .A2(n4481), .ZN(n4534) );
  NAND2_X1 U6280 ( .A1(n4760), .A2(n4759), .ZN(n4535) );
  NAND3_X1 U6281 ( .A1(n9405), .A2(n9449), .A3(n4538), .ZN(n4537) );
  OAI21_X1 U6282 ( .B1(n5121), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4541), .ZN(
        n5362) );
  AND2_X1 U6283 ( .A1(n6712), .A2(n4562), .ZN(n4561) );
  AND2_X1 U6284 ( .A1(n7116), .A2(n7115), .ZN(n5082) );
  NAND2_X1 U6285 ( .A1(n9777), .A2(n5015), .ZN(n5012) );
  NAND2_X1 U6286 ( .A1(n9729), .A2(n9524), .ZN(n4691) );
  NAND2_X1 U6287 ( .A1(n5941), .A2(n4559), .ZN(n5276) );
  INV_X1 U6288 ( .A(n6466), .ZN(n9722) );
  INV_X1 U6289 ( .A(n7996), .ZN(n4543) );
  NAND2_X1 U6290 ( .A1(n4543), .A2(n5024), .ZN(n4567) );
  INV_X1 U6291 ( .A(n7475), .ZN(n6761) );
  NAND2_X1 U6292 ( .A1(n7617), .A2(n4641), .ZN(n4913) );
  NAND2_X1 U6293 ( .A1(n4729), .A2(n4561), .ZN(P2_U3201) );
  INV_X1 U6294 ( .A(n6150), .ZN(n6762) );
  NAND2_X1 U6295 ( .A1(n5386), .A2(n5389), .ZN(n4803) );
  XNOR2_X2 U6296 ( .A(n5544), .B(n5540), .ZN(n7366) );
  OAI21_X2 U6297 ( .B1(n5936), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n4550), .ZN(
        n5118) );
  NAND2_X1 U6298 ( .A1(n8235), .A2(n6829), .ZN(n8113) );
  NOR2_X1 U6299 ( .A1(n7379), .A2(n6914), .ZN(n7530) );
  NAND2_X1 U6300 ( .A1(n8169), .A2(n8170), .ZN(n6841) );
  NAND2_X1 U6301 ( .A1(n4554), .A2(n4552), .ZN(P1_U3262) );
  OAI21_X1 U6302 ( .B1(n10332), .B2(n8078), .A(n8859), .ZN(n4553) );
  NAND2_X1 U6303 ( .A1(n8077), .A2(n9540), .ZN(n4554) );
  NAND2_X1 U6304 ( .A1(n6762), .A2(n7475), .ZN(n5281) );
  NAND4_X1 U6305 ( .A1(n9448), .A2(n9479), .A3(n9552), .A4(n9470), .ZN(n9477)
         );
  NOR2_X2 U6306 ( .A1(n5919), .A2(n4939), .ZN(n5191) );
  NAND3_X1 U6307 ( .A1(n5177), .A2(n5183), .A3(n5176), .ZN(n5919) );
  NAND2_X1 U6308 ( .A1(n4560), .A2(n5927), .ZN(P2_U3296) );
  NAND3_X1 U6309 ( .A1(n4655), .A2(n5911), .A3(n4789), .ZN(n4560) );
  XNOR2_X1 U6310 ( .A(n6604), .B(n7637), .ZN(n7634) );
  NAND3_X1 U6311 ( .A1(n5825), .A2(n5827), .A3(n4470), .ZN(n5828) );
  NAND3_X1 U6312 ( .A1(n4466), .A2(n5878), .A3(n4565), .ZN(n5831) );
  NAND2_X1 U6313 ( .A1(n4815), .A2(n5141), .ZN(n5490) );
  OAI21_X2 U6314 ( .B1(n9911), .B2(n9312), .A(n9514), .ZN(n9891) );
  NAND3_X1 U6315 ( .A1(n6355), .A2(n4567), .A3(n5022), .ZN(n9923) );
  NAND3_X1 U6316 ( .A1(n4573), .A2(n6719), .A3(n10014), .ZN(n6721) );
  NAND2_X1 U6317 ( .A1(n6718), .A2(n9445), .ZN(n4573) );
  NAND2_X1 U6318 ( .A1(n4691), .A2(n5009), .ZN(n6717) );
  NAND2_X1 U6319 ( .A1(n5024), .A2(n5023), .ZN(n5022) );
  INV_X8 U6320 ( .A(n7132), .ZN(n5936) );
  NOR2_X2 U6321 ( .A1(n6348), .A2(n6347), .ZN(n6356) );
  AOI21_X1 U6322 ( .B1(n4582), .B2(n4580), .A(n4578), .ZN(n9474) );
  AND2_X1 U6323 ( .A1(n9467), .A2(n9468), .ZN(n4584) );
  NAND3_X1 U6324 ( .A1(n4591), .A2(n4590), .A3(n4485), .ZN(n4594) );
  NAND2_X1 U6325 ( .A1(n5597), .A2(n4478), .ZN(n4591) );
  NAND2_X1 U6326 ( .A1(n5155), .A2(n5154), .ZN(n4597) );
  NAND2_X1 U6327 ( .A1(n5155), .A2(n4596), .ZN(n4595) );
  XNOR2_X1 U6328 ( .A(n4597), .B(n5513), .ZN(n7209) );
  NAND2_X1 U6329 ( .A1(n5211), .A2(n4602), .ZN(n4600) );
  OR2_X2 U6330 ( .A1(n5211), .A2(n5210), .ZN(n4844) );
  OAI21_X1 U6331 ( .B1(n5806), .B2(n5811), .A(n5815), .ZN(n5843) );
  AOI21_X1 U6332 ( .B1(n5843), .B2(n6225), .A(n4603), .ZN(n4655) );
  AND2_X2 U6333 ( .A1(n5026), .A2(n6023), .ZN(n6117) );
  AND2_X2 U6334 ( .A1(n4917), .A2(n5978), .ZN(n6023) );
  AND2_X2 U6335 ( .A1(n5929), .A2(n5027), .ZN(n5026) );
  NAND3_X1 U6336 ( .A1(n9722), .A2(n9718), .A3(n4611), .ZN(n7113) );
  NAND2_X1 U6337 ( .A1(n9922), .A2(n4617), .ZN(n4615) );
  NAND2_X1 U6338 ( .A1(n6510), .A2(n4627), .ZN(n4626) );
  INV_X1 U6339 ( .A(n6581), .ZN(n8357) );
  NAND2_X1 U6340 ( .A1(n8357), .A2(n8356), .ZN(n4898) );
  NAND3_X1 U6341 ( .A1(n4630), .A2(n4629), .A3(n4490), .ZN(n4631) );
  INV_X1 U6342 ( .A(n4631), .ZN(n6576) );
  OAI21_X1 U6343 ( .B1(n8384), .B2(n8661), .A(n4722), .ZN(n4640) );
  INV_X1 U6344 ( .A(n8395), .ZN(n4635) );
  NAND2_X1 U6345 ( .A1(n8397), .A2(n8396), .ZN(n4637) );
  NAND2_X1 U6346 ( .A1(n4634), .A2(n4633), .ZN(n4636) );
  NAND4_X1 U6347 ( .A1(n8410), .A2(n4637), .A3(n4638), .A4(n4636), .ZN(
        P2_U3200) );
  NAND2_X1 U6348 ( .A1(n7561), .A2(n6570), .ZN(n6571) );
  INV_X1 U6349 ( .A(n7157), .ZN(n4642) );
  NAND2_X1 U6350 ( .A1(n4643), .A2(n4644), .ZN(n4910) );
  NAND2_X1 U6351 ( .A1(n7927), .A2(n4407), .ZN(n4643) );
  INV_X1 U6352 ( .A(n4912), .ZN(n8326) );
  INV_X1 U6353 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4650) );
  NAND2_X1 U6354 ( .A1(n4854), .A2(n5308), .ZN(n5380) );
  NAND2_X1 U6355 ( .A1(n5904), .A2(n5903), .ZN(n5908) );
  NAND2_X1 U6356 ( .A1(n8561), .A2(n4430), .ZN(n4657) );
  NAND2_X1 U6357 ( .A1(n4657), .A2(n4658), .ZN(n8533) );
  NAND2_X1 U6358 ( .A1(n6207), .A2(n4473), .ZN(n4664) );
  NAND2_X1 U6359 ( .A1(n4667), .A2(n4736), .ZN(n4666) );
  NAND2_X1 U6360 ( .A1(n5850), .A2(n4674), .ZN(n4673) );
  OAI21_X1 U6361 ( .B1(n5851), .B2(n4675), .A(n7681), .ZN(n4672) );
  NAND2_X1 U6362 ( .A1(n4673), .A2(n4671), .ZN(n7674) );
  NAND2_X1 U6363 ( .A1(n7537), .A2(n5851), .ZN(n7538) );
  NAND2_X1 U6364 ( .A1(n8428), .A2(n4680), .ZN(n4679) );
  NOR2_X2 U6365 ( .A1(n4688), .A2(n4687), .ZN(n5929) );
  NAND4_X1 U6366 ( .A1(n6040), .A2(n6107), .A3(n6105), .A4(n5035), .ZN(n4687)
         );
  NAND4_X1 U6367 ( .A1(n4690), .A2(n4689), .A3(n8934), .A4(n6031), .ZN(n4688)
         );
  AOI21_X2 U6368 ( .B1(n6547), .B2(n10014), .A(n6546), .ZN(n8028) );
  NAND3_X1 U6369 ( .A1(n5026), .A2(n6023), .A3(n5932), .ZN(n6086) );
  NOR2_X1 U6370 ( .A1(n4812), .A2(n5763), .ZN(n5787) );
  OR2_X1 U6371 ( .A1(n5748), .A2(n4791), .ZN(n4697) );
  NAND3_X1 U6372 ( .A1(n7355), .A2(n4701), .A3(n5196), .ZN(n5368) );
  NAND2_X1 U6373 ( .A1(n5204), .A2(n4489), .ZN(n5226) );
  NAND2_X1 U6374 ( .A1(n7551), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U6375 ( .A1(n7564), .A2(n7565), .ZN(n4711) );
  XNOR2_X1 U6376 ( .A(n6613), .B(n6688), .ZN(n8351) );
  AOI21_X1 U6377 ( .B1(n8369), .B2(n8370), .A(n8368), .ZN(n8372) );
  OR2_X1 U6378 ( .A1(n8384), .A2(n4497), .ZN(n4718) );
  NAND3_X1 U6379 ( .A1(n4719), .A2(n4718), .A3(n4717), .ZN(n4730) );
  NAND3_X1 U6380 ( .A1(n8384), .A2(n4724), .A3(n6705), .ZN(n4717) );
  INV_X1 U6381 ( .A(n6614), .ZN(n4723) );
  OAI21_X1 U6382 ( .B1(n6614), .B2(n4726), .A(n4731), .ZN(n4725) );
  OR2_X1 U6383 ( .A1(n6696), .A2(n4727), .ZN(n4726) );
  NOR2_X1 U6384 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4747) );
  NOR2_X1 U6385 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4746) );
  NAND3_X1 U6386 ( .A1(n9088), .A2(n4745), .A3(n4744), .ZN(n5949) );
  AND4_X2 U6387 ( .A1(n5943), .A2(n4748), .A3(n4747), .A4(n4746), .ZN(n5978)
         );
  OAI211_X1 U6388 ( .C1(n9342), .C2(n4751), .A(n9991), .B(n4749), .ZN(n9348)
         );
  INV_X1 U6389 ( .A(n4752), .ZN(n4751) );
  NAND2_X1 U6390 ( .A1(n9346), .A2(n9315), .ZN(n4758) );
  NAND2_X1 U6391 ( .A1(n9417), .A2(n9450), .ZN(n4759) );
  NAND2_X1 U6392 ( .A1(n4762), .A2(n4483), .ZN(n4761) );
  NAND2_X1 U6393 ( .A1(n4764), .A2(n4763), .ZN(n4762) );
  NOR2_X1 U6394 ( .A1(n9473), .A2(n9471), .ZN(n4763) );
  NAND2_X1 U6395 ( .A1(n4766), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U6396 ( .A1(n4772), .A2(n4768), .ZN(n4767) );
  OAI211_X2 U6397 ( .C1(n6390), .C2(n4778), .A(n4455), .B(n6309), .ZN(n9568)
         );
  OAI21_X1 U6398 ( .B1(n5581), .B2(n4785), .A(n5580), .ZN(n5596) );
  NAND2_X1 U6399 ( .A1(n5581), .A2(n4784), .ZN(n4782) );
  NAND3_X1 U6400 ( .A1(n4783), .A2(n4782), .A3(n4787), .ZN(n5597) );
  NAND2_X1 U6401 ( .A1(n5568), .A2(n7134), .ZN(n5422) );
  NAND2_X1 U6402 ( .A1(n7161), .A2(n5568), .ZN(n5443) );
  NAND2_X1 U6403 ( .A1(n7144), .A2(n5568), .ZN(n5394) );
  NAND2_X1 U6404 ( .A1(n7165), .A2(n5568), .ZN(n5256) );
  NAND2_X1 U6405 ( .A1(n7729), .A2(n5568), .ZN(n5613) );
  NAND2_X1 U6406 ( .A1(n7790), .A2(n5568), .ZN(n5636) );
  NAND2_X1 U6407 ( .A1(n7900), .A2(n5568), .ZN(n5653) );
  NAND2_X1 U6408 ( .A1(n7959), .A2(n5568), .ZN(n5674) );
  NAND2_X1 U6409 ( .A1(n7786), .A2(n5568), .ZN(n5588) );
  NAND2_X1 U6410 ( .A1(n7970), .A2(n5568), .ZN(n5716) );
  NAND2_X1 U6411 ( .A1(n7976), .A2(n5568), .ZN(n5698) );
  NAND2_X1 U6412 ( .A1(n8103), .A2(n5568), .ZN(n5761) );
  NAND2_X1 U6413 ( .A1(n8006), .A2(n5568), .ZN(n5775) );
  NAND2_X1 U6414 ( .A1(n8797), .A2(n5568), .ZN(n5798) );
  NAND2_X1 U6415 ( .A1(n5512), .A2(n4796), .ZN(n4792) );
  NAND2_X1 U6416 ( .A1(n4792), .A2(n4793), .ZN(n5538) );
  INV_X1 U6417 ( .A(n5510), .ZN(n4799) );
  NAND2_X1 U6418 ( .A1(n5191), .A2(n5190), .ZN(n5194) );
  NAND2_X1 U6419 ( .A1(n5191), .A2(n4800), .ZN(n8798) );
  NAND2_X1 U6420 ( .A1(n7780), .A2(n7770), .ZN(n5856) );
  INV_X1 U6421 ( .A(n5111), .ZN(n4802) );
  NAND2_X4 U6422 ( .A1(n4805), .A2(n4804), .ZN(n5121) );
  NAND3_X2 U6423 ( .A1(n8078), .A2(n4807), .A3(n4806), .ZN(n4805) );
  NAND2_X1 U6424 ( .A1(n5762), .A2(n4811), .ZN(n4810) );
  INV_X1 U6425 ( .A(n4810), .ZN(n4809) );
  XNOR2_X1 U6426 ( .A(n5766), .B(n4819), .ZN(n8806) );
  XNOR2_X1 U6427 ( .A(n5764), .B(SI_29_), .ZN(n4819) );
  NAND2_X1 U6428 ( .A1(n5729), .A2(n5728), .ZN(n5766) );
  NAND2_X1 U6429 ( .A1(n5713), .A2(n4825), .ZN(n4821) );
  NAND2_X1 U6430 ( .A1(n4821), .A2(n4822), .ZN(n5758) );
  NAND2_X1 U6431 ( .A1(n5713), .A2(n5714), .ZN(n4824) );
  NAND2_X1 U6432 ( .A1(n5211), .A2(n4832), .ZN(n4831) );
  AOI211_X1 U6433 ( .C1(n9478), .C2(n9477), .A(n9476), .B(n9539), .ZN(n9561)
         );
  NAND2_X1 U6434 ( .A1(n5099), .A2(n5098), .ZN(n5307) );
  AND2_X1 U6435 ( .A1(n7349), .A2(n6775), .ZN(n6777) );
  NAND2_X1 U6436 ( .A1(n5237), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4858) );
  OAI21_X2 U6437 ( .B1(n8113), .B2(n6830), .A(n6836), .ZN(n8169) );
  NAND2_X1 U6438 ( .A1(n8283), .A2(n4865), .ZN(n4863) );
  NAND2_X1 U6439 ( .A1(n4863), .A2(n4864), .ZN(n8136) );
  NOR2_X2 U6440 ( .A1(n6815), .A2(n4866), .ZN(n4865) );
  INV_X1 U6441 ( .A(n7713), .ZN(n4876) );
  NAND3_X1 U6442 ( .A1(n5958), .A2(n4395), .A3(n4477), .ZN(n10344) );
  NAND3_X1 U6443 ( .A1(n4879), .A2(n10122), .A3(n10385), .ZN(n10099) );
  INV_X2 U6444 ( .A(n7518), .ZN(n4880) );
  NAND4_X1 U6445 ( .A1(n4890), .A2(n4889), .A3(n4888), .A4(n4887), .ZN(n5928)
         );
  NAND3_X1 U6446 ( .A1(n4898), .A2(n4896), .A3(n6582), .ZN(n6583) );
  NAND3_X1 U6447 ( .A1(n4899), .A2(n6581), .A3(n4897), .ZN(n4896) );
  NAND2_X1 U6448 ( .A1(n4899), .A2(n6581), .ZN(n8342) );
  NAND2_X1 U6449 ( .A1(n4900), .A2(n6688), .ZN(n4899) );
  INV_X1 U6450 ( .A(n6580), .ZN(n4900) );
  NAND2_X1 U6451 ( .A1(n8392), .A2(n4903), .ZN(n4902) );
  NOR2_X1 U6452 ( .A1(n6703), .A2(n4909), .ZN(n4907) );
  NAND2_X1 U6453 ( .A1(n6703), .A2(n4909), .ZN(n4908) );
  INV_X1 U6454 ( .A(n6586), .ZN(n4909) );
  NAND2_X1 U6455 ( .A1(n4910), .A2(n8325), .ZN(n8324) );
  INV_X2 U6456 ( .A(n5264), .ZN(n5315) );
  NAND2_X1 U6457 ( .A1(n8437), .A2(n5894), .ZN(n4915) );
  AND2_X2 U6458 ( .A1(n5281), .A2(n5846), .ZN(n5845) );
  NOR2_X1 U6459 ( .A1(n5928), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n4917) );
  NAND3_X1 U6460 ( .A1(n4919), .A2(n4918), .A3(n5856), .ZN(n7869) );
  NAND2_X1 U6461 ( .A1(n4921), .A2(n4925), .ZN(n4918) );
  NAND2_X1 U6462 ( .A1(n4921), .A2(n7505), .ZN(n4919) );
  AOI21_X2 U6463 ( .B1(n4924), .B2(n4923), .A(n4922), .ZN(n4921) );
  NAND2_X1 U6464 ( .A1(n9961), .A2(n4930), .ZN(n4929) );
  NAND2_X1 U6465 ( .A1(n4935), .A2(n4933), .ZN(n9841) );
  NAND2_X1 U6466 ( .A1(n4938), .A2(n5178), .ZN(n5923) );
  INV_X1 U6467 ( .A(n5919), .ZN(n4938) );
  NAND2_X1 U6468 ( .A1(n4946), .A2(n4945), .ZN(n5872) );
  OR2_X2 U6469 ( .A1(n7947), .A2(n5868), .ZN(n4946) );
  NOR2_X1 U6470 ( .A1(n9444), .A2(n4962), .ZN(n4956) );
  NAND2_X1 U6471 ( .A1(n9758), .A2(n4951), .ZN(n4950) );
  OR2_X1 U6472 ( .A1(n10153), .A2(n9762), .ZN(n4964) );
  NAND3_X1 U6473 ( .A1(n4966), .A2(n4965), .A3(n5077), .ZN(P2_U3488) );
  NAND2_X1 U6474 ( .A1(n6739), .A2(n7126), .ZN(n4965) );
  NOR2_X1 U6475 ( .A1(n6739), .A2(n6738), .ZN(n7123) );
  NAND2_X1 U6476 ( .A1(n4967), .A2(n4476), .ZN(n8030) );
  NAND2_X1 U6477 ( .A1(n4969), .A2(n4968), .ZN(n7664) );
  NAND2_X1 U6478 ( .A1(n6168), .A2(n4971), .ZN(n4970) );
  NAND2_X1 U6479 ( .A1(n4970), .A2(n6173), .ZN(n6176) );
  NAND2_X1 U6480 ( .A1(n6189), .A2(n4978), .ZN(n4977) );
  NAND2_X1 U6481 ( .A1(n4998), .A2(n4429), .ZN(n4997) );
  NAND2_X1 U6482 ( .A1(n5002), .A2(n4443), .ZN(n6334) );
  NAND3_X1 U6483 ( .A1(n6321), .A2(n10013), .A3(n6320), .ZN(n5002) );
  NAND2_X1 U6484 ( .A1(n6450), .A2(n5009), .ZN(n5005) );
  NAND2_X1 U6485 ( .A1(n6450), .A2(n6449), .ZN(n9727) );
  OAI211_X1 U6486 ( .C1(n6450), .C2(n5008), .A(n5006), .B(n5005), .ZN(n6451)
         );
  NAND2_X1 U6487 ( .A1(n5012), .A2(n5013), .ZN(n9745) );
  NAND2_X1 U6488 ( .A1(n5018), .A2(n5016), .ZN(n10352) );
  AOI21_X1 U6489 ( .B1(n5017), .B2(n9484), .A(n5020), .ZN(n5016) );
  INV_X1 U6490 ( .A(n9489), .ZN(n5017) );
  NAND2_X1 U6491 ( .A1(n9488), .A2(n4440), .ZN(n5018) );
  NAND2_X1 U6492 ( .A1(n9488), .A2(n9485), .ZN(n7757) );
  NAND2_X1 U6493 ( .A1(n6023), .A2(n5929), .ZN(n6115) );
  NAND2_X1 U6494 ( .A1(n5031), .A2(n5028), .ZN(P1_U3266) );
  NAND2_X1 U6495 ( .A1(n6466), .A2(n10112), .ZN(n5031) );
  NOR2_X2 U6496 ( .A1(n7530), .A2(n7529), .ZN(n9211) );
  NAND3_X1 U6497 ( .A1(n9542), .A2(n9541), .A3(n5032), .ZN(n9560) );
  NAND2_X2 U6498 ( .A1(n9187), .A2(n5036), .ZN(n9276) );
  NAND2_X1 U6499 ( .A1(n9200), .A2(n7040), .ZN(n8882) );
  AOI21_X2 U6500 ( .B1(n9201), .B2(n4412), .A(n5038), .ZN(n8816) );
  INV_X1 U6501 ( .A(n5043), .ZN(n8840) );
  INV_X1 U6502 ( .A(n5061), .ZN(n5059) );
  CLKBUF_X1 U6503 ( .A(n5065), .Z(n5062) );
  INV_X1 U6504 ( .A(n6933), .ZN(n7795) );
  INV_X1 U6505 ( .A(n7794), .ZN(n5069) );
  INV_X1 U6506 ( .A(n10099), .ZN(n5958) );
  INV_X1 U6507 ( .A(n5419), .ZN(n5235) );
  AOI21_X1 U6508 ( .B1(n5785), .B2(n6752), .A(n6751), .ZN(n6753) );
  NAND2_X1 U6509 ( .A1(n7113), .A2(n10442), .ZN(n6530) );
  NAND2_X1 U6510 ( .A1(n7113), .A2(n10430), .ZN(n7116) );
  AOI21_X1 U6511 ( .B1(n6853), .B2(n6852), .A(n8281), .ZN(n6854) );
  INV_X1 U6512 ( .A(n8086), .ZN(n6727) );
  AOI21_X2 U6513 ( .B1(n8148), .B2(n6827), .A(n4423), .ZN(n8235) );
  OR2_X1 U6514 ( .A1(n6222), .A2(n6759), .ZN(n6224) );
  NAND4_X2 U6515 ( .A1(n6278), .A2(n6277), .A3(n6276), .A4(n6275), .ZN(n9570)
         );
  NAND2_X1 U6516 ( .A1(n6177), .A2(n5080), .ZN(n6179) );
  OAI21_X1 U6517 ( .B1(n6716), .B2(n7114), .A(n6715), .ZN(P1_U3519) );
  NAND2_X1 U6518 ( .A1(n8881), .A2(n9283), .ZN(n9285) );
  INV_X1 U6519 ( .A(n5207), .ZN(n8807) );
  NAND2_X1 U6520 ( .A1(n6469), .A2(n9572), .ZN(n6470) );
  NAND2_X1 U6521 ( .A1(n5194), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5195) );
  OAI21_X1 U6522 ( .B1(n7479), .B2(n9572), .A(n10122), .ZN(n6271) );
  INV_X1 U6523 ( .A(n6245), .ZN(n8007) );
  AND2_X1 U6524 ( .A1(n6900), .A2(n6899), .ZN(n6901) );
  NAND2_X1 U6525 ( .A1(n7732), .A2(n6881), .ZN(n6883) );
  OAI22_X1 U6526 ( .A1(n6897), .A2(n10122), .B1(n9480), .B2(n7070), .ZN(n6898)
         );
  NAND2_X1 U6527 ( .A1(n8801), .A2(n8807), .ZN(n5297) );
  INV_X2 U6528 ( .A(n10499), .ZN(n10501) );
  INV_X1 U6529 ( .A(n8793), .ZN(n6752) );
  INV_X1 U6530 ( .A(n6236), .ZN(n10457) );
  AND2_X1 U6531 ( .A1(n6263), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5070) );
  INV_X1 U6532 ( .A(n6413), .ZN(n6433) );
  AND2_X1 U6533 ( .A1(n6374), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5071) );
  OR2_X1 U6534 ( .A1(n8023), .A2(n10194), .ZN(n5072) );
  INV_X1 U6535 ( .A(n10194), .ZN(n6526) );
  NAND2_X1 U6536 ( .A1(n8255), .A2(n8190), .ZN(n5073) );
  AND2_X1 U6537 ( .A1(n9472), .A2(n6095), .ZN(n10017) );
  AND2_X1 U6538 ( .A1(n5129), .A2(n5128), .ZN(n5074) );
  AND2_X1 U6539 ( .A1(n8821), .A2(n6526), .ZN(n5075) );
  OR2_X1 U6540 ( .A1(n7127), .A2(n8686), .ZN(n5077) );
  AND4_X1 U6541 ( .A1(n8934), .A2(n6105), .A3(n6104), .A4(n9087), .ZN(n5078)
         );
  AND2_X1 U6542 ( .A1(n9472), .A2(n7280), .ZN(n10356) );
  NAND2_X1 U6543 ( .A1(n9425), .A2(n9547), .ZN(n10014) );
  INV_X1 U6544 ( .A(n6016), .ZN(n9952) );
  AND2_X1 U6545 ( .A1(n8029), .A2(n8032), .ZN(n5079) );
  CLKBUF_X3 U6546 ( .A(n5297), .Z(n5336) );
  OR2_X1 U6547 ( .A1(n8785), .A2(n8296), .ZN(n5080) );
  AND2_X2 U6548 ( .A1(n8012), .A2(n6525), .ZN(n10430) );
  INV_X1 U6549 ( .A(n10430), .ZN(n7114) );
  INV_X1 U6550 ( .A(n5785), .ZN(n7127) );
  AND2_X1 U6551 ( .A1(n5376), .A2(n5361), .ZN(n5083) );
  AND2_X1 U6552 ( .A1(n8892), .A2(n5076), .ZN(n5084) );
  OR2_X1 U6553 ( .A1(n6912), .A2(n6911), .ZN(n5085) );
  INV_X1 U6554 ( .A(n7476), .ZN(n6469) );
  AND2_X1 U6555 ( .A1(n6879), .A2(n6878), .ZN(n5087) );
  NAND2_X1 U6556 ( .A1(n8627), .A2(n7850), .ZN(n5088) );
  AND3_X1 U6557 ( .A1(n5906), .A2(n5909), .A3(n7787), .ZN(n5089) );
  OR2_X1 U6558 ( .A1(n9209), .A2(n9210), .ZN(n5090) );
  OR2_X1 U6559 ( .A1(n8602), .A2(n8298), .ZN(n5091) );
  INV_X1 U6560 ( .A(n9322), .ZN(n9323) );
  AND2_X1 U6561 ( .A1(n9395), .A2(n9759), .ZN(n9396) );
  NAND2_X1 U6562 ( .A1(n9400), .A2(n9399), .ZN(n9410) );
  NAND2_X1 U6563 ( .A1(n5901), .A2(n6846), .ZN(n5782) );
  INV_X1 U6564 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5169) );
  AND2_X1 U6565 ( .A1(n5088), .A2(n5782), .ZN(n5783) );
  OR2_X1 U6566 ( .A1(n6754), .A2(n7690), .ZN(n6758) );
  INV_X1 U6567 ( .A(n7696), .ZN(n6162) );
  NAND2_X1 U6568 ( .A1(n10236), .A2(n4380), .ZN(n9420) );
  INV_X1 U6569 ( .A(n9776), .ZN(n6419) );
  INV_X1 U6570 ( .A(n10064), .ZN(n5986) );
  INV_X1 U6571 ( .A(n7352), .ZN(n6772) );
  INV_X1 U6572 ( .A(n7783), .ZN(n5841) );
  NAND2_X1 U6573 ( .A1(n9952), .A2(n9935), .ZN(n9895) );
  INV_X1 U6574 ( .A(n6462), .ZN(n6463) );
  OR2_X1 U6575 ( .A1(n10105), .A2(n7756), .ZN(n6474) );
  INV_X1 U6576 ( .A(n5598), .ZN(n5604) );
  INV_X1 U6577 ( .A(n5152), .ZN(n5153) );
  XNOR2_X1 U6578 ( .A(n6770), .B(n7344), .ZN(n6774) );
  INV_X1 U6579 ( .A(n8448), .ZN(n6843) );
  OR2_X1 U6580 ( .A1(n6680), .A2(n6678), .ZN(n6579) );
  INV_X1 U6581 ( .A(n5749), .ZN(n5732) );
  OR2_X1 U6582 ( .A1(n8796), .A2(n6746), .ZN(n6867) );
  INV_X1 U6583 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5914) );
  OR2_X1 U6584 ( .A1(n5440), .A2(n5214), .ZN(n5497) );
  INV_X1 U6585 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6296) );
  INV_X1 U6586 ( .A(n9282), .ZN(n9283) );
  INV_X1 U6587 ( .A(n6722), .ZN(n9445) );
  INV_X1 U6588 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7603) );
  INV_X1 U6589 ( .A(n10074), .ZN(n10070) );
  OR2_X1 U6590 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  AND2_X1 U6591 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  NOR2_X1 U6592 ( .A1(n5081), .A2(n5153), .ZN(n5154) );
  NAND2_X1 U6593 ( .A1(n5138), .A2(n5137), .ZN(n5141) );
  NAND2_X1 U6594 ( .A1(n5121), .A2(n7131), .ZN(n5100) );
  INV_X1 U6595 ( .A(n8474), .ZN(n8119) );
  AND2_X1 U6596 ( .A1(n8266), .A2(n6840), .ZN(n8171) );
  INV_X1 U6597 ( .A(n8290), .ZN(n8248) );
  NAND2_X1 U6598 ( .A1(n6857), .A2(n6873), .ZN(n8288) );
  INV_X1 U6599 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5190) );
  INV_X1 U6600 ( .A(n8457), .ZN(n8484) );
  OR2_X1 U6601 ( .A1(n10488), .A2(n10457), .ZN(n8567) );
  INV_X1 U6602 ( .A(n6867), .ZN(n6873) );
  INV_X1 U6603 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5238) );
  INV_X1 U6604 ( .A(n9746), .ZN(n9402) );
  AND2_X1 U6605 ( .A1(n7004), .A2(n7003), .ZN(n8868) );
  INV_X1 U6606 ( .A(n9305), .ZN(n9292) );
  INV_X1 U6607 ( .A(n6380), .ZN(n6423) );
  OR2_X1 U6608 ( .A1(n4377), .A2(n8020), .ZN(n10123) );
  OR2_X1 U6609 ( .A1(n7190), .A2(n4488), .ZN(n6523) );
  INV_X1 U6610 ( .A(n10266), .ZN(n6140) );
  INV_X1 U6611 ( .A(n8821), .ZN(n9721) );
  XNOR2_X1 U6612 ( .A(n5541), .B(SI_18_), .ZN(n5540) );
  NAND2_X1 U6613 ( .A1(n5152), .A2(n5147), .ZN(n5495) );
  OAI21_X1 U6614 ( .B1(n5121), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5100), .ZN(
        n5101) );
  AND2_X1 U6615 ( .A1(n6874), .A2(n6873), .ZN(n8286) );
  INV_X1 U6616 ( .A(n8288), .ZN(n8258) );
  NAND2_X1 U6617 ( .A1(n6870), .A2(n6869), .ZN(n8290) );
  AND2_X1 U6618 ( .A1(n5560), .A2(n5559), .ZN(n8214) );
  OAI21_X1 U6619 ( .B1(n6737), .B2(n7673), .A(n6241), .ZN(n6242) );
  INV_X1 U6620 ( .A(n8686), .ZN(n8673) );
  AND3_X1 U6621 ( .A1(n7120), .A2(n7119), .A3(n7118), .ZN(n7121) );
  AND2_X2 U6622 ( .A1(n6206), .A2(n6871), .ZN(n8692) );
  AND2_X1 U6623 ( .A1(n10457), .A2(n7730), .ZN(n10493) );
  AND2_X1 U6624 ( .A1(n5473), .A2(n5244), .ZN(n6671) );
  OAI222_X1 U6625 ( .A1(n7070), .A2(n7277), .B1(n7076), .B2(n7361), .C1(n4744), 
        .C2(n7175), .ZN(n7273) );
  INV_X1 U6626 ( .A(n9277), .ZN(n9299) );
  INV_X1 U6627 ( .A(n7732), .ZN(n9557) );
  OR2_X1 U6628 ( .A1(n6265), .A2(n6253), .ZN(n6256) );
  INV_X1 U6629 ( .A(n10316), .ZN(n10286) );
  AND2_X1 U6630 ( .A1(n7245), .A2(n6095), .ZN(n10312) );
  INV_X1 U6631 ( .A(n10302), .ZN(n10319) );
  XNOR2_X1 U6632 ( .A(n9711), .B(n9707), .ZN(n6084) );
  NOR2_X1 U6633 ( .A1(n4377), .A2(n8018), .ZN(n10373) );
  OAI22_X1 U6634 ( .A1(n9707), .A2(n10194), .B1(n10442), .B2(n6558), .ZN(n6559) );
  OR2_X1 U6635 ( .A1(n10430), .A2(n9108), .ZN(n6142) );
  AND2_X1 U6636 ( .A1(n9939), .A2(n10401), .ZN(n10225) );
  INV_X1 U6637 ( .A(n10225), .ZN(n10424) );
  INV_X1 U6638 ( .A(n6129), .ZN(n7189) );
  OR2_X1 U6639 ( .A1(n6861), .A2(n6562), .ZN(n6617) );
  INV_X1 U6640 ( .A(n8271), .ZN(n8281) );
  INV_X1 U6641 ( .A(n8263), .ZN(n8293) );
  AND2_X1 U6642 ( .A1(n5805), .A2(n5780), .ZN(n7850) );
  INV_X1 U6643 ( .A(n8496), .ZN(n8473) );
  INV_X1 U6644 ( .A(n8402), .ZN(n8305) );
  INV_X1 U6645 ( .A(n10443), .ZN(n7916) );
  INV_X1 U6646 ( .A(n8396), .ZN(n8389) );
  INV_X1 U6647 ( .A(n6242), .ZN(n6243) );
  NAND2_X1 U6648 ( .A1(n10464), .A2(n7426), .ZN(n8553) );
  NAND2_X1 U6649 ( .A1(n10508), .A2(n10487), .ZN(n8667) );
  NAND2_X1 U6650 ( .A1(n10508), .A2(n10473), .ZN(n8686) );
  OR2_X1 U6651 ( .A1(n10499), .A2(n10497), .ZN(n8775) );
  OR2_X1 U6652 ( .A1(n10499), .A2(n10488), .ZN(n8793) );
  AND2_X1 U6653 ( .A1(n6749), .A2(n6748), .ZN(n10499) );
  AND2_X1 U6654 ( .A1(n7160), .A2(n6219), .ZN(n7193) );
  INV_X1 U6655 ( .A(n7160), .ZN(n8795) );
  INV_X1 U6656 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7300) );
  INV_X1 U6657 ( .A(n7455), .ZN(n7149) );
  AOI21_X1 U6658 ( .B1(n8816), .B2(n7110), .A(n7109), .ZN(n7111) );
  INV_X1 U6659 ( .A(n9256), .ZN(n9302) );
  INV_X1 U6660 ( .A(n7104), .ZN(n9732) );
  INV_X1 U6661 ( .A(n10072), .ZN(n9567) );
  NAND2_X1 U6662 ( .A1(n7177), .A2(n7181), .ZN(n10332) );
  INV_X1 U6663 ( .A(n10372), .ZN(n10101) );
  INV_X1 U6664 ( .A(n10373), .ZN(n10124) );
  INV_X1 U6665 ( .A(n6559), .ZN(n6560) );
  NAND2_X1 U6666 ( .A1(n10442), .A2(n10228), .ZN(n10194) );
  AND2_X2 U6667 ( .A1(n6525), .A2(n6524), .ZN(n10442) );
  INV_X1 U6668 ( .A(n9864), .ZN(n10262) );
  NAND2_X1 U6669 ( .A1(n10430), .A2(n10228), .ZN(n10266) );
  OR2_X1 U6670 ( .A1(n7190), .A2(n7189), .ZN(n10381) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7302) );
  NOR2_X2 U6672 ( .A1(n6617), .A2(P2_U3151), .ZN(P2_U3893) );
  OAI21_X1 U6673 ( .B1(n6561), .B2(n10440), .A(n6560), .ZN(P1_U3553) );
  OAI21_X1 U6674 ( .B1(n6561), .B2(n7114), .A(n6144), .ZN(P1_U3521) );
  INV_X1 U6675 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5092) );
  INV_X1 U6676 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7171) );
  NAND2_X1 U6677 ( .A1(n5121), .A2(n7171), .ZN(n5093) );
  OAI211_X1 U6678 ( .C1(n5121), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n5093), .B(
        SI_1_), .ZN(n5099) );
  INV_X1 U6679 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5094) );
  AND2_X1 U6680 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6681 ( .A1(n5121), .A2(n5095), .ZN(n5941) );
  INV_X1 U6682 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U6683 ( .A1(n5121), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5096) );
  INV_X1 U6684 ( .A(SI_1_), .ZN(n5275) );
  OAI211_X1 U6685 ( .C1(n5121), .C2(n7133), .A(n5096), .B(n5275), .ZN(n5097)
         );
  NAND2_X1 U6686 ( .A1(n5276), .A2(n5097), .ZN(n5098) );
  INV_X1 U6687 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7156) );
  INV_X1 U6688 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7131) );
  XNOR2_X1 U6689 ( .A(n5101), .B(SI_2_), .ZN(n5306) );
  NAND2_X1 U6690 ( .A1(n5307), .A2(n5306), .ZN(n5321) );
  INV_X1 U6691 ( .A(n5101), .ZN(n5102) );
  NAND2_X1 U6692 ( .A1(n5102), .A2(SI_2_), .ZN(n5320) );
  INV_X1 U6693 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7159) );
  INV_X1 U6694 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9094) );
  MUX2_X1 U6695 ( .A(n7159), .B(n9094), .S(n5121), .Z(n5322) );
  NAND2_X1 U6696 ( .A1(n5103), .A2(SI_3_), .ZN(n5344) );
  NAND3_X1 U6697 ( .A1(n5321), .A2(n5320), .A3(n5344), .ZN(n5106) );
  NOR2_X1 U6698 ( .A1(n5103), .A2(SI_3_), .ZN(n5104) );
  NOR2_X1 U6699 ( .A1(n5346), .A2(n5104), .ZN(n5105) );
  INV_X1 U6700 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7154) );
  INV_X1 U6701 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7130) );
  INV_X1 U6702 ( .A(n5362), .ZN(n5109) );
  NAND2_X1 U6703 ( .A1(n5109), .A2(SI_5_), .ZN(n5376) );
  NAND2_X1 U6704 ( .A1(n5107), .A2(SI_4_), .ZN(n5361) );
  NAND2_X1 U6705 ( .A1(n5108), .A2(SI_6_), .ZN(n5415) );
  NAND3_X1 U6706 ( .A1(n5413), .A2(n5083), .A3(n5415), .ZN(n5113) );
  XNOR2_X1 U6707 ( .A(n5108), .B(SI_6_), .ZN(n5378) );
  NOR2_X1 U6708 ( .A1(n5109), .A2(SI_5_), .ZN(n5110) );
  MUX2_X1 U6709 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5121), .Z(n5114) );
  XNOR2_X1 U6710 ( .A(n5114), .B(SI_7_), .ZN(n5417) );
  AOI21_X1 U6711 ( .B1(n5111), .B2(n5415), .A(n5417), .ZN(n5112) );
  NAND2_X1 U6712 ( .A1(n5113), .A2(n5112), .ZN(n5116) );
  NAND2_X1 U6713 ( .A1(n5114), .A2(SI_7_), .ZN(n5115) );
  INV_X1 U6714 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7141) );
  INV_X1 U6715 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7170) );
  INV_X2 U6716 ( .A(n5121), .ZN(n7132) );
  INV_X1 U6717 ( .A(SI_8_), .ZN(n5117) );
  INV_X1 U6718 ( .A(n5118), .ZN(n5119) );
  NAND2_X1 U6719 ( .A1(n5119), .A2(SI_8_), .ZN(n5120) );
  INV_X1 U6720 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7148) );
  INV_X1 U6721 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5122) );
  MUX2_X1 U6722 ( .A(n7148), .B(n5122), .S(n5121), .Z(n5124) );
  INV_X1 U6723 ( .A(SI_9_), .ZN(n5123) );
  NAND2_X1 U6724 ( .A1(n5124), .A2(n5123), .ZN(n5128) );
  INV_X1 U6725 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6726 ( .A1(n5125), .A2(SI_9_), .ZN(n5126) );
  NAND2_X1 U6727 ( .A1(n5128), .A2(n5126), .ZN(n5127) );
  INV_X1 U6728 ( .A(n5127), .ZN(n5389) );
  INV_X1 U6729 ( .A(n5439), .ZN(n5131) );
  INV_X1 U6730 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7162) );
  INV_X1 U6731 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5130) );
  MUX2_X1 U6732 ( .A(n7162), .B(n5130), .S(n5936), .Z(n5132) );
  XNOR2_X1 U6733 ( .A(n5132), .B(SI_10_), .ZN(n5438) );
  INV_X1 U6734 ( .A(n5132), .ZN(n5133) );
  NAND2_X1 U6735 ( .A1(n5133), .A2(SI_10_), .ZN(n5134) );
  INV_X1 U6736 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5136) );
  INV_X1 U6737 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5135) );
  MUX2_X1 U6738 ( .A(n5136), .B(n5135), .S(n5936), .Z(n5138) );
  INV_X1 U6739 ( .A(SI_11_), .ZN(n5137) );
  INV_X1 U6740 ( .A(n5138), .ZN(n5139) );
  NAND2_X1 U6741 ( .A1(n5139), .A2(SI_11_), .ZN(n5140) );
  NAND2_X1 U6742 ( .A1(n5141), .A2(n5140), .ZN(n5252) );
  INV_X1 U6743 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7188) );
  INV_X1 U6744 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7186) );
  MUX2_X1 U6745 ( .A(n7188), .B(n7186), .S(n5936), .Z(n5142) );
  INV_X1 U6746 ( .A(n5142), .ZN(n5143) );
  NAND2_X1 U6747 ( .A1(n5143), .A2(SI_12_), .ZN(n5469) );
  MUX2_X1 U6748 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5936), .Z(n5151) );
  NAND2_X1 U6749 ( .A1(n5151), .A2(SI_13_), .ZN(n5150) );
  AND2_X1 U6750 ( .A1(n5469), .A2(n5150), .ZN(n5491) );
  MUX2_X1 U6751 ( .A(n7205), .B(n9171), .S(n5936), .Z(n5145) );
  INV_X1 U6752 ( .A(SI_14_), .ZN(n5144) );
  INV_X1 U6753 ( .A(n5145), .ZN(n5146) );
  NAND2_X1 U6754 ( .A1(n5146), .A2(SI_14_), .ZN(n5147) );
  INV_X1 U6755 ( .A(n5495), .ZN(n5148) );
  NAND2_X1 U6756 ( .A1(n5470), .A2(n5149), .ZN(n5155) );
  MUX2_X1 U6757 ( .A(n9107), .B(n8944), .S(n5936), .Z(n5156) );
  INV_X1 U6758 ( .A(n5156), .ZN(n5157) );
  NAND2_X1 U6759 ( .A1(n5157), .A2(SI_15_), .ZN(n5158) );
  MUX2_X1 U6760 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n5936), .Z(n5160) );
  NAND2_X1 U6761 ( .A1(n5526), .A2(n5159), .ZN(n5162) );
  NAND2_X1 U6762 ( .A1(n5160), .A2(SI_16_), .ZN(n5161) );
  MUX2_X1 U6763 ( .A(n7300), .B(n7302), .S(n5936), .Z(n5164) );
  INV_X1 U6764 ( .A(SI_17_), .ZN(n5163) );
  INV_X1 U6765 ( .A(n5164), .ZN(n5165) );
  NAND2_X1 U6766 ( .A1(n5165), .A2(SI_17_), .ZN(n5166) );
  MUX2_X1 U6767 ( .A(n9074), .B(n8948), .S(n5936), .Z(n5541) );
  INV_X1 U6768 ( .A(n5380), .ZN(n5177) );
  NOR2_X1 U6769 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5173) );
  NAND4_X1 U6770 ( .A1(n5173), .A2(n5172), .A3(n5186), .A4(n5182), .ZN(n5232)
         );
  NAND4_X1 U6771 ( .A1(n5174), .A2(n9055), .A3(n5915), .A4(n5914), .ZN(n5175)
         );
  NOR2_X1 U6772 ( .A1(n5232), .A2(n5175), .ZN(n5176) );
  INV_X1 U6773 ( .A(n5191), .ZN(n5181) );
  NAND2_X1 U6774 ( .A1(n5181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5179) );
  XNOR2_X2 U6775 ( .A(n5179), .B(n5190), .ZN(n6708) );
  INV_X4 U6776 ( .A(n4379), .ZN(n5568) );
  NOR2_X2 U6777 ( .A1(n5419), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5402) );
  AND2_X2 U6778 ( .A1(n5402), .A2(n5182), .ZN(n5212) );
  BUF_X1 U6779 ( .A(n5183), .Z(n5233) );
  AND2_X2 U6780 ( .A1(n5212), .A2(n5233), .ZN(n5187) );
  INV_X1 U6781 ( .A(n5187), .ZN(n5184) );
  NAND2_X1 U6782 ( .A1(n5184), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5185) );
  MUX2_X1 U6783 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5185), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n5188) );
  NAND2_X1 U6784 ( .A1(n5188), .A2(n5549), .ZN(n8406) );
  INV_X1 U6785 ( .A(n8406), .ZN(n6615) );
  AOI22_X1 U6786 ( .A1(n5569), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6564), .B2(
        n6615), .ZN(n5189) );
  XNOR2_X2 U6787 ( .A(n5195), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5207) );
  INV_X1 U6788 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8529) );
  INV_X1 U6789 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6790 ( .A1(n5226), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6791 ( .A1(n5554), .A2(n5205), .ZN(n8530) );
  INV_X1 U6792 ( .A(n8801), .ZN(n5206) );
  NAND2_X1 U6793 ( .A1(n8530), .A2(n5751), .ZN(n5209) );
  AOI22_X1 U6794 ( .A1(n5752), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n5799), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n5208) );
  OAI211_X1 U6795 ( .C1(n5800), .C2(n8529), .A(n5209), .B(n5208), .ZN(n8536)
         );
  INV_X1 U6796 ( .A(n8536), .ZN(n8139) );
  NAND2_X1 U6797 ( .A1(n8761), .A2(n8139), .ZN(n8520) );
  NAND2_X1 U6798 ( .A1(n7299), .A2(n5568), .ZN(n5224) );
  INV_X1 U6799 ( .A(n5212), .ZN(n5391) );
  INV_X1 U6800 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9170) );
  INV_X1 U6801 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9053) );
  NAND4_X1 U6802 ( .A1(n5241), .A2(n9170), .A3(n9053), .A4(n5213), .ZN(n5214)
         );
  INV_X1 U6803 ( .A(n5497), .ZN(n5216) );
  NAND2_X1 U6804 ( .A1(n5216), .A2(n5215), .ZN(n5514) );
  INV_X1 U6805 ( .A(n5514), .ZN(n5218) );
  NAND2_X1 U6806 ( .A1(n5218), .A2(n5217), .ZN(n5219) );
  NAND2_X1 U6807 ( .A1(n5219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U6808 ( .A1(n5527), .A2(n5220), .ZN(n5221) );
  NAND2_X1 U6809 ( .A1(n5221), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5222) );
  XNOR2_X1 U6810 ( .A(n5222), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6696) );
  AOI22_X1 U6811 ( .A1(n6696), .A2(n6564), .B1(n5569), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6812 ( .A1(n5532), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6813 ( .A1(n5226), .A2(n5225), .ZN(n8541) );
  NAND2_X1 U6814 ( .A1(n8541), .A2(n5751), .ZN(n5229) );
  AOI22_X1 U6815 ( .A1(n5752), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n5799), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6816 ( .A1(n5776), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6817 ( .A1(n8767), .A2(n8261), .ZN(n5877) );
  NAND2_X1 U6818 ( .A1(n8520), .A2(n5877), .ZN(n5832) );
  OAI21_X2 U6819 ( .B1(n5549), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5807) );
  INV_X1 U6820 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6821 ( .A1(n5807), .A2(n5230), .ZN(n5809) );
  INV_X1 U6822 ( .A(n5232), .ZN(n5234) );
  NAND2_X1 U6823 ( .A1(n5237), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5236) );
  MUX2_X1 U6824 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5236), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n5239) );
  INV_X2 U6825 ( .A(n6846), .ZN(n6206) );
  NAND2_X1 U6826 ( .A1(n5832), .A2(n6206), .ZN(n5539) );
  NAND2_X1 U6827 ( .A1(n7185), .A2(n5568), .ZN(n5246) );
  OAI21_X1 U6828 ( .B1(n5440), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6829 ( .A1(n5254), .A2(n5241), .ZN(n5242) );
  NAND2_X1 U6830 ( .A1(n5242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6831 ( .A1(n5243), .A2(n9170), .ZN(n5473) );
  OR2_X1 U6832 ( .A1(n5243), .A2(n9170), .ZN(n5244) );
  AOI22_X1 U6833 ( .A1(n6671), .A2(n6564), .B1(n5569), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6834 ( .A1(n5799), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6835 ( .A1(n5776), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6836 ( .A1(n5257), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5247) );
  AND2_X1 U6837 ( .A1(n5478), .A2(n5247), .ZN(n8586) );
  OR2_X1 U6838 ( .A1(n5733), .A2(n8586), .ZN(n5249) );
  INV_X1 U6839 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6669) );
  OR2_X1 U6840 ( .A1(n5315), .A2(n6669), .ZN(n5248) );
  NAND4_X1 U6841 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n8297)
         );
  NAND2_X1 U6842 ( .A1(n8677), .A2(n8246), .ZN(n5466) );
  XNOR2_X1 U6843 ( .A(n5253), .B(n5252), .ZN(n7165) );
  XNOR2_X1 U6844 ( .A(n5254), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7914) );
  AOI22_X1 U6845 ( .A1(n5569), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7914), .B2(
        n6564), .ZN(n5255) );
  NAND2_X1 U6846 ( .A1(n5752), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5262) );
  INV_X1 U6847 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7897) );
  OR2_X1 U6848 ( .A1(n5336), .A2(n7897), .ZN(n5261) );
  OAI21_X1 U6849 ( .B1(n5444), .B2(P2_REG3_REG_10__SCAN_IN), .A(
        P2_REG3_REG_11__SCAN_IN), .ZN(n5258) );
  AND2_X1 U6850 ( .A1(n5258), .A2(n5257), .ZN(n8247) );
  OR2_X1 U6851 ( .A1(n5733), .A2(n8247), .ZN(n5260) );
  INV_X1 U6852 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7903) );
  OR2_X1 U6853 ( .A1(n5800), .A2(n7903), .ZN(n5259) );
  NAND2_X1 U6854 ( .A1(n8579), .A2(n8157), .ZN(n5863) );
  NAND2_X1 U6855 ( .A1(n5466), .A2(n5863), .ZN(n5263) );
  NAND2_X1 U6856 ( .A1(n5263), .A2(n5867), .ZN(n5486) );
  NAND2_X1 U6857 ( .A1(n5486), .A2(n6206), .ZN(n5468) );
  INV_X1 U6858 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7468) );
  INV_X1 U6859 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7473) );
  INV_X1 U6860 ( .A(n5297), .ZN(n5265) );
  NAND2_X1 U6861 ( .A1(n5265), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5266) );
  AND4_X2 U6862 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n6150)
         );
  INV_X1 U6863 ( .A(n6708), .ZN(n6204) );
  AND2_X1 U6864 ( .A1(n5936), .A2(n7133), .ZN(n5270) );
  OAI21_X1 U6865 ( .B1(n6204), .B2(n6203), .A(n5270), .ZN(n5274) );
  NAND2_X1 U6866 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5272) );
  INV_X1 U6867 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5271) );
  XNOR2_X2 U6868 ( .A(n5272), .B(n5271), .ZN(n7386) );
  NAND3_X1 U6869 ( .A1(n6708), .A2(n4383), .A3(n7386), .ZN(n5273) );
  AND2_X1 U6870 ( .A1(n5274), .A2(n5273), .ZN(n5280) );
  XNOR2_X1 U6871 ( .A(n5276), .B(n5275), .ZN(n5278) );
  XNOR2_X1 U6872 ( .A(n5278), .B(n5277), .ZN(n7172) );
  NAND2_X1 U6873 ( .A1(n5305), .A2(n7172), .ZN(n5279) );
  INV_X1 U6874 ( .A(n5281), .ZN(n5290) );
  INV_X1 U6875 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5282) );
  INV_X1 U6876 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10447) );
  OR2_X1 U6877 ( .A1(n5298), .A2(n10447), .ZN(n5285) );
  INV_X1 U6878 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5283) );
  OR2_X1 U6879 ( .A1(n5300), .A2(n5283), .ZN(n5284) );
  INV_X1 U6880 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10446) );
  INV_X1 U6881 ( .A(SI_0_), .ZN(n5940) );
  NOR2_X1 U6882 ( .A1(n5936), .A2(n5940), .ZN(n5287) );
  XNOR2_X1 U6883 ( .A(n5287), .B(n5094), .ZN(n8813) );
  INV_X1 U6884 ( .A(n10472), .ZN(n5291) );
  AND2_X1 U6885 ( .A1(n8306), .A2(n5291), .ZN(n5820) );
  MUX2_X1 U6886 ( .A(n5290), .B(n5289), .S(n6206), .Z(n5334) );
  NAND2_X1 U6887 ( .A1(n7337), .A2(n10472), .ZN(n7415) );
  NAND2_X1 U6888 ( .A1(n7415), .A2(n7787), .ZN(n5293) );
  NAND3_X1 U6889 ( .A1(n8306), .A2(n5291), .A3(n7730), .ZN(n5292) );
  NAND2_X1 U6890 ( .A1(n5293), .A2(n5292), .ZN(n5295) );
  NAND2_X1 U6891 ( .A1(n5295), .A2(n5294), .ZN(n5312) );
  NAND2_X1 U6892 ( .A1(n5264), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5304) );
  INV_X1 U6893 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5296) );
  INV_X1 U6894 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6566) );
  OR2_X1 U6895 ( .A1(n5298), .A2(n6566), .ZN(n5302) );
  INV_X1 U6896 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5299) );
  OR2_X1 U6897 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  AND4_X2 U6898 ( .A1(n5304), .A2(n5303), .A3(n5302), .A4(n5301), .ZN(n7336)
         );
  XNOR2_X1 U6899 ( .A(n5306), .B(n5307), .ZN(n7155) );
  INV_X1 U6900 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6901 ( .A1(n5308), .A2(n5309), .ZN(n5349) );
  NAND2_X2 U6902 ( .A1(n5349), .A2(n5310), .ZN(n6567) );
  INV_X1 U6903 ( .A(n6567), .ZN(n6628) );
  NAND2_X1 U6904 ( .A1(n7336), .A2(n5311), .ZN(n5847) );
  INV_X1 U6905 ( .A(n7336), .ZN(n7345) );
  NAND2_X1 U6906 ( .A1(n7345), .A2(n7328), .ZN(n5328) );
  NAND2_X1 U6907 ( .A1(n5312), .A2(n8687), .ZN(n5333) );
  INV_X1 U6908 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5313) );
  INV_X1 U6909 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5314) );
  OR2_X1 U6910 ( .A1(n5315), .A2(n5314), .ZN(n5318) );
  INV_X1 U6911 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7550) );
  OR2_X1 U6912 ( .A1(n5298), .A2(n7550), .ZN(n5317) );
  OR2_X1 U6913 ( .A1(n5300), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6914 ( .A1(n5321), .A2(n5320), .ZN(n5343) );
  XNOR2_X1 U6915 ( .A(n5322), .B(SI_3_), .ZN(n5342) );
  XNOR2_X1 U6916 ( .A(n5343), .B(n5342), .ZN(n7158) );
  NOR2_X1 U6917 ( .A1(n7158), .A2(n4379), .ZN(n5327) );
  NAND2_X1 U6918 ( .A1(n5349), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5324) );
  INV_X1 U6919 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5323) );
  XNOR2_X2 U6920 ( .A(n5324), .B(n5323), .ZN(n7157) );
  OAI22_X1 U6921 ( .A1(n5325), .A2(n7159), .B1(n6207), .B2(n7157), .ZN(n5326)
         );
  OR2_X1 U6922 ( .A1(n5327), .A2(n5326), .ZN(n7431) );
  NAND2_X1 U6923 ( .A1(n6771), .A2(n7344), .ZN(n5819) );
  NAND2_X1 U6924 ( .A1(n5819), .A2(n5328), .ZN(n5330) );
  NAND2_X1 U6925 ( .A1(n7329), .A2(n7431), .ZN(n5849) );
  NAND2_X1 U6926 ( .A1(n5849), .A2(n5847), .ZN(n5329) );
  MUX2_X1 U6927 ( .A(n5330), .B(n5329), .S(n6846), .Z(n5331) );
  INV_X1 U6928 ( .A(n5331), .ZN(n5332) );
  OAI21_X1 U6929 ( .B1(n5334), .B2(n5333), .A(n5332), .ZN(n5353) );
  NAND2_X1 U6930 ( .A1(n5752), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5341) );
  INV_X1 U6931 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5335) );
  OR2_X1 U6932 ( .A1(n5336), .A2(n5335), .ZN(n5340) );
  NAND2_X1 U6933 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5337) );
  AND2_X1 U6934 ( .A1(n5354), .A2(n5337), .ZN(n7368) );
  OR2_X1 U6935 ( .A1(n5300), .A2(n7368), .ZN(n5339) );
  INV_X1 U6936 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9140) );
  OR2_X1 U6937 ( .A1(n5298), .A2(n9140), .ZN(n5338) );
  AND4_X2 U6938 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n7348)
         );
  NAND2_X1 U6939 ( .A1(n5343), .A2(n5342), .ZN(n5345) );
  NAND2_X1 U6940 ( .A1(n5345), .A2(n5344), .ZN(n5348) );
  INV_X1 U6941 ( .A(n5346), .ZN(n5347) );
  XNOR2_X1 U6942 ( .A(n5348), .B(n5347), .ZN(n7151) );
  OR2_X1 U6943 ( .A1(n7151), .A2(n4379), .ZN(n5352) );
  NAND2_X1 U6944 ( .A1(n5363), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5350) );
  AOI22_X1 U6945 ( .A1(n5569), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6564), .B2(
        n6631), .ZN(n5351) );
  NAND2_X1 U6946 ( .A1(n5352), .A2(n5351), .ZN(n7545) );
  NAND2_X1 U6947 ( .A1(n7348), .A2(n7545), .ZN(n7675) );
  INV_X1 U6948 ( .A(n7545), .ZN(n6776) );
  NAND2_X1 U6949 ( .A1(n6776), .A2(n8303), .ZN(n5431) );
  NAND2_X1 U6950 ( .A1(n7675), .A2(n5431), .ZN(n7542) );
  INV_X1 U6951 ( .A(n7542), .ZN(n5851) );
  NAND2_X1 U6952 ( .A1(n5353), .A2(n5851), .ZN(n5432) );
  INV_X1 U6953 ( .A(n5819), .ZN(n5367) );
  NAND2_X1 U6954 ( .A1(n5752), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6955 ( .A1(n5776), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6956 ( .A1(n5354), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5355) );
  AND2_X1 U6957 ( .A1(n5368), .A2(n5355), .ZN(n7678) );
  OR2_X1 U6958 ( .A1(n5733), .A2(n7678), .ZN(n5358) );
  INV_X1 U6959 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5356) );
  OR2_X1 U6960 ( .A1(n5336), .A2(n5356), .ZN(n5357) );
  NAND2_X1 U6961 ( .A1(n5413), .A2(n5361), .ZN(n5375) );
  XNOR2_X1 U6962 ( .A(n5362), .B(SI_5_), .ZN(n5374) );
  XNOR2_X1 U6963 ( .A(n5375), .B(n5374), .ZN(n7153) );
  OR2_X1 U6964 ( .A1(n7153), .A2(n4379), .ZN(n5366) );
  OAI21_X1 U6965 ( .B1(n5363), .B2(P2_IR_REG_4__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5364) );
  XNOR2_X1 U6966 ( .A(n5364), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7400) );
  AOI22_X1 U6967 ( .A1(n5569), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6564), .B2(
        n7400), .ZN(n5365) );
  NAND2_X1 U6968 ( .A1(n5366), .A2(n5365), .ZN(n7440) );
  OAI211_X1 U6969 ( .C1(n5432), .C2(n5367), .A(n5852), .B(n7675), .ZN(n5385)
         );
  NAND2_X1 U6970 ( .A1(n5799), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5373) );
  INV_X1 U6971 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6639) );
  OR2_X1 U6972 ( .A1(n5315), .A2(n6639), .ZN(n5372) );
  NAND2_X1 U6973 ( .A1(n5368), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5369) );
  AND2_X1 U6974 ( .A1(n5423), .A2(n5369), .ZN(n7510) );
  OR2_X1 U6975 ( .A1(n5733), .A2(n7510), .ZN(n5371) );
  INV_X1 U6976 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7509) );
  OR2_X1 U6977 ( .A1(n5800), .A2(n7509), .ZN(n5370) );
  NAND2_X1 U6978 ( .A1(n5375), .A2(n5374), .ZN(n5377) );
  NAND2_X1 U6979 ( .A1(n5377), .A2(n5376), .ZN(n5379) );
  XNOR2_X1 U6980 ( .A(n5379), .B(n5378), .ZN(n7142) );
  NAND2_X1 U6981 ( .A1(n7142), .A2(n5568), .ZN(n5384) );
  NAND2_X1 U6982 ( .A1(n5380), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5381) );
  MUX2_X1 U6983 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5381), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5382) );
  AOI22_X1 U6984 ( .A1(n5569), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6564), .B2(
        n7455), .ZN(n5383) );
  NAND2_X1 U6985 ( .A1(n5384), .A2(n5383), .ZN(n7512) );
  INV_X1 U6986 ( .A(n7440), .ZN(n10489) );
  NAND2_X1 U6987 ( .A1(n10489), .A2(n8302), .ZN(n5823) );
  NAND3_X1 U6988 ( .A1(n5385), .A2(n5854), .A3(n5823), .ZN(n5430) );
  NAND2_X1 U6989 ( .A1(n5388), .A2(n5387), .ZN(n5390) );
  NAND2_X1 U6990 ( .A1(n5391), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5392) );
  XNOR2_X1 U6991 ( .A(n5392), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7656) );
  AOI22_X1 U6992 ( .A1(n5569), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6564), .B2(
        n7656), .ZN(n5393) );
  NAND2_X1 U6993 ( .A1(n5394), .A2(n5393), .ZN(n7868) );
  NAND2_X1 U6994 ( .A1(n5799), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5399) );
  INV_X1 U6995 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7883) );
  OR2_X1 U6996 ( .A1(n5315), .A2(n7883), .ZN(n5398) );
  NAND2_X1 U6997 ( .A1(n5408), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5395) );
  AND2_X1 U6998 ( .A1(n5444), .A2(n5395), .ZN(n8616) );
  OR2_X1 U6999 ( .A1(n5733), .A2(n8616), .ZN(n5397) );
  INV_X1 U7000 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6653) );
  OR2_X1 U7001 ( .A1(n5800), .A2(n6653), .ZN(n5396) );
  NAND2_X1 U7002 ( .A1(n7868), .A2(n7776), .ZN(n5857) );
  XNOR2_X1 U7003 ( .A(n5401), .B(n5400), .ZN(n7139) );
  INV_X1 U7004 ( .A(n5402), .ZN(n5403) );
  NAND2_X1 U7005 ( .A1(n5403), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5404) );
  AOI22_X1 U7006 ( .A1(n5569), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6564), .B2(
        n7583), .ZN(n5405) );
  NAND2_X1 U7007 ( .A1(n5752), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U7008 ( .A1(n5425), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5407) );
  AND2_X1 U7009 ( .A1(n5408), .A2(n5407), .ZN(n7777) );
  OR2_X1 U7010 ( .A1(n5733), .A2(n7777), .ZN(n5410) );
  INV_X1 U7011 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7724) );
  OR2_X1 U7012 ( .A1(n5800), .A2(n7724), .ZN(n5409) );
  NAND2_X1 U7013 ( .A1(n5857), .A2(n5856), .ZN(n5412) );
  OR2_X1 U7014 ( .A1(n7770), .A2(n7780), .ZN(n5456) );
  NAND2_X1 U7015 ( .A1(n5413), .A2(n5083), .ZN(n5414) );
  NAND2_X1 U7016 ( .A1(n5416), .A2(n5415), .ZN(n5418) );
  XNOR2_X1 U7017 ( .A(n5418), .B(n5417), .ZN(n7134) );
  NAND2_X1 U7018 ( .A1(n5419), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5420) );
  XNOR2_X1 U7019 ( .A(n5420), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7637) );
  AOI22_X1 U7020 ( .A1(n5569), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6564), .B2(
        n7637), .ZN(n5421) );
  NAND2_X1 U7021 ( .A1(n5752), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5429) );
  INV_X1 U7022 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8902) );
  OR2_X1 U7023 ( .A1(n5336), .A2(n8902), .ZN(n5428) );
  NAND2_X1 U7024 ( .A1(n5423), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5424) );
  AND2_X1 U7025 ( .A1(n5425), .A2(n5424), .ZN(n7813) );
  OR2_X1 U7026 ( .A1(n5733), .A2(n7813), .ZN(n5427) );
  INV_X1 U7027 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9035) );
  OR2_X1 U7028 ( .A1(n5800), .A2(n9035), .ZN(n5426) );
  NAND4_X1 U7029 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n8300)
         );
  NAND2_X1 U7030 ( .A1(n7814), .A2(n8300), .ZN(n7668) );
  INV_X1 U7031 ( .A(n7814), .ZN(n7719) );
  INV_X1 U7032 ( .A(n8300), .ZN(n6163) );
  NAND2_X1 U7033 ( .A1(n7719), .A2(n6163), .ZN(n5450) );
  NOR2_X1 U7034 ( .A1(n5453), .A2(n6162), .ZN(n5434) );
  NAND2_X1 U7035 ( .A1(n7512), .A2(n7700), .ZN(n5853) );
  NAND3_X1 U7036 ( .A1(n5430), .A2(n5434), .A3(n5853), .ZN(n5437) );
  OAI211_X1 U7037 ( .C1(n5432), .C2(n4676), .A(n5823), .B(n5431), .ZN(n5433)
         );
  NAND3_X1 U7038 ( .A1(n5433), .A2(n5853), .A3(n5852), .ZN(n5435) );
  NAND3_X1 U7039 ( .A1(n5435), .A2(n5434), .A3(n5854), .ZN(n5436) );
  MUX2_X1 U7040 ( .A(n5437), .B(n5436), .S(n6206), .Z(n5465) );
  XNOR2_X1 U7041 ( .A(n5439), .B(n5438), .ZN(n7161) );
  NAND2_X1 U7042 ( .A1(n5440), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5441) );
  XNOR2_X1 U7043 ( .A(n5441), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6660) );
  AOI22_X1 U7044 ( .A1(n5569), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6564), .B2(
        n6660), .ZN(n5442) );
  NAND2_X1 U7045 ( .A1(n5443), .A2(n5442), .ZN(n8602) );
  NAND2_X1 U7046 ( .A1(n5752), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U7047 ( .A1(n5776), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5447) );
  INV_X1 U7048 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n8923) );
  OR2_X1 U7049 ( .A1(n5336), .A2(n8923), .ZN(n5446) );
  XNOR2_X1 U7050 ( .A(n5444), .B(n4709), .ZN(n8603) );
  OR2_X1 U7051 ( .A1(n5733), .A2(n8603), .ZN(n5445) );
  NAND4_X1 U7052 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(n8298)
         );
  NAND2_X1 U7053 ( .A1(n8602), .A2(n8156), .ZN(n7892) );
  AND2_X1 U7054 ( .A1(n5857), .A2(n6206), .ZN(n5449) );
  NAND2_X1 U7055 ( .A1(n7892), .A2(n5449), .ZN(n5460) );
  INV_X1 U7056 ( .A(n5856), .ZN(n5452) );
  INV_X1 U7057 ( .A(n5450), .ZN(n5451) );
  OR3_X1 U7058 ( .A1(n5460), .A2(n5452), .A3(n5451), .ZN(n5455) );
  INV_X1 U7059 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U7060 ( .A1(n5455), .A2(n5454), .ZN(n5458) );
  INV_X1 U7061 ( .A(n5458), .ZN(n5461) );
  AND2_X1 U7062 ( .A1(n5456), .A2(n7668), .ZN(n5855) );
  OR2_X1 U7063 ( .A1(n8602), .A2(n8156), .ZN(n5858) );
  AND3_X1 U7064 ( .A1(n5858), .A2(n6846), .A3(n8597), .ZN(n5457) );
  OAI21_X1 U7065 ( .B1(n5458), .B2(n5855), .A(n5457), .ZN(n5459) );
  OAI21_X1 U7066 ( .B1(n5461), .B2(n5460), .A(n5459), .ZN(n5464) );
  MUX2_X1 U7067 ( .A(n7892), .B(n5858), .S(n6206), .Z(n5462) );
  INV_X1 U7068 ( .A(n5462), .ZN(n5463) );
  AOI21_X1 U7069 ( .B1(n5465), .B2(n5464), .A(n5463), .ZN(n5467) );
  NAND2_X1 U7070 ( .A1(n5867), .A2(n5466), .ZN(n8591) );
  XNOR2_X1 U7071 ( .A(n8579), .B(n8607), .ZN(n7893) );
  INV_X1 U7072 ( .A(n7893), .ZN(n8580) );
  NOR2_X1 U7073 ( .A1(n8591), .A2(n8580), .ZN(n5818) );
  MUX2_X1 U7074 ( .A(n5468), .B(n5467), .S(n5818), .Z(n5485) );
  NAND2_X1 U7075 ( .A1(n5470), .A2(n5469), .ZN(n5472) );
  XNOR2_X1 U7076 ( .A(n5472), .B(n5471), .ZN(n7199) );
  NAND2_X1 U7077 ( .A1(n7199), .A2(n5568), .ZN(n5477) );
  NAND2_X1 U7078 ( .A1(n5473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5474) );
  XNOR2_X1 U7079 ( .A(n5474), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6674) );
  INV_X1 U7080 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9141) );
  NOR2_X1 U7081 ( .A1(n5325), .A2(n9141), .ZN(n5475) );
  AOI21_X1 U7082 ( .B1(n6674), .B2(n6564), .A(n5475), .ZN(n5476) );
  INV_X1 U7083 ( .A(n8227), .ZN(n7953) );
  NAND2_X1 U7084 ( .A1(n5752), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U7085 ( .A1(n5776), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5482) );
  INV_X1 U7086 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8946) );
  OR2_X1 U7087 ( .A1(n5336), .A2(n8946), .ZN(n5481) );
  NAND2_X1 U7088 ( .A1(n5478), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5479) );
  AND2_X1 U7089 ( .A1(n5501), .A2(n5479), .ZN(n8225) );
  OR2_X1 U7090 ( .A1(n5733), .A2(n8225), .ZN(n5480) );
  NAND4_X1 U7091 ( .A1(n5483), .A2(n5482), .A3(n5481), .A4(n5480), .ZN(n8583)
         );
  AND2_X1 U7092 ( .A1(n7953), .A2(n8583), .ZN(n5868) );
  INV_X1 U7093 ( .A(n8583), .ZN(n8163) );
  NAND2_X1 U7094 ( .A1(n8227), .A2(n8163), .ZN(n5869) );
  INV_X1 U7095 ( .A(n5869), .ZN(n5507) );
  OR2_X1 U7096 ( .A1(n5868), .A2(n5507), .ZN(n7946) );
  INV_X1 U7097 ( .A(n7946), .ZN(n5484) );
  INV_X1 U7098 ( .A(n5487), .ZN(n5492) );
  OR2_X1 U7099 ( .A1(n5488), .A2(n5492), .ZN(n5489) );
  OR2_X1 U7100 ( .A1(n5490), .A2(n5489), .ZN(n5494) );
  OR2_X1 U7101 ( .A1(n5492), .A2(n5491), .ZN(n5493) );
  NAND2_X1 U7102 ( .A1(n7204), .A2(n5568), .ZN(n5500) );
  NAND2_X1 U7103 ( .A1(n5497), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5498) );
  XNOR2_X1 U7104 ( .A(n5498), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6680) );
  AOI22_X1 U7105 ( .A1(n5569), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6564), .B2(
        n6680), .ZN(n5499) );
  NAND2_X1 U7106 ( .A1(n5799), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7107 ( .A1(n5501), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7108 ( .A1(n5518), .A2(n5502), .ZN(n8574) );
  NAND2_X1 U7109 ( .A1(n5751), .A2(n8574), .ZN(n5505) );
  INV_X1 U7110 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6678) );
  OR2_X1 U7111 ( .A1(n5800), .A2(n6678), .ZN(n5504) );
  INV_X1 U7112 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8672) );
  OR2_X1 U7113 ( .A1(n5315), .A2(n8672), .ZN(n5503) );
  NAND4_X1 U7114 ( .A1(n5506), .A2(n5505), .A3(n5504), .A4(n5503), .ZN(n8296)
         );
  OR2_X1 U7115 ( .A1(n8785), .A2(n8556), .ZN(n5871) );
  INV_X1 U7116 ( .A(n5871), .ZN(n5509) );
  MUX2_X1 U7117 ( .A(n5507), .B(n5868), .S(n6846), .Z(n5508) );
  NOR2_X1 U7118 ( .A1(n8575), .A2(n5508), .ZN(n5511) );
  MUX2_X1 U7119 ( .A(n5870), .B(n5509), .S(n6206), .Z(n5510) );
  NAND2_X1 U7120 ( .A1(n7209), .A2(n5568), .ZN(n5517) );
  NAND2_X1 U7121 ( .A1(n5514), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5515) );
  XNOR2_X1 U7122 ( .A(n5515), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6688) );
  AOI22_X1 U7123 ( .A1(n6688), .A2(n6564), .B1(n5569), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5516) );
  INV_X1 U7124 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U7125 ( .A1(n5518), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7126 ( .A1(n5530), .A2(n5519), .ZN(n8559) );
  NAND2_X1 U7127 ( .A1(n8559), .A2(n5751), .ZN(n5523) );
  INV_X1 U7128 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8669) );
  OR2_X1 U7129 ( .A1(n5315), .A2(n8669), .ZN(n5521) );
  INV_X1 U7130 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8778) );
  OR2_X1 U7131 ( .A1(n5336), .A2(n8778), .ZN(n5520) );
  AND2_X1 U7132 ( .A1(n5521), .A2(n5520), .ZN(n5522) );
  OAI211_X1 U7133 ( .C1(n5800), .C2(n8562), .A(n5523), .B(n5522), .ZN(n8570)
         );
  AND2_X1 U7134 ( .A1(n8779), .A2(n8570), .ZN(n6180) );
  INV_X1 U7135 ( .A(n6180), .ZN(n5524) );
  OR2_X1 U7136 ( .A1(n8779), .A2(n8570), .ZN(n6181) );
  XNOR2_X1 U7137 ( .A(n5526), .B(n5525), .ZN(n7270) );
  NAND2_X1 U7138 ( .A1(n7270), .A2(n5568), .ZN(n5529) );
  XNOR2_X1 U7139 ( .A(n5527), .B(P2_IR_REG_16__SCAN_IN), .ZN(n6692) );
  AOI22_X1 U7140 ( .A1(n6692), .A2(n6564), .B1(n5569), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U7141 ( .A1(n5530), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7142 ( .A1(n5532), .A2(n5531), .ZN(n8550) );
  NAND2_X1 U7143 ( .A1(n8550), .A2(n5751), .ZN(n5535) );
  AOI22_X1 U7144 ( .A1(n5799), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n5776), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7145 ( .A1(n5752), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7146 ( .A1(n8772), .A2(n8557), .ZN(n5875) );
  INV_X1 U7147 ( .A(n8570), .ZN(n6805) );
  OR2_X1 U7148 ( .A1(n8779), .A2(n6805), .ZN(n5874) );
  NAND2_X1 U7149 ( .A1(n8779), .A2(n6805), .ZN(n5873) );
  MUX2_X1 U7150 ( .A(n5874), .B(n5873), .S(n6846), .Z(n5536) );
  MUX2_X1 U7151 ( .A(n5876), .B(n5875), .S(n6206), .Z(n5537) );
  NAND2_X1 U7152 ( .A1(n8522), .A2(n5877), .ZN(n6182) );
  NAND2_X1 U7153 ( .A1(n5539), .A2(n5538), .ZN(n5563) );
  INV_X1 U7154 ( .A(n5541), .ZN(n5542) );
  MUX2_X1 U7155 ( .A(n9061), .B(n7502), .S(n5936), .Z(n5546) );
  INV_X1 U7156 ( .A(SI_19_), .ZN(n5545) );
  INV_X1 U7157 ( .A(n5546), .ZN(n5547) );
  NAND2_X1 U7158 ( .A1(n5547), .A2(SI_19_), .ZN(n5548) );
  NAND2_X1 U7159 ( .A1(n5564), .A2(n5548), .ZN(n5565) );
  XNOR2_X1 U7160 ( .A(n5566), .B(n5565), .ZN(n7501) );
  NAND2_X1 U7161 ( .A1(n7501), .A2(n5568), .ZN(n5553) );
  NAND2_X1 U7162 ( .A1(n5549), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5551) );
  INV_X1 U7163 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5550) );
  XNOR2_X2 U7164 ( .A(n5551), .B(n5550), .ZN(n7503) );
  AOI22_X1 U7165 ( .A1(n5569), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6587), .B2(
        n6564), .ZN(n5552) );
  NAND2_X1 U7166 ( .A1(n5554), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U7167 ( .A1(n5572), .A2(n5555), .ZN(n8517) );
  NAND2_X1 U7168 ( .A1(n8517), .A2(n5751), .ZN(n5560) );
  INV_X1 U7169 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U7170 ( .A1(n5776), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7171 ( .A1(n5799), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5556) );
  OAI211_X1 U7172 ( .C1(n5315), .C2(n8655), .A(n5557), .B(n5556), .ZN(n5558)
         );
  INV_X1 U7173 ( .A(n5558), .ZN(n5559) );
  OR2_X1 U7174 ( .A1(n8761), .A2(n8139), .ZN(n8521) );
  INV_X1 U7175 ( .A(n8520), .ZN(n5561) );
  AND2_X2 U7176 ( .A1(n8521), .A2(n8522), .ZN(n5878) );
  INV_X1 U7177 ( .A(n5878), .ZN(n5562) );
  NAND2_X1 U7178 ( .A1(n8755), .A2(n8214), .ZN(n5880) );
  OAI21_X1 U7179 ( .B1(n5563), .B2(n5562), .A(n5880), .ZN(n5581) );
  INV_X1 U7180 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7692) );
  MUX2_X1 U7181 ( .A(n7692), .B(n7707), .S(n5936), .Z(n5601) );
  XNOR2_X1 U7182 ( .A(n5601), .B(SI_20_), .ZN(n5567) );
  NAND2_X1 U7183 ( .A1(n7689), .A2(n5568), .ZN(n5571) );
  NAND2_X1 U7184 ( .A1(n5569), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5570) );
  INV_X1 U7185 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7186 ( .A1(n5572), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7187 ( .A1(n5590), .A2(n5573), .ZN(n8211) );
  NAND2_X1 U7188 ( .A1(n8211), .A2(n5751), .ZN(n5578) );
  INV_X1 U7189 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U7190 ( .A1(n5776), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7191 ( .A1(n5799), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5574) );
  OAI211_X1 U7192 ( .C1(n5315), .C2(n9132), .A(n5575), .B(n5574), .ZN(n5576)
         );
  INV_X1 U7193 ( .A(n5576), .ZN(n5577) );
  NAND2_X1 U7194 ( .A1(n8041), .A2(n8515), .ZN(n5883) );
  NAND2_X1 U7195 ( .A1(n5883), .A2(n5881), .ZN(n5579) );
  NAND2_X1 U7196 ( .A1(n5579), .A2(n6846), .ZN(n5580) );
  INV_X1 U7197 ( .A(SI_20_), .ZN(n5600) );
  OAI21_X1 U7198 ( .B1(n5582), .B2(n5600), .A(n5601), .ZN(n5584) );
  NAND2_X1 U7199 ( .A1(n5582), .A2(n5600), .ZN(n5583) );
  NAND2_X1 U7200 ( .A1(n5584), .A2(n5583), .ZN(n5586) );
  INV_X1 U7201 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7788) );
  INV_X1 U7202 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7793) );
  MUX2_X1 U7203 ( .A(n7788), .B(n7793), .S(n5936), .Z(n5598) );
  XNOR2_X1 U7204 ( .A(n5598), .B(SI_21_), .ZN(n5585) );
  NAND2_X1 U7205 ( .A1(n5569), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5587) );
  INV_X1 U7206 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U7207 ( .A1(n5590), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7208 ( .A1(n5614), .A2(n5591), .ZN(n8498) );
  INV_X1 U7209 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U7210 ( .A1(n5776), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7211 ( .A1(n5752), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5592) );
  OAI211_X1 U7212 ( .C1(n5336), .C2(n8906), .A(n5593), .B(n5592), .ZN(n5594)
         );
  AOI21_X2 U7213 ( .B1(n8498), .B2(n5751), .A(n5594), .ZN(n8483) );
  NAND2_X1 U7214 ( .A1(n8499), .A2(n8483), .ZN(n5817) );
  INV_X1 U7215 ( .A(n8515), .ZN(n8497) );
  NAND2_X1 U7216 ( .A1(n8216), .A2(n8497), .ZN(n8502) );
  AND2_X1 U7217 ( .A1(n5817), .A2(n8502), .ZN(n5885) );
  NAND2_X1 U7218 ( .A1(n5596), .A2(n5885), .ZN(n5595) );
  INV_X1 U7219 ( .A(n5601), .ZN(n5603) );
  OAI22_X1 U7220 ( .A1(SI_20_), .A2(n5603), .B1(n5604), .B2(SI_21_), .ZN(n5607) );
  INV_X1 U7221 ( .A(SI_21_), .ZN(n5599) );
  OAI21_X1 U7222 ( .B1(n5601), .B2(n5600), .A(n5599), .ZN(n5605) );
  AND2_X1 U7223 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5602) );
  AOI22_X1 U7224 ( .A1(n5605), .A2(n5604), .B1(n5603), .B2(n5602), .ZN(n5606)
         );
  INV_X1 U7225 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7731) );
  MUX2_X1 U7226 ( .A(n7731), .B(n7734), .S(n5936), .Z(n5609) );
  INV_X1 U7227 ( .A(SI_22_), .ZN(n5608) );
  NAND2_X1 U7228 ( .A1(n5609), .A2(n5608), .ZN(n5628) );
  INV_X1 U7229 ( .A(n5609), .ZN(n5610) );
  NAND2_X1 U7230 ( .A1(n5610), .A2(SI_22_), .ZN(n5611) );
  NAND2_X1 U7231 ( .A1(n5628), .A2(n5611), .ZN(n5625) );
  XNOR2_X1 U7232 ( .A(n5624), .B(n5625), .ZN(n7729) );
  NAND2_X1 U7233 ( .A1(n5569), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7234 ( .A1(n5614), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7235 ( .A1(n5637), .A2(n5615), .ZN(n8486) );
  NAND2_X1 U7236 ( .A1(n8486), .A2(n5751), .ZN(n5620) );
  INV_X1 U7237 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U7238 ( .A1(n5752), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7239 ( .A1(n5776), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5616) );
  OAI211_X1 U7240 ( .C1(n5336), .C2(n8745), .A(n5617), .B(n5616), .ZN(n5618)
         );
  INV_X1 U7241 ( .A(n5618), .ZN(n5619) );
  XNOR2_X1 U7242 ( .A(n8230), .B(n8496), .ZN(n8485) );
  NOR2_X1 U7243 ( .A1(n8496), .A2(n6206), .ZN(n5622) );
  AND2_X1 U7244 ( .A1(n8496), .A2(n6206), .ZN(n5621) );
  MUX2_X1 U7245 ( .A(n5622), .B(n5621), .S(n8230), .Z(n5623) );
  INV_X1 U7246 ( .A(n5624), .ZN(n5627) );
  INV_X1 U7247 ( .A(n5625), .ZN(n5626) );
  NAND2_X1 U7248 ( .A1(n5627), .A2(n5626), .ZN(n5629) );
  NAND2_X1 U7249 ( .A1(n5629), .A2(n5628), .ZN(n5645) );
  INV_X1 U7250 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5630) );
  MUX2_X1 U7251 ( .A(n5630), .B(n9062), .S(n5936), .Z(n5632) );
  INV_X1 U7252 ( .A(SI_23_), .ZN(n5631) );
  NAND2_X1 U7253 ( .A1(n5632), .A2(n5631), .ZN(n5646) );
  INV_X1 U7254 ( .A(n5632), .ZN(n5633) );
  NAND2_X1 U7255 ( .A1(n5633), .A2(SI_23_), .ZN(n5634) );
  XNOR2_X1 U7256 ( .A(n5645), .B(n5644), .ZN(n7790) );
  NAND2_X1 U7257 ( .A1(n5569), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7258 ( .A1(n5637), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7259 ( .A1(n5656), .A2(n5638), .ZN(n8477) );
  NAND2_X1 U7260 ( .A1(n8477), .A2(n5751), .ZN(n5643) );
  INV_X1 U7261 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U7262 ( .A1(n5799), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U7263 ( .A1(n5776), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5639) );
  OAI211_X1 U7264 ( .C1(n5315), .C2(n8645), .A(n5640), .B(n5639), .ZN(n5641)
         );
  INV_X1 U7265 ( .A(n5641), .ZN(n5642) );
  NAND2_X1 U7266 ( .A1(n8740), .A2(n8484), .ZN(n8463) );
  NAND2_X1 U7267 ( .A1(n5887), .A2(n8463), .ZN(n8472) );
  NAND2_X1 U7268 ( .A1(n5645), .A2(n5644), .ZN(n5647) );
  NAND2_X1 U7269 ( .A1(n5647), .A2(n5646), .ZN(n5666) );
  INV_X1 U7270 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9073) );
  MUX2_X1 U7271 ( .A(n9073), .B(n9037), .S(n5936), .Z(n5649) );
  INV_X1 U7272 ( .A(SI_24_), .ZN(n5648) );
  NAND2_X1 U7273 ( .A1(n5649), .A2(n5648), .ZN(n5667) );
  INV_X1 U7274 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U7275 ( .A1(n5650), .A2(SI_24_), .ZN(n5651) );
  XNOR2_X1 U7276 ( .A(n5666), .B(n5665), .ZN(n7900) );
  NAND2_X1 U7277 ( .A1(n5569), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5652) );
  INV_X1 U7278 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7279 ( .A1(n5656), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7280 ( .A1(n5675), .A2(n5657), .ZN(n8460) );
  NAND2_X1 U7281 ( .A1(n8460), .A2(n5751), .ZN(n5662) );
  INV_X1 U7282 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U7283 ( .A1(n5799), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5659) );
  INV_X1 U7284 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8467) );
  OR2_X1 U7285 ( .A1(n5800), .A2(n8467), .ZN(n5658) );
  OAI211_X1 U7286 ( .C1(n5315), .C2(n9056), .A(n5659), .B(n5658), .ZN(n5660)
         );
  INV_X1 U7287 ( .A(n5660), .ZN(n5661) );
  AND2_X1 U7288 ( .A1(n5889), .A2(n5887), .ZN(n5663) );
  NAND2_X1 U7289 ( .A1(n8734), .A2(n8119), .ZN(n5816) );
  AND2_X1 U7290 ( .A1(n5816), .A2(n8463), .ZN(n5888) );
  MUX2_X1 U7291 ( .A(n5663), .B(n5888), .S(n6206), .Z(n5664) );
  MUX2_X1 U7292 ( .A(n5816), .B(n5889), .S(n6206), .Z(n5682) );
  NAND2_X1 U7293 ( .A1(n5666), .A2(n5665), .ZN(n5668) );
  NAND2_X1 U7294 ( .A1(n5668), .A2(n5667), .ZN(n5684) );
  INV_X1 U7295 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8009) );
  MUX2_X1 U7296 ( .A(n8009), .B(n9063), .S(n5936), .Z(n5670) );
  INV_X1 U7297 ( .A(SI_25_), .ZN(n5669) );
  NAND2_X1 U7298 ( .A1(n5670), .A2(n5669), .ZN(n5685) );
  INV_X1 U7299 ( .A(n5670), .ZN(n5671) );
  NAND2_X1 U7300 ( .A1(n5671), .A2(SI_25_), .ZN(n5672) );
  XNOR2_X1 U7301 ( .A(n5684), .B(n5683), .ZN(n7959) );
  NAND2_X1 U7302 ( .A1(n5569), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7303 ( .A1(n5675), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7304 ( .A1(n5705), .A2(n5676), .ZN(n8175) );
  NAND2_X1 U7305 ( .A1(n8175), .A2(n5751), .ZN(n5681) );
  INV_X1 U7306 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U7307 ( .A1(n5799), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7308 ( .A1(n5776), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5677) );
  OAI211_X1 U7309 ( .C1(n8640), .C2(n5315), .A(n5678), .B(n5677), .ZN(n5679)
         );
  INV_X1 U7310 ( .A(n5679), .ZN(n5680) );
  NAND2_X1 U7311 ( .A1(n8728), .A2(n8275), .ZN(n5891) );
  NAND2_X1 U7312 ( .A1(n5892), .A2(n5891), .ZN(n8447) );
  NAND2_X1 U7313 ( .A1(n5684), .A2(n5683), .ZN(n5686) );
  INV_X1 U7314 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7972) );
  INV_X1 U7315 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7973) );
  MUX2_X1 U7316 ( .A(n7972), .B(n7973), .S(n5936), .Z(n5688) );
  INV_X1 U7317 ( .A(SI_26_), .ZN(n5687) );
  NAND2_X1 U7318 ( .A1(n5688), .A2(n5687), .ZN(n5691) );
  INV_X1 U7319 ( .A(n5688), .ZN(n5689) );
  NAND2_X1 U7320 ( .A1(n5689), .A2(SI_26_), .ZN(n5690) );
  INV_X1 U7321 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5692) );
  INV_X1 U7322 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7990) );
  MUX2_X1 U7323 ( .A(n5692), .B(n7990), .S(n5936), .Z(n5694) );
  INV_X1 U7324 ( .A(SI_27_), .ZN(n5693) );
  NAND2_X1 U7325 ( .A1(n5694), .A2(n5693), .ZN(n5724) );
  INV_X1 U7326 ( .A(n5694), .ZN(n5695) );
  NAND2_X1 U7327 ( .A1(n5695), .A2(SI_27_), .ZN(n5696) );
  NAND2_X1 U7328 ( .A1(n4529), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5697) );
  NAND2_X2 U7329 ( .A1(n5698), .A2(n5697), .ZN(n8717) );
  INV_X1 U7330 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U7331 ( .A1(n5707), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U7332 ( .A1(n5749), .A2(n5699), .ZN(n8434) );
  NAND2_X1 U7333 ( .A1(n8434), .A2(n5751), .ZN(n5704) );
  INV_X1 U7334 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U7335 ( .A1(n5776), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U7336 ( .A1(n5799), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5700) );
  OAI211_X1 U7337 ( .C1(n5315), .C2(n8634), .A(n5701), .B(n5700), .ZN(n5702)
         );
  INV_X1 U7338 ( .A(n5702), .ZN(n5703) );
  OR2_X2 U7339 ( .A1(n8717), .A2(n8421), .ZN(n5896) );
  NAND2_X1 U7340 ( .A1(n8717), .A2(n8421), .ZN(n5719) );
  NAND2_X1 U7341 ( .A1(n5705), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U7342 ( .A1(n5707), .A2(n5706), .ZN(n8442) );
  NAND2_X1 U7343 ( .A1(n8442), .A2(n5751), .ZN(n5712) );
  INV_X1 U7344 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U7345 ( .A1(n5752), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5709) );
  INV_X1 U7346 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8441) );
  OR2_X1 U7347 ( .A1(n5800), .A2(n8441), .ZN(n5708) );
  OAI211_X1 U7348 ( .C1(n5336), .C2(n9109), .A(n5709), .B(n5708), .ZN(n5710)
         );
  INV_X1 U7349 ( .A(n5710), .ZN(n5711) );
  XNOR2_X1 U7350 ( .A(n5713), .B(n5714), .ZN(n7970) );
  NAND2_X1 U7351 ( .A1(n5569), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5715) );
  NAND2_X2 U7352 ( .A1(n5716), .A2(n5715), .ZN(n8722) );
  INV_X1 U7353 ( .A(n8722), .ZN(n8280) );
  MUX2_X1 U7354 ( .A(n6843), .B(n8280), .S(n6206), .Z(n5744) );
  AND2_X1 U7355 ( .A1(n8448), .A2(n6206), .ZN(n5717) );
  AOI21_X1 U7356 ( .B1(n8722), .B2(n6846), .A(n5717), .ZN(n5718) );
  NAND3_X1 U7357 ( .A1(n5896), .A2(n5719), .A3(n5718), .ZN(n5745) );
  OAI21_X1 U7358 ( .B1(n8430), .B2(n5744), .A(n5745), .ZN(n5721) );
  MUX2_X1 U7359 ( .A(n5892), .B(n5891), .S(n6846), .Z(n5720) );
  NAND2_X1 U7360 ( .A1(n5721), .A2(n5720), .ZN(n5748) );
  INV_X1 U7361 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5725) );
  INV_X1 U7362 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8104) );
  MUX2_X1 U7363 ( .A(n5725), .B(n8104), .S(n5936), .Z(n5727) );
  XNOR2_X1 U7364 ( .A(n5727), .B(SI_28_), .ZN(n5759) );
  NAND2_X1 U7365 ( .A1(n5758), .A2(n5759), .ZN(n5729) );
  INV_X1 U7366 ( .A(SI_28_), .ZN(n5726) );
  NAND2_X1 U7367 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  MUX2_X1 U7368 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5936), .Z(n5764) );
  NAND2_X1 U7369 ( .A1(n5569), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5730) );
  INV_X1 U7370 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5731) );
  INV_X1 U7371 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7124) );
  NAND2_X1 U7372 ( .A1(n5776), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7373 ( .A1(n5799), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5734) );
  OAI211_X1 U7374 ( .C1(n5315), .C2(n7124), .A(n5735), .B(n5734), .ZN(n5736)
         );
  INV_X1 U7375 ( .A(n5736), .ZN(n5737) );
  NAND2_X1 U7376 ( .A1(n8422), .A2(n6206), .ZN(n5738) );
  NAND2_X1 U7377 ( .A1(n6146), .A2(n5738), .ZN(n5740) );
  OR2_X1 U7378 ( .A1(n5785), .A2(n6846), .ZN(n5739) );
  NAND2_X1 U7379 ( .A1(n5740), .A2(n5739), .ZN(n5762) );
  NOR2_X1 U7380 ( .A1(n8421), .A2(n6206), .ZN(n5742) );
  OAI21_X1 U7381 ( .B1(n8440), .B2(n6846), .A(n8717), .ZN(n5741) );
  OAI21_X1 U7382 ( .B1(n5742), .B2(n8717), .A(n5741), .ZN(n5743) );
  OAI21_X1 U7383 ( .B1(n5745), .B2(n5744), .A(n5743), .ZN(n5746) );
  INV_X1 U7384 ( .A(n5746), .ZN(n5747) );
  NAND2_X1 U7385 ( .A1(n5749), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7386 ( .A1(n6237), .A2(n5750), .ZN(n8425) );
  NAND2_X1 U7387 ( .A1(n8425), .A2(n5751), .ZN(n5757) );
  INV_X1 U7388 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9054) );
  NAND2_X1 U7389 ( .A1(n5752), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5754) );
  INV_X1 U7390 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8932) );
  OR2_X1 U7391 ( .A1(n5800), .A2(n8932), .ZN(n5753) );
  OAI211_X1 U7392 ( .C1(n5336), .C2(n9054), .A(n5754), .B(n5753), .ZN(n5755)
         );
  INV_X1 U7393 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U7394 ( .A1(n4529), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5760) );
  MUX2_X1 U7395 ( .A(n8090), .B(n8092), .S(n6846), .Z(n5763) );
  INV_X1 U7396 ( .A(n5764), .ZN(n5765) );
  INV_X1 U7397 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n5769) );
  INV_X1 U7398 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8008) );
  MUX2_X1 U7399 ( .A(n5769), .B(n8008), .S(n5936), .Z(n5771) );
  INV_X1 U7400 ( .A(SI_30_), .ZN(n5770) );
  NAND2_X1 U7401 ( .A1(n5771), .A2(n5770), .ZN(n5791) );
  INV_X1 U7402 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7403 ( .A1(n5772), .A2(SI_30_), .ZN(n5773) );
  NAND2_X1 U7404 ( .A1(n5791), .A2(n5773), .ZN(n5792) );
  NAND2_X1 U7405 ( .A1(n4529), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U7406 ( .A1(n5775), .A2(n5774), .ZN(n8627) );
  INV_X1 U7407 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U7408 ( .A1(n5776), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7409 ( .A1(n5799), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5777) );
  OAI211_X1 U7410 ( .C1(n5315), .C2(n8630), .A(n5778), .B(n5777), .ZN(n5779)
         );
  INV_X1 U7411 ( .A(n5779), .ZN(n5780) );
  OR2_X2 U7412 ( .A1(n8627), .A2(n7850), .ZN(n5901) );
  NAND2_X1 U7413 ( .A1(n5901), .A2(n6146), .ZN(n5838) );
  INV_X1 U7414 ( .A(n5838), .ZN(n5781) );
  NAND2_X1 U7415 ( .A1(n5784), .A2(n5783), .ZN(n5790) );
  NAND2_X1 U7416 ( .A1(n5785), .A2(n8422), .ZN(n6145) );
  NAND2_X1 U7417 ( .A1(n5088), .A2(n6145), .ZN(n5812) );
  AOI21_X1 U7418 ( .B1(n5786), .B2(n8090), .A(n5812), .ZN(n5789) );
  NOR2_X1 U7419 ( .A1(n5787), .A2(n6206), .ZN(n5788) );
  MUX2_X1 U7420 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n5936), .Z(n5794) );
  INV_X1 U7421 ( .A(SI_31_), .ZN(n8908) );
  XNOR2_X1 U7422 ( .A(n5794), .B(n8908), .ZN(n5795) );
  NAND2_X1 U7423 ( .A1(n5569), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5797) );
  NAND2_X2 U7424 ( .A1(n5798), .A2(n5797), .ZN(n8703) );
  INV_X1 U7425 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U7426 ( .A1(n5799), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5802) );
  INV_X1 U7427 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9066) );
  OR2_X1 U7428 ( .A1(n5800), .A2(n9066), .ZN(n5801) );
  OAI211_X1 U7429 ( .C1(n5315), .C2(n8626), .A(n5802), .B(n5801), .ZN(n5803)
         );
  INV_X1 U7430 ( .A(n5803), .ZN(n5804) );
  NOR2_X1 U7431 ( .A1(n8703), .A2(n8413), .ZN(n5811) );
  NAND2_X1 U7432 ( .A1(n8703), .A2(n8413), .ZN(n5815) );
  INV_X1 U7433 ( .A(n5807), .ZN(n5808) );
  NAND2_X1 U7434 ( .A1(n5808), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n5810) );
  NAND2_X2 U7435 ( .A1(n5809), .A2(n5810), .ZN(n7690) );
  NAND2_X1 U7436 ( .A1(n7690), .A2(n6587), .ZN(n6236) );
  INV_X1 U7437 ( .A(n5811), .ZN(n5814) );
  INV_X1 U7438 ( .A(n5812), .ZN(n5813) );
  NAND2_X1 U7439 ( .A1(n5814), .A2(n5813), .ZN(n5898) );
  INV_X1 U7440 ( .A(n5815), .ZN(n5839) );
  NAND2_X1 U7441 ( .A1(n5889), .A2(n5816), .ZN(n8465) );
  INV_X1 U7442 ( .A(n8472), .ZN(n5834) );
  NAND2_X1 U7443 ( .A1(n5884), .A2(n5817), .ZN(n8493) );
  INV_X1 U7444 ( .A(n8493), .ZN(n8504) );
  NAND2_X1 U7445 ( .A1(n5883), .A2(n8502), .ZN(n8029) );
  INV_X1 U7446 ( .A(n8512), .ZN(n8509) );
  INV_X1 U7447 ( .A(n5818), .ZN(n5829) );
  INV_X1 U7448 ( .A(n7429), .ZN(n5848) );
  INV_X1 U7449 ( .A(n5820), .ZN(n5821) );
  NAND2_X1 U7450 ( .A1(n7415), .A2(n5821), .ZN(n10467) );
  NAND4_X1 U7451 ( .A1(n5848), .A2(n5851), .A3(n5822), .A4(n8687), .ZN(n5824)
         );
  AND2_X2 U7452 ( .A1(n5852), .A2(n5823), .ZN(n7681) );
  INV_X1 U7453 ( .A(n7681), .ZN(n7676) );
  NOR2_X1 U7454 ( .A1(n5824), .A2(n7676), .ZN(n5827) );
  NAND2_X1 U7455 ( .A1(n8597), .A2(n5857), .ZN(n7873) );
  INV_X1 U7456 ( .A(n7873), .ZN(n5826) );
  NAND2_X1 U7457 ( .A1(n7780), .A2(n8299), .ZN(n7871) );
  AND2_X1 U7458 ( .A1(n6164), .A2(n7871), .ZN(n7669) );
  NAND2_X1 U7459 ( .A1(n5854), .A2(n5853), .ZN(n7506) );
  NOR2_X1 U7460 ( .A1(n7669), .A2(n7506), .ZN(n5825) );
  NAND2_X1 U7461 ( .A1(n5858), .A2(n7892), .ZN(n8604) );
  INV_X1 U7462 ( .A(n8560), .ZN(n5830) );
  NOR4_X1 U7463 ( .A1(n8029), .A2(n8509), .A3(n5832), .A4(n5831), .ZN(n5833)
         );
  NAND4_X1 U7464 ( .A1(n5834), .A2(n8504), .A3(n5833), .A4(n8481), .ZN(n5835)
         );
  NOR4_X1 U7465 ( .A1(n8430), .A2(n8447), .A3(n8465), .A4(n5835), .ZN(n5836)
         );
  XNOR2_X1 U7466 ( .A(n8722), .B(n8448), .ZN(n8438) );
  NAND3_X1 U7467 ( .A1(n5836), .A2(n8420), .A3(n8438), .ZN(n5837) );
  NOR2_X1 U7468 ( .A1(n7690), .A2(n7503), .ZN(n5909) );
  XNOR2_X1 U7469 ( .A(n5912), .B(n9055), .ZN(n6860) );
  NOR2_X1 U7470 ( .A1(n6860), .A2(P2_U3151), .ZN(n7783) );
  NOR2_X1 U7471 ( .A1(n5089), .A2(n5841), .ZN(n5842) );
  INV_X1 U7472 ( .A(n7690), .ZN(n6199) );
  NAND2_X1 U7473 ( .A1(n6199), .A2(n7503), .ZN(n5905) );
  NOR2_X1 U7474 ( .A1(n7787), .A2(n5905), .ZN(n5907) );
  INV_X1 U7475 ( .A(n8627), .ZN(n8709) );
  INV_X1 U7476 ( .A(n7415), .ZN(n5844) );
  NAND2_X1 U7477 ( .A1(n5845), .A2(n5844), .ZN(n7414) );
  NAND2_X1 U7478 ( .A1(n7414), .A2(n5846), .ZN(n8688) );
  NAND2_X1 U7479 ( .A1(n7427), .A2(n5848), .ZN(n5850) );
  NAND2_X1 U7480 ( .A1(n7674), .A2(n5852), .ZN(n7505) );
  NAND2_X1 U7481 ( .A1(n7892), .A2(n5857), .ZN(n5862) );
  NAND2_X1 U7482 ( .A1(n5858), .A2(n8597), .ZN(n5859) );
  NAND2_X1 U7483 ( .A1(n5859), .A2(n7892), .ZN(n5860) );
  AND2_X1 U7484 ( .A1(n5860), .A2(n7893), .ZN(n5861) );
  OAI21_X1 U7485 ( .B1(n7869), .B2(n5862), .A(n5861), .ZN(n5864) );
  NAND2_X1 U7486 ( .A1(n5864), .A2(n5863), .ZN(n8592) );
  INV_X1 U7487 ( .A(n8592), .ZN(n5866) );
  INV_X1 U7488 ( .A(n8591), .ZN(n5865) );
  NAND2_X1 U7489 ( .A1(n5866), .A2(n5865), .ZN(n8590) );
  NAND2_X1 U7490 ( .A1(n8590), .A2(n5867), .ZN(n7947) );
  NAND2_X1 U7491 ( .A1(n8533), .A2(n5877), .ZN(n8523) );
  NAND2_X1 U7492 ( .A1(n8523), .A2(n5878), .ZN(n5879) );
  INV_X1 U7493 ( .A(n5880), .ZN(n5882) );
  INV_X1 U7494 ( .A(n5883), .ZN(n8500) );
  NAND2_X1 U7495 ( .A1(n5890), .A2(n5889), .ZN(n8445) );
  NAND2_X1 U7496 ( .A1(n8445), .A2(n5891), .ZN(n5893) );
  NAND2_X1 U7497 ( .A1(n5893), .A2(n5892), .ZN(n8437) );
  NAND2_X1 U7498 ( .A1(n8722), .A2(n6843), .ZN(n5894) );
  OR2_X1 U7499 ( .A1(n8722), .A2(n6843), .ZN(n5895) );
  NOR2_X1 U7500 ( .A1(n8711), .A2(n8090), .ZN(n5897) );
  INV_X1 U7501 ( .A(n5898), .ZN(n5899) );
  OAI211_X1 U7502 ( .C1(n8709), .C2(n8703), .A(n5900), .B(n5899), .ZN(n5904)
         );
  INV_X1 U7503 ( .A(n8413), .ZN(n7960) );
  NAND2_X1 U7504 ( .A1(n5901), .A2(n7960), .ZN(n5902) );
  NAND2_X1 U7505 ( .A1(n5902), .A2(n8703), .ZN(n5903) );
  INV_X1 U7506 ( .A(n5908), .ZN(n5910) );
  NAND3_X1 U7507 ( .A1(n5910), .A2(n6200), .A3(n5909), .ZN(n5911) );
  INV_X1 U7508 ( .A(n6225), .ZN(n6755) );
  INV_X1 U7509 ( .A(n6216), .ZN(n5925) );
  NAND2_X1 U7510 ( .A1(n5920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5921) );
  MUX2_X1 U7511 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5921), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5922) );
  AND2_X1 U7512 ( .A1(n5923), .A2(n5922), .ZN(n6217) );
  NOR2_X1 U7513 ( .A1(n6214), .A2(n7971), .ZN(n5924) );
  NAND2_X1 U7514 ( .A1(n5925), .A2(n5924), .ZN(n6861) );
  INV_X1 U7515 ( .A(n6872), .ZN(n6868) );
  NAND3_X1 U7516 ( .A1(n6868), .A2(n6204), .A3(n4383), .ZN(n5926) );
  OAI211_X1 U7517 ( .C1(n6201), .C2(n5841), .A(n5926), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5927) );
  NAND2_X1 U7518 ( .A1(n6086), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7519 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5933) );
  MUX2_X1 U7520 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5933), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5935) );
  INV_X1 U7521 ( .A(n5943), .ZN(n5934) );
  INV_X1 U7522 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5939) );
  OAI21_X1 U7523 ( .B1(n7132), .B2(n5940), .A(n5939), .ZN(n5942) );
  AND2_X1 U7524 ( .A1(n5942), .A2(n5941), .ZN(n10285) );
  MUX2_X1 U7525 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10285), .S(n7173), .Z(n10137)
         );
  INV_X1 U7526 ( .A(n10137), .ZN(n7277) );
  OR2_X1 U7527 ( .A1(n5943), .A2(n10278), .ZN(n5944) );
  XNOR2_X1 U7528 ( .A(n5944), .B(n9088), .ZN(n7230) );
  OR2_X1 U7529 ( .A1(n7173), .A2(n7230), .ZN(n5946) );
  OR2_X1 U7530 ( .A1(n6067), .A2(n7158), .ZN(n5953) );
  OR2_X1 U7531 ( .A1(n4385), .A2(n9094), .ZN(n5952) );
  NAND2_X1 U7532 ( .A1(n5949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5948) );
  MUX2_X1 U7533 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5948), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n5950) );
  OR2_X1 U7534 ( .A1(n5949), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7535 ( .A1(n5950), .A2(n5959), .ZN(n7232) );
  OR2_X1 U7536 ( .A1(n7173), .A2(n7232), .ZN(n5951) );
  AND3_X2 U7537 ( .A1(n5953), .A2(n5952), .A3(n5951), .ZN(n10385) );
  NAND2_X1 U7538 ( .A1(n5959), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U7539 ( .A(n5954), .B(n5960), .ZN(n9599) );
  OR2_X1 U7540 ( .A1(n6067), .A2(n7151), .ZN(n5956) );
  INV_X1 U7541 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7129) );
  OR2_X1 U7542 ( .A1(n4385), .A2(n7129), .ZN(n5955) );
  INV_X2 U7543 ( .A(n9216), .ZN(n5957) );
  INV_X1 U7544 ( .A(n5959), .ZN(n5961) );
  NAND2_X1 U7545 ( .A1(n5961), .A2(n5960), .ZN(n5963) );
  NAND2_X1 U7546 ( .A1(n5963), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5962) );
  MUX2_X1 U7547 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5962), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5966) );
  INV_X1 U7548 ( .A(n5963), .ZN(n5965) );
  INV_X1 U7549 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7550 ( .A1(n5965), .A2(n5964), .ZN(n5973) );
  NAND2_X1 U7551 ( .A1(n5966), .A2(n5973), .ZN(n9614) );
  OR2_X1 U7552 ( .A1(n6067), .A2(n7153), .ZN(n5968) );
  OR2_X1 U7553 ( .A1(n4385), .A2(n7130), .ZN(n5967) );
  NAND2_X1 U7554 ( .A1(n5973), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5970) );
  XNOR2_X1 U7555 ( .A(n5970), .B(n5969), .ZN(n9628) );
  NAND2_X1 U7556 ( .A1(n7142), .A2(n5983), .ZN(n5972) );
  INV_X1 U7557 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7143) );
  OR2_X1 U7558 ( .A1(n4385), .A2(n7143), .ZN(n5971) );
  OAI211_X1 U7559 ( .C1(n7173), .C2(n9628), .A(n5972), .B(n5971), .ZN(n6319)
         );
  OAI21_X1 U7560 ( .B1(n5973), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5975) );
  INV_X1 U7561 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5974) );
  XNOR2_X1 U7562 ( .A(n5975), .B(n5974), .ZN(n9642) );
  NAND2_X1 U7563 ( .A1(n5983), .A2(n7134), .ZN(n5977) );
  INV_X1 U7564 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7135) );
  OR2_X1 U7565 ( .A1(n4384), .A2(n7135), .ZN(n5976) );
  OAI211_X1 U7566 ( .C1(n7173), .C2(n9642), .A(n5977), .B(n5976), .ZN(n10343)
         );
  OR2_X1 U7567 ( .A1(n5978), .A2(n10278), .ZN(n5980) );
  MUX2_X1 U7568 ( .A(n5980), .B(P1_IR_REG_31__SCAN_IN), .S(n5979), .Z(n5982)
         );
  NAND2_X1 U7569 ( .A1(n5982), .A2(n5981), .ZN(n7241) );
  NAND2_X1 U7570 ( .A1(n7139), .A2(n5983), .ZN(n5985) );
  OR2_X1 U7571 ( .A1(n4384), .A2(n7170), .ZN(n5984) );
  OAI211_X1 U7572 ( .C1(n7173), .C2(n7241), .A(n5985), .B(n5984), .ZN(n10064)
         );
  NAND2_X1 U7573 ( .A1(n7144), .A2(n5983), .ZN(n5989) );
  NAND2_X1 U7574 ( .A1(n5981), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5987) );
  XNOR2_X1 U7575 ( .A(n5987), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7259) );
  AOI22_X1 U7576 ( .A1(n6047), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6046), .B2(
        n7259), .ZN(n5988) );
  NAND2_X1 U7577 ( .A1(n7161), .A2(n5983), .ZN(n5991) );
  OR2_X1 U7578 ( .A1(n5981), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7579 ( .A1(n6000), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U7580 ( .A(n5992), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7313) );
  AOI22_X1 U7581 ( .A1(n6047), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6046), .B2(
        n7313), .ZN(n5990) );
  NAND2_X1 U7582 ( .A1(n5991), .A2(n5990), .ZN(n10023) );
  INV_X1 U7583 ( .A(n10023), .ZN(n10423) );
  NAND2_X1 U7584 ( .A1(n7165), .A2(n5983), .ZN(n5996) );
  NAND2_X1 U7585 ( .A1(n5992), .A2(n5997), .ZN(n5993) );
  NAND2_X1 U7586 ( .A1(n5993), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5994) );
  XNOR2_X1 U7587 ( .A(n5994), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9678) );
  AOI22_X1 U7588 ( .A1(n6047), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6046), .B2(
        n9678), .ZN(n5995) );
  NAND2_X1 U7589 ( .A1(n7185), .A2(n5983), .ZN(n6007) );
  NAND2_X1 U7590 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  NAND2_X1 U7591 ( .A1(n6003), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6002) );
  MUX2_X1 U7592 ( .A(n6002), .B(P1_IR_REG_31__SCAN_IN), .S(n6001), .Z(n6005)
         );
  INV_X1 U7593 ( .A(n6012), .ZN(n6004) );
  NAND2_X1 U7594 ( .A1(n6005), .A2(n6004), .ZN(n7597) );
  INV_X1 U7595 ( .A(n7597), .ZN(n7323) );
  AOI22_X1 U7596 ( .A1(n6047), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6046), .B2(
        n7323), .ZN(n6006) );
  NAND2_X1 U7597 ( .A1(n7199), .A2(n5983), .ZN(n6010) );
  OR2_X1 U7598 ( .A1(n6012), .A2(n10278), .ZN(n6008) );
  XNOR2_X1 U7599 ( .A(n6008), .B(P1_IR_REG_13__SCAN_IN), .ZN(n8057) );
  AOI22_X1 U7600 ( .A1(n6047), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6046), .B2(
        n8057), .ZN(n6009) );
  NAND2_X2 U7601 ( .A1(n6010), .A2(n6009), .ZN(n10222) );
  NAND2_X1 U7602 ( .A1(n7204), .A2(n5983), .ZN(n6015) );
  NAND2_X1 U7603 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  NAND2_X1 U7604 ( .A1(n6013), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6018) );
  XNOR2_X1 U7605 ( .A(n6018), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U7606 ( .A1(n6047), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6046), .B2(
        n10293), .ZN(n6014) );
  NAND2_X2 U7607 ( .A1(n6015), .A2(n6014), .ZN(n9955) );
  NAND2_X1 U7608 ( .A1(n9951), .A2(n10213), .ZN(n6016) );
  NAND2_X1 U7609 ( .A1(n7209), .A2(n5983), .ZN(n6022) );
  NAND2_X1 U7610 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  NAND2_X1 U7611 ( .A1(n6019), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6020) );
  XNOR2_X1 U7612 ( .A(n6020), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U7613 ( .A1(n6047), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6046), .B2(
        n10311), .ZN(n6021) );
  INV_X1 U7614 ( .A(n10208), .ZN(n9935) );
  NAND2_X1 U7615 ( .A1(n7299), .A2(n5983), .ZN(n6025) );
  CLKBUF_X3 U7616 ( .A(n6023), .Z(n6080) );
  XNOR2_X1 U7617 ( .A(n6030), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8066) );
  AOI22_X1 U7618 ( .A1(n6047), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6046), .B2(
        n8066), .ZN(n6024) );
  NAND2_X1 U7619 ( .A1(n7270), .A2(n5983), .ZN(n6028) );
  XNOR2_X1 U7620 ( .A(n6026), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8064) );
  AOI22_X1 U7621 ( .A1(n6047), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6046), .B2(
        n8064), .ZN(n6027) );
  OR2_X1 U7622 ( .A1(n10197), .A2(n10271), .ZN(n6029) );
  NOR2_X2 U7623 ( .A1(n9895), .A2(n6029), .ZN(n9878) );
  NAND2_X1 U7624 ( .A1(n7366), .A2(n5983), .ZN(n6036) );
  INV_X1 U7625 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U7626 ( .A1(n6030), .A2(n8905), .ZN(n6042) );
  NAND2_X1 U7627 ( .A1(n6042), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6032) );
  OR2_X1 U7628 ( .A1(n6032), .A2(n6031), .ZN(n6034) );
  NAND2_X1 U7629 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  AOI22_X1 U7630 ( .A1(n6047), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6046), .B2(
        n8068), .ZN(n6035) );
  NAND2_X1 U7631 ( .A1(n7501), .A2(n5983), .ZN(n6049) );
  INV_X1 U7632 ( .A(n6042), .ZN(n6037) );
  NAND2_X1 U7633 ( .A1(n6037), .A2(n6078), .ZN(n6045) );
  NAND2_X1 U7634 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n6038) );
  NAND2_X1 U7635 ( .A1(n6038), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6039) );
  OAI21_X1 U7636 ( .B1(n6040), .B2(P1_IR_REG_31__SCAN_IN), .A(n6039), .ZN(
        n6044) );
  AND2_X1 U7637 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6041) );
  NAND2_X1 U7638 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  NAND3_X2 U7639 ( .A1(n6045), .A2(n6044), .A3(n6043), .ZN(n9551) );
  AOI22_X1 U7640 ( .A1(n6047), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6046), .B2(
        n9540), .ZN(n6048) );
  NAND2_X1 U7641 ( .A1(n7689), .A2(n5983), .ZN(n6051) );
  OR2_X1 U7642 ( .A1(n4384), .A2(n7707), .ZN(n6050) );
  OR2_X1 U7643 ( .A1(n4385), .A2(n7793), .ZN(n6052) );
  NAND2_X1 U7644 ( .A1(n7729), .A2(n5983), .ZN(n6054) );
  OR2_X1 U7645 ( .A1(n4385), .A2(n7734), .ZN(n6053) );
  NAND2_X1 U7646 ( .A1(n7790), .A2(n5983), .ZN(n6056) );
  OR2_X1 U7647 ( .A1(n4384), .A2(n9062), .ZN(n6055) );
  NAND2_X1 U7648 ( .A1(n7900), .A2(n5983), .ZN(n6058) );
  OR2_X1 U7649 ( .A1(n4385), .A2(n9037), .ZN(n6057) );
  NAND2_X1 U7650 ( .A1(n7959), .A2(n5983), .ZN(n6060) );
  OR2_X1 U7651 ( .A1(n4384), .A2(n9063), .ZN(n6059) );
  NAND2_X1 U7652 ( .A1(n7970), .A2(n5983), .ZN(n6062) );
  OR2_X1 U7653 ( .A1(n4384), .A2(n7973), .ZN(n6061) );
  NAND2_X1 U7654 ( .A1(n7976), .A2(n5983), .ZN(n6064) );
  OR2_X1 U7655 ( .A1(n4385), .A2(n7990), .ZN(n6063) );
  NAND2_X2 U7656 ( .A1(n6064), .A2(n6063), .ZN(n8821) );
  NAND2_X1 U7657 ( .A1(n6521), .A2(n9721), .ZN(n6522) );
  NAND2_X1 U7658 ( .A1(n8103), .A2(n5983), .ZN(n6066) );
  OR2_X1 U7659 ( .A1(n4385), .A2(n8104), .ZN(n6065) );
  INV_X1 U7660 ( .A(n8806), .ZN(n6068) );
  INV_X1 U7661 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8005) );
  OR2_X1 U7662 ( .A1(n4384), .A2(n8005), .ZN(n6069) );
  NAND2_X1 U7663 ( .A1(n8006), .A2(n5983), .ZN(n6072) );
  OR2_X1 U7664 ( .A1(n4385), .A2(n8008), .ZN(n6071) );
  NAND2_X1 U7665 ( .A1(n9712), .A2(n10236), .ZN(n9711) );
  NAND2_X1 U7666 ( .A1(n8797), .A2(n5983), .ZN(n6076) );
  INV_X1 U7667 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6073) );
  OR2_X1 U7668 ( .A1(n4384), .A2(n6073), .ZN(n6075) );
  NOR2_X1 U7669 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6077) );
  NAND2_X1 U7670 ( .A1(n6023), .A2(n6079), .ZN(n6103) );
  NAND2_X1 U7671 ( .A1(n6082), .A2(n6104), .ZN(n6081) );
  INV_X2 U7672 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7673 ( .A1(n6103), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7674 ( .A1(n6084), .A2(n10369), .ZN(n9710) );
  NAND2_X1 U7675 ( .A1(n6088), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7676 ( .A1(n6533), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7677 ( .A1(n6403), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7678 ( .A1(n6541), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6092) );
  NAND3_X1 U7679 ( .A1(n6094), .A2(n6093), .A3(n6092), .ZN(n9562) );
  INV_X1 U7680 ( .A(P1_B_REG_SCAN_IN), .ZN(n6097) );
  OR2_X1 U7681 ( .A1(n7989), .A2(n6097), .ZN(n6098) );
  NAND2_X1 U7682 ( .A1(n10017), .A2(n6098), .ZN(n6545) );
  INV_X1 U7683 ( .A(n6545), .ZN(n6099) );
  NAND2_X1 U7684 ( .A1(n9562), .A2(n6099), .ZN(n10142) );
  NAND2_X1 U7685 ( .A1(n6100), .A2(n6105), .ZN(n6101) );
  NAND2_X1 U7686 ( .A1(n6101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6102) );
  INV_X1 U7687 ( .A(n6103), .ZN(n6106) );
  INV_X1 U7688 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6107) );
  INV_X1 U7689 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6109) );
  INV_X1 U7690 ( .A(n6125), .ZN(n6121) );
  NAND2_X1 U7691 ( .A1(n6111), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7692 ( .A1(n6115), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6116) );
  MUX2_X1 U7693 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6116), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6119) );
  INV_X1 U7694 ( .A(n6117), .ZN(n6118) );
  AND2_X1 U7695 ( .A1(n6119), .A2(n6118), .ZN(n6123) );
  INV_X1 U7696 ( .A(n6523), .ZN(n6128) );
  OAI21_X1 U7697 ( .B1(n6122), .B2(P1_B_REG_SCAN_IN), .A(n6123), .ZN(n6124) );
  INV_X1 U7698 ( .A(n6124), .ZN(n6127) );
  NAND3_X1 U7699 ( .A1(n6125), .A2(P1_B_REG_SCAN_IN), .A3(n6122), .ZN(n6126)
         );
  NAND2_X1 U7700 ( .A1(n6122), .A2(n7975), .ZN(n10277) );
  OAI21_X1 U7701 ( .B1(n6129), .B2(P1_D_REG_0__SCAN_IN), .A(n10277), .ZN(n7082) );
  NAND2_X1 U7702 ( .A1(n6125), .A2(n7975), .ZN(n7191) );
  OAI21_X1 U7703 ( .B1(n6129), .B2(P1_D_REG_1__SCAN_IN), .A(n7191), .ZN(n7080)
         );
  NAND2_X1 U7704 ( .A1(n10369), .A2(n9540), .ZN(n7088) );
  NOR2_X1 U7705 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .ZN(
        n9105) );
  NOR4_X1 U7706 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6132) );
  NOR4_X1 U7707 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6131) );
  NOR4_X1 U7708 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6130) );
  AND4_X1 U7709 ( .A1(n9105), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n6138)
         );
  NOR4_X1 U7710 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6136) );
  NOR4_X1 U7711 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6135) );
  NOR4_X1 U7712 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6134) );
  NOR4_X1 U7713 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6133) );
  AND4_X1 U7714 ( .A1(n6136), .A2(n6135), .A3(n6134), .A4(n6133), .ZN(n6137)
         );
  NAND2_X1 U7715 ( .A1(n6138), .A2(n6137), .ZN(n6139) );
  NAND2_X1 U7716 ( .A1(n7189), .A2(n6139), .ZN(n7079) );
  NAND2_X1 U7717 ( .A1(n6141), .A2(n6140), .ZN(n6143) );
  INV_X1 U7718 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U7719 ( .A1(n6146), .A2(n6145), .ZN(n6197) );
  NAND2_X1 U7720 ( .A1(n6754), .A2(n7690), .ZN(n6756) );
  NAND2_X1 U7721 ( .A1(n6756), .A2(n7730), .ZN(n6148) );
  NAND2_X1 U7722 ( .A1(n6148), .A2(n7503), .ZN(n6212) );
  INV_X1 U7723 ( .A(n6212), .ZN(n6149) );
  NAND2_X1 U7724 ( .A1(n6149), .A2(n7462), .ZN(n7878) );
  NAND2_X1 U7725 ( .A1(n6150), .A2(n7475), .ZN(n6151) );
  NAND2_X1 U7726 ( .A1(n6152), .A2(n6151), .ZN(n8690) );
  NAND2_X1 U7727 ( .A1(n8690), .A2(n8691), .ZN(n6154) );
  NAND2_X1 U7728 ( .A1(n7336), .A2(n7328), .ZN(n6153) );
  NAND2_X1 U7729 ( .A1(n6154), .A2(n6153), .ZN(n7428) );
  NAND2_X1 U7730 ( .A1(n7428), .A2(n7429), .ZN(n6156) );
  NAND2_X1 U7731 ( .A1(n7329), .A2(n7344), .ZN(n6155) );
  NAND2_X1 U7732 ( .A1(n6156), .A2(n6155), .ZN(n7541) );
  NAND2_X1 U7733 ( .A1(n7541), .A2(n7542), .ZN(n7680) );
  NAND2_X1 U7734 ( .A1(n7348), .A2(n6776), .ZN(n7679) );
  OR2_X1 U7735 ( .A1(n8302), .A2(n7440), .ZN(n6157) );
  AND2_X1 U7736 ( .A1(n7679), .A2(n6157), .ZN(n6158) );
  NAND2_X1 U7737 ( .A1(n7680), .A2(n6158), .ZN(n6160) );
  NAND2_X1 U7738 ( .A1(n8302), .A2(n7440), .ZN(n6159) );
  NAND2_X1 U7739 ( .A1(n6160), .A2(n6159), .ZN(n7507) );
  INV_X1 U7740 ( .A(n7700), .ZN(n8301) );
  NAND2_X1 U7741 ( .A1(n7512), .A2(n8301), .ZN(n6161) );
  NAND2_X1 U7742 ( .A1(n7814), .A2(n6163), .ZN(n7665) );
  AND2_X1 U7743 ( .A1(n7665), .A2(n6164), .ZN(n6165) );
  NAND2_X1 U7744 ( .A1(n7664), .A2(n6165), .ZN(n7872) );
  AND2_X1 U7745 ( .A1(n7873), .A2(n7871), .ZN(n6166) );
  OR2_X1 U7746 ( .A1(n7868), .A2(n8608), .ZN(n6167) );
  OR2_X1 U7747 ( .A1(n8677), .A2(n8297), .ZN(n7940) );
  OR2_X1 U7748 ( .A1(n8579), .A2(n8607), .ZN(n7938) );
  NAND2_X1 U7749 ( .A1(n7940), .A2(n7938), .ZN(n6174) );
  NAND2_X1 U7750 ( .A1(n8677), .A2(n8297), .ZN(n6172) );
  NAND2_X1 U7751 ( .A1(n8602), .A2(n8298), .ZN(n7887) );
  NAND2_X1 U7752 ( .A1(n7887), .A2(n8157), .ZN(n6170) );
  INV_X1 U7753 ( .A(n7887), .ZN(n6169) );
  AOI22_X1 U7754 ( .A1(n8579), .A2(n6170), .B1(n6169), .B2(n8607), .ZN(n6171)
         );
  NAND2_X1 U7755 ( .A1(n6172), .A2(n6171), .ZN(n7941) );
  AOI22_X1 U7756 ( .A1(n8583), .A2(n8227), .B1(n7941), .B2(n7940), .ZN(n6173)
         );
  OR2_X1 U7757 ( .A1(n8227), .A2(n8583), .ZN(n6175) );
  INV_X1 U7758 ( .A(n8569), .ZN(n6177) );
  NAND2_X1 U7759 ( .A1(n8785), .A2(n8296), .ZN(n6178) );
  INV_X1 U7760 ( .A(n8772), .ZN(n8182) );
  NAND2_X1 U7761 ( .A1(n8535), .A2(n6182), .ZN(n6184) );
  NAND2_X1 U7762 ( .A1(n8767), .A2(n8547), .ZN(n6183) );
  NAND2_X1 U7763 ( .A1(n6184), .A2(n6183), .ZN(n8525) );
  INV_X1 U7764 ( .A(n8525), .ZN(n6185) );
  OR2_X1 U7765 ( .A1(n8761), .A2(n8536), .ZN(n6186) );
  NAND2_X1 U7766 ( .A1(n8755), .A2(n8527), .ZN(n8032) );
  NOR2_X1 U7767 ( .A1(n8216), .A2(n8515), .ZN(n8491) );
  INV_X1 U7768 ( .A(n8499), .ZN(n8749) );
  AOI22_X1 U7769 ( .A1(n8493), .A2(n8491), .B1(n8483), .B2(n8749), .ZN(n6188)
         );
  OR2_X1 U7770 ( .A1(n8230), .A2(n8473), .ZN(n6190) );
  NOR2_X1 U7771 ( .A1(n8740), .A2(n8457), .ZN(n6191) );
  INV_X1 U7772 ( .A(n8740), .ZN(n8123) );
  AND2_X1 U7773 ( .A1(n8734), .A2(n8474), .ZN(n6193) );
  OR2_X1 U7774 ( .A1(n8734), .A2(n8474), .ZN(n6192) );
  NAND2_X1 U7775 ( .A1(n8728), .A2(n8458), .ZN(n6194) );
  AND2_X1 U7776 ( .A1(n8722), .A2(n8448), .ZN(n6195) );
  NAND2_X1 U7777 ( .A1(n8092), .A2(n8090), .ZN(n6196) );
  XNOR2_X1 U7778 ( .A(n6198), .B(n6197), .ZN(n6210) );
  NAND2_X1 U7779 ( .A1(n6200), .A2(n6199), .ZN(n6202) );
  NAND2_X1 U7780 ( .A1(n6587), .A2(n6201), .ZN(n6742) );
  NAND2_X1 U7781 ( .A1(n6204), .A2(n6203), .ZN(n6205) );
  NAND2_X1 U7782 ( .A1(n6207), .A2(n6205), .ZN(n6871) );
  NAND2_X1 U7783 ( .A1(n6207), .A2(P2_B_REG_SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7784 ( .A1(n8692), .A2(n6208), .ZN(n8412) );
  OAI22_X1 U7785 ( .A1(n8090), .A2(n8694), .B1(n7850), .B2(n8412), .ZN(n6209)
         );
  AOI21_X1 U7786 ( .B1(n6210), .B2(n8696), .A(n6209), .ZN(n6211) );
  OR2_X1 U7787 ( .A1(n6212), .A2(n7690), .ZN(n6213) );
  NAND2_X1 U7788 ( .A1(n6213), .A2(n6846), .ZN(n6222) );
  NAND2_X1 U7789 ( .A1(n6216), .A2(n6215), .ZN(n6218) );
  NAND2_X1 U7790 ( .A1(n6214), .A2(n7971), .ZN(n7194) );
  OAI21_X2 U7791 ( .B1(n6219), .B2(P2_D_REG_0__SCAN_IN), .A(n7194), .ZN(n6759)
         );
  NAND2_X1 U7792 ( .A1(n6216), .A2(n7971), .ZN(n6220) );
  NAND2_X1 U7793 ( .A1(n6222), .A2(n8796), .ZN(n6223) );
  NAND2_X1 U7794 ( .A1(n6224), .A2(n6223), .ZN(n7122) );
  INV_X1 U7795 ( .A(n6759), .ZN(n6740) );
  OR2_X1 U7796 ( .A1(n6846), .A2(n6225), .ZN(n6859) );
  NOR4_X1 U7797 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6233) );
  INV_X1 U7798 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n8968) );
  INV_X1 U7799 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n8967) );
  INV_X1 U7800 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n8915) );
  INV_X1 U7801 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9026) );
  NAND4_X1 U7802 ( .A1(n8968), .A2(n8967), .A3(n8915), .A4(n9026), .ZN(n9067)
         );
  NOR4_X1 U7803 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6229) );
  NOR4_X1 U7804 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6228) );
  NOR4_X1 U7805 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6227) );
  NOR4_X1 U7806 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6226) );
  NAND4_X1 U7807 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .ZN(n6230)
         );
  NOR4_X1 U7808 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        n9067), .A4(n6230), .ZN(n6232) );
  NOR4_X1 U7809 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6231) );
  AND3_X1 U7810 ( .A1(n6233), .A2(n6232), .A3(n6231), .ZN(n6234) );
  AND3_X1 U7811 ( .A1(n6859), .A2(n7160), .A3(n6745), .ZN(n7120) );
  OAI21_X1 U7812 ( .B1(n6740), .B2(n8796), .A(n7120), .ZN(n6235) );
  NOR2_X1 U7813 ( .A1(n6756), .A2(n7503), .ZN(n10463) );
  NAND2_X1 U7814 ( .A1(n10464), .A2(n10463), .ZN(n7673) );
  NOR2_X1 U7815 ( .A1(n6237), .A2(n10458), .ZN(n8414) );
  INV_X1 U7816 ( .A(n6238), .ZN(n6239) );
  INV_X1 U7817 ( .A(n8567), .ZN(n8461) );
  NOR2_X1 U7818 ( .A1(n7127), .A2(n8618), .ZN(n6240) );
  AOI211_X1 U7819 ( .C1(n10466), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8414), .B(
        n6240), .ZN(n6241) );
  NAND2_X1 U7820 ( .A1(n6244), .A2(n6243), .ZN(P2_U3204) );
  NAND2_X1 U7821 ( .A1(n4381), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6252) );
  INV_X1 U7822 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9138) );
  AND2_X2 U7823 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6285) );
  NOR2_X2 U7824 ( .A1(n6305), .A2(n6304), .ZN(n6307) );
  NAND2_X1 U7825 ( .A1(n6307), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6297) );
  NOR2_X2 U7826 ( .A1(n6312), .A2(n7225), .ZN(n6322) );
  AND2_X2 U7827 ( .A1(n6322), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6328) );
  INV_X1 U7828 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6347) );
  INV_X1 U7829 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8896) );
  OR2_X2 U7830 ( .A1(n6363), .A2(n8896), .ZN(n6368) );
  INV_X1 U7831 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6367) );
  NOR2_X2 U7832 ( .A1(n6368), .A2(n6367), .ZN(n6372) );
  AND2_X2 U7833 ( .A1(n6372), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6378) );
  INV_X1 U7834 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6393) );
  INV_X1 U7835 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8875) );
  INV_X1 U7836 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U7837 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n6431), .ZN(n6443) );
  INV_X1 U7838 ( .A(n6443), .ZN(n6247) );
  NAND2_X1 U7839 ( .A1(n6247), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6454) );
  INV_X1 U7840 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U7841 ( .A1(n8935), .A2(n6443), .ZN(n6248) );
  NAND2_X1 U7842 ( .A1(n4388), .A2(n9719), .ZN(n6251) );
  NAND2_X1 U7843 ( .A1(n6403), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7844 ( .A1(n6404), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6249) );
  OR2_X1 U7845 ( .A1(n8821), .A2(n7104), .ZN(n9407) );
  NAND2_X1 U7846 ( .A1(n8821), .A2(n7104), .ZN(n9411) );
  NAND2_X1 U7847 ( .A1(n4388), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6257) );
  INV_X1 U7848 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7849 ( .A1(n4378), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7850 ( .A1(n6423), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6254) );
  NAND4_X2 U7851 ( .A1(n6257), .A2(n6256), .A3(n6255), .A4(n6254), .ZN(n9571)
         );
  NAND2_X1 U7852 ( .A1(n10108), .A2(n7518), .ZN(n6273) );
  NOR2_X1 U7853 ( .A1(n5070), .A2(n5071), .ZN(n6262) );
  INV_X1 U7854 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6258) );
  OR2_X1 U7855 ( .A1(n6259), .A2(n6258), .ZN(n6261) );
  NAND2_X1 U7856 ( .A1(n6274), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6260) );
  AND3_X2 U7857 ( .A1(n6262), .A2(n6261), .A3(n6260), .ZN(n7361) );
  NAND2_X1 U7858 ( .A1(n7361), .A2(n10137), .ZN(n7479) );
  NAND2_X1 U7859 ( .A1(n4378), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7860 ( .A1(n6263), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6268) );
  INV_X1 U7861 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6264) );
  OR2_X1 U7862 ( .A1(n6265), .A2(n6264), .ZN(n6267) );
  NAND2_X1 U7863 ( .A1(n6374), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6266) );
  AND4_X4 U7864 ( .A1(n6269), .A2(n6268), .A3(n6267), .A4(n6266), .ZN(n9480)
         );
  NAND2_X1 U7865 ( .A1(n7479), .A2(n9572), .ZN(n6270) );
  NAND3_X1 U7866 ( .A1(n6271), .A2(n9482), .A3(n6270), .ZN(n6272) );
  INV_X1 U7867 ( .A(n10106), .ZN(n6279) );
  NAND2_X1 U7868 ( .A1(n6533), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6278) );
  INV_X1 U7869 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U7870 ( .A1(n6413), .A2(n7533), .ZN(n6277) );
  NAND2_X1 U7871 ( .A1(n4378), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7872 ( .A1(n6541), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6275) );
  INV_X2 U7873 ( .A(n9570), .ZN(n9214) );
  INV_X1 U7874 ( .A(n10385), .ZN(n10104) );
  NAND2_X1 U7875 ( .A1(n6279), .A2(n9322), .ZN(n9488) );
  NAND2_X1 U7876 ( .A1(n9570), .A2(n10385), .ZN(n9485) );
  NOR2_X1 U7877 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6280) );
  NOR2_X1 U7878 ( .A1(n6285), .A2(n6280), .ZN(n10087) );
  NAND2_X1 U7879 ( .A1(n4389), .A2(n10087), .ZN(n6283) );
  NAND2_X1 U7880 ( .A1(n4378), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7881 ( .A1(n6404), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7882 ( .A1(n4381), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6290) );
  OAI21_X1 U7883 ( .B1(n6285), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6305), .ZN(
        n6286) );
  INV_X1 U7884 ( .A(n6286), .ZN(n10357) );
  NAND2_X1 U7885 ( .A1(n6413), .A2(n10357), .ZN(n6289) );
  NAND2_X1 U7886 ( .A1(n4378), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7887 ( .A1(n6541), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6287) );
  AND4_X2 U7888 ( .A1(n6290), .A2(n6289), .A3(n6288), .A4(n6287), .ZN(n10073)
         );
  NAND2_X1 U7889 ( .A1(n10073), .A2(n10360), .ZN(n9490) );
  NAND2_X2 U7890 ( .A1(n9569), .A2(n10392), .ZN(n6472) );
  NAND2_X1 U7891 ( .A1(n10352), .A2(n6472), .ZN(n10029) );
  OR2_X1 U7892 ( .A1(n6307), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6291) );
  AND2_X1 U7893 ( .A1(n6297), .A2(n6291), .ZN(n10342) );
  NAND2_X1 U7894 ( .A1(n6413), .A2(n10342), .ZN(n6295) );
  NAND2_X1 U7895 ( .A1(n4381), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7896 ( .A1(n6403), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7897 ( .A1(n6541), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U7898 ( .A1(n10072), .A2(n10343), .ZN(n10055) );
  NAND2_X1 U7899 ( .A1(n6533), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7900 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  AND2_X1 U7901 ( .A1(n6312), .A2(n6298), .ZN(n10063) );
  NAND2_X1 U7902 ( .A1(n6413), .A2(n10063), .ZN(n6301) );
  NAND2_X1 U7903 ( .A1(n6403), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7904 ( .A1(n6541), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6299) );
  AND4_X2 U7905 ( .A1(n6302), .A2(n6301), .A3(n6300), .A4(n6299), .ZN(n10334)
         );
  NAND2_X1 U7906 ( .A1(n10334), .A2(n10064), .ZN(n9344) );
  NAND2_X1 U7907 ( .A1(n10055), .A2(n9344), .ZN(n10034) );
  NAND2_X1 U7908 ( .A1(n4381), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6310) );
  AND2_X1 U7909 ( .A1(n6305), .A2(n6304), .ZN(n6306) );
  NOR2_X1 U7910 ( .A1(n6307), .A2(n6306), .ZN(n10078) );
  NAND2_X1 U7911 ( .A1(n6413), .A2(n10078), .ZN(n6309) );
  NAND2_X1 U7912 ( .A1(n6541), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6308) );
  INV_X1 U7913 ( .A(n9492), .ZN(n10030) );
  NOR2_X1 U7914 ( .A1(n10034), .A2(n10030), .ZN(n6311) );
  INV_X1 U7915 ( .A(n10050), .ZN(n10416) );
  NAND2_X1 U7916 ( .A1(n6533), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6317) );
  AND2_X1 U7917 ( .A1(n6312), .A2(n7225), .ZN(n6313) );
  NOR2_X1 U7918 ( .A1(n6322), .A2(n6313), .ZN(n10046) );
  NAND2_X1 U7919 ( .A1(n6413), .A2(n10046), .ZN(n6316) );
  NAND2_X1 U7920 ( .A1(n6403), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7921 ( .A1(n6404), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U7922 ( .A1(n6318), .A2(n10034), .ZN(n9498) );
  INV_X1 U7923 ( .A(n6319), .ZN(n10397) );
  NAND2_X1 U7924 ( .A1(n9568), .A2(n10397), .ZN(n10031) );
  NAND2_X1 U7925 ( .A1(n9567), .A2(n10403), .ZN(n9343) );
  NAND2_X1 U7926 ( .A1(n9498), .A2(n9497), .ZN(n6320) );
  NAND2_X1 U7927 ( .A1(n4381), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6327) );
  NOR2_X1 U7928 ( .A1(n6322), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U7929 ( .A1(n4389), .A2(n4392), .ZN(n6326) );
  NAND2_X1 U7930 ( .A1(n6403), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7931 ( .A1(n6404), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6324) );
  OR2_X1 U7932 ( .A1(n10023), .A2(n10043), .ZN(n9500) );
  NAND2_X1 U7933 ( .A1(n10023), .A2(n10043), .ZN(n9991) );
  NAND2_X1 U7934 ( .A1(n9500), .A2(n9991), .ZN(n10009) );
  INV_X1 U7935 ( .A(n10009), .ZN(n10013) );
  NAND2_X1 U7936 ( .A1(n4381), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6333) );
  OR2_X1 U7937 ( .A1(n6328), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6329) );
  AND2_X1 U7938 ( .A1(n6335), .A2(n6329), .ZN(n10003) );
  NAND2_X1 U7939 ( .A1(n4389), .A2(n10003), .ZN(n6332) );
  NAND2_X1 U7940 ( .A1(n6403), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7941 ( .A1(n6541), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6330) );
  NAND4_X1 U7942 ( .A1(n6333), .A2(n6332), .A3(n6331), .A4(n6330), .ZN(n10016)
         );
  INV_X1 U7943 ( .A(n10016), .ZN(n8853) );
  NAND2_X1 U7944 ( .A1(n10227), .A2(n8853), .ZN(n9349) );
  AND2_X1 U7945 ( .A1(n9349), .A2(n9991), .ZN(n9504) );
  OR2_X1 U7946 ( .A1(n10227), .A2(n8853), .ZN(n9359) );
  NAND2_X1 U7947 ( .A1(n6334), .A2(n9359), .ZN(n7996) );
  NAND2_X1 U7948 ( .A1(n6533), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7949 ( .A1(n6335), .A2(n7310), .ZN(n6336) );
  AND2_X1 U7950 ( .A1(n6341), .A2(n6336), .ZN(n9978) );
  NAND2_X1 U7951 ( .A1(n6413), .A2(n9978), .ZN(n6339) );
  NAND2_X1 U7952 ( .A1(n6403), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U7953 ( .A1(n6404), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7954 ( .A1(n7994), .A2(n9968), .ZN(n9506) );
  NAND2_X1 U7955 ( .A1(n6533), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U7956 ( .A1(n6341), .A2(n7603), .ZN(n6342) );
  AND2_X1 U7957 ( .A1(n6348), .A2(n6342), .ZN(n9971) );
  NAND2_X1 U7958 ( .A1(n4389), .A2(n9971), .ZN(n6345) );
  NAND2_X1 U7959 ( .A1(n4386), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U7960 ( .A1(n6404), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6343) );
  OR2_X1 U7961 ( .A1(n10222), .A2(n9941), .ZN(n9507) );
  NAND2_X1 U7962 ( .A1(n10222), .A2(n9941), .ZN(n9944) );
  NAND2_X1 U7963 ( .A1(n4381), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6353) );
  AND2_X1 U7964 ( .A1(n6348), .A2(n6347), .ZN(n6349) );
  NOR2_X1 U7965 ( .A1(n6356), .A2(n6349), .ZN(n9954) );
  NAND2_X1 U7966 ( .A1(n6413), .A2(n9954), .ZN(n6352) );
  NAND2_X1 U7967 ( .A1(n4386), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U7968 ( .A1(n6541), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6350) );
  NAND4_X1 U7969 ( .A1(n6353), .A2(n6352), .A3(n6351), .A4(n6350), .ZN(n9929)
         );
  INV_X1 U7970 ( .A(n9929), .ZN(n9967) );
  NAND2_X1 U7971 ( .A1(n9955), .A2(n9967), .ZN(n9354) );
  INV_X1 U7972 ( .A(n9944), .ZN(n6354) );
  NOR2_X1 U7973 ( .A1(n9947), .A2(n6354), .ZN(n6355) );
  OR2_X1 U7974 ( .A1(n6356), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6357) );
  AND2_X1 U7975 ( .A1(n6357), .A2(n6363), .ZN(n9932) );
  NAND2_X1 U7976 ( .A1(n6413), .A2(n9932), .ZN(n6361) );
  NAND2_X1 U7977 ( .A1(n4381), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U7978 ( .A1(n4386), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U7979 ( .A1(n6541), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6358) );
  OR2_X1 U7980 ( .A1(n10208), .A2(n9942), .ZN(n9513) );
  NAND2_X1 U7981 ( .A1(n10208), .A2(n9942), .ZN(n9370) );
  NAND2_X1 U7982 ( .A1(n9513), .A2(n9370), .ZN(n9924) );
  INV_X1 U7983 ( .A(n9508), .ZN(n9925) );
  NOR2_X1 U7984 ( .A1(n9924), .A2(n9925), .ZN(n6362) );
  NAND2_X1 U7985 ( .A1(n9923), .A2(n6362), .ZN(n9926) );
  NAND2_X1 U7986 ( .A1(n6363), .A2(n8896), .ZN(n6364) );
  AND2_X1 U7987 ( .A1(n6368), .A2(n6364), .ZN(n9917) );
  AOI22_X1 U7988 ( .A1(n9917), .A2(n4389), .B1(n6533), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n6366) );
  AOI22_X1 U7989 ( .A1(n4386), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n6404), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U7990 ( .A1(n10271), .A2(n9894), .ZN(n9516) );
  INV_X1 U7991 ( .A(n9516), .ZN(n9312) );
  AND2_X1 U7992 ( .A1(n6368), .A2(n6367), .ZN(n6369) );
  OR2_X1 U7993 ( .A1(n6369), .A2(n6372), .ZN(n9897) );
  AOI22_X1 U7994 ( .A1(n4381), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n4386), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U7995 ( .A1(n6541), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6370) );
  OAI211_X1 U7996 ( .C1(n9897), .C2(n6303), .A(n6371), .B(n6370), .ZN(n9914)
         );
  INV_X1 U7997 ( .A(n9914), .ZN(n9877) );
  NAND2_X1 U7998 ( .A1(n10197), .A2(n9877), .ZN(n9429) );
  NAND2_X1 U7999 ( .A1(n9891), .A2(n9429), .ZN(n9872) );
  NOR2_X1 U8000 ( .A1(n6372), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6373) );
  OR2_X1 U8001 ( .A1(n6378), .A2(n6373), .ZN(n9882) );
  AOI22_X1 U8002 ( .A1(n4381), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n4386), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U8003 ( .A1(n6541), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6375) );
  OAI211_X1 U8004 ( .C1(n9882), .C2(n6303), .A(n6376), .B(n6375), .ZN(n9860)
         );
  INV_X1 U8005 ( .A(n9860), .ZN(n9893) );
  OR2_X1 U8006 ( .A1(n9881), .A2(n9893), .ZN(n9428) );
  AND2_X1 U8007 ( .A1(n9428), .A2(n9871), .ZN(n9519) );
  NAND2_X1 U8008 ( .A1(n9872), .A2(n9519), .ZN(n6377) );
  NAND2_X1 U8009 ( .A1(n9881), .A2(n9893), .ZN(n9427) );
  NAND2_X1 U8010 ( .A1(n6377), .A2(n9427), .ZN(n9858) );
  OR2_X1 U8011 ( .A1(n6378), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6379) );
  AND2_X1 U8012 ( .A1(n6394), .A2(n6379), .ZN(n9863) );
  NAND2_X1 U8013 ( .A1(n9863), .A2(n4389), .ZN(n6385) );
  INV_X1 U8014 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U8015 ( .A1(n4386), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U8016 ( .A1(n6404), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6381) );
  OAI211_X1 U8017 ( .C1(n6436), .C2(n10187), .A(n6382), .B(n6381), .ZN(n6383)
         );
  INV_X1 U8018 ( .A(n6383), .ZN(n6384) );
  NAND2_X1 U8019 ( .A1(n6385), .A2(n6384), .ZN(n9845) );
  INV_X1 U8020 ( .A(n9845), .ZN(n9876) );
  OR2_X1 U8021 ( .A1(n9864), .A2(n9876), .ZN(n9380) );
  NAND2_X1 U8022 ( .A1(n9864), .A2(n9876), .ZN(n9520) );
  NAND2_X1 U8023 ( .A1(n9858), .A2(n9857), .ZN(n6386) );
  AND2_X1 U8024 ( .A1(n4471), .A2(n8875), .ZN(n6387) );
  OR2_X1 U8025 ( .A1(n6387), .A2(n6401), .ZN(n9833) );
  INV_X1 U8026 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U8027 ( .A1(n6533), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U8028 ( .A1(n6404), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6388) );
  OAI211_X1 U8029 ( .C1(n6390), .C2(n9145), .A(n6389), .B(n6388), .ZN(n6391)
         );
  INV_X1 U8030 ( .A(n6391), .ZN(n6392) );
  OAI21_X2 U8031 ( .B1(n9833), .B2(n6433), .A(n6392), .ZN(n9846) );
  INV_X1 U8032 ( .A(n9846), .ZN(n9237) );
  OR2_X1 U8033 ( .A1(n10256), .A2(n9237), .ZN(n6505) );
  NAND2_X1 U8034 ( .A1(n6394), .A2(n6393), .ZN(n6395) );
  AND2_X1 U8035 ( .A1(n4471), .A2(n6395), .ZN(n9850) );
  NAND2_X1 U8036 ( .A1(n9850), .A2(n6413), .ZN(n6400) );
  INV_X1 U8037 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9045) );
  NAND2_X1 U8038 ( .A1(n4381), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U8039 ( .A1(n6541), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6396) );
  OAI211_X1 U8040 ( .C1(n6390), .C2(n9045), .A(n6397), .B(n6396), .ZN(n6398)
         );
  INV_X1 U8041 ( .A(n6398), .ZN(n6399) );
  NAND2_X1 U8042 ( .A1(n6400), .A2(n6399), .ZN(n9861) );
  NAND2_X1 U8043 ( .A1(n9853), .A2(n9861), .ZN(n9820) );
  NOR2_X1 U8044 ( .A1(n6401), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6402) );
  OR2_X1 U8045 ( .A1(n6411), .A2(n6402), .ZN(n9809) );
  INV_X1 U8046 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U8047 ( .A1(n6403), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U8048 ( .A1(n6423), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6405) );
  OAI211_X1 U8049 ( .C1(n10169), .C2(n6436), .A(n6406), .B(n6405), .ZN(n6407)
         );
  INV_X1 U8050 ( .A(n6407), .ZN(n6408) );
  OAI21_X2 U8051 ( .B1(n9809), .B2(n6433), .A(n6408), .ZN(n9826) );
  INV_X1 U8052 ( .A(n9826), .ZN(n6409) );
  OR2_X1 U8053 ( .A1(n9808), .A2(n6409), .ZN(n9310) );
  NAND2_X1 U8054 ( .A1(n9808), .A2(n6409), .ZN(n9377) );
  NAND2_X1 U8055 ( .A1(n10256), .A2(n9237), .ZN(n9376) );
  INV_X1 U8056 ( .A(n9861), .ZN(n8876) );
  NAND2_X1 U8057 ( .A1(n10180), .A2(n8876), .ZN(n9821) );
  NAND2_X1 U8058 ( .A1(n9376), .A2(n9821), .ZN(n6410) );
  NAND2_X1 U8059 ( .A1(n6410), .A2(n6505), .ZN(n9798) );
  AND2_X1 U8060 ( .A1(n9801), .A2(n9798), .ZN(n9386) );
  OR2_X1 U8061 ( .A1(n6411), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6412) );
  AND2_X1 U8062 ( .A1(n6421), .A2(n6412), .ZN(n9788) );
  NAND2_X1 U8063 ( .A1(n9788), .A2(n4388), .ZN(n6418) );
  INV_X1 U8064 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U8065 ( .A1(n4386), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8066 ( .A1(n6404), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6414) );
  OAI211_X1 U8067 ( .C1(n6436), .C2(n10164), .A(n6415), .B(n6414), .ZN(n6416)
         );
  INV_X1 U8068 ( .A(n6416), .ZN(n6417) );
  INV_X1 U8069 ( .A(n9803), .ZN(n9309) );
  XNOR2_X1 U8070 ( .A(n9787), .B(n9309), .ZN(n9776) );
  NAND2_X1 U8071 ( .A1(n9787), .A2(n9309), .ZN(n9451) );
  NAND2_X1 U8072 ( .A1(n6421), .A2(n9204), .ZN(n6422) );
  NAND2_X1 U8073 ( .A1(n6430), .A2(n6422), .ZN(n9768) );
  INV_X1 U8074 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U8075 ( .A1(n6423), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U8076 ( .A1(n4386), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6424) );
  OAI211_X1 U8077 ( .C1(n6436), .C2(n10159), .A(n6425), .B(n6424), .ZN(n6426)
         );
  INV_X1 U8078 ( .A(n6426), .ZN(n6427) );
  INV_X1 U8079 ( .A(n9781), .ZN(n6429) );
  NAND2_X1 U8080 ( .A1(n9767), .A2(n6429), .ZN(n9459) );
  NAND2_X1 U8081 ( .A1(n9454), .A2(n9459), .ZN(n9757) );
  NAND2_X1 U8082 ( .A1(n6430), .A2(n9138), .ZN(n6432) );
  NAND2_X1 U8083 ( .A1(n6432), .A2(n6441), .ZN(n9751) );
  INV_X1 U8084 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U8085 ( .A1(n4386), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U8086 ( .A1(n6541), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6434) );
  OAI211_X1 U8087 ( .C1(n9071), .C2(n6436), .A(n6435), .B(n6434), .ZN(n6437)
         );
  INV_X1 U8088 ( .A(n6437), .ZN(n6438) );
  INV_X1 U8089 ( .A(n9762), .ZN(n6440) );
  NAND2_X1 U8090 ( .A1(n10153), .A2(n6440), .ZN(n9460) );
  NAND2_X1 U8091 ( .A1(n6533), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6448) );
  INV_X1 U8092 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8093 ( .A1(n6413), .A2(n9736), .ZN(n6447) );
  NAND2_X1 U8094 ( .A1(n4386), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U8095 ( .A1(n6423), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6445) );
  XNOR2_X1 U8096 ( .A(n9735), .B(n9402), .ZN(n9728) );
  INV_X1 U8097 ( .A(n9728), .ZN(n6449) );
  NAND2_X1 U8098 ( .A1(n9735), .A2(n9402), .ZN(n9524) );
  INV_X1 U8099 ( .A(n6451), .ZN(n6465) );
  NAND2_X1 U8100 ( .A1(n9557), .A2(n9540), .ZN(n9425) );
  INV_X1 U8101 ( .A(n9539), .ZN(n7087) );
  NAND2_X1 U8102 ( .A1(n6518), .A2(n7087), .ZN(n9547) );
  INV_X1 U8103 ( .A(n10014), .ZN(n6464) );
  NAND2_X1 U8104 ( .A1(n6274), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6459) );
  INV_X1 U8105 ( .A(n6454), .ZN(n6452) );
  NAND2_X1 U8106 ( .A1(n6452), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6534) );
  INV_X1 U8107 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U8108 ( .A1(n6454), .A2(n6453), .ZN(n6455) );
  NAND2_X1 U8109 ( .A1(n4389), .A2(n8081), .ZN(n6458) );
  NAND2_X1 U8110 ( .A1(n4386), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U8111 ( .A1(n6423), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6456) );
  INV_X1 U8112 ( .A(n10017), .ZN(n6461) );
  INV_X1 U8113 ( .A(n6095), .ZN(n7280) );
  INV_X1 U8114 ( .A(n10356), .ZN(n6460) );
  OAI21_X1 U8115 ( .B1(n6465), .B2(n6464), .A(n6463), .ZN(n6466) );
  INV_X1 U8116 ( .A(n7361), .ZN(n7481) );
  NAND2_X1 U8117 ( .A1(n7481), .A2(n10137), .ZN(n7476) );
  NAND2_X1 U8118 ( .A1(n7476), .A2(n9480), .ZN(n6468) );
  NAND2_X1 U8119 ( .A1(n6468), .A2(n4391), .ZN(n6471) );
  NAND3_X1 U8120 ( .A1(n6471), .A2(n7520), .A3(n6470), .ZN(n7755) );
  NAND2_X1 U8121 ( .A1(n9214), .A2(n10385), .ZN(n6473) );
  NAND3_X1 U8122 ( .A1(n7755), .A2(n6473), .A3(n7754), .ZN(n6475) );
  NAND2_X1 U8123 ( .A1(n10364), .A2(n9216), .ZN(n9314) );
  NAND2_X1 U8124 ( .A1(n9322), .A2(n9485), .ZN(n10105) );
  INV_X1 U8125 ( .A(n6473), .ZN(n7756) );
  NAND4_X1 U8126 ( .A1(n6475), .A2(n10366), .A3(n9314), .A4(n6474), .ZN(n6478)
         );
  NOR2_X1 U8127 ( .A1(n10364), .A2(n9216), .ZN(n9320) );
  NOR2_X1 U8128 ( .A1(n9569), .A2(n10360), .ZN(n6476) );
  NAND2_X1 U8129 ( .A1(n6478), .A2(n6477), .ZN(n10075) );
  NAND2_X1 U8130 ( .A1(n10075), .A2(n10074), .ZN(n6480) );
  NAND2_X1 U8131 ( .A1(n10350), .A2(n10397), .ZN(n6479) );
  NAND2_X1 U8132 ( .A1(n10055), .A2(n9343), .ZN(n10336) );
  NAND2_X1 U8133 ( .A1(n9344), .A2(n10033), .ZN(n10061) );
  NAND2_X1 U8134 ( .A1(n10334), .A2(n5986), .ZN(n6481) );
  NAND2_X1 U8135 ( .A1(n6482), .A2(n6481), .ZN(n10037) );
  NAND2_X1 U8136 ( .A1(n9496), .A2(n9347), .ZN(n10038) );
  NAND2_X1 U8137 ( .A1(n10037), .A2(n10038), .ZN(n9987) );
  NAND2_X1 U8138 ( .A1(n10058), .A2(n10416), .ZN(n9986) );
  NAND2_X1 U8139 ( .A1(n10227), .A2(n10016), .ZN(n6487) );
  INV_X1 U8140 ( .A(n6487), .ZN(n9437) );
  NOR2_X1 U8141 ( .A1(n10227), .A2(n10016), .ZN(n9438) );
  INV_X1 U8142 ( .A(n9438), .ZN(n6483) );
  INV_X1 U8143 ( .A(n10043), .ZN(n9994) );
  OR2_X1 U8144 ( .A1(n10023), .A2(n9994), .ZN(n9988) );
  AND2_X1 U8145 ( .A1(n6483), .A2(n9988), .ZN(n6484) );
  OR2_X1 U8146 ( .A1(n9437), .A2(n6484), .ZN(n6486) );
  AND2_X1 U8147 ( .A1(n9986), .A2(n6486), .ZN(n6485) );
  NAND2_X1 U8148 ( .A1(n9987), .A2(n6485), .ZN(n7992) );
  INV_X1 U8149 ( .A(n6486), .ZN(n6489) );
  AND2_X1 U8150 ( .A1(n10009), .A2(n6487), .ZN(n6488) );
  OR2_X1 U8151 ( .A1(n6489), .A2(n6488), .ZN(n7991) );
  AND2_X1 U8152 ( .A1(n7991), .A2(n5023), .ZN(n6490) );
  NAND2_X1 U8153 ( .A1(n7992), .A2(n6490), .ZN(n6492) );
  INV_X1 U8154 ( .A(n9968), .ZN(n9995) );
  OR2_X1 U8155 ( .A1(n7994), .A2(n9995), .ZN(n6491) );
  NAND2_X1 U8156 ( .A1(n6492), .A2(n6491), .ZN(n9961) );
  INV_X1 U8157 ( .A(n9941), .ZN(n9565) );
  OR2_X1 U8158 ( .A1(n10222), .A2(n9565), .ZN(n6493) );
  NAND2_X1 U8159 ( .A1(n9955), .A2(n9929), .ZN(n6494) );
  INV_X1 U8160 ( .A(n9942), .ZN(n9913) );
  OR2_X1 U8161 ( .A1(n10208), .A2(n9913), .ZN(n6495) );
  AND2_X2 U8162 ( .A1(n9514), .A2(n9516), .ZN(n9910) );
  INV_X1 U8163 ( .A(n9894), .ZN(n9928) );
  NAND2_X1 U8164 ( .A1(n10271), .A2(n9928), .ZN(n6497) );
  OR2_X1 U8165 ( .A1(n10197), .A2(n9914), .ZN(n6498) );
  NAND2_X1 U8166 ( .A1(n10197), .A2(n9914), .ZN(n6499) );
  NAND2_X1 U8167 ( .A1(n6500), .A2(n6499), .ZN(n9870) );
  OR2_X1 U8168 ( .A1(n9881), .A2(n9860), .ZN(n6501) );
  NAND2_X1 U8169 ( .A1(n9881), .A2(n9860), .ZN(n6502) );
  INV_X1 U8170 ( .A(n9843), .ZN(n6503) );
  OR2_X1 U8171 ( .A1(n9864), .A2(n9845), .ZN(n9840) );
  AND2_X1 U8172 ( .A1(n6503), .A2(n9840), .ZN(n6504) );
  NAND2_X1 U8173 ( .A1(n9841), .A2(n6504), .ZN(n9794) );
  NAND2_X1 U8174 ( .A1(n10180), .A2(n9861), .ZN(n9795) );
  NAND2_X1 U8175 ( .A1(n10256), .A2(n9846), .ZN(n9796) );
  NAND3_X1 U8176 ( .A1(n9794), .A2(n9795), .A3(n9796), .ZN(n6508) );
  NOR2_X1 U8177 ( .A1(n9808), .A2(n9826), .ZN(n6506) );
  AOI21_X1 U8178 ( .B1(n9823), .B2(n9796), .A(n6506), .ZN(n6507) );
  NAND2_X1 U8179 ( .A1(n6508), .A2(n6507), .ZN(n6510) );
  NAND2_X1 U8180 ( .A1(n9808), .A2(n9826), .ZN(n6509) );
  AND2_X1 U8181 ( .A1(n9787), .A2(n9803), .ZN(n6512) );
  NOR2_X1 U8182 ( .A1(n9767), .A2(n9781), .ZN(n6514) );
  NAND2_X1 U8183 ( .A1(n9767), .A2(n9781), .ZN(n6513) );
  AND2_X1 U8184 ( .A1(n10153), .A2(n9762), .ZN(n6515) );
  NOR2_X1 U8185 ( .A1(n9735), .A2(n9746), .ZN(n6517) );
  NAND2_X1 U8186 ( .A1(n9735), .A2(n9746), .ZN(n6516) );
  NAND2_X1 U8187 ( .A1(n6518), .A2(n9539), .ZN(n6882) );
  OR2_X1 U8188 ( .A1(n6884), .A2(n6882), .ZN(n10131) );
  INV_X1 U8189 ( .A(n10133), .ZN(n6520) );
  NAND3_X1 U8190 ( .A1(n10131), .A2(n6520), .A3(n6519), .ZN(n9939) );
  NAND2_X1 U8191 ( .A1(n7732), .A2(n9540), .ZN(n9315) );
  OAI211_X1 U8192 ( .C1(n6521), .C2(n9721), .A(n6522), .B(n10369), .ZN(n9718)
         );
  NOR2_X1 U8193 ( .A1(n7082), .A2(n6523), .ZN(n6524) );
  INV_X1 U8194 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6527) );
  NOR2_X1 U8195 ( .A1(n10442), .A2(n6527), .ZN(n6528) );
  NAND2_X1 U8196 ( .A1(n7106), .A2(n8818), .ZN(n9412) );
  INV_X1 U8197 ( .A(n9411), .ZN(n6531) );
  NOR2_X1 U8198 ( .A1(n9445), .A2(n6531), .ZN(n6532) );
  NAND2_X1 U8199 ( .A1(n6717), .A2(n6532), .ZN(n6719) );
  NAND2_X1 U8200 ( .A1(n6719), .A2(n9449), .ZN(n6540) );
  NAND2_X1 U8201 ( .A1(n4381), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6538) );
  INV_X1 U8202 ( .A(n6534), .ZN(n8021) );
  NAND2_X1 U8203 ( .A1(n6413), .A2(n8021), .ZN(n6537) );
  NAND2_X1 U8204 ( .A1(n4386), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8205 ( .A1(n6423), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6535) );
  NAND4_X1 U8206 ( .A1(n6538), .A2(n6537), .A3(n6536), .A4(n6535), .ZN(n9563)
         );
  INV_X1 U8207 ( .A(n9563), .ZN(n6539) );
  XNOR2_X1 U8208 ( .A(n6540), .B(n9446), .ZN(n6547) );
  NAND2_X1 U8209 ( .A1(n6274), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U8210 ( .A1(n4386), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U8211 ( .A1(n6404), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6542) );
  AND3_X1 U8212 ( .A1(n6544), .A2(n6543), .A3(n6542), .ZN(n9447) );
  OAI22_X1 U8213 ( .A1(n8818), .A2(n6460), .B1(n9447), .B2(n6545), .ZN(n6546)
         );
  OR2_X2 U8214 ( .A1(n6723), .A2(n6722), .ZN(n8015) );
  INV_X1 U8215 ( .A(n8015), .ZN(n6549) );
  NAND3_X1 U8216 ( .A1(n6549), .A2(n8016), .A3(n10424), .ZN(n6552) );
  INV_X1 U8217 ( .A(n8818), .ZN(n9564) );
  NAND2_X1 U8218 ( .A1(n7106), .A2(n9564), .ZN(n8014) );
  NAND4_X1 U8219 ( .A1(n8015), .A2(n9446), .A3(n10424), .A4(n8014), .ZN(n6551)
         );
  AOI211_X1 U8220 ( .C1(n6556), .C2(n5086), .A(n10214), .B(n9712), .ZN(n8025)
         );
  NOR3_X1 U8221 ( .A1(n9446), .A2(n10225), .A3(n8014), .ZN(n6550) );
  INV_X1 U8222 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U8223 ( .A1(n10440), .A2(n6553), .ZN(n6554) );
  NAND2_X1 U8224 ( .A1(n6555), .A2(n6554), .ZN(n6557) );
  INV_X1 U8225 ( .A(n6556), .ZN(n8023) );
  NAND2_X1 U8226 ( .A1(n6557), .A2(n5072), .ZN(P1_U3551) );
  INV_X1 U8227 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6558) );
  INV_X1 U8228 ( .A(n6860), .ZN(n6562) );
  OR2_X1 U8229 ( .A1(n6846), .A2(n6562), .ZN(n6563) );
  NAND2_X1 U8230 ( .A1(n6563), .A2(n6617), .ZN(n6619) );
  OR2_X1 U8231 ( .A1(n6619), .A2(n6564), .ZN(n6565) );
  NAND2_X1 U8232 ( .A1(n6565), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8233 ( .A(n6660), .ZN(n7737) );
  INV_X1 U8234 ( .A(n7583), .ZN(n7140) );
  XNOR2_X1 U8235 ( .A(n6567), .B(n6566), .ZN(n7563) );
  NOR2_X1 U8236 ( .A1(n10447), .A2(n10448), .ZN(n6568) );
  NAND2_X1 U8237 ( .A1(n5308), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6569) );
  OAI21_X1 U8238 ( .B1(n7386), .B2(n6568), .A(n6569), .ZN(n7389) );
  NAND2_X1 U8239 ( .A1(n7563), .A2(n7562), .ZN(n7561) );
  NAND2_X1 U8240 ( .A1(n6567), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U8241 ( .A1(n6571), .A2(n7157), .ZN(n7617) );
  XNOR2_X1 U8242 ( .A(n6631), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7616) );
  OR2_X1 U8243 ( .A1(n6631), .A2(n9140), .ZN(n6573) );
  INV_X1 U8244 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7401) );
  XNOR2_X1 U8245 ( .A(n7455), .B(n7509), .ZN(n7451) );
  XNOR2_X1 U8246 ( .A(n7583), .B(n7724), .ZN(n7578) );
  AOI21_X1 U8247 ( .B1(n6576), .B2(n7656), .A(n6577), .ZN(n7651) );
  NAND2_X1 U8248 ( .A1(n7651), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7741) );
  INV_X1 U8249 ( .A(n6577), .ZN(n7739) );
  INV_X1 U8250 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6659) );
  XNOR2_X1 U8251 ( .A(n6660), .B(n6659), .ZN(n7740) );
  AOI21_X1 U8252 ( .B1(n7741), .B2(n7739), .A(n7740), .ZN(n7738) );
  INV_X1 U8253 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8585) );
  XNOR2_X1 U8254 ( .A(n6671), .B(n8585), .ZN(n7924) );
  INV_X1 U8255 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8308) );
  XNOR2_X1 U8256 ( .A(n6680), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n8325) );
  INV_X1 U8257 ( .A(n6688), .ZN(n8348) );
  XNOR2_X1 U8258 ( .A(n6692), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8356) );
  INV_X1 U8259 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8549) );
  OR2_X1 U8260 ( .A1(n6692), .A2(n8549), .ZN(n6582) );
  INV_X1 U8261 ( .A(n6696), .ZN(n8378) );
  NAND2_X1 U8262 ( .A1(n6583), .A2(n8378), .ZN(n6584) );
  OAI21_X1 U8263 ( .B1(n6583), .B2(n8378), .A(n6584), .ZN(n8376) );
  INV_X1 U8264 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8540) );
  INV_X1 U8265 ( .A(n6584), .ZN(n8394) );
  NAND2_X1 U8266 ( .A1(n8406), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6586) );
  OAI21_X1 U8267 ( .B1(n8406), .B2(P2_REG2_REG_18__SCAN_IN), .A(n6586), .ZN(
        n6585) );
  INV_X1 U8268 ( .A(n6585), .ZN(n8393) );
  XNOR2_X1 U8269 ( .A(n6587), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6703) );
  OR2_X1 U8270 ( .A1(n6708), .A2(P2_U3151), .ZN(n6620) );
  INV_X1 U8271 ( .A(n6692), .ZN(n8360) );
  INV_X1 U8272 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U8273 ( .A1(n5308), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6592) );
  NAND2_X1 U8274 ( .A1(n7386), .A2(n6592), .ZN(n6591) );
  INV_X1 U8275 ( .A(n10448), .ZN(n9052) );
  NAND2_X1 U8276 ( .A1(n9052), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6589) );
  OR2_X1 U8277 ( .A1(n6589), .A2(n5308), .ZN(n6590) );
  NAND2_X1 U8278 ( .A1(n6591), .A2(n6590), .ZN(n7390) );
  NAND2_X1 U8279 ( .A1(n7390), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U8280 ( .A1(n6593), .A2(n6592), .ZN(n7565) );
  NAND2_X1 U8281 ( .A1(n6567), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U8282 ( .A1(n6595), .A2(n7157), .ZN(n6596) );
  NAND2_X1 U8283 ( .A1(n6597), .A2(n6596), .ZN(n7611) );
  INV_X1 U8284 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6598) );
  MUX2_X1 U8285 ( .A(n6598), .B(P2_REG1_REG_4__SCAN_IN), .S(n6631), .Z(n7612)
         );
  NAND2_X1 U8286 ( .A1(n7611), .A2(n7612), .ZN(n7610) );
  OR2_X1 U8287 ( .A1(n6631), .A2(n6598), .ZN(n6599) );
  XNOR2_X1 U8288 ( .A(n6600), .B(n7400), .ZN(n7399) );
  NAND2_X1 U8289 ( .A1(n7399), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U8290 ( .A1(n6600), .A2(n7152), .ZN(n6601) );
  NAND2_X1 U8291 ( .A1(n6602), .A2(n6601), .ZN(n7447) );
  MUX2_X1 U8292 ( .A(n6639), .B(P2_REG1_REG_6__SCAN_IN), .S(n7455), .Z(n7448)
         );
  NAND2_X1 U8293 ( .A1(n7447), .A2(n7448), .ZN(n7446) );
  NAND2_X1 U8294 ( .A1(n7149), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6603) );
  INV_X1 U8295 ( .A(n7637), .ZN(n7136) );
  NAND2_X1 U8296 ( .A1(n6604), .A2(n7136), .ZN(n6605) );
  XNOR2_X1 U8297 ( .A(n7583), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7576) );
  INV_X1 U8298 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7708) );
  OR2_X1 U8299 ( .A1(n7583), .A2(n7708), .ZN(n6606) );
  NAND2_X1 U8300 ( .A1(n6607), .A2(n6606), .ZN(n6608) );
  INV_X1 U8301 ( .A(n7656), .ZN(n7146) );
  NAND2_X1 U8302 ( .A1(n6608), .A2(n7146), .ZN(n6609) );
  XNOR2_X1 U8303 ( .A(n6660), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7736) );
  INV_X1 U8304 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8684) );
  INV_X1 U8305 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7889) );
  OAI22_X1 U8306 ( .A1(n7908), .A2(n7889), .B1(n7914), .B2(n6610), .ZN(n7922)
         );
  XNOR2_X1 U8307 ( .A(n6671), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7923) );
  INV_X1 U8308 ( .A(n6611), .ZN(n6612) );
  XOR2_X1 U8309 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n6680), .Z(n8323) );
  NAND2_X1 U8310 ( .A1(n6613), .A2(n8348), .ZN(n8370) );
  INV_X1 U8311 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8664) );
  XNOR2_X1 U8312 ( .A(n6692), .B(n8664), .ZN(n8368) );
  XNOR2_X1 U8313 ( .A(n6614), .B(n6696), .ZN(n8384) );
  INV_X1 U8314 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8661) );
  XNOR2_X1 U8315 ( .A(n6615), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8391) );
  XNOR2_X1 U8316 ( .A(n7503), .B(n8655), .ZN(n6702) );
  INV_X1 U8317 ( .A(n6616), .ZN(n10453) );
  INV_X1 U8318 ( .A(n6617), .ZN(n6621) );
  NOR2_X2 U8319 ( .A1(P2_U3150), .A2(n6621), .ZN(n10443) );
  NOR2_X1 U8320 ( .A1(n4383), .A2(P2_U3151), .ZN(n7977) );
  NAND2_X1 U8321 ( .A1(n7977), .A2(n6708), .ZN(n6618) );
  OR2_X1 U8322 ( .A1(n6619), .A2(n6618), .ZN(n6623) );
  INV_X1 U8323 ( .A(n6620), .ZN(n8808) );
  NAND2_X1 U8324 ( .A1(n6621), .A2(n8808), .ZN(n6622) );
  NAND2_X1 U8325 ( .A1(n6623), .A2(n6622), .ZN(n10444) );
  NAND2_X1 U8326 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8137) );
  OAI21_X1 U8327 ( .B1(n8401), .B2(n7503), .A(n8137), .ZN(n6711) );
  XNOR2_X1 U8328 ( .A(n6625), .B(n7386), .ZN(n7385) );
  NOR2_X1 U8329 ( .A1(n6624), .A2(n9052), .ZN(n10451) );
  NAND2_X1 U8330 ( .A1(n6625), .A2(n7386), .ZN(n6626) );
  MUX2_X1 U8331 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n4383), .Z(n6627) );
  XNOR2_X1 U8332 ( .A(n6627), .B(n6628), .ZN(n7571) );
  INV_X1 U8333 ( .A(n6627), .ZN(n6629) );
  NOR2_X1 U8334 ( .A1(n6629), .A2(n6628), .ZN(n6630) );
  MUX2_X1 U8335 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n4383), .Z(n6632) );
  XNOR2_X1 U8336 ( .A(n6632), .B(n4642), .ZN(n7556) );
  NAND2_X1 U8337 ( .A1(n7557), .A2(n7556), .ZN(n7625) );
  MUX2_X1 U8338 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4383), .Z(n6634) );
  INV_X1 U8339 ( .A(n6631), .ZN(n7615) );
  XNOR2_X1 U8340 ( .A(n6634), .B(n7615), .ZN(n7626) );
  NOR2_X1 U8341 ( .A1(n6632), .A2(n7157), .ZN(n7627) );
  NOR2_X1 U8342 ( .A1(n7626), .A2(n7627), .ZN(n6633) );
  NAND2_X1 U8343 ( .A1(n7625), .A2(n6633), .ZN(n7629) );
  NAND2_X1 U8344 ( .A1(n6634), .A2(n7615), .ZN(n6635) );
  NAND2_X1 U8345 ( .A1(n7629), .A2(n6635), .ZN(n7398) );
  MUX2_X1 U8346 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n4383), .Z(n6636) );
  XNOR2_X1 U8347 ( .A(n6636), .B(n7400), .ZN(n7397) );
  NAND2_X1 U8348 ( .A1(n7398), .A2(n7397), .ZN(n6638) );
  NAND2_X1 U8349 ( .A1(n6636), .A2(n7152), .ZN(n6637) );
  NAND2_X1 U8350 ( .A1(n6638), .A2(n6637), .ZN(n7445) );
  MUX2_X1 U8351 ( .A(n7509), .B(n6639), .S(n4383), .Z(n6640) );
  NAND2_X1 U8352 ( .A1(n6640), .A2(n7455), .ZN(n7641) );
  INV_X1 U8353 ( .A(n6640), .ZN(n6641) );
  NAND2_X1 U8354 ( .A1(n6641), .A2(n7149), .ZN(n6642) );
  NAND2_X1 U8355 ( .A1(n7641), .A2(n6642), .ZN(n7444) );
  NAND2_X1 U8356 ( .A1(n7642), .A2(n7641), .ZN(n6647) );
  INV_X1 U8357 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7768) );
  MUX2_X1 U8358 ( .A(n9035), .B(n7768), .S(n4383), .Z(n6643) );
  NAND2_X1 U8359 ( .A1(n6643), .A2(n7637), .ZN(n7581) );
  INV_X1 U8360 ( .A(n6643), .ZN(n6644) );
  NAND2_X1 U8361 ( .A1(n6644), .A2(n7136), .ZN(n6645) );
  NAND2_X1 U8362 ( .A1(n7581), .A2(n6645), .ZN(n7640) );
  INV_X1 U8363 ( .A(n7640), .ZN(n6646) );
  NAND2_X1 U8364 ( .A1(n7644), .A2(n7581), .ZN(n6652) );
  MUX2_X1 U8365 ( .A(n7724), .B(n7708), .S(n4383), .Z(n6648) );
  NAND2_X1 U8366 ( .A1(n6648), .A2(n7583), .ZN(n7653) );
  INV_X1 U8367 ( .A(n6648), .ZN(n6649) );
  NAND2_X1 U8368 ( .A1(n6649), .A2(n7140), .ZN(n6650) );
  NAND2_X1 U8369 ( .A1(n7653), .A2(n6650), .ZN(n7580) );
  INV_X1 U8370 ( .A(n7580), .ZN(n6651) );
  NAND2_X1 U8371 ( .A1(n6652), .A2(n6651), .ZN(n7654) );
  NAND2_X1 U8372 ( .A1(n7654), .A2(n7653), .ZN(n6658) );
  MUX2_X1 U8373 ( .A(n6653), .B(n7883), .S(n4383), .Z(n6654) );
  NAND2_X1 U8374 ( .A1(n6654), .A2(n7656), .ZN(n7747) );
  INV_X1 U8375 ( .A(n6654), .ZN(n6655) );
  NAND2_X1 U8376 ( .A1(n6655), .A2(n7146), .ZN(n6656) );
  NAND2_X1 U8377 ( .A1(n7747), .A2(n6656), .ZN(n7652) );
  INV_X1 U8378 ( .A(n7652), .ZN(n6657) );
  NAND2_X1 U8379 ( .A1(n6658), .A2(n6657), .ZN(n7748) );
  NAND2_X1 U8380 ( .A1(n7748), .A2(n7747), .ZN(n6665) );
  MUX2_X1 U8381 ( .A(n6659), .B(n8684), .S(n4383), .Z(n6661) );
  NAND2_X1 U8382 ( .A1(n6661), .A2(n6660), .ZN(n7911) );
  INV_X1 U8383 ( .A(n6661), .ZN(n6662) );
  NAND2_X1 U8384 ( .A1(n6662), .A2(n7737), .ZN(n6663) );
  NAND2_X1 U8385 ( .A1(n7911), .A2(n6663), .ZN(n7746) );
  INV_X1 U8386 ( .A(n7746), .ZN(n6664) );
  NAND2_X1 U8387 ( .A1(n7912), .A2(n7911), .ZN(n6668) );
  MUX2_X1 U8388 ( .A(n7903), .B(n7889), .S(n4383), .Z(n6666) );
  NAND2_X1 U8389 ( .A1(n6666), .A2(n7914), .ZN(n7930) );
  OAI21_X1 U8390 ( .B1(n7914), .B2(n6666), .A(n7930), .ZN(n7910) );
  INV_X1 U8391 ( .A(n7910), .ZN(n6667) );
  NAND2_X1 U8392 ( .A1(n6668), .A2(n6667), .ZN(n7931) );
  NAND2_X1 U8393 ( .A1(n7931), .A2(n7930), .ZN(n6673) );
  MUX2_X1 U8394 ( .A(n8585), .B(n6669), .S(n4383), .Z(n6670) );
  NAND2_X1 U8395 ( .A1(n6671), .A2(n6670), .ZN(n8312) );
  OAI21_X1 U8396 ( .B1(n6671), .B2(n6670), .A(n8312), .ZN(n7929) );
  INV_X1 U8397 ( .A(n7929), .ZN(n6672) );
  NAND2_X1 U8398 ( .A1(n6673), .A2(n6672), .ZN(n8313) );
  NAND2_X1 U8399 ( .A1(n8313), .A2(n8312), .ZN(n6677) );
  INV_X1 U8400 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7945) );
  MUX2_X1 U8401 ( .A(n8308), .B(n7945), .S(n4383), .Z(n6675) );
  NAND2_X1 U8402 ( .A1(n6674), .A2(n6675), .ZN(n8333) );
  OR2_X1 U8403 ( .A1(n6675), .A2(n6674), .ZN(n6676) );
  AND2_X1 U8404 ( .A1(n8333), .A2(n6676), .ZN(n8310) );
  NAND2_X1 U8405 ( .A1(n8334), .A2(n8333), .ZN(n6684) );
  MUX2_X1 U8406 ( .A(n6678), .B(n8672), .S(n4383), .Z(n6679) );
  NAND2_X1 U8407 ( .A1(n6679), .A2(n6680), .ZN(n6685) );
  INV_X1 U8408 ( .A(n6679), .ZN(n6681) );
  INV_X1 U8409 ( .A(n6680), .ZN(n8331) );
  NAND2_X1 U8410 ( .A1(n6681), .A2(n8331), .ZN(n6682) );
  NAND2_X1 U8411 ( .A1(n6685), .A2(n6682), .ZN(n8332) );
  INV_X1 U8412 ( .A(n8332), .ZN(n6683) );
  NAND2_X1 U8413 ( .A1(n6684), .A2(n6683), .ZN(n8336) );
  NAND2_X1 U8414 ( .A1(n8336), .A2(n6685), .ZN(n8345) );
  MUX2_X1 U8415 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n4383), .Z(n6686) );
  XNOR2_X1 U8416 ( .A(n6688), .B(n6686), .ZN(n8344) );
  NAND2_X1 U8417 ( .A1(n8345), .A2(n8344), .ZN(n8343) );
  INV_X1 U8418 ( .A(n6686), .ZN(n6687) );
  NAND2_X1 U8419 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  NAND2_X1 U8420 ( .A1(n8343), .A2(n6689), .ZN(n8364) );
  MUX2_X1 U8421 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n4383), .Z(n6690) );
  NAND2_X1 U8422 ( .A1(n8360), .A2(n6690), .ZN(n8362) );
  NAND2_X1 U8423 ( .A1(n8364), .A2(n8362), .ZN(n6693) );
  INV_X1 U8424 ( .A(n6690), .ZN(n6691) );
  NAND2_X1 U8425 ( .A1(n6692), .A2(n6691), .ZN(n8361) );
  NAND2_X1 U8426 ( .A1(n6693), .A2(n8361), .ZN(n8379) );
  MUX2_X1 U8427 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n4383), .Z(n6694) );
  XNOR2_X1 U8428 ( .A(n6696), .B(n6694), .ZN(n8380) );
  INV_X1 U8429 ( .A(n6694), .ZN(n6695) );
  AND2_X1 U8430 ( .A1(n6696), .A2(n6695), .ZN(n6697) );
  INV_X1 U8431 ( .A(n6701), .ZN(n6699) );
  MUX2_X1 U8432 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n4383), .Z(n6700) );
  INV_X1 U8433 ( .A(n6700), .ZN(n6698) );
  NAND2_X1 U8434 ( .A1(n6699), .A2(n6698), .ZN(n8398) );
  AND2_X1 U8435 ( .A1(n6701), .A2(n6700), .ZN(n8400) );
  INV_X1 U8436 ( .A(n6702), .ZN(n6705) );
  INV_X1 U8437 ( .A(n6703), .ZN(n6704) );
  MUX2_X1 U8438 ( .A(n6705), .B(n6704), .S(n6203), .Z(n6706) );
  XNOR2_X1 U8439 ( .A(n6707), .B(n6706), .ZN(n6709) );
  NAND2_X1 U8440 ( .A1(n8305), .A2(n6708), .ZN(n8404) );
  NOR2_X1 U8441 ( .A1(n6709), .A2(n8404), .ZN(n6710) );
  AOI211_X1 U8442 ( .C1(P2_ADDR_REG_19__SCAN_IN), .C2(n10443), .A(n6711), .B(
        n6710), .ZN(n6712) );
  NAND2_X1 U8443 ( .A1(n7114), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U8444 ( .A1(n6717), .A2(n9411), .ZN(n6718) );
  AOI22_X1 U8445 ( .A1(n10017), .A2(n9563), .B1(n9732), .B2(n10356), .ZN(n6720) );
  NAND2_X1 U8446 ( .A1(n6721), .A2(n6720), .ZN(n8086) );
  NAND2_X1 U8447 ( .A1(n6723), .A2(n6722), .ZN(n6724) );
  AOI21_X1 U8448 ( .B1(n6522), .B2(n7106), .A(n10214), .ZN(n6725) );
  AND2_X1 U8449 ( .A1(n6725), .A2(n5086), .ZN(n8080) );
  OR2_X1 U8450 ( .A1(n6732), .A2(n7114), .ZN(n6729) );
  OR2_X1 U8451 ( .A1(n10430), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U8452 ( .A1(n6729), .A2(n6728), .ZN(n6731) );
  INV_X1 U8453 ( .A(n7106), .ZN(n8084) );
  NAND2_X1 U8454 ( .A1(n7106), .A2(n6140), .ZN(n6730) );
  NAND2_X1 U8455 ( .A1(n6731), .A2(n6730), .ZN(P1_U3518) );
  OR2_X1 U8456 ( .A1(n10442), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U8457 ( .A1(n7106), .A2(n6526), .ZN(n6734) );
  NAND2_X1 U8458 ( .A1(n6735), .A2(n6734), .ZN(P1_U3550) );
  INV_X1 U8459 ( .A(n10493), .ZN(n6736) );
  NOR2_X1 U8460 ( .A1(n6737), .A2(n6736), .ZN(n6738) );
  NAND2_X1 U8461 ( .A1(n6740), .A2(n8796), .ZN(n7119) );
  INV_X1 U8462 ( .A(n6745), .ZN(n6741) );
  OR2_X1 U8463 ( .A1(n7690), .A2(n6742), .ZN(n6743) );
  OAI21_X1 U8464 ( .B1(n8795), .B2(n6848), .A(n6872), .ZN(n6744) );
  NAND2_X1 U8465 ( .A1(n6865), .A2(n6744), .ZN(n6749) );
  NAND2_X1 U8466 ( .A1(n6759), .A2(n6745), .ZN(n6746) );
  NAND3_X1 U8467 ( .A1(n6848), .A2(n6846), .A3(n10488), .ZN(n6747) );
  NAND2_X1 U8468 ( .A1(n8567), .A2(n6747), .ZN(n6858) );
  NAND3_X1 U8469 ( .A1(n6873), .A2(n7160), .A3(n6858), .ZN(n6748) );
  INV_X1 U8470 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6750) );
  NOR2_X1 U8471 ( .A1(n10501), .A2(n6750), .ZN(n6751) );
  OAI21_X1 U8472 ( .B1(n7123), .B2(n10499), .A(n6753), .ZN(P2_U3456) );
  AND2_X1 U8473 ( .A1(n6756), .A2(n6755), .ZN(n6757) );
  OAI21_X2 U8474 ( .B1(n6759), .B2(n6758), .A(n6757), .ZN(n6770) );
  OR2_X1 U8475 ( .A1(n6770), .A2(n10472), .ZN(n6760) );
  NAND2_X1 U8476 ( .A1(n6760), .A2(n7415), .ZN(n7335) );
  XNOR2_X1 U8477 ( .A(n4376), .B(n6761), .ZN(n6763) );
  XNOR2_X1 U8478 ( .A(n6763), .B(n8304), .ZN(n7334) );
  NAND2_X1 U8479 ( .A1(n7335), .A2(n7334), .ZN(n6765) );
  NAND2_X1 U8480 ( .A1(n6763), .A2(n6150), .ZN(n6764) );
  NAND2_X1 U8481 ( .A1(n6765), .A2(n6764), .ZN(n7327) );
  XNOR2_X1 U8482 ( .A(n6770), .B(n7328), .ZN(n6766) );
  XNOR2_X1 U8483 ( .A(n6766), .B(n7336), .ZN(n7326) );
  NAND2_X1 U8484 ( .A1(n7327), .A2(n7326), .ZN(n6769) );
  INV_X1 U8485 ( .A(n6766), .ZN(n6767) );
  NAND2_X1 U8486 ( .A1(n6767), .A2(n7336), .ZN(n6768) );
  NAND2_X1 U8487 ( .A1(n6769), .A2(n6768), .ZN(n7351) );
  INV_X1 U8488 ( .A(n7351), .ZN(n6773) );
  INV_X2 U8489 ( .A(n6770), .ZN(n8089) );
  INV_X4 U8490 ( .A(n8089), .ZN(n6837) );
  XNOR2_X1 U8491 ( .A(n6774), .B(n6771), .ZN(n7352) );
  NAND2_X1 U8492 ( .A1(n6774), .A2(n6771), .ZN(n6775) );
  XNOR2_X1 U8493 ( .A(n6776), .B(n6837), .ZN(n6778) );
  INV_X1 U8494 ( .A(n6778), .ZN(n6779) );
  NAND2_X1 U8495 ( .A1(n6779), .A2(n7348), .ZN(n6780) );
  XNOR2_X1 U8496 ( .A(n6837), .B(n10489), .ZN(n6781) );
  XNOR2_X1 U8497 ( .A(n6781), .B(n7495), .ZN(n7434) );
  INV_X1 U8498 ( .A(n6781), .ZN(n6782) );
  NAND2_X1 U8499 ( .A1(n6782), .A2(n7495), .ZN(n6783) );
  XNOR2_X1 U8500 ( .A(n6837), .B(n7512), .ZN(n6784) );
  XNOR2_X1 U8501 ( .A(n6784), .B(n7700), .ZN(n7490) );
  INV_X1 U8502 ( .A(n6784), .ZN(n6785) );
  NAND2_X1 U8503 ( .A1(n6785), .A2(n8301), .ZN(n6786) );
  NAND2_X1 U8504 ( .A1(n7492), .A2(n6786), .ZN(n7713) );
  XNOR2_X1 U8505 ( .A(n6837), .B(n7814), .ZN(n6787) );
  XNOR2_X1 U8506 ( .A(n6787), .B(n8300), .ZN(n7714) );
  OR2_X1 U8507 ( .A1(n6787), .A2(n8300), .ZN(n6788) );
  XNOR2_X1 U8508 ( .A(n6837), .B(n7780), .ZN(n7771) );
  XNOR2_X1 U8509 ( .A(n7868), .B(n6837), .ZN(n6789) );
  XNOR2_X1 U8510 ( .A(n6789), .B(n8608), .ZN(n7804) );
  INV_X1 U8511 ( .A(n6789), .ZN(n6790) );
  NAND2_X1 U8512 ( .A1(n6790), .A2(n8608), .ZN(n6791) );
  XNOR2_X1 U8513 ( .A(n8602), .B(n6837), .ZN(n8124) );
  XNOR2_X1 U8514 ( .A(n8579), .B(n8089), .ZN(n8158) );
  NAND2_X1 U8515 ( .A1(n8158), .A2(n8607), .ZN(n8159) );
  OAI21_X1 U8516 ( .B1(n8156), .B2(n8124), .A(n8159), .ZN(n6797) );
  XNOR2_X1 U8517 ( .A(n8677), .B(n6837), .ZN(n6798) );
  XNOR2_X1 U8518 ( .A(n6798), .B(n8246), .ZN(n8161) );
  AOI21_X1 U8519 ( .B1(n8124), .B2(n8156), .A(n8157), .ZN(n6794) );
  NAND3_X1 U8520 ( .A1(n8124), .A2(n8156), .A3(n8157), .ZN(n6793) );
  OAI21_X1 U8521 ( .B1(n8158), .B2(n6794), .A(n6793), .ZN(n6795) );
  INV_X1 U8522 ( .A(n6798), .ZN(n6799) );
  NAND2_X1 U8523 ( .A1(n6799), .A2(n8297), .ZN(n6800) );
  XNOR2_X1 U8524 ( .A(n8227), .B(n6837), .ZN(n6801) );
  NAND2_X1 U8525 ( .A1(n6801), .A2(n8163), .ZN(n8219) );
  INV_X1 U8526 ( .A(n6801), .ZN(n6802) );
  NAND2_X1 U8527 ( .A1(n6802), .A2(n8583), .ZN(n8220) );
  XNOR2_X1 U8528 ( .A(n8785), .B(n6837), .ZN(n6803) );
  XNOR2_X1 U8529 ( .A(n6803), .B(n8556), .ZN(n8107) );
  NAND2_X1 U8530 ( .A1(n6803), .A2(n8556), .ZN(n6804) );
  XNOR2_X1 U8531 ( .A(n8779), .B(n6837), .ZN(n6806) );
  XNOR2_X1 U8532 ( .A(n6806), .B(n6805), .ZN(n8282) );
  INV_X1 U8533 ( .A(n6806), .ZN(n6807) );
  NAND2_X1 U8534 ( .A1(n6807), .A2(n8570), .ZN(n6808) );
  XNOR2_X1 U8535 ( .A(n8772), .B(n6837), .ZN(n6811) );
  XNOR2_X1 U8536 ( .A(n6811), .B(n8557), .ZN(n8180) );
  XNOR2_X1 U8537 ( .A(n8767), .B(n6837), .ZN(n6810) );
  OR2_X1 U8538 ( .A1(n8180), .A2(n6812), .ZN(n8188) );
  XNOR2_X1 U8539 ( .A(n8761), .B(n6837), .ZN(n6809) );
  XNOR2_X1 U8540 ( .A(n6809), .B(n8536), .ZN(n8257) );
  INV_X1 U8541 ( .A(n8257), .ZN(n6814) );
  NAND2_X1 U8542 ( .A1(n6810), .A2(n8261), .ZN(n6813) );
  AND2_X1 U8543 ( .A1(n6813), .A2(n8190), .ZN(n8254) );
  XNOR2_X1 U8544 ( .A(n8755), .B(n6837), .ZN(n8134) );
  AND2_X1 U8545 ( .A1(n8134), .A2(n8214), .ZN(n6816) );
  INV_X1 U8546 ( .A(n8134), .ZN(n6817) );
  NAND2_X1 U8547 ( .A1(n6817), .A2(n8527), .ZN(n6818) );
  XNOR2_X1 U8548 ( .A(n8041), .B(n8089), .ZN(n6820) );
  NAND2_X1 U8549 ( .A1(n6820), .A2(n8497), .ZN(n8145) );
  INV_X1 U8550 ( .A(n6820), .ZN(n6821) );
  NAND2_X1 U8551 ( .A1(n6821), .A2(n8515), .ZN(n6822) );
  NAND2_X1 U8552 ( .A1(n8145), .A2(n6822), .ZN(n8210) );
  OR2_X2 U8553 ( .A1(n8209), .A2(n8210), .ZN(n8144) );
  NAND2_X1 U8554 ( .A1(n8144), .A2(n8145), .ZN(n8148) );
  XNOR2_X1 U8555 ( .A(n8499), .B(n6837), .ZN(n6823) );
  NAND2_X1 U8556 ( .A1(n6823), .A2(n8483), .ZN(n8231) );
  INV_X1 U8557 ( .A(n6823), .ZN(n6824) );
  INV_X1 U8558 ( .A(n8483), .ZN(n8294) );
  NAND2_X1 U8559 ( .A1(n6824), .A2(n8294), .ZN(n6825) );
  AND2_X1 U8560 ( .A1(n8231), .A2(n6825), .ZN(n8147) );
  XNOR2_X1 U8561 ( .A(n8230), .B(n6837), .ZN(n6828) );
  XNOR2_X1 U8562 ( .A(n6828), .B(n8473), .ZN(n8232) );
  AND2_X1 U8563 ( .A1(n8147), .A2(n8232), .ZN(n6827) );
  INV_X1 U8564 ( .A(n8232), .ZN(n6826) );
  NAND2_X1 U8565 ( .A1(n6828), .A2(n8496), .ZN(n6829) );
  XNOR2_X1 U8566 ( .A(n8740), .B(n6837), .ZN(n6834) );
  AND2_X1 U8567 ( .A1(n6834), .A2(n8484), .ZN(n6830) );
  XNOR2_X1 U8568 ( .A(n8734), .B(n6837), .ZN(n6831) );
  NAND2_X1 U8569 ( .A1(n6831), .A2(n8119), .ZN(n8170) );
  INV_X1 U8570 ( .A(n6831), .ZN(n6832) );
  NAND2_X1 U8571 ( .A1(n6832), .A2(n8474), .ZN(n6833) );
  NAND2_X1 U8572 ( .A1(n8170), .A2(n6833), .ZN(n8199) );
  INV_X1 U8573 ( .A(n6834), .ZN(n8114) );
  AND2_X1 U8574 ( .A1(n8114), .A2(n8457), .ZN(n6835) );
  NOR2_X1 U8575 ( .A1(n8199), .A2(n6835), .ZN(n6836) );
  XNOR2_X1 U8576 ( .A(n8728), .B(n6837), .ZN(n6838) );
  NAND2_X1 U8577 ( .A1(n6838), .A2(n8275), .ZN(n8266) );
  INV_X1 U8578 ( .A(n6838), .ZN(n6839) );
  NAND2_X1 U8579 ( .A1(n6839), .A2(n8458), .ZN(n6840) );
  NAND2_X1 U8580 ( .A1(n6841), .A2(n8171), .ZN(n8173) );
  NAND2_X1 U8581 ( .A1(n8173), .A2(n8266), .ZN(n6842) );
  XNOR2_X1 U8582 ( .A(n8722), .B(n6837), .ZN(n6844) );
  XNOR2_X1 U8583 ( .A(n6844), .B(n8448), .ZN(n8267) );
  NAND2_X1 U8584 ( .A1(n6844), .A2(n6843), .ZN(n6845) );
  XNOR2_X1 U8585 ( .A(n8717), .B(n6837), .ZN(n8096) );
  XNOR2_X1 U8586 ( .A(n8096), .B(n8421), .ZN(n6852) );
  NOR2_X2 U8587 ( .A1(n6853), .A2(n6852), .ZN(n8102) );
  NAND3_X1 U8588 ( .A1(n6865), .A2(n6846), .A3(n10488), .ZN(n6847) );
  NAND2_X1 U8589 ( .A1(n6847), .A2(n6848), .ZN(n6851) );
  INV_X1 U8590 ( .A(n6848), .ZN(n6849) );
  NAND2_X1 U8591 ( .A1(n6867), .A2(n6849), .ZN(n6862) );
  AND2_X1 U8592 ( .A1(n6862), .A2(n7160), .ZN(n6850) );
  INV_X1 U8593 ( .A(n6854), .ZN(n6880) );
  OR2_X1 U8594 ( .A1(n6865), .A2(n10457), .ZN(n6855) );
  NAND2_X1 U8595 ( .A1(n8717), .A2(n8263), .ZN(n6879) );
  INV_X1 U8596 ( .A(n6871), .ZN(n6856) );
  NOR2_X1 U8597 ( .A1(n6872), .A2(n6856), .ZN(n6857) );
  INV_X1 U8598 ( .A(n6858), .ZN(n6864) );
  AND4_X1 U8599 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6863)
         );
  OAI21_X1 U8600 ( .B1(n6865), .B2(n6864), .A(n6863), .ZN(n6866) );
  NAND2_X1 U8601 ( .A1(n6866), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6870) );
  NAND2_X1 U8602 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  AOI22_X1 U8603 ( .A1(n8434), .A2(n8290), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6876) );
  NOR2_X1 U8604 ( .A1(n6872), .A2(n6871), .ZN(n6874) );
  NAND2_X1 U8605 ( .A1(n8448), .A2(n8286), .ZN(n6875) );
  OAI211_X1 U8606 ( .C1(n8090), .C2(n8288), .A(n6876), .B(n6875), .ZN(n6877)
         );
  INV_X1 U8607 ( .A(n6877), .ZN(n6878) );
  OAI21_X1 U8608 ( .B1(n8102), .B2(n6880), .A(n5087), .ZN(P2_U3154) );
  OR2_X1 U8609 ( .A1(n9551), .A2(n6882), .ZN(n9950) );
  NAND3_X1 U8610 ( .A1(n6886), .A2(n6884), .A3(n6882), .ZN(n6934) );
  NAND2_X1 U8611 ( .A1(n10208), .A2(n7045), .ZN(n6888) );
  INV_X1 U8612 ( .A(n6882), .ZN(n6885) );
  OR2_X1 U8613 ( .A1(n9942), .A2(n7070), .ZN(n6887) );
  NAND2_X1 U8614 ( .A1(n6888), .A2(n6887), .ZN(n6889) );
  XNOR2_X1 U8615 ( .A(n6889), .B(n7043), .ZN(n6983) );
  NAND2_X1 U8616 ( .A1(n10208), .A2(n7002), .ZN(n6891) );
  OR2_X1 U8617 ( .A1(n9942), .A2(n7076), .ZN(n6890) );
  NAND2_X1 U8618 ( .A1(n6891), .A2(n6890), .ZN(n9298) );
  NAND2_X1 U8619 ( .A1(n10364), .A2(n7002), .ZN(n6893) );
  NAND2_X1 U8620 ( .A1(n9216), .A2(n7045), .ZN(n6892) );
  NAND2_X1 U8621 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  XNOR2_X1 U8622 ( .A(n6894), .B(n7073), .ZN(n6923) );
  INV_X2 U8623 ( .A(n7076), .ZN(n7049) );
  AND2_X1 U8624 ( .A1(n9216), .A2(n7002), .ZN(n6895) );
  AOI21_X1 U8625 ( .B1(n10364), .B2(n7049), .A(n6895), .ZN(n6924) );
  XNOR2_X1 U8626 ( .A(n6923), .B(n6924), .ZN(n9209) );
  OAI22_X1 U8627 ( .A1(n9214), .A2(n7070), .B1(n10385), .B2(n6897), .ZN(n6896)
         );
  XNOR2_X1 U8628 ( .A(n6896), .B(n7043), .ZN(n6916) );
  OAI22_X1 U8629 ( .A1(n9214), .A2(n7076), .B1(n10385), .B2(n7070), .ZN(n6915)
         );
  NOR2_X1 U8630 ( .A1(n6916), .A2(n6915), .ZN(n9210) );
  OAI22_X1 U8631 ( .A1(n9480), .A2(n7076), .B1(n10122), .B2(n7070), .ZN(n6899)
         );
  XNOR2_X1 U8632 ( .A(n6898), .B(n7043), .ZN(n6900) );
  NOR2_X1 U8633 ( .A1(n6899), .A2(n6900), .ZN(n6904) );
  INV_X1 U8634 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7178) );
  AOI21_X1 U8635 ( .B1(n7002), .B2(n7481), .A(n6902), .ZN(n6903) );
  OAI21_X1 U8636 ( .B1(n7175), .B2(n7178), .A(n6903), .ZN(n7274) );
  AOI22_X1 U8637 ( .A1(n7273), .A2(n7274), .B1(n7073), .B2(n6903), .ZN(n7359)
         );
  NAND2_X1 U8638 ( .A1(n7358), .A2(n7359), .ZN(n7357) );
  INV_X1 U8639 ( .A(n6904), .ZN(n7377) );
  NAND2_X1 U8640 ( .A1(n9571), .A2(n7002), .ZN(n6907) );
  NAND2_X1 U8641 ( .A1(n7518), .A2(n6905), .ZN(n6906) );
  NAND2_X1 U8642 ( .A1(n6907), .A2(n6906), .ZN(n6908) );
  XNOR2_X1 U8643 ( .A(n6908), .B(n7073), .ZN(n6912) );
  NAND2_X1 U8644 ( .A1(n9571), .A2(n7049), .ZN(n6910) );
  NAND2_X1 U8645 ( .A1(n7518), .A2(n7002), .ZN(n6909) );
  AND2_X1 U8646 ( .A1(n6910), .A2(n6909), .ZN(n6911) );
  NAND2_X1 U8647 ( .A1(n6912), .A2(n6911), .ZN(n6913) );
  NAND2_X1 U8648 ( .A1(n6913), .A2(n5085), .ZN(n7376) );
  AOI21_X2 U8649 ( .B1(n7357), .B2(n7377), .A(n7376), .ZN(n7379) );
  INV_X1 U8650 ( .A(n6913), .ZN(n6914) );
  XNOR2_X1 U8651 ( .A(n6916), .B(n6915), .ZN(n7529) );
  OAI22_X1 U8652 ( .A1(n10073), .A2(n7070), .B1(n10392), .B2(n6897), .ZN(n6917) );
  XNOR2_X1 U8653 ( .A(n6917), .B(n7043), .ZN(n7822) );
  INV_X1 U8654 ( .A(n7822), .ZN(n7820) );
  OR2_X1 U8655 ( .A1(n10073), .A2(n7076), .ZN(n6919) );
  NAND2_X1 U8656 ( .A1(n10360), .A2(n7002), .ZN(n6918) );
  NAND2_X1 U8657 ( .A1(n6919), .A2(n6918), .ZN(n6927) );
  INV_X1 U8658 ( .A(n6927), .ZN(n7853) );
  OAI22_X1 U8659 ( .A1(n10350), .A2(n7070), .B1(n10397), .B2(n6897), .ZN(n6920) );
  XNOR2_X1 U8660 ( .A(n6920), .B(n7073), .ZN(n6930) );
  INV_X1 U8661 ( .A(n6930), .ZN(n7857) );
  OR2_X1 U8662 ( .A1(n10350), .A2(n7076), .ZN(n6922) );
  NAND2_X1 U8663 ( .A1(n10079), .A2(n7002), .ZN(n6921) );
  NAND2_X1 U8664 ( .A1(n6922), .A2(n6921), .ZN(n7856) );
  NAND2_X1 U8665 ( .A1(n7857), .A2(n7856), .ZN(n7855) );
  INV_X1 U8666 ( .A(n6923), .ZN(n6926) );
  INV_X1 U8667 ( .A(n6924), .ZN(n6925) );
  NAND2_X1 U8668 ( .A1(n6926), .A2(n6925), .ZN(n7821) );
  OAI211_X1 U8669 ( .C1(n7820), .C2(n7853), .A(n7855), .B(n7821), .ZN(n6932)
         );
  OAI21_X1 U8670 ( .B1(n7822), .B2(n6927), .A(n7856), .ZN(n6929) );
  NOR3_X1 U8671 ( .A1(n7822), .A2(n7856), .A3(n6927), .ZN(n6928) );
  AOI21_X1 U8672 ( .B1(n6930), .B2(n6929), .A(n6928), .ZN(n6931) );
  OAI21_X1 U8673 ( .B1(n7824), .B2(n6932), .A(n6931), .ZN(n6933) );
  OAI22_X1 U8674 ( .A1(n10072), .A2(n7076), .B1(n10403), .B2(n7070), .ZN(n6937) );
  AOI22_X1 U8675 ( .A1(n9567), .A2(n7002), .B1(n10343), .B2(n7045), .ZN(n6935)
         );
  XNOR2_X1 U8676 ( .A(n6935), .B(n7043), .ZN(n6936) );
  XOR2_X1 U8677 ( .A(n6937), .B(n6936), .Z(n7794) );
  AOI22_X1 U8678 ( .A1(n10018), .A2(n7002), .B1(n10050), .B2(n7045), .ZN(n6938) );
  XOR2_X1 U8679 ( .A(n7043), .B(n6938), .Z(n9222) );
  OR2_X1 U8680 ( .A1(n10058), .A2(n7076), .ZN(n6940) );
  NAND2_X1 U8681 ( .A1(n10050), .A2(n7002), .ZN(n6939) );
  NAND2_X1 U8682 ( .A1(n6940), .A2(n6939), .ZN(n9223) );
  OAI22_X1 U8683 ( .A1(n10334), .A2(n7070), .B1(n5986), .B2(n6897), .ZN(n6941)
         );
  XNOR2_X1 U8684 ( .A(n6941), .B(n7043), .ZN(n6944) );
  OR2_X1 U8685 ( .A1(n10334), .A2(n7076), .ZN(n6943) );
  NAND2_X1 U8686 ( .A1(n10064), .A2(n7002), .ZN(n6942) );
  NAND2_X1 U8687 ( .A1(n6943), .A2(n6942), .ZN(n7963) );
  OAI22_X1 U8688 ( .A1(n9222), .A2(n9223), .B1(n6944), .B2(n7963), .ZN(n6948)
         );
  INV_X1 U8689 ( .A(n6944), .ZN(n9221) );
  INV_X1 U8690 ( .A(n7963), .ZN(n6945) );
  NOR2_X1 U8691 ( .A1(n9221), .A2(n6945), .ZN(n6946) );
  OAI21_X1 U8692 ( .B1(n6946), .B2(n9223), .A(n9222), .ZN(n6947) );
  NAND2_X1 U8693 ( .A1(n10227), .A2(n7045), .ZN(n6950) );
  NAND2_X1 U8694 ( .A1(n10016), .A2(n7002), .ZN(n6949) );
  NAND2_X1 U8695 ( .A1(n6950), .A2(n6949), .ZN(n6951) );
  XNOR2_X1 U8696 ( .A(n6951), .B(n7043), .ZN(n9263) );
  INV_X1 U8697 ( .A(n9263), .ZN(n6959) );
  NAND2_X1 U8698 ( .A1(n10227), .A2(n7002), .ZN(n6953) );
  NAND2_X1 U8699 ( .A1(n10016), .A2(n7049), .ZN(n6952) );
  NAND2_X1 U8700 ( .A1(n6953), .A2(n6952), .ZN(n9262) );
  INV_X1 U8701 ( .A(n9262), .ZN(n6964) );
  NAND2_X1 U8702 ( .A1(n10023), .A2(n7045), .ZN(n6955) );
  OR2_X1 U8703 ( .A1(n10043), .A2(n7070), .ZN(n6954) );
  NAND2_X1 U8704 ( .A1(n6955), .A2(n6954), .ZN(n6956) );
  XNOR2_X1 U8705 ( .A(n6956), .B(n7043), .ZN(n9261) );
  INV_X1 U8706 ( .A(n9261), .ZN(n8847) );
  NAND2_X1 U8707 ( .A1(n10023), .A2(n7002), .ZN(n6958) );
  OR2_X1 U8708 ( .A1(n10043), .A2(n7076), .ZN(n6957) );
  NAND2_X1 U8709 ( .A1(n6958), .A2(n6957), .ZN(n6960) );
  INV_X1 U8710 ( .A(n6960), .ZN(n8849) );
  AOI22_X1 U8711 ( .A1(n6959), .A2(n6964), .B1(n8847), .B2(n8849), .ZN(n6966)
         );
  AND2_X1 U8712 ( .A1(n9261), .A2(n6960), .ZN(n6961) );
  INV_X1 U8713 ( .A(n6961), .ZN(n6963) );
  OAI21_X1 U8714 ( .B1(n6961), .B2(n9262), .A(n9263), .ZN(n6962) );
  OAI21_X1 U8715 ( .B1(n6964), .B2(n6963), .A(n6962), .ZN(n6965) );
  AOI22_X1 U8716 ( .A1(n7994), .A2(n7045), .B1(n7002), .B2(n9995), .ZN(n6967)
         );
  XOR2_X1 U8717 ( .A(n7043), .B(n6967), .Z(n6969) );
  OAI22_X1 U8718 ( .A1(n9981), .A2(n7070), .B1(n9968), .B2(n7076), .ZN(n6968)
         );
  NOR2_X1 U8719 ( .A1(n6969), .A2(n6968), .ZN(n6970) );
  AOI21_X1 U8720 ( .B1(n6969), .B2(n6968), .A(n6970), .ZN(n7981) );
  NAND2_X1 U8721 ( .A1(n7980), .A2(n7981), .ZN(n7979) );
  INV_X1 U8722 ( .A(n6970), .ZN(n6971) );
  NAND2_X1 U8723 ( .A1(n10222), .A2(n7045), .ZN(n6973) );
  OR2_X1 U8724 ( .A1(n9941), .A2(n7070), .ZN(n6972) );
  NAND2_X1 U8725 ( .A1(n6973), .A2(n6972), .ZN(n6974) );
  XNOR2_X1 U8726 ( .A(n6974), .B(n7043), .ZN(n6977) );
  AOI22_X1 U8727 ( .A1(n10222), .A2(n7002), .B1(n7049), .B2(n9565), .ZN(n6975)
         );
  XNOR2_X1 U8728 ( .A(n6977), .B(n6975), .ZN(n9243) );
  INV_X1 U8729 ( .A(n6975), .ZN(n6976) );
  OR2_X1 U8730 ( .A1(n6977), .A2(n6976), .ZN(n6978) );
  AOI22_X1 U8731 ( .A1(n9955), .A2(n7045), .B1(n7002), .B2(n9929), .ZN(n6979)
         );
  AOI22_X1 U8732 ( .A1(n9955), .A2(n7002), .B1(n7049), .B2(n9929), .ZN(n8826)
         );
  AOI22_X1 U8733 ( .A1(n10271), .A2(n7045), .B1(n7002), .B2(n9928), .ZN(n6980)
         );
  XOR2_X1 U8734 ( .A(n7043), .B(n6980), .Z(n6982) );
  INV_X1 U8735 ( .A(n10271), .ZN(n9909) );
  OAI22_X1 U8736 ( .A1(n9909), .A2(n7070), .B1(n9894), .B2(n7076), .ZN(n6981)
         );
  NOR2_X1 U8737 ( .A1(n6982), .A2(n6981), .ZN(n6986) );
  AOI21_X1 U8738 ( .B1(n6982), .B2(n6981), .A(n6986), .ZN(n8892) );
  INV_X1 U8739 ( .A(n6983), .ZN(n8889) );
  INV_X1 U8740 ( .A(n9298), .ZN(n6984) );
  NAND2_X1 U8741 ( .A1(n6985), .A2(n5084), .ZN(n8893) );
  INV_X1 U8742 ( .A(n6986), .ZN(n6987) );
  NAND2_X1 U8743 ( .A1(n10197), .A2(n7045), .ZN(n6989) );
  NAND2_X1 U8744 ( .A1(n9914), .A2(n7002), .ZN(n6988) );
  NAND2_X1 U8745 ( .A1(n6989), .A2(n6988), .ZN(n6990) );
  XNOR2_X1 U8746 ( .A(n6990), .B(n7043), .ZN(n6991) );
  AOI22_X1 U8747 ( .A1(n10197), .A2(n7002), .B1(n7049), .B2(n9914), .ZN(n6992)
         );
  XNOR2_X1 U8748 ( .A(n6991), .B(n6992), .ZN(n9189) );
  INV_X1 U8749 ( .A(n6991), .ZN(n6993) );
  NAND2_X1 U8750 ( .A1(n6993), .A2(n6992), .ZN(n6994) );
  NAND2_X1 U8751 ( .A1(n9881), .A2(n7045), .ZN(n6996) );
  NAND2_X1 U8752 ( .A1(n9860), .A2(n7002), .ZN(n6995) );
  NAND2_X1 U8753 ( .A1(n6996), .A2(n6995), .ZN(n6997) );
  XNOR2_X1 U8754 ( .A(n6997), .B(n7043), .ZN(n7001) );
  NAND2_X1 U8755 ( .A1(n9881), .A2(n7002), .ZN(n6999) );
  NAND2_X1 U8756 ( .A1(n9860), .A2(n7049), .ZN(n6998) );
  NAND2_X1 U8757 ( .A1(n6999), .A2(n6998), .ZN(n7000) );
  NOR2_X1 U8758 ( .A1(n7001), .A2(n7000), .ZN(n9273) );
  NAND2_X1 U8759 ( .A1(n7001), .A2(n7000), .ZN(n9271) );
  NAND2_X1 U8760 ( .A1(n9864), .A2(n7002), .ZN(n7004) );
  NAND2_X1 U8761 ( .A1(n9845), .A2(n7049), .ZN(n7003) );
  NAND2_X1 U8762 ( .A1(n9864), .A2(n7045), .ZN(n7006) );
  NAND2_X1 U8763 ( .A1(n9845), .A2(n7002), .ZN(n7005) );
  NAND2_X1 U8764 ( .A1(n7006), .A2(n7005), .ZN(n7007) );
  XNOR2_X1 U8765 ( .A(n7007), .B(n7073), .ZN(n8866) );
  OAI22_X1 U8766 ( .A1(n9853), .A2(n6897), .B1(n8876), .B2(n7070), .ZN(n7008)
         );
  XNOR2_X1 U8767 ( .A(n7008), .B(n7043), .ZN(n7010) );
  OAI22_X1 U8768 ( .A1(n9853), .A2(n7070), .B1(n8876), .B2(n7076), .ZN(n7009)
         );
  NAND2_X1 U8769 ( .A1(n7010), .A2(n7009), .ZN(n8870) );
  OAI21_X1 U8770 ( .B1(n8868), .B2(n8866), .A(n8870), .ZN(n7012) );
  NAND3_X1 U8771 ( .A1(n8870), .A2(n8868), .A3(n8866), .ZN(n7011) );
  OR2_X1 U8772 ( .A1(n7010), .A2(n7009), .ZN(n8871) );
  NAND2_X1 U8773 ( .A1(n10256), .A2(n7045), .ZN(n7014) );
  NAND2_X1 U8774 ( .A1(n9846), .A2(n7002), .ZN(n7013) );
  NAND2_X1 U8775 ( .A1(n7014), .A2(n7013), .ZN(n7015) );
  XNOR2_X1 U8776 ( .A(n7015), .B(n7043), .ZN(n7017) );
  AND2_X1 U8777 ( .A1(n9846), .A2(n7049), .ZN(n7016) );
  AOI21_X1 U8778 ( .B1(n10256), .B2(n7002), .A(n7016), .ZN(n7018) );
  XNOR2_X1 U8779 ( .A(n7017), .B(n7018), .ZN(n8872) );
  INV_X1 U8780 ( .A(n7017), .ZN(n7019) );
  NAND2_X1 U8781 ( .A1(n7019), .A2(n7018), .ZN(n7020) );
  NAND2_X1 U8782 ( .A1(n9808), .A2(n7045), .ZN(n7022) );
  NAND2_X1 U8783 ( .A1(n9826), .A2(n7002), .ZN(n7021) );
  NAND2_X1 U8784 ( .A1(n7022), .A2(n7021), .ZN(n7023) );
  XNOR2_X1 U8785 ( .A(n7023), .B(n7043), .ZN(n8834) );
  NAND2_X1 U8786 ( .A1(n9808), .A2(n7002), .ZN(n7025) );
  NAND2_X1 U8787 ( .A1(n9826), .A2(n7049), .ZN(n7024) );
  NAND2_X1 U8788 ( .A1(n7025), .A2(n7024), .ZN(n9252) );
  AOI22_X1 U8789 ( .A1(n9787), .A2(n7045), .B1(n7002), .B2(n9803), .ZN(n7026)
         );
  XNOR2_X1 U8790 ( .A(n7026), .B(n7043), .ZN(n7028) );
  AOI22_X1 U8791 ( .A1(n9787), .A2(n7002), .B1(n7049), .B2(n9803), .ZN(n7027)
         );
  NAND2_X1 U8792 ( .A1(n7028), .A2(n7027), .ZN(n9197) );
  OAI21_X1 U8793 ( .B1(n7028), .B2(n7027), .A(n9197), .ZN(n8836) );
  AOI21_X1 U8794 ( .B1(n8834), .B2(n9252), .A(n8836), .ZN(n7029) );
  NAND2_X1 U8795 ( .A1(n8840), .A2(n9197), .ZN(n7039) );
  NAND2_X1 U8796 ( .A1(n9767), .A2(n7045), .ZN(n7031) );
  NAND2_X1 U8797 ( .A1(n9781), .A2(n7002), .ZN(n7030) );
  NAND2_X1 U8798 ( .A1(n7031), .A2(n7030), .ZN(n7032) );
  XNOR2_X1 U8799 ( .A(n7032), .B(n7073), .ZN(n7034) );
  AND2_X1 U8800 ( .A1(n9781), .A2(n7049), .ZN(n7033) );
  AOI21_X1 U8801 ( .B1(n9767), .B2(n7002), .A(n7033), .ZN(n7035) );
  NAND2_X1 U8802 ( .A1(n7034), .A2(n7035), .ZN(n7040) );
  INV_X1 U8803 ( .A(n7034), .ZN(n7037) );
  INV_X1 U8804 ( .A(n7035), .ZN(n7036) );
  NAND2_X1 U8805 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  NAND2_X1 U8806 ( .A1(n7039), .A2(n9198), .ZN(n9200) );
  NAND2_X1 U8807 ( .A1(n10153), .A2(n7045), .ZN(n7042) );
  NAND2_X1 U8808 ( .A1(n9762), .A2(n7002), .ZN(n7041) );
  NAND2_X1 U8809 ( .A1(n7042), .A2(n7041), .ZN(n7044) );
  XNOR2_X1 U8810 ( .A(n7044), .B(n7043), .ZN(n7053) );
  AOI22_X1 U8811 ( .A1(n10153), .A2(n7002), .B1(n7049), .B2(n9762), .ZN(n7051)
         );
  XNOR2_X1 U8812 ( .A(n7053), .B(n7051), .ZN(n8883) );
  NAND2_X1 U8813 ( .A1(n9735), .A2(n7045), .ZN(n7047) );
  NAND2_X1 U8814 ( .A1(n9746), .A2(n7002), .ZN(n7046) );
  NAND2_X1 U8815 ( .A1(n7047), .A2(n7046), .ZN(n7048) );
  XNOR2_X1 U8816 ( .A(n7048), .B(n7073), .ZN(n7063) );
  AND2_X1 U8817 ( .A1(n9746), .A2(n7049), .ZN(n7050) );
  AOI21_X1 U8818 ( .B1(n9735), .B2(n7002), .A(n7050), .ZN(n7064) );
  XNOR2_X1 U8819 ( .A(n7063), .B(n7064), .ZN(n9284) );
  INV_X1 U8820 ( .A(n7051), .ZN(n7052) );
  NOR2_X1 U8821 ( .A1(n7053), .A2(n7052), .ZN(n9282) );
  NOR2_X1 U8822 ( .A1(n9284), .A2(n9282), .ZN(n7054) );
  NAND2_X1 U8823 ( .A1(n8821), .A2(n7045), .ZN(n7056) );
  OR2_X1 U8824 ( .A1(n7104), .A2(n7070), .ZN(n7055) );
  NAND2_X1 U8825 ( .A1(n7056), .A2(n7055), .ZN(n7057) );
  XNOR2_X1 U8826 ( .A(n7057), .B(n7073), .ZN(n7060) );
  INV_X1 U8827 ( .A(n7060), .ZN(n7062) );
  NOR2_X1 U8828 ( .A1(n7104), .A2(n7076), .ZN(n7058) );
  AOI21_X1 U8829 ( .B1(n8821), .B2(n7002), .A(n7058), .ZN(n7059) );
  INV_X1 U8830 ( .A(n7059), .ZN(n7061) );
  AOI21_X1 U8831 ( .B1(n7062), .B2(n7061), .A(n7085), .ZN(n8814) );
  INV_X1 U8832 ( .A(n8814), .ZN(n7068) );
  INV_X1 U8833 ( .A(n7063), .ZN(n7066) );
  INV_X1 U8834 ( .A(n7064), .ZN(n7065) );
  NAND2_X1 U8835 ( .A1(n7066), .A2(n7065), .ZN(n8815) );
  INV_X1 U8836 ( .A(n8815), .ZN(n7067) );
  NOR2_X1 U8837 ( .A1(n7068), .A2(n7067), .ZN(n7069) );
  NAND2_X1 U8838 ( .A1(n7106), .A2(n7045), .ZN(n7072) );
  OR2_X1 U8839 ( .A1(n8818), .A2(n7070), .ZN(n7071) );
  NAND2_X1 U8840 ( .A1(n7072), .A2(n7071), .ZN(n7074) );
  XNOR2_X1 U8841 ( .A(n7074), .B(n7073), .ZN(n7078) );
  NAND2_X1 U8842 ( .A1(n7106), .A2(n7002), .ZN(n7075) );
  OAI21_X1 U8843 ( .B1(n8818), .B2(n7076), .A(n7075), .ZN(n7077) );
  XNOR2_X1 U8844 ( .A(n7078), .B(n7077), .ZN(n7086) );
  INV_X1 U8845 ( .A(n7079), .ZN(n7081) );
  NOR2_X1 U8846 ( .A1(n7081), .A2(n7080), .ZN(n8011) );
  INV_X1 U8847 ( .A(n7082), .ZN(n7083) );
  NAND2_X1 U8848 ( .A1(n8011), .A2(n7083), .ZN(n7099) );
  OR2_X1 U8849 ( .A1(n10228), .A2(n9472), .ZN(n7092) );
  NAND3_X1 U8850 ( .A1(n7086), .A2(n7085), .A3(n9287), .ZN(n7108) );
  NAND2_X1 U8851 ( .A1(n10133), .A2(n7087), .ZN(n8020) );
  OR3_X1 U8852 ( .A1(n7099), .A2(n7190), .A3(n8020), .ZN(n7089) );
  NOR2_X1 U8853 ( .A1(n7190), .A2(n10131), .ZN(n9554) );
  INV_X1 U8854 ( .A(n9554), .ZN(n7090) );
  OR2_X1 U8855 ( .A1(n7099), .A2(n7090), .ZN(n7091) );
  AOI22_X1 U8856 ( .A1(n9289), .A2(n9563), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n7103) );
  INV_X1 U8857 ( .A(n7092), .ZN(n7093) );
  NAND2_X1 U8858 ( .A1(n7099), .A2(n7093), .ZN(n7096) );
  NAND2_X1 U8859 ( .A1(n9548), .A2(n7175), .ZN(n7094) );
  NOR2_X1 U8860 ( .A1(n4488), .A2(n7094), .ZN(n7095) );
  AOI21_X1 U8861 ( .B1(n7096), .B2(n7095), .A(P1_U3086), .ZN(n7101) );
  NOR2_X1 U8862 ( .A1(n8020), .A2(P1_U3086), .ZN(n7097) );
  OR2_X1 U8863 ( .A1(n9554), .A2(n7097), .ZN(n7098) );
  AND2_X1 U8864 ( .A1(n7099), .A2(n7098), .ZN(n7100) );
  NAND2_X1 U8865 ( .A1(n9305), .A2(n8081), .ZN(n7102) );
  OAI211_X1 U8866 ( .C1(n7104), .C2(n9277), .A(n7103), .B(n7102), .ZN(n7105)
         );
  AOI21_X1 U8867 ( .B1(n7106), .B2(n9256), .A(n7105), .ZN(n7107) );
  NAND2_X1 U8868 ( .A1(n7108), .A2(n7107), .ZN(n7109) );
  NAND2_X1 U8869 ( .A1(n7112), .A2(n7111), .ZN(P1_U3220) );
  NAND2_X1 U8870 ( .A1(n7114), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7115) );
  NAND2_X1 U8871 ( .A1(n8821), .A2(n6140), .ZN(n7117) );
  NAND2_X1 U8872 ( .A1(n5082), .A2(n7117), .ZN(P1_U3517) );
  INV_X1 U8873 ( .A(n10508), .ZN(n7125) );
  NAND2_X1 U8874 ( .A1(n7125), .A2(n7124), .ZN(n7126) );
  NOR2_X1 U8875 ( .A1(n7175), .A2(P1_U3086), .ZN(n7128) );
  AND2_X2 U8876 ( .A1(n7128), .A2(n9548), .ZN(P1_U3973) );
  NOR2_X1 U8877 ( .A1(n5936), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10281) );
  NAND2_X1 U8878 ( .A1(n5936), .A2(P1_U3086), .ZN(n10283) );
  OAI222_X1 U8879 ( .A1(n8105), .A2(n7129), .B1(n10283), .B2(n7151), .C1(
        P1_U3086), .C2(n9599), .ZN(P1_U3351) );
  OAI222_X1 U8880 ( .A1(n8105), .A2(n7130), .B1(n10283), .B2(n7153), .C1(
        P1_U3086), .C2(n9614), .ZN(P1_U3350) );
  OAI222_X1 U8881 ( .A1(n8105), .A2(n9094), .B1(n10283), .B2(n7158), .C1(
        P1_U3086), .C2(n7232), .ZN(P1_U3352) );
  OAI222_X1 U8882 ( .A1(n8105), .A2(n7131), .B1(n10283), .B2(n7155), .C1(
        P1_U3086), .C2(n7230), .ZN(P1_U3353) );
  NAND2_X1 U8883 ( .A1(n7132), .A2(P2_U3151), .ZN(n7691) );
  AND2_X1 U8884 ( .A1(n5936), .A2(P2_U3151), .ZN(n8809) );
  INV_X1 U8885 ( .A(n8809), .ZN(n8804) );
  OAI222_X1 U8886 ( .A1(n7386), .A2(P2_U3151), .B1(n7691), .B2(n7172), .C1(
        n7133), .C2(n8804), .ZN(P2_U3294) );
  INV_X1 U8887 ( .A(n7134), .ZN(n7137) );
  OAI222_X1 U8888 ( .A1(n8105), .A2(n7135), .B1(n10283), .B2(n7137), .C1(
        P1_U3086), .C2(n9642), .ZN(P1_U3348) );
  INV_X1 U8889 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7138) );
  OAI222_X1 U8890 ( .A1(n8804), .A2(n7138), .B1(n7691), .B2(n7137), .C1(
        P2_U3151), .C2(n7136), .ZN(P2_U3288) );
  INV_X1 U8891 ( .A(n7139), .ZN(n7169) );
  OAI222_X1 U8892 ( .A1(n8804), .A2(n7141), .B1(n7691), .B2(n7169), .C1(
        P2_U3151), .C2(n7140), .ZN(P2_U3287) );
  INV_X1 U8893 ( .A(n7142), .ZN(n7150) );
  OAI222_X1 U8894 ( .A1(n8105), .A2(n7143), .B1(n10283), .B2(n7150), .C1(
        P1_U3086), .C2(n9628), .ZN(P1_U3349) );
  INV_X1 U8895 ( .A(n7144), .ZN(n7147) );
  AOI22_X1 U8896 ( .A1(n7259), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10281), .ZN(n7145) );
  OAI21_X1 U8897 ( .B1(n7147), .B2(n10283), .A(n7145), .ZN(P1_U3346) );
  OAI222_X1 U8898 ( .A1(n8804), .A2(n7148), .B1(n7691), .B2(n7147), .C1(n7146), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  CLKBUF_X1 U8899 ( .A(n7691), .Z(n8811) );
  OAI222_X1 U8900 ( .A1(n8804), .A2(n4569), .B1(n8811), .B2(n7150), .C1(
        P2_U3151), .C2(n7149), .ZN(P2_U3289) );
  OAI222_X1 U8901 ( .A1(n8804), .A2(n4531), .B1(n8811), .B2(n7151), .C1(
        P2_U3151), .C2(n7615), .ZN(P2_U3291) );
  OAI222_X1 U8902 ( .A1(n8804), .A2(n7154), .B1(n8811), .B2(n7153), .C1(
        P2_U3151), .C2(n7152), .ZN(P2_U3290) );
  OAI222_X1 U8903 ( .A1(n8804), .A2(n7156), .B1(n8811), .B2(n7155), .C1(
        P2_U3151), .C2(n6567), .ZN(P2_U3293) );
  OAI222_X1 U8904 ( .A1(n8804), .A2(n7159), .B1(n8811), .B2(n7158), .C1(
        P2_U3151), .C2(n7157), .ZN(P2_U3292) );
  NOR2_X1 U8905 ( .A1(n7193), .A2(n8968), .ZN(P2_U3252) );
  INV_X1 U8906 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n8955) );
  NOR2_X1 U8907 ( .A1(n7193), .A2(n8955), .ZN(P2_U3246) );
  INV_X1 U8908 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9177) );
  NOR2_X1 U8909 ( .A1(n7193), .A2(n9177), .ZN(P2_U3263) );
  NOR2_X1 U8910 ( .A1(n7193), .A2(n9026), .ZN(P2_U3256) );
  INV_X1 U8911 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9178) );
  NOR2_X1 U8912 ( .A1(n7193), .A2(n9178), .ZN(P2_U3251) );
  INV_X1 U8913 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n8918) );
  NOR2_X1 U8914 ( .A1(n7193), .A2(n8918), .ZN(P2_U3250) );
  NOR2_X1 U8915 ( .A1(n7193), .A2(n8915), .ZN(P2_U3244) );
  NOR2_X1 U8916 ( .A1(n7193), .A2(n8967), .ZN(P2_U3243) );
  INV_X1 U8917 ( .A(n7161), .ZN(n7164) );
  OAI222_X1 U8918 ( .A1(n8804), .A2(n7162), .B1(n7691), .B2(n7164), .C1(n7737), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U8919 ( .A(n10283), .ZN(n7789) );
  INV_X1 U8920 ( .A(n7789), .ZN(n8004) );
  AOI22_X1 U8921 ( .A1(n7313), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10281), .ZN(n7163) );
  OAI21_X1 U8922 ( .B1(n7164), .B2(n8004), .A(n7163), .ZN(P1_U3345) );
  INV_X1 U8923 ( .A(n7165), .ZN(n7168) );
  AOI22_X1 U8924 ( .A1(n7914), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8809), .ZN(n7166) );
  OAI21_X1 U8925 ( .B1(n7168), .B2(n8811), .A(n7166), .ZN(P2_U3284) );
  AOI22_X1 U8926 ( .A1(n9678), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10281), .ZN(n7167) );
  OAI21_X1 U8927 ( .B1(n7168), .B2(n10283), .A(n7167), .ZN(P1_U3344) );
  OAI222_X1 U8928 ( .A1(n8105), .A2(n7170), .B1(n8004), .B2(n7169), .C1(
        P1_U3086), .C2(n7241), .ZN(P1_U3347) );
  NAND2_X1 U8929 ( .A1(n9472), .A2(n9548), .ZN(n7174) );
  AND2_X1 U8930 ( .A1(n7174), .A2(n7173), .ZN(n7180) );
  INV_X1 U8931 ( .A(n7180), .ZN(n7177) );
  INV_X1 U8932 ( .A(n7175), .ZN(n7176) );
  AOI21_X1 U8933 ( .B1(n7176), .B2(n9548), .A(P1_U3086), .ZN(n7181) );
  INV_X1 U8934 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7184) );
  OAI21_X1 U8935 ( .B1(n7989), .B2(P1_REG2_REG_0__SCAN_IN), .A(n7280), .ZN(
        n7282) );
  AOI21_X1 U8936 ( .B1(n7989), .B2(n7178), .A(n7282), .ZN(n7179) );
  XNOR2_X1 U8937 ( .A(n7179), .B(n4744), .ZN(n7182) );
  AOI22_X1 U8938 ( .A1(n7182), .A2(n7245), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n7183) );
  OAI21_X1 U8939 ( .B1(n10332), .B2(n7184), .A(n7183), .ZN(P1_U3243) );
  INV_X1 U8940 ( .A(n10332), .ZN(n9699) );
  NOR2_X1 U8941 ( .A1(n9699), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8942 ( .A(n7185), .ZN(n7187) );
  OAI222_X1 U8943 ( .A1(n8105), .A2(n7186), .B1(n8004), .B2(n7187), .C1(n7597), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  OAI222_X1 U8944 ( .A1(n8804), .A2(n7188), .B1(n7691), .B2(n7187), .C1(n7928), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U8945 ( .A(n10381), .ZN(n10380) );
  INV_X1 U8946 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U8947 ( .A1(n10380), .A2(n7191), .ZN(n7192) );
  OAI21_X1 U8948 ( .B1(n10380), .B2(n8924), .A(n7192), .ZN(P1_U3440) );
  AND2_X1 U8949 ( .A1(n7198), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8950 ( .A1(n7198), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8951 ( .A1(n7198), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8952 ( .A1(n7198), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8953 ( .A1(n7198), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8954 ( .A1(n7198), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8955 ( .A1(n7198), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8956 ( .A1(n7198), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8957 ( .A1(n7198), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8958 ( .A1(n7198), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8959 ( .A1(n7198), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8960 ( .A1(n7198), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8961 ( .A1(n7198), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8962 ( .A1(n7198), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8963 ( .A1(n7198), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8964 ( .A1(n7198), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8965 ( .A1(n7198), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8966 ( .A1(n7198), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8967 ( .A1(n7198), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8968 ( .A1(n7198), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8969 ( .A1(n7198), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8970 ( .A1(n7198), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8971 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7197) );
  INV_X1 U8972 ( .A(n7194), .ZN(n7196) );
  AOI22_X1 U8973 ( .A1(n7198), .A2(n7197), .B1(n7196), .B2(n7195), .ZN(
        P2_U3376) );
  INV_X1 U8974 ( .A(n7199), .ZN(n7208) );
  AOI22_X1 U8975 ( .A1(n8057), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10281), .ZN(n7200) );
  OAI21_X1 U8976 ( .B1(n7208), .B2(n10283), .A(n7200), .ZN(P1_U3342) );
  NAND2_X1 U8977 ( .A1(n7481), .A2(P1_U3973), .ZN(n7201) );
  OAI21_X1 U8978 ( .B1(P1_U3973), .B2(n5094), .A(n7201), .ZN(P1_U3554) );
  INV_X1 U8979 ( .A(P1_U3973), .ZN(n7203) );
  NAND2_X1 U8980 ( .A1(n7203), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7202) );
  OAI21_X1 U8981 ( .B1(n9447), .B2(n7203), .A(n7202), .ZN(P1_U3584) );
  INV_X1 U8982 ( .A(n7204), .ZN(n7207) );
  OAI222_X1 U8983 ( .A1(n8804), .A2(n7205), .B1(n7691), .B2(n7207), .C1(
        P2_U3151), .C2(n8331), .ZN(P2_U3281) );
  INV_X1 U8984 ( .A(n10293), .ZN(n7206) );
  OAI222_X1 U8985 ( .A1(n8105), .A2(n9171), .B1(n8004), .B2(n7207), .C1(
        P1_U3086), .C2(n7206), .ZN(P1_U3341) );
  OAI222_X1 U8986 ( .A1(n8804), .A2(n9141), .B1(n7691), .B2(n7208), .C1(
        P2_U3151), .C2(n4647), .ZN(P2_U3282) );
  INV_X1 U8987 ( .A(n7209), .ZN(n7210) );
  OAI222_X1 U8988 ( .A1(n8804), .A2(n9107), .B1(n7691), .B2(n7210), .C1(n8348), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  INV_X1 U8989 ( .A(n10311), .ZN(n8062) );
  OAI222_X1 U8990 ( .A1(n8105), .A2(n8944), .B1(n8004), .B2(n7210), .C1(n8062), 
        .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U8991 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10048) );
  MUX2_X1 U8992 ( .A(n10048), .B(P1_REG2_REG_9__SCAN_IN), .S(n7259), .Z(n7224)
         );
  XNOR2_X1 U8993 ( .A(n7228), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9579) );
  AND2_X1 U8994 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9578) );
  NAND2_X1 U8995 ( .A1(n9579), .A2(n9578), .ZN(n9577) );
  INV_X1 U8996 ( .A(n7228), .ZN(n9576) );
  NAND2_X1 U8997 ( .A1(n9576), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7211) );
  NAND2_X1 U8998 ( .A1(n9577), .A2(n7211), .ZN(n7288) );
  XNOR2_X1 U8999 ( .A(n7230), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n7289) );
  NAND2_X1 U9000 ( .A1(n7288), .A2(n7289), .ZN(n7287) );
  INV_X1 U9001 ( .A(n7230), .ZN(n7297) );
  NAND2_X1 U9002 ( .A1(n7297), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7212) );
  NAND2_X1 U9003 ( .A1(n7287), .A2(n7212), .ZN(n9594) );
  XNOR2_X1 U9004 ( .A(n7232), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U9005 ( .A1(n9594), .A2(n9595), .ZN(n9593) );
  INV_X1 U9006 ( .A(n7232), .ZN(n9589) );
  NAND2_X1 U9007 ( .A1(n9589), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7213) );
  NAND2_X1 U9008 ( .A1(n9593), .A2(n7213), .ZN(n9605) );
  INV_X1 U9009 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9051) );
  MUX2_X1 U9010 ( .A(n9051), .B(P1_REG2_REG_4__SCAN_IN), .S(n9599), .Z(n9606)
         );
  NAND2_X1 U9011 ( .A1(n9605), .A2(n9606), .ZN(n9604) );
  OR2_X1 U9012 ( .A1(n9599), .A2(n9051), .ZN(n7214) );
  NAND2_X1 U9013 ( .A1(n9604), .A2(n7214), .ZN(n9623) );
  XNOR2_X1 U9014 ( .A(n9614), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U9015 ( .A1(n9623), .A2(n9624), .ZN(n9622) );
  INV_X1 U9016 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7215) );
  OR2_X1 U9017 ( .A1(n9614), .A2(n7215), .ZN(n7216) );
  NAND2_X1 U9018 ( .A1(n9622), .A2(n7216), .ZN(n9634) );
  XNOR2_X1 U9019 ( .A(n9628), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U9020 ( .A1(n9634), .A2(n9635), .ZN(n9633) );
  INV_X1 U9021 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7217) );
  OR2_X1 U9022 ( .A1(n9628), .A2(n7217), .ZN(n7218) );
  NAND2_X1 U9023 ( .A1(n9633), .A2(n7218), .ZN(n9648) );
  XNOR2_X1 U9024 ( .A(n9642), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U9025 ( .A1(n9648), .A2(n9649), .ZN(n9647) );
  INV_X1 U9026 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7219) );
  OR2_X1 U9027 ( .A1(n9642), .A2(n7219), .ZN(n7220) );
  NAND2_X1 U9028 ( .A1(n9647), .A2(n7220), .ZN(n9664) );
  XNOR2_X1 U9029 ( .A(n7241), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n9665) );
  NAND2_X1 U9030 ( .A1(n9664), .A2(n9665), .ZN(n9663) );
  INV_X1 U9031 ( .A(n7241), .ZN(n9659) );
  NAND2_X1 U9032 ( .A1(n9659), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7221) );
  NAND2_X1 U9033 ( .A1(n9663), .A2(n7221), .ZN(n7223) );
  INV_X1 U9034 ( .A(n7261), .ZN(n7222) );
  AOI21_X1 U9035 ( .B1(n7224), .B2(n7223), .A(n7222), .ZN(n7250) );
  NOR2_X1 U9036 ( .A1(n6095), .A2(n7989), .ZN(n9553) );
  NAND2_X1 U9037 ( .A1(n7245), .A2(n9553), .ZN(n10316) );
  INV_X1 U9038 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7227) );
  NOR2_X1 U9039 ( .A1(n7225), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9226) );
  INV_X1 U9040 ( .A(n9226), .ZN(n7226) );
  OAI21_X1 U9041 ( .B1(n10332), .B2(n7227), .A(n7226), .ZN(n7248) );
  XNOR2_X1 U9042 ( .A(n7228), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9582) );
  AND2_X1 U9043 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9581) );
  NAND2_X1 U9044 ( .A1(n9582), .A2(n9581), .ZN(n9580) );
  NAND2_X1 U9045 ( .A1(n9576), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7229) );
  NAND2_X1 U9046 ( .A1(n9580), .A2(n7229), .ZN(n7291) );
  XNOR2_X1 U9047 ( .A(n7230), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U9048 ( .A1(n7291), .A2(n7292), .ZN(n7290) );
  NAND2_X1 U9049 ( .A1(n7297), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7231) );
  NAND2_X1 U9050 ( .A1(n7290), .A2(n7231), .ZN(n9591) );
  XNOR2_X1 U9051 ( .A(n7232), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9592) );
  NAND2_X1 U9052 ( .A1(n9591), .A2(n9592), .ZN(n9590) );
  NAND2_X1 U9053 ( .A1(n9589), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7233) );
  NAND2_X1 U9054 ( .A1(n9590), .A2(n7233), .ZN(n9608) );
  INV_X1 U9055 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9168) );
  MUX2_X1 U9056 ( .A(n9168), .B(P1_REG1_REG_4__SCAN_IN), .S(n9599), .Z(n9609)
         );
  NAND2_X1 U9057 ( .A1(n9608), .A2(n9609), .ZN(n9607) );
  OR2_X1 U9058 ( .A1(n9599), .A2(n9168), .ZN(n7234) );
  NAND2_X1 U9059 ( .A1(n9607), .A2(n7234), .ZN(n9620) );
  XNOR2_X1 U9060 ( .A(n9614), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U9061 ( .A1(n9620), .A2(n9621), .ZN(n9619) );
  INV_X1 U9062 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7235) );
  OR2_X1 U9063 ( .A1(n9614), .A2(n7235), .ZN(n7236) );
  NAND2_X1 U9064 ( .A1(n9619), .A2(n7236), .ZN(n9637) );
  XNOR2_X1 U9065 ( .A(n9628), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U9066 ( .A1(n9637), .A2(n9638), .ZN(n9636) );
  INV_X1 U9067 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7237) );
  OR2_X1 U9068 ( .A1(n9628), .A2(n7237), .ZN(n7238) );
  NAND2_X1 U9069 ( .A1(n9636), .A2(n7238), .ZN(n9651) );
  XNOR2_X1 U9070 ( .A(n9642), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n9652) );
  NAND2_X1 U9071 ( .A1(n9651), .A2(n9652), .ZN(n9650) );
  INV_X1 U9072 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7239) );
  OR2_X1 U9073 ( .A1(n9642), .A2(n7239), .ZN(n7240) );
  NAND2_X1 U9074 ( .A1(n9650), .A2(n7240), .ZN(n9661) );
  INV_X1 U9075 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10436) );
  MUX2_X1 U9076 ( .A(n10436), .B(P1_REG1_REG_8__SCAN_IN), .S(n7241), .Z(n9662)
         );
  NAND2_X1 U9077 ( .A1(n9661), .A2(n9662), .ZN(n9660) );
  NAND2_X1 U9078 ( .A1(n9659), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7242) );
  NAND2_X1 U9079 ( .A1(n9660), .A2(n7242), .ZN(n7244) );
  INV_X1 U9080 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10438) );
  MUX2_X1 U9081 ( .A(n10438), .B(P1_REG1_REG_9__SCAN_IN), .S(n7259), .Z(n7243)
         );
  NAND2_X1 U9082 ( .A1(n7244), .A2(n7243), .ZN(n7246) );
  NAND2_X1 U9083 ( .A1(n7245), .A2(n7989), .ZN(n10302) );
  AOI21_X1 U9084 ( .B1(n7255), .B2(n7246), .A(n10302), .ZN(n7247) );
  AOI211_X1 U9085 ( .C1(n10312), .C2(n7259), .A(n7248), .B(n7247), .ZN(n7249)
         );
  OAI21_X1 U9086 ( .B1(n7250), .B2(n10316), .A(n7249), .ZN(P1_U3252) );
  NOR2_X1 U9087 ( .A1(n8290), .A2(P2_U3151), .ZN(n7338) );
  AOI22_X1 U9088 ( .A1(n8271), .A2(n10467), .B1(n8258), .B2(n8304), .ZN(n7252)
         );
  NAND2_X1 U9089 ( .A1(n8263), .A2(n10472), .ZN(n7251) );
  OAI211_X1 U9090 ( .C1(n7338), .C2(n5283), .A(n7252), .B(n7251), .ZN(P2_U3172) );
  INV_X1 U9091 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7253) );
  MUX2_X1 U9092 ( .A(n7253), .B(P1_REG1_REG_10__SCAN_IN), .S(n7313), .Z(n7258)
         );
  OR2_X1 U9093 ( .A1(n7259), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7254) );
  NAND2_X1 U9094 ( .A1(n7255), .A2(n7254), .ZN(n7257) );
  INV_X1 U9095 ( .A(n7315), .ZN(n7256) );
  AOI211_X1 U9096 ( .C1(n7258), .C2(n7257), .A(n10302), .B(n7256), .ZN(n7269)
         );
  XNOR2_X1 U9097 ( .A(n7313), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7264) );
  OR2_X1 U9098 ( .A1(n7259), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7260) );
  NAND2_X1 U9099 ( .A1(n7261), .A2(n7260), .ZN(n7263) );
  INV_X1 U9100 ( .A(n7304), .ZN(n7262) );
  AOI211_X1 U9101 ( .C1(n7264), .C2(n7263), .A(n10316), .B(n7262), .ZN(n7268)
         );
  INV_X1 U9102 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7266) );
  NAND2_X1 U9103 ( .A1(n10312), .A2(n7313), .ZN(n7265) );
  NAND2_X1 U9104 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8851) );
  OAI211_X1 U9105 ( .C1(n7266), .C2(n10332), .A(n7265), .B(n8851), .ZN(n7267)
         );
  OR3_X1 U9106 ( .A1(n7269), .A2(n7268), .A3(n7267), .ZN(P1_U3253) );
  INV_X1 U9107 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9106) );
  INV_X1 U9108 ( .A(n7270), .ZN(n7271) );
  INV_X1 U9109 ( .A(n8064), .ZN(n9687) );
  OAI222_X1 U9110 ( .A1(n8105), .A2(n9106), .B1(n8004), .B2(n7271), .C1(
        P1_U3086), .C2(n9687), .ZN(P1_U3339) );
  INV_X1 U9111 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7272) );
  OAI222_X1 U9112 ( .A1(n8804), .A2(n7272), .B1(n7691), .B2(n7271), .C1(
        P2_U3151), .C2(n8360), .ZN(P2_U3279) );
  XNOR2_X1 U9113 ( .A(n7274), .B(n7273), .ZN(n7281) );
  NAND2_X1 U9114 ( .A1(n9292), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7382) );
  OAI22_X1 U9115 ( .A1(n9302), .A2(n7277), .B1(n9301), .B2(n9480), .ZN(n7275)
         );
  AOI21_X1 U9116 ( .B1(n7382), .B2(P1_REG3_REG_0__SCAN_IN), .A(n7275), .ZN(
        n7276) );
  OAI21_X1 U9117 ( .B1(n9307), .B2(n7281), .A(n7276), .ZN(P1_U3232) );
  NOR2_X1 U9118 ( .A1(n9480), .A2(n6461), .ZN(n10136) );
  NAND2_X1 U9119 ( .A1(n7481), .A2(n7277), .ZN(n9481) );
  AND2_X1 U9120 ( .A1(n7479), .A2(n9481), .ZN(n10134) );
  AOI21_X1 U9121 ( .B1(n6464), .B2(n10225), .A(n10134), .ZN(n7278) );
  AOI211_X1 U9122 ( .C1(n10137), .C2(n10133), .A(n10136), .B(n7278), .ZN(
        n10382) );
  NAND2_X1 U9123 ( .A1(n10440), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7279) );
  OAI21_X1 U9124 ( .B1(n10382), .B2(n10440), .A(n7279), .ZN(P1_U3522) );
  NAND3_X1 U9125 ( .A1(n7281), .A2(n7280), .A3(n7989), .ZN(n7284) );
  AOI22_X1 U9126 ( .A1(n4744), .A2(n7282), .B1(n9553), .B2(n9578), .ZN(n7283)
         );
  NAND3_X1 U9127 ( .A1(n7284), .A2(P1_U3973), .A3(n7283), .ZN(n9613) );
  INV_X1 U9128 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7286) );
  INV_X1 U9129 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7285) );
  OAI22_X1 U9130 ( .A1(n10332), .A2(n7286), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7285), .ZN(n7296) );
  OAI21_X1 U9131 ( .B1(n7289), .B2(n7288), .A(n7287), .ZN(n7294) );
  OAI21_X1 U9132 ( .B1(n7292), .B2(n7291), .A(n7290), .ZN(n7293) );
  OAI22_X1 U9133 ( .A1(n10316), .A2(n7294), .B1(n10302), .B2(n7293), .ZN(n7295) );
  AOI211_X1 U9134 ( .C1(n7297), .C2(n10312), .A(n7296), .B(n7295), .ZN(n7298)
         );
  NAND2_X1 U9135 ( .A1(n9613), .A2(n7298), .ZN(P1_U3245) );
  INV_X1 U9136 ( .A(n7299), .ZN(n7301) );
  OAI222_X1 U9137 ( .A1(n8804), .A2(n7300), .B1(n7691), .B2(n7301), .C1(
        P2_U3151), .C2(n8378), .ZN(P2_U3278) );
  INV_X1 U9138 ( .A(n8066), .ZN(n9702) );
  OAI222_X1 U9139 ( .A1(n8105), .A2(n7302), .B1(n8004), .B2(n7301), .C1(
        P1_U3086), .C2(n9702), .ZN(P1_U3338) );
  INV_X1 U9140 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7596) );
  XNOR2_X1 U9141 ( .A(n7597), .B(n7596), .ZN(n7309) );
  NAND2_X1 U9142 ( .A1(n7313), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7303) );
  NAND2_X1 U9143 ( .A1(n7304), .A2(n7303), .ZN(n9674) );
  INV_X1 U9144 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7305) );
  XNOR2_X1 U9145 ( .A(n9678), .B(n7305), .ZN(n9673) );
  NAND2_X1 U9146 ( .A1(n9674), .A2(n9673), .ZN(n9672) );
  NAND2_X1 U9147 ( .A1(n9678), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7306) );
  NAND2_X1 U9148 ( .A1(n9672), .A2(n7306), .ZN(n7308) );
  INV_X1 U9149 ( .A(n7599), .ZN(n7307) );
  AOI21_X1 U9150 ( .B1(n7309), .B2(n7308), .A(n7307), .ZN(n7325) );
  INV_X1 U9151 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7312) );
  NOR2_X1 U9152 ( .A1(n7310), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7983) );
  INV_X1 U9153 ( .A(n7983), .ZN(n7311) );
  OAI21_X1 U9154 ( .B1(n10332), .B2(n7312), .A(n7311), .ZN(n7322) );
  NAND2_X1 U9155 ( .A1(n7313), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7314) );
  NAND2_X1 U9156 ( .A1(n7315), .A2(n7314), .ZN(n9671) );
  INV_X1 U9157 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7316) );
  XNOR2_X1 U9158 ( .A(n9678), .B(n7316), .ZN(n9670) );
  NAND2_X1 U9159 ( .A1(n9671), .A2(n9670), .ZN(n9669) );
  NAND2_X1 U9160 ( .A1(n9678), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7317) );
  NAND2_X1 U9161 ( .A1(n9669), .A2(n7317), .ZN(n7319) );
  INV_X1 U9162 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8002) );
  XNOR2_X1 U9163 ( .A(n7597), .B(n8002), .ZN(n7318) );
  NAND2_X1 U9164 ( .A1(n7319), .A2(n7318), .ZN(n7320) );
  AOI21_X1 U9165 ( .B1(n7592), .B2(n7320), .A(n10302), .ZN(n7321) );
  AOI211_X1 U9166 ( .C1(n10312), .C2(n7323), .A(n7322), .B(n7321), .ZN(n7324)
         );
  OAI21_X1 U9167 ( .B1(n7325), .B2(n10316), .A(n7324), .ZN(P1_U3255) );
  XOR2_X1 U9168 ( .A(n7327), .B(n7326), .Z(n7333) );
  OR2_X1 U9169 ( .A1(n7328), .A2(n10488), .ZN(n10456) );
  INV_X1 U9170 ( .A(n10456), .ZN(n8700) );
  OAI22_X1 U9171 ( .A1(n8274), .A2(n6150), .B1(n7329), .B2(n8288), .ZN(n7331)
         );
  NOR2_X1 U9172 ( .A1(n7338), .A2(n5299), .ZN(n7330) );
  AOI211_X1 U9173 ( .C1(n7489), .C2(n8700), .A(n7331), .B(n7330), .ZN(n7332)
         );
  OAI21_X1 U9174 ( .B1(n7333), .B2(n8281), .A(n7332), .ZN(P2_U3177) );
  XOR2_X1 U9175 ( .A(n7334), .B(n7335), .Z(n7343) );
  OR2_X1 U9176 ( .A1(n7475), .A2(n10488), .ZN(n7420) );
  INV_X1 U9177 ( .A(n7420), .ZN(n7341) );
  OAI22_X1 U9178 ( .A1(n8274), .A2(n7337), .B1(n7336), .B2(n8288), .ZN(n7340)
         );
  NOR2_X1 U9179 ( .A1(n7338), .A2(n7468), .ZN(n7339) );
  AOI211_X1 U9180 ( .C1(n7489), .C2(n7341), .A(n7340), .B(n7339), .ZN(n7342)
         );
  OAI21_X1 U9181 ( .B1(n8281), .B2(n7343), .A(n7342), .ZN(P2_U3162) );
  NOR2_X1 U9182 ( .A1(n7344), .A2(n10488), .ZN(n10480) );
  NAND2_X1 U9183 ( .A1(n7489), .A2(n10480), .ZN(n7347) );
  NOR2_X1 U9184 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7355), .ZN(n7555) );
  AOI21_X1 U9185 ( .B1(n8286), .B2(n7345), .A(n7555), .ZN(n7346) );
  OAI211_X1 U9186 ( .C1(n7348), .C2(n8288), .A(n7347), .B(n7346), .ZN(n7354)
         );
  INV_X1 U9187 ( .A(n7349), .ZN(n7350) );
  AOI211_X1 U9188 ( .C1(n7352), .C2(n7351), .A(n8281), .B(n7350), .ZN(n7353)
         );
  AOI211_X1 U9189 ( .C1(n7355), .C2(n8290), .A(n7354), .B(n7353), .ZN(n7356)
         );
  INV_X1 U9190 ( .A(n7356), .ZN(P2_U3158) );
  INV_X1 U9191 ( .A(n7382), .ZN(n7365) );
  INV_X1 U9192 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9573) );
  OAI21_X1 U9193 ( .B1(n7359), .B2(n7358), .A(n7357), .ZN(n7360) );
  NAND2_X1 U9194 ( .A1(n7360), .A2(n9287), .ZN(n7364) );
  OAI22_X1 U9195 ( .A1(n9302), .A2(n10122), .B1(n9277), .B2(n7361), .ZN(n7362)
         );
  AOI21_X1 U9196 ( .B1(n9289), .B2(n9571), .A(n7362), .ZN(n7363) );
  OAI211_X1 U9197 ( .C1(n7365), .C2(n9573), .A(n7364), .B(n7363), .ZN(P1_U3222) );
  INV_X1 U9198 ( .A(n7366), .ZN(n7367) );
  INV_X1 U9199 ( .A(n8068), .ZN(n10324) );
  OAI222_X1 U9200 ( .A1(n8105), .A2(n8948), .B1(n8004), .B2(n7367), .C1(n10324), .C2(P1_U3086), .ZN(P1_U3337) );
  OAI222_X1 U9201 ( .A1(P2_U3151), .A2(n8406), .B1(n7691), .B2(n7367), .C1(
        n9074), .C2(n8804), .ZN(P2_U3277) );
  INV_X1 U9202 ( .A(n7368), .ZN(n7544) );
  AND2_X1 U9203 ( .A1(n10473), .A2(n7545), .ZN(n10485) );
  NAND2_X1 U9204 ( .A1(n7489), .A2(n10485), .ZN(n7370) );
  AND2_X1 U9205 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7613) );
  AOI21_X1 U9206 ( .B1(n8286), .B2(n6771), .A(n7613), .ZN(n7369) );
  OAI211_X1 U9207 ( .C1(n7495), .C2(n8288), .A(n7370), .B(n7369), .ZN(n7374)
         );
  AOI21_X1 U9208 ( .B1(n7372), .B2(n7371), .A(n8281), .ZN(n7373) );
  AOI211_X1 U9209 ( .C1(n7544), .C2(n8290), .A(n7374), .B(n7373), .ZN(n7375)
         );
  INV_X1 U9210 ( .A(n7375), .ZN(P2_U3170) );
  AND3_X1 U9211 ( .A1(n7357), .A2(n7377), .A3(n7376), .ZN(n7378) );
  OAI21_X1 U9212 ( .B1(n7379), .B2(n7378), .A(n9287), .ZN(n7384) );
  AOI22_X1 U9213 ( .A1(n9299), .A2(n9572), .B1(n7518), .B2(n9256), .ZN(n7380)
         );
  OAI21_X1 U9214 ( .B1(n9214), .B2(n9301), .A(n7380), .ZN(n7381) );
  AOI21_X1 U9215 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7382), .A(n7381), .ZN(
        n7383) );
  NAND2_X1 U9216 ( .A1(n7384), .A2(n7383), .ZN(P1_U3237) );
  XNOR2_X1 U9217 ( .A(n7385), .B(n10451), .ZN(n7396) );
  OAI22_X1 U9218 ( .A1(n8401), .A2(n7386), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7468), .ZN(n7394) );
  INV_X1 U9219 ( .A(n7387), .ZN(n7388) );
  AOI21_X1 U9220 ( .B1(n7473), .B2(n7389), .A(n7388), .ZN(n7392) );
  INV_X1 U9221 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7423) );
  XNOR2_X1 U9222 ( .A(n7390), .B(n7423), .ZN(n7391) );
  OAI22_X1 U9223 ( .A1(n8389), .A2(n7392), .B1(n8411), .B2(n7391), .ZN(n7393)
         );
  AOI211_X1 U9224 ( .C1(n10443), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7394), .B(
        n7393), .ZN(n7395) );
  OAI21_X1 U9225 ( .B1(n8404), .B2(n7396), .A(n7395), .ZN(P2_U3183) );
  XNOR2_X1 U9226 ( .A(n7398), .B(n7397), .ZN(n7411) );
  XNOR2_X1 U9227 ( .A(n7399), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U9228 ( .A1(n10443), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n7407) );
  AND2_X1 U9229 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7436) );
  AOI21_X1 U9230 ( .B1(n10444), .B2(n7400), .A(n7436), .ZN(n7406) );
  NAND2_X1 U9231 ( .A1(n7402), .A2(n7401), .ZN(n7403) );
  NAND2_X1 U9232 ( .A1(n7452), .A2(n7403), .ZN(n7404) );
  NAND2_X1 U9233 ( .A1(n8396), .A2(n7404), .ZN(n7405) );
  NAND3_X1 U9234 ( .A1(n7407), .A2(n7406), .A3(n7405), .ZN(n7408) );
  AOI21_X1 U9235 ( .B1(n8385), .B2(n7409), .A(n7408), .ZN(n7410) );
  OAI21_X1 U9236 ( .B1(n8404), .B2(n7411), .A(n7410), .ZN(P2_U3187) );
  INV_X1 U9237 ( .A(n7412), .ZN(n7413) );
  NAND2_X1 U9238 ( .A1(n7414), .A2(n7416), .ZN(n7471) );
  INV_X1 U9239 ( .A(n7878), .ZN(n8689) );
  NAND2_X1 U9240 ( .A1(n7471), .A2(n8689), .ZN(n7418) );
  AOI22_X1 U9241 ( .A1(n8692), .A2(n7345), .B1(n8609), .B2(n8306), .ZN(n7417)
         );
  OAI211_X1 U9242 ( .C1(n7419), .C2(n10469), .A(n7418), .B(n7417), .ZN(n7469)
         );
  NAND2_X1 U9243 ( .A1(n7471), .A2(n10493), .ZN(n7421) );
  NAND2_X1 U9244 ( .A1(n7421), .A2(n7420), .ZN(n7422) );
  NOR2_X1 U9245 ( .A1(n7469), .A2(n7422), .ZN(n10475) );
  MUX2_X1 U9246 ( .A(n7423), .B(n10475), .S(n10508), .Z(n7424) );
  INV_X1 U9247 ( .A(n7424), .ZN(P2_U3460) );
  INV_X1 U9248 ( .A(n10463), .ZN(n7425) );
  NAND2_X1 U9249 ( .A1(n7878), .A2(n7425), .ZN(n7426) );
  XNOR2_X1 U9250 ( .A(n7427), .B(n7429), .ZN(n10477) );
  XNOR2_X1 U9251 ( .A(n7428), .B(n7429), .ZN(n7430) );
  AOI222_X1 U9252 ( .A1(n8696), .A2(n7430), .B1(n8303), .B2(n8692), .C1(n7345), 
        .C2(n8609), .ZN(n10478) );
  MUX2_X1 U9253 ( .A(n7550), .B(n10478), .S(n10464), .Z(n7433) );
  AOI22_X1 U9254 ( .A1(n8589), .A2(n7431), .B1(n7355), .B2(n8588), .ZN(n7432)
         );
  OAI211_X1 U9255 ( .C1(n8553), .C2(n10477), .A(n7433), .B(n7432), .ZN(
        P2_U3230) );
  XOR2_X1 U9256 ( .A(n7435), .B(n7434), .Z(n7442) );
  AOI21_X1 U9257 ( .B1(n8286), .B2(n8303), .A(n7436), .ZN(n7437) );
  OAI21_X1 U9258 ( .B1(n7700), .B2(n8288), .A(n7437), .ZN(n7439) );
  NOR2_X1 U9259 ( .A1(n8248), .A2(n7678), .ZN(n7438) );
  AOI211_X1 U9260 ( .C1(n8263), .C2(n7440), .A(n7439), .B(n7438), .ZN(n7441)
         );
  OAI21_X1 U9261 ( .B1(n7442), .B2(n8281), .A(n7441), .ZN(P2_U3167) );
  INV_X1 U9262 ( .A(n7642), .ZN(n7443) );
  AOI21_X1 U9263 ( .B1(n7445), .B2(n7444), .A(n7443), .ZN(n7461) );
  OAI21_X1 U9264 ( .B1(n7448), .B2(n7447), .A(n7446), .ZN(n7459) );
  INV_X1 U9265 ( .A(n7449), .ZN(n7454) );
  NAND3_X1 U9266 ( .A1(n7452), .A2(n7451), .A3(n7450), .ZN(n7453) );
  AOI21_X1 U9267 ( .B1(n7454), .B2(n7453), .A(n8389), .ZN(n7458) );
  INV_X1 U9268 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U9269 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U9270 ( .A1(n10444), .A2(n7455), .ZN(n7456) );
  OAI211_X1 U9271 ( .C1(n7916), .C2(n9146), .A(n7494), .B(n7456), .ZN(n7457)
         );
  AOI211_X1 U9272 ( .C1(n8385), .C2(n7459), .A(n7458), .B(n7457), .ZN(n7460)
         );
  OAI21_X1 U9273 ( .B1(n7461), .B2(n8404), .A(n7460), .ZN(P2_U3188) );
  AOI22_X1 U9274 ( .A1(n8589), .A2(n10472), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8588), .ZN(n7467) );
  INV_X1 U9275 ( .A(n7462), .ZN(n7463) );
  NOR2_X1 U9276 ( .A1(n7463), .A2(n10473), .ZN(n7464) );
  INV_X1 U9277 ( .A(n8692), .ZN(n8558) );
  NOR2_X1 U9278 ( .A1(n8558), .A2(n6150), .ZN(n10471) );
  AOI21_X1 U9279 ( .B1(n7464), .B2(n10467), .A(n10471), .ZN(n7465) );
  MUX2_X1 U9280 ( .A(n10447), .B(n7465), .S(n10464), .Z(n7466) );
  NAND2_X1 U9281 ( .A1(n7467), .A2(n7466), .ZN(P2_U3233) );
  NOR2_X1 U9282 ( .A1(n10458), .A2(n7468), .ZN(n7470) );
  AOI211_X1 U9283 ( .C1(n10463), .C2(n7471), .A(n7470), .B(n7469), .ZN(n7472)
         );
  MUX2_X1 U9284 ( .A(n7473), .B(n7472), .S(n10464), .Z(n7474) );
  OAI21_X1 U9285 ( .B1(n8618), .B2(n7475), .A(n7474), .ZN(P2_U3232) );
  XNOR2_X1 U9286 ( .A(n9480), .B(n10122), .ZN(n9430) );
  INV_X1 U9287 ( .A(n9430), .ZN(n7477) );
  NAND2_X1 U9288 ( .A1(n7477), .A2(n7476), .ZN(n7515) );
  INV_X1 U9289 ( .A(n7515), .ZN(n7478) );
  AOI21_X1 U9290 ( .B1(n6469), .B2(n9430), .A(n7478), .ZN(n10125) );
  INV_X1 U9291 ( .A(n7479), .ZN(n7480) );
  NAND2_X1 U9292 ( .A1(n9430), .A2(n7480), .ZN(n7519) );
  OAI21_X1 U9293 ( .B1(n7480), .B2(n9430), .A(n7519), .ZN(n7482) );
  AOI222_X1 U9294 ( .A1(n10014), .A2(n7482), .B1(n7481), .B2(n10356), .C1(
        n9571), .C2(n10017), .ZN(n10130) );
  AOI21_X1 U9295 ( .B1(n4391), .B2(n10137), .A(n10214), .ZN(n7483) );
  NAND2_X1 U9296 ( .A1(n7483), .A2(n7517), .ZN(n10120) );
  OAI211_X1 U9297 ( .C1(n10125), .C2(n10225), .A(n10130), .B(n10120), .ZN(
        n7487) );
  OAI22_X1 U9298 ( .A1(n10194), .A2(n10122), .B1(n10442), .B2(n6264), .ZN(
        n7484) );
  AOI21_X1 U9299 ( .B1(n7487), .B2(n10442), .A(n7484), .ZN(n7485) );
  INV_X1 U9300 ( .A(n7485), .ZN(P1_U3523) );
  INV_X1 U9301 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9126) );
  OAI22_X1 U9302 ( .A1(n10266), .A2(n10122), .B1(n10430), .B2(n9126), .ZN(
        n7486) );
  AOI21_X1 U9303 ( .B1(n7487), .B2(n10430), .A(n7486), .ZN(n7488) );
  INV_X1 U9304 ( .A(n7488), .ZN(P1_U3456) );
  INV_X1 U9305 ( .A(n7489), .ZN(n7500) );
  NAND2_X1 U9306 ( .A1(n7512), .A2(n10473), .ZN(n10494) );
  AOI21_X1 U9307 ( .B1(n7491), .B2(n7490), .A(n8281), .ZN(n7493) );
  NAND2_X1 U9308 ( .A1(n7493), .A2(n7492), .ZN(n7499) );
  OAI21_X1 U9309 ( .B1(n8274), .B2(n7495), .A(n7494), .ZN(n7497) );
  NOR2_X1 U9310 ( .A1(n8248), .A2(n7510), .ZN(n7496) );
  AOI211_X1 U9311 ( .C1(n8258), .C2(n8300), .A(n7497), .B(n7496), .ZN(n7498)
         );
  OAI211_X1 U9312 ( .C1(n7500), .C2(n10494), .A(n7499), .B(n7498), .ZN(
        P2_U3179) );
  INV_X1 U9313 ( .A(n7501), .ZN(n7504) );
  OAI222_X1 U9314 ( .A1(n8105), .A2(n7502), .B1(n8004), .B2(n7504), .C1(
        P1_U3086), .C2(n9551), .ZN(P1_U3336) );
  OAI222_X1 U9315 ( .A1(n8804), .A2(n9061), .B1(n7691), .B2(n7504), .C1(
        P2_U3151), .C2(n7503), .ZN(P2_U3276) );
  XNOR2_X1 U9316 ( .A(n7505), .B(n7506), .ZN(n10496) );
  XOR2_X1 U9317 ( .A(n7507), .B(n7506), .Z(n7508) );
  AOI222_X1 U9318 ( .A1(n8696), .A2(n7508), .B1(n8300), .B2(n8692), .C1(n8302), 
        .C2(n8609), .ZN(n10495) );
  MUX2_X1 U9319 ( .A(n7509), .B(n10495), .S(n10464), .Z(n7514) );
  INV_X1 U9320 ( .A(n7510), .ZN(n7511) );
  AOI22_X1 U9321 ( .A1(n8589), .A2(n7512), .B1(n8588), .B2(n7511), .ZN(n7513)
         );
  OAI211_X1 U9322 ( .C1(n8553), .C2(n10496), .A(n7514), .B(n7513), .ZN(
        P2_U3227) );
  INV_X1 U9323 ( .A(n7520), .ZN(n9432) );
  OAI211_X1 U9324 ( .C1(n4391), .C2(n9572), .A(n7515), .B(n9432), .ZN(n7516)
         );
  NAND2_X1 U9325 ( .A1(n7516), .A2(n7755), .ZN(n10111) );
  AOI211_X1 U9326 ( .C1(n7518), .C2(n7517), .A(n10214), .B(n10100), .ZN(n10116) );
  OAI21_X1 U9327 ( .B1(n10122), .B2(n9572), .A(n7519), .ZN(n7521) );
  XNOR2_X1 U9328 ( .A(n7521), .B(n7520), .ZN(n7522) );
  OAI222_X1 U9329 ( .A1(n6460), .A2(n9480), .B1(n6461), .B2(n9214), .C1(n6464), 
        .C2(n7522), .ZN(n10113) );
  AOI211_X1 U9330 ( .C1(n10424), .C2(n10111), .A(n10116), .B(n10113), .ZN(
        n7528) );
  INV_X1 U9331 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7523) );
  INV_X1 U9332 ( .A(n7524), .ZN(n7525) );
  OAI21_X1 U9333 ( .B1(n7528), .B2(n7114), .A(n7525), .ZN(P1_U3459) );
  INV_X1 U9334 ( .A(n7526), .ZN(n7527) );
  OAI21_X1 U9335 ( .B1(n7528), .B2(n10440), .A(n7527), .ZN(P1_U3524) );
  AOI21_X1 U9336 ( .B1(n7530), .B2(n7529), .A(n9211), .ZN(n7536) );
  NAND2_X1 U9337 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9586) );
  INV_X1 U9338 ( .A(n9586), .ZN(n7532) );
  OAI22_X1 U9339 ( .A1(n10108), .A2(n9277), .B1(n9301), .B2(n10361), .ZN(n7531) );
  AOI211_X1 U9340 ( .C1(n10104), .C2(n9256), .A(n7532), .B(n7531), .ZN(n7535)
         );
  NAND2_X1 U9341 ( .A1(n9305), .A2(n7533), .ZN(n7534) );
  OAI211_X1 U9342 ( .C1(n7536), .C2(n9307), .A(n7535), .B(n7534), .ZN(P1_U3218) );
  INV_X1 U9343 ( .A(n7537), .ZN(n7540) );
  INV_X1 U9344 ( .A(n7538), .ZN(n7539) );
  AOI21_X1 U9345 ( .B1(n7540), .B2(n7542), .A(n7539), .ZN(n10482) );
  XNOR2_X1 U9346 ( .A(n7542), .B(n7541), .ZN(n7543) );
  AOI222_X1 U9347 ( .A1(n8696), .A2(n7543), .B1(n6771), .B2(n8609), .C1(n8302), 
        .C2(n8692), .ZN(n10483) );
  MUX2_X1 U9348 ( .A(n9140), .B(n10483), .S(n10464), .Z(n7547) );
  AOI22_X1 U9349 ( .A1(n8589), .A2(n7545), .B1(n8588), .B2(n7544), .ZN(n7546)
         );
  OAI211_X1 U9350 ( .C1(n10482), .C2(n8553), .A(n7547), .B(n7546), .ZN(
        P2_U3229) );
  INV_X1 U9351 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n8962) );
  INV_X1 U9352 ( .A(n7619), .ZN(n7548) );
  AOI21_X1 U9353 ( .B1(n7550), .B2(n7549), .A(n7548), .ZN(n7553) );
  XOR2_X1 U9354 ( .A(n7551), .B(P2_REG1_REG_3__SCAN_IN), .Z(n7552) );
  OAI22_X1 U9355 ( .A1(n8389), .A2(n7553), .B1(n7552), .B2(n8411), .ZN(n7554)
         );
  AOI211_X1 U9356 ( .C1(n4642), .C2(n10444), .A(n7555), .B(n7554), .ZN(n7560)
         );
  OAI21_X1 U9357 ( .B1(n7557), .B2(n7556), .A(n7625), .ZN(n7558) );
  INV_X1 U9358 ( .A(n8404), .ZN(n10452) );
  NAND2_X1 U9359 ( .A1(n7558), .A2(n10452), .ZN(n7559) );
  OAI211_X1 U9360 ( .C1(n8962), .C2(n7916), .A(n7560), .B(n7559), .ZN(P2_U3185) );
  INV_X1 U9361 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7575) );
  OAI21_X1 U9362 ( .B1(n7563), .B2(n7562), .A(n7561), .ZN(n7569) );
  XOR2_X1 U9363 ( .A(n7565), .B(n7564), .Z(n7566) );
  NOR2_X1 U9364 ( .A1(n8411), .A2(n7566), .ZN(n7568) );
  OAI22_X1 U9365 ( .A1(n8401), .A2(n6567), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5299), .ZN(n7567) );
  AOI211_X1 U9366 ( .C1(n8396), .C2(n7569), .A(n7568), .B(n7567), .ZN(n7574)
         );
  XOR2_X1 U9367 ( .A(n7571), .B(n7570), .Z(n7572) );
  NAND2_X1 U9368 ( .A1(n7572), .A2(n10452), .ZN(n7573) );
  OAI211_X1 U9369 ( .C1(n7575), .C2(n7916), .A(n7574), .B(n7573), .ZN(P2_U3184) );
  XOR2_X1 U9370 ( .A(n7577), .B(n7576), .Z(n7590) );
  NAND3_X1 U9371 ( .A1(n7635), .A2(n7578), .A3(n4393), .ZN(n7579) );
  AOI21_X1 U9372 ( .B1(n4495), .B2(n7579), .A(n8389), .ZN(n7588) );
  NAND3_X1 U9373 ( .A1(n7644), .A2(n7581), .A3(n7580), .ZN(n7582) );
  AOI21_X1 U9374 ( .B1(n7654), .B2(n7582), .A(n8404), .ZN(n7587) );
  INV_X1 U9375 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U9376 ( .A1(n10444), .A2(n7583), .ZN(n7584) );
  NAND2_X1 U9377 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7774) );
  OAI211_X1 U9378 ( .C1(n7916), .C2(n7585), .A(n7584), .B(n7774), .ZN(n7586)
         );
  NOR3_X1 U9379 ( .A1(n7588), .A2(n7587), .A3(n7586), .ZN(n7589) );
  OAI21_X1 U9380 ( .B1(n7590), .B2(n8411), .A(n7589), .ZN(P2_U3190) );
  XNOR2_X1 U9381 ( .A(n8057), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U9382 ( .A1(n7597), .A2(n8002), .ZN(n7591) );
  NAND2_X1 U9383 ( .A1(n7592), .A2(n7591), .ZN(n7594) );
  INV_X1 U9384 ( .A(n8059), .ZN(n7593) );
  AOI211_X1 U9385 ( .C1(n7595), .C2(n7594), .A(n10302), .B(n7593), .ZN(n7609)
         );
  XNOR2_X1 U9386 ( .A(n8057), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9387 ( .A1(n7597), .A2(n7596), .ZN(n7598) );
  NAND2_X1 U9388 ( .A1(n7599), .A2(n7598), .ZN(n7601) );
  INV_X1 U9389 ( .A(n8047), .ZN(n7600) );
  AOI211_X1 U9390 ( .C1(n7602), .C2(n7601), .A(n10316), .B(n7600), .ZN(n7608)
         );
  INV_X1 U9391 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7606) );
  NAND2_X1 U9392 ( .A1(n10312), .A2(n8057), .ZN(n7605) );
  NOR2_X1 U9393 ( .A1(n7603), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9245) );
  INV_X1 U9394 ( .A(n9245), .ZN(n7604) );
  OAI211_X1 U9395 ( .C1(n7606), .C2(n10332), .A(n7605), .B(n7604), .ZN(n7607)
         );
  OR3_X1 U9396 ( .A1(n7609), .A2(n7608), .A3(n7607), .ZN(P1_U3256) );
  INV_X1 U9397 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7633) );
  OAI21_X1 U9398 ( .B1(n7612), .B2(n7611), .A(n7610), .ZN(n7624) );
  INV_X1 U9399 ( .A(n7613), .ZN(n7614) );
  OAI21_X1 U9400 ( .B1(n8401), .B2(n7615), .A(n7614), .ZN(n7623) );
  INV_X1 U9401 ( .A(n7616), .ZN(n7618) );
  NAND3_X1 U9402 ( .A1(n7619), .A2(n7618), .A3(n7617), .ZN(n7620) );
  AOI21_X1 U9403 ( .B1(n7621), .B2(n7620), .A(n8389), .ZN(n7622) );
  AOI211_X1 U9404 ( .C1(n8385), .C2(n7624), .A(n7623), .B(n7622), .ZN(n7632)
         );
  INV_X1 U9405 ( .A(n7625), .ZN(n7628) );
  OAI21_X1 U9406 ( .B1(n7628), .B2(n7627), .A(n7626), .ZN(n7630) );
  NAND3_X1 U9407 ( .A1(n7630), .A2(n10452), .A3(n7629), .ZN(n7631) );
  OAI211_X1 U9408 ( .C1(n7916), .C2(n7633), .A(n7632), .B(n7631), .ZN(P2_U3186) );
  XNOR2_X1 U9409 ( .A(n7634), .B(n7768), .ZN(n7649) );
  OAI21_X1 U9410 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7636), .A(n7635), .ZN(
        n7647) );
  INV_X1 U9411 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7639) );
  AND2_X1 U9412 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7715) );
  AOI21_X1 U9413 ( .B1(n10444), .B2(n7637), .A(n7715), .ZN(n7638) );
  OAI21_X1 U9414 ( .B1(n7916), .B2(n7639), .A(n7638), .ZN(n7646) );
  NAND3_X1 U9415 ( .A1(n7642), .A2(n7641), .A3(n7640), .ZN(n7643) );
  AOI21_X1 U9416 ( .B1(n7644), .B2(n7643), .A(n8404), .ZN(n7645) );
  AOI211_X1 U9417 ( .C1(n7647), .C2(n8396), .A(n7646), .B(n7645), .ZN(n7648)
         );
  OAI21_X1 U9418 ( .B1(n7649), .B2(n8411), .A(n7648), .ZN(P2_U3189) );
  XNOR2_X1 U9419 ( .A(n7650), .B(n7883), .ZN(n7663) );
  OAI21_X1 U9420 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7651), .A(n7741), .ZN(
        n7661) );
  NAND3_X1 U9421 ( .A1(n7654), .A2(n7653), .A3(n7652), .ZN(n7655) );
  AOI21_X1 U9422 ( .B1(n7748), .B2(n7655), .A(n8404), .ZN(n7660) );
  INV_X1 U9423 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7658) );
  AND2_X1 U9424 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7807) );
  AOI21_X1 U9425 ( .B1(n10444), .B2(n7656), .A(n7807), .ZN(n7657) );
  OAI21_X1 U9426 ( .B1(n7916), .B2(n7658), .A(n7657), .ZN(n7659) );
  AOI211_X1 U9427 ( .C1(n7661), .C2(n8396), .A(n7660), .B(n7659), .ZN(n7662)
         );
  OAI21_X1 U9428 ( .B1(n7663), .B2(n8411), .A(n7662), .ZN(P2_U3191) );
  NAND2_X1 U9429 ( .A1(n7664), .A2(n7665), .ZN(n7666) );
  XNOR2_X1 U9430 ( .A(n7666), .B(n7669), .ZN(n7667) );
  AOI222_X1 U9431 ( .A1(n8696), .A2(n7667), .B1(n8300), .B2(n8609), .C1(n8608), 
        .C2(n8692), .ZN(n7723) );
  AOI22_X1 U9432 ( .A1(n6752), .A2(n7780), .B1(P2_REG0_REG_8__SCAN_IN), .B2(
        n10499), .ZN(n7672) );
  NAND2_X1 U9433 ( .A1(n7695), .A2(n7668), .ZN(n7670) );
  XNOR2_X1 U9434 ( .A(n7670), .B(n7669), .ZN(n7722) );
  NAND2_X1 U9435 ( .A1(n7878), .A2(n6736), .ZN(n10487) );
  INV_X1 U9436 ( .A(n10487), .ZN(n10497) );
  INV_X1 U9437 ( .A(n8775), .ZN(n8786) );
  NAND2_X1 U9438 ( .A1(n7722), .A2(n8786), .ZN(n7671) );
  OAI211_X1 U9439 ( .C1(n7723), .C2(n10499), .A(n7672), .B(n7671), .ZN(
        P2_U3414) );
  INV_X1 U9440 ( .A(n7673), .ZN(n8622) );
  NAND3_X1 U9441 ( .A1(n7538), .A2(n7676), .A3(n7675), .ZN(n7677) );
  NAND2_X1 U9442 ( .A1(n7674), .A2(n7677), .ZN(n10492) );
  OAI22_X1 U9443 ( .A1(n8618), .A2(n10489), .B1(n7678), .B2(n10458), .ZN(n7687) );
  NAND2_X1 U9444 ( .A1(n7680), .A2(n7679), .ZN(n7682) );
  XNOR2_X1 U9445 ( .A(n7682), .B(n7681), .ZN(n7685) );
  NAND2_X1 U9446 ( .A1(n10492), .A2(n8689), .ZN(n7684) );
  AOI22_X1 U9447 ( .A1(n8609), .A2(n8303), .B1(n8301), .B2(n8692), .ZN(n7683)
         );
  OAI211_X1 U9448 ( .C1(n7685), .C2(n10469), .A(n7684), .B(n7683), .ZN(n10490)
         );
  MUX2_X1 U9449 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10490), .S(n10464), .Z(n7686) );
  AOI211_X1 U9450 ( .C1(n8622), .C2(n10492), .A(n7687), .B(n7686), .ZN(n7688)
         );
  INV_X1 U9451 ( .A(n7688), .ZN(P2_U3228) );
  INV_X1 U9452 ( .A(n7689), .ZN(n7706) );
  OAI222_X1 U9453 ( .A1(n8804), .A2(n7692), .B1(n7691), .B2(n7706), .C1(n7690), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  OR2_X1 U9454 ( .A1(n7693), .A2(n7696), .ZN(n7694) );
  NAND2_X1 U9455 ( .A1(n7695), .A2(n7694), .ZN(n7704) );
  INV_X1 U9456 ( .A(n7704), .ZN(n7818) );
  NAND2_X1 U9457 ( .A1(n7697), .A2(n7696), .ZN(n7698) );
  NAND2_X1 U9458 ( .A1(n7664), .A2(n7698), .ZN(n7702) );
  NAND2_X1 U9459 ( .A1(n8692), .A2(n8299), .ZN(n7699) );
  OAI21_X1 U9460 ( .B1(n7700), .B2(n8694), .A(n7699), .ZN(n7701) );
  AOI21_X1 U9461 ( .B1(n7702), .B2(n8696), .A(n7701), .ZN(n7703) );
  OAI21_X1 U9462 ( .B1(n7704), .B2(n7878), .A(n7703), .ZN(n7815) );
  AOI21_X1 U9463 ( .B1(n10493), .B2(n7818), .A(n7815), .ZN(n7767) );
  AOI22_X1 U9464 ( .A1(n6752), .A2(n7719), .B1(P2_REG0_REG_7__SCAN_IN), .B2(
        n10499), .ZN(n7705) );
  OAI21_X1 U9465 ( .B1(n7767), .B2(n10499), .A(n7705), .ZN(P2_U3411) );
  OAI222_X1 U9466 ( .A1(n8105), .A2(n7707), .B1(P1_U3086), .B2(n9539), .C1(
        n10283), .C2(n7706), .ZN(P1_U3335) );
  MUX2_X1 U9467 ( .A(n7708), .B(n7723), .S(n10508), .Z(n7710) );
  INV_X1 U9468 ( .A(n8667), .ZN(n8674) );
  AOI22_X1 U9469 ( .A1(n7722), .A2(n8674), .B1(n8673), .B2(n7780), .ZN(n7709)
         );
  NAND2_X1 U9470 ( .A1(n7710), .A2(n7709), .ZN(P2_U3467) );
  INV_X1 U9471 ( .A(n7711), .ZN(n7712) );
  AOI21_X1 U9472 ( .B1(n7714), .B2(n7713), .A(n7712), .ZN(n7721) );
  AOI21_X1 U9473 ( .B1(n8286), .B2(n8301), .A(n7715), .ZN(n7716) );
  OAI21_X1 U9474 ( .B1(n7770), .B2(n8288), .A(n7716), .ZN(n7718) );
  NOR2_X1 U9475 ( .A1(n8248), .A2(n7813), .ZN(n7717) );
  AOI211_X1 U9476 ( .C1(n8263), .C2(n7719), .A(n7718), .B(n7717), .ZN(n7720)
         );
  OAI21_X1 U9477 ( .B1(n7721), .B2(n8281), .A(n7720), .ZN(P2_U3153) );
  INV_X1 U9478 ( .A(n7722), .ZN(n7728) );
  MUX2_X1 U9479 ( .A(n7724), .B(n7723), .S(n10464), .Z(n7727) );
  INV_X1 U9480 ( .A(n7777), .ZN(n7725) );
  AOI22_X1 U9481 ( .A1(n8589), .A2(n7780), .B1(n8588), .B2(n7725), .ZN(n7726)
         );
  OAI211_X1 U9482 ( .C1(n7728), .C2(n8553), .A(n7727), .B(n7726), .ZN(P2_U3225) );
  INV_X1 U9483 ( .A(n7729), .ZN(n7733) );
  OAI222_X1 U9484 ( .A1(n8804), .A2(n7731), .B1(n8811), .B2(n7733), .C1(
        P2_U3151), .C2(n7730), .ZN(P2_U3273) );
  OAI222_X1 U9485 ( .A1(n8105), .A2(n7734), .B1(n8004), .B2(n7733), .C1(n7732), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  XOR2_X1 U9486 ( .A(n7736), .B(n7735), .Z(n7753) );
  NAND2_X1 U9487 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8128) );
  OAI21_X1 U9488 ( .B1(n8401), .B2(n7737), .A(n8128), .ZN(n7745) );
  INV_X1 U9489 ( .A(n7738), .ZN(n7743) );
  NAND3_X1 U9490 ( .A1(n7741), .A2(n7740), .A3(n7739), .ZN(n7742) );
  AOI21_X1 U9491 ( .B1(n7743), .B2(n7742), .A(n8389), .ZN(n7744) );
  AOI211_X1 U9492 ( .C1(n10443), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7745), .B(
        n7744), .ZN(n7752) );
  INV_X1 U9493 ( .A(n7912), .ZN(n7750) );
  AND3_X1 U9494 ( .A1(n7748), .A2(n7747), .A3(n7746), .ZN(n7749) );
  OAI21_X1 U9495 ( .B1(n7750), .B2(n7749), .A(n10452), .ZN(n7751) );
  OAI211_X1 U9496 ( .C1(n7753), .C2(n8411), .A(n7752), .B(n7751), .ZN(P2_U3192) );
  AND2_X1 U9497 ( .A1(n7755), .A2(n7754), .ZN(n10096) );
  INV_X1 U9498 ( .A(n10105), .ZN(n10095) );
  NOR2_X1 U9499 ( .A1(n10096), .A2(n10095), .ZN(n10094) );
  NOR2_X1 U9500 ( .A1(n10094), .A2(n7756), .ZN(n10365) );
  XNOR2_X1 U9501 ( .A(n10364), .B(n5957), .ZN(n9435) );
  XNOR2_X1 U9502 ( .A(n10365), .B(n9435), .ZN(n10093) );
  XNOR2_X1 U9503 ( .A(n7757), .B(n9435), .ZN(n7758) );
  AOI222_X1 U9504 ( .A1(n9569), .A2(n10017), .B1(n9570), .B2(n10356), .C1(
        n10014), .C2(n7758), .ZN(n10085) );
  AOI21_X1 U9505 ( .B1(n10099), .B2(n9216), .A(n10214), .ZN(n7760) );
  NAND2_X1 U9506 ( .A1(n7760), .A2(n7759), .ZN(n10086) );
  OAI211_X1 U9507 ( .C1(n10225), .C2(n10093), .A(n10085), .B(n10086), .ZN(
        n7765) );
  INV_X1 U9508 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7761) );
  OAI22_X1 U9509 ( .A1(n10266), .A2(n5957), .B1(n10430), .B2(n7761), .ZN(n7762) );
  AOI21_X1 U9510 ( .B1(n7765), .B2(n10430), .A(n7762), .ZN(n7763) );
  INV_X1 U9511 ( .A(n7763), .ZN(P1_U3465) );
  OAI22_X1 U9512 ( .A1(n10194), .A2(n5957), .B1(n10442), .B2(n9168), .ZN(n7764) );
  AOI21_X1 U9513 ( .B1(n7765), .B2(n10442), .A(n7764), .ZN(n7766) );
  INV_X1 U9514 ( .A(n7766), .ZN(P1_U3526) );
  MUX2_X1 U9515 ( .A(n7768), .B(n7767), .S(n10508), .Z(n7769) );
  OAI21_X1 U9516 ( .B1(n7814), .B2(n8686), .A(n7769), .ZN(P2_U3466) );
  XNOR2_X1 U9517 ( .A(n7771), .B(n7770), .ZN(n7772) );
  XNOR2_X1 U9518 ( .A(n7773), .B(n7772), .ZN(n7782) );
  NAND2_X1 U9519 ( .A1(n8286), .A2(n8300), .ZN(n7775) );
  OAI211_X1 U9520 ( .C1(n7776), .C2(n8288), .A(n7775), .B(n7774), .ZN(n7779)
         );
  NOR2_X1 U9521 ( .A1(n8248), .A2(n7777), .ZN(n7778) );
  AOI211_X1 U9522 ( .C1(n8263), .C2(n7780), .A(n7779), .B(n7778), .ZN(n7781)
         );
  OAI21_X1 U9523 ( .B1(n7782), .B2(n8281), .A(n7781), .ZN(P2_U3161) );
  INV_X1 U9524 ( .A(n7790), .ZN(n7785) );
  AOI21_X1 U9525 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8809), .A(n7783), .ZN(
        n7784) );
  OAI21_X1 U9526 ( .B1(n7785), .B2(n8811), .A(n7784), .ZN(P2_U3272) );
  INV_X1 U9527 ( .A(n7786), .ZN(n7792) );
  OAI222_X1 U9528 ( .A1(n8804), .A2(n7788), .B1(n8811), .B2(n7792), .C1(n7787), 
        .C2(P2_U3151), .ZN(P2_U3274) );
  NAND2_X1 U9529 ( .A1(n7790), .A2(n7789), .ZN(n7791) );
  OR2_X1 U9530 ( .A1(n9548), .A2(P1_U3086), .ZN(n9556) );
  OAI211_X1 U9531 ( .C1(n9062), .C2(n8105), .A(n7791), .B(n9556), .ZN(P1_U3332) );
  XNOR2_X1 U9532 ( .A(n7795), .B(n7794), .ZN(n7802) );
  NAND2_X1 U9533 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9643) );
  INV_X1 U9534 ( .A(n9643), .ZN(n7796) );
  AOI21_X1 U9535 ( .B1(n9299), .B2(n9568), .A(n7796), .ZN(n7800) );
  NAND2_X1 U9536 ( .A1(n9256), .A2(n10343), .ZN(n7799) );
  NAND2_X1 U9537 ( .A1(n9305), .A2(n10342), .ZN(n7798) );
  NAND2_X1 U9538 ( .A1(n9289), .A2(n9566), .ZN(n7797) );
  NAND4_X1 U9539 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n7801)
         );
  AOI21_X1 U9540 ( .B1(n7802), .B2(n9287), .A(n7801), .ZN(n7803) );
  INV_X1 U9541 ( .A(n7803), .ZN(P1_U3213) );
  XNOR2_X1 U9542 ( .A(n7805), .B(n7804), .ZN(n7812) );
  INV_X1 U9543 ( .A(n8616), .ZN(n7806) );
  NAND2_X1 U9544 ( .A1(n8290), .A2(n7806), .ZN(n7809) );
  AOI21_X1 U9545 ( .B1(n8286), .B2(n8299), .A(n7807), .ZN(n7808) );
  OAI211_X1 U9546 ( .C1(n8156), .C2(n8288), .A(n7809), .B(n7808), .ZN(n7810)
         );
  AOI21_X1 U9547 ( .B1(n8263), .B2(n7868), .A(n7810), .ZN(n7811) );
  OAI21_X1 U9548 ( .B1(n7812), .B2(n8281), .A(n7811), .ZN(P2_U3171) );
  OAI22_X1 U9549 ( .A1(n8618), .A2(n7814), .B1(n7813), .B2(n10458), .ZN(n7817)
         );
  MUX2_X1 U9550 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7815), .S(n10464), .Z(n7816)
         );
  AOI211_X1 U9551 ( .C1(n7818), .C2(n8622), .A(n7817), .B(n7816), .ZN(n7819)
         );
  INV_X1 U9552 ( .A(n7819), .ZN(P2_U3226) );
  INV_X1 U9553 ( .A(n7824), .ZN(n9213) );
  NAND3_X1 U9554 ( .A1(n9213), .A2(n7820), .A3(n7821), .ZN(n7851) );
  INV_X1 U9555 ( .A(n7821), .ZN(n7823) );
  OAI21_X1 U9556 ( .B1(n7824), .B2(n7823), .A(n7822), .ZN(n7852) );
  NAND2_X1 U9557 ( .A1(n7851), .A2(n7852), .ZN(n7825) );
  XNOR2_X1 U9558 ( .A(n7825), .B(n7853), .ZN(n7830) );
  NAND2_X1 U9559 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9615) );
  INV_X1 U9560 ( .A(n9615), .ZN(n7827) );
  NOR2_X1 U9561 ( .A1(n9277), .A2(n10361), .ZN(n7826) );
  AOI211_X1 U9562 ( .C1(n9289), .C2(n9568), .A(n7827), .B(n7826), .ZN(n7829)
         );
  AOI22_X1 U9563 ( .A1(n9305), .A2(n10357), .B1(n10360), .B2(n9256), .ZN(n7828) );
  OAI211_X1 U9564 ( .C1(n7830), .C2(n9307), .A(n7829), .B(n7828), .ZN(P1_U3227) );
  INV_X1 U9565 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10518) );
  INV_X1 U9566 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10331) );
  NOR2_X1 U9567 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7831) );
  AOI21_X1 U9568 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7831), .ZN(n10521) );
  INV_X1 U9569 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9124) );
  INV_X1 U9570 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9122) );
  AOI22_X1 U9571 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n9124), .B2(n9122), .ZN(n10524) );
  INV_X1 U9572 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9072) );
  INV_X1 U9573 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U9574 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .B1(n9072), .B2(n10315), .ZN(n10527) );
  NOR2_X1 U9575 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n7832) );
  AOI21_X1 U9576 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n7832), .ZN(n10530) );
  NOR2_X1 U9577 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7833) );
  AOI21_X1 U9578 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7833), .ZN(n10533) );
  NOR2_X1 U9579 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7834) );
  AOI21_X1 U9580 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7834), .ZN(n10536) );
  NOR2_X1 U9581 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7835) );
  AOI21_X1 U9582 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7835), .ZN(n10539) );
  NOR2_X1 U9583 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7836) );
  AOI21_X1 U9584 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7836), .ZN(n10542) );
  NOR2_X1 U9585 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7837) );
  AOI21_X1 U9586 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7837), .ZN(n10551) );
  NOR2_X1 U9587 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7838) );
  AOI21_X1 U9588 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7838), .ZN(n10557) );
  NOR2_X1 U9589 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7839) );
  AOI21_X1 U9590 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7839), .ZN(n10554) );
  NOR2_X1 U9591 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7840) );
  AOI21_X1 U9592 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7840), .ZN(n10548) );
  NOR2_X1 U9593 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7841) );
  AOI21_X1 U9594 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7841), .ZN(n10545) );
  AND2_X1 U9595 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7842) );
  NOR2_X1 U9596 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7842), .ZN(n10510) );
  INV_X1 U9597 ( .A(n10510), .ZN(n10511) );
  INV_X1 U9598 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10513) );
  NAND3_X1 U9599 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10512) );
  NAND2_X1 U9600 ( .A1(n10513), .A2(n10512), .ZN(n10509) );
  NAND2_X1 U9601 ( .A1(n10511), .A2(n10509), .ZN(n10560) );
  NAND2_X1 U9602 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7843) );
  OAI21_X1 U9603 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7843), .ZN(n10559) );
  NOR2_X1 U9604 ( .A1(n10560), .A2(n10559), .ZN(n10558) );
  AOI21_X1 U9605 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10558), .ZN(n10563) );
  NAND2_X1 U9606 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7844) );
  OAI21_X1 U9607 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7844), .ZN(n10562) );
  NOR2_X1 U9608 ( .A1(n10563), .A2(n10562), .ZN(n10561) );
  AOI21_X1 U9609 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10561), .ZN(n10566) );
  NOR2_X1 U9610 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7845) );
  AOI21_X1 U9611 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7845), .ZN(n10565) );
  NAND2_X1 U9612 ( .A1(n10566), .A2(n10565), .ZN(n10564) );
  OAI21_X1 U9613 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10564), .ZN(n10544) );
  NAND2_X1 U9614 ( .A1(n10545), .A2(n10544), .ZN(n10543) );
  OAI21_X1 U9615 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10543), .ZN(n10547) );
  NAND2_X1 U9616 ( .A1(n10548), .A2(n10547), .ZN(n10546) );
  OAI21_X1 U9617 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10546), .ZN(n10553) );
  NAND2_X1 U9618 ( .A1(n10554), .A2(n10553), .ZN(n10552) );
  OAI21_X1 U9619 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10552), .ZN(n10556) );
  NAND2_X1 U9620 ( .A1(n10557), .A2(n10556), .ZN(n10555) );
  OAI21_X1 U9621 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10555), .ZN(n10550) );
  NAND2_X1 U9622 ( .A1(n10551), .A2(n10550), .ZN(n10549) );
  OAI21_X1 U9623 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10549), .ZN(n10541) );
  NAND2_X1 U9624 ( .A1(n10542), .A2(n10541), .ZN(n10540) );
  OAI21_X1 U9625 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10540), .ZN(n10538) );
  NAND2_X1 U9626 ( .A1(n10539), .A2(n10538), .ZN(n10537) );
  OAI21_X1 U9627 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10537), .ZN(n10535) );
  NAND2_X1 U9628 ( .A1(n10536), .A2(n10535), .ZN(n10534) );
  OAI21_X1 U9629 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10534), .ZN(n10532) );
  NAND2_X1 U9630 ( .A1(n10533), .A2(n10532), .ZN(n10531) );
  OAI21_X1 U9631 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10531), .ZN(n10529) );
  NAND2_X1 U9632 ( .A1(n10530), .A2(n10529), .ZN(n10528) );
  OAI21_X1 U9633 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10528), .ZN(n10526) );
  NAND2_X1 U9634 ( .A1(n10527), .A2(n10526), .ZN(n10525) );
  OAI21_X1 U9635 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10525), .ZN(n10523) );
  NAND2_X1 U9636 ( .A1(n10524), .A2(n10523), .ZN(n10522) );
  OAI21_X1 U9637 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10522), .ZN(n10520) );
  NAND2_X1 U9638 ( .A1(n10521), .A2(n10520), .ZN(n10519) );
  OAI21_X1 U9639 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10519), .ZN(n7846) );
  OR2_X1 U9640 ( .A1(n10331), .A2(n7846), .ZN(n10517) );
  NAND2_X1 U9641 ( .A1(n10518), .A2(n10517), .ZN(n10514) );
  NAND2_X1 U9642 ( .A1(n10331), .A2(n7846), .ZN(n10516) );
  NAND2_X1 U9643 ( .A1(n10514), .A2(n10516), .ZN(n7848) );
  XNOR2_X1 U9644 ( .A(n8078), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7847) );
  XNOR2_X1 U9645 ( .A(n7848), .B(n7847), .ZN(ADD_1068_U4) );
  NAND2_X1 U9646 ( .A1(n8402), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7849) );
  OAI21_X1 U9647 ( .B1(n7850), .B2(n8402), .A(n7849), .ZN(P2_U3521) );
  INV_X1 U9648 ( .A(n7851), .ZN(n7854) );
  OAI21_X1 U9649 ( .B1(n7854), .B2(n7853), .A(n7852), .ZN(n7859) );
  OAI21_X1 U9650 ( .B1(n7857), .B2(n7856), .A(n7855), .ZN(n7858) );
  XNOR2_X1 U9651 ( .A(n7859), .B(n7858), .ZN(n7866) );
  NAND2_X1 U9652 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9629) );
  INV_X1 U9653 ( .A(n9629), .ZN(n7860) );
  AOI21_X1 U9654 ( .B1(n9299), .B2(n9569), .A(n7860), .ZN(n7864) );
  NAND2_X1 U9655 ( .A1(n9256), .A2(n10079), .ZN(n7863) );
  NAND2_X1 U9656 ( .A1(n9305), .A2(n10078), .ZN(n7862) );
  NAND2_X1 U9657 ( .A1(n9289), .A2(n9567), .ZN(n7861) );
  NAND4_X1 U9658 ( .A1(n7864), .A2(n7863), .A3(n7862), .A4(n7861), .ZN(n7865)
         );
  AOI21_X1 U9659 ( .B1(n7866), .B2(n9287), .A(n7865), .ZN(n7867) );
  INV_X1 U9660 ( .A(n7867), .ZN(P1_U3239) );
  INV_X1 U9661 ( .A(n7868), .ZN(n8617) );
  INV_X1 U9662 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7880) );
  NAND2_X1 U9663 ( .A1(n7869), .A2(n7873), .ZN(n7870) );
  NAND2_X1 U9664 ( .A1(n8598), .A2(n7870), .ZN(n7879) );
  INV_X1 U9665 ( .A(n7879), .ZN(n8623) );
  AOI22_X1 U9666 ( .A1(n8609), .A2(n8299), .B1(n8692), .B2(n8298), .ZN(n7877)
         );
  AND2_X1 U9667 ( .A1(n7872), .A2(n7871), .ZN(n7874) );
  XNOR2_X1 U9668 ( .A(n7874), .B(n7873), .ZN(n7875) );
  NAND2_X1 U9669 ( .A1(n7875), .A2(n8696), .ZN(n7876) );
  OAI211_X1 U9670 ( .C1(n7879), .C2(n7878), .A(n7877), .B(n7876), .ZN(n8619)
         );
  AOI21_X1 U9671 ( .B1(n10493), .B2(n8623), .A(n8619), .ZN(n7882) );
  MUX2_X1 U9672 ( .A(n7880), .B(n7882), .S(n10501), .Z(n7881) );
  OAI21_X1 U9673 ( .B1(n8617), .B2(n8793), .A(n7881), .ZN(P2_U3417) );
  MUX2_X1 U9674 ( .A(n7883), .B(n7882), .S(n10508), .Z(n7884) );
  OAI21_X1 U9675 ( .B1(n8617), .B2(n8686), .A(n7884), .ZN(P2_U3468) );
  NAND2_X1 U9676 ( .A1(n8402), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7885) );
  OAI21_X1 U9677 ( .B1(n8422), .B2(n8402), .A(n7885), .ZN(P2_U3520) );
  NAND2_X1 U9678 ( .A1(n7886), .A2(n7887), .ZN(n8581) );
  XNOR2_X1 U9679 ( .A(n8581), .B(n7893), .ZN(n7888) );
  AOI222_X1 U9680 ( .A1(n8696), .A2(n7888), .B1(n8298), .B2(n8609), .C1(n8297), 
        .C2(n8692), .ZN(n7902) );
  MUX2_X1 U9681 ( .A(n7889), .B(n7902), .S(n10508), .Z(n7896) );
  INV_X1 U9682 ( .A(n8597), .ZN(n7890) );
  NOR2_X1 U9683 ( .A1(n8604), .A2(n7890), .ZN(n7891) );
  NAND2_X1 U9684 ( .A1(n8598), .A2(n7891), .ZN(n8600) );
  NAND2_X1 U9685 ( .A1(n8600), .A2(n7892), .ZN(n7894) );
  XNOR2_X1 U9686 ( .A(n7894), .B(n7893), .ZN(n7901) );
  AOI22_X1 U9687 ( .A1(n7901), .A2(n8674), .B1(n8673), .B2(n8579), .ZN(n7895)
         );
  NAND2_X1 U9688 ( .A1(n7896), .A2(n7895), .ZN(P2_U3470) );
  MUX2_X1 U9689 ( .A(n7897), .B(n7902), .S(n10501), .Z(n7899) );
  AOI22_X1 U9690 ( .A1(n7901), .A2(n8786), .B1(n6752), .B2(n8579), .ZN(n7898)
         );
  NAND2_X1 U9691 ( .A1(n7899), .A2(n7898), .ZN(P2_U3423) );
  INV_X1 U9692 ( .A(n7900), .ZN(n8079) );
  OAI222_X1 U9693 ( .A1(P1_U3086), .A2(n6122), .B1(n8004), .B2(n8079), .C1(
        n9037), .C2(n8105), .ZN(P1_U3331) );
  INV_X1 U9694 ( .A(n7901), .ZN(n7907) );
  MUX2_X1 U9695 ( .A(n7903), .B(n7902), .S(n10464), .Z(n7906) );
  INV_X1 U9696 ( .A(n8247), .ZN(n7904) );
  AOI22_X1 U9697 ( .A1(n8589), .A2(n8579), .B1(n8588), .B2(n7904), .ZN(n7905)
         );
  OAI211_X1 U9698 ( .C1(n7907), .C2(n8553), .A(n7906), .B(n7905), .ZN(P2_U3222) );
  XNOR2_X1 U9699 ( .A(n7908), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n7921) );
  OAI21_X1 U9700 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n7909), .A(n7925), .ZN(
        n7919) );
  NAND3_X1 U9701 ( .A1(n7912), .A2(n7911), .A3(n7910), .ZN(n7913) );
  AOI21_X1 U9702 ( .B1(n7931), .B2(n7913), .A(n8404), .ZN(n7918) );
  INV_X1 U9703 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8960) );
  NAND2_X1 U9704 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U9705 ( .A1(n10444), .A2(n7914), .ZN(n7915) );
  OAI211_X1 U9706 ( .C1(n7916), .C2(n8960), .A(n8245), .B(n7915), .ZN(n7917)
         );
  AOI211_X1 U9707 ( .C1(n7919), .C2(n8396), .A(n7918), .B(n7917), .ZN(n7920)
         );
  OAI21_X1 U9708 ( .B1(n7921), .B2(n8411), .A(n7920), .ZN(P2_U3193) );
  XOR2_X1 U9709 ( .A(n7923), .B(n7922), .Z(n7937) );
  AND3_X1 U9710 ( .A1(n7925), .A2(n7924), .A3(n4411), .ZN(n7926) );
  OAI21_X1 U9711 ( .B1(n7927), .B2(n7926), .A(n8396), .ZN(n7936) );
  NAND2_X1 U9712 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8162) );
  OAI21_X1 U9713 ( .B1(n8401), .B2(n7928), .A(n8162), .ZN(n7934) );
  NAND3_X1 U9714 ( .A1(n7931), .A2(n7930), .A3(n7929), .ZN(n7932) );
  AOI21_X1 U9715 ( .B1(n8313), .B2(n7932), .A(n8404), .ZN(n7933) );
  AOI211_X1 U9716 ( .C1(n10443), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7934), .B(
        n7933), .ZN(n7935) );
  OAI211_X1 U9717 ( .C1(n7937), .C2(n8411), .A(n7936), .B(n7935), .ZN(P2_U3194) );
  INV_X1 U9718 ( .A(n7938), .ZN(n7939) );
  NOR2_X1 U9719 ( .A1(n7886), .A2(n7939), .ZN(n7942) );
  OAI21_X1 U9720 ( .B1(n7942), .B2(n7941), .A(n7940), .ZN(n7943) );
  XNOR2_X1 U9721 ( .A(n7943), .B(n7946), .ZN(n7944) );
  AOI222_X1 U9722 ( .A1(n8696), .A2(n7944), .B1(n8296), .B2(n8692), .C1(n8297), 
        .C2(n8609), .ZN(n7952) );
  MUX2_X1 U9723 ( .A(n7945), .B(n7952), .S(n10508), .Z(n7949) );
  XNOR2_X1 U9724 ( .A(n7947), .B(n7946), .ZN(n7956) );
  AOI22_X1 U9725 ( .A1(n7956), .A2(n8674), .B1(n8673), .B2(n8227), .ZN(n7948)
         );
  NAND2_X1 U9726 ( .A1(n7949), .A2(n7948), .ZN(P2_U3472) );
  MUX2_X1 U9727 ( .A(n8946), .B(n7952), .S(n10501), .Z(n7951) );
  AOI22_X1 U9728 ( .A1(n7956), .A2(n8786), .B1(n6752), .B2(n8227), .ZN(n7950)
         );
  NAND2_X1 U9729 ( .A1(n7951), .A2(n7950), .ZN(P2_U3429) );
  INV_X1 U9730 ( .A(n7952), .ZN(n7955) );
  OAI22_X1 U9731 ( .A1(n7953), .A2(n8567), .B1(n8225), .B2(n10458), .ZN(n7954)
         );
  OAI21_X1 U9732 ( .B1(n7955), .B2(n7954), .A(n10464), .ZN(n7958) );
  INV_X1 U9733 ( .A(n8553), .ZN(n8593) );
  AOI22_X1 U9734 ( .A1(n7956), .A2(n8593), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10466), .ZN(n7957) );
  NAND2_X1 U9735 ( .A1(n7958), .A2(n7957), .ZN(P2_U3220) );
  INV_X1 U9736 ( .A(n7959), .ZN(n8010) );
  NAND2_X1 U9737 ( .A1(n7960), .A2(n8305), .ZN(n7961) );
  OAI21_X1 U9738 ( .B1(n8305), .B2(n6073), .A(n7961), .ZN(P2_U3522) );
  XNOR2_X1 U9739 ( .A(n7962), .B(n9221), .ZN(n7964) );
  NOR2_X1 U9740 ( .A1(n7964), .A2(n7963), .ZN(n9220) );
  AOI21_X1 U9741 ( .B1(n7964), .B2(n7963), .A(n9220), .ZN(n7969) );
  NOR2_X1 U9742 ( .A1(n9302), .A2(n5986), .ZN(n7967) );
  NAND2_X1 U9743 ( .A1(n9299), .A2(n9567), .ZN(n7965) );
  NAND2_X1 U9744 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9656) );
  OAI211_X1 U9745 ( .C1(n10058), .C2(n9301), .A(n7965), .B(n9656), .ZN(n7966)
         );
  AOI211_X1 U9746 ( .C1(n10063), .C2(n9305), .A(n7967), .B(n7966), .ZN(n7968)
         );
  OAI21_X1 U9747 ( .B1(n7969), .B2(n9307), .A(n7968), .ZN(P1_U3221) );
  INV_X1 U9748 ( .A(n7970), .ZN(n7974) );
  OAI222_X1 U9749 ( .A1(n8804), .A2(n7972), .B1(n8811), .B2(n7974), .C1(n7971), 
        .C2(P2_U3151), .ZN(P2_U3269) );
  OAI222_X1 U9750 ( .A1(P1_U3086), .A2(n7975), .B1(n8004), .B2(n7974), .C1(
        n7973), .C2(n8105), .ZN(P1_U3329) );
  INV_X1 U9751 ( .A(n7976), .ZN(n7988) );
  AOI21_X1 U9752 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n8809), .A(n7977), .ZN(
        n7978) );
  OAI21_X1 U9753 ( .B1(n7988), .B2(n8811), .A(n7978), .ZN(P2_U3268) );
  OAI21_X1 U9754 ( .B1(n7981), .B2(n7980), .A(n7979), .ZN(n7982) );
  NAND2_X1 U9755 ( .A1(n7982), .A2(n9287), .ZN(n7987) );
  AOI21_X1 U9756 ( .B1(n9289), .B2(n9565), .A(n7983), .ZN(n7984) );
  OAI21_X1 U9757 ( .B1(n8853), .B2(n9277), .A(n7984), .ZN(n7985) );
  AOI21_X1 U9758 ( .B1(n9978), .B2(n9305), .A(n7985), .ZN(n7986) );
  OAI211_X1 U9759 ( .C1(n9981), .C2(n9302), .A(n7987), .B(n7986), .ZN(P1_U3224) );
  OAI222_X1 U9760 ( .A1(n8105), .A2(n7990), .B1(P1_U3086), .B2(n7989), .C1(
        n10283), .C2(n7988), .ZN(P1_U3328) );
  INV_X1 U9761 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U9762 ( .A1(n7992), .A2(n7991), .ZN(n7993) );
  XNOR2_X1 U9763 ( .A(n7993), .B(n9439), .ZN(n9976) );
  INV_X1 U9764 ( .A(n10227), .ZN(n10006) );
  NAND2_X1 U9765 ( .A1(n10021), .A2(n10006), .ZN(n9999) );
  AOI21_X1 U9766 ( .B1(n9999), .B2(n7994), .A(n10214), .ZN(n7995) );
  AND2_X1 U9767 ( .A1(n4491), .A2(n7995), .ZN(n9977) );
  XNOR2_X1 U9768 ( .A(n7997), .B(n9439), .ZN(n7998) );
  OAI222_X1 U9769 ( .A1(n6460), .A2(n8853), .B1(n6461), .B2(n9941), .C1(n6464), 
        .C2(n7998), .ZN(n9983) );
  AOI211_X1 U9770 ( .C1(n9976), .C2(n10424), .A(n9977), .B(n9983), .ZN(n8001)
         );
  MUX2_X1 U9771 ( .A(n7999), .B(n8001), .S(n10430), .Z(n8000) );
  OAI21_X1 U9772 ( .B1(n9981), .B2(n10266), .A(n8000), .ZN(P1_U3489) );
  MUX2_X1 U9773 ( .A(n8002), .B(n8001), .S(n10442), .Z(n8003) );
  OAI21_X1 U9774 ( .B1(n9981), .B2(n10194), .A(n8003), .ZN(P1_U3534) );
  INV_X1 U9775 ( .A(n8006), .ZN(n8803) );
  OAI222_X1 U9776 ( .A1(n8105), .A2(n8008), .B1(n10283), .B2(n8803), .C1(n8007), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U9777 ( .A1(P2_U3151), .A2(n6216), .B1(n8811), .B2(n8010), .C1(
        n8009), .C2(n8804), .ZN(P2_U3270) );
  NAND2_X1 U9778 ( .A1(n8012), .A2(n8011), .ZN(n8013) );
  NAND2_X1 U9779 ( .A1(n8015), .A2(n8014), .ZN(n8017) );
  XNOR2_X1 U9780 ( .A(n8017), .B(n8016), .ZN(n8019) );
  AND2_X1 U9781 ( .A1(n9939), .A2(n9950), .ZN(n8018) );
  NAND2_X1 U9782 ( .A1(n8019), .A2(n10373), .ZN(n8027) );
  NOR2_X4 U9783 ( .A1(n4377), .A2(n9540), .ZN(n10372) );
  INV_X2 U9784 ( .A(n10097), .ZN(n10358) );
  AOI22_X1 U9785 ( .A1(n4377), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8021), .B2(
        n10358), .ZN(n8022) );
  OAI21_X1 U9786 ( .B1(n8023), .B2(n10123), .A(n8022), .ZN(n8024) );
  AOI21_X1 U9787 ( .B1(n8025), .B2(n10372), .A(n8024), .ZN(n8026) );
  OAI211_X1 U9788 ( .C1(n8028), .C2(n4377), .A(n8027), .B(n8026), .ZN(P1_U3356) );
  INV_X1 U9789 ( .A(n8029), .ZN(n8034) );
  XNOR2_X1 U9790 ( .A(n8501), .B(n8034), .ZN(n8045) );
  INV_X1 U9791 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U9792 ( .A1(n8031), .A2(n8032), .ZN(n8033) );
  NOR2_X1 U9793 ( .A1(n8033), .A2(n8034), .ZN(n8492) );
  AOI21_X1 U9794 ( .B1(n8034), .B2(n8033), .A(n8492), .ZN(n8035) );
  OAI222_X1 U9795 ( .A1(n8558), .A2(n8483), .B1(n8694), .B2(n8214), .C1(n10469), .C2(n8035), .ZN(n8043) );
  AOI21_X1 U9796 ( .B1(n10473), .B2(n8216), .A(n8043), .ZN(n8038) );
  MUX2_X1 U9797 ( .A(n8036), .B(n8038), .S(n10501), .Z(n8037) );
  OAI21_X1 U9798 ( .B1(n8045), .B2(n8775), .A(n8037), .ZN(P2_U3447) );
  MUX2_X1 U9799 ( .A(n9132), .B(n8038), .S(n10508), .Z(n8039) );
  OAI21_X1 U9800 ( .B1(n8045), .B2(n8667), .A(n8039), .ZN(P2_U3479) );
  AOI22_X1 U9801 ( .A1(n10466), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8588), .B2(
        n8211), .ZN(n8040) );
  OAI21_X1 U9802 ( .B1(n8041), .B2(n8618), .A(n8040), .ZN(n8042) );
  AOI21_X1 U9803 ( .B1(n8043), .B2(n10464), .A(n8042), .ZN(n8044) );
  OAI21_X1 U9804 ( .B1(n8045), .B2(n8553), .A(n8044), .ZN(P2_U3213) );
  NAND2_X1 U9805 ( .A1(n8057), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U9806 ( .A1(n8047), .A2(n8046), .ZN(n10288) );
  INV_X1 U9807 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9120) );
  MUX2_X1 U9808 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n9120), .S(n10293), .Z(
        n10287) );
  NOR2_X1 U9809 ( .A1(n8048), .A2(n8062), .ZN(n8049) );
  INV_X1 U9810 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10307) );
  XOR2_X1 U9811 ( .A(n10311), .B(n8048), .Z(n10308) );
  NOR2_X1 U9812 ( .A1(n10307), .A2(n10308), .ZN(n10306) );
  NAND2_X1 U9813 ( .A1(n8064), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8050) );
  OAI21_X1 U9814 ( .B1(n8064), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8050), .ZN(
        n9689) );
  NOR2_X1 U9815 ( .A1(n9690), .A2(n9689), .ZN(n9688) );
  INV_X1 U9816 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9898) );
  XNOR2_X1 U9817 ( .A(n8066), .B(n9898), .ZN(n9696) );
  NAND2_X1 U9818 ( .A1(n9695), .A2(n9696), .ZN(n8052) );
  OR2_X1 U9819 ( .A1(n8066), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8051) );
  NAND2_X1 U9820 ( .A1(n8052), .A2(n8051), .ZN(n10318) );
  NAND2_X1 U9821 ( .A1(n8068), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8054) );
  OR2_X1 U9822 ( .A1(n8068), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8053) );
  NAND2_X1 U9823 ( .A1(n8054), .A2(n8053), .ZN(n10317) );
  NAND2_X1 U9824 ( .A1(n10327), .A2(n8054), .ZN(n8055) );
  XNOR2_X1 U9825 ( .A(n8055), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n8075) );
  INV_X1 U9826 ( .A(n8075), .ZN(n8073) );
  INV_X1 U9827 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8056) );
  AOI22_X1 U9828 ( .A1(n8064), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8056), .B2(
        n9687), .ZN(n9683) );
  NAND2_X1 U9829 ( .A1(n8057), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U9830 ( .A1(n8059), .A2(n8058), .ZN(n10290) );
  INV_X1 U9831 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8060) );
  XNOR2_X1 U9832 ( .A(n10293), .B(n8060), .ZN(n10289) );
  AND2_X1 U9833 ( .A1(n10290), .A2(n10289), .ZN(n10292) );
  AOI21_X1 U9834 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n10293), .A(n10292), .ZN(
        n8061) );
  NOR2_X1 U9835 ( .A1(n8061), .A2(n8062), .ZN(n8063) );
  INV_X1 U9836 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10304) );
  XNOR2_X1 U9837 ( .A(n8062), .B(n8061), .ZN(n10305) );
  NOR2_X1 U9838 ( .A1(n10304), .A2(n10305), .ZN(n10303) );
  NOR2_X1 U9839 ( .A1(n8063), .A2(n10303), .ZN(n9684) );
  NAND2_X1 U9840 ( .A1(n9683), .A2(n9684), .ZN(n9682) );
  OAI21_X1 U9841 ( .B1(n8064), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9682), .ZN(
        n9698) );
  INV_X1 U9842 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8065) );
  XNOR2_X1 U9843 ( .A(n8066), .B(n8065), .ZN(n9697) );
  NOR2_X1 U9844 ( .A1(n8066), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8067) );
  AOI21_X1 U9845 ( .B1(n9698), .B2(n9697), .A(n8067), .ZN(n10322) );
  OR2_X1 U9846 ( .A1(n8068), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U9847 ( .A1(n8068), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8070) );
  AND2_X1 U9848 ( .A1(n8069), .A2(n8070), .ZN(n10321) );
  NAND2_X1 U9849 ( .A1(n10322), .A2(n10321), .ZN(n10320) );
  NAND2_X1 U9850 ( .A1(n10320), .A2(n8070), .ZN(n8071) );
  XNOR2_X1 U9851 ( .A(n8071), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8074) );
  AOI21_X1 U9852 ( .B1(n8074), .B2(n10319), .A(n10312), .ZN(n8072) );
  OAI21_X1 U9853 ( .B1(n8073), .B2(n10316), .A(n8072), .ZN(n8077) );
  OAI22_X1 U9854 ( .A1(n8075), .A2(n10316), .B1(n8074), .B2(n10302), .ZN(n8076) );
  NAND2_X1 U9855 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8859) );
  OAI222_X1 U9856 ( .A1(n8804), .A2(n9073), .B1(n8811), .B2(n8079), .C1(n6214), 
        .C2(P2_U3151), .ZN(P2_U3271) );
  NAND2_X1 U9857 ( .A1(n8080), .A2(n10372), .ZN(n8083) );
  AOI22_X1 U9858 ( .A1(n4377), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8081), .B2(
        n10358), .ZN(n8082) );
  OAI211_X1 U9859 ( .C1(n8084), .C2(n10123), .A(n8083), .B(n8082), .ZN(n8085)
         );
  AOI21_X1 U9860 ( .B1(n8086), .B2(n10112), .A(n8085), .ZN(n8087) );
  OAI21_X1 U9861 ( .B1(n8088), .B2(n10124), .A(n8087), .ZN(P1_U3265) );
  XNOR2_X1 U9862 ( .A(n8090), .B(n8089), .ZN(n8091) );
  XNOR2_X1 U9863 ( .A(n8092), .B(n8091), .ZN(n8093) );
  INV_X1 U9864 ( .A(n8093), .ZN(n8097) );
  OAI211_X1 U9865 ( .C1(n8421), .C2(n8096), .A(n8097), .B(n8271), .ZN(n8101)
         );
  AOI22_X1 U9866 ( .A1(n8425), .A2(n8290), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8095) );
  NAND2_X1 U9867 ( .A1(n8440), .A2(n8286), .ZN(n8094) );
  OAI211_X1 U9868 ( .C1(n8422), .C2(n8288), .A(n8095), .B(n8094), .ZN(n8099)
         );
  NOR4_X1 U9869 ( .A1(n8097), .A2(n8421), .A3(n8096), .A4(n8281), .ZN(n8098)
         );
  AOI211_X1 U9870 ( .C1(n8263), .C2(n8711), .A(n8099), .B(n8098), .ZN(n8100)
         );
  INV_X1 U9871 ( .A(n8103), .ZN(n8812) );
  OAI222_X1 U9872 ( .A1(n8105), .A2(n8104), .B1(P1_U3086), .B2(n6095), .C1(
        n10283), .C2(n8812), .ZN(P1_U3327) );
  XOR2_X1 U9873 ( .A(n8107), .B(n8106), .Z(n8112) );
  NAND2_X1 U9874 ( .A1(n8290), .A2(n8574), .ZN(n8109) );
  INV_X1 U9875 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9079) );
  NOR2_X1 U9876 ( .A1(n9079), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8329) );
  AOI21_X1 U9877 ( .B1(n8258), .B2(n8570), .A(n8329), .ZN(n8108) );
  OAI211_X1 U9878 ( .C1(n8163), .C2(n8274), .A(n8109), .B(n8108), .ZN(n8110)
         );
  AOI21_X1 U9879 ( .B1(n8785), .B2(n8263), .A(n8110), .ZN(n8111) );
  OAI21_X1 U9880 ( .B1(n8112), .B2(n8281), .A(n8111), .ZN(P2_U3155) );
  INV_X1 U9881 ( .A(n8113), .ZN(n8115) );
  AOI21_X1 U9882 ( .B1(n8115), .B2(n8114), .A(n8197), .ZN(n8116) );
  NAND2_X1 U9883 ( .A1(n8116), .A2(n8484), .ZN(n8200) );
  OAI21_X1 U9884 ( .B1(n8484), .B2(n8116), .A(n8200), .ZN(n8117) );
  NAND2_X1 U9885 ( .A1(n8117), .A2(n8271), .ZN(n8122) );
  AOI22_X1 U9886 ( .A1(n8473), .A2(n8286), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8118) );
  OAI21_X1 U9887 ( .B1(n8119), .B2(n8288), .A(n8118), .ZN(n8120) );
  AOI21_X1 U9888 ( .B1(n8477), .B2(n8290), .A(n8120), .ZN(n8121) );
  OAI211_X1 U9889 ( .C1(n8123), .C2(n8293), .A(n8122), .B(n8121), .ZN(P2_U3156) );
  INV_X1 U9890 ( .A(n8124), .ZN(n8127) );
  XNOR2_X1 U9891 ( .A(n8125), .B(n8298), .ZN(n8126) );
  NOR2_X1 U9892 ( .A1(n8126), .A2(n8127), .ZN(n8154) );
  AOI21_X1 U9893 ( .B1(n8127), .B2(n8126), .A(n8154), .ZN(n8133) );
  OAI21_X1 U9894 ( .B1(n8288), .B2(n8157), .A(n8128), .ZN(n8129) );
  AOI21_X1 U9895 ( .B1(n8286), .B2(n8608), .A(n8129), .ZN(n8130) );
  OAI21_X1 U9896 ( .B1(n8248), .B2(n8603), .A(n8130), .ZN(n8131) );
  AOI21_X1 U9897 ( .B1(n8263), .B2(n8602), .A(n8131), .ZN(n8132) );
  OAI21_X1 U9898 ( .B1(n8133), .B2(n8281), .A(n8132), .ZN(P2_U3157) );
  XNOR2_X1 U9899 ( .A(n8134), .B(n8214), .ZN(n8135) );
  XNOR2_X1 U9900 ( .A(n8136), .B(n8135), .ZN(n8143) );
  NAND2_X1 U9901 ( .A1(n8515), .A2(n8258), .ZN(n8138) );
  OAI211_X1 U9902 ( .C1(n8139), .C2(n8274), .A(n8138), .B(n8137), .ZN(n8140)
         );
  AOI21_X1 U9903 ( .B1(n8517), .B2(n8290), .A(n8140), .ZN(n8142) );
  NAND2_X1 U9904 ( .A1(n8755), .A2(n8263), .ZN(n8141) );
  OAI211_X1 U9905 ( .C1(n8143), .C2(n8281), .A(n8142), .B(n8141), .ZN(P2_U3159) );
  INV_X1 U9906 ( .A(n8144), .ZN(n8208) );
  INV_X1 U9907 ( .A(n8145), .ZN(n8146) );
  NOR3_X1 U9908 ( .A1(n8208), .A2(n8146), .A3(n8147), .ZN(n8149) );
  AND2_X1 U9909 ( .A1(n8148), .A2(n8147), .ZN(n8234) );
  OAI21_X1 U9910 ( .B1(n8149), .B2(n8234), .A(n8271), .ZN(n8153) );
  AOI22_X1 U9911 ( .A1(n8515), .A2(n8286), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8150) );
  OAI21_X1 U9912 ( .B1(n8496), .B2(n8288), .A(n8150), .ZN(n8151) );
  AOI21_X1 U9913 ( .B1(n8498), .B2(n8290), .A(n8151), .ZN(n8152) );
  OAI211_X1 U9914 ( .C1(n8749), .C2(n8293), .A(n8153), .B(n8152), .ZN(P2_U3163) );
  INV_X1 U9915 ( .A(n8125), .ZN(n8155) );
  AOI21_X1 U9916 ( .B1(n8156), .B2(n8155), .A(n8154), .ZN(n8244) );
  XNOR2_X1 U9917 ( .A(n8158), .B(n8157), .ZN(n8243) );
  NAND2_X1 U9918 ( .A1(n8244), .A2(n8243), .ZN(n8242) );
  NAND2_X1 U9919 ( .A1(n8242), .A2(n8159), .ZN(n8160) );
  XOR2_X1 U9920 ( .A(n8161), .B(n8160), .Z(n8168) );
  OAI21_X1 U9921 ( .B1(n8288), .B2(n8163), .A(n8162), .ZN(n8164) );
  AOI21_X1 U9922 ( .B1(n8286), .B2(n8607), .A(n8164), .ZN(n8165) );
  OAI21_X1 U9923 ( .B1(n8248), .B2(n8586), .A(n8165), .ZN(n8166) );
  AOI21_X1 U9924 ( .B1(n8263), .B2(n8677), .A(n8166), .ZN(n8167) );
  OAI21_X1 U9925 ( .B1(n8168), .B2(n8281), .A(n8167), .ZN(P2_U3164) );
  INV_X1 U9926 ( .A(n8728), .ZN(n8451) );
  INV_X1 U9927 ( .A(n8169), .ZN(n8201) );
  INV_X1 U9928 ( .A(n8170), .ZN(n8172) );
  NOR3_X1 U9929 ( .A1(n8201), .A2(n8172), .A3(n8171), .ZN(n8174) );
  INV_X1 U9930 ( .A(n8173), .ZN(n8269) );
  OAI21_X1 U9931 ( .B1(n8174), .B2(n8269), .A(n8271), .ZN(n8179) );
  INV_X1 U9932 ( .A(n8175), .ZN(n8450) );
  AOI22_X1 U9933 ( .A1(n8474), .A2(n8286), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8176) );
  OAI21_X1 U9934 ( .B1(n8450), .B2(n8248), .A(n8176), .ZN(n8177) );
  AOI21_X1 U9935 ( .B1(n8258), .B2(n8448), .A(n8177), .ZN(n8178) );
  OAI211_X1 U9936 ( .C1(n8451), .C2(n8293), .A(n8179), .B(n8178), .ZN(P2_U3165) );
  AOI21_X1 U9937 ( .B1(n8180), .B2(n8189), .A(n4413), .ZN(n8186) );
  NAND2_X1 U9938 ( .A1(n8286), .A2(n8570), .ZN(n8181) );
  NAND2_X1 U9939 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8359) );
  OAI211_X1 U9940 ( .C1(n8261), .C2(n8288), .A(n8181), .B(n8359), .ZN(n8184)
         );
  NOR2_X1 U9941 ( .A1(n8182), .A2(n8293), .ZN(n8183) );
  AOI211_X1 U9942 ( .C1(n8550), .C2(n8290), .A(n8184), .B(n8183), .ZN(n8185)
         );
  OAI21_X1 U9943 ( .B1(n8186), .B2(n8281), .A(n8185), .ZN(P2_U3166) );
  INV_X1 U9944 ( .A(n8767), .ZN(n8196) );
  NOR3_X1 U9945 ( .A1(n4413), .A2(n4494), .A3(n8187), .ZN(n8191) );
  OR2_X1 U9946 ( .A1(n8189), .A2(n8188), .ZN(n8255) );
  OAI21_X1 U9947 ( .B1(n8191), .B2(n5073), .A(n8271), .ZN(n8195) );
  NAND2_X1 U9948 ( .A1(n8258), .A2(n8536), .ZN(n8192) );
  NAND2_X1 U9949 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8377) );
  OAI211_X1 U9950 ( .C1(n8274), .C2(n8557), .A(n8192), .B(n8377), .ZN(n8193)
         );
  AOI21_X1 U9951 ( .B1(n8541), .B2(n8290), .A(n8193), .ZN(n8194) );
  OAI211_X1 U9952 ( .C1(n8196), .C2(n8293), .A(n8195), .B(n8194), .ZN(P2_U3168) );
  INV_X1 U9953 ( .A(n8734), .ZN(n8207) );
  INV_X1 U9954 ( .A(n8197), .ZN(n8198) );
  AND3_X1 U9955 ( .A1(n8200), .A2(n8199), .A3(n8198), .ZN(n8202) );
  OAI21_X1 U9956 ( .B1(n8202), .B2(n8201), .A(n8271), .ZN(n8206) );
  AOI22_X1 U9957 ( .A1(n8457), .A2(n8286), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8203) );
  OAI21_X1 U9958 ( .B1(n8275), .B2(n8288), .A(n8203), .ZN(n8204) );
  AOI21_X1 U9959 ( .B1(n8460), .B2(n8290), .A(n8204), .ZN(n8205) );
  OAI211_X1 U9960 ( .C1(n8207), .C2(n8293), .A(n8206), .B(n8205), .ZN(P2_U3169) );
  AOI21_X1 U9961 ( .B1(n8210), .B2(n8209), .A(n8208), .ZN(n8218) );
  AOI22_X1 U9962 ( .A1(n8294), .A2(n8258), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8213) );
  NAND2_X1 U9963 ( .A1(n8290), .A2(n8211), .ZN(n8212) );
  OAI211_X1 U9964 ( .C1(n8214), .C2(n8274), .A(n8213), .B(n8212), .ZN(n8215)
         );
  AOI21_X1 U9965 ( .B1(n8216), .B2(n8263), .A(n8215), .ZN(n8217) );
  OAI21_X1 U9966 ( .B1(n8218), .B2(n8281), .A(n8217), .ZN(P2_U3173) );
  NAND2_X1 U9967 ( .A1(n8220), .A2(n8219), .ZN(n8222) );
  XOR2_X1 U9968 ( .A(n8222), .B(n8221), .Z(n8229) );
  NAND2_X1 U9969 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8309) );
  OAI21_X1 U9970 ( .B1(n8288), .B2(n8556), .A(n8309), .ZN(n8223) );
  AOI21_X1 U9971 ( .B1(n8286), .B2(n8297), .A(n8223), .ZN(n8224) );
  OAI21_X1 U9972 ( .B1(n8248), .B2(n8225), .A(n8224), .ZN(n8226) );
  AOI21_X1 U9973 ( .B1(n8227), .B2(n8263), .A(n8226), .ZN(n8228) );
  OAI21_X1 U9974 ( .B1(n8229), .B2(n8281), .A(n8228), .ZN(P2_U3174) );
  INV_X1 U9975 ( .A(n8230), .ZN(n8747) );
  INV_X1 U9976 ( .A(n8231), .ZN(n8233) );
  NOR3_X1 U9977 ( .A1(n8234), .A2(n8233), .A3(n8232), .ZN(n8237) );
  INV_X1 U9978 ( .A(n8235), .ZN(n8236) );
  OAI21_X1 U9979 ( .B1(n8237), .B2(n8236), .A(n8271), .ZN(n8241) );
  AOI22_X1 U9980 ( .A1(n8294), .A2(n8286), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8238) );
  OAI21_X1 U9981 ( .B1(n8484), .B2(n8288), .A(n8238), .ZN(n8239) );
  AOI21_X1 U9982 ( .B1(n8486), .B2(n8290), .A(n8239), .ZN(n8240) );
  OAI211_X1 U9983 ( .C1(n8747), .C2(n8293), .A(n8241), .B(n8240), .ZN(P2_U3175) );
  INV_X1 U9984 ( .A(n8579), .ZN(n8253) );
  OAI211_X1 U9985 ( .C1(n8244), .C2(n8243), .A(n8242), .B(n8271), .ZN(n8252)
         );
  OAI21_X1 U9986 ( .B1(n8288), .B2(n8246), .A(n8245), .ZN(n8250) );
  NOR2_X1 U9987 ( .A1(n8248), .A2(n8247), .ZN(n8249) );
  AOI211_X1 U9988 ( .C1(n8286), .C2(n8298), .A(n8250), .B(n8249), .ZN(n8251)
         );
  OAI211_X1 U9989 ( .C1(n8253), .C2(n8293), .A(n8252), .B(n8251), .ZN(P2_U3176) );
  NAND2_X1 U9990 ( .A1(n8255), .A2(n8254), .ZN(n8256) );
  XOR2_X1 U9991 ( .A(n8257), .B(n8256), .Z(n8265) );
  AND2_X1 U9992 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8409) );
  AOI21_X1 U9993 ( .B1(n8527), .B2(n8258), .A(n8409), .ZN(n8260) );
  NAND2_X1 U9994 ( .A1(n8290), .A2(n8530), .ZN(n8259) );
  OAI211_X1 U9995 ( .C1(n8261), .C2(n8274), .A(n8260), .B(n8259), .ZN(n8262)
         );
  AOI21_X1 U9996 ( .B1(n8761), .B2(n8263), .A(n8262), .ZN(n8264) );
  OAI21_X1 U9997 ( .B1(n8265), .B2(n8281), .A(n8264), .ZN(P2_U3178) );
  INV_X1 U9998 ( .A(n8266), .ZN(n8268) );
  NOR3_X1 U9999 ( .A1(n8269), .A2(n8268), .A3(n8267), .ZN(n8273) );
  INV_X1 U10000 ( .A(n8270), .ZN(n8272) );
  OAI21_X1 U10001 ( .B1(n8273), .B2(n8272), .A(n8271), .ZN(n8279) );
  OAI22_X1 U10002 ( .A1(n8275), .A2(n8274), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8970), .ZN(n8277) );
  NOR2_X1 U10003 ( .A1(n8421), .A2(n8288), .ZN(n8276) );
  AOI211_X1 U10004 ( .C1(n8442), .C2(n8290), .A(n8277), .B(n8276), .ZN(n8278)
         );
  OAI211_X1 U10005 ( .C1(n8280), .C2(n8293), .A(n8279), .B(n8278), .ZN(
        P2_U3180) );
  INV_X1 U10006 ( .A(n8779), .ZN(n8563) );
  AOI21_X1 U10007 ( .B1(n8283), .B2(n8282), .A(n8281), .ZN(n8285) );
  NAND2_X1 U10008 ( .A1(n8285), .A2(n8284), .ZN(n8292) );
  NAND2_X1 U10009 ( .A1(n8286), .A2(n8296), .ZN(n8287) );
  NAND2_X1 U10010 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8346) );
  OAI211_X1 U10011 ( .C1(n8557), .C2(n8288), .A(n8287), .B(n8346), .ZN(n8289)
         );
  AOI21_X1 U10012 ( .B1(n8290), .B2(n8559), .A(n8289), .ZN(n8291) );
  OAI211_X1 U10013 ( .C1(n8563), .C2(n8293), .A(n8292), .B(n8291), .ZN(
        P2_U3181) );
  MUX2_X1 U10014 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8432), .S(n8305), .Z(
        P2_U3519) );
  MUX2_X1 U10015 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8440), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10016 ( .A(n8448), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8402), .Z(
        P2_U3517) );
  MUX2_X1 U10017 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8458), .S(n8305), .Z(
        P2_U3516) );
  MUX2_X1 U10018 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8474), .S(n8305), .Z(
        P2_U3515) );
  MUX2_X1 U10019 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8457), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10020 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8473), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10021 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8294), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10022 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8515), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10023 ( .A(n8527), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8402), .Z(
        P2_U3510) );
  MUX2_X1 U10024 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8536), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10025 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8547), .S(P2_U3893), .Z(
        P2_U3508) );
  INV_X1 U10026 ( .A(n8557), .ZN(n8295) );
  MUX2_X1 U10027 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8295), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8570), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8296), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10030 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8583), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8297), .S(n8305), .Z(
        P2_U3503) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8607), .S(n8305), .Z(
        P2_U3502) );
  MUX2_X1 U10033 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8298), .S(n8305), .Z(
        P2_U3501) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8608), .S(n8305), .Z(
        P2_U3500) );
  MUX2_X1 U10035 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8299), .S(n8305), .Z(
        P2_U3499) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8300), .S(n8305), .Z(
        P2_U3498) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8301), .S(n8305), .Z(
        P2_U3497) );
  MUX2_X1 U10038 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8302), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10039 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8303), .S(n8305), .Z(
        P2_U3495) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n6771), .S(n8305), .Z(
        P2_U3494) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n7345), .S(n8305), .Z(
        P2_U3493) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8304), .S(n8305), .Z(
        P2_U3492) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8306), .S(n8305), .Z(
        P2_U3491) );
  AOI21_X1 U10044 ( .B1(n8308), .B2(n8307), .A(n4414), .ZN(n8321) );
  OAI21_X1 U10045 ( .B1(n8401), .B2(n4647), .A(n8309), .ZN(n8316) );
  INV_X1 U10046 ( .A(n8310), .ZN(n8311) );
  NAND3_X1 U10047 ( .A1(n8313), .A2(n8312), .A3(n8311), .ZN(n8314) );
  AOI21_X1 U10048 ( .B1(n8334), .B2(n8314), .A(n8404), .ZN(n8315) );
  AOI211_X1 U10049 ( .C1(n10443), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n8316), .B(
        n8315), .ZN(n8320) );
  XNOR2_X1 U10050 ( .A(n8317), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10051 ( .A1(n8318), .A2(n8385), .ZN(n8319) );
  OAI211_X1 U10052 ( .C1(n8321), .C2(n8389), .A(n8320), .B(n8319), .ZN(
        P2_U3195) );
  XOR2_X1 U10053 ( .A(n8323), .B(n8322), .Z(n8341) );
  INV_X1 U10054 ( .A(n8324), .ZN(n8328) );
  NOR3_X1 U10055 ( .A1(n8326), .A2(n4414), .A3(n8325), .ZN(n8327) );
  OAI21_X1 U10056 ( .B1(n8328), .B2(n8327), .A(n8396), .ZN(n8340) );
  INV_X1 U10057 ( .A(n8329), .ZN(n8330) );
  OAI21_X1 U10058 ( .B1(n8401), .B2(n8331), .A(n8330), .ZN(n8338) );
  NAND3_X1 U10059 ( .A1(n8334), .A2(n8333), .A3(n8332), .ZN(n8335) );
  AOI21_X1 U10060 ( .B1(n8336), .B2(n8335), .A(n8404), .ZN(n8337) );
  AOI211_X1 U10061 ( .C1(n10443), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8338), .B(
        n8337), .ZN(n8339) );
  OAI211_X1 U10062 ( .C1(n8341), .C2(n8411), .A(n8340), .B(n8339), .ZN(
        P2_U3196) );
  AOI21_X1 U10063 ( .B1(n8562), .B2(n8342), .A(n4394), .ZN(n8355) );
  OAI21_X1 U10064 ( .B1(n8345), .B2(n8344), .A(n8343), .ZN(n8350) );
  NAND2_X1 U10065 ( .A1(n10443), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8347) );
  OAI211_X1 U10066 ( .C1(n8401), .C2(n8348), .A(n8347), .B(n8346), .ZN(n8349)
         );
  AOI21_X1 U10067 ( .B1(n8350), .B2(n10452), .A(n8349), .ZN(n8354) );
  OAI21_X1 U10068 ( .B1(n8351), .B2(P2_REG1_REG_15__SCAN_IN), .A(n8369), .ZN(
        n8352) );
  NAND2_X1 U10069 ( .A1(n8352), .A2(n8385), .ZN(n8353) );
  OAI211_X1 U10070 ( .C1(n8355), .C2(n8389), .A(n8354), .B(n8353), .ZN(
        P2_U3197) );
  NOR3_X1 U10071 ( .A1(n4394), .A2(n8357), .A3(n8356), .ZN(n8358) );
  OAI21_X1 U10072 ( .B1(n4448), .B2(n8358), .A(n8396), .ZN(n8375) );
  OAI21_X1 U10073 ( .B1(n8401), .B2(n8360), .A(n8359), .ZN(n8367) );
  NAND2_X1 U10074 ( .A1(n8362), .A2(n8361), .ZN(n8363) );
  XNOR2_X1 U10075 ( .A(n8364), .B(n8363), .ZN(n8365) );
  NOR2_X1 U10076 ( .A1(n8365), .A2(n8404), .ZN(n8366) );
  AOI211_X1 U10077 ( .C1(n10443), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n8367), .B(
        n8366), .ZN(n8374) );
  AND3_X1 U10078 ( .A1(n8370), .A2(n8369), .A3(n8368), .ZN(n8371) );
  OAI21_X1 U10079 ( .B1(n8372), .B2(n8371), .A(n8385), .ZN(n8373) );
  NAND3_X1 U10080 ( .A1(n8375), .A2(n8374), .A3(n8373), .ZN(P2_U3198) );
  AOI21_X1 U10081 ( .B1(n8540), .B2(n8376), .A(n8395), .ZN(n8390) );
  OAI21_X1 U10082 ( .B1(n8401), .B2(n8378), .A(n8377), .ZN(n8383) );
  XOR2_X1 U10083 ( .A(n8380), .B(n8379), .Z(n8381) );
  NOR2_X1 U10084 ( .A1(n8381), .A2(n8404), .ZN(n8382) );
  AOI211_X1 U10085 ( .C1(n10443), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8383), .B(
        n8382), .ZN(n8388) );
  XOR2_X1 U10086 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8384), .Z(n8386) );
  NAND2_X1 U10087 ( .A1(n8386), .A2(n8385), .ZN(n8387) );
  OAI211_X1 U10088 ( .C1(n8390), .C2(n8389), .A(n8388), .B(n8387), .ZN(
        P2_U3199) );
  NOR3_X1 U10089 ( .A1(n8395), .A2(n8394), .A3(n8393), .ZN(n8397) );
  INV_X1 U10090 ( .A(n8398), .ZN(n8399) );
  INV_X1 U10091 ( .A(n8405), .ZN(n8403) );
  OAI21_X1 U10092 ( .B1(n8403), .B2(n8402), .A(n8401), .ZN(n8407) );
  AOI211_X1 U10093 ( .C1(n10443), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8409), .B(
        n8408), .ZN(n8410) );
  NAND2_X1 U10094 ( .A1(n8703), .A2(n8589), .ZN(n8415) );
  AOI21_X1 U10095 ( .B1(n8704), .B2(n10464), .A(n8414), .ZN(n8417) );
  OAI211_X1 U10096 ( .C1(n10464), .C2(n9066), .A(n8415), .B(n8417), .ZN(
        P2_U3202) );
  NAND2_X1 U10097 ( .A1(n10466), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8416) );
  OAI211_X1 U10098 ( .C1(n8709), .C2(n8618), .A(n8417), .B(n8416), .ZN(
        P2_U3203) );
  XNOR2_X1 U10099 ( .A(n8418), .B(n8420), .ZN(n8714) );
  XNOR2_X1 U10100 ( .A(n8419), .B(n8420), .ZN(n8424) );
  OAI22_X1 U10101 ( .A1(n8422), .A2(n8558), .B1(n8421), .B2(n8694), .ZN(n8423)
         );
  AOI21_X1 U10102 ( .B1(n8424), .B2(n8696), .A(n8423), .ZN(n8710) );
  MUX2_X1 U10103 ( .A(n8932), .B(n8710), .S(n10464), .Z(n8427) );
  AOI22_X1 U10104 ( .A1(n8711), .A2(n8589), .B1(n8588), .B2(n8425), .ZN(n8426)
         );
  OAI211_X1 U10105 ( .C1(n8714), .C2(n8553), .A(n8427), .B(n8426), .ZN(
        P2_U3205) );
  XNOR2_X1 U10106 ( .A(n8428), .B(n8429), .ZN(n8720) );
  INV_X1 U10107 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8433) );
  MUX2_X1 U10108 ( .A(n8433), .B(n8715), .S(n10464), .Z(n8436) );
  AOI22_X1 U10109 ( .A1(n8717), .A2(n8589), .B1(n8588), .B2(n8434), .ZN(n8435)
         );
  OAI211_X1 U10110 ( .C1(n8720), .C2(n8553), .A(n8436), .B(n8435), .ZN(
        P2_U3206) );
  XNOR2_X1 U10111 ( .A(n8437), .B(n8438), .ZN(n8725) );
  MUX2_X1 U10112 ( .A(n8441), .B(n8721), .S(n10464), .Z(n8444) );
  AOI22_X1 U10113 ( .A1(n8722), .A2(n8589), .B1(n8588), .B2(n8442), .ZN(n8443)
         );
  OAI211_X1 U10114 ( .C1(n8725), .C2(n8553), .A(n8444), .B(n8443), .ZN(
        P2_U3207) );
  XOR2_X1 U10115 ( .A(n8445), .B(n8447), .Z(n8731) );
  XNOR2_X1 U10116 ( .A(n8446), .B(n8447), .ZN(n8449) );
  AOI222_X1 U10117 ( .A1(n8696), .A2(n8449), .B1(n8474), .B2(n8609), .C1(n8448), .C2(n8692), .ZN(n8726) );
  INV_X1 U10118 ( .A(n8726), .ZN(n8453) );
  OAI22_X1 U10119 ( .A1(n8451), .A2(n8567), .B1(n8450), .B2(n10458), .ZN(n8452) );
  OAI21_X1 U10120 ( .B1(n8453), .B2(n8452), .A(n10464), .ZN(n8455) );
  NAND2_X1 U10121 ( .A1(n10466), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8454) );
  OAI211_X1 U10122 ( .C1(n8731), .C2(n8553), .A(n8455), .B(n8454), .ZN(
        P2_U3208) );
  XOR2_X1 U10123 ( .A(n8465), .B(n8456), .Z(n8459) );
  AOI222_X1 U10124 ( .A1(n8696), .A2(n8459), .B1(n8458), .B2(n8692), .C1(n8457), .C2(n8609), .ZN(n8732) );
  AOI22_X1 U10125 ( .A1(n8734), .A2(n8461), .B1(n8588), .B2(n8460), .ZN(n8462)
         );
  AOI21_X1 U10126 ( .B1(n8732), .B2(n8462), .A(n10466), .ZN(n8469) );
  NAND2_X1 U10127 ( .A1(n8464), .A2(n8463), .ZN(n8466) );
  XNOR2_X1 U10128 ( .A(n8466), .B(n8465), .ZN(n8737) );
  OAI22_X1 U10129 ( .A1(n8737), .A2(n8553), .B1(n8467), .B2(n10464), .ZN(n8468) );
  OR2_X1 U10130 ( .A1(n8469), .A2(n8468), .ZN(P2_U3209) );
  XNOR2_X1 U10131 ( .A(n8470), .B(n8472), .ZN(n8743) );
  INV_X1 U10132 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8476) );
  XNOR2_X1 U10133 ( .A(n8471), .B(n8472), .ZN(n8475) );
  AOI222_X1 U10134 ( .A1(n8696), .A2(n8475), .B1(n8474), .B2(n8692), .C1(n8473), .C2(n8609), .ZN(n8738) );
  MUX2_X1 U10135 ( .A(n8476), .B(n8738), .S(n10464), .Z(n8479) );
  AOI22_X1 U10136 ( .A1(n8740), .A2(n8589), .B1(n8588), .B2(n8477), .ZN(n8478)
         );
  OAI211_X1 U10137 ( .C1(n8743), .C2(n8553), .A(n8479), .B(n8478), .ZN(
        P2_U3210) );
  XNOR2_X1 U10138 ( .A(n8480), .B(n8481), .ZN(n8482) );
  OAI222_X1 U10139 ( .A1(n8558), .A2(n8484), .B1(n8694), .B2(n8483), .C1(n8482), .C2(n10469), .ZN(n8648) );
  INV_X1 U10140 ( .A(n8648), .ZN(n8490) );
  XNOR2_X1 U10141 ( .A(n4446), .B(n8485), .ZN(n8649) );
  AOI22_X1 U10142 ( .A1(n10466), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8486), 
        .B2(n8588), .ZN(n8487) );
  OAI21_X1 U10143 ( .B1(n8747), .B2(n8618), .A(n8487), .ZN(n8488) );
  AOI21_X1 U10144 ( .B1(n8649), .B2(n8593), .A(n8488), .ZN(n8489) );
  OAI21_X1 U10145 ( .B1(n8490), .B2(n10466), .A(n8489), .ZN(P2_U3211) );
  NOR2_X1 U10146 ( .A1(n8492), .A2(n8491), .ZN(n8494) );
  XNOR2_X1 U10147 ( .A(n8494), .B(n8493), .ZN(n8495) );
  OAI222_X1 U10148 ( .A1(n8694), .A2(n8497), .B1(n8558), .B2(n8496), .C1(
        n10469), .C2(n8495), .ZN(n8748) );
  AOI21_X1 U10149 ( .B1(n8588), .B2(n8498), .A(n8748), .ZN(n8508) );
  AOI22_X1 U10150 ( .A1(n8499), .A2(n8589), .B1(P2_REG2_REG_21__SCAN_IN), .B2(
        n10466), .ZN(n8507) );
  OR2_X1 U10151 ( .A1(n8501), .A2(n8500), .ZN(n8503) );
  NAND2_X1 U10152 ( .A1(n8503), .A2(n8502), .ZN(n8505) );
  XNOR2_X1 U10153 ( .A(n8505), .B(n8504), .ZN(n8652) );
  NAND2_X1 U10154 ( .A1(n8652), .A2(n8593), .ZN(n8506) );
  OAI211_X1 U10155 ( .C1(n8508), .C2(n10466), .A(n8507), .B(n8506), .ZN(
        P2_U3212) );
  XNOR2_X1 U10156 ( .A(n4669), .B(n8509), .ZN(n8758) );
  INV_X1 U10157 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8516) );
  AND2_X1 U10158 ( .A1(n8536), .A2(n8609), .ZN(n8514) );
  INV_X1 U10159 ( .A(n8031), .ZN(n8510) );
  AOI211_X1 U10160 ( .C1(n8512), .C2(n8511), .A(n10469), .B(n8510), .ZN(n8513)
         );
  AOI211_X1 U10161 ( .C1(n8692), .C2(n8515), .A(n8514), .B(n8513), .ZN(n8753)
         );
  MUX2_X1 U10162 ( .A(n8516), .B(n8753), .S(n10464), .Z(n8519) );
  AOI22_X1 U10163 ( .A1(n8755), .A2(n8589), .B1(n8588), .B2(n8517), .ZN(n8518)
         );
  OAI211_X1 U10164 ( .C1(n8758), .C2(n8553), .A(n8519), .B(n8518), .ZN(
        P2_U3214) );
  NAND2_X1 U10165 ( .A1(n8521), .A2(n8520), .ZN(n8526) );
  NAND2_X1 U10166 ( .A1(n8523), .A2(n8522), .ZN(n8524) );
  XOR2_X1 U10167 ( .A(n8526), .B(n8524), .Z(n8764) );
  XOR2_X1 U10168 ( .A(n8526), .B(n8525), .Z(n8528) );
  AOI222_X1 U10169 ( .A1(n8696), .A2(n8528), .B1(n8527), .B2(n8692), .C1(n8547), .C2(n8609), .ZN(n8759) );
  MUX2_X1 U10170 ( .A(n8529), .B(n8759), .S(n10464), .Z(n8532) );
  AOI22_X1 U10171 ( .A1(n8761), .A2(n8589), .B1(n8588), .B2(n8530), .ZN(n8531)
         );
  OAI211_X1 U10172 ( .C1(n8764), .C2(n8553), .A(n8532), .B(n8531), .ZN(
        P2_U3215) );
  XNOR2_X1 U10173 ( .A(n8533), .B(n8534), .ZN(n8770) );
  XNOR2_X1 U10174 ( .A(n8535), .B(n8534), .ZN(n8539) );
  NAND2_X1 U10175 ( .A1(n8536), .A2(n8692), .ZN(n8537) );
  OAI21_X1 U10176 ( .B1(n8557), .B2(n8694), .A(n8537), .ZN(n8538) );
  AOI21_X1 U10177 ( .B1(n8539), .B2(n8696), .A(n8538), .ZN(n8765) );
  MUX2_X1 U10178 ( .A(n8540), .B(n8765), .S(n10464), .Z(n8543) );
  AOI22_X1 U10179 ( .A1(n8767), .A2(n8589), .B1(n8588), .B2(n8541), .ZN(n8542)
         );
  OAI211_X1 U10180 ( .C1(n8770), .C2(n8553), .A(n8543), .B(n8542), .ZN(
        P2_U3216) );
  XNOR2_X1 U10181 ( .A(n8544), .B(n8545), .ZN(n8776) );
  XOR2_X1 U10182 ( .A(n8546), .B(n8545), .Z(n8548) );
  AOI222_X1 U10183 ( .A1(n8696), .A2(n8548), .B1(n8547), .B2(n8692), .C1(n8570), .C2(n8609), .ZN(n8771) );
  MUX2_X1 U10184 ( .A(n8549), .B(n8771), .S(n10464), .Z(n8552) );
  AOI22_X1 U10185 ( .A1(n8772), .A2(n8589), .B1(n8588), .B2(n8550), .ZN(n8551)
         );
  OAI211_X1 U10186 ( .C1(n8776), .C2(n8553), .A(n8552), .B(n8551), .ZN(
        P2_U3217) );
  XNOR2_X1 U10187 ( .A(n8554), .B(n8560), .ZN(n8555) );
  OAI222_X1 U10188 ( .A1(n8558), .A2(n8557), .B1(n8694), .B2(n8556), .C1(
        n10469), .C2(n8555), .ZN(n8668) );
  AOI21_X1 U10189 ( .B1(n8588), .B2(n8559), .A(n8668), .ZN(n8566) );
  XNOR2_X1 U10190 ( .A(n8561), .B(n8560), .ZN(n8780) );
  OAI22_X1 U10191 ( .A1(n8563), .A2(n8618), .B1(n8562), .B2(n10464), .ZN(n8564) );
  AOI21_X1 U10192 ( .B1(n8780), .B2(n8593), .A(n8564), .ZN(n8565) );
  OAI21_X1 U10193 ( .B1(n8566), .B2(n10466), .A(n8565), .ZN(P2_U3218) );
  INV_X1 U10194 ( .A(n8785), .ZN(n8568) );
  NOR2_X1 U10195 ( .A1(n8568), .A2(n8567), .ZN(n8573) );
  XNOR2_X1 U10196 ( .A(n8569), .B(n8575), .ZN(n8571) );
  AOI222_X1 U10197 ( .A1(n8696), .A2(n8571), .B1(n8570), .B2(n8692), .C1(n8583), .C2(n8609), .ZN(n8783) );
  INV_X1 U10198 ( .A(n8783), .ZN(n8572) );
  AOI211_X1 U10199 ( .C1(n8588), .C2(n8574), .A(n8573), .B(n8572), .ZN(n8578)
         );
  XOR2_X1 U10200 ( .A(n8576), .B(n8575), .Z(n8787) );
  AOI22_X1 U10201 ( .A1(n8787), .A2(n8593), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n10466), .ZN(n8577) );
  OAI21_X1 U10202 ( .B1(n8578), .B2(n10466), .A(n8577), .ZN(P2_U3219) );
  AOI22_X1 U10203 ( .A1(n8581), .A2(n8580), .B1(n8607), .B2(n8579), .ZN(n8582)
         );
  XNOR2_X1 U10204 ( .A(n8582), .B(n8591), .ZN(n8584) );
  AOI222_X1 U10205 ( .A1(n8696), .A2(n8584), .B1(n8583), .B2(n8692), .C1(n8607), .C2(n8609), .ZN(n8680) );
  MUX2_X1 U10206 ( .A(n8585), .B(n8680), .S(n10464), .Z(n8596) );
  INV_X1 U10207 ( .A(n8586), .ZN(n8587) );
  AOI22_X1 U10208 ( .A1(n8677), .A2(n8589), .B1(n8588), .B2(n8587), .ZN(n8595)
         );
  NAND2_X1 U10209 ( .A1(n8592), .A2(n8591), .ZN(n8678) );
  NAND3_X1 U10210 ( .A1(n8590), .A2(n8678), .A3(n8593), .ZN(n8594) );
  NAND3_X1 U10211 ( .A1(n8596), .A2(n8595), .A3(n8594), .ZN(P2_U3221) );
  NAND2_X1 U10212 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U10213 ( .A1(n8599), .A2(n8604), .ZN(n8601) );
  NAND2_X1 U10214 ( .A1(n8601), .A2(n8600), .ZN(n8683) );
  INV_X1 U10215 ( .A(n8602), .ZN(n8794) );
  OAI22_X1 U10216 ( .A1(n8618), .A2(n8794), .B1(n8603), .B2(n10458), .ZN(n8614) );
  XNOR2_X1 U10217 ( .A(n8605), .B(n8604), .ZN(n8606) );
  NAND2_X1 U10218 ( .A1(n8606), .A2(n8696), .ZN(n8612) );
  AOI22_X1 U10219 ( .A1(n8609), .A2(n8608), .B1(n8607), .B2(n8692), .ZN(n8611)
         );
  NAND2_X1 U10220 ( .A1(n8683), .A2(n8689), .ZN(n8610) );
  NAND3_X1 U10221 ( .A1(n8612), .A2(n8611), .A3(n8610), .ZN(n8682) );
  MUX2_X1 U10222 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8682), .S(n10464), .Z(
        n8613) );
  AOI211_X1 U10223 ( .C1(n8622), .C2(n8683), .A(n8614), .B(n8613), .ZN(n8615)
         );
  INV_X1 U10224 ( .A(n8615), .ZN(P2_U3223) );
  OAI22_X1 U10225 ( .A1(n8618), .A2(n8617), .B1(n8616), .B2(n10458), .ZN(n8621) );
  MUX2_X1 U10226 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8619), .S(n10464), .Z(n8620) );
  AOI211_X1 U10227 ( .C1(n8623), .C2(n8622), .A(n8621), .B(n8620), .ZN(n8624)
         );
  INV_X1 U10228 ( .A(n8624), .ZN(P2_U3224) );
  NAND2_X1 U10229 ( .A1(n8703), .A2(n8673), .ZN(n8625) );
  NAND2_X1 U10230 ( .A1(n8704), .A2(n10508), .ZN(n8628) );
  OAI211_X1 U10231 ( .C1(n10508), .C2(n8626), .A(n8625), .B(n8628), .ZN(
        P2_U3490) );
  NAND2_X1 U10232 ( .A1(n8627), .A2(n8673), .ZN(n8629) );
  OAI211_X1 U10233 ( .C1(n10508), .C2(n8630), .A(n8629), .B(n8628), .ZN(
        P2_U3489) );
  INV_X1 U10234 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8631) );
  MUX2_X1 U10235 ( .A(n8631), .B(n8710), .S(n10508), .Z(n8633) );
  NAND2_X1 U10236 ( .A1(n8711), .A2(n8673), .ZN(n8632) );
  OAI211_X1 U10237 ( .C1(n8714), .C2(n8667), .A(n8633), .B(n8632), .ZN(
        P2_U3487) );
  MUX2_X1 U10238 ( .A(n8634), .B(n8715), .S(n10508), .Z(n8636) );
  NAND2_X1 U10239 ( .A1(n8717), .A2(n8673), .ZN(n8635) );
  OAI211_X1 U10240 ( .C1(n8720), .C2(n8667), .A(n8636), .B(n8635), .ZN(
        P2_U3486) );
  INV_X1 U10241 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8637) );
  MUX2_X1 U10242 ( .A(n8637), .B(n8721), .S(n10508), .Z(n8639) );
  NAND2_X1 U10243 ( .A1(n8722), .A2(n8673), .ZN(n8638) );
  OAI211_X1 U10244 ( .C1(n8667), .C2(n8725), .A(n8639), .B(n8638), .ZN(
        P2_U3485) );
  MUX2_X1 U10245 ( .A(n8640), .B(n8726), .S(n10508), .Z(n8642) );
  NAND2_X1 U10246 ( .A1(n8728), .A2(n8673), .ZN(n8641) );
  OAI211_X1 U10247 ( .C1(n8731), .C2(n8667), .A(n8642), .B(n8641), .ZN(
        P2_U3484) );
  MUX2_X1 U10248 ( .A(n9056), .B(n8732), .S(n10508), .Z(n8644) );
  NAND2_X1 U10249 ( .A1(n8734), .A2(n8673), .ZN(n8643) );
  OAI211_X1 U10250 ( .C1(n8667), .C2(n8737), .A(n8644), .B(n8643), .ZN(
        P2_U3483) );
  MUX2_X1 U10251 ( .A(n8645), .B(n8738), .S(n10508), .Z(n8647) );
  NAND2_X1 U10252 ( .A1(n8740), .A2(n8673), .ZN(n8646) );
  OAI211_X1 U10253 ( .C1(n8743), .C2(n8667), .A(n8647), .B(n8646), .ZN(
        P2_U3482) );
  INV_X1 U10254 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8650) );
  AOI21_X1 U10255 ( .B1(n8649), .B2(n10487), .A(n8648), .ZN(n8744) );
  MUX2_X1 U10256 ( .A(n8650), .B(n8744), .S(n10508), .Z(n8651) );
  OAI21_X1 U10257 ( .B1(n8747), .B2(n8686), .A(n8651), .ZN(P2_U3481) );
  MUX2_X1 U10258 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8748), .S(n10508), .Z(
        n8654) );
  INV_X1 U10259 ( .A(n8652), .ZN(n8750) );
  OAI22_X1 U10260 ( .A1(n8750), .A2(n8667), .B1(n8749), .B2(n8686), .ZN(n8653)
         );
  OR2_X1 U10261 ( .A1(n8654), .A2(n8653), .ZN(P2_U3480) );
  MUX2_X1 U10262 ( .A(n8655), .B(n8753), .S(n10508), .Z(n8657) );
  NAND2_X1 U10263 ( .A1(n8755), .A2(n8673), .ZN(n8656) );
  OAI211_X1 U10264 ( .C1(n8667), .C2(n8758), .A(n8657), .B(n8656), .ZN(
        P2_U3478) );
  INV_X1 U10265 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8658) );
  MUX2_X1 U10266 ( .A(n8658), .B(n8759), .S(n10508), .Z(n8660) );
  NAND2_X1 U10267 ( .A1(n8761), .A2(n8673), .ZN(n8659) );
  OAI211_X1 U10268 ( .C1(n8764), .C2(n8667), .A(n8660), .B(n8659), .ZN(
        P2_U3477) );
  MUX2_X1 U10269 ( .A(n8661), .B(n8765), .S(n10508), .Z(n8663) );
  NAND2_X1 U10270 ( .A1(n8767), .A2(n8673), .ZN(n8662) );
  OAI211_X1 U10271 ( .C1(n8770), .C2(n8667), .A(n8663), .B(n8662), .ZN(
        P2_U3476) );
  MUX2_X1 U10272 ( .A(n8664), .B(n8771), .S(n10508), .Z(n8666) );
  NAND2_X1 U10273 ( .A1(n8772), .A2(n8673), .ZN(n8665) );
  OAI211_X1 U10274 ( .C1(n8776), .C2(n8667), .A(n8666), .B(n8665), .ZN(
        P2_U3475) );
  INV_X1 U10275 ( .A(n8668), .ZN(n8777) );
  MUX2_X1 U10276 ( .A(n8669), .B(n8777), .S(n10508), .Z(n8671) );
  AOI22_X1 U10277 ( .A1(n8780), .A2(n8674), .B1(n8673), .B2(n8779), .ZN(n8670)
         );
  NAND2_X1 U10278 ( .A1(n8671), .A2(n8670), .ZN(P2_U3474) );
  MUX2_X1 U10279 ( .A(n8672), .B(n8783), .S(n10508), .Z(n8676) );
  AOI22_X1 U10280 ( .A1(n8787), .A2(n8674), .B1(n8673), .B2(n8785), .ZN(n8675)
         );
  NAND2_X1 U10281 ( .A1(n8676), .A2(n8675), .ZN(P2_U3473) );
  INV_X1 U10282 ( .A(n8677), .ZN(n8681) );
  NAND3_X1 U10283 ( .A1(n8590), .A2(n8678), .A3(n10487), .ZN(n8679) );
  OAI211_X1 U10284 ( .C1(n8681), .C2(n10488), .A(n8680), .B(n8679), .ZN(n8790)
         );
  MUX2_X1 U10285 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8790), .S(n10508), .Z(
        P2_U3471) );
  AOI21_X1 U10286 ( .B1(n10493), .B2(n8683), .A(n8682), .ZN(n8791) );
  MUX2_X1 U10287 ( .A(n8684), .B(n8791), .S(n10508), .Z(n8685) );
  OAI21_X1 U10288 ( .B1(n8794), .B2(n8686), .A(n8685), .ZN(P2_U3469) );
  XNOR2_X1 U10289 ( .A(n8688), .B(n8687), .ZN(n10462) );
  NAND2_X1 U10290 ( .A1(n10462), .A2(n8689), .ZN(n8699) );
  XNOR2_X1 U10291 ( .A(n8691), .B(n8690), .ZN(n8697) );
  NAND2_X1 U10292 ( .A1(n6771), .A2(n8692), .ZN(n8693) );
  OAI21_X1 U10293 ( .B1(n6150), .B2(n8694), .A(n8693), .ZN(n8695) );
  AOI21_X1 U10294 ( .B1(n8697), .B2(n8696), .A(n8695), .ZN(n8698) );
  AND2_X1 U10295 ( .A1(n8699), .A2(n8698), .ZN(n10459) );
  AOI21_X1 U10296 ( .B1(n10462), .B2(n10493), .A(n8700), .ZN(n8701) );
  AND2_X1 U10297 ( .A1(n10459), .A2(n8701), .ZN(n10476) );
  INV_X1 U10298 ( .A(n10476), .ZN(n8702) );
  MUX2_X1 U10299 ( .A(n8702), .B(P2_REG1_REG_2__SCAN_IN), .S(n7125), .Z(
        P2_U3461) );
  INV_X1 U10300 ( .A(n8703), .ZN(n8706) );
  NAND2_X1 U10301 ( .A1(n10499), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U10302 ( .A1(n8704), .A2(n10501), .ZN(n8708) );
  OAI211_X1 U10303 ( .C1(n8706), .C2(n8793), .A(n8705), .B(n8708), .ZN(
        P2_U3458) );
  NAND2_X1 U10304 ( .A1(n10499), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8707) );
  OAI211_X1 U10305 ( .C1(n8709), .C2(n8793), .A(n8708), .B(n8707), .ZN(
        P2_U3457) );
  MUX2_X1 U10306 ( .A(n9054), .B(n8710), .S(n10501), .Z(n8713) );
  NAND2_X1 U10307 ( .A1(n8711), .A2(n6752), .ZN(n8712) );
  OAI211_X1 U10308 ( .C1(n8714), .C2(n8775), .A(n8713), .B(n8712), .ZN(
        P2_U3455) );
  INV_X1 U10309 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8716) );
  MUX2_X1 U10310 ( .A(n8716), .B(n8715), .S(n10501), .Z(n8719) );
  NAND2_X1 U10311 ( .A1(n8717), .A2(n6752), .ZN(n8718) );
  OAI211_X1 U10312 ( .C1(n8720), .C2(n8775), .A(n8719), .B(n8718), .ZN(
        P2_U3454) );
  MUX2_X1 U10313 ( .A(n9109), .B(n8721), .S(n10501), .Z(n8724) );
  NAND2_X1 U10314 ( .A1(n8722), .A2(n6752), .ZN(n8723) );
  OAI211_X1 U10315 ( .C1(n8725), .C2(n8775), .A(n8724), .B(n8723), .ZN(
        P2_U3453) );
  INV_X1 U10316 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8727) );
  MUX2_X1 U10317 ( .A(n8727), .B(n8726), .S(n10501), .Z(n8730) );
  NAND2_X1 U10318 ( .A1(n8728), .A2(n6752), .ZN(n8729) );
  OAI211_X1 U10319 ( .C1(n8731), .C2(n8775), .A(n8730), .B(n8729), .ZN(
        P2_U3452) );
  INV_X1 U10320 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8733) );
  MUX2_X1 U10321 ( .A(n8733), .B(n8732), .S(n10501), .Z(n8736) );
  NAND2_X1 U10322 ( .A1(n8734), .A2(n6752), .ZN(n8735) );
  OAI211_X1 U10323 ( .C1(n8737), .C2(n8775), .A(n8736), .B(n8735), .ZN(
        P2_U3451) );
  INV_X1 U10324 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8739) );
  MUX2_X1 U10325 ( .A(n8739), .B(n8738), .S(n10501), .Z(n8742) );
  NAND2_X1 U10326 ( .A1(n8740), .A2(n6752), .ZN(n8741) );
  OAI211_X1 U10327 ( .C1(n8743), .C2(n8775), .A(n8742), .B(n8741), .ZN(
        P2_U3450) );
  MUX2_X1 U10328 ( .A(n8745), .B(n8744), .S(n10501), .Z(n8746) );
  OAI21_X1 U10329 ( .B1(n8747), .B2(n8793), .A(n8746), .ZN(P2_U3449) );
  MUX2_X1 U10330 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8748), .S(n10501), .Z(
        n8752) );
  OAI22_X1 U10331 ( .A1(n8750), .A2(n8775), .B1(n8749), .B2(n8793), .ZN(n8751)
         );
  OR2_X1 U10332 ( .A1(n8752), .A2(n8751), .ZN(P2_U3448) );
  INV_X1 U10333 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8754) );
  MUX2_X1 U10334 ( .A(n8754), .B(n8753), .S(n10501), .Z(n8757) );
  NAND2_X1 U10335 ( .A1(n8755), .A2(n6752), .ZN(n8756) );
  OAI211_X1 U10336 ( .C1(n8758), .C2(n8775), .A(n8757), .B(n8756), .ZN(
        P2_U3446) );
  INV_X1 U10337 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8760) );
  MUX2_X1 U10338 ( .A(n8760), .B(n8759), .S(n10501), .Z(n8763) );
  NAND2_X1 U10339 ( .A1(n8761), .A2(n6752), .ZN(n8762) );
  OAI211_X1 U10340 ( .C1(n8764), .C2(n8775), .A(n8763), .B(n8762), .ZN(
        P2_U3444) );
  INV_X1 U10341 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8766) );
  MUX2_X1 U10342 ( .A(n8766), .B(n8765), .S(n10501), .Z(n8769) );
  NAND2_X1 U10343 ( .A1(n8767), .A2(n6752), .ZN(n8768) );
  OAI211_X1 U10344 ( .C1(n8770), .C2(n8775), .A(n8769), .B(n8768), .ZN(
        P2_U3441) );
  INV_X1 U10345 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9103) );
  MUX2_X1 U10346 ( .A(n9103), .B(n8771), .S(n10501), .Z(n8774) );
  NAND2_X1 U10347 ( .A1(n8772), .A2(n6752), .ZN(n8773) );
  OAI211_X1 U10348 ( .C1(n8776), .C2(n8775), .A(n8774), .B(n8773), .ZN(
        P2_U3438) );
  MUX2_X1 U10349 ( .A(n8778), .B(n8777), .S(n10501), .Z(n8782) );
  AOI22_X1 U10350 ( .A1(n8780), .A2(n8786), .B1(n6752), .B2(n8779), .ZN(n8781)
         );
  NAND2_X1 U10351 ( .A1(n8782), .A2(n8781), .ZN(P2_U3435) );
  INV_X1 U10352 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8784) );
  MUX2_X1 U10353 ( .A(n8784), .B(n8783), .S(n10501), .Z(n8789) );
  AOI22_X1 U10354 ( .A1(n8787), .A2(n8786), .B1(n6752), .B2(n8785), .ZN(n8788)
         );
  NAND2_X1 U10355 ( .A1(n8789), .A2(n8788), .ZN(P2_U3432) );
  MUX2_X1 U10356 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8790), .S(n10501), .Z(
        P2_U3426) );
  MUX2_X1 U10357 ( .A(n8923), .B(n8791), .S(n10501), .Z(n8792) );
  OAI21_X1 U10358 ( .B1(n8794), .B2(n8793), .A(n8792), .ZN(P2_U3420) );
  MUX2_X1 U10359 ( .A(n8796), .B(P2_D_REG_1__SCAN_IN), .S(n8795), .Z(P2_U3377)
         );
  INV_X1 U10360 ( .A(n8797), .ZN(n10284) );
  NOR4_X1 U10361 ( .A1(n8798), .A2(P2_IR_REG_30__SCAN_IN), .A3(n4859), .A4(
        P2_U3151), .ZN(n8799) );
  AOI21_X1 U10362 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n8809), .A(n8799), .ZN(
        n8800) );
  OAI21_X1 U10363 ( .B1(n10284), .B2(n8811), .A(n8800), .ZN(P2_U3264) );
  AOI22_X1 U10364 ( .A1(n5206), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8809), .ZN(n8802) );
  OAI21_X1 U10365 ( .B1(n8803), .B2(n8811), .A(n8802), .ZN(P2_U3265) );
  INV_X1 U10366 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8805) );
  OAI222_X1 U10367 ( .A1(n8807), .A2(P2_U3151), .B1(n8811), .B2(n8806), .C1(
        n8805), .C2(n8804), .ZN(P2_U3266) );
  AOI21_X1 U10368 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n8809), .A(n8808), .ZN(
        n8810) );
  OAI21_X1 U10369 ( .B1(n8812), .B2(n8811), .A(n8810), .ZN(P2_U3267) );
  MUX2_X1 U10370 ( .A(n8813), .B(n10448), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3295) );
  AOI21_X1 U10371 ( .B1(n9286), .B2(n8815), .A(n8814), .ZN(n8817) );
  OAI21_X1 U10372 ( .B1(n8817), .B2(n8816), .A(n9287), .ZN(n8824) );
  NOR2_X1 U10373 ( .A1(n9301), .A2(n8818), .ZN(n8820) );
  OAI22_X1 U10374 ( .A1(n9277), .A2(n9402), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8935), .ZN(n8819) );
  AOI211_X1 U10375 ( .C1(n9719), .C2(n9305), .A(n8820), .B(n8819), .ZN(n8823)
         );
  NAND2_X1 U10376 ( .A1(n8821), .A2(n9256), .ZN(n8822) );
  NAND3_X1 U10377 ( .A1(n8824), .A2(n8823), .A3(n8822), .ZN(P1_U3214) );
  NAND2_X1 U10378 ( .A1(n8825), .A2(n5059), .ZN(n8827) );
  XNOR2_X1 U10379 ( .A(n8827), .B(n8826), .ZN(n8832) );
  NAND2_X1 U10380 ( .A1(n9299), .A2(n9565), .ZN(n8828) );
  NAND2_X1 U10381 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10299)
         );
  OAI211_X1 U10382 ( .C1(n9942), .C2(n9301), .A(n8828), .B(n10299), .ZN(n8830)
         );
  INV_X1 U10383 ( .A(n9955), .ZN(n10213) );
  NOR2_X1 U10384 ( .A1(n10213), .A2(n9302), .ZN(n8829) );
  AOI211_X1 U10385 ( .C1(n9954), .C2(n9305), .A(n8830), .B(n8829), .ZN(n8831)
         );
  OAI21_X1 U10386 ( .B1(n8832), .B2(n9307), .A(n8831), .ZN(P1_U3215) );
  INV_X1 U10387 ( .A(n8834), .ZN(n8835) );
  NAND2_X1 U10388 ( .A1(n8833), .A2(n8835), .ZN(n8837) );
  OAI21_X1 U10389 ( .B1(n8833), .B2(n8835), .A(n8837), .ZN(n9251) );
  NOR2_X1 U10390 ( .A1(n9251), .A2(n9252), .ZN(n9250) );
  INV_X1 U10391 ( .A(n8836), .ZN(n8839) );
  INV_X1 U10392 ( .A(n8837), .ZN(n8838) );
  OAI21_X1 U10393 ( .B1(n8841), .B2(n5043), .A(n9287), .ZN(n8846) );
  INV_X1 U10394 ( .A(n9788), .ZN(n8843) );
  AOI22_X1 U10395 ( .A1(n9826), .A2(n9299), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8842) );
  OAI21_X1 U10396 ( .B1(n9292), .B2(n8843), .A(n8842), .ZN(n8844) );
  AOI21_X1 U10397 ( .B1(n9289), .B2(n9781), .A(n8844), .ZN(n8845) );
  OAI211_X1 U10398 ( .C1(n10249), .C2(n9302), .A(n8846), .B(n8845), .ZN(
        P1_U3216) );
  XNOR2_X1 U10399 ( .A(n9260), .B(n8847), .ZN(n8848) );
  NAND2_X1 U10400 ( .A1(n8848), .A2(n8849), .ZN(n9259) );
  OAI21_X1 U10401 ( .B1(n8849), .B2(n8848), .A(n9259), .ZN(n8850) );
  NAND2_X1 U10402 ( .A1(n8850), .A2(n9287), .ZN(n8856) );
  NAND2_X1 U10403 ( .A1(n9299), .A2(n10018), .ZN(n8852) );
  OAI211_X1 U10404 ( .C1(n8853), .C2(n9301), .A(n8852), .B(n8851), .ZN(n8854)
         );
  AOI21_X1 U10405 ( .B1(n4392), .B2(n9305), .A(n8854), .ZN(n8855) );
  OAI211_X1 U10406 ( .C1(n10423), .C2(n9302), .A(n8856), .B(n8855), .ZN(
        P1_U3217) );
  INV_X1 U10407 ( .A(n8866), .ZN(n8865) );
  XNOR2_X1 U10408 ( .A(n8865), .B(n8868), .ZN(n8858) );
  XNOR2_X1 U10409 ( .A(n8857), .B(n8858), .ZN(n8864) );
  NAND2_X1 U10410 ( .A1(n9861), .A2(n9289), .ZN(n8860) );
  OAI211_X1 U10411 ( .C1(n9893), .C2(n9277), .A(n8860), .B(n8859), .ZN(n8862)
         );
  NOR2_X1 U10412 ( .A1(n10262), .A2(n9302), .ZN(n8861) );
  AOI211_X1 U10413 ( .C1(n9863), .C2(n9305), .A(n8862), .B(n8861), .ZN(n8863)
         );
  OAI21_X1 U10414 ( .B1(n8864), .B2(n9307), .A(n8863), .ZN(P1_U3219) );
  INV_X1 U10415 ( .A(n10256), .ZN(n9837) );
  NOR2_X1 U10416 ( .A1(n8857), .A2(n8865), .ZN(n8869) );
  INV_X1 U10417 ( .A(n8857), .ZN(n8867) );
  OAI22_X1 U10418 ( .A1(n8869), .A2(n8868), .B1(n8867), .B2(n8866), .ZN(n9233)
         );
  NAND2_X1 U10419 ( .A1(n8871), .A2(n8870), .ZN(n9234) );
  NOR2_X1 U10420 ( .A1(n9233), .A2(n9234), .ZN(n9232) );
  INV_X1 U10421 ( .A(n8871), .ZN(n8873) );
  NOR3_X1 U10422 ( .A1(n9232), .A2(n8873), .A3(n8872), .ZN(n8874) );
  OAI21_X1 U10423 ( .B1(n8874), .B2(n5046), .A(n9287), .ZN(n8880) );
  NOR2_X1 U10424 ( .A1(n9833), .A2(n9292), .ZN(n8878) );
  OAI22_X1 U10425 ( .A1(n8876), .A2(n9277), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8875), .ZN(n8877) );
  AOI211_X1 U10426 ( .C1(n9289), .C2(n9826), .A(n8878), .B(n8877), .ZN(n8879)
         );
  OAI211_X1 U10427 ( .C1(n9837), .C2(n9302), .A(n8880), .B(n8879), .ZN(
        P1_U3223) );
  OAI21_X1 U10428 ( .B1(n8883), .B2(n8882), .A(n8881), .ZN(n8884) );
  NAND2_X1 U10429 ( .A1(n8884), .A2(n9287), .ZN(n8888) );
  AOI22_X1 U10430 ( .A1(n9289), .A2(n9746), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8885) );
  OAI21_X1 U10431 ( .B1(n9751), .B2(n9292), .A(n8885), .ZN(n8886) );
  AOI21_X1 U10432 ( .B1(n9299), .B2(n9781), .A(n8886), .ZN(n8887) );
  OAI211_X1 U10433 ( .C1(n4891), .C2(n9302), .A(n8888), .B(n8887), .ZN(
        P1_U3225) );
  NAND2_X1 U10434 ( .A1(n4439), .A2(n8889), .ZN(n8890) );
  OAI21_X1 U10435 ( .B1(n4439), .B2(n8889), .A(n8890), .ZN(n9297) );
  NOR2_X1 U10436 ( .A1(n9297), .A2(n9298), .ZN(n9296) );
  INV_X1 U10437 ( .A(n8890), .ZN(n8891) );
  NOR3_X1 U10438 ( .A1(n9296), .A2(n8892), .A3(n8891), .ZN(n8895) );
  INV_X1 U10439 ( .A(n8893), .ZN(n8894) );
  OAI21_X1 U10440 ( .B1(n8895), .B2(n8894), .A(n9287), .ZN(n8900) );
  NOR2_X1 U10441 ( .A1(n8896), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9685) );
  AOI21_X1 U10442 ( .B1(n9289), .B2(n9914), .A(n9685), .ZN(n8897) );
  OAI21_X1 U10443 ( .B1(n9942), .B2(n9277), .A(n8897), .ZN(n8898) );
  AOI21_X1 U10444 ( .B1(n9917), .B2(n9305), .A(n8898), .ZN(n8899) );
  OAI211_X1 U10445 ( .C1(n9909), .C2(n9302), .A(n8900), .B(n8899), .ZN(
        P1_U3226) );
  AOI22_X1 U10446 ( .A1(n8902), .A2(keyinput51), .B1(n9107), .B2(keyinput83), 
        .ZN(n8901) );
  OAI221_X1 U10447 ( .B1(n8902), .B2(keyinput51), .C1(n9107), .C2(keyinput83), 
        .A(n8901), .ZN(n8913) );
  AOI22_X1 U10448 ( .A1(n9109), .A2(keyinput4), .B1(n10187), .B2(keyinput27), 
        .ZN(n8903) );
  OAI221_X1 U10449 ( .B1(n9109), .B2(keyinput4), .C1(n10187), .C2(keyinput27), 
        .A(n8903), .ZN(n8912) );
  AOI22_X1 U10450 ( .A1(n8906), .A2(keyinput84), .B1(n8905), .B2(keyinput120), 
        .ZN(n8904) );
  OAI221_X1 U10451 ( .B1(n8906), .B2(keyinput84), .C1(n8905), .C2(keyinput120), 
        .A(n8904), .ZN(n8911) );
  INV_X1 U10452 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8909) );
  AOI22_X1 U10453 ( .A1(n8909), .A2(keyinput7), .B1(n8908), .B2(keyinput32), 
        .ZN(n8907) );
  OAI221_X1 U10454 ( .B1(n8909), .B2(keyinput7), .C1(n8908), .C2(keyinput32), 
        .A(n8907), .ZN(n8910) );
  NOR4_X1 U10455 ( .A1(n8913), .A2(n8912), .A3(n8911), .A4(n8910), .ZN(n8942)
         );
  AOI22_X1 U10456 ( .A1(n8916), .A2(keyinput26), .B1(n8915), .B2(keyinput98), 
        .ZN(n8914) );
  OAI221_X1 U10457 ( .B1(n8916), .B2(keyinput26), .C1(n8915), .C2(keyinput98), 
        .A(n8914), .ZN(n8920) );
  AOI22_X1 U10458 ( .A1(n8441), .A2(keyinput38), .B1(n8918), .B2(keyinput103), 
        .ZN(n8917) );
  OAI221_X1 U10459 ( .B1(n8441), .B2(keyinput38), .C1(n8918), .C2(keyinput103), 
        .A(n8917), .ZN(n8919) );
  NOR2_X1 U10460 ( .A1(n8920), .A2(n8919), .ZN(n8941) );
  AOI22_X1 U10461 ( .A1(n9051), .A2(keyinput102), .B1(keyinput33), .B2(n8467), 
        .ZN(n8921) );
  OAI221_X1 U10462 ( .B1(n9051), .B2(keyinput102), .C1(n8467), .C2(keyinput33), 
        .A(n8921), .ZN(n8928) );
  AOI22_X1 U10463 ( .A1(n8923), .A2(keyinput125), .B1(n9103), .B2(keyinput36), 
        .ZN(n8922) );
  OAI221_X1 U10464 ( .B1(n8923), .B2(keyinput125), .C1(n9103), .C2(keyinput36), 
        .A(n8922), .ZN(n8927) );
  XNOR2_X1 U10465 ( .A(keyinput46), .B(n8924), .ZN(n8926) );
  XNOR2_X1 U10466 ( .A(keyinput15), .B(n7253), .ZN(n8925) );
  NOR4_X1 U10467 ( .A1(n8928), .A2(n8927), .A3(n8926), .A4(n8925), .ZN(n8940)
         );
  AOI22_X1 U10468 ( .A1(n9072), .A2(keyinput0), .B1(n5094), .B2(keyinput43), 
        .ZN(n8929) );
  OAI221_X1 U10469 ( .B1(n9072), .B2(keyinput0), .C1(n5094), .C2(keyinput43), 
        .A(n8929), .ZN(n8938) );
  AOI22_X1 U10470 ( .A1(n8932), .A2(keyinput106), .B1(n8931), .B2(keyinput57), 
        .ZN(n8930) );
  OAI221_X1 U10471 ( .B1(n8932), .B2(keyinput106), .C1(n8931), .C2(keyinput57), 
        .A(n8930), .ZN(n8937) );
  AOI22_X1 U10472 ( .A1(n8935), .A2(keyinput9), .B1(n8934), .B2(keyinput126), 
        .ZN(n8933) );
  OAI221_X1 U10473 ( .B1(n8935), .B2(keyinput9), .C1(n8934), .C2(keyinput126), 
        .A(n8933), .ZN(n8936) );
  NOR3_X1 U10474 ( .A1(n8938), .A2(n8937), .A3(n8936), .ZN(n8939) );
  NAND4_X1 U10475 ( .A1(n8942), .A2(n8941), .A3(n8940), .A4(n8939), .ZN(n8980)
         );
  AOI22_X1 U10476 ( .A1(n8944), .A2(keyinput41), .B1(keyinput22), .B2(n10169), 
        .ZN(n8943) );
  OAI221_X1 U10477 ( .B1(n8944), .B2(keyinput41), .C1(n10169), .C2(keyinput22), 
        .A(n8943), .ZN(n8953) );
  AOI22_X1 U10478 ( .A1(n9106), .A2(keyinput122), .B1(keyinput39), .B2(n8946), 
        .ZN(n8945) );
  OAI221_X1 U10479 ( .B1(n9106), .B2(keyinput122), .C1(n8946), .C2(keyinput39), 
        .A(n8945), .ZN(n8952) );
  AOI22_X1 U10480 ( .A1(n8948), .A2(keyinput61), .B1(keyinput3), .B2(n9108), 
        .ZN(n8947) );
  OAI221_X1 U10481 ( .B1(n8948), .B2(keyinput61), .C1(n9108), .C2(keyinput3), 
        .A(n8947), .ZN(n8951) );
  AOI22_X1 U10482 ( .A1(n9045), .A2(keyinput81), .B1(n4589), .B2(keyinput114), 
        .ZN(n8949) );
  OAI221_X1 U10483 ( .B1(n9045), .B2(keyinput81), .C1(n4589), .C2(keyinput114), 
        .A(n8949), .ZN(n8950) );
  NOR4_X1 U10484 ( .A1(n8953), .A2(n8952), .A3(n8951), .A4(n8950), .ZN(n8978)
         );
  INV_X1 U10485 ( .A(SI_18_), .ZN(n9064) );
  AOI22_X1 U10486 ( .A1(n9064), .A2(keyinput66), .B1(keyinput108), .B2(n8955), 
        .ZN(n8954) );
  OAI221_X1 U10487 ( .B1(n9064), .B2(keyinput66), .C1(n8955), .C2(keyinput108), 
        .A(n8954), .ZN(n8958) );
  INV_X1 U10488 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U10489 ( .A1(n9074), .A2(keyinput73), .B1(keyinput88), .B2(n10409), 
        .ZN(n8956) );
  OAI221_X1 U10490 ( .B1(n9074), .B2(keyinput73), .C1(n10409), .C2(keyinput88), 
        .A(n8956), .ZN(n8957) );
  NOR2_X1 U10491 ( .A1(n8958), .A2(n8957), .ZN(n8977) );
  INV_X1 U10492 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9092) );
  AOI22_X1 U10493 ( .A1(n9092), .A2(keyinput30), .B1(keyinput110), .B2(n8960), 
        .ZN(n8959) );
  OAI221_X1 U10494 ( .B1(n9092), .B2(keyinput30), .C1(n8960), .C2(keyinput110), 
        .A(n8959), .ZN(n8965) );
  INV_X1 U10495 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8963) );
  AOI22_X1 U10496 ( .A1(n8963), .A2(keyinput79), .B1(keyinput87), .B2(n8962), 
        .ZN(n8961) );
  OAI221_X1 U10497 ( .B1(n8963), .B2(keyinput79), .C1(n8962), .C2(keyinput87), 
        .A(n8961), .ZN(n8964) );
  NOR2_X1 U10498 ( .A1(n8965), .A2(n8964), .ZN(n8976) );
  AOI22_X1 U10499 ( .A1(n8968), .A2(keyinput44), .B1(keyinput35), .B2(n8967), 
        .ZN(n8966) );
  OAI221_X1 U10500 ( .B1(n8968), .B2(keyinput44), .C1(n8967), .C2(keyinput35), 
        .A(n8966), .ZN(n8974) );
  INV_X1 U10501 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9065) );
  AOI22_X1 U10502 ( .A1(n8970), .A2(keyinput58), .B1(keyinput67), .B2(n9065), 
        .ZN(n8969) );
  OAI221_X1 U10503 ( .B1(n8970), .B2(keyinput58), .C1(n9065), .C2(keyinput67), 
        .A(n8969), .ZN(n8973) );
  AOI22_X1 U10504 ( .A1(n9062), .A2(keyinput95), .B1(keyinput76), .B2(n9071), 
        .ZN(n8971) );
  OAI221_X1 U10505 ( .B1(n9062), .B2(keyinput95), .C1(n9071), .C2(keyinput76), 
        .A(n8971), .ZN(n8972) );
  NOR3_X1 U10506 ( .A1(n8974), .A2(n8973), .A3(n8972), .ZN(n8975) );
  NAND4_X1 U10507 ( .A1(n8978), .A2(n8977), .A3(n8976), .A4(n8975), .ZN(n8979)
         );
  NOR2_X1 U10508 ( .A1(n8980), .A2(n8979), .ZN(n9044) );
  XNOR2_X1 U10509 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput92), .ZN(n8984) );
  XNOR2_X1 U10510 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(keyinput97), .ZN(n8983)
         );
  XNOR2_X1 U10511 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput25), .ZN(n8982) );
  XNOR2_X1 U10512 ( .A(P2_REG0_REG_22__SCAN_IN), .B(keyinput23), .ZN(n8981) );
  NAND4_X1 U10513 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), .ZN(n8990)
         );
  XNOR2_X1 U10514 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput19), .ZN(n8988) );
  XNOR2_X1 U10515 ( .A(P2_REG2_REG_31__SCAN_IN), .B(keyinput1), .ZN(n8987) );
  XNOR2_X1 U10516 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput20), .ZN(n8986) );
  XNOR2_X1 U10517 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(keyinput117), .ZN(n8985)
         );
  NAND4_X1 U10518 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(n8989)
         );
  NOR2_X1 U10519 ( .A1(n8990), .A2(n8989), .ZN(n9024) );
  XNOR2_X1 U10520 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput127), .ZN(n8994) );
  XNOR2_X1 U10521 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput123), .ZN(n8993)
         );
  XNOR2_X1 U10522 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput124), .ZN(n8992) );
  XNOR2_X1 U10523 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(keyinput115), .ZN(n8991)
         );
  NAND4_X1 U10524 ( .A1(n8994), .A2(n8993), .A3(n8992), .A4(n8991), .ZN(n9000)
         );
  XNOR2_X1 U10525 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput118), .ZN(n8998) );
  XNOR2_X1 U10526 ( .A(P1_REG1_REG_28__SCAN_IN), .B(keyinput112), .ZN(n8997)
         );
  XNOR2_X1 U10527 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput107), .ZN(n8996) );
  XNOR2_X1 U10528 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput111), .ZN(n8995) );
  NAND4_X1 U10529 ( .A1(n8998), .A2(n8997), .A3(n8996), .A4(n8995), .ZN(n8999)
         );
  NOR2_X1 U10530 ( .A1(n9000), .A2(n8999), .ZN(n9023) );
  XNOR2_X1 U10531 ( .A(P2_REG1_REG_10__SCAN_IN), .B(keyinput104), .ZN(n9004)
         );
  XNOR2_X1 U10532 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput90), .ZN(n9003) );
  XNOR2_X1 U10533 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput96), .ZN(n9002) );
  XNOR2_X1 U10534 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput78), .ZN(n9001) );
  NAND4_X1 U10535 ( .A1(n9004), .A2(n9003), .A3(n9002), .A4(n9001), .ZN(n9010)
         );
  XNOR2_X1 U10536 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput60), .ZN(n9008) );
  XNOR2_X1 U10537 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(keyinput62), .ZN(n9007)
         );
  XNOR2_X1 U10538 ( .A(SI_7_), .B(keyinput52), .ZN(n9006) );
  XNOR2_X1 U10539 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput56), .ZN(n9005) );
  NAND4_X1 U10540 ( .A1(n9008), .A2(n9007), .A3(n9006), .A4(n9005), .ZN(n9009)
         );
  NOR2_X1 U10541 ( .A1(n9010), .A2(n9009), .ZN(n9022) );
  XNOR2_X1 U10542 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput50), .ZN(n9014) );
  XNOR2_X1 U10543 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput34), .ZN(n9013) );
  XNOR2_X1 U10544 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput45), .ZN(n9012) );
  XNOR2_X1 U10545 ( .A(P2_D_REG_0__SCAN_IN), .B(keyinput31), .ZN(n9011) );
  NAND4_X1 U10546 ( .A1(n9014), .A2(n9013), .A3(n9012), .A4(n9011), .ZN(n9020)
         );
  XNOR2_X1 U10547 ( .A(P2_REG0_REG_28__SCAN_IN), .B(keyinput18), .ZN(n9018) );
  XNOR2_X1 U10548 ( .A(n10448), .B(keyinput29), .ZN(n9017) );
  XNOR2_X1 U10549 ( .A(P1_REG0_REG_15__SCAN_IN), .B(keyinput17), .ZN(n9016) );
  XNOR2_X1 U10550 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput8), .ZN(n9015) );
  NAND4_X1 U10551 ( .A1(n9018), .A2(n9017), .A3(n9016), .A4(n9015), .ZN(n9019)
         );
  NOR2_X1 U10552 ( .A1(n9020), .A2(n9019), .ZN(n9021) );
  AND4_X1 U10553 ( .A1(n9024), .A2(n9023), .A3(n9022), .A4(n9021), .ZN(n9043)
         );
  AOI22_X1 U10554 ( .A1(n9026), .A2(keyinput71), .B1(keyinput63), .B2(n9056), 
        .ZN(n9025) );
  OAI221_X1 U10555 ( .B1(n9026), .B2(keyinput71), .C1(n9056), .C2(keyinput63), 
        .A(n9025), .ZN(n9033) );
  INV_X1 U10556 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10379) );
  XNOR2_X1 U10557 ( .A(n10379), .B(keyinput86), .ZN(n9032) );
  XNOR2_X1 U10558 ( .A(keyinput119), .B(P2_REG0_REG_5__SCAN_IN), .ZN(n9030) );
  XNOR2_X1 U10559 ( .A(keyinput100), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9029)
         );
  XNOR2_X1 U10560 ( .A(keyinput89), .B(P1_REG0_REG_5__SCAN_IN), .ZN(n9028) );
  XNOR2_X1 U10561 ( .A(keyinput94), .B(P1_D_REG_23__SCAN_IN), .ZN(n9027) );
  NAND4_X1 U10562 ( .A1(n9030), .A2(n9029), .A3(n9028), .A4(n9027), .ZN(n9031)
         );
  NOR3_X1 U10563 ( .A1(n9033), .A2(n9032), .A3(n9031), .ZN(n9042) );
  AOI22_X1 U10564 ( .A1(n9035), .A2(keyinput13), .B1(n6258), .B2(keyinput65), 
        .ZN(n9034) );
  OAI221_X1 U10565 ( .B1(n9035), .B2(keyinput13), .C1(n6258), .C2(keyinput65), 
        .A(n9034), .ZN(n9040) );
  AOI22_X1 U10566 ( .A1(n10315), .A2(keyinput2), .B1(n9037), .B2(keyinput11), 
        .ZN(n9036) );
  OAI221_X1 U10567 ( .B1(n10315), .B2(keyinput2), .C1(n9037), .C2(keyinput11), 
        .A(n9036), .ZN(n9039) );
  INV_X1 U10568 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10301) );
  XNOR2_X1 U10569 ( .A(n10301), .B(keyinput113), .ZN(n9038) );
  NOR3_X1 U10570 ( .A1(n9040), .A2(n9039), .A3(n9038), .ZN(n9041) );
  AND4_X1 U10571 ( .A1(n9044), .A2(n9043), .A3(n9042), .A4(n9041), .ZN(n9186)
         );
  NAND4_X1 U10572 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), 
        .A3(P2_REG3_REG_13__SCAN_IN), .A4(P2_REG2_REG_28__SCAN_IN), .ZN(n9050)
         );
  NAND4_X1 U10573 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P2_DATAO_REG_24__SCAN_IN), .A3(P1_ADDR_REG_15__SCAN_IN), .A4(n9045), .ZN(n9049) );
  INV_X1 U10574 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9046) );
  NAND4_X1 U10575 ( .A1(n9046), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_IR_REG_17__SCAN_IN), .ZN(n9048) );
  NAND4_X1 U10576 ( .A1(n8960), .A2(P2_REG1_REG_1__SCAN_IN), .A3(
        P2_D_REG_0__SCAN_IN), .A4(P1_DATAO_REG_10__SCAN_IN), .ZN(n9047) );
  OR4_X1 U10577 ( .A1(n9050), .A2(n9049), .A3(n9048), .A4(n9047), .ZN(n9102)
         );
  INV_X1 U10578 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10376) );
  NAND4_X1 U10579 ( .A1(n10376), .A2(n9126), .A3(n9124), .A4(
        P2_REG3_REG_3__SCAN_IN), .ZN(n9101) );
  NAND4_X1 U10580 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), 
        .A3(P2_REG2_REG_24__SCAN_IN), .A4(n9051), .ZN(n9100) );
  INV_X1 U10581 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10260) );
  NAND4_X1 U10582 ( .A1(n9168), .A2(n10260), .A3(n9145), .A4(
        P1_REG1_REG_28__SCAN_IN), .ZN(n9060) );
  NAND4_X1 U10583 ( .A1(n9053), .A2(n9052), .A3(n5238), .A4(
        P2_IR_REG_2__SCAN_IN), .ZN(n9059) );
  NAND4_X1 U10584 ( .A1(n9055), .A2(n9054), .A3(n4710), .A4(
        P2_IR_REG_20__SCAN_IN), .ZN(n9058) );
  NAND4_X1 U10585 ( .A1(n9056), .A2(P2_REG3_REG_21__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .A4(P2_REG1_REG_10__SCAN_IN), .ZN(n9057) );
  NOR4_X1 U10586 ( .A1(n9060), .A2(n9059), .A3(n9058), .A4(n9057), .ZN(n9098)
         );
  NAND4_X1 U10587 ( .A1(n9063), .A2(n9062), .A3(n9061), .A4(
        P1_D_REG_1__SCAN_IN), .ZN(n9090) );
  NAND4_X1 U10588 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .A3(P1_REG3_REG_27__SCAN_IN), .A4(n9064), .ZN(n9070) );
  INV_X1 U10589 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10395) );
  OR4_X1 U10590 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_27__SCAN_IN), 
        .A3(n10395), .A4(n9065), .ZN(n9069) );
  NAND4_X1 U10591 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .A3(n9170), .A4(n9066), .ZN(n9068) );
  NOR4_X1 U10592 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .ZN(n9086)
         );
  NAND4_X1 U10593 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(SI_31_), .A3(
        P2_ADDR_REG_13__SCAN_IN), .A4(n9071), .ZN(n9078) );
  NAND4_X1 U10594 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(P2_ADDR_REG_18__SCAN_IN), 
        .A3(n9073), .A4(n9072), .ZN(n9077) );
  NAND4_X1 U10595 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .A3(P1_REG3_REG_13__SCAN_IN), .A4(n5094), .ZN(n9076) );
  NAND4_X1 U10596 ( .A1(P1_REG0_REG_7__SCAN_IN), .A2(P2_REG0_REG_21__SCAN_IN), 
        .A3(n9074), .A4(n6073), .ZN(n9075) );
  NOR4_X1 U10597 ( .A1(n9078), .A2(n9077), .A3(n9076), .A4(n9075), .ZN(n9085)
         );
  NAND4_X1 U10598 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(P1_REG2_REG_14__SCAN_IN), 
        .A3(P2_ADDR_REG_16__SCAN_IN), .A4(n9140), .ZN(n9083) );
  NAND4_X1 U10599 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(P2_DATAO_REG_15__SCAN_IN), .A3(P2_IR_REG_25__SCAN_IN), .A4(n7253), .ZN(n9082) );
  NAND4_X1 U10600 ( .A1(P1_REG1_REG_1__SCAN_IN), .A2(n10159), .A3(n9079), .A4(
        n9132), .ZN(n9081) );
  NAND4_X1 U10601 ( .A1(SI_15_), .A2(P1_REG0_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_7__SCAN_IN), .A4(P2_REG0_REG_5__SCAN_IN), .ZN(n9080) );
  NOR4_X1 U10602 ( .A1(n9083), .A2(n9082), .A3(n9081), .A4(n9080), .ZN(n9084)
         );
  NAND4_X1 U10603 ( .A1(n9087), .A2(n9086), .A3(n9085), .A4(n9084), .ZN(n9089)
         );
  NOR4_X1 U10604 ( .A1(n9090), .A2(n9089), .A3(P1_IR_REG_26__SCAN_IN), .A4(
        n9088), .ZN(n9097) );
  INV_X1 U10605 ( .A(SI_7_), .ZN(n9091) );
  NOR4_X1 U10606 ( .A1(n9092), .A2(n9091), .A3(P2_DATAO_REG_7__SCAN_IN), .A4(
        P1_REG3_REG_18__SCAN_IN), .ZN(n9096) );
  INV_X1 U10607 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9093) );
  NOR4_X1 U10608 ( .A1(n9094), .A2(n9093), .A3(P1_REG0_REG_15__SCAN_IN), .A4(
        P1_REG3_REG_6__SCAN_IN), .ZN(n9095) );
  NAND4_X1 U10609 ( .A1(n9098), .A2(n9097), .A3(n9096), .A4(n9095), .ZN(n9099)
         );
  OR4_X1 U10610 ( .A1(n9102), .A2(n9101), .A3(n9100), .A4(n9099), .ZN(n9116)
         );
  NOR4_X1 U10611 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P2_REG0_REG_10__SCAN_IN), 
        .A3(P2_ADDR_REG_6__SCAN_IN), .A4(n9103), .ZN(n9104) );
  NAND4_X1 U10612 ( .A1(n9105), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_REG2_REG_26__SCAN_IN), .A4(n9104), .ZN(n9115) );
  NOR4_X1 U10613 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(P2_REG0_REG_7__SCAN_IN), 
        .A3(n9107), .A4(n9106), .ZN(n9113) );
  NOR4_X1 U10614 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_REG1_REG_17__SCAN_IN), 
        .A3(P2_IR_REG_3__SCAN_IN), .A4(P2_REG0_REG_22__SCAN_IN), .ZN(n9112) );
  INV_X1 U10615 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10233) );
  NOR4_X1 U10616 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(P1_DATAO_REG_3__SCAN_IN), 
        .A3(n10233), .A4(n9108), .ZN(n9111) );
  NOR4_X1 U10617 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .A3(n10187), .A4(n9109), .ZN(n9110) );
  NAND4_X1 U10618 ( .A1(n9113), .A2(n9112), .A3(n9111), .A4(n9110), .ZN(n9114)
         );
  NOR3_X1 U10619 ( .A1(n9116), .A2(n9115), .A3(n9114), .ZN(n9118) );
  INV_X1 U10620 ( .A(keyinput37), .ZN(n9117) );
  OAI21_X1 U10621 ( .B1(n9118), .B2(P2_IR_REG_27__SCAN_IN), .A(n9117), .ZN(
        n9185) );
  AOI22_X1 U10622 ( .A1(n9120), .A2(keyinput55), .B1(keyinput72), .B2(n7355), 
        .ZN(n9119) );
  OAI221_X1 U10623 ( .B1(n9120), .B2(keyinput55), .C1(n7355), .C2(keyinput72), 
        .A(n9119), .ZN(n9130) );
  AOI22_X1 U10624 ( .A1(n10376), .A2(keyinput82), .B1(keyinput105), .B2(n9122), 
        .ZN(n9121) );
  OAI221_X1 U10625 ( .B1(n10376), .B2(keyinput82), .C1(n9122), .C2(keyinput105), .A(n9121), .ZN(n9129) );
  INV_X1 U10626 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U10627 ( .A1(n10429), .A2(keyinput21), .B1(keyinput91), .B2(n9124), 
        .ZN(n9123) );
  OAI221_X1 U10628 ( .B1(n10429), .B2(keyinput21), .C1(n9124), .C2(keyinput91), 
        .A(n9123), .ZN(n9128) );
  AOI22_X1 U10629 ( .A1(n9126), .A2(keyinput59), .B1(keyinput80), .B2(n6073), 
        .ZN(n9125) );
  OAI221_X1 U10630 ( .B1(n9126), .B2(keyinput59), .C1(n6073), .C2(keyinput80), 
        .A(n9125), .ZN(n9127) );
  NOR4_X1 U10631 ( .A1(n9130), .A2(n9129), .A3(n9128), .A4(n9127), .ZN(n9184)
         );
  INV_X1 U10632 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U10633 ( .A1(n10378), .A2(keyinput6), .B1(keyinput10), .B2(n9132), 
        .ZN(n9131) );
  OAI221_X1 U10634 ( .B1(n10378), .B2(keyinput6), .C1(n9132), .C2(keyinput10), 
        .A(n9131), .ZN(n9136) );
  INV_X1 U10635 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9134) );
  AOI22_X1 U10636 ( .A1(n9046), .A2(keyinput74), .B1(n9134), .B2(keyinput70), 
        .ZN(n9133) );
  OAI221_X1 U10637 ( .B1(n9046), .B2(keyinput74), .C1(n9134), .C2(keyinput70), 
        .A(n9133), .ZN(n9135) );
  NOR2_X1 U10638 ( .A1(n9136), .A2(n9135), .ZN(n9166) );
  AOI22_X1 U10639 ( .A1(n7603), .A2(keyinput116), .B1(n9138), .B2(keyinput93), 
        .ZN(n9137) );
  OAI221_X1 U10640 ( .B1(n7603), .B2(keyinput116), .C1(n9138), .C2(keyinput93), 
        .A(n9137), .ZN(n9143) );
  AOI22_X1 U10641 ( .A1(n9141), .A2(keyinput48), .B1(keyinput75), .B2(n9140), 
        .ZN(n9139) );
  OAI221_X1 U10642 ( .B1(n9141), .B2(keyinput48), .C1(n9140), .C2(keyinput75), 
        .A(n9139), .ZN(n9142) );
  NOR2_X1 U10643 ( .A1(n9143), .A2(n9142), .ZN(n9165) );
  AOI22_X1 U10644 ( .A1(n9146), .A2(keyinput54), .B1(n9145), .B2(keyinput24), 
        .ZN(n9144) );
  OAI221_X1 U10645 ( .B1(n9146), .B2(keyinput54), .C1(n9145), .C2(keyinput24), 
        .A(n9144), .ZN(n9152) );
  XNOR2_X1 U10646 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput5), .ZN(n9150) );
  XNOR2_X1 U10647 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput53), .ZN(n9149) );
  XNOR2_X1 U10648 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput109), .ZN(n9148) );
  NAND2_X1 U10649 ( .A1(n5180), .A2(keyinput37), .ZN(n9147) );
  NAND4_X1 U10650 ( .A1(n9150), .A2(n9149), .A3(n9148), .A4(n9147), .ZN(n9151)
         );
  NOR2_X1 U10651 ( .A1(n9152), .A2(n9151), .ZN(n9164) );
  XNOR2_X1 U10652 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput28), .ZN(n9156) );
  XNOR2_X1 U10653 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput14), .ZN(n9155) );
  XNOR2_X1 U10654 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput121), .ZN(n9154) );
  XNOR2_X1 U10655 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput101), .ZN(n9153) );
  NAND4_X1 U10656 ( .A1(n9156), .A2(n9155), .A3(n9154), .A4(n9153), .ZN(n9162)
         );
  XNOR2_X1 U10657 ( .A(P1_REG0_REG_30__SCAN_IN), .B(keyinput49), .ZN(n9160) );
  XNOR2_X1 U10658 ( .A(P1_REG1_REG_17__SCAN_IN), .B(keyinput85), .ZN(n9159) );
  XNOR2_X1 U10659 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput99), .ZN(n9158) );
  XNOR2_X1 U10660 ( .A(P1_REG1_REG_24__SCAN_IN), .B(keyinput16), .ZN(n9157) );
  NAND4_X1 U10661 ( .A1(n9160), .A2(n9159), .A3(n9158), .A4(n9157), .ZN(n9161)
         );
  NOR2_X1 U10662 ( .A1(n9162), .A2(n9161), .ZN(n9163) );
  NAND4_X1 U10663 ( .A1(n9166), .A2(n9165), .A3(n9164), .A4(n9163), .ZN(n9182)
         );
  AOI22_X1 U10664 ( .A1(n10260), .A2(keyinput47), .B1(keyinput68), .B2(n9168), 
        .ZN(n9167) );
  OAI221_X1 U10665 ( .B1(n10260), .B2(keyinput47), .C1(n9168), .C2(keyinput68), 
        .A(n9167), .ZN(n9176) );
  AOI22_X1 U10666 ( .A1(n9171), .A2(keyinput64), .B1(keyinput69), .B2(n9170), 
        .ZN(n9169) );
  OAI221_X1 U10667 ( .B1(n9171), .B2(keyinput64), .C1(n9170), .C2(keyinput69), 
        .A(n9169), .ZN(n9175) );
  INV_X1 U10668 ( .A(SI_15_), .ZN(n9173) );
  AOI22_X1 U10669 ( .A1(n9173), .A2(keyinput42), .B1(keyinput77), .B2(n4710), 
        .ZN(n9172) );
  OAI221_X1 U10670 ( .B1(n9173), .B2(keyinput42), .C1(n4710), .C2(keyinput77), 
        .A(n9172), .ZN(n9174) );
  OR3_X1 U10671 ( .A1(n9176), .A2(n9175), .A3(n9174), .ZN(n9181) );
  XNOR2_X1 U10672 ( .A(n9177), .B(keyinput40), .ZN(n9180) );
  XNOR2_X1 U10673 ( .A(n9178), .B(keyinput12), .ZN(n9179) );
  NOR4_X1 U10674 ( .A1(n9182), .A2(n9181), .A3(n9180), .A4(n9179), .ZN(n9183)
         );
  NAND4_X1 U10675 ( .A1(n9186), .A2(n9185), .A3(n9184), .A4(n9183), .ZN(n9196)
         );
  OAI21_X1 U10676 ( .B1(n9189), .B2(n9188), .A(n9187), .ZN(n9194) );
  NAND2_X1 U10677 ( .A1(n10197), .A2(n9256), .ZN(n9192) );
  NAND2_X1 U10678 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9701) );
  OAI21_X1 U10679 ( .B1(n9277), .B2(n9894), .A(n9701), .ZN(n9190) );
  AOI21_X1 U10680 ( .B1(n9289), .B2(n9860), .A(n9190), .ZN(n9191) );
  OAI211_X1 U10681 ( .C1(n9292), .C2(n9897), .A(n9192), .B(n9191), .ZN(n9193)
         );
  AOI21_X1 U10682 ( .B1(n9194), .B2(n9287), .A(n9193), .ZN(n9195) );
  XOR2_X1 U10683 ( .A(n9196), .B(n9195), .Z(P1_U3228) );
  INV_X1 U10684 ( .A(n9767), .ZN(n10245) );
  INV_X1 U10685 ( .A(n9197), .ZN(n9199) );
  NOR3_X1 U10686 ( .A1(n5043), .A2(n9199), .A3(n9198), .ZN(n9203) );
  INV_X1 U10687 ( .A(n9201), .ZN(n9202) );
  OAI21_X1 U10688 ( .B1(n9203), .B2(n9202), .A(n9287), .ZN(n9208) );
  OAI22_X1 U10689 ( .A1(n9768), .A2(n9292), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9204), .ZN(n9206) );
  NOR2_X1 U10690 ( .A1(n9309), .A2(n9277), .ZN(n9205) );
  AOI211_X1 U10691 ( .C1(n9289), .C2(n9762), .A(n9206), .B(n9205), .ZN(n9207)
         );
  OAI211_X1 U10692 ( .C1(n10245), .C2(n9302), .A(n9208), .B(n9207), .ZN(
        P1_U3229) );
  OAI21_X1 U10693 ( .B1(n9211), .B2(n9210), .A(n9209), .ZN(n9212) );
  NAND3_X1 U10694 ( .A1(n9213), .A2(n9287), .A3(n9212), .ZN(n9219) );
  NAND2_X1 U10695 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9600) );
  OAI21_X1 U10696 ( .B1(n9277), .B2(n9214), .A(n9600), .ZN(n9215) );
  AOI21_X1 U10697 ( .B1(n9289), .B2(n9569), .A(n9215), .ZN(n9218) );
  AOI22_X1 U10698 ( .A1(n9305), .A2(n10087), .B1(n9216), .B2(n9256), .ZN(n9217) );
  NAND3_X1 U10699 ( .A1(n9219), .A2(n9218), .A3(n9217), .ZN(P1_U3230) );
  AOI21_X1 U10700 ( .B1(n9221), .B2(n7962), .A(n9220), .ZN(n9225) );
  XOR2_X1 U10701 ( .A(n9223), .B(n9222), .Z(n9224) );
  XNOR2_X1 U10702 ( .A(n9225), .B(n9224), .ZN(n9231) );
  AOI21_X1 U10703 ( .B1(n9299), .B2(n9566), .A(n9226), .ZN(n9228) );
  NAND2_X1 U10704 ( .A1(n9305), .A2(n10046), .ZN(n9227) );
  OAI211_X1 U10705 ( .C1(n10043), .C2(n9301), .A(n9228), .B(n9227), .ZN(n9229)
         );
  AOI21_X1 U10706 ( .B1(n10050), .B2(n9256), .A(n9229), .ZN(n9230) );
  OAI21_X1 U10707 ( .B1(n9231), .B2(n9307), .A(n9230), .ZN(P1_U3231) );
  AOI21_X1 U10708 ( .B1(n9234), .B2(n9233), .A(n9232), .ZN(n9240) );
  AOI22_X1 U10709 ( .A1(n9299), .A2(n9845), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9236) );
  NAND2_X1 U10710 ( .A1(n9305), .A2(n9850), .ZN(n9235) );
  OAI211_X1 U10711 ( .C1(n9237), .C2(n9301), .A(n9236), .B(n9235), .ZN(n9238)
         );
  AOI21_X1 U10712 ( .B1(n10180), .B2(n9256), .A(n9238), .ZN(n9239) );
  OAI21_X1 U10713 ( .B1(n9240), .B2(n9307), .A(n9239), .ZN(P1_U3233) );
  OAI21_X1 U10714 ( .B1(n9243), .B2(n9242), .A(n9241), .ZN(n9244) );
  NAND2_X1 U10715 ( .A1(n9244), .A2(n9287), .ZN(n9249) );
  AOI21_X1 U10716 ( .B1(n9289), .B2(n9929), .A(n9245), .ZN(n9246) );
  OAI21_X1 U10717 ( .B1(n9968), .B2(n9277), .A(n9246), .ZN(n9247) );
  AOI21_X1 U10718 ( .B1(n9971), .B2(n9305), .A(n9247), .ZN(n9248) );
  OAI211_X1 U10719 ( .C1(n4882), .C2(n9302), .A(n9249), .B(n9248), .ZN(
        P1_U3234) );
  AOI21_X1 U10720 ( .B1(n9252), .B2(n9251), .A(n9250), .ZN(n9258) );
  NAND2_X1 U10721 ( .A1(n9803), .A2(n9289), .ZN(n9254) );
  AOI22_X1 U10722 ( .A1(n9846), .A2(n9299), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9253) );
  OAI211_X1 U10723 ( .C1(n9292), .C2(n9809), .A(n9254), .B(n9253), .ZN(n9255)
         );
  AOI21_X1 U10724 ( .B1(n9808), .B2(n9256), .A(n9255), .ZN(n9257) );
  OAI21_X1 U10725 ( .B1(n9258), .B2(n9307), .A(n9257), .ZN(P1_U3235) );
  OAI21_X1 U10726 ( .B1(n9261), .B2(n9260), .A(n9259), .ZN(n9265) );
  XNOR2_X1 U10727 ( .A(n9263), .B(n9262), .ZN(n9264) );
  XNOR2_X1 U10728 ( .A(n9265), .B(n9264), .ZN(n9270) );
  NAND2_X1 U10729 ( .A1(n9299), .A2(n9994), .ZN(n9266) );
  NAND2_X1 U10730 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9675) );
  OAI211_X1 U10731 ( .C1(n9968), .C2(n9301), .A(n9266), .B(n9675), .ZN(n9268)
         );
  NOR2_X1 U10732 ( .A1(n10006), .A2(n9302), .ZN(n9267) );
  AOI211_X1 U10733 ( .C1(n10003), .C2(n9305), .A(n9268), .B(n9267), .ZN(n9269)
         );
  OAI21_X1 U10734 ( .B1(n9270), .B2(n9307), .A(n9269), .ZN(P1_U3236) );
  INV_X1 U10735 ( .A(n9271), .ZN(n9275) );
  OAI21_X1 U10736 ( .B1(n9275), .B2(n9273), .A(n9272), .ZN(n9274) );
  OAI211_X1 U10737 ( .C1(n9276), .C2(n9275), .A(n9287), .B(n9274), .ZN(n9281)
         );
  NAND2_X1 U10738 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10329)
         );
  OAI21_X1 U10739 ( .B1(n9277), .B2(n9877), .A(n10329), .ZN(n9279) );
  NOR2_X1 U10740 ( .A1(n9292), .A2(n9882), .ZN(n9278) );
  AOI211_X1 U10741 ( .C1(n9289), .C2(n9845), .A(n9279), .B(n9278), .ZN(n9280)
         );
  OAI211_X1 U10742 ( .C1(n10267), .C2(n9302), .A(n9281), .B(n9280), .ZN(
        P1_U3238) );
  NAND2_X1 U10743 ( .A1(n9285), .A2(n9284), .ZN(n9288) );
  NAND3_X1 U10744 ( .A1(n9288), .A2(n9287), .A3(n9286), .ZN(n9295) );
  INV_X1 U10745 ( .A(n9736), .ZN(n9291) );
  AOI22_X1 U10746 ( .A1(n9289), .A2(n9732), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9290) );
  OAI21_X1 U10747 ( .B1(n9292), .B2(n9291), .A(n9290), .ZN(n9293) );
  AOI21_X1 U10748 ( .B1(n9762), .B2(n9299), .A(n9293), .ZN(n9294) );
  OAI211_X1 U10749 ( .C1(n10240), .C2(n9302), .A(n9295), .B(n9294), .ZN(
        P1_U3240) );
  AOI21_X1 U10750 ( .B1(n9298), .B2(n9297), .A(n9296), .ZN(n9308) );
  NAND2_X1 U10751 ( .A1(n9299), .A2(n9929), .ZN(n9300) );
  NAND2_X1 U10752 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10313)
         );
  OAI211_X1 U10753 ( .C1(n9894), .C2(n9301), .A(n9300), .B(n10313), .ZN(n9304)
         );
  NOR2_X1 U10754 ( .A1(n9935), .A2(n9302), .ZN(n9303) );
  AOI211_X1 U10755 ( .C1(n9932), .C2(n9305), .A(n9304), .B(n9303), .ZN(n9306)
         );
  OAI21_X1 U10756 ( .B1(n9308), .B2(n9307), .A(n9306), .ZN(P1_U3241) );
  OR2_X1 U10757 ( .A1(n9787), .A2(n9309), .ZN(n9391) );
  NAND2_X1 U10758 ( .A1(n9391), .A2(n9310), .ZN(n9452) );
  NAND2_X1 U10759 ( .A1(n9871), .A2(n9514), .ZN(n9311) );
  MUX2_X1 U10760 ( .A(n9312), .B(n9311), .S(n9315), .Z(n9373) );
  AND2_X1 U10761 ( .A1(n9485), .A2(n4380), .ZN(n9313) );
  AOI21_X1 U10762 ( .B1(n10106), .B2(n9313), .A(n10366), .ZN(n9326) );
  INV_X1 U10763 ( .A(n9314), .ZN(n9319) );
  OR2_X1 U10764 ( .A1(n9322), .A2(n9315), .ZN(n9318) );
  INV_X1 U10765 ( .A(n9485), .ZN(n9316) );
  NAND2_X1 U10766 ( .A1(n9316), .A2(n9546), .ZN(n9317) );
  OAI211_X1 U10767 ( .C1(n9320), .C2(n9319), .A(n9318), .B(n9317), .ZN(n9321)
         );
  INV_X1 U10768 ( .A(n9321), .ZN(n9325) );
  OR3_X1 U10769 ( .A1(n10106), .A2(n9323), .A3(n4380), .ZN(n9324) );
  NAND4_X1 U10770 ( .A1(n9326), .A2(n10070), .A3(n9325), .A4(n9324), .ZN(n9340) );
  NAND2_X1 U10771 ( .A1(n10073), .A2(n9546), .ZN(n9335) );
  OAI21_X1 U10772 ( .B1(n9335), .B2(n9568), .A(n10360), .ZN(n9330) );
  OR2_X1 U10773 ( .A1(n10073), .A2(n9315), .ZN(n9327) );
  OAI21_X1 U10774 ( .B1(n9327), .B2(n10350), .A(n10392), .ZN(n9329) );
  OAI22_X1 U10775 ( .A1(n9327), .A2(n10360), .B1(n10350), .B2(n9315), .ZN(
        n9328) );
  AOI22_X1 U10776 ( .A1(n9330), .A2(n9329), .B1(n9328), .B2(n10397), .ZN(n9339) );
  NAND4_X1 U10777 ( .A1(n5017), .A2(n10031), .A3(n6472), .A4(n9315), .ZN(n9333) );
  INV_X1 U10778 ( .A(n9484), .ZN(n9331) );
  NAND4_X1 U10779 ( .A1(n9492), .A2(n9490), .A3(n9331), .A4(n4380), .ZN(n9332)
         );
  AND2_X1 U10780 ( .A1(n9333), .A2(n9332), .ZN(n9338) );
  NAND2_X1 U10781 ( .A1(n10350), .A2(n9546), .ZN(n9334) );
  OAI21_X1 U10782 ( .B1(n9335), .B2(n10392), .A(n9334), .ZN(n9336) );
  NAND2_X1 U10783 ( .A1(n9336), .A2(n10079), .ZN(n9337) );
  NAND4_X1 U10784 ( .A1(n9340), .A2(n9339), .A3(n9338), .A4(n9337), .ZN(n9342)
         );
  INV_X1 U10785 ( .A(n10336), .ZN(n9341) );
  NAND2_X1 U10786 ( .A1(n9496), .A2(n9344), .ZN(n9345) );
  NAND3_X1 U10787 ( .A1(n9348), .A2(n9500), .A3(n9359), .ZN(n9350) );
  NAND3_X1 U10788 ( .A1(n9350), .A2(n9506), .A3(n9349), .ZN(n9353) );
  MUX2_X1 U10789 ( .A(n9507), .B(n9944), .S(n9315), .Z(n9351) );
  INV_X1 U10790 ( .A(n9351), .ZN(n9352) );
  NOR2_X1 U10791 ( .A1(n9947), .A2(n9352), .ZN(n9363) );
  NAND3_X1 U10792 ( .A1(n9353), .A2(n9363), .A3(n9360), .ZN(n9355) );
  AND2_X1 U10793 ( .A1(n9370), .A2(n9354), .ZN(n9512) );
  AOI21_X1 U10794 ( .B1(n9355), .B2(n9512), .A(n9546), .ZN(n9368) );
  INV_X1 U10795 ( .A(n9496), .ZN(n9356) );
  OAI21_X1 U10796 ( .B1(n9357), .B2(n9356), .A(n9500), .ZN(n9358) );
  NAND2_X1 U10797 ( .A1(n9358), .A2(n9504), .ZN(n9361) );
  AND2_X1 U10798 ( .A1(n9360), .A2(n9359), .ZN(n9502) );
  NAND2_X1 U10799 ( .A1(n9361), .A2(n9502), .ZN(n9362) );
  NAND3_X1 U10800 ( .A1(n9362), .A2(n9506), .A3(n9315), .ZN(n9366) );
  INV_X1 U10801 ( .A(n9965), .ZN(n9365) );
  INV_X1 U10802 ( .A(n9363), .ZN(n9364) );
  AOI21_X1 U10803 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9367) );
  NAND2_X1 U10804 ( .A1(n9513), .A2(n9508), .ZN(n9369) );
  OAI21_X1 U10805 ( .B1(n4380), .B2(n9370), .A(n9910), .ZN(n9371) );
  INV_X1 U10806 ( .A(n9429), .ZN(n9372) );
  NAND2_X1 U10807 ( .A1(n9378), .A2(n9519), .ZN(n9374) );
  NOR2_X1 U10808 ( .A1(n9452), .A2(n9375), .ZN(n9385) );
  NAND2_X1 U10809 ( .A1(n9376), .A2(n9546), .ZN(n9387) );
  INV_X1 U10810 ( .A(n9387), .ZN(n9384) );
  AND2_X1 U10811 ( .A1(n9451), .A2(n9377), .ZN(n9458) );
  NAND3_X1 U10812 ( .A1(n9379), .A2(n9821), .A3(n9520), .ZN(n9382) );
  AOI21_X1 U10813 ( .B1(n9820), .B2(n9380), .A(n9546), .ZN(n9381) );
  AOI21_X1 U10814 ( .B1(n9382), .B2(n9546), .A(n9381), .ZN(n9383) );
  OAI211_X1 U10815 ( .C1(n9385), .C2(n9384), .A(n9458), .B(n9383), .ZN(n9398)
         );
  NOR2_X1 U10816 ( .A1(n9452), .A2(n9546), .ZN(n9390) );
  INV_X1 U10817 ( .A(n9386), .ZN(n9389) );
  OAI22_X1 U10818 ( .A1(n9801), .A2(n4380), .B1(n9523), .B2(n9387), .ZN(n9388)
         );
  AOI22_X1 U10819 ( .A1(n9390), .A2(n9389), .B1(n9388), .B2(n9458), .ZN(n9397)
         );
  INV_X1 U10820 ( .A(n9391), .ZN(n9393) );
  INV_X1 U10821 ( .A(n9451), .ZN(n9392) );
  MUX2_X1 U10822 ( .A(n9393), .B(n9392), .S(n4380), .Z(n9394) );
  INV_X1 U10823 ( .A(n9394), .ZN(n9395) );
  INV_X1 U10824 ( .A(n9757), .ZN(n9759) );
  MUX2_X1 U10825 ( .A(n9454), .B(n9459), .S(n9315), .Z(n9399) );
  AND2_X1 U10826 ( .A1(n9524), .A2(n9460), .ZN(n9408) );
  INV_X1 U10827 ( .A(n9408), .ZN(n9401) );
  AOI21_X1 U10828 ( .B1(n9410), .B2(n9457), .A(n9401), .ZN(n9404) );
  OR2_X1 U10829 ( .A1(n9735), .A2(n9402), .ZN(n9406) );
  INV_X1 U10830 ( .A(n9406), .ZN(n9403) );
  OAI21_X1 U10831 ( .B1(n9404), .B2(n9403), .A(n9411), .ZN(n9405) );
  AND2_X1 U10832 ( .A1(n9407), .A2(n9406), .ZN(n9468) );
  INV_X1 U10833 ( .A(n9457), .ZN(n9409) );
  NAND2_X1 U10834 ( .A1(n9412), .A2(n9411), .ZN(n9466) );
  INV_X1 U10835 ( .A(n9449), .ZN(n9414) );
  NOR2_X1 U10836 ( .A1(n9415), .A2(n9414), .ZN(n9416) );
  INV_X1 U10837 ( .A(n9469), .ZN(n9418) );
  INV_X1 U10838 ( .A(n9562), .ZN(n9423) );
  AOI21_X1 U10839 ( .B1(n10236), .B2(n9469), .A(n9546), .ZN(n9422) );
  AND2_X1 U10840 ( .A1(n9707), .A2(n9562), .ZN(n9473) );
  NOR2_X1 U10841 ( .A1(n9423), .A2(n9447), .ZN(n9471) );
  OAI22_X1 U10842 ( .A1(n9544), .A2(n9425), .B1(n6518), .B2(n9551), .ZN(n9478)
         );
  OR2_X1 U10843 ( .A1(n9715), .A2(n9447), .ZN(n9426) );
  AND2_X1 U10844 ( .A1(n4483), .A2(n9426), .ZN(n9479) );
  NAND2_X1 U10845 ( .A1(n9428), .A2(n9427), .ZN(n9874) );
  NAND2_X1 U10846 ( .A1(n9871), .A2(n9429), .ZN(n9890) );
  AND4_X1 U10847 ( .A1(n10095), .A2(n10134), .A3(n9431), .A4(n9430), .ZN(n9434) );
  NOR2_X1 U10848 ( .A1(n10366), .A2(n10030), .ZN(n9433) );
  NAND4_X1 U10849 ( .A1(n9434), .A2(n9433), .A3(n9496), .A4(n9432), .ZN(n9436)
         );
  NOR4_X1 U10850 ( .A1(n9436), .A2(n9435), .A3(n10034), .A4(n9497), .ZN(n9440)
         );
  OR2_X1 U10851 ( .A1(n9438), .A2(n9437), .ZN(n9993) );
  NOR4_X1 U10852 ( .A1(n9874), .A2(n9890), .A3(n6496), .A4(n9441), .ZN(n9442)
         );
  NAND4_X1 U10853 ( .A1(n9801), .A2(n9843), .A3(n9857), .A4(n9442), .ZN(n9443)
         );
  NOR4_X1 U10854 ( .A1(n9446), .A2(n9728), .A3(n9445), .A4(n4486), .ZN(n9448)
         );
  NAND2_X1 U10855 ( .A1(n9715), .A2(n9447), .ZN(n9470) );
  INV_X1 U10856 ( .A(n9473), .ZN(n9552) );
  NAND2_X1 U10857 ( .A1(n9450), .A2(n9449), .ZN(n9533) );
  NAND2_X1 U10858 ( .A1(n9452), .A2(n9451), .ZN(n9453) );
  NAND2_X1 U10859 ( .A1(n9454), .A2(n9453), .ZN(n9455) );
  NAND2_X1 U10860 ( .A1(n9455), .A2(n9459), .ZN(n9456) );
  AND2_X1 U10861 ( .A1(n9457), .A2(n9456), .ZN(n9463) );
  INV_X1 U10862 ( .A(n9463), .ZN(n9526) );
  OAI21_X1 U10863 ( .B1(n9526), .B2(n9799), .A(n9524), .ZN(n9467) );
  INV_X1 U10864 ( .A(n9468), .ZN(n9529) );
  NAND3_X1 U10865 ( .A1(n9459), .A2(n9458), .A3(n9798), .ZN(n9462) );
  INV_X1 U10866 ( .A(n9460), .ZN(n9461) );
  AOI21_X1 U10867 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(n9464) );
  NOR2_X1 U10868 ( .A1(n9529), .A2(n9464), .ZN(n9465) );
  OR2_X1 U10869 ( .A1(n9466), .A2(n9465), .ZN(n9531) );
  NAND2_X1 U10870 ( .A1(n9470), .A2(n9469), .ZN(n9535) );
  OAI211_X1 U10871 ( .C1(n9474), .C2(n9473), .A(n9472), .B(n4483), .ZN(n9475)
         );
  INV_X1 U10872 ( .A(n9479), .ZN(n9537) );
  OR2_X1 U10873 ( .A1(n9480), .A2(n4391), .ZN(n9483) );
  AND4_X1 U10874 ( .A1(n9483), .A2(n6518), .A3(n9482), .A4(n9481), .ZN(n9487)
         );
  AND3_X1 U10875 ( .A1(n9485), .A2(n6472), .A3(n9484), .ZN(n9486) );
  OAI21_X1 U10876 ( .B1(n9488), .B2(n9487), .A(n9486), .ZN(n9495) );
  NAND2_X1 U10877 ( .A1(n9490), .A2(n9489), .ZN(n9491) );
  NAND2_X1 U10878 ( .A1(n9491), .A2(n6472), .ZN(n9493) );
  AND2_X1 U10879 ( .A1(n9493), .A2(n9492), .ZN(n9494) );
  NAND4_X1 U10880 ( .A1(n9495), .A2(n9494), .A3(n9496), .A4(n9498), .ZN(n9501)
         );
  NAND3_X1 U10881 ( .A1(n9498), .A2(n9497), .A3(n9496), .ZN(n9499) );
  NAND3_X1 U10882 ( .A1(n9501), .A2(n9500), .A3(n9499), .ZN(n9505) );
  INV_X1 U10883 ( .A(n9502), .ZN(n9503) );
  AOI21_X1 U10884 ( .B1(n9505), .B2(n9504), .A(n9503), .ZN(n9510) );
  NAND2_X1 U10885 ( .A1(n9944), .A2(n9506), .ZN(n9509) );
  OAI211_X1 U10886 ( .C1(n9510), .C2(n9509), .A(n9508), .B(n9507), .ZN(n9511)
         );
  NAND2_X1 U10887 ( .A1(n9512), .A2(n9511), .ZN(n9515) );
  NAND3_X1 U10888 ( .A1(n9515), .A2(n9514), .A3(n9513), .ZN(n9517) );
  NAND2_X1 U10889 ( .A1(n9517), .A2(n9516), .ZN(n9518) );
  AOI21_X1 U10890 ( .B1(n9519), .B2(n9518), .A(n4447), .ZN(n9521) );
  OAI21_X1 U10891 ( .B1(n9521), .B2(n4461), .A(n9520), .ZN(n9522) );
  NAND2_X1 U10892 ( .A1(n9523), .A2(n9522), .ZN(n9525) );
  OAI21_X1 U10893 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9527) );
  INV_X1 U10894 ( .A(n9527), .ZN(n9528) );
  NOR2_X1 U10895 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  NOR2_X1 U10896 ( .A1(n9531), .A2(n9530), .ZN(n9532) );
  NOR2_X1 U10897 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  NOR2_X1 U10898 ( .A1(n9535), .A2(n9534), .ZN(n9536) );
  OR2_X1 U10899 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  NAND2_X1 U10900 ( .A1(n9538), .A2(n9552), .ZN(n9543) );
  NAND3_X1 U10901 ( .A1(n9543), .A2(n9540), .A3(n9539), .ZN(n9542) );
  INV_X1 U10902 ( .A(n9556), .ZN(n9541) );
  INV_X1 U10903 ( .A(n9544), .ZN(n9545) );
  OAI21_X1 U10904 ( .B1(n9546), .B2(n4483), .A(n9545), .ZN(n9550) );
  NOR4_X1 U10905 ( .A1(n9548), .A2(n9557), .A3(P1_U3086), .A4(n9547), .ZN(
        n9549) );
  OAI211_X1 U10906 ( .C1(n9552), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9559)
         );
  NAND2_X1 U10907 ( .A1(n9554), .A2(n9553), .ZN(n9555) );
  OAI211_X1 U10908 ( .C1(n9557), .C2(n9556), .A(n9555), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9558) );
  OAI211_X1 U10909 ( .C1(n9561), .C2(n9560), .A(n9559), .B(n9558), .ZN(
        P1_U3242) );
  MUX2_X1 U10910 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9562), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10911 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9563), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10912 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9564), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10913 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9732), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10914 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9746), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10915 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9762), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10916 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9781), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10917 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9803), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10918 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9826), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10919 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9846), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10920 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9861), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10921 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9845), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10922 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9860), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10923 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9914), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10924 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9928), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10925 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9913), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10926 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9929), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10927 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9565), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10928 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9995), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10929 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n10016), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10930 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9994), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10931 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n10018), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10932 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9566), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10933 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9567), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10934 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9568), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10935 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9569), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10936 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n10364), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10937 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9570), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10938 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9571), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10939 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9572), .S(P1_U3973), .Z(
        P1_U3555) );
  INV_X1 U10940 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9574) );
  OAI22_X1 U10941 ( .A1(n10332), .A2(n9574), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9573), .ZN(n9575) );
  AOI21_X1 U10942 ( .B1(n9576), .B2(n10312), .A(n9575), .ZN(n9585) );
  OAI211_X1 U10943 ( .C1(n9579), .C2(n9578), .A(n10286), .B(n9577), .ZN(n9584)
         );
  OAI211_X1 U10944 ( .C1(n9582), .C2(n9581), .A(n10319), .B(n9580), .ZN(n9583)
         );
  NAND3_X1 U10945 ( .A1(n9585), .A2(n9584), .A3(n9583), .ZN(P1_U3244) );
  INV_X1 U10946 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9587) );
  OAI21_X1 U10947 ( .B1(n10332), .B2(n9587), .A(n9586), .ZN(n9588) );
  AOI21_X1 U10948 ( .B1(n9589), .B2(n10312), .A(n9588), .ZN(n9598) );
  OAI211_X1 U10949 ( .C1(n9592), .C2(n9591), .A(n10319), .B(n9590), .ZN(n9597)
         );
  OAI211_X1 U10950 ( .C1(n9595), .C2(n9594), .A(n10286), .B(n9593), .ZN(n9596)
         );
  NAND3_X1 U10951 ( .A1(n9598), .A2(n9597), .A3(n9596), .ZN(P1_U3246) );
  INV_X1 U10952 ( .A(n9599), .ZN(n9603) );
  INV_X1 U10953 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9601) );
  OAI21_X1 U10954 ( .B1(n10332), .B2(n9601), .A(n9600), .ZN(n9602) );
  AOI21_X1 U10955 ( .B1(n9603), .B2(n10312), .A(n9602), .ZN(n9612) );
  OAI211_X1 U10956 ( .C1(n9606), .C2(n9605), .A(n10286), .B(n9604), .ZN(n9611)
         );
  OAI211_X1 U10957 ( .C1(n9609), .C2(n9608), .A(n10319), .B(n9607), .ZN(n9610)
         );
  NAND4_X1 U10958 ( .A1(n9613), .A2(n9612), .A3(n9611), .A4(n9610), .ZN(
        P1_U3247) );
  INV_X1 U10959 ( .A(n9614), .ZN(n9618) );
  INV_X1 U10960 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9616) );
  OAI21_X1 U10961 ( .B1(n10332), .B2(n9616), .A(n9615), .ZN(n9617) );
  AOI21_X1 U10962 ( .B1(n9618), .B2(n10312), .A(n9617), .ZN(n9627) );
  OAI211_X1 U10963 ( .C1(n9621), .C2(n9620), .A(n10319), .B(n9619), .ZN(n9626)
         );
  OAI211_X1 U10964 ( .C1(n9624), .C2(n9623), .A(n10286), .B(n9622), .ZN(n9625)
         );
  NAND3_X1 U10965 ( .A1(n9627), .A2(n9626), .A3(n9625), .ZN(P1_U3248) );
  INV_X1 U10966 ( .A(n9628), .ZN(n9632) );
  INV_X1 U10967 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9630) );
  OAI21_X1 U10968 ( .B1(n10332), .B2(n9630), .A(n9629), .ZN(n9631) );
  AOI21_X1 U10969 ( .B1(n9632), .B2(n10312), .A(n9631), .ZN(n9641) );
  OAI211_X1 U10970 ( .C1(n9635), .C2(n9634), .A(n10286), .B(n9633), .ZN(n9640)
         );
  OAI211_X1 U10971 ( .C1(n9638), .C2(n9637), .A(n10319), .B(n9636), .ZN(n9639)
         );
  NAND3_X1 U10972 ( .A1(n9641), .A2(n9640), .A3(n9639), .ZN(P1_U3249) );
  INV_X1 U10973 ( .A(n9642), .ZN(n9646) );
  INV_X1 U10974 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9644) );
  OAI21_X1 U10975 ( .B1(n10332), .B2(n9644), .A(n9643), .ZN(n9645) );
  AOI21_X1 U10976 ( .B1(n9646), .B2(n10312), .A(n9645), .ZN(n9655) );
  OAI211_X1 U10977 ( .C1(n9649), .C2(n9648), .A(n10286), .B(n9647), .ZN(n9654)
         );
  OAI211_X1 U10978 ( .C1(n9652), .C2(n9651), .A(n10319), .B(n9650), .ZN(n9653)
         );
  NAND3_X1 U10979 ( .A1(n9655), .A2(n9654), .A3(n9653), .ZN(P1_U3250) );
  INV_X1 U10980 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9657) );
  OAI21_X1 U10981 ( .B1(n10332), .B2(n9657), .A(n9656), .ZN(n9658) );
  AOI21_X1 U10982 ( .B1(n9659), .B2(n10312), .A(n9658), .ZN(n9668) );
  OAI211_X1 U10983 ( .C1(n9662), .C2(n9661), .A(n10319), .B(n9660), .ZN(n9667)
         );
  OAI211_X1 U10984 ( .C1(n9665), .C2(n9664), .A(n10286), .B(n9663), .ZN(n9666)
         );
  NAND3_X1 U10985 ( .A1(n9668), .A2(n9667), .A3(n9666), .ZN(P1_U3251) );
  OAI211_X1 U10986 ( .C1(n9671), .C2(n9670), .A(n9669), .B(n10319), .ZN(n9681)
         );
  OAI211_X1 U10987 ( .C1(n9674), .C2(n9673), .A(n9672), .B(n10286), .ZN(n9680)
         );
  INV_X1 U10988 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9676) );
  OAI21_X1 U10989 ( .B1(n10332), .B2(n9676), .A(n9675), .ZN(n9677) );
  AOI21_X1 U10990 ( .B1(n9678), .B2(n10312), .A(n9677), .ZN(n9679) );
  NAND3_X1 U10991 ( .A1(n9681), .A2(n9680), .A3(n9679), .ZN(P1_U3254) );
  OAI21_X1 U10992 ( .B1(n9684), .B2(n9683), .A(n9682), .ZN(n9693) );
  INV_X1 U10993 ( .A(n10312), .ZN(n10325) );
  AOI21_X1 U10994 ( .B1(n9699), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9685), .ZN(
        n9686) );
  OAI21_X1 U10995 ( .B1(n10325), .B2(n9687), .A(n9686), .ZN(n9692) );
  AOI211_X1 U10996 ( .C1(n9690), .C2(n9689), .A(n9688), .B(n10316), .ZN(n9691)
         );
  AOI211_X1 U10997 ( .C1(n10319), .C2(n9693), .A(n9692), .B(n9691), .ZN(n9694)
         );
  INV_X1 U10998 ( .A(n9694), .ZN(P1_U3259) );
  XOR2_X1 U10999 ( .A(n9696), .B(n9695), .Z(n9706) );
  XNOR2_X1 U11000 ( .A(n9698), .B(n9697), .ZN(n9704) );
  NAND2_X1 U11001 ( .A1(n9699), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9700) );
  OAI211_X1 U11002 ( .C1(n10325), .C2(n9702), .A(n9701), .B(n9700), .ZN(n9703)
         );
  AOI21_X1 U11003 ( .B1(n9704), .B2(n10319), .A(n9703), .ZN(n9705) );
  OAI21_X1 U11004 ( .B1(n9706), .B2(n10316), .A(n9705), .ZN(P1_U3260) );
  NOR2_X1 U11005 ( .A1(n4377), .A2(n10142), .ZN(n9714) );
  NOR2_X1 U11006 ( .A1(n9707), .A2(n10123), .ZN(n9708) );
  AOI211_X1 U11007 ( .C1(n4377), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9714), .B(
        n9708), .ZN(n9709) );
  OAI21_X1 U11008 ( .B1(n9710), .B2(n10101), .A(n9709), .ZN(P1_U3263) );
  OAI211_X1 U11009 ( .C1(n10236), .C2(n9712), .A(n10369), .B(n9711), .ZN(
        n10143) );
  AND2_X1 U11010 ( .A1(n4377), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9713) );
  NOR2_X1 U11011 ( .A1(n9714), .A2(n9713), .ZN(n9717) );
  NAND2_X1 U11012 ( .A1(n9715), .A2(n10359), .ZN(n9716) );
  OAI211_X1 U11013 ( .C1(n10143), .C2(n10101), .A(n9717), .B(n9716), .ZN(
        P1_U3264) );
  INV_X1 U11014 ( .A(n9718), .ZN(n9724) );
  AOI22_X1 U11015 ( .A1(n4377), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9719), .B2(
        n10358), .ZN(n9720) );
  OAI21_X1 U11016 ( .B1(n9721), .B2(n10123), .A(n9720), .ZN(n9723) );
  XNOR2_X1 U11017 ( .A(n9726), .B(n9728), .ZN(n10148) );
  INV_X1 U11018 ( .A(n10148), .ZN(n9741) );
  NAND2_X1 U11019 ( .A1(n9729), .A2(n9728), .ZN(n9730) );
  NAND2_X1 U11020 ( .A1(n9727), .A2(n9730), .ZN(n9731) );
  NAND2_X1 U11021 ( .A1(n9731), .A2(n10014), .ZN(n9734) );
  AOI22_X1 U11022 ( .A1(n9762), .A2(n10356), .B1(n10017), .B2(n9732), .ZN(
        n9733) );
  AOI211_X1 U11023 ( .C1(n9735), .C2(n9749), .A(n10214), .B(n6521), .ZN(n10147) );
  NAND2_X1 U11024 ( .A1(n10147), .A2(n10372), .ZN(n9738) );
  AOI22_X1 U11025 ( .A1(n4377), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9736), .B2(
        n10358), .ZN(n9737) );
  OAI211_X1 U11026 ( .C1(n10240), .C2(n10123), .A(n9738), .B(n9737), .ZN(n9739) );
  AOI21_X1 U11027 ( .B1(n10112), .B2(n10146), .A(n9739), .ZN(n9740) );
  OAI21_X1 U11028 ( .B1(n9741), .B2(n10124), .A(n9740), .ZN(P1_U3267) );
  XOR2_X1 U11029 ( .A(n9742), .B(n9744), .Z(n10155) );
  OAI211_X1 U11030 ( .C1(n9745), .C2(n9744), .A(n9743), .B(n10014), .ZN(n9748)
         );
  AOI22_X1 U11031 ( .A1(n9781), .A2(n10356), .B1(n10017), .B2(n9746), .ZN(
        n9747) );
  NAND2_X1 U11032 ( .A1(n9748), .A2(n9747), .ZN(n10152) );
  INV_X1 U11033 ( .A(n9749), .ZN(n9750) );
  AOI211_X1 U11034 ( .C1(n10153), .C2(n9765), .A(n10214), .B(n9750), .ZN(
        n10151) );
  NAND2_X1 U11035 ( .A1(n10151), .A2(n10372), .ZN(n9754) );
  INV_X1 U11036 ( .A(n9751), .ZN(n9752) );
  AOI22_X1 U11037 ( .A1(n9752), .A2(n10358), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n4377), .ZN(n9753) );
  OAI211_X1 U11038 ( .C1(n4891), .C2(n10123), .A(n9754), .B(n9753), .ZN(n9755)
         );
  AOI21_X1 U11039 ( .B1(n10112), .B2(n10152), .A(n9755), .ZN(n9756) );
  OAI21_X1 U11040 ( .B1(n10155), .B2(n10124), .A(n9756), .ZN(P1_U3268) );
  XNOR2_X1 U11041 ( .A(n9758), .B(n9757), .ZN(n10158) );
  INV_X1 U11042 ( .A(n10158), .ZN(n9774) );
  XNOR2_X1 U11043 ( .A(n9760), .B(n9759), .ZN(n9761) );
  NAND2_X1 U11044 ( .A1(n9761), .A2(n10014), .ZN(n9764) );
  AOI22_X1 U11045 ( .A1(n9762), .A2(n10017), .B1(n10356), .B2(n9803), .ZN(
        n9763) );
  NAND2_X1 U11046 ( .A1(n9764), .A2(n9763), .ZN(n10157) );
  INV_X1 U11047 ( .A(n9765), .ZN(n9766) );
  AOI211_X1 U11048 ( .C1(n9767), .C2(n9784), .A(n10214), .B(n9766), .ZN(n10156) );
  NAND2_X1 U11049 ( .A1(n10156), .A2(n10372), .ZN(n9771) );
  INV_X1 U11050 ( .A(n9768), .ZN(n9769) );
  AOI22_X1 U11051 ( .A1(n9769), .A2(n10358), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n4377), .ZN(n9770) );
  OAI211_X1 U11052 ( .C1(n10245), .C2(n10123), .A(n9771), .B(n9770), .ZN(n9772) );
  AOI21_X1 U11053 ( .B1(n10112), .B2(n10157), .A(n9772), .ZN(n9773) );
  OAI21_X1 U11054 ( .B1(n9774), .B2(n10124), .A(n9773), .ZN(P1_U3269) );
  XOR2_X1 U11055 ( .A(n9775), .B(n9776), .Z(n10163) );
  INV_X1 U11056 ( .A(n10163), .ZN(n9793) );
  NAND2_X1 U11057 ( .A1(n9777), .A2(n9776), .ZN(n9778) );
  NAND2_X1 U11058 ( .A1(n9779), .A2(n9778), .ZN(n9780) );
  NAND2_X1 U11059 ( .A1(n9780), .A2(n10014), .ZN(n9783) );
  AOI22_X1 U11060 ( .A1(n9781), .A2(n10017), .B1(n10356), .B2(n9826), .ZN(
        n9782) );
  NAND2_X1 U11061 ( .A1(n9783), .A2(n9782), .ZN(n10162) );
  INV_X1 U11062 ( .A(n9806), .ZN(n9786) );
  INV_X1 U11063 ( .A(n9784), .ZN(n9785) );
  AOI211_X1 U11064 ( .C1(n9787), .C2(n9786), .A(n10214), .B(n9785), .ZN(n10161) );
  NAND2_X1 U11065 ( .A1(n10161), .A2(n10372), .ZN(n9790) );
  AOI22_X1 U11066 ( .A1(n9788), .A2(n10358), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n4377), .ZN(n9789) );
  OAI211_X1 U11067 ( .C1(n10249), .C2(n10123), .A(n9790), .B(n9789), .ZN(n9791) );
  AOI21_X1 U11068 ( .B1(n10112), .B2(n10162), .A(n9791), .ZN(n9792) );
  OAI21_X1 U11069 ( .B1(n9793), .B2(n10124), .A(n9792), .ZN(P1_U3270) );
  NAND2_X1 U11070 ( .A1(n9794), .A2(n9795), .ZN(n9818) );
  NAND2_X1 U11071 ( .A1(n9818), .A2(n9817), .ZN(n9816) );
  NAND2_X1 U11072 ( .A1(n9816), .A2(n9796), .ZN(n9797) );
  XNOR2_X1 U11073 ( .A(n9797), .B(n9801), .ZN(n10168) );
  INV_X1 U11074 ( .A(n10168), .ZN(n9815) );
  AND2_X1 U11075 ( .A1(n9799), .A2(n9798), .ZN(n9802) );
  OAI211_X1 U11076 ( .C1(n9802), .C2(n9801), .A(n9800), .B(n10014), .ZN(n9805)
         );
  AOI22_X1 U11077 ( .A1(n9803), .A2(n10017), .B1(n10356), .B2(n9846), .ZN(
        n9804) );
  NAND2_X1 U11078 ( .A1(n9805), .A2(n9804), .ZN(n10166) );
  INV_X1 U11079 ( .A(n9832), .ZN(n9807) );
  AOI211_X1 U11080 ( .C1(n9808), .C2(n9807), .A(n10214), .B(n9806), .ZN(n10167) );
  NAND2_X1 U11081 ( .A1(n10167), .A2(n10372), .ZN(n9812) );
  INV_X1 U11082 ( .A(n9809), .ZN(n9810) );
  AOI22_X1 U11083 ( .A1(n9810), .A2(n10358), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n4377), .ZN(n9811) );
  OAI211_X1 U11084 ( .C1(n10253), .C2(n10123), .A(n9812), .B(n9811), .ZN(n9813) );
  AOI21_X1 U11085 ( .B1(n10112), .B2(n10166), .A(n9813), .ZN(n9814) );
  OAI21_X1 U11086 ( .B1(n10124), .B2(n9815), .A(n9814), .ZN(P1_U3271) );
  OAI21_X1 U11087 ( .B1(n9818), .B2(n9817), .A(n9816), .ZN(n10171) );
  NAND2_X1 U11088 ( .A1(n9819), .A2(n9820), .ZN(n9822) );
  NAND2_X1 U11089 ( .A1(n9822), .A2(n9821), .ZN(n9824) );
  XNOR2_X1 U11090 ( .A(n9824), .B(n9823), .ZN(n9825) );
  NAND2_X1 U11091 ( .A1(n9825), .A2(n10014), .ZN(n9828) );
  AOI22_X1 U11092 ( .A1(n9826), .A2(n10017), .B1(n10356), .B2(n9861), .ZN(
        n9827) );
  NAND2_X1 U11093 ( .A1(n9828), .A2(n9827), .ZN(n10173) );
  INV_X1 U11094 ( .A(n9829), .ZN(n9849) );
  NAND2_X1 U11095 ( .A1(n9849), .A2(n10256), .ZN(n9830) );
  NAND2_X1 U11096 ( .A1(n9830), .A2(n10369), .ZN(n9831) );
  NOR2_X1 U11097 ( .A1(n9832), .A2(n9831), .ZN(n10172) );
  NAND2_X1 U11098 ( .A1(n10172), .A2(n10372), .ZN(n9836) );
  INV_X1 U11099 ( .A(n9833), .ZN(n9834) );
  AOI22_X1 U11100 ( .A1(n9834), .A2(n10358), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n4377), .ZN(n9835) );
  OAI211_X1 U11101 ( .C1(n9837), .C2(n10123), .A(n9836), .B(n9835), .ZN(n9838)
         );
  AOI21_X1 U11102 ( .B1(n10173), .B2(n10112), .A(n9838), .ZN(n9839) );
  OAI21_X1 U11103 ( .B1(n10171), .B2(n10124), .A(n9839), .ZN(P1_U3272) );
  AND2_X1 U11104 ( .A1(n9841), .A2(n9840), .ZN(n9842) );
  OAI21_X1 U11105 ( .B1(n9842), .B2(n6503), .A(n9794), .ZN(n10182) );
  XNOR2_X1 U11106 ( .A(n9819), .B(n9843), .ZN(n9844) );
  NAND2_X1 U11107 ( .A1(n9844), .A2(n10014), .ZN(n9848) );
  AOI22_X1 U11108 ( .A1(n9846), .A2(n10017), .B1(n10356), .B2(n9845), .ZN(
        n9847) );
  NAND2_X1 U11109 ( .A1(n9848), .A2(n9847), .ZN(n10179) );
  AOI211_X1 U11110 ( .C1(n10180), .C2(n9862), .A(n10214), .B(n9829), .ZN(
        n10178) );
  NAND2_X1 U11111 ( .A1(n10178), .A2(n10372), .ZN(n9852) );
  AOI22_X1 U11112 ( .A1(n9850), .A2(n10358), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n4377), .ZN(n9851) );
  OAI211_X1 U11113 ( .C1(n9853), .C2(n10123), .A(n9852), .B(n9851), .ZN(n9854)
         );
  AOI21_X1 U11114 ( .B1(n10112), .B2(n10179), .A(n9854), .ZN(n9855) );
  OAI21_X1 U11115 ( .B1(n10124), .B2(n10182), .A(n9855), .ZN(P1_U3273) );
  XOR2_X1 U11116 ( .A(n9856), .B(n9857), .Z(n10185) );
  XNOR2_X1 U11117 ( .A(n9858), .B(n9857), .ZN(n9859) );
  AOI222_X1 U11118 ( .A1(n9861), .A2(n10017), .B1(n9860), .B2(n10356), .C1(
        n10014), .C2(n9859), .ZN(n10184) );
  INV_X1 U11119 ( .A(n10184), .ZN(n9868) );
  OAI211_X1 U11120 ( .C1(n9879), .C2(n10262), .A(n10369), .B(n9862), .ZN(
        n10183) );
  AOI22_X1 U11121 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(n4377), .B1(n9863), .B2(
        n10358), .ZN(n9866) );
  NAND2_X1 U11122 ( .A1(n9864), .A2(n10359), .ZN(n9865) );
  OAI211_X1 U11123 ( .C1(n10183), .C2(n10101), .A(n9866), .B(n9865), .ZN(n9867) );
  AOI21_X1 U11124 ( .B1(n9868), .B2(n10112), .A(n9867), .ZN(n9869) );
  OAI21_X1 U11125 ( .B1(n10124), .B2(n10185), .A(n9869), .ZN(P1_U3274) );
  XOR2_X1 U11126 ( .A(n9870), .B(n9874), .Z(n10191) );
  INV_X1 U11127 ( .A(n10191), .ZN(n9888) );
  NAND2_X1 U11128 ( .A1(n9872), .A2(n9871), .ZN(n9873) );
  XOR2_X1 U11129 ( .A(n9874), .B(n9873), .Z(n9875) );
  OAI222_X1 U11130 ( .A1(n6460), .A2(n9877), .B1(n6461), .B2(n9876), .C1(n6464), .C2(n9875), .ZN(n10189) );
  INV_X1 U11131 ( .A(n9878), .ZN(n9880) );
  AOI211_X1 U11132 ( .C1(n9881), .C2(n9880), .A(n10214), .B(n9879), .ZN(n10190) );
  NAND2_X1 U11133 ( .A1(n10190), .A2(n10372), .ZN(n9885) );
  INV_X1 U11134 ( .A(n9882), .ZN(n9883) );
  AOI22_X1 U11135 ( .A1(n4377), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9883), .B2(
        n10358), .ZN(n9884) );
  OAI211_X1 U11136 ( .C1(n10267), .C2(n10123), .A(n9885), .B(n9884), .ZN(n9886) );
  AOI21_X1 U11137 ( .B1(n10189), .B2(n10112), .A(n9886), .ZN(n9887) );
  OAI21_X1 U11138 ( .B1(n10124), .B2(n9888), .A(n9887), .ZN(P1_U3275) );
  XNOR2_X1 U11139 ( .A(n9889), .B(n9890), .ZN(n10199) );
  XOR2_X1 U11140 ( .A(n9891), .B(n9890), .Z(n9892) );
  OAI222_X1 U11141 ( .A1(n6460), .A2(n9894), .B1(n6461), .B2(n9893), .C1(n6464), .C2(n9892), .ZN(n10195) );
  NAND2_X1 U11142 ( .A1(n10195), .A2(n10112), .ZN(n9902) );
  OR2_X1 U11143 ( .A1(n9895), .A2(n10271), .ZN(n9906) );
  AOI211_X1 U11144 ( .C1(n10197), .C2(n9906), .A(n10214), .B(n9878), .ZN(
        n10196) );
  INV_X1 U11145 ( .A(n10197), .ZN(n9896) );
  NOR2_X1 U11146 ( .A1(n9896), .A2(n10123), .ZN(n9900) );
  OAI22_X1 U11147 ( .A1(n10112), .A2(n9898), .B1(n9897), .B2(n10097), .ZN(
        n9899) );
  AOI211_X1 U11148 ( .C1(n10196), .C2(n10372), .A(n9900), .B(n9899), .ZN(n9901) );
  OAI211_X1 U11149 ( .C1(n10199), .C2(n10124), .A(n9902), .B(n9901), .ZN(
        P1_U3276) );
  NAND2_X1 U11150 ( .A1(n9903), .A2(n9910), .ZN(n9904) );
  NAND2_X1 U11151 ( .A1(n9905), .A2(n9904), .ZN(n10200) );
  AOI21_X1 U11152 ( .B1(n9895), .B2(n10271), .A(n10214), .ZN(n9907) );
  AND2_X1 U11153 ( .A1(n9907), .A2(n9906), .ZN(n10201) );
  INV_X1 U11154 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9908) );
  OAI22_X1 U11155 ( .A1(n9909), .A2(n10123), .B1(n10112), .B2(n9908), .ZN(
        n9920) );
  XNOR2_X1 U11156 ( .A(n9911), .B(n9910), .ZN(n9912) );
  NAND2_X1 U11157 ( .A1(n9912), .A2(n10014), .ZN(n9916) );
  AOI22_X1 U11158 ( .A1(n9914), .A2(n10017), .B1(n9913), .B2(n10356), .ZN(
        n9915) );
  NAND2_X1 U11159 ( .A1(n9916), .A2(n9915), .ZN(n10202) );
  AOI21_X1 U11160 ( .B1(n9917), .B2(n10358), .A(n10202), .ZN(n9918) );
  NOR2_X1 U11161 ( .A1(n9918), .A2(n4377), .ZN(n9919) );
  AOI211_X1 U11162 ( .C1(n10201), .C2(n10372), .A(n9920), .B(n9919), .ZN(n9921) );
  OAI21_X1 U11163 ( .B1(n10124), .B2(n10200), .A(n9921), .ZN(P1_U3277) );
  XOR2_X1 U11164 ( .A(n9922), .B(n9924), .Z(n10211) );
  INV_X1 U11165 ( .A(n9923), .ZN(n9945) );
  OAI21_X1 U11166 ( .B1(n9945), .B2(n9925), .A(n9924), .ZN(n9927) );
  NAND2_X1 U11167 ( .A1(n9927), .A2(n9926), .ZN(n9930) );
  AOI222_X1 U11168 ( .A1(n10014), .A2(n9930), .B1(n9929), .B2(n10356), .C1(
        n9928), .C2(n10017), .ZN(n10210) );
  INV_X1 U11169 ( .A(n10210), .ZN(n9937) );
  INV_X1 U11170 ( .A(n9895), .ZN(n9931) );
  AOI211_X1 U11171 ( .C1(n10208), .C2(n6016), .A(n10214), .B(n9931), .ZN(
        n10207) );
  NAND2_X1 U11172 ( .A1(n10207), .A2(n10372), .ZN(n9934) );
  AOI22_X1 U11173 ( .A1(n4377), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9932), .B2(
        n10358), .ZN(n9933) );
  OAI211_X1 U11174 ( .C1(n9935), .C2(n10123), .A(n9934), .B(n9933), .ZN(n9936)
         );
  AOI21_X1 U11175 ( .B1(n9937), .B2(n10112), .A(n9936), .ZN(n9938) );
  OAI21_X1 U11176 ( .B1(n10211), .B2(n10124), .A(n9938), .ZN(P1_U3278) );
  INV_X1 U11177 ( .A(n9939), .ZN(n10341) );
  XNOR2_X1 U11178 ( .A(n9940), .B(n9947), .ZN(n10212) );
  OAI22_X1 U11179 ( .A1(n9942), .A2(n6461), .B1(n9941), .B2(n6460), .ZN(n9949)
         );
  NAND2_X1 U11180 ( .A1(n9943), .A2(n9944), .ZN(n9946) );
  AOI211_X1 U11181 ( .C1(n9947), .C2(n9946), .A(n6464), .B(n9945), .ZN(n9948)
         );
  AOI211_X1 U11182 ( .C1(n10341), .C2(n10212), .A(n9949), .B(n9948), .ZN(
        n10218) );
  NOR2_X1 U11183 ( .A1(n4377), .A2(n9950), .ZN(n10346) );
  INV_X1 U11184 ( .A(n9951), .ZN(n9970) );
  AND2_X1 U11185 ( .A1(n9970), .A2(n9955), .ZN(n9953) );
  OR2_X1 U11186 ( .A1(n9953), .A2(n9952), .ZN(n10215) );
  NAND2_X1 U11187 ( .A1(n10372), .A2(n10369), .ZN(n10002) );
  AOI22_X1 U11188 ( .A1(n4377), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9954), .B2(
        n10358), .ZN(n9957) );
  NAND2_X1 U11189 ( .A1(n9955), .A2(n10359), .ZN(n9956) );
  OAI211_X1 U11190 ( .C1(n10215), .C2(n10002), .A(n9957), .B(n9956), .ZN(n9958) );
  AOI21_X1 U11191 ( .B1(n10212), .B2(n10346), .A(n9958), .ZN(n9959) );
  OAI21_X1 U11192 ( .B1(n10218), .B2(n4377), .A(n9959), .ZN(P1_U3279) );
  OAI21_X1 U11193 ( .B1(n9961), .B2(n9965), .A(n9960), .ZN(n9962) );
  INV_X1 U11194 ( .A(n9962), .ZN(n10224) );
  INV_X1 U11195 ( .A(n9943), .ZN(n9963) );
  AOI21_X1 U11196 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(n9966) );
  OAI222_X1 U11197 ( .A1(n6460), .A2(n9968), .B1(n6461), .B2(n9967), .C1(n6464), .C2(n9966), .ZN(n10220) );
  AOI21_X1 U11198 ( .B1(n4491), .B2(n10222), .A(n10214), .ZN(n9969) );
  AND2_X1 U11199 ( .A1(n9970), .A2(n9969), .ZN(n10221) );
  NAND2_X1 U11200 ( .A1(n10221), .A2(n10372), .ZN(n9973) );
  AOI22_X1 U11201 ( .A1(n4377), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9971), .B2(
        n10358), .ZN(n9972) );
  OAI211_X1 U11202 ( .C1(n4882), .C2(n10123), .A(n9973), .B(n9972), .ZN(n9974)
         );
  AOI21_X1 U11203 ( .B1(n10220), .B2(n10112), .A(n9974), .ZN(n9975) );
  OAI21_X1 U11204 ( .B1(n10224), .B2(n10124), .A(n9975), .ZN(P1_U3280) );
  INV_X1 U11205 ( .A(n9976), .ZN(n9985) );
  NAND2_X1 U11206 ( .A1(n9977), .A2(n10372), .ZN(n9980) );
  AOI22_X1 U11207 ( .A1(n4377), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9978), .B2(
        n10358), .ZN(n9979) );
  OAI211_X1 U11208 ( .C1(n9981), .C2(n10123), .A(n9980), .B(n9979), .ZN(n9982)
         );
  AOI21_X1 U11209 ( .B1(n9983), .B2(n10112), .A(n9982), .ZN(n9984) );
  OAI21_X1 U11210 ( .B1(n10124), .B2(n9985), .A(n9984), .ZN(P1_U3281) );
  NAND2_X1 U11211 ( .A1(n9987), .A2(n9986), .ZN(n10010) );
  NAND2_X1 U11212 ( .A1(n10010), .A2(n10009), .ZN(n9989) );
  NAND2_X1 U11213 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  XOR2_X1 U11214 ( .A(n9990), .B(n9993), .Z(n10226) );
  NAND2_X1 U11215 ( .A1(n10011), .A2(n9991), .ZN(n9992) );
  XOR2_X1 U11216 ( .A(n9993), .B(n9992), .Z(n9997) );
  AOI22_X1 U11217 ( .A1(n10017), .A2(n9995), .B1(n9994), .B2(n10356), .ZN(
        n9996) );
  OAI21_X1 U11218 ( .B1(n9997), .B2(n6464), .A(n9996), .ZN(n9998) );
  AOI21_X1 U11219 ( .B1(n10341), .B2(n10226), .A(n9998), .ZN(n10231) );
  INV_X1 U11220 ( .A(n10021), .ZN(n10001) );
  INV_X1 U11221 ( .A(n9999), .ZN(n10000) );
  AOI21_X1 U11222 ( .B1(n10227), .B2(n10001), .A(n10000), .ZN(n10229) );
  INV_X1 U11223 ( .A(n10002), .ZN(n10138) );
  NAND2_X1 U11224 ( .A1(n10229), .A2(n10138), .ZN(n10005) );
  AOI22_X1 U11225 ( .A1(n4377), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n10003), 
        .B2(n10358), .ZN(n10004) );
  OAI211_X1 U11226 ( .C1(n10006), .C2(n10123), .A(n10005), .B(n10004), .ZN(
        n10007) );
  AOI21_X1 U11227 ( .B1(n10346), .B2(n10226), .A(n10007), .ZN(n10008) );
  OAI21_X1 U11228 ( .B1(n10231), .B2(n4377), .A(n10008), .ZN(P1_U3282) );
  XNOR2_X1 U11229 ( .A(n10010), .B(n10009), .ZN(n10425) );
  INV_X1 U11230 ( .A(n10425), .ZN(n10028) );
  OAI21_X1 U11231 ( .B1(n10013), .B2(n10012), .A(n10011), .ZN(n10015) );
  NAND2_X1 U11232 ( .A1(n10015), .A2(n10014), .ZN(n10020) );
  AOI22_X1 U11233 ( .A1(n10018), .A2(n10356), .B1(n10017), .B2(n10016), .ZN(
        n10019) );
  NAND2_X1 U11234 ( .A1(n10020), .A2(n10019), .ZN(n10426) );
  OAI21_X1 U11235 ( .B1(n10041), .B2(n10423), .A(n10369), .ZN(n10022) );
  OR2_X1 U11236 ( .A1(n10022), .A2(n10021), .ZN(n10421) );
  AOI22_X1 U11237 ( .A1(n4377), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n4392), .B2(
        n10358), .ZN(n10025) );
  NAND2_X1 U11238 ( .A1(n10359), .A2(n10023), .ZN(n10024) );
  OAI211_X1 U11239 ( .C1(n10421), .C2(n10101), .A(n10025), .B(n10024), .ZN(
        n10026) );
  AOI21_X1 U11240 ( .B1(n10426), .B2(n10112), .A(n10026), .ZN(n10027) );
  OAI21_X1 U11241 ( .B1(n10028), .B2(n10124), .A(n10027), .ZN(P1_U3283) );
  INV_X1 U11242 ( .A(n10029), .ZN(n10032) );
  AOI21_X1 U11243 ( .B1(n10032), .B2(n10031), .A(n10030), .ZN(n10337) );
  NOR2_X1 U11244 ( .A1(n10337), .A2(n10336), .ZN(n10335) );
  OAI21_X1 U11245 ( .B1(n10335), .B2(n10034), .A(n10033), .ZN(n10035) );
  XOR2_X1 U11246 ( .A(n10038), .B(n10035), .Z(n10036) );
  OAI22_X1 U11247 ( .A1(n10036), .A2(n6464), .B1(n10334), .B2(n6460), .ZN(
        n10417) );
  INV_X1 U11248 ( .A(n10417), .ZN(n10054) );
  XNOR2_X1 U11249 ( .A(n10037), .B(n10038), .ZN(n10419) );
  NAND2_X1 U11250 ( .A1(n10039), .A2(n10050), .ZN(n10040) );
  NAND2_X1 U11251 ( .A1(n10040), .A2(n10369), .ZN(n10042) );
  OR2_X1 U11252 ( .A1(n10042), .A2(n10041), .ZN(n10045) );
  OR2_X1 U11253 ( .A1(n10043), .A2(n6461), .ZN(n10044) );
  AND2_X1 U11254 ( .A1(n10045), .A2(n10044), .ZN(n10415) );
  INV_X1 U11255 ( .A(n10046), .ZN(n10047) );
  OAI22_X1 U11256 ( .A1(n10112), .A2(n10048), .B1(n10047), .B2(n10097), .ZN(
        n10049) );
  AOI21_X1 U11257 ( .B1(n10359), .B2(n10050), .A(n10049), .ZN(n10051) );
  OAI21_X1 U11258 ( .B1(n10415), .B2(n10101), .A(n10051), .ZN(n10052) );
  AOI21_X1 U11259 ( .B1(n10373), .B2(n10419), .A(n10052), .ZN(n10053) );
  OAI21_X1 U11260 ( .B1(n10054), .B2(n4377), .A(n10053), .ZN(P1_U3284) );
  INV_X1 U11261 ( .A(n10335), .ZN(n10056) );
  NAND2_X1 U11262 ( .A1(n10056), .A2(n10055), .ZN(n10057) );
  XNOR2_X1 U11263 ( .A(n10057), .B(n10061), .ZN(n10059) );
  OAI222_X1 U11264 ( .A1(n6460), .A2(n10072), .B1(n10059), .B2(n6464), .C1(
        n6461), .C2(n10058), .ZN(n10411) );
  INV_X1 U11265 ( .A(n10411), .ZN(n10069) );
  XNOR2_X1 U11266 ( .A(n10060), .B(n10061), .ZN(n10413) );
  INV_X1 U11267 ( .A(n10344), .ZN(n10062) );
  OAI211_X1 U11268 ( .C1(n10062), .C2(n5986), .A(n10369), .B(n10039), .ZN(
        n10410) );
  AOI22_X1 U11269 ( .A1(n4377), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n10063), .B2(
        n10358), .ZN(n10066) );
  NAND2_X1 U11270 ( .A1(n10359), .A2(n10064), .ZN(n10065) );
  OAI211_X1 U11271 ( .C1(n10410), .C2(n10101), .A(n10066), .B(n10065), .ZN(
        n10067) );
  AOI21_X1 U11272 ( .B1(n10373), .B2(n10413), .A(n10067), .ZN(n10068) );
  OAI21_X1 U11273 ( .B1(n10069), .B2(n4377), .A(n10068), .ZN(P1_U3285) );
  XNOR2_X1 U11274 ( .A(n10029), .B(n10070), .ZN(n10071) );
  OAI222_X1 U11275 ( .A1(n6460), .A2(n10073), .B1(n6461), .B2(n10072), .C1(
        n6464), .C2(n10071), .ZN(n10398) );
  INV_X1 U11276 ( .A(n10398), .ZN(n10084) );
  XNOR2_X1 U11277 ( .A(n10075), .B(n10074), .ZN(n10400) );
  INV_X1 U11278 ( .A(n10368), .ZN(n10077) );
  INV_X1 U11279 ( .A(n10345), .ZN(n10076) );
  OAI211_X1 U11280 ( .C1(n10397), .C2(n10077), .A(n10076), .B(n10369), .ZN(
        n10396) );
  AOI22_X1 U11281 ( .A1(n4377), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n10078), .B2(
        n10358), .ZN(n10081) );
  NAND2_X1 U11282 ( .A1(n10359), .A2(n10079), .ZN(n10080) );
  OAI211_X1 U11283 ( .C1(n10396), .C2(n10101), .A(n10081), .B(n10080), .ZN(
        n10082) );
  AOI21_X1 U11284 ( .B1(n10373), .B2(n10400), .A(n10082), .ZN(n10083) );
  OAI21_X1 U11285 ( .B1(n10084), .B2(n4377), .A(n10083), .ZN(P1_U3287) );
  MUX2_X1 U11286 ( .A(n9051), .B(n10085), .S(n10112), .Z(n10092) );
  INV_X1 U11287 ( .A(n10086), .ZN(n10090) );
  INV_X1 U11288 ( .A(n10087), .ZN(n10088) );
  OAI22_X1 U11289 ( .A1(n10123), .A2(n5957), .B1(n10097), .B2(n10088), .ZN(
        n10089) );
  AOI21_X1 U11290 ( .B1(n10090), .B2(n10372), .A(n10089), .ZN(n10091) );
  OAI211_X1 U11291 ( .C1(n10124), .C2(n10093), .A(n10092), .B(n10091), .ZN(
        P1_U3289) );
  AOI21_X1 U11292 ( .B1(n10096), .B2(n10095), .A(n10094), .ZN(n10383) );
  INV_X1 U11293 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10098) );
  OAI22_X1 U11294 ( .A1(n10112), .A2(n10098), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n10097), .ZN(n10103) );
  OAI211_X1 U11295 ( .C1(n10100), .C2(n10385), .A(n10099), .B(n10369), .ZN(
        n10384) );
  NOR2_X1 U11296 ( .A1(n10101), .A2(n10384), .ZN(n10102) );
  AOI211_X1 U11297 ( .C1(n10359), .C2(n10104), .A(n10103), .B(n10102), .ZN(
        n10110) );
  XNOR2_X1 U11298 ( .A(n10106), .B(n10105), .ZN(n10107) );
  OAI222_X1 U11299 ( .A1(n6460), .A2(n10108), .B1(n10107), .B2(n6464), .C1(
        n6461), .C2(n10361), .ZN(n10386) );
  NAND2_X1 U11300 ( .A1(n10386), .A2(n10112), .ZN(n10109) );
  OAI211_X1 U11301 ( .C1(n10383), .C2(n10124), .A(n10110), .B(n10109), .ZN(
        P1_U3290) );
  INV_X1 U11302 ( .A(n10111), .ZN(n10119) );
  NAND2_X1 U11303 ( .A1(n10113), .A2(n10112), .ZN(n10118) );
  AOI22_X1 U11304 ( .A1(n4377), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10358), .ZN(n10114) );
  AOI21_X1 U11305 ( .B1(n10116), .B2(n10372), .A(n10115), .ZN(n10117) );
  OAI211_X1 U11306 ( .C1(n10119), .C2(n10124), .A(n10118), .B(n10117), .ZN(
        P1_U3291) );
  INV_X1 U11307 ( .A(n10120), .ZN(n10128) );
  AOI22_X1 U11308 ( .A1(n4377), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n10358), .ZN(n10121) );
  OAI21_X1 U11309 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(n10127) );
  NOR2_X1 U11310 ( .A1(n10125), .A2(n10124), .ZN(n10126) );
  AOI211_X1 U11311 ( .C1(n10128), .C2(n10372), .A(n10127), .B(n10126), .ZN(
        n10129) );
  OAI21_X1 U11312 ( .B1(n4377), .B2(n10130), .A(n10129), .ZN(P1_U3292) );
  INV_X1 U11313 ( .A(n10131), .ZN(n10132) );
  NOR3_X1 U11314 ( .A1(n10134), .A2(n10133), .A3(n10132), .ZN(n10135) );
  AOI211_X1 U11315 ( .C1(n10358), .C2(P1_REG3_REG_0__SCAN_IN), .A(n10136), .B(
        n10135), .ZN(n10141) );
  NAND2_X1 U11316 ( .A1(n4377), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10140) );
  OAI21_X1 U11317 ( .B1(n10138), .B2(n10359), .A(n10137), .ZN(n10139) );
  OAI211_X1 U11318 ( .C1(n10141), .C2(n4377), .A(n10140), .B(n10139), .ZN(
        P1_U3293) );
  AND2_X1 U11319 ( .A1(n10143), .A2(n10142), .ZN(n10234) );
  INV_X1 U11320 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10144) );
  MUX2_X1 U11321 ( .A(n10234), .B(n10144), .S(n10440), .Z(n10145) );
  OAI21_X1 U11322 ( .B1(n10236), .B2(n10194), .A(n10145), .ZN(P1_U3552) );
  INV_X1 U11323 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10149) );
  MUX2_X1 U11324 ( .A(n10149), .B(n10237), .S(n10442), .Z(n10150) );
  OAI21_X1 U11325 ( .B1(n10240), .B2(n10194), .A(n10150), .ZN(P1_U3548) );
  AOI211_X1 U11326 ( .C1(n10228), .C2(n10153), .A(n10152), .B(n10151), .ZN(
        n10154) );
  OAI21_X1 U11327 ( .B1(n10155), .B2(n10225), .A(n10154), .ZN(n10241) );
  MUX2_X1 U11328 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10241), .S(n10442), .Z(
        P1_U3547) );
  AOI211_X1 U11329 ( .C1(n10158), .C2(n10424), .A(n10157), .B(n10156), .ZN(
        n10242) );
  MUX2_X1 U11330 ( .A(n10159), .B(n10242), .S(n10442), .Z(n10160) );
  OAI21_X1 U11331 ( .B1(n10245), .B2(n10194), .A(n10160), .ZN(P1_U3546) );
  AOI211_X1 U11332 ( .C1(n10163), .C2(n10424), .A(n10162), .B(n10161), .ZN(
        n10246) );
  MUX2_X1 U11333 ( .A(n10164), .B(n10246), .S(n10442), .Z(n10165) );
  OAI21_X1 U11334 ( .B1(n10249), .B2(n10194), .A(n10165), .ZN(P1_U3545) );
  AOI211_X1 U11335 ( .C1(n10168), .C2(n10424), .A(n10167), .B(n10166), .ZN(
        n10250) );
  MUX2_X1 U11336 ( .A(n10169), .B(n10250), .S(n10442), .Z(n10170) );
  OAI21_X1 U11337 ( .B1(n10253), .B2(n10194), .A(n10170), .ZN(P1_U3544) );
  OR2_X1 U11338 ( .A1(n10171), .A2(n10225), .ZN(n10175) );
  NOR2_X1 U11339 ( .A1(n10173), .A2(n10172), .ZN(n10174) );
  NAND2_X1 U11340 ( .A1(n10175), .A2(n10174), .ZN(n10254) );
  MUX2_X1 U11341 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10254), .S(n10442), .Z(
        n10176) );
  AOI21_X1 U11342 ( .B1(n6526), .B2(n10256), .A(n10176), .ZN(n10177) );
  INV_X1 U11343 ( .A(n10177), .ZN(P1_U3543) );
  AOI211_X1 U11344 ( .C1(n10228), .C2(n10180), .A(n10179), .B(n10178), .ZN(
        n10181) );
  OAI21_X1 U11345 ( .B1(n10225), .B2(n10182), .A(n10181), .ZN(n10258) );
  MUX2_X1 U11346 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10258), .S(n10442), .Z(
        P1_U3542) );
  OAI211_X1 U11347 ( .C1(n10225), .C2(n10185), .A(n10184), .B(n10183), .ZN(
        n10186) );
  INV_X1 U11348 ( .A(n10186), .ZN(n10259) );
  MUX2_X1 U11349 ( .A(n10187), .B(n10259), .S(n10442), .Z(n10188) );
  OAI21_X1 U11350 ( .B1(n10262), .B2(n10194), .A(n10188), .ZN(P1_U3541) );
  INV_X1 U11351 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10192) );
  AOI211_X1 U11352 ( .C1(n10191), .C2(n10424), .A(n10190), .B(n10189), .ZN(
        n10263) );
  MUX2_X1 U11353 ( .A(n10192), .B(n10263), .S(n10442), .Z(n10193) );
  OAI21_X1 U11354 ( .B1(n10267), .B2(n10194), .A(n10193), .ZN(P1_U3540) );
  AOI211_X1 U11355 ( .C1(n10228), .C2(n10197), .A(n10196), .B(n10195), .ZN(
        n10198) );
  OAI21_X1 U11356 ( .B1(n10225), .B2(n10199), .A(n10198), .ZN(n10268) );
  MUX2_X1 U11357 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10268), .S(n10442), .Z(
        P1_U3539) );
  OR2_X1 U11358 ( .A1(n10200), .A2(n10225), .ZN(n10204) );
  NOR2_X1 U11359 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  NAND2_X1 U11360 ( .A1(n10204), .A2(n10203), .ZN(n10269) );
  MUX2_X1 U11361 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10269), .S(n10442), .Z(
        n10205) );
  AOI21_X1 U11362 ( .B1(n6526), .B2(n10271), .A(n10205), .ZN(n10206) );
  INV_X1 U11363 ( .A(n10206), .ZN(P1_U3538) );
  AOI21_X1 U11364 ( .B1(n10228), .B2(n10208), .A(n10207), .ZN(n10209) );
  OAI211_X1 U11365 ( .C1(n10225), .C2(n10211), .A(n10210), .B(n10209), .ZN(
        n10273) );
  MUX2_X1 U11366 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10273), .S(n10442), .Z(
        P1_U3537) );
  INV_X1 U11367 ( .A(n10212), .ZN(n10219) );
  INV_X1 U11368 ( .A(n10228), .ZN(n10422) );
  OAI22_X1 U11369 ( .A1(n10215), .A2(n10214), .B1(n10213), .B2(n10422), .ZN(
        n10216) );
  INV_X1 U11370 ( .A(n10216), .ZN(n10217) );
  OAI211_X1 U11371 ( .C1(n10219), .C2(n10401), .A(n10218), .B(n10217), .ZN(
        n10274) );
  MUX2_X1 U11372 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10274), .S(n10442), .Z(
        P1_U3536) );
  AOI211_X1 U11373 ( .C1(n10228), .C2(n10222), .A(n10221), .B(n10220), .ZN(
        n10223) );
  OAI21_X1 U11374 ( .B1(n10225), .B2(n10224), .A(n10223), .ZN(n10275) );
  MUX2_X1 U11375 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10275), .S(n10442), .Z(
        P1_U3535) );
  INV_X1 U11376 ( .A(n10226), .ZN(n10232) );
  AOI22_X1 U11377 ( .A1(n10229), .A2(n10369), .B1(n10228), .B2(n10227), .ZN(
        n10230) );
  OAI211_X1 U11378 ( .C1(n10401), .C2(n10232), .A(n10231), .B(n10230), .ZN(
        n10276) );
  MUX2_X1 U11379 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10276), .S(n10442), .Z(
        P1_U3533) );
  MUX2_X1 U11380 ( .A(n10234), .B(n10233), .S(n7114), .Z(n10235) );
  OAI21_X1 U11381 ( .B1(n10236), .B2(n10266), .A(n10235), .ZN(P1_U3520) );
  INV_X1 U11382 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10238) );
  MUX2_X1 U11383 ( .A(n10238), .B(n10237), .S(n10430), .Z(n10239) );
  OAI21_X1 U11384 ( .B1(n10240), .B2(n10266), .A(n10239), .ZN(P1_U3516) );
  MUX2_X1 U11385 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10241), .S(n10430), .Z(
        P1_U3515) );
  INV_X1 U11386 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10243) );
  MUX2_X1 U11387 ( .A(n10243), .B(n10242), .S(n10430), .Z(n10244) );
  OAI21_X1 U11388 ( .B1(n10245), .B2(n10266), .A(n10244), .ZN(P1_U3514) );
  INV_X1 U11389 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10247) );
  MUX2_X1 U11390 ( .A(n10247), .B(n10246), .S(n10430), .Z(n10248) );
  OAI21_X1 U11391 ( .B1(n10249), .B2(n10266), .A(n10248), .ZN(P1_U3513) );
  INV_X1 U11392 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10251) );
  MUX2_X1 U11393 ( .A(n10251), .B(n10250), .S(n10430), .Z(n10252) );
  OAI21_X1 U11394 ( .B1(n10253), .B2(n10266), .A(n10252), .ZN(P1_U3512) );
  MUX2_X1 U11395 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10254), .S(n10430), .Z(
        n10255) );
  AOI21_X1 U11396 ( .B1(n6140), .B2(n10256), .A(n10255), .ZN(n10257) );
  INV_X1 U11397 ( .A(n10257), .ZN(P1_U3511) );
  MUX2_X1 U11398 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10258), .S(n10430), .Z(
        P1_U3510) );
  MUX2_X1 U11399 ( .A(n10260), .B(n10259), .S(n10430), .Z(n10261) );
  OAI21_X1 U11400 ( .B1(n10262), .B2(n10266), .A(n10261), .ZN(P1_U3509) );
  INV_X1 U11401 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10264) );
  MUX2_X1 U11402 ( .A(n10264), .B(n10263), .S(n10430), .Z(n10265) );
  OAI21_X1 U11403 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(P1_U3507) );
  MUX2_X1 U11404 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10268), .S(n10430), .Z(
        P1_U3504) );
  MUX2_X1 U11405 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10269), .S(n10430), .Z(
        n10270) );
  AOI21_X1 U11406 ( .B1(n6140), .B2(n10271), .A(n10270), .ZN(n10272) );
  INV_X1 U11407 ( .A(n10272), .ZN(P1_U3501) );
  MUX2_X1 U11408 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10273), .S(n10430), .Z(
        P1_U3498) );
  MUX2_X1 U11409 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10274), .S(n10430), .Z(
        P1_U3495) );
  MUX2_X1 U11410 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10275), .S(n10430), .Z(
        P1_U3492) );
  MUX2_X1 U11411 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10276), .S(n10430), .Z(
        P1_U3486) );
  MUX2_X1 U11412 ( .A(n10277), .B(P1_D_REG_0__SCAN_IN), .S(n10381), .Z(
        P1_U3439) );
  NOR4_X1 U11413 ( .A1(n10279), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10278), .A4(
        P1_U3086), .ZN(n10280) );
  AOI21_X1 U11414 ( .B1(n10281), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10280), 
        .ZN(n10282) );
  OAI21_X1 U11415 ( .B1(n10284), .B2(n10283), .A(n10282), .ZN(P1_U3324) );
  MUX2_X1 U11416 ( .A(n10285), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11417 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11418 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11419 ( .B1(n10288), .B2(n10287), .A(n10286), .ZN(n10297) );
  OAI21_X1 U11420 ( .B1(n10290), .B2(n10289), .A(n10319), .ZN(n10291) );
  OR2_X1 U11421 ( .A1(n10292), .A2(n10291), .ZN(n10295) );
  NAND2_X1 U11422 ( .A1(n10312), .A2(n10293), .ZN(n10294) );
  OAI211_X1 U11423 ( .C1(n10297), .C2(n10296), .A(n10295), .B(n10294), .ZN(
        n10298) );
  INV_X1 U11424 ( .A(n10298), .ZN(n10300) );
  OAI211_X1 U11425 ( .C1(n10301), .C2(n10332), .A(n10300), .B(n10299), .ZN(
        P1_U3257) );
  AOI211_X1 U11426 ( .C1(n10305), .C2(n10304), .A(n10303), .B(n10302), .ZN(
        n10310) );
  AOI211_X1 U11427 ( .C1(n10308), .C2(n10307), .A(n10306), .B(n10316), .ZN(
        n10309) );
  AOI211_X1 U11428 ( .C1(n10312), .C2(n10311), .A(n10310), .B(n10309), .ZN(
        n10314) );
  OAI211_X1 U11429 ( .C1(n10315), .C2(n10332), .A(n10314), .B(n10313), .ZN(
        P1_U3258) );
  AOI21_X1 U11430 ( .B1(n10318), .B2(n10317), .A(n10316), .ZN(n10328) );
  OAI211_X1 U11431 ( .C1(n10322), .C2(n10321), .A(n10320), .B(n10319), .ZN(
        n10323) );
  OAI21_X1 U11432 ( .B1(n10325), .B2(n10324), .A(n10323), .ZN(n10326) );
  AOI21_X1 U11433 ( .B1(n10328), .B2(n10327), .A(n10326), .ZN(n10330) );
  OAI211_X1 U11434 ( .C1(n10332), .C2(n10331), .A(n10330), .B(n10329), .ZN(
        P1_U3261) );
  XNOR2_X1 U11435 ( .A(n10333), .B(n10336), .ZN(n10407) );
  OAI22_X1 U11436 ( .A1(n10334), .A2(n6461), .B1(n10350), .B2(n6460), .ZN(
        n10340) );
  AOI21_X1 U11437 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(n10338) );
  NOR2_X1 U11438 ( .A1(n10338), .A2(n6464), .ZN(n10339) );
  AOI211_X1 U11439 ( .C1(n10341), .C2(n10407), .A(n10340), .B(n10339), .ZN(
        n10404) );
  AOI222_X1 U11440 ( .A1(n10343), .A2(n10359), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n4377), .C1(n10358), .C2(n10342), .ZN(n10349) );
  OAI211_X1 U11441 ( .C1(n10345), .C2(n10403), .A(n10344), .B(n10369), .ZN(
        n10402) );
  INV_X1 U11442 ( .A(n10402), .ZN(n10347) );
  AOI22_X1 U11443 ( .A1(n10372), .A2(n10347), .B1(n10407), .B2(n10346), .ZN(
        n10348) );
  OAI211_X1 U11444 ( .C1(n4377), .C2(n10404), .A(n10349), .B(n10348), .ZN(
        P1_U3286) );
  NOR2_X1 U11445 ( .A1(n10350), .A2(n6461), .ZN(n10355) );
  INV_X1 U11446 ( .A(n6472), .ZN(n10351) );
  NOR2_X1 U11447 ( .A1(n10352), .A2(n10351), .ZN(n10353) );
  AOI211_X1 U11448 ( .C1(n5019), .C2(n10366), .A(n6464), .B(n10353), .ZN(
        n10354) );
  AOI211_X1 U11449 ( .C1(n10356), .C2(n10364), .A(n10355), .B(n10354), .ZN(
        n10391) );
  AOI222_X1 U11450 ( .A1(n10360), .A2(n10359), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n4377), .C1(n10358), .C2(n10357), .ZN(n10375) );
  INV_X1 U11451 ( .A(n10365), .ZN(n10362) );
  OAI21_X1 U11452 ( .B1(n10362), .B2(n10361), .A(n5957), .ZN(n10363) );
  OAI21_X1 U11453 ( .B1(n10365), .B2(n10364), .A(n10363), .ZN(n10367) );
  XNOR2_X1 U11454 ( .A(n10367), .B(n10366), .ZN(n10394) );
  INV_X1 U11455 ( .A(n7759), .ZN(n10370) );
  OAI211_X1 U11456 ( .C1(n10370), .C2(n10392), .A(n10369), .B(n10368), .ZN(
        n10390) );
  INV_X1 U11457 ( .A(n10390), .ZN(n10371) );
  AOI22_X1 U11458 ( .A1(n10394), .A2(n10373), .B1(n10372), .B2(n10371), .ZN(
        n10374) );
  OAI211_X1 U11459 ( .C1(n4377), .C2(n10391), .A(n10375), .B(n10374), .ZN(
        P1_U3288) );
  AND2_X1 U11460 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10381), .ZN(P1_U3294) );
  AND2_X1 U11461 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10381), .ZN(P1_U3295) );
  AND2_X1 U11462 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10381), .ZN(P1_U3296) );
  AND2_X1 U11463 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10381), .ZN(P1_U3297) );
  NOR2_X1 U11464 ( .A1(n10380), .A2(n10376), .ZN(P1_U3298) );
  AND2_X1 U11465 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10381), .ZN(P1_U3299) );
  AND2_X1 U11466 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10381), .ZN(P1_U3300) );
  AND2_X1 U11467 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10381), .ZN(P1_U3301) );
  INV_X1 U11468 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10377) );
  NOR2_X1 U11469 ( .A1(n10380), .A2(n10377), .ZN(P1_U3302) );
  NOR2_X1 U11470 ( .A1(n10380), .A2(n10378), .ZN(P1_U3303) );
  AND2_X1 U11471 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10381), .ZN(P1_U3304) );
  AND2_X1 U11472 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10381), .ZN(P1_U3305) );
  AND2_X1 U11473 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10381), .ZN(P1_U3306) );
  AND2_X1 U11474 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10381), .ZN(P1_U3307) );
  AND2_X1 U11475 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10381), .ZN(P1_U3308) );
  AND2_X1 U11476 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10381), .ZN(P1_U3309) );
  AND2_X1 U11477 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10381), .ZN(P1_U3310) );
  AND2_X1 U11478 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10381), .ZN(P1_U3311) );
  AND2_X1 U11479 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10381), .ZN(P1_U3312) );
  AND2_X1 U11480 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10381), .ZN(P1_U3313) );
  AND2_X1 U11481 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10381), .ZN(P1_U3314) );
  AND2_X1 U11482 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10381), .ZN(P1_U3315) );
  AND2_X1 U11483 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10381), .ZN(P1_U3316) );
  AND2_X1 U11484 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10381), .ZN(P1_U3317) );
  AND2_X1 U11485 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10381), .ZN(P1_U3318) );
  NOR2_X1 U11486 ( .A1(n10380), .A2(n10379), .ZN(P1_U3319) );
  AND2_X1 U11487 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10381), .ZN(P1_U3320) );
  AND2_X1 U11488 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10381), .ZN(P1_U3321) );
  AND2_X1 U11489 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10381), .ZN(P1_U3322) );
  AND2_X1 U11490 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10381), .ZN(P1_U3323) );
  AOI22_X1 U11491 ( .A1(n10430), .A2(n10382), .B1(n6258), .B2(n7114), .ZN(
        P1_U3453) );
  INV_X1 U11492 ( .A(n10383), .ZN(n10388) );
  OAI21_X1 U11493 ( .B1(n10385), .B2(n10422), .A(n10384), .ZN(n10387) );
  AOI211_X1 U11494 ( .C1(n10424), .C2(n10388), .A(n10387), .B(n10386), .ZN(
        n10432) );
  INV_X1 U11495 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U11496 ( .A1(n10430), .A2(n10432), .B1(n10389), .B2(n7114), .ZN(
        P1_U3462) );
  OAI211_X1 U11497 ( .C1(n10392), .C2(n10422), .A(n10391), .B(n10390), .ZN(
        n10393) );
  AOI21_X1 U11498 ( .B1(n10424), .B2(n10394), .A(n10393), .ZN(n10433) );
  AOI22_X1 U11499 ( .A1(n10430), .A2(n10433), .B1(n10395), .B2(n7114), .ZN(
        P1_U3468) );
  OAI21_X1 U11500 ( .B1(n10397), .B2(n10422), .A(n10396), .ZN(n10399) );
  AOI211_X1 U11501 ( .C1(n10424), .C2(n10400), .A(n10399), .B(n10398), .ZN(
        n10434) );
  AOI22_X1 U11502 ( .A1(n10430), .A2(n10434), .B1(n4778), .B2(n7114), .ZN(
        P1_U3471) );
  INV_X1 U11503 ( .A(n10401), .ZN(n10408) );
  OAI21_X1 U11504 ( .B1(n10403), .B2(n10422), .A(n10402), .ZN(n10406) );
  INV_X1 U11505 ( .A(n10404), .ZN(n10405) );
  AOI211_X1 U11506 ( .C1(n10408), .C2(n10407), .A(n10406), .B(n10405), .ZN(
        n10435) );
  AOI22_X1 U11507 ( .A1(n10430), .A2(n10435), .B1(n10409), .B2(n7114), .ZN(
        P1_U3474) );
  OAI21_X1 U11508 ( .B1(n5986), .B2(n10422), .A(n10410), .ZN(n10412) );
  AOI211_X1 U11509 ( .C1(n10424), .C2(n10413), .A(n10412), .B(n10411), .ZN(
        n10437) );
  INV_X1 U11510 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U11511 ( .A1(n10430), .A2(n10437), .B1(n10414), .B2(n7114), .ZN(
        P1_U3477) );
  OAI21_X1 U11512 ( .B1(n10416), .B2(n10422), .A(n10415), .ZN(n10418) );
  AOI211_X1 U11513 ( .C1(n10424), .C2(n10419), .A(n10418), .B(n10417), .ZN(
        n10439) );
  INV_X1 U11514 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U11515 ( .A1(n10430), .A2(n10439), .B1(n10420), .B2(n7114), .ZN(
        P1_U3480) );
  OAI21_X1 U11516 ( .B1(n10423), .B2(n10422), .A(n10421), .ZN(n10428) );
  AND2_X1 U11517 ( .A1(n10425), .A2(n10424), .ZN(n10427) );
  NOR3_X1 U11518 ( .A1(n10428), .A2(n10427), .A3(n10426), .ZN(n10441) );
  AOI22_X1 U11519 ( .A1(n10430), .A2(n10441), .B1(n10429), .B2(n7114), .ZN(
        P1_U3483) );
  INV_X1 U11520 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U11521 ( .A1(n10442), .A2(n10432), .B1(n10431), .B2(n10440), .ZN(
        P1_U3525) );
  AOI22_X1 U11522 ( .A1(n10442), .A2(n10433), .B1(n7235), .B2(n10440), .ZN(
        P1_U3527) );
  AOI22_X1 U11523 ( .A1(n10442), .A2(n10434), .B1(n7237), .B2(n10440), .ZN(
        P1_U3528) );
  AOI22_X1 U11524 ( .A1(n10442), .A2(n10435), .B1(n7239), .B2(n10440), .ZN(
        P1_U3529) );
  AOI22_X1 U11525 ( .A1(n10442), .A2(n10437), .B1(n10436), .B2(n10440), .ZN(
        P1_U3530) );
  AOI22_X1 U11526 ( .A1(n10442), .A2(n10439), .B1(n10438), .B2(n10440), .ZN(
        P1_U3531) );
  AOI22_X1 U11527 ( .A1(n10442), .A2(n10441), .B1(n7253), .B2(n10440), .ZN(
        P1_U3532) );
  AOI22_X1 U11528 ( .A1(n10448), .A2(n10444), .B1(n10443), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n10455) );
  MUX2_X1 U11529 ( .A(n10447), .B(n10446), .S(n4383), .Z(n10449) );
  NOR2_X1 U11530 ( .A1(n10449), .A2(n10448), .ZN(n10450) );
  OAI22_X1 U11531 ( .A1(n10453), .A2(n10452), .B1(n10451), .B2(n10450), .ZN(
        n10454) );
  OAI211_X1 U11532 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5283), .A(n10455), .B(
        n10454), .ZN(P2_U3182) );
  OAI22_X1 U11533 ( .A1(n10458), .A2(n5299), .B1(n10457), .B2(n10456), .ZN(
        n10461) );
  INV_X1 U11534 ( .A(n10459), .ZN(n10460) );
  AOI211_X1 U11535 ( .C1(n10463), .C2(n10462), .A(n10461), .B(n10460), .ZN(
        n10465) );
  AOI22_X1 U11536 ( .A1(n10466), .A2(n6566), .B1(n10465), .B2(n10464), .ZN(
        P2_U3231) );
  INV_X1 U11537 ( .A(n10467), .ZN(n10468) );
  AOI21_X1 U11538 ( .B1(n10497), .B2(n10469), .A(n10468), .ZN(n10470) );
  AOI211_X1 U11539 ( .C1(n10473), .C2(n10472), .A(n10471), .B(n10470), .ZN(
        n10502) );
  AOI22_X1 U11540 ( .A1(n10501), .A2(n10502), .B1(n5282), .B2(n10499), .ZN(
        P2_U3390) );
  INV_X1 U11541 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U11542 ( .A1(n10501), .A2(n10475), .B1(n10474), .B2(n10499), .ZN(
        P2_U3393) );
  AOI22_X1 U11543 ( .A1(n10501), .A2(n10476), .B1(n5296), .B2(n10499), .ZN(
        P2_U3396) );
  INV_X1 U11544 ( .A(n10477), .ZN(n10481) );
  INV_X1 U11545 ( .A(n10478), .ZN(n10479) );
  AOI211_X1 U11546 ( .C1(n10481), .C2(n10487), .A(n10480), .B(n10479), .ZN(
        n10503) );
  AOI22_X1 U11547 ( .A1(n10501), .A2(n10503), .B1(n5313), .B2(n10499), .ZN(
        P2_U3399) );
  INV_X1 U11548 ( .A(n10482), .ZN(n10486) );
  INV_X1 U11549 ( .A(n10483), .ZN(n10484) );
  AOI211_X1 U11550 ( .C1(n10487), .C2(n10486), .A(n10485), .B(n10484), .ZN(
        n10504) );
  AOI22_X1 U11551 ( .A1(n10501), .A2(n10504), .B1(n5335), .B2(n10499), .ZN(
        P2_U3402) );
  NOR2_X1 U11552 ( .A1(n10489), .A2(n10488), .ZN(n10491) );
  AOI211_X1 U11553 ( .C1(n10493), .C2(n10492), .A(n10491), .B(n10490), .ZN(
        n10506) );
  AOI22_X1 U11554 ( .A1(n10501), .A2(n10506), .B1(n5356), .B2(n10499), .ZN(
        P2_U3405) );
  OAI211_X1 U11555 ( .C1(n10497), .C2(n10496), .A(n10495), .B(n10494), .ZN(
        n10498) );
  INV_X1 U11556 ( .A(n10498), .ZN(n10507) );
  INV_X1 U11557 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U11558 ( .A1(n10501), .A2(n10507), .B1(n10500), .B2(n10499), .ZN(
        P2_U3408) );
  AOI22_X1 U11559 ( .A1(n10508), .A2(n10502), .B1(n10446), .B2(n7125), .ZN(
        P2_U3459) );
  AOI22_X1 U11560 ( .A1(n10508), .A2(n10503), .B1(n5314), .B2(n7125), .ZN(
        P2_U3462) );
  AOI22_X1 U11561 ( .A1(n10508), .A2(n10504), .B1(n6598), .B2(n7125), .ZN(
        P2_U3463) );
  INV_X1 U11562 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10505) );
  AOI22_X1 U11563 ( .A1(n10508), .A2(n10506), .B1(n10505), .B2(n7125), .ZN(
        P2_U3464) );
  AOI22_X1 U11564 ( .A1(n10508), .A2(n10507), .B1(n6639), .B2(n7125), .ZN(
        P2_U3465) );
  OAI222_X1 U11565 ( .A1(n10513), .A2(n10512), .B1(n10513), .B2(n10511), .C1(
        n10510), .C2(n10509), .ZN(ADD_1068_U5) );
  XOR2_X1 U11566 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  INV_X1 U11567 ( .A(n10516), .ZN(n10515) );
  OAI222_X1 U11568 ( .A1(n10518), .A2(n10517), .B1(n10518), .B2(n10516), .C1(
        n10515), .C2(n10514), .ZN(ADD_1068_U55) );
  OAI21_X1 U11569 ( .B1(n10521), .B2(n10520), .A(n10519), .ZN(ADD_1068_U56) );
  OAI21_X1 U11570 ( .B1(n10524), .B2(n10523), .A(n10522), .ZN(ADD_1068_U57) );
  OAI21_X1 U11571 ( .B1(n10527), .B2(n10526), .A(n10525), .ZN(ADD_1068_U58) );
  OAI21_X1 U11572 ( .B1(n10530), .B2(n10529), .A(n10528), .ZN(ADD_1068_U59) );
  OAI21_X1 U11573 ( .B1(n10533), .B2(n10532), .A(n10531), .ZN(ADD_1068_U60) );
  OAI21_X1 U11574 ( .B1(n10536), .B2(n10535), .A(n10534), .ZN(ADD_1068_U61) );
  OAI21_X1 U11575 ( .B1(n10539), .B2(n10538), .A(n10537), .ZN(ADD_1068_U62) );
  OAI21_X1 U11576 ( .B1(n10542), .B2(n10541), .A(n10540), .ZN(ADD_1068_U63) );
  OAI21_X1 U11577 ( .B1(n10545), .B2(n10544), .A(n10543), .ZN(ADD_1068_U51) );
  OAI21_X1 U11578 ( .B1(n10548), .B2(n10547), .A(n10546), .ZN(ADD_1068_U50) );
  OAI21_X1 U11579 ( .B1(n10551), .B2(n10550), .A(n10549), .ZN(ADD_1068_U47) );
  OAI21_X1 U11580 ( .B1(n10554), .B2(n10553), .A(n10552), .ZN(ADD_1068_U49) );
  OAI21_X1 U11581 ( .B1(n10557), .B2(n10556), .A(n10555), .ZN(ADD_1068_U48) );
  AOI21_X1 U11582 ( .B1(n10560), .B2(n10559), .A(n10558), .ZN(ADD_1068_U54) );
  AOI21_X1 U11583 ( .B1(n10563), .B2(n10562), .A(n10561), .ZN(ADD_1068_U53) );
  OAI21_X1 U11584 ( .B1(n10566), .B2(n10565), .A(n10564), .ZN(ADD_1068_U52) );
  CLKBUF_X2 U5043 ( .A(n6467), .Z(n4391) );
endmodule

