

module b21_C_AntiSAT_k_128_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067;

  INV_X4 U4810 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  XNOR2_X1 U4811 ( .A(n9141), .B(n9140), .ZN(n7314) );
  AOI21_X1 U4812 ( .B1(n5839), .B2(P1_REG1_REG_2__SCAN_IN), .A(n9580), .ZN(
        n5842) );
  CLKBUF_X2 U4813 ( .A(n5117), .Z(n8240) );
  INV_X1 U4814 ( .A(n8442), .ZN(n8435) );
  INV_X2 U4816 ( .A(n6095), .ZN(n8482) );
  OAI21_X1 U4817 ( .B1(n9659), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9663), .ZN(
        n9140) );
  INV_X1 U4818 ( .A(n5614), .ZN(n8173) );
  INV_X1 U4819 ( .A(n5147), .ZN(n5464) );
  OR2_X1 U4820 ( .A1(n7558), .A2(n8927), .ZN(n7616) );
  INV_X1 U4821 ( .A(n7750), .ZN(n7822) );
  NOR2_X1 U4822 ( .A1(n9582), .A2(n9581), .ZN(n9580) );
  AND2_X1 U4823 ( .A1(n9625), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9614) );
  INV_X1 U4824 ( .A(n6169), .ZN(n9695) );
  NAND2_X1 U4825 ( .A1(n6417), .A2(n6457), .ZN(n8028) );
  NAND2_X1 U4826 ( .A1(n4760), .A2(n4761), .ZN(n5024) );
  INV_X1 U4828 ( .A(n5929), .ZN(n8109) );
  OAI22_X1 U4829 ( .A1(n9614), .A2(n9628), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n9625), .ZN(n9640) );
  XNOR2_X1 U4830 ( .A(n5661), .B(n5660), .ZN(n9591) );
  INV_X2 U4831 ( .A(n4469), .ZN(n5419) );
  AOI21_X2 U4832 ( .B1(n7024), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6592), .ZN(
        n6595) );
  OAI21_X2 U4833 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n4903), .ZN(n4761) );
  AND2_X4 U4834 ( .A1(n9491), .A2(n5707), .ZN(n7244) );
  OAI222_X1 U4835 ( .A1(P2_U3152), .A2(n4894), .B1(n8980), .B2(n9492), .C1(
        n9989), .C2(n8979), .ZN(P2_U3328) );
  AND2_X4 U4836 ( .A1(n4894), .A2(n4895), .ZN(n5086) );
  XNOR2_X2 U4837 ( .A(n4890), .B(n8974), .ZN(n4894) );
  AND2_X1 U4838 ( .A1(n4749), .A2(n4747), .ZN(n8545) );
  AND2_X1 U4839 ( .A1(n4809), .A2(n4796), .ZN(n4795) );
  AOI21_X1 U4840 ( .B1(n4380), .B2(n8817), .A(n5515), .ZN(n7709) );
  AND3_X1 U4841 ( .A1(n4815), .A2(n4322), .A3(n4810), .ZN(n8982) );
  NAND2_X1 U4842 ( .A1(n4440), .A2(n9078), .ZN(n8993) );
  OAI22_X1 U4843 ( .A1(n9245), .A2(n4613), .B1(n4615), .B2(n4612), .ZN(n9203)
         );
  NAND2_X1 U4844 ( .A1(n4826), .A2(n8512), .ZN(n4825) );
  NOR2_X1 U4845 ( .A1(n7502), .A2(n8390), .ZN(n7501) );
  NAND2_X1 U4846 ( .A1(n8512), .A2(n4828), .ZN(n4827) );
  NAND2_X1 U4847 ( .A1(n7385), .A2(n7384), .ZN(n7386) );
  OAI22_X2 U4848 ( .A1(n9361), .A2(n8125), .B1(n4517), .B2(n8124), .ZN(n9340)
         );
  NAND2_X1 U4849 ( .A1(n4383), .A2(n7366), .ZN(n7385) );
  NAND2_X1 U4850 ( .A1(n4633), .A2(n4367), .ZN(n8123) );
  NAND2_X1 U4851 ( .A1(n4439), .A2(n4343), .ZN(n7182) );
  NAND2_X1 U4852 ( .A1(n6984), .A2(n6983), .ZN(n4383) );
  NAND2_X1 U4853 ( .A1(n6886), .A2(n6885), .ZN(n6984) );
  NAND2_X1 U4854 ( .A1(n7454), .A2(n4634), .ZN(n4633) );
  INV_X1 U4855 ( .A(n7337), .ZN(n4637) );
  NAND2_X1 U4856 ( .A1(n7107), .A2(n8267), .ZN(n7170) );
  NAND2_X1 U4857 ( .A1(n4838), .A2(n4837), .ZN(n6659) );
  AND2_X1 U4858 ( .A1(n6817), .A2(n5193), .ZN(n7650) );
  OR2_X1 U4859 ( .A1(n7496), .A2(n9105), .ZN(n4634) );
  NOR2_X1 U4860 ( .A1(n9106), .A2(n7832), .ZN(n4635) );
  NAND2_X1 U4861 ( .A1(n7140), .A2(n7139), .ZN(n7236) );
  NAND2_X1 U4862 ( .A1(n7026), .A2(n7025), .ZN(n9464) );
  NAND2_X1 U4863 ( .A1(n5201), .A2(n5200), .ZN(n5207) );
  INV_X1 U4864 ( .A(n6697), .ZN(n6677) );
  NAND2_X1 U4865 ( .A1(n5634), .A2(n9742), .ZN(n8583) );
  NAND2_X2 U4866 ( .A1(n8298), .A2(n8321), .ZN(n8255) );
  OR2_X1 U4867 ( .A1(n6024), .A2(n6023), .ZN(n4530) );
  NAND2_X1 U4868 ( .A1(n9695), .A2(n9117), .ZN(n6457) );
  AND3_X1 U4869 ( .A1(n5113), .A2(n5112), .A3(n5111), .ZN(n6555) );
  INV_X2 U4870 ( .A(n8250), .ZN(n8187) );
  NAND2_X1 U4871 ( .A1(n4716), .A2(n6216), .ZN(n5614) );
  INV_X1 U4872 ( .A(n9117), .ZN(n6456) );
  XNOR2_X1 U4873 ( .A(n5583), .B(n5582), .ZN(n5929) );
  INV_X2 U4874 ( .A(n6067), .ZN(n7896) );
  NAND4_X1 U4875 ( .A1(n5107), .A2(n5106), .A3(n5105), .A4(n5104), .ZN(n8638)
         );
  INV_X1 U4876 ( .A(n7676), .ZN(n6391) );
  INV_X2 U4877 ( .A(n4680), .ZN(n7869) );
  AND4_X1 U4878 ( .A1(n5068), .A2(n5067), .A3(n5066), .A4(n5065), .ZN(n6771)
         );
  INV_X1 U4879 ( .A(n4680), .ZN(n4305) );
  XNOR2_X1 U4880 ( .A(n5566), .B(n5565), .ZN(n7400) );
  INV_X1 U4881 ( .A(n5706), .ZN(n9491) );
  XNOR2_X1 U4882 ( .A(n5592), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U4883 ( .A1(n5699), .A2(n5698), .ZN(n7639) );
  XNOR2_X1 U4884 ( .A(n5695), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5706) );
  MUX2_X1 U4885 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5697), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5699) );
  NAND2_X1 U4886 ( .A1(n5698), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5695) );
  NAND2_X2 U4887 ( .A1(n7725), .A2(P1_U3084), .ZN(n9495) );
  AND3_X1 U4889 ( .A1(n4710), .A2(n5561), .A3(n4317), .ZN(n5696) );
  NOR2_X1 U4890 ( .A1(n4346), .A2(n4840), .ZN(n4839) );
  AND3_X1 U4891 ( .A1(n4359), .A2(n5564), .A3(n4855), .ZN(n4710) );
  AND2_X1 U4892 ( .A1(n5570), .A2(n5574), .ZN(n4847) );
  AND2_X1 U4893 ( .A1(n4876), .A2(n4875), .ZN(n5123) );
  NOR3_X1 U4894 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n5559) );
  INV_X1 U4895 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5478) );
  INV_X1 U4896 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6245) );
  INV_X1 U4897 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5886) );
  INV_X1 U4898 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5584) );
  INV_X1 U4899 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5574) );
  INV_X1 U4900 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10016) );
  INV_X1 U4901 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5224) );
  INV_X1 U4902 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5225) );
  INV_X1 U4903 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5166) );
  INV_X1 U4904 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6153) );
  NOR2_X1 U4905 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4876) );
  NOR2_X1 U4906 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4875) );
  INV_X4 U4907 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U4908 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5558) );
  NOR2_X1 U4909 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5557) );
  INV_X4 U4910 ( .A(n7868), .ZN(n7346) );
  OAI21_X2 U4911 ( .B1(n6119), .B2(n6067), .A(n4353), .ZN(n6515) );
  XNOR2_X2 U4912 ( .A(n4381), .B(n5021), .ZN(n5509) );
  NAND2_X1 U4913 ( .A1(n5944), .A2(n7725), .ZN(n4306) );
  AND2_X4 U4914 ( .A1(n5925), .A2(n6132), .ZN(n5930) );
  XNOR2_X2 U4915 ( .A(n9118), .B(n9071), .ZN(n8033) );
  OAI211_X1 U4916 ( .C1(n5944), .C2(n9591), .A(n5991), .B(n5990), .ZN(n9071)
         );
  OAI22_X2 U4917 ( .A1(n6863), .A2(n6862), .B1(n9111), .B2(n6861), .ZN(n7022)
         );
  NAND2_X2 U4918 ( .A1(n6778), .A2(n6777), .ZN(n6863) );
  NOR2_X1 U4919 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4879) );
  XNOR2_X1 U4920 ( .A(n5391), .B(SI_24_), .ZN(n5386) );
  OAI21_X1 U4921 ( .B1(n5046), .B2(n4991), .A(n4990), .ZN(n5035) );
  NAND2_X1 U4922 ( .A1(n5996), .A2(n5995), .ZN(n9355) );
  AOI21_X1 U4923 ( .B1(n9191), .B2(n7346), .A(n7893), .ZN(n9208) );
  AOI21_X1 U4924 ( .B1(n8340), .B2(n8442), .A(n4480), .ZN(n4479) );
  AND2_X1 U4925 ( .A1(n8341), .A2(n8435), .ZN(n4480) );
  NOR2_X1 U4926 ( .A1(n4653), .A2(n4652), .ZN(n4651) );
  INV_X1 U4927 ( .A(SI_16_), .ZN(n4981) );
  NAND2_X1 U4928 ( .A1(n4572), .A2(n4333), .ZN(n4940) );
  INV_X1 U4929 ( .A(n5162), .ZN(n4571) );
  NOR2_X1 U4930 ( .A1(n7372), .A2(n7371), .ZN(n7373) );
  INV_X1 U4931 ( .A(n6885), .ZN(n4726) );
  NOR2_X1 U4932 ( .A1(n4662), .A2(n4791), .ZN(n4790) );
  INV_X1 U4933 ( .A(n4852), .ZN(n4791) );
  AND2_X1 U4934 ( .A1(n4779), .A2(n4778), .ZN(n4776) );
  NAND2_X1 U4935 ( .A1(n8927), .A2(n8623), .ZN(n4783) );
  NAND2_X1 U4936 ( .A1(n7128), .A2(n7108), .ZN(n8362) );
  OR2_X1 U4937 ( .A1(n5207), .A2(n6819), .ZN(n8337) );
  AND2_X1 U4938 ( .A1(n6479), .A2(n6741), .ZN(n5487) );
  AND2_X1 U4939 ( .A1(n8317), .A2(n8316), .ZN(n8253) );
  OR2_X1 U4940 ( .A1(n8519), .A2(n4812), .ZN(n4811) );
  NOR2_X1 U4941 ( .A1(n9059), .A2(n4812), .ZN(n4798) );
  NAND2_X1 U4942 ( .A1(n9237), .A2(n9250), .ZN(n4622) );
  OR2_X1 U4943 ( .A1(n9418), .A2(n9034), .ZN(n8149) );
  INV_X1 U4944 ( .A(n4604), .ZN(n4603) );
  OAI21_X1 U4945 ( .B1(n4607), .B2(n4605), .A(n8126), .ZN(n4604) );
  AND2_X1 U4946 ( .A1(n5899), .A2(n8097), .ZN(n5960) );
  NAND2_X1 U4947 ( .A1(n5461), .A2(n5460), .ZN(n7711) );
  NAND2_X1 U4948 ( .A1(n5428), .A2(n5427), .ZN(n5441) );
  AND4_X1 U4949 ( .A1(n5578), .A2(n5584), .A3(n6153), .A4(n5577), .ZN(n5564)
         );
  NAND2_X1 U4950 ( .A1(n5005), .A2(n5004), .ZN(n5346) );
  INV_X1 U4951 ( .A(n5576), .ZN(n4841) );
  OAI21_X1 U4952 ( .B1(n6635), .B2(n4396), .A(n4393), .ZN(n6734) );
  AND2_X1 U4953 ( .A1(n4752), .A2(n4394), .ZN(n4393) );
  AND2_X1 U4954 ( .A1(n5628), .A2(n5621), .ZN(n4752) );
  NAND2_X1 U4955 ( .A1(n4395), .A2(n6636), .ZN(n4394) );
  AND2_X1 U4956 ( .A1(n6806), .A2(n5610), .ZN(n4721) );
  NAND2_X1 U4957 ( .A1(n9763), .A2(n4382), .ZN(n8250) );
  INV_X1 U4958 ( .A(n8453), .ZN(n4382) );
  NAND2_X1 U4959 ( .A1(n4476), .A2(n8282), .ZN(n4475) );
  NAND2_X1 U4960 ( .A1(n4478), .A2(n4477), .ZN(n4476) );
  INV_X1 U4961 ( .A(n8445), .ZN(n4477) );
  NAND2_X1 U4962 ( .A1(n8446), .A2(n8447), .ZN(n4478) );
  AND2_X1 U4963 ( .A1(n4901), .A2(n4900), .ZN(n8586) );
  INV_X1 U4964 ( .A(n5215), .ZN(n8237) );
  INV_X1 U4965 ( .A(n4894), .ZN(n4893) );
  NAND2_X1 U4966 ( .A1(n4894), .A2(n7500), .ZN(n5215) );
  AND2_X1 U4967 ( .A1(n8683), .A2(n8682), .ZN(n8684) );
  AOI21_X1 U4968 ( .B1(n8973), .B2(n5464), .A(n8244), .ZN(n8246) );
  AOI21_X1 U4969 ( .B1(n8978), .B2(n5464), .A(n8236), .ZN(n8731) );
  OAI21_X1 U4970 ( .B1(n4787), .B2(n4323), .A(n4452), .ZN(n8737) );
  INV_X1 U4971 ( .A(n4453), .ZN(n4452) );
  OAI21_X1 U4972 ( .B1(n4313), .B2(n4323), .A(n4457), .ZN(n4453) );
  OR2_X1 U4973 ( .A1(n8616), .A2(n8883), .ZN(n4457) );
  OR2_X1 U4974 ( .A1(n5218), .A2(n4864), .ZN(n5236) );
  INV_X1 U4975 ( .A(n5097), .ZN(n5326) );
  INV_X1 U4976 ( .A(n5749), .ZN(n5325) );
  OR2_X1 U4977 ( .A1(n5510), .A2(n5721), .ZN(n8861) );
  NAND2_X1 U4978 ( .A1(n5026), .A2(n5025), .ZN(n8898) );
  INV_X1 U4979 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4882) );
  INV_X1 U4980 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5021) );
  AND2_X1 U4981 ( .A1(n5472), .A2(n5324), .ZN(n7547) );
  OAI22_X1 U4982 ( .A1(n6292), .A2(n4447), .B1(n6293), .B2(n4448), .ZN(n6649)
         );
  AND2_X1 U4983 ( .A1(n6293), .A2(n4448), .ZN(n4447) );
  INV_X1 U4984 ( .A(n9059), .ZN(n4815) );
  NAND2_X1 U4985 ( .A1(n6649), .A2(n6648), .ZN(n4838) );
  OR2_X1 U4986 ( .A1(n8525), .A2(n8524), .ZN(n4813) );
  NAND2_X1 U4987 ( .A1(n4435), .A2(n4434), .ZN(n7529) );
  OR2_X1 U4988 ( .A1(n7490), .A2(n7518), .ZN(n4434) );
  NOR2_X1 U4989 ( .A1(n9190), .A2(n9392), .ZN(n8131) );
  AOI21_X1 U4990 ( .B1(n9203), .B2(n9205), .A(n4620), .ZN(n9189) );
  NOR2_X1 U4991 ( .A1(n9403), .A2(n9226), .ZN(n4620) );
  INV_X1 U4992 ( .A(n9227), .ZN(n9250) );
  AOI22_X1 U4993 ( .A1(n9279), .A2(n8127), .B1(n9026), .B2(n9284), .ZN(n9261)
         );
  NAND2_X1 U4994 ( .A1(n4358), .A2(n4610), .ZN(n4606) );
  AND2_X1 U4995 ( .A1(n9448), .A2(n9371), .ZN(n4611) );
  INV_X1 U4996 ( .A(n6120), .ZN(n7804) );
  NAND2_X1 U4997 ( .A1(n5929), .A2(n8092), .ZN(n5963) );
  NAND2_X1 U4998 ( .A1(n5394), .A2(n5393), .ZN(n5407) );
  NAND2_X1 U4999 ( .A1(n4592), .A2(n4994), .ZN(n5320) );
  NAND2_X1 U5000 ( .A1(n5035), .A2(n4992), .ZN(n4592) );
  BUF_X1 U5001 ( .A(n5024), .Z(n7725) );
  OR2_X1 U5002 ( .A1(n5721), .A2(n5508), .ZN(n8859) );
  AND2_X1 U5003 ( .A1(n5742), .A2(n5741), .ZN(n9686) );
  INV_X1 U5004 ( .A(n8097), .ZN(n9178) );
  AND2_X1 U5005 ( .A1(n8164), .A2(n8163), .ZN(n9394) );
  AOI22_X1 U5006 ( .A1(n9104), .A2(n9380), .B1(n8162), .B2(n9103), .ZN(n8163)
         );
  NAND2_X1 U5007 ( .A1(n8322), .A2(n8319), .ZN(n4467) );
  NAND2_X1 U5008 ( .A1(n7948), .A2(n4413), .ZN(n7958) );
  NOR2_X1 U5009 ( .A1(n4411), .A2(n8047), .ZN(n4410) );
  INV_X1 U5010 ( .A(n7964), .ZN(n4411) );
  NAND2_X1 U5011 ( .A1(n8049), .A2(n7968), .ZN(n4409) );
  AND2_X1 U5012 ( .A1(n4487), .A2(n8404), .ZN(n4486) );
  NAND2_X1 U5013 ( .A1(n4483), .A2(n4490), .ZN(n4487) );
  NAND2_X1 U5014 ( .A1(n8393), .A2(n8402), .ZN(n4483) );
  NAND2_X1 U5015 ( .A1(n4423), .A2(n4421), .ZN(n7983) );
  NAND2_X1 U5016 ( .A1(n4422), .A2(n8016), .ZN(n4421) );
  NAND2_X1 U5017 ( .A1(n4424), .A2(n8010), .ZN(n4423) );
  NAND2_X1 U5018 ( .A1(n7979), .A2(n7978), .ZN(n4422) );
  OAI21_X1 U5019 ( .B1(n8399), .B2(n8821), .A(n4349), .ZN(n4498) );
  INV_X1 U5020 ( .A(n8417), .ZN(n4496) );
  INV_X1 U5021 ( .A(n4946), .ZN(n4773) );
  INV_X1 U5022 ( .A(n4853), .ZN(n4655) );
  OAI21_X1 U5023 ( .B1(n4495), .B2(n4494), .A(n4492), .ZN(n4491) );
  NAND2_X1 U5024 ( .A1(n5439), .A2(n4365), .ZN(n4494) );
  NOR2_X1 U5025 ( .A1(n8744), .A2(n4493), .ZN(n4492) );
  AOI21_X1 U5026 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n4495) );
  NAND2_X1 U5027 ( .A1(n8285), .A2(n5517), .ZN(n8442) );
  OAI21_X1 U5028 ( .B1(n7711), .B2(n7710), .A(n7713), .ZN(n7722) );
  AND2_X1 U5029 ( .A1(n4594), .A2(n5384), .ZN(n4593) );
  AND2_X1 U5030 ( .A1(n5383), .A2(n5386), .ZN(n5384) );
  NAND2_X1 U5031 ( .A1(n4597), .A2(n4595), .ZN(n4594) );
  INV_X1 U5032 ( .A(n5345), .ZN(n4595) );
  INV_X1 U5033 ( .A(n4597), .ZN(n4596) );
  INV_X1 U5034 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5578) );
  NOR2_X1 U5035 ( .A1(n4769), .A2(n4773), .ZN(n4768) );
  INV_X1 U5036 ( .A(n4939), .ZN(n4769) );
  OAI21_X1 U5037 ( .B1(n4319), .B2(n4773), .A(n4856), .ZN(n4772) );
  NAND2_X1 U5038 ( .A1(n8179), .A2(n4388), .ZN(n4387) );
  INV_X1 U5039 ( .A(n8563), .ZN(n4388) );
  OR2_X1 U5040 ( .A1(n8577), .A2(n8576), .ZN(n4750) );
  NAND2_X1 U5041 ( .A1(n7380), .A2(n7377), .ZN(n7378) );
  NAND2_X1 U5042 ( .A1(n4328), .A2(n4727), .ZN(n4723) );
  OAI21_X1 U5043 ( .B1(n4654), .B2(n4649), .A(n4325), .ZN(n4648) );
  OAI21_X1 U5044 ( .B1(n4647), .B2(n4649), .A(n4646), .ZN(n4645) );
  AOI21_X1 U5045 ( .B1(n4650), .B2(n4652), .A(n4310), .ZN(n4646) );
  INV_X1 U5046 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U5047 ( .A1(n8781), .A2(n8761), .ZN(n4458) );
  OR2_X1 U5048 ( .A1(n8883), .A2(n8747), .ZN(n8428) );
  NAND2_X1 U5049 ( .A1(n4666), .A2(n5505), .ZN(n4660) );
  OR2_X1 U5050 ( .A1(n8807), .A2(n4661), .ZN(n4659) );
  NAND2_X1 U5051 ( .A1(n4666), .A2(n4662), .ZN(n4661) );
  AND2_X1 U5052 ( .A1(n8910), .A2(n8860), .ZN(n8411) );
  AND2_X1 U5053 ( .A1(n8842), .A2(n8621), .ZN(n8396) );
  NAND2_X1 U5054 ( .A1(n7623), .A2(n4672), .ZN(n4673) );
  NOR2_X1 U5055 ( .A1(n8855), .A2(n8395), .ZN(n4672) );
  NOR2_X1 U5056 ( .A1(n7618), .A2(n8858), .ZN(n4775) );
  OR2_X1 U5057 ( .A1(n5318), .A2(n7565), .ZN(n8289) );
  OR2_X1 U5058 ( .A1(n7501), .A2(n4369), .ZN(n4459) );
  NOR2_X1 U5059 ( .A1(n8947), .A2(n8941), .ZN(n4552) );
  NOR2_X1 U5060 ( .A1(n8376), .A2(n4668), .ZN(n4667) );
  INV_X1 U5061 ( .A(n8378), .ZN(n4668) );
  AND2_X1 U5062 ( .A1(n7175), .A2(n9527), .ZN(n7174) );
  NAND2_X1 U5063 ( .A1(n6543), .A2(n4339), .ZN(n4642) );
  INV_X1 U5064 ( .A(n5486), .ZN(n8298) );
  NAND2_X1 U5065 ( .A1(n8282), .A2(n8303), .ZN(n6216) );
  AOI21_X1 U5066 ( .B1(n9753), .B2(n9759), .A(n9761), .ZN(n6206) );
  INV_X1 U5067 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5038) );
  INV_X1 U5068 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5037) );
  INV_X1 U5069 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4674) );
  AND2_X1 U5070 ( .A1(n5037), .A2(n5038), .ZN(n4759) );
  INV_X1 U5071 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5477) );
  INV_X1 U5072 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5476) );
  INV_X2 U5073 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U5074 ( .A1(n4817), .A2(n4816), .ZN(n8476) );
  AOI21_X1 U5075 ( .B1(n4818), .B2(n4821), .A(n4318), .ZN(n4816) );
  INV_X1 U5076 ( .A(n8094), .ZN(n4427) );
  OR2_X1 U5077 ( .A1(n8011), .A2(n8016), .ZN(n4430) );
  OR2_X1 U5078 ( .A1(n8012), .A2(n8010), .ZN(n4429) );
  INV_X1 U5079 ( .A(n6132), .ZN(n5932) );
  OR2_X1 U5080 ( .A1(n9403), .A2(n9096), .ZN(n8155) );
  INV_X1 U5081 ( .A(n4618), .ZN(n4616) );
  NAND2_X1 U5082 ( .A1(n9406), .A2(n9240), .ZN(n4621) );
  AND2_X1 U5083 ( .A1(n9426), .A2(n9026), .ZN(n8145) );
  OR2_X1 U5084 ( .A1(n9426), .A2(n9026), .ZN(n8144) );
  OR2_X1 U5085 ( .A1(n9432), .A2(n9049), .ZN(n8024) );
  NOR2_X1 U5086 ( .A1(n9316), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U5087 ( .A1(n9337), .A2(n9082), .ZN(n4610) );
  OR2_X1 U5088 ( .A1(n9436), .A2(n9328), .ZN(n8141) );
  NAND2_X1 U5089 ( .A1(n8047), .A2(n7966), .ZN(n4709) );
  INV_X1 U5090 ( .A(n8137), .ZN(n4705) );
  OR2_X1 U5091 ( .A1(n9375), .A2(n9376), .ZN(n9347) );
  OR2_X1 U5092 ( .A1(n9459), .A2(n7610), .ZN(n8135) );
  OR2_X1 U5093 ( .A1(n7832), .A2(n7831), .ZN(n7960) );
  NAND2_X1 U5094 ( .A1(n6319), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7242) );
  NAND2_X1 U5095 ( .A1(n7141), .A2(n8042), .ZN(n4693) );
  NOR2_X1 U5096 ( .A1(n4692), .A2(n8045), .ZN(n4691) );
  INV_X1 U5097 ( .A(n7954), .ZN(n4692) );
  OR2_X1 U5098 ( .A1(n6928), .A2(n6927), .ZN(n7029) );
  NOR2_X1 U5099 ( .A1(n6423), .A2(n6488), .ZN(n6499) );
  NAND2_X1 U5100 ( .A1(n4703), .A2(n4701), .ZN(n6458) );
  NOR2_X1 U5101 ( .A1(n8065), .A2(n4702), .ZN(n4701) );
  INV_X1 U5102 ( .A(n6409), .ZN(n4702) );
  NAND2_X1 U5103 ( .A1(n6408), .A2(n8033), .ZN(n4703) );
  XNOR2_X1 U5104 ( .A(n7722), .B(n7721), .ZN(n7719) );
  NOR2_X1 U5105 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5692) );
  NAND2_X1 U5106 ( .A1(n4575), .A2(n5409), .ZN(n5426) );
  NOR2_X1 U5107 ( .A1(n5408), .A2(n4577), .ZN(n4576) );
  INV_X1 U5108 ( .A(n5393), .ZN(n4577) );
  NAND2_X1 U5109 ( .A1(n4599), .A2(n5008), .ZN(n5367) );
  NAND2_X1 U5110 ( .A1(n5581), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5585) );
  AOI21_X1 U5111 ( .B1(n5034), .B2(n4590), .A(n4588), .ZN(n4587) );
  INV_X1 U5112 ( .A(n4590), .ZN(n4589) );
  INV_X1 U5113 ( .A(n4999), .ZN(n4588) );
  AND2_X1 U5114 ( .A1(n5004), .A2(n5003), .ZN(n5336) );
  OAI21_X1 U5115 ( .B1(n4586), .B2(n4582), .A(n4579), .ZN(n5302) );
  NAND2_X1 U5116 ( .A1(n4584), .A2(n4583), .ZN(n4582) );
  AOI21_X1 U5117 ( .B1(n4584), .B2(n4581), .A(n4580), .ZN(n4579) );
  INV_X1 U5118 ( .A(n5285), .ZN(n4583) );
  AND2_X1 U5119 ( .A1(n4985), .A2(n4984), .ZN(n5301) );
  AND2_X1 U5120 ( .A1(n5577), .A2(n5815), .ZN(n4842) );
  INV_X1 U5121 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5560) );
  AOI21_X1 U5122 ( .B1(n5145), .B2(n4763), .A(n4355), .ZN(n4762) );
  INV_X1 U5123 ( .A(n4931), .ZN(n4763) );
  OAI21_X1 U5124 ( .B1(n5942), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4920), .ZN(
        n4921) );
  NAND2_X1 U5125 ( .A1(n4641), .A2(n5657), .ZN(n4640) );
  NAND2_X1 U5126 ( .A1(n5897), .A2(n4906), .ZN(n4908) );
  NOR2_X1 U5127 ( .A1(n8209), .A2(n4748), .ZN(n4747) );
  AND2_X1 U5128 ( .A1(n8577), .A2(n8576), .ZN(n4748) );
  AND2_X1 U5129 ( .A1(n4750), .A2(n8186), .ZN(n4744) );
  AND2_X1 U5130 ( .A1(n4738), .A2(n4732), .ZN(n4731) );
  NAND2_X1 U5131 ( .A1(n8567), .A2(n4733), .ZN(n4732) );
  NAND2_X1 U5132 ( .A1(n8177), .A2(n8603), .ZN(n4391) );
  INV_X1 U5133 ( .A(n4399), .ZN(n4398) );
  OAI21_X1 U5134 ( .B1(n4401), .B2(n4400), .A(n7572), .ZN(n4399) );
  INV_X1 U5135 ( .A(n4404), .ZN(n4400) );
  NAND2_X1 U5136 ( .A1(n7474), .A2(n7475), .ZN(n4404) );
  OR2_X1 U5137 ( .A1(n8577), .A2(n8576), .ZN(n4742) );
  NOR2_X1 U5138 ( .A1(n4756), .A2(n4368), .ZN(n4755) );
  INV_X1 U5139 ( .A(n7387), .ZN(n4756) );
  OR2_X1 U5140 ( .A1(n5279), .A2(n5278), .ZN(n5293) );
  NOR2_X1 U5141 ( .A1(n5804), .A2(n4560), .ZN(n5758) );
  AND2_X1 U5142 ( .A1(n5761), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4560) );
  OR2_X1 U5143 ( .A1(n5758), .A2(n5757), .ZN(n4559) );
  OR2_X1 U5144 ( .A1(n6187), .A2(n6186), .ZN(n4557) );
  AND2_X1 U5145 ( .A1(n4557), .A2(n4556), .ZN(n6378) );
  NAND2_X1 U5146 ( .A1(n6375), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4556) );
  OR2_X1 U5147 ( .A1(n6378), .A2(n6377), .ZN(n4555) );
  NOR2_X1 U5148 ( .A1(n6962), .A2(n4563), .ZN(n6964) );
  AND2_X1 U5149 ( .A1(n6963), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4563) );
  NAND2_X1 U5150 ( .A1(n7410), .A2(n4561), .ZN(n8648) );
  INV_X1 U5151 ( .A(n7412), .ZN(n4561) );
  AND2_X1 U5152 ( .A1(n8698), .A2(n8701), .ZN(n4569) );
  NAND2_X1 U5153 ( .A1(n8684), .A2(n8685), .ZN(n8699) );
  INV_X1 U5154 ( .A(n8699), .ZN(n4568) );
  OAI21_X1 U5155 ( .B1(n8684), .B2(n4566), .A(n4564), .ZN(n8709) );
  INV_X1 U5156 ( .A(n4569), .ZN(n4566) );
  AOI21_X1 U5157 ( .B1(n4565), .B2(n4569), .A(n4373), .ZN(n4564) );
  NAND2_X1 U5158 ( .A1(n4545), .A2(n8731), .ZN(n4544) );
  INV_X1 U5159 ( .A(n4545), .ZN(n4543) );
  NOR2_X1 U5160 ( .A1(n4327), .A2(n4853), .ZN(n8235) );
  AND2_X1 U5161 ( .A1(n4377), .A2(n4376), .ZN(n8758) );
  NOR2_X1 U5162 ( .A1(n8759), .A2(n8760), .ZN(n4376) );
  AND2_X1 U5163 ( .A1(n5453), .A2(n5452), .ZN(n8762) );
  NAND2_X1 U5164 ( .A1(n4665), .A2(n4458), .ZN(n4456) );
  INV_X1 U5165 ( .A(n4786), .ZN(n4785) );
  OAI22_X1 U5166 ( .A1(n4666), .A2(n4792), .B1(n8894), .B2(n8618), .ZN(n4786)
         );
  NOR2_X1 U5167 ( .A1(n4666), .A2(n4789), .ZN(n4788) );
  INV_X1 U5168 ( .A(n4790), .ZN(n4789) );
  NAND2_X1 U5169 ( .A1(n8805), .A2(n8586), .ZN(n4792) );
  OR2_X1 U5170 ( .A1(n8807), .A2(n8808), .ZN(n4663) );
  NAND2_X1 U5171 ( .A1(n8903), .A2(n4790), .ZN(n4793) );
  NAND2_X1 U5172 ( .A1(n8862), .A2(n8842), .ZN(n8836) );
  INV_X1 U5173 ( .A(n5330), .ZN(n4869) );
  INV_X1 U5174 ( .A(n8621), .ZN(n8860) );
  AOI21_X1 U5175 ( .B1(n7542), .B2(n8273), .A(n5504), .ZN(n7619) );
  NAND2_X1 U5176 ( .A1(n7619), .A2(n7620), .ZN(n7623) );
  NAND2_X1 U5177 ( .A1(n4780), .A2(n4783), .ZN(n4779) );
  INV_X1 U5178 ( .A(n8272), .ZN(n4780) );
  NAND2_X1 U5179 ( .A1(n4781), .A2(n4783), .ZN(n4778) );
  NAND2_X1 U5180 ( .A1(n5335), .A2(n4782), .ZN(n4781) );
  INV_X1 U5181 ( .A(n4784), .ZN(n4782) );
  INV_X1 U5182 ( .A(n4459), .ZN(n7556) );
  OR2_X1 U5183 ( .A1(n7329), .A2(n7509), .ZN(n4850) );
  NAND2_X1 U5184 ( .A1(n4866), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5310) );
  INV_X1 U5185 ( .A(n5293), .ZN(n4866) );
  NAND2_X1 U5186 ( .A1(n4867), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5312) );
  INV_X1 U5187 ( .A(n5310), .ZN(n4867) );
  OR2_X1 U5188 ( .A1(n7214), .A2(n7261), .ZN(n8378) );
  OR2_X1 U5189 ( .A1(n5255), .A2(n7227), .ZN(n5279) );
  NOR2_X2 U5190 ( .A1(n7116), .A2(n8952), .ZN(n7175) );
  AND2_X1 U5191 ( .A1(n5493), .A2(n4332), .ZN(n4669) );
  AND2_X1 U5192 ( .A1(n8359), .A2(n8362), .ZN(n8266) );
  NAND2_X1 U5193 ( .A1(n4332), .A2(n8338), .ZN(n8264) );
  NAND2_X1 U5194 ( .A1(n4379), .A2(n4671), .ZN(n4670) );
  INV_X1 U5195 ( .A(n6821), .ZN(n4379) );
  AND4_X1 U5196 ( .A1(n5223), .A2(n5222), .A3(n5221), .A4(n5220), .ZN(n7656)
         );
  AND2_X1 U5197 ( .A1(n6560), .A2(n5180), .ZN(n6818) );
  NOR2_X1 U5198 ( .A1(n6975), .A2(n9802), .ZN(n4548) );
  OR2_X1 U5199 ( .A1(n5174), .A2(n5173), .ZN(n5187) );
  AND2_X1 U5200 ( .A1(n8344), .A2(n8331), .ZN(n8259) );
  INV_X1 U5201 ( .A(n6357), .ZN(n5128) );
  NAND2_X1 U5202 ( .A1(n6441), .A2(n6443), .ZN(n5085) );
  INV_X1 U5203 ( .A(n8859), .ZN(n7566) );
  INV_X1 U5204 ( .A(n8817), .ZN(n8857) );
  NAND2_X1 U5205 ( .A1(n5466), .A2(n5465), .ZN(n7700) );
  AND2_X1 U5206 ( .A1(n5144), .A2(n5143), .ZN(n9794) );
  INV_X1 U5207 ( .A(n9786), .ZN(n9810) );
  INV_X1 U5208 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U5209 ( .A1(n5521), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5548) );
  XNOR2_X1 U5210 ( .A(n5548), .B(P2_IR_REG_23__SCAN_IN), .ZN(n5722) );
  OAI21_X1 U5211 ( .B1(n5480), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5520) );
  NOR2_X1 U5212 ( .A1(n4801), .A2(n4445), .ZN(n4444) );
  NAND2_X1 U5213 ( .A1(n6655), .A2(n6654), .ZN(n6657) );
  NAND2_X1 U5214 ( .A1(n7090), .A2(n7089), .ZN(n4439) );
  XNOR2_X1 U5215 ( .A(n6081), .B(n6095), .ZN(n6263) );
  AND2_X1 U5216 ( .A1(n7603), .A2(n4819), .ZN(n4818) );
  NAND2_X1 U5217 ( .A1(n7600), .A2(n4820), .ZN(n4819) );
  INV_X1 U5218 ( .A(n7530), .ZN(n4820) );
  NAND2_X1 U5219 ( .A1(n7529), .A2(n7530), .ZN(n7601) );
  OR2_X1 U5220 ( .A1(n7820), .A2(n8986), .ZN(n7865) );
  INV_X1 U5221 ( .A(n8519), .ZN(n4810) );
  INV_X1 U5222 ( .A(n7809), .ZN(n6323) );
  NAND2_X1 U5223 ( .A1(n4824), .A2(n4829), .ZN(n8513) );
  AND2_X1 U5224 ( .A1(n4804), .A2(n4802), .ZN(n4801) );
  NAND2_X1 U5225 ( .A1(n4803), .A2(n4364), .ZN(n4802) );
  NAND2_X1 U5226 ( .A1(n4805), .A2(n9040), .ZN(n4804) );
  INV_X1 U5227 ( .A(n9032), .ZN(n4803) );
  NOR2_X1 U5228 ( .A1(n4806), .A2(n4797), .ZN(n4796) );
  INV_X1 U5229 ( .A(n4811), .ZN(n4797) );
  NAND2_X1 U5230 ( .A1(n8109), .A2(n5900), .ZN(n8061) );
  INV_X1 U5231 ( .A(n7490), .ZN(n4437) );
  NAND2_X1 U5232 ( .A1(n7485), .A2(n7484), .ZN(n4438) );
  NAND2_X1 U5233 ( .A1(n7427), .A2(n7426), .ZN(n7486) );
  OAI21_X1 U5234 ( .B1(n7868), .B2(n4681), .A(n4679), .ZN(n4678) );
  AND2_X1 U5235 ( .A1(n5706), .A2(n7639), .ZN(n6114) );
  NAND2_X1 U5236 ( .A1(n5862), .A2(n5863), .ZN(n9599) );
  AND2_X1 U5237 ( .A1(n4521), .A2(n4520), .ZN(n9598) );
  NAND2_X1 U5238 ( .A1(n6056), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U5239 ( .A1(n9602), .A2(n5864), .ZN(n4520) );
  NAND2_X1 U5240 ( .A1(n9662), .A2(n9661), .ZN(n9660) );
  NAND2_X1 U5241 ( .A1(n4525), .A2(n4524), .ZN(n4523) );
  INV_X1 U5242 ( .A(n9138), .ZN(n4524) );
  NAND2_X1 U5243 ( .A1(n7731), .A2(n7730), .ZN(n8114) );
  INV_X1 U5244 ( .A(n9240), .ZN(n9209) );
  NOR2_X1 U5245 ( .A1(n4687), .A2(n9218), .ZN(n4685) );
  INV_X1 U5246 ( .A(n8151), .ZN(n4683) );
  INV_X1 U5247 ( .A(n4685), .ZN(n4684) );
  NAND2_X1 U5248 ( .A1(n8155), .A2(n8022), .ZN(n9205) );
  NAND2_X1 U5249 ( .A1(n4686), .A2(n4685), .ZN(n9225) );
  AND2_X1 U5250 ( .A1(n4622), .A2(n8129), .ZN(n4618) );
  NAND2_X1 U5251 ( .A1(n8130), .A2(n8129), .ZN(n4619) );
  NOR2_X1 U5252 ( .A1(n9309), .A2(n9432), .ZN(n9293) );
  NAND2_X1 U5253 ( .A1(n4601), .A2(n4600), .ZN(n9292) );
  AOI21_X1 U5254 ( .B1(n4603), .B2(n4605), .A(n4348), .ZN(n4600) );
  NAND2_X1 U5255 ( .A1(n9326), .A2(n9324), .ZN(n4700) );
  AND2_X1 U5256 ( .A1(n4610), .A2(n9348), .ZN(n4607) );
  NAND2_X1 U5257 ( .A1(n6321), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7808) );
  INV_X1 U5258 ( .A(n7459), .ZN(n6321) );
  OR2_X1 U5259 ( .A1(n7469), .A2(n9459), .ZN(n9363) );
  INV_X1 U5260 ( .A(n9353), .ZN(n8124) );
  OAI21_X1 U5261 ( .B1(n7342), .B2(n8046), .A(n7960), .ZN(n7465) );
  OR2_X1 U5262 ( .A1(n8061), .A2(n5736), .ZN(n9331) );
  INV_X1 U5263 ( .A(n9355), .ZN(n9374) );
  INV_X1 U5264 ( .A(n9329), .ZN(n9372) );
  INV_X1 U5265 ( .A(n9331), .ZN(n9380) );
  NAND2_X1 U5266 ( .A1(n7900), .A2(n7899), .ZN(n9392) );
  OR2_X1 U5267 ( .A1(n5963), .A2(n5960), .ZN(n9710) );
  OR3_X1 U5268 ( .A1(n7400), .A2(n7272), .A3(n7079), .ZN(n6132) );
  XNOR2_X1 U5269 ( .A(n5575), .B(n5574), .ZN(n6130) );
  XNOR2_X1 U5270 ( .A(n7719), .B(SI_30_), .ZN(n8978) );
  NAND2_X1 U5271 ( .A1(n5693), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5590) );
  INV_X1 U5272 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5570) );
  NOR2_X1 U5273 ( .A1(n5366), .A2(n4598), .ZN(n4597) );
  INV_X1 U5274 ( .A(n5008), .ZN(n4598) );
  OR2_X1 U5275 ( .A1(n6246), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U5276 ( .A1(n4578), .A2(n4584), .ZN(n5286) );
  NAND2_X1 U5277 ( .A1(n4586), .A2(n4308), .ZN(n4578) );
  AOI21_X1 U5278 ( .B1(n5268), .B2(n5267), .A(n5266), .ZN(n5270) );
  XNOR2_X1 U5279 ( .A(n5249), .B(n5248), .ZN(n7138) );
  OR2_X1 U5280 ( .A1(n5683), .A2(n9486), .ZN(n5686) );
  NAND2_X1 U5281 ( .A1(n4928), .A2(n4927), .ZN(n5137) );
  NAND2_X1 U5282 ( .A1(n4735), .A2(n8170), .ZN(n8568) );
  NAND2_X1 U5283 ( .A1(n7629), .A2(n4736), .ZN(n4735) );
  NAND2_X1 U5284 ( .A1(n5348), .A2(n5347), .ZN(n8916) );
  NAND2_X1 U5285 ( .A1(n5235), .A2(n5234), .ZN(n7128) );
  AND2_X1 U5286 ( .A1(n8184), .A2(n8183), .ZN(n8575) );
  AND4_X1 U5287 ( .A1(n5136), .A2(n5135), .A3(n5134), .A4(n5133), .ZN(n8218)
         );
  NAND2_X1 U5288 ( .A1(n6734), .A2(n6733), .ZN(n6736) );
  AND3_X1 U5289 ( .A1(n5354), .A2(n5353), .A3(n5352), .ZN(n8844) );
  INV_X1 U5290 ( .A(n8842), .ZN(n8910) );
  AND4_X1 U5291 ( .A1(n5206), .A2(n5205), .A3(n5204), .A4(n5203), .ZN(n6819)
         );
  AND4_X1 U5292 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n7108)
         );
  NAND2_X1 U5293 ( .A1(n5213), .A2(n5212), .ZN(n7007) );
  NAND2_X1 U5294 ( .A1(n4469), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U5295 ( .A1(n6635), .A2(n5617), .ZN(n4392) );
  NAND2_X1 U5296 ( .A1(n8452), .A2(n8451), .ZN(n4470) );
  NAND2_X1 U5297 ( .A1(n4475), .A2(n4472), .ZN(n4471) );
  INV_X1 U5298 ( .A(n8449), .ZN(n4472) );
  OR2_X1 U5299 ( .A1(n4475), .A2(n4474), .ZN(n4473) );
  NAND2_X1 U5300 ( .A1(n4717), .A2(n5595), .ZN(n4474) );
  NAND2_X1 U5301 ( .A1(n5637), .A2(n9760), .ZN(n9754) );
  INV_X1 U5302 ( .A(n8762), .ZN(n8615) );
  AND2_X1 U5303 ( .A1(n7077), .A2(n7365), .ZN(n9757) );
  NOR2_X1 U5304 ( .A1(n5722), .A2(P2_U3152), .ZN(n9760) );
  INV_X1 U5305 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8974) );
  XNOR2_X1 U5306 ( .A(n5023), .B(n5022), .ZN(n5508) );
  INV_X1 U5307 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U5308 ( .A1(n4541), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5023) );
  NAND2_X1 U5309 ( .A1(n5534), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4381) );
  INV_X1 U5310 ( .A(n7547), .ZN(n9744) );
  NAND2_X1 U5311 ( .A1(n7819), .A2(n7818), .ZN(n9421) );
  NAND2_X1 U5312 ( .A1(n7806), .A2(n7805), .ZN(n9444) );
  NAND2_X1 U5313 ( .A1(n9089), .A2(n4843), .ZN(n9011) );
  AND2_X1 U5314 ( .A1(n9001), .A2(n8537), .ZN(n4843) );
  OR2_X1 U5315 ( .A1(n9015), .A2(n9086), .ZN(n4844) );
  NAND2_X1 U5316 ( .A1(n7884), .A2(n7883), .ZN(n9396) );
  NAND2_X1 U5317 ( .A1(n9046), .A2(n9047), .ZN(n9022) );
  NAND2_X1 U5318 ( .A1(n7759), .A2(n7758), .ZN(n9411) );
  NAND2_X1 U5319 ( .A1(n7864), .A2(n7863), .ZN(n9418) );
  INV_X1 U5320 ( .A(n9099), .ZN(n9050) );
  NAND2_X1 U5321 ( .A1(n7801), .A2(n7800), .ZN(n9448) );
  NAND2_X1 U5322 ( .A1(n9091), .A2(n9090), .ZN(n9089) );
  INV_X1 U5323 ( .A(n9086), .ZN(n9088) );
  NAND2_X1 U5324 ( .A1(n7767), .A2(n7766), .ZN(n9227) );
  NAND2_X1 U5325 ( .A1(n7875), .A2(n7874), .ZN(n9273) );
  OAI21_X1 U5326 ( .B1(n9176), .B2(n9623), .A(n4534), .ZN(n4533) );
  AOI21_X1 U5327 ( .B1(n9177), .B2(n9686), .A(n9678), .ZN(n4534) );
  NAND2_X1 U5328 ( .A1(n9367), .A2(n6277), .ZN(n9364) );
  INV_X1 U5329 ( .A(n4624), .ZN(n4623) );
  OAI21_X1 U5330 ( .B1(n9394), .B2(n9717), .A(n4372), .ZN(n4624) );
  INV_X1 U5331 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4631) );
  AOI21_X1 U5332 ( .B1(n9465), .B2(n9392), .A(n9391), .ZN(n9393) );
  NAND2_X1 U5333 ( .A1(n8159), .A2(n4363), .ZN(n4629) );
  NOR2_X1 U5334 ( .A1(n8159), .A2(n4363), .ZN(n4628) );
  XNOR2_X1 U5335 ( .A(n5889), .B(n5888), .ZN(n8097) );
  INV_X1 U5336 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5888) );
  INV_X1 U5337 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4903) );
  OAI21_X1 U5338 ( .B1(n4466), .B2(n4331), .A(n8330), .ZN(n8350) );
  AOI21_X1 U5339 ( .B1(n8311), .B2(n8310), .A(n4467), .ZN(n4466) );
  NOR2_X1 U5340 ( .A1(n7942), .A2(n7935), .ZN(n4418) );
  NAND2_X1 U5341 ( .A1(n7934), .A2(n7933), .ZN(n4417) );
  AOI21_X1 U5342 ( .B1(n4415), .B2(n8016), .A(n4414), .ZN(n4413) );
  OAI211_X1 U5343 ( .C1(n8016), .C2(n7938), .A(n7949), .B(n8040), .ZN(n4414)
         );
  NAND2_X1 U5344 ( .A1(n4416), .A2(n7937), .ZN(n4415) );
  OAI21_X1 U5345 ( .B1(n4418), .B2(n4417), .A(n4715), .ZN(n4416) );
  AOI21_X1 U5346 ( .B1(n8365), .B2(n8361), .A(n8360), .ZN(n8367) );
  OAI21_X1 U5347 ( .B1(n4408), .B2(n4407), .A(n7975), .ZN(n7980) );
  NAND2_X1 U5348 ( .A1(n9360), .A2(n7969), .ZN(n4407) );
  AOI21_X1 U5349 ( .B1(n7965), .B2(n4410), .A(n4409), .ZN(n4408) );
  AND2_X1 U5350 ( .A1(n4482), .A2(n4362), .ZN(n4481) );
  OR2_X1 U5351 ( .A1(n4486), .A2(n8395), .ZN(n4482) );
  INV_X1 U5352 ( .A(n4485), .ZN(n4484) );
  AOI21_X1 U5353 ( .B1(n4486), .B2(n4488), .A(n8395), .ZN(n4485) );
  NAND2_X1 U5354 ( .A1(n4419), .A2(n8143), .ZN(n7982) );
  NAND2_X1 U5355 ( .A1(n7983), .A2(n4420), .ZN(n4419) );
  AND2_X1 U5356 ( .A1(n8024), .A2(n8141), .ZN(n4420) );
  AND2_X1 U5357 ( .A1(n4497), .A2(n4496), .ZN(n8422) );
  INV_X1 U5358 ( .A(n8430), .ZN(n4493) );
  INV_X1 U5359 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n4878) );
  INV_X1 U5360 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4877) );
  NOR2_X1 U5361 ( .A1(n5319), .A2(n4591), .ZN(n4590) );
  INV_X1 U5362 ( .A(n4994), .ZN(n4591) );
  INV_X1 U5363 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4987) );
  NOR2_X1 U5364 ( .A1(n4308), .A2(n5285), .ZN(n4581) );
  INV_X1 U5365 ( .A(n4980), .ZN(n4580) );
  INV_X1 U5366 ( .A(n8170), .ZN(n4733) );
  NOR2_X1 U5367 ( .A1(n4734), .A2(n4730), .ZN(n4729) );
  INV_X1 U5368 ( .A(n4736), .ZN(n4730) );
  INV_X1 U5369 ( .A(n8567), .ZN(n4734) );
  INV_X1 U5370 ( .A(n4739), .ZN(n4738) );
  OAI21_X1 U5371 ( .B1(n8177), .B2(n8603), .A(n8597), .ZN(n4739) );
  INV_X1 U5372 ( .A(n5617), .ZN(n4395) );
  NAND2_X1 U5373 ( .A1(n8246), .A2(n8727), .ZN(n8441) );
  NAND2_X1 U5374 ( .A1(n4491), .A2(n4338), .ZN(n8438) );
  NAND2_X1 U5375 ( .A1(n4574), .A2(n4573), .ZN(n8447) );
  NAND2_X1 U5376 ( .A1(n8287), .A2(n8435), .ZN(n4573) );
  NAND2_X1 U5377 ( .A1(n8286), .A2(n8442), .ZN(n4574) );
  NAND2_X1 U5378 ( .A1(n8648), .A2(n8647), .ZN(n8655) );
  INV_X1 U5379 ( .A(n8685), .ZN(n4565) );
  NOR2_X1 U5380 ( .A1(n4546), .A2(n7700), .ZN(n4545) );
  NAND2_X1 U5381 ( .A1(n8743), .A2(n4547), .ZN(n4546) );
  INV_X1 U5382 ( .A(n4456), .ZN(n4454) );
  OR2_X1 U5383 ( .A1(n5501), .A2(n8385), .ZN(n7505) );
  NAND2_X1 U5384 ( .A1(n7319), .A2(n5499), .ZN(n7506) );
  NOR2_X1 U5385 ( .A1(n7663), .A2(n5207), .ZN(n6898) );
  NAND2_X1 U5386 ( .A1(n5207), .A2(n6819), .ZN(n8294) );
  AND2_X1 U5387 ( .A1(n8343), .A2(n8353), .ZN(n7651) );
  NAND2_X1 U5388 ( .A1(n9780), .A2(n8639), .ZN(n8320) );
  NAND2_X1 U5389 ( .A1(n4374), .A2(n7676), .ZN(n8315) );
  NAND2_X1 U5390 ( .A1(n7263), .A2(n4342), .ZN(n7324) );
  NAND2_X1 U5391 ( .A1(n8368), .A2(n7169), .ZN(n8374) );
  INV_X1 U5392 ( .A(n4765), .ZN(n7109) );
  OAI21_X1 U5393 ( .B1(n8266), .B2(n6990), .A(n5262), .ZN(n4765) );
  NOR2_X1 U5394 ( .A1(n9778), .A2(n8303), .ZN(n5633) );
  INV_X1 U5395 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U5396 ( .A1(n5036), .A2(n4759), .ZN(n5474) );
  AND2_X1 U5397 ( .A1(n5036), .A2(n5037), .ZN(n5304) );
  INV_X1 U5398 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5273) );
  OR2_X1 U5399 ( .A1(n5168), .A2(n5167), .ZN(n5182) );
  INV_X1 U5400 ( .A(n7518), .ZN(n4436) );
  AND2_X1 U5401 ( .A1(n8501), .A2(n4830), .ZN(n4829) );
  NAND2_X1 U5402 ( .A1(n9047), .A2(n4833), .ZN(n4830) );
  INV_X1 U5403 ( .A(n4806), .ZN(n4805) );
  NAND2_X1 U5404 ( .A1(n4364), .A2(n4813), .ZN(n4806) );
  NOR2_X1 U5405 ( .A1(n7422), .A2(n4823), .ZN(n4822) );
  INV_X1 U5406 ( .A(n7181), .ZN(n4823) );
  NOR2_X1 U5407 ( .A1(n7306), .A2(n4535), .ZN(n7307) );
  NOR2_X1 U5408 ( .A1(n4537), .A2(n4536), .ZN(n4535) );
  INV_X1 U5409 ( .A(n7313), .ZN(n4537) );
  NAND2_X1 U5410 ( .A1(n4511), .A2(n9215), .ZN(n4510) );
  NOR2_X1 U5411 ( .A1(n9406), .A2(n9411), .ZN(n4511) );
  NAND2_X1 U5412 ( .A1(n6324), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7820) );
  INV_X1 U5413 ( .A(n7785), .ZN(n6324) );
  OR2_X1 U5414 ( .A1(n9421), .A2(n9249), .ZN(n8147) );
  INV_X1 U5415 ( .A(n4606), .ZN(n4605) );
  NAND2_X1 U5416 ( .A1(n4515), .A2(n9337), .ZN(n4514) );
  INV_X1 U5417 ( .A(n4516), .ZN(n4515) );
  NAND2_X1 U5418 ( .A1(n9346), .A2(n4517), .ZN(n4516) );
  NOR2_X1 U5419 ( .A1(n9464), .A2(n7835), .ZN(n4505) );
  NOR2_X1 U5420 ( .A1(n7236), .A2(n4504), .ZN(n4503) );
  INV_X1 U5421 ( .A(n4505), .ZN(n4504) );
  INV_X1 U5422 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7028) );
  OR2_X1 U5423 ( .A1(n7029), .A2(n7028), .ZN(n7149) );
  INV_X1 U5424 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6927) );
  INV_X1 U5425 ( .A(n6851), .ZN(n6318) );
  NOR2_X1 U5426 ( .A1(n7941), .A2(n4714), .ZN(n4713) );
  INV_X1 U5427 ( .A(n7926), .ZN(n4714) );
  INV_X1 U5428 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6716) );
  OR2_X1 U5429 ( .A1(n6717), .A2(n6716), .ZN(n6851) );
  NAND2_X1 U5430 ( .A1(n6317), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6717) );
  INV_X1 U5431 ( .A(n6662), .ZN(n6317) );
  INV_X1 U5432 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6305) );
  OR2_X1 U5433 ( .A1(n6306), .A2(n6305), .ZN(n6662) );
  AND2_X1 U5434 ( .A1(n6677), .A2(n6605), .ZN(n4519) );
  OR2_X1 U5435 ( .A1(n9396), .A2(n9208), .ZN(n8158) );
  NAND2_X1 U5436 ( .A1(n5998), .A2(n5997), .ZN(n6408) );
  OAI21_X1 U5437 ( .B1(n5572), .B2(n9486), .A(n4845), .ZN(n5593) );
  INV_X1 U5438 ( .A(n4846), .ZN(n4845) );
  OAI21_X1 U5439 ( .B1(n4847), .B2(n9486), .A(n5589), .ZN(n4846) );
  AND2_X1 U5440 ( .A1(n5442), .A2(n5432), .ZN(n5440) );
  AND2_X1 U5441 ( .A1(n5427), .A2(n5413), .ZN(n5425) );
  AND2_X1 U5442 ( .A1(n5390), .A2(n5389), .ZN(n5394) );
  NAND2_X1 U5443 ( .A1(n4986), .A2(n4985), .ZN(n5046) );
  OR2_X1 U5444 ( .A1(n5245), .A2(n5244), .ZN(n5268) );
  INV_X1 U5445 ( .A(n4772), .ZN(n4771) );
  AND2_X1 U5446 ( .A1(n5674), .A2(n5556), .ZN(n5682) );
  INV_X1 U5447 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5556) );
  INV_X1 U5448 ( .A(n5024), .ZN(n4919) );
  NAND2_X1 U5449 ( .A1(n4412), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4760) );
  NAND2_X1 U5450 ( .A1(n4904), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4412) );
  OR2_X1 U5451 ( .A1(n5312), .A2(n4868), .ZN(n5330) );
  NAND2_X1 U5452 ( .A1(n4718), .A2(n4717), .ZN(n4716) );
  NOR2_X1 U5453 ( .A1(n9763), .A2(n8303), .ZN(n4718) );
  NOR2_X1 U5454 ( .A1(n8171), .A2(n4737), .ZN(n4736) );
  INV_X1 U5455 ( .A(n7628), .ZN(n4737) );
  OR2_X1 U5456 ( .A1(n5375), .A2(n5374), .ZN(n5377) );
  INV_X1 U5457 ( .A(n4386), .ZN(n4385) );
  OAI21_X1 U5458 ( .B1(n4330), .B2(n4391), .A(n4387), .ZN(n4386) );
  AND2_X1 U5459 ( .A1(n6757), .A2(n6752), .ZN(n4751) );
  NAND2_X1 U5460 ( .A1(n6391), .A2(n8250), .ZN(n5598) );
  NOR2_X1 U5461 ( .A1(n7476), .A2(n4402), .ZN(n4401) );
  INV_X1 U5462 ( .A(n7392), .ZN(n4402) );
  AND2_X1 U5463 ( .A1(n7378), .A2(n4723), .ZN(n4722) );
  OR2_X1 U5464 ( .A1(n5641), .A2(n9754), .ZN(n5632) );
  AOI21_X1 U5465 ( .B1(n8745), .B2(n4653), .A(n4648), .ZN(n8241) );
  AND2_X1 U5466 ( .A1(n8439), .A2(n8441), .ZN(n8287) );
  NOR2_X1 U5467 ( .A1(n9498), .A2(n9499), .ZN(n9497) );
  NOR2_X1 U5468 ( .A1(n9497), .A2(n4570), .ZN(n9511) );
  NOR2_X1 U5469 ( .A1(n5764), .A2(n5751), .ZN(n4570) );
  AND2_X1 U5470 ( .A1(n4559), .A2(n4558), .ZN(n5795) );
  NAND2_X1 U5471 ( .A1(n5775), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4558) );
  NOR2_X1 U5472 ( .A1(n5795), .A2(n5794), .ZN(n5793) );
  AND2_X1 U5473 ( .A1(n4555), .A2(n4554), .ZN(n6581) );
  NAND2_X1 U5474 ( .A1(n6580), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4554) );
  NOR2_X1 U5475 ( .A1(n6964), .A2(n6965), .ZN(n7053) );
  NOR2_X1 U5476 ( .A1(n7053), .A2(n4562), .ZN(n7057) );
  AND2_X1 U5477 ( .A1(n7054), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4562) );
  NAND2_X1 U5478 ( .A1(n7057), .A2(n7056), .ZN(n7224) );
  XNOR2_X1 U5479 ( .A(n8655), .B(n8671), .ZN(n8649) );
  AND2_X1 U5480 ( .A1(n5447), .A2(n7703), .ZN(n8741) );
  OR2_X1 U5481 ( .A1(n8754), .A2(n4546), .ZN(n8738) );
  AND2_X1 U5482 ( .A1(n5424), .A2(n5423), .ZN(n8761) );
  NOR2_X1 U5483 ( .A1(n4664), .A2(n4658), .ZN(n4657) );
  NAND2_X1 U5484 ( .A1(n4665), .A2(n5506), .ZN(n4664) );
  INV_X1 U5485 ( .A(n4660), .ZN(n4658) );
  NAND2_X1 U5486 ( .A1(n4659), .A2(n4660), .ZN(n8788) );
  NOR2_X1 U5487 ( .A1(n8836), .A2(n8905), .ZN(n8819) );
  NAND2_X1 U5488 ( .A1(n4673), .A2(n4336), .ZN(n8847) );
  NOR2_X1 U5489 ( .A1(n8863), .A2(n8916), .ZN(n8862) );
  NOR2_X1 U5490 ( .A1(n8396), .A2(n8411), .ZN(n8834) );
  OR2_X1 U5491 ( .A1(n5349), .A2(n4870), .ZN(n5358) );
  OAI21_X1 U5492 ( .B1(n4459), .B2(n4344), .A(n4774), .ZN(n8852) );
  AOI21_X1 U5493 ( .B1(n4776), .B2(n8275), .A(n4775), .ZN(n4774) );
  INV_X1 U5494 ( .A(n4778), .ZN(n4777) );
  NOR2_X1 U5495 ( .A1(n8932), .A2(n8624), .ZN(n4784) );
  AND2_X1 U5496 ( .A1(n7563), .A2(n4309), .ZN(n4550) );
  NOR2_X1 U5497 ( .A1(n7556), .A2(n8272), .ZN(n7555) );
  INV_X1 U5498 ( .A(n8270), .ZN(n8390) );
  NAND2_X1 U5499 ( .A1(n7174), .A2(n8383), .ZN(n7328) );
  NAND2_X1 U5500 ( .A1(n7174), .A2(n4552), .ZN(n7504) );
  AND2_X1 U5501 ( .A1(n8388), .A2(n8387), .ZN(n8385) );
  NAND2_X1 U5502 ( .A1(n7170), .A2(n5496), .ZN(n7168) );
  NAND2_X1 U5503 ( .A1(n4865), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5255) );
  INV_X1 U5504 ( .A(n5236), .ZN(n4865) );
  NAND2_X1 U5505 ( .A1(n4378), .A2(n8364), .ZN(n5495) );
  OAI21_X1 U5506 ( .B1(n6821), .B2(n5494), .A(n4669), .ZN(n4378) );
  INV_X1 U5507 ( .A(n8374), .ZN(n8267) );
  OR2_X1 U5508 ( .A1(n6997), .A2(n7128), .ZN(n7116) );
  NAND2_X1 U5509 ( .A1(n4766), .A2(n5261), .ZN(n6990) );
  INV_X1 U5510 ( .A(n8264), .ZN(n4766) );
  NAND2_X1 U5511 ( .A1(n4863), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5218) );
  AND2_X1 U5512 ( .A1(n8346), .A2(n5161), .ZN(n4460) );
  OAI21_X1 U5513 ( .B1(n6474), .B2(n5487), .A(n8344), .ZN(n6821) );
  NAND2_X1 U5514 ( .A1(n6403), .A2(n4311), .ZN(n6567) );
  NAND2_X1 U5515 ( .A1(n6399), .A2(n8327), .ZN(n6474) );
  AND2_X1 U5516 ( .A1(n6403), .A2(n9794), .ZN(n6476) );
  NAND2_X1 U5517 ( .A1(n4375), .A2(n8299), .ZN(n6400) );
  NAND2_X1 U5518 ( .A1(n4642), .A2(n4315), .ZN(n4375) );
  NAND2_X1 U5519 ( .A1(n6400), .A2(n8258), .ZN(n6399) );
  OR2_X1 U5520 ( .A1(n6554), .A2(n9785), .ZN(n6359) );
  AOI21_X1 U5521 ( .B1(n4450), .B2(n8255), .A(n4351), .ZN(n4449) );
  INV_X1 U5522 ( .A(n5101), .ZN(n4450) );
  NAND2_X1 U5523 ( .A1(n8323), .A2(n8299), .ZN(n8256) );
  AND4_X1 U5524 ( .A1(n5121), .A2(n5120), .A3(n5119), .A4(n5118), .ZN(n6632)
         );
  NAND2_X1 U5525 ( .A1(n8297), .A2(n8320), .ZN(n8254) );
  NAND2_X1 U5526 ( .A1(n5483), .A2(n5482), .ZN(n7660) );
  OR2_X1 U5527 ( .A1(n5097), .A2(n5657), .ZN(n5080) );
  NOR2_X1 U5528 ( .A1(n6450), .A2(n9771), .ZN(n6539) );
  NAND2_X1 U5529 ( .A1(n6389), .A2(n8315), .ZN(n8305) );
  NAND2_X1 U5530 ( .A1(n6205), .A2(n6391), .ZN(n8313) );
  NOR2_X1 U5531 ( .A1(n6771), .A2(n6770), .ZN(n6217) );
  OR2_X1 U5532 ( .A1(n6208), .A2(n6207), .ZN(n6218) );
  NAND2_X1 U5533 ( .A1(n5415), .A2(n5414), .ZN(n8889) );
  NAND2_X1 U5534 ( .A1(n5184), .A2(n5183), .ZN(n6975) );
  OR3_X1 U5535 ( .A1(n6206), .A2(n5633), .A3(n6207), .ZN(n6370) );
  AND2_X1 U5536 ( .A1(n4542), .A2(n4887), .ZN(n4539) );
  AND2_X1 U5537 ( .A1(n4314), .A2(n5021), .ZN(n4542) );
  AND2_X1 U5538 ( .A1(n5036), .A2(n4887), .ZN(n5526) );
  NAND2_X1 U5539 ( .A1(n5036), .A2(n4757), .ZN(n5480) );
  NOR2_X1 U5540 ( .A1(n4758), .A2(n4347), .ZN(n4757) );
  INV_X1 U5541 ( .A(n4759), .ZN(n4758) );
  AND2_X1 U5542 ( .A1(n5199), .A2(n5210), .ZN(n6963) );
  AND2_X1 U5543 ( .A1(n5148), .A2(n5142), .ZN(n5830) );
  INV_X1 U5544 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U5545 ( .A1(n9077), .A2(n9080), .ZN(n4440) );
  INV_X1 U5546 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9025) );
  NOR2_X1 U5547 ( .A1(n5936), .A2(n5935), .ZN(n7687) );
  NAND2_X1 U5548 ( .A1(n5934), .A2(n5933), .ZN(n5935) );
  INV_X1 U5549 ( .A(n9047), .ZN(n4831) );
  INV_X1 U5550 ( .A(n4829), .ZN(n4826) );
  NAND2_X1 U5551 ( .A1(n6843), .A2(n6842), .ZN(n6919) );
  NAND2_X1 U5552 ( .A1(n8479), .A2(n8478), .ZN(n9078) );
  NAND2_X1 U5553 ( .A1(n4428), .A2(n4425), .ZN(n8101) );
  AND2_X1 U5554 ( .A1(n8020), .A2(n4426), .ZN(n4425) );
  NAND2_X1 U5555 ( .A1(n4427), .A2(n8010), .ZN(n4426) );
  AND2_X1 U5556 ( .A1(n9386), .A2(n8119), .ZN(n8091) );
  AND2_X1 U5557 ( .A1(n4530), .A2(n4529), .ZN(n9625) );
  NAND2_X1 U5558 ( .A1(n6346), .A2(n6022), .ZN(n4529) );
  AOI21_X1 U5559 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9125), .A(n9121), .ZN(
        n9651) );
  NOR2_X1 U5560 ( .A1(n6595), .A2(n6594), .ZN(n7306) );
  XNOR2_X1 U5561 ( .A(n7307), .B(n9659), .ZN(n9662) );
  OR2_X1 U5562 ( .A1(n9135), .A2(n9136), .ZN(n4525) );
  AND2_X1 U5563 ( .A1(n4523), .A2(n4522), .ZN(n9161) );
  NAND2_X1 U5564 ( .A1(n9158), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4522) );
  NOR2_X1 U5565 ( .A1(n9161), .A2(n9160), .ZN(n9165) );
  INV_X1 U5566 ( .A(n4621), .ZN(n4612) );
  NAND2_X1 U5567 ( .A1(n4617), .A2(n4621), .ZN(n4613) );
  AOI21_X1 U5568 ( .B1(n4617), .B2(n4616), .A(n4352), .ZN(n4615) );
  NOR2_X1 U5569 ( .A1(n9251), .A2(n4509), .ZN(n9220) );
  INV_X1 U5570 ( .A(n4511), .ZN(n4509) );
  OR2_X1 U5571 ( .A1(n9262), .A2(n9418), .ZN(n9251) );
  NOR2_X1 U5572 ( .A1(n9251), .A2(n9411), .ZN(n9233) );
  OR2_X1 U5573 ( .A1(n8023), .A2(n8130), .ZN(n9246) );
  AND2_X1 U5574 ( .A1(n9293), .A2(n9284), .ZN(n9280) );
  AND2_X1 U5575 ( .A1(n9268), .A2(n8144), .ZN(n9285) );
  OAI21_X1 U5576 ( .B1(n9326), .B2(n4697), .A(n4694), .ZN(n9300) );
  INV_X1 U5577 ( .A(n4698), .ZN(n4697) );
  AND2_X1 U5578 ( .A1(n8142), .A2(n4695), .ZN(n4694) );
  NAND2_X1 U5579 ( .A1(n4698), .A2(n4696), .ZN(n4695) );
  OR2_X1 U5580 ( .A1(n7808), .A2(n6322), .ZN(n7809) );
  NAND2_X1 U5581 ( .A1(n9347), .A2(n8138), .ZN(n9350) );
  NOR2_X1 U5582 ( .A1(n9363), .A2(n4516), .ZN(n9341) );
  NOR2_X1 U5583 ( .A1(n9363), .A2(n9453), .ZN(n9362) );
  INV_X1 U5584 ( .A(n4708), .ZN(n4707) );
  AOI21_X1 U5585 ( .B1(n4708), .B2(n4706), .A(n4705), .ZN(n4704) );
  AND2_X1 U5586 ( .A1(n4709), .A2(n8135), .ZN(n4708) );
  NAND2_X1 U5587 ( .A1(n6320), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7344) );
  INV_X1 U5588 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7343) );
  OR2_X1 U5589 ( .A1(n7344), .A2(n7343), .ZN(n7459) );
  AND2_X1 U5590 ( .A1(n6949), .A2(n4502), .ZN(n7357) );
  AND2_X1 U5591 ( .A1(n4503), .A2(n9544), .ZN(n4502) );
  AOI21_X1 U5592 ( .B1(n4691), .B2(n7136), .A(n4689), .ZN(n4688) );
  INV_X1 U5593 ( .A(n4691), .ZN(n4690) );
  INV_X1 U5594 ( .A(n7833), .ZN(n4689) );
  NAND2_X1 U5595 ( .A1(n6949), .A2(n4503), .ZN(n7251) );
  AOI21_X1 U5596 ( .B1(n7137), .B2(n7136), .A(n7135), .ZN(n7239) );
  NAND2_X1 U5597 ( .A1(n4693), .A2(n4691), .ZN(n4857) );
  NAND2_X1 U5598 ( .A1(n4693), .A2(n7954), .ZN(n7145) );
  INV_X1 U5599 ( .A(n9107), .ZN(n7237) );
  NAND2_X1 U5600 ( .A1(n6949), .A2(n9554), .ZN(n7037) );
  AND2_X1 U5601 ( .A1(n6944), .A2(n7848), .ZN(n6945) );
  NAND2_X1 U5602 ( .A1(n4712), .A2(n4711), .ZN(n6944) );
  AND2_X1 U5603 ( .A1(n4715), .A2(n7940), .ZN(n4711) );
  NAND2_X1 U5604 ( .A1(n4712), .A2(n7940), .ZN(n6943) );
  AND3_X1 U5605 ( .A1(n6499), .A2(n4519), .A3(n4518), .ZN(n6869) );
  NOR2_X1 U5606 ( .A1(n6907), .A2(n6861), .ZN(n4518) );
  NAND2_X1 U5607 ( .A1(n6680), .A2(n6679), .ZN(n6683) );
  AND2_X1 U5608 ( .A1(n7940), .A2(n7933), .ZN(n8036) );
  NAND2_X1 U5609 ( .A1(n6675), .A2(n7926), .ZN(n6780) );
  NAND2_X1 U5610 ( .A1(n6499), .A2(n4519), .ZN(n6689) );
  AND2_X1 U5611 ( .A1(n6499), .A2(n6605), .ZN(n6620) );
  OAI21_X1 U5612 ( .B1(n6068), .B2(n6067), .A(n4431), .ZN(n6488) );
  NOR2_X1 U5613 ( .A1(n4337), .A2(n4432), .ZN(n4431) );
  NOR2_X1 U5614 ( .A1(n5944), .A2(n6070), .ZN(n4432) );
  OR2_X1 U5615 ( .A1(n6609), .A2(n6607), .ZN(n6490) );
  AOI21_X1 U5616 ( .B1(n6458), .B2(n8063), .A(n6410), .ZN(n6493) );
  NAND2_X1 U5617 ( .A1(n4703), .A2(n6409), .ZN(n8064) );
  NOR2_X1 U5618 ( .A1(n6161), .A2(n4307), .ZN(n6432) );
  NAND2_X1 U5619 ( .A1(n6240), .A2(n6239), .ZN(n6241) );
  NAND2_X1 U5620 ( .A1(n7841), .A2(n5923), .ZN(n6161) );
  NAND2_X1 U5621 ( .A1(n7771), .A2(n7770), .ZN(n9426) );
  NAND2_X1 U5622 ( .A1(n7457), .A2(n7456), .ZN(n9459) );
  OAI211_X1 U5623 ( .C1(n5944), .C2(n6056), .A(n6055), .B(n6054), .ZN(n6526)
         );
  AND2_X1 U5624 ( .A1(n5891), .A2(n5890), .ZN(n5907) );
  OR2_X1 U5625 ( .A1(n5963), .A2(n8104), .ZN(n9696) );
  INV_X1 U5626 ( .A(n9696), .ZN(n9437) );
  INV_X1 U5627 ( .A(n9710), .ZN(n9465) );
  INV_X1 U5628 ( .A(SI_21_), .ZN(n9873) );
  XNOR2_X1 U5629 ( .A(n7728), .B(n7727), .ZN(n8973) );
  XNOR2_X1 U5630 ( .A(n7711), .B(n5463), .ZN(n7897) );
  XNOR2_X1 U5631 ( .A(n5441), .B(n5440), .ZN(n7733) );
  XNOR2_X1 U5632 ( .A(n5020), .B(n5386), .ZN(n7861) );
  INV_X1 U5633 ( .A(n4842), .ZN(n4840) );
  XNOR2_X1 U5634 ( .A(n5046), .B(n5045), .ZN(n7593) );
  XNOR2_X1 U5635 ( .A(n5209), .B(n5208), .ZN(n6920) );
  NAND2_X1 U5636 ( .A1(n4770), .A2(n4946), .ZN(n5194) );
  NAND2_X1 U5637 ( .A1(n5181), .A2(n4319), .ZN(n4770) );
  XNOR2_X1 U5638 ( .A(n5181), .B(n4319), .ZN(n6706) );
  NAND2_X1 U5639 ( .A1(n4572), .A2(n4762), .ZN(n5163) );
  NAND2_X1 U5640 ( .A1(n4924), .A2(n4923), .ZN(n5125) );
  XNOR2_X1 U5641 ( .A(n4526), .B(P1_IR_REG_3__SCAN_IN), .ZN(n5861) );
  OAI21_X1 U5642 ( .B1(n5662), .B2(P1_IR_REG_2__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U5643 ( .A1(n4528), .A2(n4527), .ZN(n5662) );
  XNOR2_X1 U5644 ( .A(n4908), .B(n4907), .ZN(n5056) );
  AND4_X1 U5645 ( .A1(n5179), .A2(n5178), .A3(n5177), .A4(n5176), .ZN(n6820)
         );
  NAND2_X1 U5646 ( .A1(n6626), .A2(n5621), .ZN(n5631) );
  NAND2_X1 U5647 ( .A1(n4743), .A2(n4745), .ZN(n8549) );
  INV_X1 U5648 ( .A(n4746), .ZN(n4745) );
  OAI21_X1 U5649 ( .B1(n4747), .B2(n8193), .A(n8544), .ZN(n4746) );
  AND4_X1 U5650 ( .A1(n5260), .A2(n5259), .A3(n5258), .A4(n5257), .ZN(n7211)
         );
  AND4_X1 U5651 ( .A1(n5299), .A2(n5298), .A3(n5297), .A4(n5296), .ZN(n8382)
         );
  NAND2_X1 U5652 ( .A1(n5277), .A2(n5276), .ZN(n7214) );
  AND2_X1 U5653 ( .A1(n4390), .A2(n4389), .ZN(n8558) );
  AND2_X1 U5654 ( .A1(n8178), .A2(n4391), .ZN(n4390) );
  NAND2_X1 U5655 ( .A1(n6796), .A2(n6752), .ZN(n7645) );
  INV_X1 U5656 ( .A(n6542), .ZN(n9780) );
  NAND2_X1 U5657 ( .A1(n4403), .A2(n7577), .ZN(n7587) );
  OAI21_X1 U5658 ( .B1(n7448), .B2(n4400), .A(n4398), .ZN(n4403) );
  NAND2_X1 U5659 ( .A1(n5328), .A2(n5327), .ZN(n8927) );
  AOI21_X1 U5660 ( .B1(n8756), .B2(n4469), .A(n5438), .ZN(n8747) );
  NAND2_X1 U5661 ( .A1(n5445), .A2(n5444), .ZN(n8878) );
  AND4_X1 U5662 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n7655)
         );
  NAND2_X1 U5663 ( .A1(n5308), .A2(n5307), .ZN(n8941) );
  AND4_X1 U5664 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n7509)
         );
  NAND2_X1 U5665 ( .A1(n7448), .A2(n7392), .ZN(n7477) );
  NAND2_X1 U5666 ( .A1(n5609), .A2(n5647), .ZN(n6805) );
  NAND2_X1 U5667 ( .A1(n6805), .A2(n4721), .ZN(n8229) );
  NAND2_X1 U5668 ( .A1(n7629), .A2(n7628), .ZN(n8172) );
  AND4_X1 U5669 ( .A1(n5284), .A2(n5283), .A3(n5282), .A4(n5281), .ZN(n7261)
         );
  NAND2_X1 U5670 ( .A1(n5253), .A2(n5252), .ZN(n8952) );
  NAND2_X1 U5671 ( .A1(n8568), .A2(n8567), .ZN(n8598) );
  AND4_X1 U5672 ( .A1(n5044), .A2(n5043), .A3(n5042), .A4(n5041), .ZN(n7565)
         );
  AND3_X1 U5673 ( .A1(n5334), .A2(n5333), .A3(n5332), .ZN(n7633) );
  OR2_X1 U5674 ( .A1(n6888), .A2(n8859), .ZN(n8607) );
  NAND2_X1 U5675 ( .A1(n4397), .A2(n4404), .ZN(n7573) );
  NAND2_X1 U5676 ( .A1(n7448), .A2(n4401), .ZN(n4397) );
  AND4_X1 U5677 ( .A1(n5158), .A2(n5157), .A3(n5156), .A4(n5155), .ZN(n6741)
         );
  OR2_X1 U5678 ( .A1(n6888), .A2(n8861), .ZN(n8608) );
  INV_X1 U5679 ( .A(n5613), .ZN(n4720) );
  INV_X1 U5680 ( .A(n8545), .ZN(n4406) );
  NAND2_X1 U5681 ( .A1(n8208), .A2(n8209), .ZN(n4405) );
  NAND2_X1 U5682 ( .A1(n4741), .A2(n4740), .ZN(n8208) );
  NAND2_X1 U5683 ( .A1(n8577), .A2(n8576), .ZN(n4740) );
  NAND2_X1 U5684 ( .A1(n4753), .A2(n7445), .ZN(n7698) );
  INV_X1 U5685 ( .A(n4754), .ZN(n4753) );
  OR2_X1 U5686 ( .A1(n5215), .A2(n5073), .ZN(n5075) );
  INV_X1 U5687 ( .A(n4559), .ZN(n5774) );
  INV_X1 U5688 ( .A(n4557), .ZN(n6374) );
  INV_X1 U5689 ( .A(n4555), .ZN(n6579) );
  NOR2_X1 U5690 ( .A1(n5233), .A2(n5232), .ZN(n7222) );
  INV_X1 U5691 ( .A(n7410), .ZN(n7411) );
  NAND2_X1 U5692 ( .A1(n8699), .A2(n4569), .ZN(n8708) );
  NOR2_X1 U5693 ( .A1(n4568), .A2(n4567), .ZN(n8700) );
  INV_X1 U5694 ( .A(n8698), .ZN(n4567) );
  AND2_X1 U5695 ( .A1(n5769), .A2(n5768), .ZN(n9728) );
  NAND2_X1 U5696 ( .A1(n5769), .A2(n5508), .ZN(n9731) );
  INV_X1 U5697 ( .A(n8246), .ZN(n8874) );
  OR3_X1 U5698 ( .A1(n5446), .A2(n8551), .A3(n8200), .ZN(n7703) );
  INV_X1 U5699 ( .A(n5514), .ZN(n5515) );
  XNOR2_X1 U5700 ( .A(n8235), .B(n8434), .ZN(n4380) );
  AOI22_X1 U5701 ( .A1(n8615), .A2(n7566), .B1(n8726), .B2(n8614), .ZN(n5514)
         );
  INV_X1 U5702 ( .A(n8878), .ZN(n8743) );
  NAND2_X1 U5703 ( .A1(n4455), .A2(n4456), .ZN(n8753) );
  NAND2_X1 U5704 ( .A1(n4787), .A2(n4313), .ZN(n4455) );
  NAND2_X1 U5705 ( .A1(n4787), .A2(n4785), .ZN(n8769) );
  NAND2_X1 U5706 ( .A1(n5400), .A2(n5399), .ZN(n8894) );
  AND2_X1 U5707 ( .A1(n4793), .A2(n4792), .ZN(n8785) );
  INV_X1 U5708 ( .A(n4663), .ZN(n8806) );
  NAND2_X1 U5709 ( .A1(n8903), .A2(n4852), .ZN(n8798) );
  AND2_X1 U5710 ( .A1(n5357), .A2(n5356), .ZN(n8842) );
  NAND2_X1 U5711 ( .A1(n7623), .A2(n8407), .ZN(n8854) );
  OAI21_X1 U5712 ( .B1(n7556), .B2(n4779), .A(n4778), .ZN(n7615) );
  NAND2_X1 U5713 ( .A1(n4670), .A2(n4669), .ZN(n6993) );
  NAND2_X1 U5714 ( .A1(n4670), .A2(n5493), .ZN(n6896) );
  AND2_X1 U5715 ( .A1(n4461), .A2(n5159), .ZN(n6473) );
  BUF_X1 U5716 ( .A(n5516), .Z(n9771) );
  NOR2_X1 U5717 ( .A1(n9752), .A2(n9749), .ZN(n8823) );
  INV_X1 U5718 ( .A(n8869), .ZN(n8828) );
  INV_X1 U5719 ( .A(n8736), .ZN(n8864) );
  INV_X1 U5720 ( .A(n8823), .ZN(n8873) );
  AOI211_X1 U5721 ( .C1(n9772), .C2(n9525), .A(n9524), .B(n9523), .ZN(n9533)
         );
  OR2_X1 U5722 ( .A1(n6370), .A2(n5627), .ZN(n9816) );
  NAND2_X1 U5723 ( .A1(n4465), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4890) );
  NAND2_X1 U5724 ( .A1(n4891), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4892) );
  NAND2_X1 U5725 ( .A1(n5036), .A2(n4463), .ZN(n4891) );
  INV_X1 U5726 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7275) );
  INV_X1 U5727 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7076) );
  XNOR2_X1 U5728 ( .A(n5525), .B(n5524), .ZN(n7077) );
  INV_X1 U5729 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U5730 ( .A1(n5523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5525) );
  INV_X1 U5731 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9886) );
  INV_X1 U5732 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7006) );
  INV_X1 U5733 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8207) );
  INV_X1 U5734 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6271) );
  INV_X1 U5735 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9884) );
  INV_X1 U5736 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6181) );
  INV_X1 U5737 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5984) );
  INV_X1 U5738 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5820) );
  INV_X1 U5739 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5720) );
  NOR2_X1 U5740 ( .A1(n4444), .A2(n4443), .ZN(n4442) );
  INV_X1 U5741 ( .A(n8537), .ZN(n4443) );
  INV_X1 U5742 ( .A(n9303), .ZN(n9026) );
  NAND2_X1 U5743 ( .A1(n4814), .A2(n8519), .ZN(n8983) );
  NAND2_X1 U5744 ( .A1(n4322), .A2(n4815), .ZN(n4814) );
  AND2_X1 U5745 ( .A1(n6650), .A2(n6653), .ZN(n4837) );
  AND2_X1 U5746 ( .A1(n6658), .A2(n6657), .ZN(n6713) );
  NAND2_X1 U5747 ( .A1(n7783), .A2(n7782), .ZN(n9432) );
  NAND2_X1 U5748 ( .A1(n8982), .A2(n4807), .ZN(n4799) );
  NAND2_X1 U5749 ( .A1(n4808), .A2(n4807), .ZN(n4800) );
  INV_X1 U5750 ( .A(n9379), .ZN(n7610) );
  NAND2_X1 U5751 ( .A1(n7601), .A2(n7600), .ZN(n7602) );
  NOR2_X1 U5752 ( .A1(n4808), .A2(n8982), .ZN(n9039) );
  NAND2_X1 U5753 ( .A1(n4836), .A2(n4835), .ZN(n4834) );
  NAND2_X1 U5754 ( .A1(n7790), .A2(n7789), .ZN(n9436) );
  NAND2_X1 U5755 ( .A1(n7182), .A2(n7181), .ZN(n7421) );
  NAND2_X1 U5756 ( .A1(n5941), .A2(n6028), .ZN(n4638) );
  AND2_X1 U5757 ( .A1(n5974), .A2(n5973), .ZN(n9092) );
  AND2_X1 U5758 ( .A1(n7887), .A2(n7747), .ZN(n9222) );
  OR2_X1 U5759 ( .A1(n6136), .A2(n6135), .ZN(n9099) );
  NAND2_X1 U5760 ( .A1(n5962), .A2(n5961), .ZN(n9086) );
  INV_X1 U5761 ( .A(n9092), .ZN(n9051) );
  NAND2_X1 U5762 ( .A1(n4433), .A2(n7490), .ZN(n7517) );
  NAND2_X1 U5763 ( .A1(n4438), .A2(n7486), .ZN(n4433) );
  INV_X1 U5764 ( .A(n5899), .ZN(n8104) );
  INV_X1 U5765 ( .A(n9694), .ZN(n8107) );
  NAND2_X1 U5766 ( .A1(n7828), .A2(n7827), .ZN(n9287) );
  NAND4_X1 U5767 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n9115)
         );
  NAND4_X1 U5768 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n9116)
         );
  NAND4_X1 U5769 ( .A1(n6008), .A2(n6007), .A3(n6006), .A4(n6005), .ZN(n9117)
         );
  NAND3_X2 U5770 ( .A1(n4675), .A2(n5901), .A3(n4676), .ZN(n9120) );
  INV_X1 U5771 ( .A(n4678), .ZN(n4675) );
  AND2_X1 U5772 ( .A1(n5681), .A2(n5680), .ZN(n5918) );
  NOR2_X1 U5773 ( .A1(n9597), .A2(n5865), .ZN(n5913) );
  NOR2_X1 U5774 ( .A1(n5913), .A2(n5912), .ZN(n5911) );
  INV_X1 U5775 ( .A(n4530), .ZN(n6345) );
  AND2_X1 U5776 ( .A1(n5819), .A2(n5818), .ZN(n9646) );
  INV_X1 U5777 ( .A(n4523), .ZN(n9157) );
  INV_X1 U5778 ( .A(n4525), .ZN(n9139) );
  INV_X1 U5779 ( .A(n9676), .ZN(n9637) );
  AND2_X1 U5780 ( .A1(n5848), .A2(n5736), .ZN(n9678) );
  INV_X1 U5781 ( .A(n8114), .ZN(n9386) );
  NAND2_X1 U5782 ( .A1(n7715), .A2(n7714), .ZN(n9387) );
  OAI21_X1 U5783 ( .B1(n9238), .B2(n4684), .A(n4682), .ZN(n9206) );
  AOI21_X1 U5784 ( .B1(n4685), .B2(n4683), .A(n8154), .ZN(n4682) );
  AND2_X1 U5785 ( .A1(n4686), .A2(n8152), .ZN(n4858) );
  NAND2_X1 U5786 ( .A1(n4614), .A2(n4617), .ZN(n9219) );
  NAND2_X1 U5787 ( .A1(n9245), .A2(n4618), .ZN(n4614) );
  OAI21_X1 U5788 ( .B1(n9245), .B2(n8130), .A(n8129), .ZN(n9232) );
  INV_X1 U5789 ( .A(n9421), .ZN(n9267) );
  INV_X1 U5790 ( .A(n9426), .ZN(n9284) );
  NAND2_X1 U5791 ( .A1(n4700), .A2(n8140), .ZN(n9315) );
  NAND2_X1 U5792 ( .A1(n4602), .A2(n4606), .ZN(n9308) );
  NAND2_X1 U5793 ( .A1(n9340), .A2(n4607), .ZN(n4602) );
  AND2_X1 U5794 ( .A1(n4609), .A2(n4608), .ZN(n9325) );
  INV_X1 U5795 ( .A(n4611), .ZN(n4608) );
  NAND2_X1 U5796 ( .A1(n9340), .A2(n9348), .ZN(n4609) );
  NAND2_X1 U5797 ( .A1(n7341), .A2(n7340), .ZN(n7496) );
  INV_X1 U5798 ( .A(n6515), .ZN(n6605) );
  INV_X1 U5799 ( .A(n9364), .ZN(n9183) );
  AND2_X1 U5800 ( .A1(n9370), .A2(n9437), .ZN(n9322) );
  INV_X1 U5801 ( .A(n9692), .ZN(n9860) );
  INV_X1 U5802 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5694) );
  CLKBUF_X1 U5803 ( .A(n5735), .Z(n5736) );
  CLKBUF_X1 U5804 ( .A(n5594), .Z(n8117) );
  INV_X1 U5805 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U5806 ( .A1(n5569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5566) );
  INV_X1 U5807 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7757) );
  INV_X1 U5808 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7862) );
  XNOR2_X1 U5809 ( .A(n5571), .B(n5570), .ZN(n7079) );
  INV_X1 U5810 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7817) );
  XNOR2_X1 U5811 ( .A(n5371), .B(n5370), .ZN(n7816) );
  NAND2_X1 U5812 ( .A1(n4599), .A2(n4597), .ZN(n5385) );
  INV_X1 U5813 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5582) );
  INV_X1 U5814 ( .A(n5900), .ZN(n8092) );
  INV_X1 U5815 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7788) );
  INV_X1 U5816 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6589) );
  AND2_X1 U5817 ( .A1(n6229), .A2(n6484), .ZN(n9172) );
  INV_X1 U5818 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6180) );
  INV_X1 U5819 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6155) );
  INV_X1 U5820 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5982) );
  OR2_X1 U5821 ( .A1(n5981), .A2(n5980), .ZN(n6349) );
  INV_X1 U5822 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9865) );
  NAND2_X1 U5823 ( .A1(n4764), .A2(n4931), .ZN(n5146) );
  XNOR2_X1 U5824 ( .A(n5137), .B(n5138), .ZN(n6119) );
  XNOR2_X1 U5825 ( .A(n5125), .B(n5124), .ZN(n6068) );
  INV_X1 U5826 ( .A(n9602), .ZN(n6056) );
  NOR2_X1 U5827 ( .A1(n7299), .A2(n10057), .ZN(n9859) );
  AOI21_X1 U5828 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9857), .ZN(n9856) );
  NOR2_X1 U5829 ( .A1(n9856), .A2(n9855), .ZN(n9854) );
  AOI21_X1 U5830 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9854), .ZN(n9853) );
  OAI21_X1 U5831 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9851), .ZN(n9849) );
  AND3_X1 U5832 ( .A1(n4473), .A2(n4471), .A3(n4470), .ZN(n8458) );
  INV_X1 U5833 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4902) );
  OR2_X1 U5834 ( .A1(n9011), .A2(n4844), .ZN(n9019) );
  OAI21_X1 U5835 ( .B1(n9179), .B2(n9178), .A(n4531), .ZN(P1_U3260) );
  AOI21_X1 U5836 ( .B1(n4533), .B2(n9178), .A(n4532), .ZN(n4531) );
  OAI21_X1 U5837 ( .B1(n9671), .B2(n4903), .A(n9180), .ZN(n4532) );
  AOI211_X1 U5838 ( .C1(n9391), .C2(n9370), .A(n8166), .B(n8165), .ZN(n8167)
         );
  AND2_X1 U5839 ( .A1(n9393), .A2(n9394), .ZN(n4632) );
  NAND2_X1 U5840 ( .A1(n9719), .A2(n9706), .ZN(n4630) );
  INV_X1 U5841 ( .A(n4626), .ZN(n4625) );
  OAI21_X1 U5842 ( .B1(n9393), .B2(n9717), .A(n4623), .ZN(n4626) );
  INV_X1 U5843 ( .A(n8744), .ZN(n4649) );
  INV_X1 U5844 ( .A(n6092), .ZN(n9007) );
  INV_X2 U5845 ( .A(n9007), .ZN(n8508) );
  AND2_X1 U5846 ( .A1(n4324), .A2(n5208), .ZN(n4308) );
  AND2_X1 U5847 ( .A1(n4552), .A2(n4551), .ZN(n4309) );
  AND2_X1 U5848 ( .A1(n4656), .A2(n8303), .ZN(n4310) );
  INV_X1 U5849 ( .A(n7244), .ZN(n5700) );
  INV_X1 U5850 ( .A(n5086), .ZN(n5309) );
  NAND2_X1 U5851 ( .A1(n9491), .A2(n7639), .ZN(n4680) );
  NAND2_X1 U5852 ( .A1(n5049), .A2(n5048), .ZN(n5318) );
  NAND2_X1 U5853 ( .A1(n4841), .A2(n4842), .ZN(n5979) );
  NAND2_X1 U5854 ( .A1(n4585), .A2(n4324), .ZN(n4584) );
  AND2_X1 U5855 ( .A1(n6509), .A2(n9794), .ZN(n4311) );
  NAND2_X1 U5856 ( .A1(n6632), .A2(n9740), .ZN(n4312) );
  INV_X1 U5857 ( .A(n8789), .ZN(n4666) );
  AND2_X1 U5858 ( .A1(n4785), .A2(n4458), .ZN(n4313) );
  INV_X1 U5859 ( .A(n8771), .ZN(n4665) );
  AND2_X1 U5860 ( .A1(n4888), .A2(n4674), .ZN(n4314) );
  INV_X1 U5861 ( .A(n8346), .ZN(n8332) );
  AND2_X1 U5862 ( .A1(n8323), .A2(n8321), .ZN(n4315) );
  INV_X1 U5863 ( .A(n8982), .ZN(n4794) );
  NAND2_X1 U5864 ( .A1(n4357), .A2(n4622), .ZN(n4617) );
  AND2_X1 U5865 ( .A1(n4663), .A2(n8419), .ZN(n4316) );
  AND2_X1 U5866 ( .A1(n5040), .A2(n5039), .ZN(n7563) );
  INV_X1 U5867 ( .A(n7563), .ZN(n8932) );
  AND2_X1 U5868 ( .A1(n4354), .A2(n4847), .ZN(n4317) );
  INV_X1 U5869 ( .A(n9403), .ZN(n9215) );
  NAND2_X1 U5870 ( .A1(n7736), .A2(n7735), .ZN(n9403) );
  AND2_X1 U5871 ( .A1(n8469), .A2(n8468), .ZN(n4318) );
  INV_X1 U5872 ( .A(n8255), .ZN(n4451) );
  NAND2_X1 U5873 ( .A1(n6949), .A2(n4505), .ZN(n4506) );
  XNOR2_X1 U5874 ( .A(n5479), .B(n5478), .ZN(n8284) );
  INV_X1 U5875 ( .A(n8284), .ZN(n8303) );
  AND2_X1 U5876 ( .A1(n5517), .A2(n8284), .ZN(n9763) );
  AND2_X1 U5877 ( .A1(n4946), .A2(n4945), .ZN(n4319) );
  INV_X1 U5878 ( .A(n6114), .ZN(n7750) );
  NAND2_X2 U5879 ( .A1(n6000), .A2(n5925), .ZN(n6095) );
  NAND2_X1 U5880 ( .A1(n4809), .A2(n4811), .ZN(n4808) );
  NAND4_X1 U5881 ( .A1(n5711), .A2(n5710), .A3(n5709), .A4(n5708), .ZN(n5931)
         );
  INV_X1 U5882 ( .A(n8639), .ZN(n5100) );
  OAI21_X1 U5883 ( .B1(n5887), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5885) );
  OR2_X1 U5884 ( .A1(n8754), .A2(n4544), .ZN(n4320) );
  INV_X1 U5885 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4527) );
  NOR2_X1 U5886 ( .A1(n5576), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5817) );
  AND2_X1 U5887 ( .A1(n4700), .A2(n4698), .ZN(n4321) );
  NAND2_X2 U5888 ( .A1(n5707), .A2(n5706), .ZN(n7868) );
  OR2_X1 U5889 ( .A1(n8515), .A2(n8514), .ZN(n4322) );
  INV_X1 U5890 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9486) );
  OR2_X1 U5891 ( .A1(n5439), .A2(n4454), .ZN(n4323) );
  NAND2_X1 U5892 ( .A1(n4974), .A2(n4973), .ZN(n4324) );
  NAND2_X1 U5893 ( .A1(n4655), .A2(n8436), .ZN(n4654) );
  NAND2_X1 U5894 ( .A1(n5900), .A2(n5899), .ZN(n5925) );
  XNOR2_X1 U5895 ( .A(n5520), .B(n5481), .ZN(n5517) );
  NAND2_X1 U5896 ( .A1(n7700), .A2(n8746), .ZN(n4325) );
  NAND2_X1 U5897 ( .A1(n8916), .A2(n8844), .ZN(n4326) );
  NOR2_X1 U5898 ( .A1(n8745), .A2(n8744), .ZN(n4327) );
  NAND2_X1 U5899 ( .A1(n4834), .A2(n4832), .ZN(n9046) );
  AND2_X1 U5900 ( .A1(n7369), .A2(n4725), .ZN(n4328) );
  AND2_X1 U5901 ( .A1(n9444), .A2(n9352), .ZN(n4329) );
  AND2_X1 U5902 ( .A1(n4389), .A2(n8563), .ZN(n4330) );
  INV_X1 U5903 ( .A(n8808), .ZN(n4662) );
  AND2_X1 U5904 ( .A1(n8326), .A2(n8435), .ZN(n4331) );
  INV_X1 U5905 ( .A(n9040), .ZN(n4807) );
  INV_X1 U5906 ( .A(n4374), .ZN(n6205) );
  XNOR2_X1 U5907 ( .A(n5057), .B(n5058), .ZN(n5764) );
  NOR2_X1 U5908 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5674) );
  NAND2_X1 U5909 ( .A1(n7235), .A2(n7234), .ZN(n7832) );
  INV_X1 U5910 ( .A(n7832), .ZN(n9544) );
  NAND2_X1 U5911 ( .A1(n7263), .A2(n5300), .ZN(n7322) );
  INV_X1 U5912 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U5913 ( .A1(n7007), .A2(n7656), .ZN(n4332) );
  NAND2_X1 U5914 ( .A1(n5290), .A2(n5289), .ZN(n8947) );
  AND2_X1 U5915 ( .A1(n4762), .A2(n4571), .ZN(n4333) );
  AND3_X1 U5916 ( .A1(n5091), .A2(n5088), .A3(n5089), .ZN(n4334) );
  OR2_X1 U5917 ( .A1(n5585), .A2(n5584), .ZN(n4335) );
  AND2_X1 U5918 ( .A1(n8834), .A2(n4326), .ZN(n4336) );
  INV_X1 U5919 ( .A(n8992), .ZN(n4835) );
  INV_X1 U5920 ( .A(n7500), .ZN(n4895) );
  XNOR2_X1 U5921 ( .A(n4892), .B(n4464), .ZN(n7500) );
  NOR2_X1 U5922 ( .A1(n6120), .A2(n6069), .ZN(n4337) );
  NAND2_X1 U5923 ( .A1(n6922), .A2(n6921), .ZN(n7835) );
  AND2_X1 U5924 ( .A1(n8434), .A2(n8433), .ZN(n4338) );
  INV_X1 U5925 ( .A(n9406), .ZN(n9224) );
  NAND2_X1 U5926 ( .A1(n7746), .A2(n7745), .ZN(n9406) );
  NOR3_X1 U5927 ( .A1(n9251), .A2(n9396), .A3(n4510), .ZN(n4507) );
  NOR2_X1 U5928 ( .A1(n5486), .A2(n4643), .ZN(n4339) );
  NOR2_X1 U5929 ( .A1(n4390), .A2(n4389), .ZN(n4340) );
  AND2_X1 U5930 ( .A1(n8026), .A2(n8140), .ZN(n9324) );
  INV_X1 U5931 ( .A(n9324), .ZN(n4696) );
  AND2_X1 U5932 ( .A1(n5138), .A2(n5145), .ZN(n4341) );
  INV_X1 U5933 ( .A(n4325), .ZN(n4652) );
  INV_X1 U5934 ( .A(n4654), .ZN(n4653) );
  AND2_X1 U5935 ( .A1(n5317), .A2(n5300), .ZN(n4342) );
  INV_X1 U5936 ( .A(n4508), .ZN(n9210) );
  NOR2_X1 U5937 ( .A1(n9251), .A2(n4510), .ZN(n4508) );
  AND2_X1 U5938 ( .A1(n7096), .A2(n7094), .ZN(n4343) );
  OR2_X1 U5939 ( .A1(n7620), .A2(n4777), .ZN(n4344) );
  NAND2_X1 U5940 ( .A1(n4673), .A2(n4326), .ZN(n4345) );
  INV_X1 U5941 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4889) );
  INV_X1 U5942 ( .A(n4377), .ZN(n8770) );
  NAND2_X1 U5943 ( .A1(n4659), .A2(n4657), .ZN(n4377) );
  OR2_X1 U5944 ( .A1(n5580), .A2(n5579), .ZN(n4346) );
  INV_X1 U5945 ( .A(n4833), .ZN(n4832) );
  NOR2_X1 U5946 ( .A1(n8487), .A2(n8488), .ZN(n4833) );
  INV_X1 U5947 ( .A(n4490), .ZN(n4488) );
  NAND3_X1 U5948 ( .A1(n5477), .A2(n5476), .A3(n5475), .ZN(n4347) );
  NOR2_X1 U5949 ( .A1(n9313), .A2(n9328), .ZN(n4348) );
  AND2_X1 U5950 ( .A1(n4662), .A2(n4499), .ZN(n4349) );
  NAND2_X1 U5951 ( .A1(n5572), .A2(n5574), .ZN(n4350) );
  INV_X1 U5952 ( .A(n8179), .ZN(n4389) );
  AND2_X1 U5953 ( .A1(n8221), .A2(n6555), .ZN(n4351) );
  AND2_X1 U5954 ( .A1(n9224), .A2(n9209), .ZN(n4352) );
  AND2_X1 U5955 ( .A1(n6122), .A2(n4638), .ZN(n4353) );
  AND2_X1 U5956 ( .A1(n5692), .A2(n5691), .ZN(n4354) );
  INV_X1 U5957 ( .A(n5494), .ZN(n4671) );
  AND2_X1 U5958 ( .A1(n4933), .A2(SI_7_), .ZN(n4355) );
  NAND2_X1 U5959 ( .A1(n5373), .A2(n5372), .ZN(n8905) );
  INV_X1 U5960 ( .A(n8905), .ZN(n4501) );
  AND4_X1 U5961 ( .A1(n5054), .A2(n5053), .A3(n5052), .A4(n5051), .ZN(n7676)
         );
  NOR2_X1 U5962 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4356) );
  INV_X1 U5963 ( .A(n9090), .ZN(n4445) );
  INV_X2 U5964 ( .A(n5944), .ZN(n5941) );
  INV_X1 U5965 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4528) );
  NAND2_X1 U5966 ( .A1(n8637), .A2(n9740), .ZN(n8323) );
  NAND2_X1 U5967 ( .A1(n9239), .A2(n4619), .ZN(n4357) );
  OR2_X1 U5968 ( .A1(n4329), .A2(n4611), .ZN(n4358) );
  INV_X1 U5969 ( .A(n7936), .ZN(n4715) );
  AND3_X1 U5970 ( .A1(n5562), .A2(n5563), .A3(n5560), .ZN(n4359) );
  NOR2_X1 U5971 ( .A1(n4968), .A2(n4967), .ZN(n4360) );
  AND2_X1 U5972 ( .A1(n4356), .A2(n4314), .ZN(n4361) );
  INV_X1 U5973 ( .A(n5930), .ZN(n5938) );
  INV_X1 U5974 ( .A(n4650), .ZN(n4647) );
  NOR2_X1 U5975 ( .A1(n8288), .A2(n4651), .ZN(n4650) );
  NOR2_X1 U5976 ( .A1(n4831), .A2(n8992), .ZN(n4828) );
  INV_X1 U5977 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5815) );
  AND2_X1 U5978 ( .A1(n4326), .A2(n8405), .ZN(n4362) );
  NAND2_X1 U5979 ( .A1(n7650), .A2(n8262), .ZN(n6893) );
  INV_X1 U5980 ( .A(n8984), .ZN(n4812) );
  NAND2_X1 U5981 ( .A1(n5526), .A2(n4888), .ZN(n5529) );
  INV_X1 U5982 ( .A(n7966), .ZN(n4706) );
  NOR2_X1 U5983 ( .A1(n9193), .A2(n9208), .ZN(n4363) );
  NAND2_X1 U5984 ( .A1(n8531), .A2(n8530), .ZN(n4364) );
  NAND2_X1 U5985 ( .A1(n5561), .A2(n5560), .ZN(n5576) );
  INV_X1 U5986 ( .A(n5318), .ZN(n4551) );
  INV_X1 U5987 ( .A(n7684), .ZN(n5923) );
  INV_X1 U5988 ( .A(n8140), .ZN(n4699) );
  NAND2_X1 U5989 ( .A1(n7168), .A2(n8378), .ZN(n7260) );
  NAND2_X1 U5990 ( .A1(n7595), .A2(n7594), .ZN(n9453) );
  INV_X1 U5991 ( .A(n9453), .ZN(n4517) );
  OR2_X1 U5992 ( .A1(n8427), .A2(n8435), .ZN(n4365) );
  INV_X1 U5993 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4464) );
  INV_X1 U5994 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U5995 ( .A1(n5434), .A2(n5433), .ZN(n8883) );
  INV_X1 U5996 ( .A(n8883), .ZN(n4547) );
  INV_X1 U5997 ( .A(n9106), .ZN(n7831) );
  NAND2_X1 U5998 ( .A1(n7168), .A2(n4667), .ZN(n7319) );
  NOR3_X1 U5999 ( .A1(n9363), .A2(n9436), .A3(n4514), .ZN(n4512) );
  NOR2_X1 U6000 ( .A1(n7209), .A2(n7372), .ZN(n4366) );
  OR2_X1 U6001 ( .A1(n9537), .A2(n7467), .ZN(n4367) );
  NOR2_X1 U6002 ( .A1(n8382), .A2(n8187), .ZN(n4368) );
  NAND2_X1 U6003 ( .A1(n7174), .A2(n4309), .ZN(n4553) );
  INV_X1 U6004 ( .A(n4513), .ZN(n9332) );
  NOR2_X1 U6005 ( .A1(n9363), .A2(n4514), .ZN(n4513) );
  OR2_X1 U6006 ( .A1(n8898), .A2(n8586), .ZN(n8419) );
  INV_X1 U6007 ( .A(n9226), .ZN(n9096) );
  NAND2_X1 U6008 ( .A1(n7742), .A2(n7741), .ZN(n9226) );
  INV_X1 U6009 ( .A(n4538), .ZN(n8863) );
  NOR2_X1 U6010 ( .A1(n7616), .A2(n5344), .ZN(n4538) );
  OR2_X1 U6011 ( .A1(n5033), .A2(n5032), .ZN(n8624) );
  AND2_X1 U6012 ( .A1(n4551), .A2(n7565), .ZN(n4369) );
  INV_X1 U6013 ( .A(n8152), .ZN(n4687) );
  OR2_X1 U6014 ( .A1(n9411), .A2(n9250), .ZN(n8152) );
  NOR2_X1 U6015 ( .A1(n5036), .A2(n4889), .ZN(n4370) );
  OR2_X1 U6016 ( .A1(n4437), .A2(n4436), .ZN(n4371) );
  AND2_X1 U6017 ( .A1(n5586), .A2(n4335), .ZN(n5900) );
  NAND2_X1 U6018 ( .A1(n6396), .A2(n5160), .ZN(n4461) );
  OAI211_X1 U6019 ( .C1(n4721), .C2(n4720), .A(n4719), .B(n8224), .ZN(n6635)
         );
  OR2_X1 U6020 ( .A1(n9719), .A2(n4631), .ZN(n4372) );
  NAND2_X1 U6021 ( .A1(n5102), .A2(n5101), .ZN(n6553) );
  NAND2_X1 U6022 ( .A1(n4642), .A2(n8321), .ZN(n6362) );
  INV_X1 U6023 ( .A(n7600), .ZN(n4821) );
  XNOR2_X1 U6024 ( .A(n5885), .B(n5886), .ZN(n5899) );
  INV_X1 U6025 ( .A(n9659), .ZN(n7311) );
  AND2_X1 U6026 ( .A1(n6154), .A2(n6176), .ZN(n9659) );
  NAND2_X1 U6027 ( .A1(n5485), .A2(n8307), .ZN(n6543) );
  NAND2_X1 U6028 ( .A1(n4439), .A2(n7094), .ZN(n7095) );
  NAND2_X1 U6029 ( .A1(n4392), .A2(n6636), .ZN(n6626) );
  AND2_X1 U6030 ( .A1(n4710), .A2(n5561), .ZN(n5572) );
  INV_X1 U6031 ( .A(n6636), .ZN(n4396) );
  INV_X1 U6032 ( .A(n9802), .ZN(n4549) );
  XNOR2_X1 U6033 ( .A(n5473), .B(n5475), .ZN(n8282) );
  INV_X1 U6034 ( .A(n8727), .ZN(n4656) );
  NAND2_X1 U6035 ( .A1(n5927), .A2(n5926), .ZN(n7685) );
  NOR2_X1 U6036 ( .A1(n8707), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4373) );
  INV_X1 U6037 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n4536) );
  AND2_X1 U6038 ( .A1(n8454), .A2(n7547), .ZN(n8450) );
  INV_X1 U6039 ( .A(n8450), .ZN(n4717) );
  INV_X1 U6040 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n4468) );
  INV_X1 U6041 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n4681) );
  INV_X1 U6042 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n4677) );
  AND2_X2 U6043 ( .A1(n8453), .A2(n9763), .ZN(n9772) );
  NAND2_X1 U6044 ( .A1(n9744), .A2(n8282), .ZN(n8453) );
  NAND2_X2 U6045 ( .A1(n5061), .A2(n5060), .ZN(n4374) );
  NAND2_X1 U6046 ( .A1(n6205), .A2(n6770), .ZN(n6450) );
  NAND2_X1 U6047 ( .A1(n4374), .A2(n9762), .ZN(n6219) );
  XNOR2_X1 U6048 ( .A(n4374), .B(n5614), .ZN(n5597) );
  NAND2_X1 U6049 ( .A1(n8583), .A2(n4374), .ZN(n6254) );
  NOR2_X2 U6050 ( .A1(n8758), .A2(n5507), .ZN(n8745) );
  NAND3_X1 U6051 ( .A1(n5519), .A2(n7709), .A3(n5518), .ZN(n8877) );
  NAND2_X1 U6052 ( .A1(n4540), .A2(n5036), .ZN(n5534) );
  OR2_X1 U6053 ( .A1(n8178), .A2(n4330), .ZN(n4384) );
  NAND2_X1 U6054 ( .A1(n4384), .A2(n4385), .ZN(n8180) );
  XNOR2_X1 U6055 ( .A(n8180), .B(n8181), .ZN(n8589) );
  NAND3_X1 U6056 ( .A1(n4406), .A2(n4405), .A3(n8604), .ZN(n8215) );
  NAND3_X1 U6057 ( .A1(n7981), .A2(n8025), .A3(n8140), .ZN(n4424) );
  NAND4_X1 U6058 ( .A1(n4430), .A2(n8094), .A3(n8088), .A4(n4429), .ZN(n4428)
         );
  NAND3_X1 U6059 ( .A1(n4438), .A2(n7486), .A3(n4437), .ZN(n7519) );
  NAND3_X1 U6060 ( .A1(n4438), .A2(n7486), .A3(n4371), .ZN(n4435) );
  NAND3_X1 U6061 ( .A1(n4440), .A2(n4828), .A3(n9078), .ZN(n4824) );
  INV_X1 U6062 ( .A(n8993), .ZN(n4836) );
  NAND2_X1 U6063 ( .A1(n4794), .A2(n4795), .ZN(n4446) );
  NAND2_X1 U6064 ( .A1(n4441), .A2(n4442), .ZN(n9000) );
  NAND3_X1 U6065 ( .A1(n4794), .A2(n4795), .A3(n9090), .ZN(n4441) );
  NAND2_X1 U6066 ( .A1(n4446), .A2(n4801), .ZN(n9091) );
  NAND3_X1 U6067 ( .A1(n6658), .A2(n6714), .A3(n6657), .ZN(n6843) );
  INV_X1 U6068 ( .A(n6291), .ZN(n4448) );
  AND2_X1 U6069 ( .A1(n5072), .A2(n5071), .ZN(n6441) );
  OAI21_X1 U6070 ( .B1(n5102), .B2(n4451), .A(n4449), .ZN(n6357) );
  NAND2_X1 U6071 ( .A1(n8737), .A2(n8744), .ZN(n5455) );
  NAND3_X1 U6072 ( .A1(n5159), .A2(n4460), .A3(n4461), .ZN(n6560) );
  NAND3_X1 U6073 ( .A1(n5159), .A2(n4461), .A3(n5161), .ZN(n6561) );
  AND2_X1 U6074 ( .A1(n4361), .A2(n4887), .ZN(n4463) );
  NAND2_X1 U6075 ( .A1(n4462), .A2(n5036), .ZN(n4465) );
  AND3_X1 U6076 ( .A1(n4361), .A2(n4464), .A3(n4887), .ZN(n4462) );
  NOR2_X2 U6077 ( .A1(n4894), .A2(n7500), .ZN(n4469) );
  NAND2_X1 U6078 ( .A1(n4469), .A2(n4468), .ZN(n5089) );
  NAND2_X1 U6079 ( .A1(n4469), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U6080 ( .A1(n4469), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6081 ( .A1(n8358), .A2(n4479), .ZN(n8365) );
  OAI21_X1 U6082 ( .B1(n8392), .B2(n4484), .A(n4481), .ZN(n4489) );
  NAND2_X1 U6083 ( .A1(n8392), .A2(n8393), .ZN(n8403) );
  NAND2_X1 U6084 ( .A1(n4489), .A2(n8406), .ZN(n8398) );
  AND2_X1 U6085 ( .A1(n8400), .A2(n8394), .ZN(n4490) );
  NOR2_X2 U6086 ( .A1(n5271), .A2(n4883), .ZN(n5036) );
  NAND4_X1 U6087 ( .A1(n5123), .A2(n4881), .A3(n4880), .A4(n4879), .ZN(n5271)
         );
  OAI211_X1 U6088 ( .C1(n8415), .C2(n8435), .A(n4498), .B(n8418), .ZN(n4497)
         );
  AOI21_X1 U6089 ( .B1(n4501), .B2(n4500), .A(n8442), .ZN(n4499) );
  INV_X1 U6090 ( .A(n8845), .ZN(n4500) );
  INV_X1 U6091 ( .A(n4506), .ZN(n7160) );
  INV_X1 U6092 ( .A(n4507), .ZN(n9190) );
  INV_X2 U6093 ( .A(n5726), .ZN(n5561) );
  INV_X1 U6094 ( .A(n4512), .ZN(n9309) );
  NAND3_X1 U6095 ( .A1(n6499), .A2(n4519), .A3(n6692), .ZN(n6786) );
  INV_X1 U6096 ( .A(n7841), .ZN(n6012) );
  AND3_X2 U6097 ( .A1(n5947), .A2(n5948), .A3(n5946), .ZN(n7841) );
  NOR2_X1 U6098 ( .A1(n9599), .A2(n9598), .ZN(n9597) );
  NAND2_X1 U6099 ( .A1(n5849), .A2(n5850), .ZN(n5862) );
  MUX2_X1 U6100 ( .A(n5846), .B(P1_REG2_REG_3__SCAN_IN), .S(n5861), .Z(n5847)
         );
  NAND2_X1 U6101 ( .A1(n5036), .A2(n4539), .ZN(n4541) );
  AND2_X1 U6102 ( .A1(n4887), .A2(n4314), .ZN(n4540) );
  NOR2_X1 U6103 ( .A1(n8754), .A2(n4543), .ZN(n8730) );
  NOR2_X1 U6104 ( .A1(n8754), .A2(n8883), .ZN(n8755) );
  NAND3_X1 U6105 ( .A1(n4548), .A2(n4311), .A3(n6403), .ZN(n7663) );
  NAND3_X1 U6106 ( .A1(n6403), .A2(n4311), .A3(n4549), .ZN(n6828) );
  NAND2_X1 U6107 ( .A1(n7174), .A2(n4550), .ZN(n7558) );
  INV_X1 U6108 ( .A(n4553), .ZN(n7557) );
  MUX2_X1 U6109 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n5751), .S(n5764), .Z(n9498)
         );
  MUX2_X1 U6110 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5024), .Z(n5055) );
  NAND2_X1 U6111 ( .A1(n4940), .A2(n4768), .ZN(n4767) );
  NAND2_X1 U6112 ( .A1(n4341), .A2(n5137), .ZN(n4572) );
  NAND2_X1 U6113 ( .A1(n5394), .A2(n4576), .ZN(n4575) );
  INV_X1 U6114 ( .A(n5209), .ZN(n4586) );
  OAI21_X1 U6115 ( .B1(n5209), .B2(n4957), .A(n4956), .ZN(n5245) );
  NAND2_X1 U6116 ( .A1(n4360), .A2(n4956), .ZN(n4585) );
  OAI21_X1 U6117 ( .B1(n5035), .B2(n4589), .A(n4587), .ZN(n5337) );
  OAI21_X1 U6118 ( .B1(n5006), .B2(n4596), .A(n4593), .ZN(n5390) );
  NAND2_X1 U6119 ( .A1(n5006), .A2(n5345), .ZN(n4599) );
  NAND2_X1 U6120 ( .A1(n4953), .A2(n4952), .ZN(n5209) );
  NAND2_X1 U6121 ( .A1(n5443), .A2(n5442), .ZN(n5457) );
  NOR2_X1 U6122 ( .A1(n6351), .A2(n6352), .ZN(n6592) );
  MUX2_X1 U6123 ( .A(n5844), .B(P1_REG2_REG_1__SCAN_IN), .S(n5939), .Z(n9574)
         );
  AOI21_X1 U6124 ( .B1(n9172), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9165), .ZN(
        n9673) );
  XNOR2_X2 U6125 ( .A(n4527), .B(n5676), .ZN(n5939) );
  NAND2_X1 U6126 ( .A1(n4918), .A2(n4917), .ZN(n5108) );
  NAND2_X1 U6127 ( .A1(n4767), .A2(n4771), .ZN(n4953) );
  NAND2_X1 U6128 ( .A1(n9340), .A2(n4603), .ZN(n4601) );
  NAND2_X1 U6129 ( .A1(n9187), .A2(n4628), .ZN(n4627) );
  OAI21_X1 U6130 ( .B1(n9395), .B2(n4630), .A(n4625), .ZN(P1_U3520) );
  OAI211_X2 U6131 ( .C1(n9187), .C2(n8055), .A(n4629), .B(n4627), .ZN(n9395)
         );
  OAI21_X1 U6132 ( .B1(n9395), .B2(n9468), .A(n4632), .ZN(n9471) );
  AOI21_X2 U6133 ( .B1(n4637), .B2(n4636), .A(n4635), .ZN(n7454) );
  NAND2_X1 U6134 ( .A1(n7832), .A2(n9106), .ZN(n4636) );
  NAND3_X1 U6135 ( .A1(n6613), .A2(n6612), .A3(n8037), .ZN(n6680) );
  INV_X1 U6136 ( .A(n6683), .ZN(n6682) );
  INV_X1 U6137 ( .A(n4760), .ZN(n4641) );
  OAI211_X1 U6138 ( .C1(n4761), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n4640), .B(
        n4639), .ZN(n4911) );
  NAND3_X1 U6139 ( .A1(n4761), .A2(n4760), .A3(n5989), .ZN(n4639) );
  NAND2_X1 U6140 ( .A1(n5090), .A2(n4334), .ZN(n8639) );
  NAND2_X1 U6141 ( .A1(n6543), .A2(n8297), .ZN(n6550) );
  INV_X1 U6142 ( .A(n8297), .ZN(n4643) );
  INV_X1 U6143 ( .A(n4644), .ZN(n8242) );
  AOI21_X1 U6144 ( .B1(n8745), .B2(n4650), .A(n4645), .ZN(n4644) );
  INV_X1 U6145 ( .A(n4673), .ZN(n8853) );
  OR2_X1 U6146 ( .A1(n4680), .A2(n4677), .ZN(n4676) );
  NAND3_X1 U6147 ( .A1(n9491), .A2(n5707), .A3(P1_REG1_REG_1__SCAN_IN), .ZN(
        n4679) );
  XNOR2_X2 U6148 ( .A(n7841), .B(n9120), .ZN(n6158) );
  NAND2_X1 U6149 ( .A1(n9238), .A2(n8151), .ZN(n4686) );
  OAI21_X1 U6150 ( .B1(n7141), .B2(n4690), .A(n4688), .ZN(n7342) );
  OAI21_X1 U6151 ( .B1(n7465), .B2(n4707), .A(n4704), .ZN(n9375) );
  OAI21_X1 U6152 ( .B1(n7465), .B2(n8047), .A(n7966), .ZN(n8136) );
  NAND3_X1 U6153 ( .A1(n4710), .A2(n5561), .A3(n4847), .ZN(n5693) );
  NAND2_X1 U6154 ( .A1(n6675), .A2(n4713), .ZN(n4712) );
  XNOR2_X1 U6155 ( .A(n5598), .B(n5597), .ZN(n6250) );
  NAND3_X1 U6156 ( .A1(n5609), .A2(n5647), .A3(n5613), .ZN(n4719) );
  NAND2_X1 U6157 ( .A1(n4724), .A2(n4722), .ZN(n7379) );
  NAND2_X1 U6158 ( .A1(n6886), .A2(n4328), .ZN(n4724) );
  NAND2_X1 U6159 ( .A1(n6983), .A2(n4726), .ZN(n4725) );
  INV_X1 U6160 ( .A(n6983), .ZN(n4727) );
  NAND2_X1 U6161 ( .A1(n4728), .A2(n4731), .ZN(n8178) );
  NAND2_X1 U6162 ( .A1(n7629), .A2(n4729), .ZN(n4728) );
  NAND2_X1 U6163 ( .A1(n8575), .A2(n4742), .ZN(n4741) );
  NAND2_X1 U6164 ( .A1(n8575), .A2(n4750), .ZN(n4749) );
  NAND2_X1 U6165 ( .A1(n8575), .A2(n4744), .ZN(n4743) );
  NAND2_X1 U6166 ( .A1(n6796), .A2(n4751), .ZN(n6761) );
  NAND2_X1 U6167 ( .A1(n6761), .A2(n6760), .ZN(n6763) );
  NAND2_X1 U6168 ( .A1(n7386), .A2(n4755), .ZN(n4754) );
  NAND2_X1 U6169 ( .A1(n4754), .A2(n7445), .ZN(n7388) );
  NAND3_X1 U6170 ( .A1(n7445), .A2(n7386), .A3(n7387), .ZN(n7695) );
  NAND3_X1 U6171 ( .A1(n4761), .A2(n4760), .A3(n4905), .ZN(n5897) );
  NAND2_X1 U6172 ( .A1(n7324), .A2(n4850), .ZN(n7502) );
  NAND2_X1 U6173 ( .A1(n5137), .A2(n5138), .ZN(n4764) );
  NAND2_X1 U6174 ( .A1(n4940), .A2(n4939), .ZN(n5181) );
  NOR2_X1 U6175 ( .A1(n7555), .A2(n4784), .ZN(n7540) );
  NAND2_X1 U6176 ( .A1(n8903), .A2(n4788), .ZN(n4787) );
  INV_X1 U6177 ( .A(n4793), .ZN(n8797) );
  NAND2_X1 U6178 ( .A1(n4322), .A2(n4798), .ZN(n4809) );
  NAND3_X1 U6179 ( .A1(n4800), .A2(n4813), .A3(n4799), .ZN(n9031) );
  NAND2_X1 U6180 ( .A1(n7529), .A2(n4818), .ZN(n4817) );
  OAI21_X1 U6181 ( .B1(n7529), .B2(n4821), .A(n4818), .ZN(n8470) );
  NAND2_X1 U6182 ( .A1(n7182), .A2(n4822), .ZN(n7431) );
  OAI21_X1 U6183 ( .B1(n8993), .B2(n4827), .A(n4825), .ZN(n8515) );
  NAND2_X1 U6184 ( .A1(n4838), .A2(n6650), .ZN(n6655) );
  NAND2_X1 U6185 ( .A1(n4841), .A2(n4839), .ZN(n5887) );
  INV_X1 U6186 ( .A(n5346), .ZN(n5006) );
  NAND2_X1 U6187 ( .A1(n4919), .A2(n6053), .ZN(n4920) );
  NAND2_X1 U6188 ( .A1(n5457), .A2(n5456), .ZN(n5461) );
  NAND2_X1 U6189 ( .A1(n5441), .A2(n5440), .ZN(n5443) );
  NOR2_X1 U6190 ( .A1(n8587), .A2(n8187), .ZN(n8601) );
  AND2_X1 U6191 ( .A1(n8282), .A2(n9763), .ZN(n9786) );
  INV_X1 U6192 ( .A(n8282), .ZN(n8448) );
  AOI21_X2 U6193 ( .B1(n7022), .B2(n7021), .A(n4851), .ZN(n7137) );
  INV_X1 U6194 ( .A(n5517), .ZN(n8454) );
  NAND2_X1 U6195 ( .A1(n4305), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5710) );
  OR2_X1 U6196 ( .A1(n9234), .A2(n7868), .ZN(n7767) );
  NAND2_X1 U6197 ( .A1(n5586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5583) );
  MUX2_X1 U6198 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9496), .S(n5944), .Z(n7684) );
  NAND2_X1 U6199 ( .A1(n5931), .A2(n6092), .ZN(n5926) );
  AND2_X1 U6200 ( .A1(n9002), .A2(n5931), .ZN(n5936) );
  OR2_X1 U6201 ( .A1(n6067), .A2(n5988), .ZN(n5991) );
  NAND2_X1 U6202 ( .A1(n5929), .A2(n5960), .ZN(n6001) );
  NAND2_X4 U6203 ( .A1(n5749), .A2(n5942), .ZN(n5097) );
  AOI21_X2 U6204 ( .B1(n5128), .B2(n4312), .A(n4854), .ZN(n6396) );
  AOI22_X1 U6205 ( .A1(n8835), .A2(n8843), .B1(n8860), .B2(n8842), .ZN(n8822)
         );
  INV_X1 U6206 ( .A(n8036), .ZN(n6681) );
  NOR2_X1 U6207 ( .A1(n5492), .A2(n5491), .ZN(n4848) );
  NAND2_X1 U6208 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n4849) );
  NOR2_X1 U6209 ( .A1(n7020), .A2(n7019), .ZN(n4851) );
  OR2_X1 U6210 ( .A1(n4501), .A2(n8845), .ZN(n4852) );
  AND2_X1 U6211 ( .A1(n8743), .A2(n8615), .ZN(n4853) );
  NOR2_X1 U6212 ( .A1(n8256), .A2(n9740), .ZN(n4854) );
  AND4_X1 U6213 ( .A1(n5886), .A2(n10016), .A3(n6245), .A4(n5815), .ZN(n4855)
         );
  AND2_X1 U6214 ( .A1(n4952), .A2(n4951), .ZN(n4856) );
  INV_X1 U6215 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5481) );
  INV_X1 U6216 ( .A(n9493), .ZN(n7045) );
  INV_X1 U6217 ( .A(n7236), .ZN(n7159) );
  NAND2_X1 U6218 ( .A1(n6106), .A2(n6197), .ZN(n4859) );
  INV_X1 U6219 ( .A(n9772), .ZN(n9808) );
  INV_X1 U6220 ( .A(n8385), .ZN(n5317) );
  AND2_X2 U6221 ( .A1(n6218), .A2(n9742), .ZN(n9752) );
  INV_X2 U6222 ( .A(n9816), .ZN(n9817) );
  INV_X2 U6223 ( .A(n9828), .ZN(n9830) );
  INV_X2 U6224 ( .A(n9717), .ZN(n9719) );
  NAND2_X1 U6225 ( .A1(n6241), .A2(n9365), .ZN(n9367) );
  INV_X2 U6226 ( .A(n9724), .ZN(n9561) );
  NOR2_X1 U6227 ( .A1(n8270), .A2(n5498), .ZN(n5500) );
  OR4_X1 U6228 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n5879) );
  INV_X1 U6229 ( .A(n8376), .ZN(n5497) );
  NAND2_X1 U6230 ( .A1(n4882), .A2(n5273), .ZN(n4883) );
  AND2_X1 U6231 ( .A1(n6107), .A2(n6168), .ZN(n6099) );
  INV_X1 U6232 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5577) );
  INV_X1 U6233 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5278) );
  INV_X1 U6234 ( .A(n5630), .ZN(n5628) );
  INV_X1 U6235 ( .A(n7646), .ZN(n6757) );
  INV_X1 U6236 ( .A(n5358), .ZN(n4871) );
  INV_X1 U6237 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6238 ( .A1(n6217), .A2(n5070), .ZN(n5071) );
  NAND2_X1 U6239 ( .A1(n6107), .A2(n4859), .ZN(n6108) );
  INV_X1 U6240 ( .A(n7865), .ZN(n6325) );
  INV_X1 U6241 ( .A(n7149), .ZN(n6319) );
  INV_X1 U6242 ( .A(n5939), .ZN(n5940) );
  INV_X1 U6243 ( .A(n9218), .ZN(n8153) );
  OR2_X1 U6244 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  INV_X1 U6245 ( .A(n5417), .ZN(n5416) );
  OR2_X1 U6246 ( .A1(n5402), .A2(n5401), .ZN(n5417) );
  NAND2_X1 U6247 ( .A1(n4871), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5375) );
  INV_X1 U6248 ( .A(n7098), .ZN(n7096) );
  NAND2_X1 U6249 ( .A1(n6080), .A2(n6079), .ZN(n6081) );
  OR2_X1 U6250 ( .A1(n7867), .A2(n9033), .ZN(n7761) );
  NAND2_X1 U6251 ( .A1(n6325), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U6252 ( .A1(n6323), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U6253 ( .A1(n6318), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6928) );
  NAND2_X1 U6254 ( .A1(n7244), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5708) );
  INV_X1 U6255 ( .A(n6349), .ZN(n7024) );
  OR2_X1 U6256 ( .A1(n9436), .A2(n9302), .ZN(n8126) );
  NAND2_X1 U6257 ( .A1(n7035), .A2(n7142), .ZN(n7141) );
  NAND2_X1 U6258 ( .A1(n5941), .A2(n5940), .ZN(n5948) );
  NAND2_X1 U6259 ( .A1(n5426), .A2(n5425), .ZN(n5428) );
  NAND2_X1 U6260 ( .A1(n5337), .A2(n5336), .ZN(n5005) );
  NAND2_X1 U6261 ( .A1(n5416), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5446) );
  INV_X1 U6262 ( .A(n8640), .ZN(n5082) );
  NAND2_X1 U6263 ( .A1(n5339), .A2(n5338), .ZN(n5344) );
  OR2_X1 U6264 ( .A1(n5632), .A2(n8453), .ZN(n6888) );
  NAND2_X1 U6265 ( .A1(n4869), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5349) );
  INV_X1 U6266 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7227) );
  AND2_X1 U6267 ( .A1(n8400), .A2(n8404), .ZN(n8273) );
  INV_X1 U6268 ( .A(n7651), .ZN(n8261) );
  INV_X1 U6269 ( .A(n9757), .ZN(n5550) );
  INV_X1 U6270 ( .A(n8372), .ZN(n8268) );
  OR3_X1 U6271 ( .A1(n7077), .A2(n7365), .A3(n7273), .ZN(n5637) );
  NAND2_X1 U6272 ( .A1(n5474), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6273 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  INV_X1 U6274 ( .A(n6654), .ZN(n6653) );
  AND2_X1 U6275 ( .A1(n9056), .A2(n9057), .ZN(n9059) );
  OR2_X1 U6276 ( .A1(n7761), .A2(n9094), .ZN(n7887) );
  OR2_X1 U6277 ( .A1(n5965), .A2(n8107), .ZN(n5968) );
  AND2_X1 U6278 ( .A1(n7889), .A2(n7888), .ZN(n9191) );
  OR2_X1 U6279 ( .A1(n7792), .A2(n9025), .ZN(n7785) );
  INV_X1 U6280 ( .A(n9623), .ZN(n5848) );
  INV_X1 U6281 ( .A(n9287), .ZN(n9249) );
  INV_X1 U6282 ( .A(n9371), .ZN(n9330) );
  INV_X1 U6283 ( .A(n9105), .ZN(n7467) );
  OR2_X1 U6284 ( .A1(n8061), .A2(n5973), .ZN(n9329) );
  OR2_X1 U6285 ( .A1(n9696), .A2(n5967), .ZN(n9365) );
  INV_X1 U6286 ( .A(n7496), .ZN(n9537) );
  AND2_X1 U6287 ( .A1(n7918), .A2(n7920), .ZN(n6607) );
  OR2_X1 U6288 ( .A1(n8061), .A2(n5960), .ZN(n6131) );
  OR2_X1 U6289 ( .A1(n8016), .A2(n8104), .ZN(n9535) );
  AND2_X1 U6290 ( .A1(n5666), .A2(n5665), .ZN(n9690) );
  INV_X1 U6291 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5567) );
  OR2_X1 U6292 ( .A1(n5637), .A2(P2_U3152), .ZN(n5747) );
  INV_X1 U6293 ( .A(n9732), .ZN(n9727) );
  NAND2_X1 U6294 ( .A1(n8428), .A2(n8429), .ZN(n8759) );
  AND2_X1 U6295 ( .A1(n8407), .A2(n8405), .ZN(n7620) );
  AND2_X1 U6296 ( .A1(n8394), .A2(n8402), .ZN(n8272) );
  NAND2_X1 U6297 ( .A1(n4717), .A2(n8249), .ZN(n8817) );
  NAND2_X1 U6298 ( .A1(n5551), .A2(n5550), .ZN(n6369) );
  INV_X1 U6299 ( .A(n9800), .ZN(n9790) );
  OR3_X1 U6300 ( .A1(n9744), .A2(n8448), .A3(n8454), .ZN(n9778) );
  NAND2_X1 U6301 ( .A1(n7660), .A2(n9778), .ZN(n9800) );
  AND2_X1 U6302 ( .A1(n5536), .A2(n5535), .ZN(n9753) );
  AND2_X1 U6303 ( .A1(n5275), .A2(n5287), .ZN(n7407) );
  AND2_X1 U6304 ( .A1(n5942), .A2(P2_U3152), .ZN(n6150) );
  INV_X1 U6305 ( .A(n9095), .ZN(n9073) );
  AND2_X1 U6306 ( .A1(n5848), .A2(n5973), .ZN(n9676) );
  INV_X1 U6307 ( .A(n9686), .ZN(n9579) );
  INV_X1 U6308 ( .A(n9671), .ZN(n9685) );
  AND2_X1 U6309 ( .A1(n8108), .A2(n6095), .ZN(n6422) );
  INV_X1 U6310 ( .A(n7354), .ZN(n7158) );
  INV_X1 U6311 ( .A(n7363), .ZN(n7165) );
  INV_X1 U6312 ( .A(n9367), .ZN(n9356) );
  NOR2_X1 U6313 ( .A1(n5893), .A2(n9693), .ZN(n5894) );
  AND2_X1 U6314 ( .A1(n7354), .A2(n9535), .ZN(n9468) );
  AND2_X1 U6315 ( .A1(n5906), .A2(n6131), .ZN(n6240) );
  AOI21_X1 U6316 ( .B1(n9690), .B2(n5669), .A(n5667), .ZN(n6238) );
  INV_X1 U6317 ( .A(n5736), .ZN(n5973) );
  INV_X1 U6318 ( .A(n8724), .ZN(n9729) );
  OR3_X1 U6319 ( .A1(n8564), .A2(n8563), .A3(n8587), .ZN(n8565) );
  INV_X1 U6320 ( .A(n8898), .ZN(n8805) );
  INV_X1 U6321 ( .A(n8889), .ZN(n8781) );
  AND2_X1 U6322 ( .A1(n5382), .A2(n5381), .ZN(n8845) );
  OR2_X1 U6323 ( .A1(n5747), .A2(n5722), .ZN(n8620) );
  INV_X1 U6324 ( .A(n9728), .ZN(n9730) );
  OR2_X1 U6325 ( .A1(n8831), .A2(n9810), .ZN(n8736) );
  NAND2_X1 U6326 ( .A1(n8826), .A2(n6209), .ZN(n8869) );
  OR2_X1 U6327 ( .A1(n6370), .A2(n6369), .ZN(n9828) );
  NOR2_X1 U6328 ( .A1(n9754), .A2(n9753), .ZN(n9755) );
  INV_X1 U6329 ( .A(n9755), .ZN(n9758) );
  NAND2_X1 U6330 ( .A1(n5534), .A2(n5533), .ZN(n7365) );
  INV_X1 U6331 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6591) );
  INV_X1 U6332 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5730) );
  INV_X1 U6333 ( .A(n7043), .ZN(n8980) );
  NAND2_X1 U6334 ( .A1(n5974), .A2(n5736), .ZN(n9095) );
  INV_X1 U6335 ( .A(n9084), .ZN(n9102) );
  NAND2_X1 U6336 ( .A1(n7754), .A2(n7753), .ZN(n9240) );
  INV_X1 U6337 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9613) );
  INV_X1 U6338 ( .A(n9678), .ZN(n9592) );
  OR2_X1 U6339 ( .A1(P1_U3083), .A2(n5733), .ZN(n9671) );
  NAND2_X1 U6340 ( .A1(n9367), .A2(n6422), .ZN(n9383) );
  OR2_X1 U6341 ( .A1(n9319), .A2(n6273), .ZN(n7363) );
  NAND2_X1 U6342 ( .A1(n5907), .A2(n5894), .ZN(n9724) );
  NAND2_X1 U6343 ( .A1(n5907), .A2(n6240), .ZN(n9717) );
  AND2_X1 U6344 ( .A1(n9691), .A2(n9694), .ZN(n9692) );
  AND2_X1 U6345 ( .A1(n6132), .A2(n5663), .ZN(n9694) );
  INV_X1 U6346 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7734) );
  INV_X1 U6347 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7769) );
  INV_X1 U6348 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6248) );
  NOR2_X1 U6349 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  INV_X2 U6350 ( .A(n8620), .ZN(P2_U3966) );
  INV_X1 U6351 ( .A(n9119), .ZN(P1_U4006) );
  NAND2_X1 U6352 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5115) );
  INV_X1 U6353 ( .A(n5115), .ZN(n4860) );
  NAND2_X1 U6354 ( .A1(n4860), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5131) );
  INV_X1 U6355 ( .A(n5131), .ZN(n4861) );
  NAND2_X1 U6356 ( .A1(n4861), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5153) );
  INV_X1 U6357 ( .A(n5153), .ZN(n4862) );
  NAND2_X1 U6358 ( .A1(n4862), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5174) );
  INV_X1 U6359 ( .A(n5187), .ZN(n4863) );
  NAND2_X1 U6360 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n4864) );
  NAND2_X1 U6361 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n4868) );
  NAND2_X1 U6362 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n4870) );
  INV_X1 U6363 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5374) );
  INV_X1 U6364 ( .A(n5377), .ZN(n4872) );
  NAND2_X1 U6365 ( .A1(n4872), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5402) );
  INV_X1 U6366 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n4873) );
  NAND2_X1 U6367 ( .A1(n5377), .A2(n4873), .ZN(n4874) );
  NAND2_X1 U6368 ( .A1(n5402), .A2(n4874), .ZN(n8802) );
  AND4_X2 U6369 ( .A1(n5166), .A2(n5225), .A3(n4877), .A4(n5224), .ZN(n4881)
         );
  NOR2_X1 U6371 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n4884) );
  NAND4_X1 U6372 ( .A1(n4884), .A2(n5477), .A3(n5038), .A4(n5522), .ZN(n4886)
         );
  NAND4_X1 U6373 ( .A1(n5475), .A2(n5037), .A3(n5476), .A4(n5478), .ZN(n4885)
         );
  NOR2_X1 U6374 ( .A1(n4886), .A2(n4885), .ZN(n4887) );
  OR2_X1 U6375 ( .A1(n8802), .A2(n5419), .ZN(n4901) );
  NAND2_X2 U6376 ( .A1(n7500), .A2(n4893), .ZN(n5117) );
  INV_X1 U6377 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n4898) );
  NAND2_X1 U6378 ( .A1(n8237), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n4897) );
  NAND2_X1 U6379 ( .A1(n5086), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n4896) );
  OAI211_X1 U6380 ( .C1(n8240), .C2(n4898), .A(n4897), .B(n4896), .ZN(n4899)
         );
  INV_X1 U6381 ( .A(n4899), .ZN(n4900) );
  INV_X1 U6382 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4904) );
  AND2_X1 U6383 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4905) );
  NAND3_X1 U6384 ( .A1(n5024), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4906) );
  INV_X1 U6385 ( .A(SI_1_), .ZN(n4907) );
  NAND2_X1 U6386 ( .A1(n5056), .A2(n5055), .ZN(n4910) );
  NAND2_X1 U6387 ( .A1(n4908), .A2(SI_1_), .ZN(n4909) );
  NAND2_X1 U6388 ( .A1(n4910), .A2(n4909), .ZN(n5078) );
  INV_X1 U6389 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5657) );
  INV_X1 U6390 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5989) );
  XNOR2_X1 U6391 ( .A(n4911), .B(SI_2_), .ZN(n5079) );
  NAND2_X1 U6392 ( .A1(n5078), .A2(n5079), .ZN(n4914) );
  INV_X1 U6393 ( .A(n4911), .ZN(n4912) );
  NAND2_X1 U6394 ( .A1(n4912), .A2(SI_2_), .ZN(n4913) );
  NAND2_X1 U6395 ( .A1(n4914), .A2(n4913), .ZN(n5095) );
  INV_X1 U6396 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5658) );
  INV_X1 U6397 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6088) );
  MUX2_X1 U6398 ( .A(n5658), .B(n6088), .S(n4919), .Z(n4915) );
  XNOR2_X1 U6399 ( .A(n4915), .B(SI_3_), .ZN(n5096) );
  NAND2_X1 U6400 ( .A1(n5095), .A2(n5096), .ZN(n4918) );
  INV_X1 U6401 ( .A(n4915), .ZN(n4916) );
  NAND2_X1 U6402 ( .A1(n4916), .A2(SI_3_), .ZN(n4917) );
  INV_X1 U6403 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5659) );
  INV_X1 U6404 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6053) );
  XNOR2_X1 U6405 ( .A(n4921), .B(SI_4_), .ZN(n5109) );
  NAND2_X1 U6406 ( .A1(n5108), .A2(n5109), .ZN(n4924) );
  INV_X1 U6407 ( .A(n4921), .ZN(n4922) );
  NAND2_X1 U6408 ( .A1(n4922), .A2(SI_4_), .ZN(n4923) );
  INV_X1 U6409 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5670) );
  INV_X1 U6410 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6069) );
  MUX2_X1 U6411 ( .A(n5670), .B(n6069), .S(n5942), .Z(n4925) );
  XNOR2_X1 U6412 ( .A(n4925), .B(SI_5_), .ZN(n5124) );
  NAND2_X1 U6413 ( .A1(n5125), .A2(n5124), .ZN(n4928) );
  INV_X1 U6414 ( .A(n4925), .ZN(n4926) );
  NAND2_X1 U6415 ( .A1(n4926), .A2(SI_5_), .ZN(n4927) );
  INV_X1 U6416 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5671) );
  INV_X1 U6417 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6121) );
  MUX2_X1 U6418 ( .A(n5671), .B(n6121), .S(n5942), .Z(n4929) );
  XNOR2_X1 U6419 ( .A(n4929), .B(SI_6_), .ZN(n5138) );
  INV_X1 U6420 ( .A(n4929), .ZN(n4930) );
  NAND2_X1 U6421 ( .A1(n4930), .A2(SI_6_), .ZN(n4931) );
  INV_X1 U6422 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5684) );
  INV_X1 U6423 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6288) );
  MUX2_X1 U6424 ( .A(n5684), .B(n6288), .S(n5942), .Z(n4932) );
  XNOR2_X1 U6425 ( .A(n4932), .B(SI_7_), .ZN(n5145) );
  INV_X1 U6426 ( .A(n4932), .ZN(n4933) );
  INV_X1 U6427 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5690) );
  INV_X1 U6428 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n4934) );
  MUX2_X1 U6429 ( .A(n5690), .B(n4934), .S(n5942), .Z(n4936) );
  INV_X1 U6430 ( .A(SI_8_), .ZN(n4935) );
  NAND2_X1 U6431 ( .A1(n4936), .A2(n4935), .ZN(n4939) );
  INV_X1 U6432 ( .A(n4936), .ZN(n4937) );
  NAND2_X1 U6433 ( .A1(n4937), .A2(SI_8_), .ZN(n4938) );
  NAND2_X1 U6434 ( .A1(n4939), .A2(n4938), .ZN(n5162) );
  INV_X1 U6435 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4941) );
  MUX2_X1 U6436 ( .A(n5720), .B(n4941), .S(n5942), .Z(n4943) );
  INV_X1 U6437 ( .A(SI_9_), .ZN(n4942) );
  NAND2_X1 U6438 ( .A1(n4943), .A2(n4942), .ZN(n4946) );
  INV_X1 U6439 ( .A(n4943), .ZN(n4944) );
  NAND2_X1 U6440 ( .A1(n4944), .A2(SI_9_), .ZN(n4945) );
  INV_X1 U6441 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4947) );
  MUX2_X1 U6442 ( .A(n5730), .B(n4947), .S(n5942), .Z(n4949) );
  INV_X1 U6443 ( .A(SI_10_), .ZN(n4948) );
  NAND2_X1 U6444 ( .A1(n4949), .A2(n4948), .ZN(n4952) );
  INV_X1 U6445 ( .A(n4949), .ZN(n4950) );
  NAND2_X1 U6446 ( .A1(n4950), .A2(SI_10_), .ZN(n4951) );
  MUX2_X1 U6447 ( .A(n5820), .B(n9865), .S(n5942), .Z(n4954) );
  XNOR2_X1 U6448 ( .A(n4954), .B(SI_11_), .ZN(n5208) );
  INV_X1 U6449 ( .A(n5208), .ZN(n4957) );
  INV_X1 U6450 ( .A(n4954), .ZN(n4955) );
  NAND2_X1 U6451 ( .A1(n4955), .A2(SI_11_), .ZN(n4956) );
  MUX2_X1 U6452 ( .A(n5984), .B(n5982), .S(n5942), .Z(n4959) );
  INV_X1 U6453 ( .A(SI_12_), .ZN(n4958) );
  NAND2_X1 U6454 ( .A1(n4959), .A2(n4958), .ZN(n5246) );
  INV_X1 U6455 ( .A(n4959), .ZN(n4960) );
  NAND2_X1 U6456 ( .A1(n4960), .A2(SI_12_), .ZN(n4961) );
  NAND2_X1 U6457 ( .A1(n5246), .A2(n4961), .ZN(n5244) );
  MUX2_X1 U6458 ( .A(n6181), .B(n6155), .S(n5942), .Z(n4965) );
  XNOR2_X1 U6459 ( .A(n4965), .B(SI_14_), .ZN(n5269) );
  INV_X1 U6460 ( .A(n5269), .ZN(n4964) );
  INV_X1 U6461 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6036) );
  INV_X1 U6462 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4962) );
  MUX2_X1 U6463 ( .A(n6036), .B(n4962), .S(n5942), .Z(n4970) );
  INV_X1 U6464 ( .A(n4970), .ZN(n4963) );
  NAND2_X1 U6465 ( .A1(n4963), .A2(SI_13_), .ZN(n5265) );
  NOR2_X1 U6466 ( .A1(n4964), .A2(n5265), .ZN(n4972) );
  OR2_X1 U6467 ( .A1(n5244), .A2(n4972), .ZN(n4968) );
  INV_X1 U6468 ( .A(n4965), .ZN(n4966) );
  NAND2_X1 U6469 ( .A1(n4966), .A2(SI_14_), .ZN(n4974) );
  INV_X1 U6470 ( .A(n4974), .ZN(n4967) );
  INV_X1 U6471 ( .A(SI_13_), .ZN(n4969) );
  NAND2_X1 U6472 ( .A1(n4970), .A2(n4969), .ZN(n5247) );
  AND2_X1 U6473 ( .A1(n5246), .A2(n5247), .ZN(n5267) );
  AND2_X1 U6474 ( .A1(n5267), .A2(n5269), .ZN(n4971) );
  NOR2_X1 U6475 ( .A1(n4972), .A2(n4971), .ZN(n4973) );
  INV_X1 U6476 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n4975) );
  MUX2_X1 U6477 ( .A(n4975), .B(n6180), .S(n5942), .Z(n4977) );
  INV_X1 U6478 ( .A(SI_15_), .ZN(n4976) );
  NAND2_X1 U6479 ( .A1(n4977), .A2(n4976), .ZN(n4980) );
  INV_X1 U6480 ( .A(n4977), .ZN(n4978) );
  NAND2_X1 U6481 ( .A1(n4978), .A2(SI_15_), .ZN(n4979) );
  NAND2_X1 U6482 ( .A1(n4980), .A2(n4979), .ZN(n5285) );
  MUX2_X1 U6483 ( .A(n9884), .B(n6248), .S(n5942), .Z(n4982) );
  NAND2_X1 U6484 ( .A1(n4982), .A2(n4981), .ZN(n4985) );
  INV_X1 U6485 ( .A(n4982), .ZN(n4983) );
  NAND2_X1 U6486 ( .A1(n4983), .A2(SI_16_), .ZN(n4984) );
  NAND2_X1 U6487 ( .A1(n5302), .A2(n5301), .ZN(n4986) );
  MUX2_X1 U6488 ( .A(n6271), .B(n4987), .S(n5942), .Z(n4988) );
  XNOR2_X1 U6489 ( .A(n4988), .B(SI_17_), .ZN(n5045) );
  INV_X1 U6490 ( .A(n5045), .ZN(n4991) );
  INV_X1 U6491 ( .A(n4988), .ZN(n4989) );
  NAND2_X1 U6492 ( .A1(n4989), .A2(SI_17_), .ZN(n4990) );
  MUX2_X1 U6493 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5942), .Z(n4993) );
  XNOR2_X1 U6494 ( .A(n4993), .B(SI_18_), .ZN(n5034) );
  INV_X1 U6495 ( .A(n5034), .ZN(n4992) );
  NAND2_X1 U6496 ( .A1(n4993), .A2(SI_18_), .ZN(n4994) );
  MUX2_X1 U6497 ( .A(n6591), .B(n6589), .S(n5942), .Z(n4996) );
  INV_X1 U6498 ( .A(SI_19_), .ZN(n4995) );
  NAND2_X1 U6499 ( .A1(n4996), .A2(n4995), .ZN(n4999) );
  INV_X1 U6500 ( .A(n4996), .ZN(n4997) );
  NAND2_X1 U6501 ( .A1(n4997), .A2(SI_19_), .ZN(n4998) );
  NAND2_X1 U6502 ( .A1(n4999), .A2(n4998), .ZN(n5319) );
  MUX2_X1 U6503 ( .A(n8207), .B(n7788), .S(n5942), .Z(n5001) );
  INV_X1 U6504 ( .A(SI_20_), .ZN(n5000) );
  NAND2_X1 U6505 ( .A1(n5001), .A2(n5000), .ZN(n5004) );
  INV_X1 U6506 ( .A(n5001), .ZN(n5002) );
  NAND2_X1 U6507 ( .A1(n5002), .A2(SI_20_), .ZN(n5003) );
  MUX2_X1 U6508 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5942), .Z(n5007) );
  XNOR2_X1 U6509 ( .A(n5007), .B(n9873), .ZN(n5345) );
  NAND2_X1 U6510 ( .A1(n5007), .A2(SI_21_), .ZN(n5008) );
  MUX2_X1 U6511 ( .A(n7006), .B(n7769), .S(n5942), .Z(n5010) );
  INV_X1 U6512 ( .A(SI_22_), .ZN(n5009) );
  NAND2_X1 U6513 ( .A1(n5010), .A2(n5009), .ZN(n5368) );
  INV_X1 U6514 ( .A(n5010), .ZN(n5011) );
  NAND2_X1 U6515 ( .A1(n5011), .A2(SI_22_), .ZN(n5012) );
  NAND2_X1 U6516 ( .A1(n5368), .A2(n5012), .ZN(n5366) );
  MUX2_X1 U6517 ( .A(n9886), .B(n7817), .S(n5942), .Z(n5016) );
  INV_X1 U6518 ( .A(n5016), .ZN(n5013) );
  NAND2_X1 U6519 ( .A1(n5013), .A2(SI_23_), .ZN(n5387) );
  INV_X1 U6520 ( .A(n5387), .ZN(n5017) );
  OR2_X1 U6521 ( .A1(n5366), .A2(n5017), .ZN(n5014) );
  OR2_X1 U6522 ( .A1(n5367), .A2(n5014), .ZN(n5019) );
  INV_X1 U6523 ( .A(SI_23_), .ZN(n5015) );
  NAND2_X1 U6524 ( .A1(n5016), .A2(n5015), .ZN(n5369) );
  AND2_X1 U6525 ( .A1(n5368), .A2(n5369), .ZN(n5383) );
  OR2_X1 U6526 ( .A1(n5017), .A2(n5383), .ZN(n5018) );
  NAND2_X1 U6527 ( .A1(n5019), .A2(n5018), .ZN(n5020) );
  MUX2_X1 U6528 ( .A(n7076), .B(n7862), .S(n5942), .Z(n5391) );
  NAND2_X4 U6529 ( .A1(n5508), .A2(n5509), .ZN(n5749) );
  NAND2_X1 U6531 ( .A1(n7861), .A2(n5464), .ZN(n5026) );
  OR2_X1 U6532 ( .A1(n5097), .A2(n7076), .ZN(n5025) );
  INV_X1 U6533 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5028) );
  INV_X1 U6534 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5027) );
  OAI21_X1 U6535 ( .B1(n5312), .B2(n5028), .A(n5027), .ZN(n5029) );
  NAND2_X1 U6536 ( .A1(n5029), .A2(n5330), .ZN(n7560) );
  INV_X1 U6537 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5030) );
  OAI22_X1 U6538 ( .A1(n7560), .A2(n5419), .B1(n5117), .B2(n5030), .ZN(n5033)
         );
  INV_X1 U6539 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U6540 ( .A1(n8237), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5031) );
  OAI21_X1 U6541 ( .B1(n5309), .B2(n8696), .A(n5031), .ZN(n5032) );
  INV_X1 U6542 ( .A(n8624), .ZN(n7394) );
  XNOR2_X1 U6543 ( .A(n5035), .B(n5034), .ZN(n7799) );
  NAND2_X1 U6544 ( .A1(n7799), .A2(n5464), .ZN(n5040) );
  XNOR2_X1 U6545 ( .A(n5321), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8707) );
  AOI22_X1 U6546 ( .A1(n5326), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5325), .B2(
        n8707), .ZN(n5039) );
  XNOR2_X1 U6547 ( .A(n5312), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n7393) );
  NAND2_X1 U6548 ( .A1(n7393), .A2(n4469), .ZN(n5044) );
  NAND2_X1 U6549 ( .A1(n5086), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6550 ( .A1(n8237), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5042) );
  INV_X1 U6551 ( .A(n8240), .ZN(n5351) );
  NAND2_X1 U6552 ( .A1(n5351), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5041) );
  NAND2_X1 U6553 ( .A1(n7593), .A2(n5464), .ZN(n5049) );
  OR2_X1 U6554 ( .A1(n5304), .A2(n4889), .ZN(n5047) );
  XNOR2_X1 U6555 ( .A(n5047), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8697) );
  AOI22_X1 U6556 ( .A1(n5326), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5325), .B2(
        n8697), .ZN(n5048) );
  INV_X1 U6557 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6215) );
  OR2_X1 U6558 ( .A1(n5117), .A2(n6215), .ZN(n5054) );
  INV_X1 U6559 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5050) );
  OR2_X1 U6560 ( .A1(n5215), .A2(n5050), .ZN(n5053) );
  INV_X1 U6561 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U6562 ( .A1(n5086), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5051) );
  XNOR2_X1 U6563 ( .A(n5056), .B(n5055), .ZN(n5943) );
  INV_X1 U6564 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6565 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5057) );
  OAI22_X1 U6566 ( .A1(n5147), .A2(n5943), .B1(n5749), .B2(n5764), .ZN(n5059)
         );
  INV_X1 U6567 ( .A(n5059), .ZN(n5061) );
  INV_X1 U6568 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5656) );
  OR2_X1 U6569 ( .A1(n5097), .A2(n5656), .ZN(n5060) );
  NAND2_X1 U6570 ( .A1(n6205), .A2(n7676), .ZN(n5070) );
  AND2_X1 U6571 ( .A1(n8315), .A2(n5070), .ZN(n5062) );
  NAND2_X1 U6572 ( .A1(n5062), .A2(n8313), .ZN(n5072) );
  INV_X1 U6573 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5063) );
  OR2_X1 U6574 ( .A1(n5215), .A2(n5063), .ZN(n5068) );
  NAND2_X1 U6575 ( .A1(n5086), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5067) );
  INV_X1 U6576 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6776) );
  INV_X1 U6577 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5064) );
  OR2_X1 U6578 ( .A1(n5117), .A2(n5064), .ZN(n5065) );
  NAND2_X1 U6579 ( .A1(n7725), .A2(SI_0_), .ZN(n5069) );
  XNOR2_X1 U6580 ( .A(n5069), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8981) );
  MUX2_X1 U6581 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8981), .S(n5749), .Z(n9762) );
  INV_X1 U6582 ( .A(n9762), .ZN(n6770) );
  INV_X1 U6583 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7677) );
  INV_X1 U6584 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5763) );
  OR2_X1 U6585 ( .A1(n5117), .A2(n5763), .ZN(n5076) );
  INV_X1 U6586 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U6587 ( .A1(n5086), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5074) );
  NAND4_X1 U6588 ( .A1(n5077), .A2(n5076), .A3(n5075), .A4(n5074), .ZN(n8640)
         );
  OAI21_X1 U6589 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(P2_IR_REG_0__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5092) );
  INV_X1 U6590 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9875) );
  XNOR2_X1 U6591 ( .A(n5092), .B(n9875), .ZN(n5765) );
  XNOR2_X1 U6592 ( .A(n5078), .B(n5079), .ZN(n5988) );
  OR2_X1 U6593 ( .A1(n5147), .A2(n5988), .ZN(n5081) );
  OAI211_X1 U6594 ( .C1(n5749), .C2(n5765), .A(n5081), .B(n5080), .ZN(n5516)
         );
  INV_X1 U6595 ( .A(n5516), .ZN(n5083) );
  NAND2_X1 U6596 ( .A1(n8640), .A2(n5083), .ZN(n8317) );
  NAND2_X1 U6597 ( .A1(n5082), .A2(n5516), .ZN(n8316) );
  INV_X1 U6598 ( .A(n8253), .ZN(n6443) );
  NAND2_X1 U6599 ( .A1(n5082), .A2(n5083), .ZN(n5084) );
  NAND2_X1 U6600 ( .A1(n5085), .A2(n5084), .ZN(n6536) );
  NAND2_X1 U6601 ( .A1(n5086), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5091) );
  INV_X1 U6602 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5087) );
  OR2_X1 U6603 ( .A1(n5215), .A2(n5087), .ZN(n5090) );
  INV_X1 U6604 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5762) );
  OR2_X1 U6605 ( .A1(n5117), .A2(n5762), .ZN(n5088) );
  NAND2_X1 U6606 ( .A1(n5092), .A2(n9875), .ZN(n5093) );
  NAND2_X1 U6607 ( .A1(n5093), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5094) );
  XNOR2_X1 U6608 ( .A(n5094), .B(P2_IR_REG_3__SCAN_IN), .ZN(n5761) );
  INV_X1 U6609 ( .A(n5761), .ZN(n5814) );
  XNOR2_X1 U6610 ( .A(n5096), .B(n5095), .ZN(n6087) );
  OR2_X1 U6611 ( .A1(n5147), .A2(n6087), .ZN(n5099) );
  OR2_X1 U6612 ( .A1(n5097), .A2(n5658), .ZN(n5098) );
  OAI211_X1 U6613 ( .C1(n5749), .C2(n5814), .A(n5099), .B(n5098), .ZN(n6542)
         );
  NAND2_X1 U6614 ( .A1(n5100), .A2(n6542), .ZN(n8297) );
  NAND2_X1 U6615 ( .A1(n6536), .A2(n8254), .ZN(n5102) );
  NAND2_X1 U6616 ( .A1(n5100), .A2(n9780), .ZN(n5101) );
  NAND2_X1 U6617 ( .A1(n5086), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5107) );
  INV_X1 U6618 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5103) );
  OR2_X1 U6619 ( .A1(n5215), .A2(n5103), .ZN(n5106) );
  OAI21_X1 U6620 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5115), .ZN(n6812) );
  OR2_X1 U6621 ( .A1(n5419), .A2(n6812), .ZN(n5105) );
  INV_X1 U6622 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5767) );
  OR2_X1 U6623 ( .A1(n8240), .A2(n5767), .ZN(n5104) );
  XNOR2_X1 U6624 ( .A(n5108), .B(n5109), .ZN(n6052) );
  OR2_X1 U6625 ( .A1(n5147), .A2(n6052), .ZN(n5113) );
  OR2_X1 U6626 ( .A1(n5097), .A2(n5659), .ZN(n5112) );
  OR2_X1 U6627 ( .A1(n5123), .A2(n4889), .ZN(n5110) );
  XNOR2_X1 U6628 ( .A(n5110), .B(n5122), .ZN(n5785) );
  OR2_X1 U6629 ( .A1(n5749), .A2(n5785), .ZN(n5111) );
  NOR2_X1 U6630 ( .A1(n8638), .A2(n6555), .ZN(n5486) );
  NAND2_X1 U6631 ( .A1(n8638), .A2(n6555), .ZN(n8321) );
  INV_X1 U6632 ( .A(n8638), .ZN(n8221) );
  NAND2_X1 U6633 ( .A1(n5086), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5121) );
  OR2_X1 U6634 ( .A1(n5215), .A2(n6368), .ZN(n5120) );
  INV_X1 U6635 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5114) );
  NAND2_X1 U6636 ( .A1(n5115), .A2(n5114), .ZN(n5116) );
  NAND2_X1 U6637 ( .A1(n5131), .A2(n5116), .ZN(n9741) );
  OR2_X1 U6638 ( .A1(n5419), .A2(n9741), .ZN(n5119) );
  INV_X1 U6639 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5783) );
  OR2_X1 U6640 ( .A1(n5117), .A2(n5783), .ZN(n5118) );
  NAND2_X1 U6641 ( .A1(n5123), .A2(n5122), .ZN(n5168) );
  NAND2_X1 U6642 ( .A1(n5168), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5139) );
  XNOR2_X1 U6643 ( .A(n5139), .B(P2_IR_REG_5__SCAN_IN), .ZN(n5782) );
  INV_X1 U6644 ( .A(n5782), .ZN(n5803) );
  OR2_X1 U6645 ( .A1(n6068), .A2(n5147), .ZN(n5127) );
  OR2_X1 U6646 ( .A1(n5097), .A2(n5670), .ZN(n5126) );
  OAI211_X1 U6647 ( .C1(n5749), .C2(n5803), .A(n5127), .B(n5126), .ZN(n8219)
         );
  INV_X1 U6648 ( .A(n8219), .ZN(n9740) );
  INV_X1 U6649 ( .A(n6632), .ZN(n8637) );
  NAND2_X1 U6650 ( .A1(n6632), .A2(n8219), .ZN(n8299) );
  NAND2_X1 U6651 ( .A1(n5086), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5136) );
  INV_X1 U6652 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5129) );
  OR2_X1 U6653 ( .A1(n5215), .A2(n5129), .ZN(n5135) );
  INV_X1 U6654 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6655 ( .A1(n5131), .A2(n5130), .ZN(n5132) );
  NAND2_X1 U6656 ( .A1(n5153), .A2(n5132), .ZN(n6627) );
  OR2_X1 U6657 ( .A1(n5419), .A2(n6627), .ZN(n5134) );
  INV_X1 U6658 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6402) );
  OR2_X1 U6659 ( .A1(n5117), .A2(n6402), .ZN(n5133) );
  INV_X1 U6660 ( .A(n8218), .ZN(n8636) );
  OR2_X1 U6661 ( .A1(n6119), .A2(n5147), .ZN(n5144) );
  NAND2_X1 U6662 ( .A1(n5139), .A2(n5166), .ZN(n5140) );
  NAND2_X1 U6663 ( .A1(n5140), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6664 ( .A1(n5141), .A2(n5165), .ZN(n5148) );
  OR2_X1 U6665 ( .A1(n5141), .A2(n5165), .ZN(n5142) );
  AOI22_X1 U6666 ( .A1(n5326), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5325), .B2(
        n5830), .ZN(n5143) );
  INV_X1 U6667 ( .A(n9794), .ZN(n6630) );
  NAND2_X1 U6668 ( .A1(n8636), .A2(n6630), .ZN(n6395) );
  XNOR2_X1 U6669 ( .A(n5146), .B(n5145), .ZN(n6287) );
  OR2_X1 U6670 ( .A1(n6287), .A2(n5147), .ZN(n5151) );
  NAND2_X1 U6671 ( .A1(n5148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5149) );
  XNOR2_X1 U6672 ( .A(n5149), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6184) );
  AOI22_X1 U6673 ( .A1(n5326), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5325), .B2(
        n6184), .ZN(n5150) );
  NAND2_X1 U6674 ( .A1(n5151), .A2(n5150), .ZN(n6479) );
  NAND2_X1 U6675 ( .A1(n5086), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5158) );
  INV_X1 U6676 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5152) );
  OR2_X1 U6677 ( .A1(n5215), .A2(n5152), .ZN(n5157) );
  INV_X1 U6678 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U6679 ( .A1(n5153), .A2(n5823), .ZN(n5154) );
  NAND2_X1 U6680 ( .A1(n5174), .A2(n5154), .ZN(n6508) );
  OR2_X1 U6681 ( .A1(n5419), .A2(n6508), .ZN(n5156) );
  INV_X1 U6682 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6507) );
  OR2_X1 U6683 ( .A1(n8240), .A2(n6507), .ZN(n5155) );
  OR2_X1 U6684 ( .A1(n6479), .A2(n6741), .ZN(n8344) );
  INV_X1 U6685 ( .A(n5487), .ZN(n8331) );
  INV_X1 U6686 ( .A(n8259), .ZN(n8329) );
  AND2_X1 U6687 ( .A1(n6395), .A2(n8329), .ZN(n5160) );
  NAND2_X1 U6688 ( .A1(n8218), .A2(n9794), .ZN(n6470) );
  OR2_X1 U6689 ( .A1(n8259), .A2(n6470), .ZN(n5159) );
  INV_X1 U6690 ( .A(n6741), .ZN(n8635) );
  OR2_X1 U6691 ( .A1(n8635), .A2(n6479), .ZN(n5161) );
  XNOR2_X1 U6692 ( .A(n5163), .B(n5162), .ZN(n6642) );
  NAND2_X1 U6693 ( .A1(n6642), .A2(n5464), .ZN(n5171) );
  NAND3_X1 U6694 ( .A1(n5166), .A2(n5165), .A3(n5164), .ZN(n5167) );
  NAND2_X1 U6695 ( .A1(n5182), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5169) );
  XNOR2_X1 U6696 ( .A(n5169), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6375) );
  AOI22_X1 U6697 ( .A1(n5326), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5325), .B2(
        n6375), .ZN(n5170) );
  NAND2_X1 U6698 ( .A1(n5171), .A2(n5170), .ZN(n9802) );
  NAND2_X1 U6699 ( .A1(n5086), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5179) );
  INV_X1 U6700 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5172) );
  OR2_X1 U6701 ( .A1(n5215), .A2(n5172), .ZN(n5178) );
  NAND2_X1 U6702 ( .A1(n5174), .A2(n5173), .ZN(n5175) );
  NAND2_X1 U6703 ( .A1(n5187), .A2(n5175), .ZN(n6740) );
  OR2_X1 U6704 ( .A1(n5419), .A2(n6740), .ZN(n5177) );
  INV_X1 U6705 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6566) );
  OR2_X1 U6706 ( .A1(n8240), .A2(n6566), .ZN(n5176) );
  OR2_X1 U6707 ( .A1(n9802), .A2(n6820), .ZN(n8342) );
  NAND2_X1 U6708 ( .A1(n9802), .A2(n6820), .ZN(n8347) );
  NAND2_X1 U6709 ( .A1(n8342), .A2(n8347), .ZN(n8346) );
  INV_X1 U6710 ( .A(n6820), .ZN(n8634) );
  NAND2_X1 U6711 ( .A1(n9802), .A2(n8634), .ZN(n5180) );
  NAND2_X1 U6712 ( .A1(n6706), .A2(n5464), .ZN(n5184) );
  NOR2_X1 U6713 ( .A1(n5182), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5228) );
  OR2_X1 U6714 ( .A1(n5228), .A2(n4889), .ZN(n5195) );
  XNOR2_X1 U6715 ( .A(n5195), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6580) );
  AOI22_X1 U6716 ( .A1(n5326), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5325), .B2(
        n6580), .ZN(n5183) );
  NAND2_X1 U6717 ( .A1(n5086), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5192) );
  INV_X1 U6718 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5185) );
  OR2_X1 U6719 ( .A1(n5215), .A2(n5185), .ZN(n5191) );
  INV_X1 U6720 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6721 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  NAND2_X1 U6722 ( .A1(n5218), .A2(n5188), .ZN(n6830) );
  OR2_X1 U6723 ( .A1(n5419), .A2(n6830), .ZN(n5190) );
  INV_X1 U6724 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6831) );
  OR2_X1 U6725 ( .A1(n8240), .A2(n6831), .ZN(n5189) );
  OR2_X1 U6726 ( .A1(n6975), .A2(n7655), .ZN(n8343) );
  NAND2_X1 U6727 ( .A1(n6975), .A2(n7655), .ZN(n8353) );
  NAND2_X1 U6728 ( .A1(n6818), .A2(n8261), .ZN(n6817) );
  INV_X1 U6729 ( .A(n7655), .ZN(n8633) );
  OR2_X1 U6730 ( .A1(n6975), .A2(n8633), .ZN(n5193) );
  XNOR2_X1 U6731 ( .A(n5194), .B(n4856), .ZN(n5725) );
  NAND2_X1 U6732 ( .A1(n5725), .A2(n5464), .ZN(n5201) );
  INV_X1 U6733 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6734 ( .A1(n5195), .A2(n5226), .ZN(n5196) );
  NAND2_X1 U6735 ( .A1(n5196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5198) );
  INV_X1 U6736 ( .A(n5198), .ZN(n5197) );
  NAND2_X1 U6737 ( .A1(n5197), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6738 ( .A1(n5198), .A2(n5225), .ZN(n5210) );
  AOI22_X1 U6739 ( .A1(n5326), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5325), .B2(
        n6963), .ZN(n5200) );
  NAND2_X1 U6740 ( .A1(n5086), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5206) );
  INV_X1 U6741 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5202) );
  OR2_X1 U6742 ( .A1(n5215), .A2(n5202), .ZN(n5205) );
  INV_X1 U6743 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5217) );
  XNOR2_X1 U6744 ( .A(n5218), .B(n5217), .ZN(n7661) );
  OR2_X1 U6745 ( .A1(n5419), .A2(n7661), .ZN(n5204) );
  INV_X1 U6746 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7662) );
  OR2_X1 U6747 ( .A1(n5117), .A2(n7662), .ZN(n5203) );
  NAND2_X1 U6748 ( .A1(n8337), .A2(n8294), .ZN(n8262) );
  INV_X1 U6749 ( .A(n6819), .ZN(n8632) );
  NAND2_X1 U6750 ( .A1(n5207), .A2(n8632), .ZN(n6894) );
  NAND2_X1 U6751 ( .A1(n6920), .A2(n5464), .ZN(n5213) );
  NAND2_X1 U6752 ( .A1(n5210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5211) );
  XNOR2_X1 U6753 ( .A(n5211), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7054) );
  AOI22_X1 U6754 ( .A1(n5326), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5325), .B2(
        n7054), .ZN(n5212) );
  NAND2_X1 U6755 ( .A1(n5086), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5223) );
  INV_X1 U6756 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5214) );
  OR2_X1 U6757 ( .A1(n5215), .A2(n5214), .ZN(n5222) );
  INV_X1 U6758 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5216) );
  OAI21_X1 U6759 ( .B1(n5218), .B2(n5217), .A(n5216), .ZN(n5219) );
  NAND2_X1 U6760 ( .A1(n5219), .A2(n5236), .ZN(n6901) );
  OR2_X1 U6761 ( .A1(n5419), .A2(n6901), .ZN(n5221) );
  INV_X1 U6762 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6902) );
  OR2_X1 U6763 ( .A1(n8240), .A2(n6902), .ZN(n5220) );
  INV_X1 U6764 ( .A(n7656), .ZN(n8631) );
  NAND2_X1 U6765 ( .A1(n7007), .A2(n8631), .ZN(n5261) );
  AND2_X1 U6766 ( .A1(n6894), .A2(n5261), .ZN(n6989) );
  XNOR2_X1 U6767 ( .A(n5245), .B(n5244), .ZN(n7023) );
  NAND2_X1 U6768 ( .A1(n7023), .A2(n5464), .ZN(n5235) );
  AND3_X1 U6769 ( .A1(n5226), .A2(n5225), .A3(n5224), .ZN(n5227) );
  AND2_X1 U6770 ( .A1(n5228), .A2(n5227), .ZN(n5231) );
  NOR2_X1 U6771 ( .A1(n5231), .A2(n4889), .ZN(n5229) );
  MUX2_X1 U6772 ( .A(n4889), .B(n5229), .S(P2_IR_REG_12__SCAN_IN), .Z(n5233)
         );
  NAND2_X1 U6773 ( .A1(n5231), .A2(n5230), .ZN(n5250) );
  INV_X1 U6774 ( .A(n5250), .ZN(n5232) );
  AOI22_X1 U6775 ( .A1(n5326), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5325), .B2(
        n7222), .ZN(n5234) );
  NAND2_X1 U6776 ( .A1(n8237), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5241) );
  INV_X1 U6777 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7050) );
  OR2_X1 U6778 ( .A1(n5117), .A2(n7050), .ZN(n5240) );
  INV_X1 U6779 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U6780 ( .A1(n5236), .A2(n7058), .ZN(n5237) );
  NAND2_X1 U6781 ( .A1(n5255), .A2(n5237), .ZN(n7000) );
  OR2_X1 U6782 ( .A1(n5419), .A2(n7000), .ZN(n5239) );
  INV_X1 U6783 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7055) );
  OR2_X1 U6784 ( .A1(n5309), .A2(n7055), .ZN(n5238) );
  OR2_X1 U6785 ( .A1(n7128), .A2(n7108), .ZN(n8359) );
  INV_X1 U6786 ( .A(n8266), .ZN(n5242) );
  AND2_X1 U6787 ( .A1(n6989), .A2(n5242), .ZN(n5243) );
  NAND2_X1 U6788 ( .A1(n6893), .A2(n5243), .ZN(n7110) );
  NAND2_X1 U6789 ( .A1(n5268), .A2(n5246), .ZN(n5249) );
  AND2_X1 U6790 ( .A1(n5247), .A2(n5265), .ZN(n5248) );
  NAND2_X1 U6791 ( .A1(n7138), .A2(n5464), .ZN(n5253) );
  NAND2_X1 U6792 ( .A1(n5250), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5251) );
  XNOR2_X1 U6793 ( .A(n5251), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7409) );
  AOI22_X1 U6794 ( .A1(n5326), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5325), .B2(
        n7409), .ZN(n5252) );
  NAND2_X1 U6795 ( .A1(n8237), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5260) );
  INV_X1 U6796 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5254) );
  OR2_X1 U6797 ( .A1(n5309), .A2(n5254), .ZN(n5259) );
  NAND2_X1 U6798 ( .A1(n5255), .A2(n7227), .ZN(n5256) );
  NAND2_X1 U6799 ( .A1(n5279), .A2(n5256), .ZN(n7119) );
  OR2_X1 U6800 ( .A1(n5419), .A2(n7119), .ZN(n5258) );
  INV_X1 U6801 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7120) );
  OR2_X1 U6802 ( .A1(n5117), .A2(n7120), .ZN(n5257) );
  OR2_X1 U6803 ( .A1(n8952), .A2(n7211), .ZN(n8368) );
  NAND2_X1 U6804 ( .A1(n8952), .A2(n7211), .ZN(n7169) );
  OR2_X1 U6805 ( .A1(n7007), .A2(n7656), .ZN(n8338) );
  INV_X1 U6806 ( .A(n7108), .ZN(n8630) );
  OR2_X1 U6807 ( .A1(n7128), .A2(n8630), .ZN(n5262) );
  AND2_X1 U6808 ( .A1(n8374), .A2(n7109), .ZN(n5263) );
  NAND2_X1 U6809 ( .A1(n7110), .A2(n5263), .ZN(n7111) );
  INV_X1 U6810 ( .A(n7211), .ZN(n8629) );
  NAND2_X1 U6811 ( .A1(n8952), .A2(n8629), .ZN(n5264) );
  NAND2_X1 U6812 ( .A1(n7111), .A2(n5264), .ZN(n7167) );
  INV_X1 U6813 ( .A(n5265), .ZN(n5266) );
  XNOR2_X1 U6814 ( .A(n5270), .B(n5269), .ZN(n7233) );
  NAND2_X1 U6815 ( .A1(n7233), .A2(n5464), .ZN(n5277) );
  AND2_X1 U6816 ( .A1(n5271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6817 ( .A1(n5272), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5275) );
  INV_X1 U6818 ( .A(n5272), .ZN(n5274) );
  NAND2_X1 U6819 ( .A1(n5274), .A2(n5273), .ZN(n5287) );
  AOI22_X1 U6820 ( .A1(n5326), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5325), .B2(
        n7407), .ZN(n5276) );
  NAND2_X1 U6821 ( .A1(n8237), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5284) );
  INV_X1 U6822 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8645) );
  OR2_X1 U6823 ( .A1(n5309), .A2(n8645), .ZN(n5283) );
  NAND2_X1 U6824 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  NAND2_X1 U6825 ( .A1(n5293), .A2(n5280), .ZN(n7210) );
  OR2_X1 U6826 ( .A1(n5419), .A2(n7210), .ZN(n5282) );
  INV_X1 U6827 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8643) );
  OR2_X1 U6828 ( .A1(n8240), .A2(n8643), .ZN(n5281) );
  NAND2_X1 U6829 ( .A1(n7214), .A2(n7261), .ZN(n8377) );
  NAND2_X1 U6830 ( .A1(n8378), .A2(n8377), .ZN(n8372) );
  INV_X1 U6831 ( .A(n7261), .ZN(n8628) );
  OAI22_X1 U6832 ( .A1(n7167), .A2(n8268), .B1(n7214), .B2(n8628), .ZN(n7264)
         );
  XNOR2_X1 U6833 ( .A(n5286), .B(n5285), .ZN(n7338) );
  NAND2_X1 U6834 ( .A1(n7338), .A2(n5464), .ZN(n5290) );
  NAND2_X1 U6835 ( .A1(n5287), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5288) );
  XNOR2_X1 U6836 ( .A(n5288), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8667) );
  AOI22_X1 U6837 ( .A1(n5326), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5325), .B2(
        n8667), .ZN(n5289) );
  NAND2_X1 U6838 ( .A1(n8237), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5299) );
  INV_X1 U6839 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5291) );
  OR2_X1 U6840 ( .A1(n5309), .A2(n5291), .ZN(n5298) );
  INV_X1 U6841 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6842 ( .A1(n5293), .A2(n5292), .ZN(n5294) );
  NAND2_X1 U6843 ( .A1(n5310), .A2(n5294), .ZN(n7693) );
  OR2_X1 U6844 ( .A1(n5419), .A2(n7693), .ZN(n5297) );
  INV_X1 U6845 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5295) );
  OR2_X1 U6846 ( .A1(n5117), .A2(n5295), .ZN(n5296) );
  XNOR2_X1 U6847 ( .A(n8947), .B(n8382), .ZN(n8376) );
  NAND2_X1 U6848 ( .A1(n7264), .A2(n8376), .ZN(n7263) );
  INV_X1 U6849 ( .A(n8382), .ZN(n8627) );
  OR2_X1 U6850 ( .A1(n8947), .A2(n8627), .ZN(n5300) );
  XNOR2_X1 U6851 ( .A(n5302), .B(n5301), .ZN(n7455) );
  NAND2_X1 U6852 ( .A1(n7455), .A2(n5464), .ZN(n5308) );
  MUX2_X1 U6853 ( .A(n4889), .B(n4370), .S(P2_IR_REG_16__SCAN_IN), .Z(n5303)
         );
  INV_X1 U6854 ( .A(n5303), .ZN(n5306) );
  INV_X1 U6855 ( .A(n5304), .ZN(n5305) );
  AND2_X1 U6856 ( .A1(n5306), .A2(n5305), .ZN(n8681) );
  AOI22_X1 U6857 ( .A1(n5326), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5325), .B2(
        n8681), .ZN(n5307) );
  NAND2_X1 U6858 ( .A1(n8237), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5316) );
  INV_X1 U6859 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8658) );
  OR2_X1 U6860 ( .A1(n5309), .A2(n8658), .ZN(n5315) );
  INV_X1 U6861 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U6862 ( .A1(n5310), .A2(n8661), .ZN(n5311) );
  NAND2_X1 U6863 ( .A1(n5312), .A2(n5311), .ZN(n7443) );
  OR2_X1 U6864 ( .A1(n5419), .A2(n7443), .ZN(n5314) );
  INV_X1 U6865 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7330) );
  OR2_X1 U6866 ( .A1(n8240), .A2(n7330), .ZN(n5313) );
  OR2_X1 U6867 ( .A1(n8941), .A2(n7509), .ZN(n8388) );
  NAND2_X1 U6868 ( .A1(n8941), .A2(n7509), .ZN(n8387) );
  INV_X1 U6869 ( .A(n8941), .ZN(n7329) );
  NAND2_X1 U6870 ( .A1(n5318), .A2(n7565), .ZN(n8290) );
  NAND2_X1 U6871 ( .A1(n8289), .A2(n8290), .ZN(n8270) );
  AND2_X1 U6872 ( .A1(n7563), .A2(n8624), .ZN(n5503) );
  INV_X1 U6873 ( .A(n5503), .ZN(n8394) );
  NAND2_X1 U6874 ( .A1(n8932), .A2(n7394), .ZN(n8402) );
  XNOR2_X1 U6875 ( .A(n5320), .B(n5319), .ZN(n7803) );
  NAND2_X1 U6876 ( .A1(n7803), .A2(n5464), .ZN(n5328) );
  NAND2_X1 U6877 ( .A1(n5321), .A2(n5477), .ZN(n5322) );
  NAND2_X1 U6878 ( .A1(n5322), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6879 ( .A1(n5323), .A2(n5476), .ZN(n5472) );
  OR2_X1 U6880 ( .A1(n5323), .A2(n5476), .ZN(n5324) );
  AOI22_X1 U6881 ( .A1(n5326), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7547), .B2(
        n5325), .ZN(n5327) );
  INV_X1 U6882 ( .A(n8927), .ZN(n7550) );
  INV_X1 U6883 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6884 ( .A1(n5330), .A2(n5329), .ZN(n5331) );
  NAND2_X1 U6885 ( .A1(n5349), .A2(n5331), .ZN(n7589) );
  OR2_X1 U6886 ( .A1(n7589), .A2(n5419), .ZN(n5334) );
  AOI22_X1 U6887 ( .A1(n5086), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n8237), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6888 ( .A1(n5351), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6889 ( .A1(n7550), .A2(n7633), .ZN(n5335) );
  INV_X1 U6890 ( .A(n7633), .ZN(n8623) );
  XNOR2_X1 U6891 ( .A(n5337), .B(n5336), .ZN(n6836) );
  NAND2_X1 U6892 ( .A1(n6836), .A2(n5464), .ZN(n5339) );
  OR2_X1 U6893 ( .A1(n5097), .A2(n8207), .ZN(n5338) );
  XNOR2_X1 U6894 ( .A(n5349), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n7630) );
  INV_X1 U6895 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6896 ( .A1(n5086), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6897 ( .A1(n8237), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5340) );
  OAI211_X1 U6898 ( .C1(n5342), .C2(n8240), .A(n5341), .B(n5340), .ZN(n5343)
         );
  AOI21_X1 U6899 ( .B1(n7630), .B2(n4469), .A(n5343), .ZN(n8858) );
  OR2_X1 U6900 ( .A1(n5344), .A2(n8858), .ZN(n8407) );
  NAND2_X1 U6901 ( .A1(n5344), .A2(n8858), .ZN(n8405) );
  INV_X1 U6902 ( .A(n5344), .ZN(n7618) );
  XNOR2_X1 U6903 ( .A(n5346), .B(n5345), .ZN(n7780) );
  NAND2_X1 U6904 ( .A1(n7780), .A2(n5464), .ZN(n5348) );
  INV_X1 U6905 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6877) );
  OR2_X1 U6906 ( .A1(n5097), .A2(n6877), .ZN(n5347) );
  INV_X1 U6907 ( .A(n8916), .ZN(n8870) );
  INV_X1 U6908 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7631) );
  INV_X1 U6909 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8569) );
  OAI21_X1 U6910 ( .B1(n5349), .B2(n7631), .A(n8569), .ZN(n5350) );
  AND2_X1 U6911 ( .A1(n5350), .A2(n5358), .ZN(n8866) );
  NAND2_X1 U6912 ( .A1(n8866), .A2(n4469), .ZN(n5354) );
  AOI22_X1 U6913 ( .A1(n5086), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n8237), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6914 ( .A1(n5351), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5352) );
  NOR2_X1 U6915 ( .A1(n8870), .A2(n8844), .ZN(n5355) );
  INV_X1 U6916 ( .A(n8844), .ZN(n8622) );
  OAI22_X1 U6917 ( .A1(n8852), .A2(n5355), .B1(n8622), .B2(n8916), .ZN(n8835)
         );
  XNOR2_X1 U6918 ( .A(n5367), .B(n5366), .ZN(n7768) );
  NAND2_X1 U6919 ( .A1(n7768), .A2(n5464), .ZN(n5357) );
  OR2_X1 U6920 ( .A1(n5097), .A2(n7006), .ZN(n5356) );
  INV_X1 U6921 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U6922 ( .A1(n5358), .A2(n10029), .ZN(n5359) );
  NAND2_X1 U6923 ( .A1(n5375), .A2(n5359), .ZN(n8839) );
  OR2_X1 U6924 ( .A1(n8839), .A2(n5419), .ZN(n5365) );
  INV_X1 U6925 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6926 ( .A1(n8237), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6927 ( .A1(n5086), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5360) );
  OAI211_X1 U6928 ( .C1(n8240), .C2(n5362), .A(n5361), .B(n5360), .ZN(n5363)
         );
  INV_X1 U6929 ( .A(n5363), .ZN(n5364) );
  NAND2_X1 U6930 ( .A1(n5365), .A2(n5364), .ZN(n8621) );
  INV_X1 U6931 ( .A(n8834), .ZN(n8843) );
  NAND2_X1 U6932 ( .A1(n5385), .A2(n5368), .ZN(n5371) );
  AND2_X1 U6933 ( .A1(n5369), .A2(n5387), .ZN(n5370) );
  NAND2_X1 U6934 ( .A1(n7816), .A2(n5464), .ZN(n5373) );
  OR2_X1 U6935 ( .A1(n5097), .A2(n9886), .ZN(n5372) );
  NAND2_X1 U6936 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  NAND2_X1 U6937 ( .A1(n5377), .A2(n5376), .ZN(n8824) );
  OR2_X1 U6938 ( .A1(n8824), .A2(n5419), .ZN(n5382) );
  INV_X1 U6939 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U6940 ( .A1(n5086), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6941 ( .A1(n8237), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5378) );
  OAI211_X1 U6942 ( .C1(n8825), .C2(n5117), .A(n5379), .B(n5378), .ZN(n5380)
         );
  INV_X1 U6943 ( .A(n5380), .ZN(n5381) );
  XNOR2_X1 U6944 ( .A(n8905), .B(n8845), .ZN(n8821) );
  NAND2_X1 U6945 ( .A1(n8822), .A2(n8821), .ZN(n8903) );
  NAND2_X1 U6946 ( .A1(n8898), .A2(n8586), .ZN(n8418) );
  NAND2_X1 U6947 ( .A1(n8419), .A2(n8418), .ZN(n8808) );
  INV_X1 U6948 ( .A(n5386), .ZN(n5388) );
  INV_X1 U6949 ( .A(n5391), .ZN(n5392) );
  NAND2_X1 U6950 ( .A1(n5392), .A2(SI_24_), .ZN(n5393) );
  MUX2_X1 U6951 ( .A(n7275), .B(n7757), .S(n5942), .Z(n5396) );
  INV_X1 U6952 ( .A(SI_25_), .ZN(n5395) );
  NAND2_X1 U6953 ( .A1(n5396), .A2(n5395), .ZN(n5409) );
  INV_X1 U6954 ( .A(n5396), .ZN(n5397) );
  NAND2_X1 U6955 ( .A1(n5397), .A2(SI_25_), .ZN(n5398) );
  NAND2_X1 U6956 ( .A1(n5409), .A2(n5398), .ZN(n5408) );
  XNOR2_X1 U6957 ( .A(n5407), .B(n5408), .ZN(n7756) );
  NAND2_X1 U6958 ( .A1(n7756), .A2(n5464), .ZN(n5400) );
  OR2_X1 U6959 ( .A1(n5097), .A2(n7275), .ZN(n5399) );
  INV_X1 U6960 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6961 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  AND2_X1 U6962 ( .A1(n5417), .A2(n5403), .ZN(n8579) );
  INV_X1 U6963 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U6964 ( .A1(n5086), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6965 ( .A1(n8237), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5404) );
  OAI211_X1 U6966 ( .C1(n8786), .C2(n5117), .A(n5405), .B(n5404), .ZN(n5406)
         );
  AOI21_X1 U6967 ( .B1(n8579), .B2(n4469), .A(n5406), .ZN(n8809) );
  OR2_X1 U6968 ( .A1(n8894), .A2(n8809), .ZN(n5506) );
  NAND2_X1 U6969 ( .A1(n8894), .A2(n8809), .ZN(n8423) );
  NAND2_X1 U6970 ( .A1(n5506), .A2(n8423), .ZN(n8789) );
  INV_X1 U6971 ( .A(n8809), .ZN(n8618) );
  INV_X1 U6972 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7364) );
  INV_X1 U6973 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7744) );
  MUX2_X1 U6974 ( .A(n7364), .B(n7744), .S(n5942), .Z(n5411) );
  INV_X1 U6975 ( .A(SI_26_), .ZN(n5410) );
  NAND2_X1 U6976 ( .A1(n5411), .A2(n5410), .ZN(n5427) );
  INV_X1 U6977 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U6978 ( .A1(n5412), .A2(SI_26_), .ZN(n5413) );
  XNOR2_X1 U6979 ( .A(n5426), .B(n5425), .ZN(n7743) );
  NAND2_X1 U6980 ( .A1(n7743), .A2(n5464), .ZN(n5415) );
  OR2_X1 U6981 ( .A1(n5097), .A2(n7364), .ZN(n5414) );
  INV_X1 U6982 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U6983 ( .A1(n5417), .A2(n8212), .ZN(n5418) );
  NAND2_X1 U6984 ( .A1(n5446), .A2(n5418), .ZN(n8779) );
  OR2_X1 U6985 ( .A1(n8779), .A2(n5419), .ZN(n5424) );
  INV_X1 U6986 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U6987 ( .A1(n5086), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6988 ( .A1(n8237), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5420) );
  OAI211_X1 U6989 ( .C1(n8780), .C2(n8240), .A(n5421), .B(n5420), .ZN(n5422)
         );
  INV_X1 U6990 ( .A(n5422), .ZN(n5423) );
  OR2_X1 U6991 ( .A1(n8889), .A2(n8761), .ZN(n8427) );
  NAND2_X1 U6992 ( .A1(n8889), .A2(n8761), .ZN(n8425) );
  NAND2_X1 U6993 ( .A1(n8427), .A2(n8425), .ZN(n8771) );
  INV_X1 U6994 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7452) );
  MUX2_X1 U6995 ( .A(n7452), .B(n7734), .S(n5942), .Z(n5430) );
  INV_X1 U6996 ( .A(SI_27_), .ZN(n5429) );
  NAND2_X1 U6997 ( .A1(n5430), .A2(n5429), .ZN(n5442) );
  INV_X1 U6998 ( .A(n5430), .ZN(n5431) );
  NAND2_X1 U6999 ( .A1(n5431), .A2(SI_27_), .ZN(n5432) );
  NAND2_X1 U7000 ( .A1(n7733), .A2(n5464), .ZN(n5434) );
  OR2_X1 U7001 ( .A1(n5097), .A2(n7452), .ZN(n5433) );
  XNOR2_X1 U7002 ( .A(n5446), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8756) );
  INV_X1 U7003 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U7004 ( .A1(n5086), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U7005 ( .A1(n8237), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5435) );
  OAI211_X1 U7006 ( .C1(n5437), .C2(n5117), .A(n5436), .B(n5435), .ZN(n5438)
         );
  NAND2_X1 U7007 ( .A1(n8883), .A2(n8747), .ZN(n8429) );
  INV_X1 U7008 ( .A(n8759), .ZN(n5439) );
  INV_X1 U7009 ( .A(n8747), .ZN(n8616) );
  INV_X1 U7010 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7882) );
  INV_X1 U7011 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8234) );
  MUX2_X1 U7012 ( .A(n7882), .B(n8234), .S(n7725), .Z(n5459) );
  XNOR2_X1 U7013 ( .A(n5459), .B(SI_28_), .ZN(n5456) );
  XNOR2_X1 U7014 ( .A(n5457), .B(n5456), .ZN(n7881) );
  NAND2_X1 U7015 ( .A1(n7881), .A2(n5464), .ZN(n5445) );
  OR2_X1 U7016 ( .A1(n5097), .A2(n8234), .ZN(n5444) );
  INV_X1 U7017 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8551) );
  INV_X1 U7018 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8200) );
  OAI21_X1 U7019 ( .B1(n5446), .B2(n8551), .A(n8200), .ZN(n5447) );
  NAND2_X1 U7020 ( .A1(n8741), .A2(n4469), .ZN(n5453) );
  INV_X1 U7021 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U7022 ( .A1(n5086), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U7023 ( .A1(n8237), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5448) );
  OAI211_X1 U7024 ( .C1(n5450), .C2(n5117), .A(n5449), .B(n5448), .ZN(n5451)
         );
  INV_X1 U7025 ( .A(n5451), .ZN(n5452) );
  XNOR2_X1 U7026 ( .A(n8878), .B(n8762), .ZN(n8744) );
  NAND2_X1 U7027 ( .A1(n8743), .A2(n8762), .ZN(n5454) );
  NAND2_X1 U7028 ( .A1(n5455), .A2(n5454), .ZN(n5471) );
  INV_X1 U7029 ( .A(SI_28_), .ZN(n5458) );
  NAND2_X1 U7030 ( .A1(n5459), .A2(n5458), .ZN(n5460) );
  MUX2_X1 U7031 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n7725), .Z(n7712) );
  INV_X1 U7032 ( .A(SI_29_), .ZN(n5462) );
  XNOR2_X1 U7033 ( .A(n7712), .B(n5462), .ZN(n5463) );
  NAND2_X1 U7034 ( .A1(n7897), .A2(n5464), .ZN(n5466) );
  INV_X1 U7035 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7499) );
  OR2_X1 U7036 ( .A1(n5097), .A2(n7499), .ZN(n5465) );
  INV_X1 U7037 ( .A(n7703), .ZN(n5470) );
  INV_X1 U7038 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7702) );
  NAND2_X1 U7039 ( .A1(n8237), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U7040 ( .A1(n5086), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5467) );
  OAI211_X1 U7041 ( .C1(n7702), .C2(n8240), .A(n5468), .B(n5467), .ZN(n5469)
         );
  AOI21_X1 U7042 ( .B1(n5470), .B2(n4469), .A(n5469), .ZN(n8746) );
  OR2_X1 U7043 ( .A1(n7700), .A2(n8746), .ZN(n8436) );
  NAND2_X1 U7044 ( .A1(n8436), .A2(n4325), .ZN(n8279) );
  INV_X1 U7045 ( .A(n8279), .ZN(n8434) );
  XNOR2_X1 U7046 ( .A(n5471), .B(n8279), .ZN(n7699) );
  NAND2_X1 U7047 ( .A1(n5472), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U7048 ( .A1(n5480), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U7049 ( .A1(n6216), .A2(n5517), .ZN(n5483) );
  NAND2_X1 U7050 ( .A1(n8454), .A2(n8303), .ZN(n5721) );
  AND2_X1 U7051 ( .A1(n5721), .A2(n9744), .ZN(n5482) );
  NAND2_X1 U7052 ( .A1(n7699), .A2(n9800), .ZN(n5519) );
  NAND2_X1 U7053 ( .A1(n6771), .A2(n9762), .ZN(n6389) );
  NAND2_X1 U7054 ( .A1(n8305), .A2(n8313), .ZN(n6444) );
  INV_X1 U7055 ( .A(n6444), .ZN(n5484) );
  NAND2_X1 U7056 ( .A1(n5484), .A2(n8253), .ZN(n6442) );
  NAND2_X1 U7057 ( .A1(n6442), .A2(n8316), .ZN(n5485) );
  INV_X1 U7058 ( .A(n8254), .ZN(n8307) );
  NAND2_X1 U7059 ( .A1(n6470), .A2(n6395), .ZN(n8258) );
  NAND2_X1 U7060 ( .A1(n8218), .A2(n6630), .ZN(n8327) );
  NAND2_X1 U7061 ( .A1(n8353), .A2(n8294), .ZN(n8333) );
  NOR2_X1 U7062 ( .A1(n8333), .A2(n7651), .ZN(n5492) );
  INV_X1 U7063 ( .A(n5492), .ZN(n5488) );
  NAND2_X1 U7064 ( .A1(n8332), .A2(n5488), .ZN(n5489) );
  OR2_X1 U7065 ( .A1(n5489), .A2(n8335), .ZN(n5494) );
  AND2_X1 U7066 ( .A1(n8353), .A2(n8294), .ZN(n5490) );
  AND2_X1 U7067 ( .A1(n8347), .A2(n5490), .ZN(n5491) );
  NAND2_X1 U7068 ( .A1(n8337), .A2(n4848), .ZN(n5493) );
  AND2_X1 U7069 ( .A1(n8359), .A2(n8338), .ZN(n8364) );
  NAND2_X1 U7070 ( .A1(n5495), .A2(n8362), .ZN(n7107) );
  INV_X1 U7071 ( .A(n7169), .ZN(n8370) );
  NOR2_X1 U7072 ( .A1(n8372), .A2(n8370), .ZN(n5496) );
  NAND2_X1 U7073 ( .A1(n8947), .A2(n8382), .ZN(n7320) );
  INV_X1 U7074 ( .A(n8387), .ZN(n5498) );
  AND2_X1 U7075 ( .A1(n7320), .A2(n5500), .ZN(n5499) );
  INV_X1 U7076 ( .A(n5500), .ZN(n5501) );
  AND2_X1 U7077 ( .A1(n7505), .A2(n8289), .ZN(n5502) );
  NAND2_X1 U7078 ( .A1(n7506), .A2(n5502), .ZN(n7564) );
  AOI21_X1 U7079 ( .B1(n7564), .B2(n8402), .A(n5503), .ZN(n7542) );
  OR2_X1 U7080 ( .A1(n8927), .A2(n7633), .ZN(n8400) );
  NAND2_X1 U7081 ( .A1(n8927), .A2(n7633), .ZN(n8404) );
  INV_X1 U7082 ( .A(n8404), .ZN(n5504) );
  XNOR2_X1 U7083 ( .A(n8916), .B(n8844), .ZN(n8855) );
  INV_X1 U7084 ( .A(n8396), .ZN(n8413) );
  NAND2_X1 U7085 ( .A1(n8847), .A2(n8413), .ZN(n8815) );
  NAND2_X1 U7086 ( .A1(n8905), .A2(n8845), .ZN(n8416) );
  OAI21_X1 U7087 ( .B1(n8815), .B2(n8821), .A(n8416), .ZN(n8807) );
  INV_X1 U7088 ( .A(n8419), .ZN(n5505) );
  INV_X1 U7089 ( .A(n5506), .ZN(n8772) );
  INV_X1 U7090 ( .A(n8425), .ZN(n8760) );
  INV_X1 U7091 ( .A(n8428), .ZN(n5507) );
  NAND2_X1 U7092 ( .A1(n8448), .A2(n8303), .ZN(n8249) );
  INV_X1 U7093 ( .A(n5509), .ZN(n5511) );
  INV_X1 U7094 ( .A(n5508), .ZN(n5510) );
  AOI21_X1 U7095 ( .B1(n5511), .B2(P2_B_REG_SCAN_IN), .A(n8861), .ZN(n8726) );
  INV_X1 U7096 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U7097 ( .A1(n5086), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7098 ( .A1(n8237), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5512) );
  OAI211_X1 U7099 ( .C1(n8240), .C2(n8732), .A(n5513), .B(n5512), .ZN(n8614)
         );
  NAND2_X1 U7100 ( .A1(n6539), .A2(n9780), .ZN(n6554) );
  INV_X1 U7101 ( .A(n6555), .ZN(n9785) );
  NOR2_X2 U7102 ( .A1(n6359), .A2(n8219), .ZN(n6403) );
  INV_X1 U7103 ( .A(n6479), .ZN(n6509) );
  INV_X1 U7104 ( .A(n7007), .ZN(n6900) );
  NAND2_X1 U7105 ( .A1(n6898), .A2(n6900), .ZN(n6997) );
  INV_X1 U7106 ( .A(n7214), .ZN(n9527) );
  INV_X1 U7107 ( .A(n8947), .ZN(n8383) );
  NAND2_X1 U7108 ( .A1(n8805), .A2(n8819), .ZN(n8799) );
  NOR2_X2 U7109 ( .A1(n8799), .A2(n8894), .ZN(n8792) );
  NAND2_X1 U7110 ( .A1(n8781), .A2(n8792), .ZN(n8754) );
  AOI21_X1 U7111 ( .B1(n7700), .B2(n8738), .A(n8730), .ZN(n7706) );
  AOI22_X1 U7112 ( .A1(n7706), .A2(n9786), .B1(n9772), .B2(n7700), .ZN(n5518)
         );
  NAND2_X1 U7113 ( .A1(n5520), .A2(n5481), .ZN(n5521) );
  NAND2_X1 U7114 ( .A1(n5548), .A2(n5522), .ZN(n5523) );
  XNOR2_X1 U7115 ( .A(n7077), .B(P2_B_REG_SCAN_IN), .ZN(n5531) );
  INV_X1 U7116 ( .A(n5526), .ZN(n5527) );
  NAND2_X1 U7117 ( .A1(n5527), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5528) );
  MUX2_X1 U7118 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5528), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5530) );
  NAND2_X1 U7119 ( .A1(n5530), .A2(n5529), .ZN(n7273) );
  NAND2_X1 U7120 ( .A1(n5531), .A2(n7273), .ZN(n5536) );
  NAND2_X1 U7121 ( .A1(n5529), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5532) );
  MUX2_X1 U7122 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5532), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5533) );
  INV_X1 U7123 ( .A(n7365), .ZN(n5535) );
  INV_X1 U7124 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9759) );
  AND2_X1 U7125 ( .A1(n7365), .A2(n7273), .ZN(n9761) );
  NOR2_X1 U7126 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .ZN(
        n5540) );
  NOR4_X1 U7127 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5539) );
  NOR4_X1 U7128 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5538) );
  NOR4_X1 U7129 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5537) );
  AND4_X1 U7130 ( .A1(n5540), .A2(n5539), .A3(n5538), .A4(n5537), .ZN(n5546)
         );
  NOR4_X1 U7131 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5544) );
  NOR4_X1 U7132 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5543) );
  NOR4_X1 U7133 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5542) );
  NOR4_X1 U7134 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5541) );
  AND4_X1 U7135 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .ZN(n5545)
         );
  NAND2_X1 U7136 ( .A1(n5546), .A2(n5545), .ZN(n5547) );
  NAND2_X1 U7137 ( .A1(n9753), .A2(n5547), .ZN(n5626) );
  INV_X1 U7138 ( .A(n5721), .ZN(n5748) );
  AND2_X1 U7139 ( .A1(n5748), .A2(n8453), .ZN(n5635) );
  NOR2_X1 U7140 ( .A1(n9754), .A2(n5635), .ZN(n5549) );
  NAND2_X1 U7141 ( .A1(n5626), .A2(n5549), .ZN(n6207) );
  INV_X1 U7142 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9756) );
  NAND2_X1 U7143 ( .A1(n9753), .A2(n9756), .ZN(n5551) );
  INV_X1 U7144 ( .A(n6369), .ZN(n5627) );
  NAND2_X1 U7145 ( .A1(n8877), .A2(n9817), .ZN(n5554) );
  INV_X1 U7146 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5552) );
  OR2_X1 U7147 ( .A1(n9817), .A2(n5552), .ZN(n5553) );
  NAND2_X1 U7148 ( .A1(n5554), .A2(n5553), .ZN(P2_U3517) );
  AND2_X2 U7149 ( .A1(n5558), .A2(n5557), .ZN(n5672) );
  NAND3_X1 U7150 ( .A1(n5682), .A2(n5672), .A3(n5559), .ZN(n5726) );
  NOR2_X1 U7151 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5563) );
  NOR2_X1 U7152 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5562) );
  NAND2_X1 U7153 ( .A1(n5590), .A2(n5567), .ZN(n5569) );
  OR2_X1 U7154 ( .A1(n5590), .A2(n5567), .ZN(n5568) );
  NAND2_X1 U7155 ( .A1(n5569), .A2(n5568), .ZN(n7272) );
  NAND2_X1 U7156 ( .A1(n4350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5571) );
  INV_X1 U7157 ( .A(n5572), .ZN(n5573) );
  NAND2_X1 U7158 ( .A1(n5573), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7159 ( .A1(n5932), .A2(n6130), .ZN(n5732) );
  OR2_X2 U7160 ( .A1(n5732), .A2(P1_U3084), .ZN(n9119) );
  INV_X1 U7161 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6227) );
  INV_X1 U7162 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6177) );
  NAND4_X1 U7163 ( .A1(n6227), .A2(n5578), .A3(n6177), .A4(n6153), .ZN(n5580)
         );
  NAND2_X1 U7164 ( .A1(n10016), .A2(n6245), .ZN(n5579) );
  NAND2_X1 U7165 ( .A1(n5885), .A2(n5886), .ZN(n5581) );
  NAND2_X1 U7166 ( .A1(n5585), .A2(n5584), .ZN(n5586) );
  INV_X1 U7167 ( .A(n6130), .ZN(n7046) );
  OR2_X1 U7168 ( .A1(n8061), .A2(n7046), .ZN(n5587) );
  NAND2_X1 U7169 ( .A1(n5587), .A2(n5732), .ZN(n5734) );
  INV_X1 U7170 ( .A(n5692), .ZN(n5588) );
  NAND2_X1 U7171 ( .A1(n5588), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5589) );
  INV_X1 U7172 ( .A(n5593), .ZN(n5591) );
  NAND2_X1 U7173 ( .A1(n5591), .A2(n4849), .ZN(n5592) );
  XNOR2_X1 U7174 ( .A(n5593), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5594) );
  NAND2_X2 U7175 ( .A1(n5735), .A2(n5594), .ZN(n5944) );
  OAI21_X1 U7176 ( .B1(n5734), .B2(n5941), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  INV_X1 U7177 ( .A(n9763), .ZN(n5595) );
  NAND2_X1 U7178 ( .A1(n6217), .A2(n8250), .ZN(n6772) );
  OR2_X1 U7179 ( .A1(n5614), .A2(n9762), .ZN(n5596) );
  AND2_X1 U7180 ( .A1(n6772), .A2(n5596), .ZN(n6251) );
  NAND2_X1 U7181 ( .A1(n6250), .A2(n6251), .ZN(n7672) );
  INV_X1 U7182 ( .A(n5597), .ZN(n7671) );
  NAND2_X1 U7183 ( .A1(n5598), .A2(n7671), .ZN(n5599) );
  NAND2_X1 U7184 ( .A1(n7672), .A2(n5599), .ZN(n5600) );
  OR2_X1 U7185 ( .A1(n5082), .A2(n8187), .ZN(n5603) );
  XNOR2_X1 U7186 ( .A(n9771), .B(n5614), .ZN(n5601) );
  XNOR2_X1 U7187 ( .A(n5603), .B(n5601), .ZN(n7673) );
  NAND2_X1 U7188 ( .A1(n5600), .A2(n7673), .ZN(n5647) );
  INV_X1 U7189 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U7190 ( .A1(n5603), .A2(n5602), .ZN(n5648) );
  NOR2_X1 U7191 ( .A1(n5100), .A2(n8187), .ZN(n5604) );
  XNOR2_X1 U7192 ( .A(n6542), .B(n5614), .ZN(n6807) );
  NAND2_X1 U7193 ( .A1(n5604), .A2(n6807), .ZN(n5610) );
  INV_X1 U7194 ( .A(n5604), .ZN(n5606) );
  INV_X1 U7195 ( .A(n6807), .ZN(n5605) );
  NAND2_X1 U7196 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  NAND2_X1 U7197 ( .A1(n5610), .A2(n5607), .ZN(n5651) );
  INV_X1 U7198 ( .A(n5651), .ZN(n5608) );
  AND2_X1 U7199 ( .A1(n5648), .A2(n5608), .ZN(n5609) );
  XNOR2_X1 U7200 ( .A(n6555), .B(n8173), .ZN(n5611) );
  NAND2_X1 U7201 ( .A1(n8638), .A2(n8250), .ZN(n5612) );
  XNOR2_X1 U7202 ( .A(n5611), .B(n5612), .ZN(n6806) );
  INV_X1 U7203 ( .A(n5611), .ZN(n8226) );
  NAND2_X1 U7204 ( .A1(n8226), .A2(n5612), .ZN(n5613) );
  OR2_X1 U7205 ( .A1(n6632), .A2(n8187), .ZN(n5616) );
  XNOR2_X1 U7206 ( .A(n8219), .B(n8195), .ZN(n5615) );
  XNOR2_X1 U7207 ( .A(n5616), .B(n5615), .ZN(n8224) );
  INV_X1 U7208 ( .A(n5615), .ZN(n6638) );
  NAND2_X1 U7209 ( .A1(n5616), .A2(n6638), .ZN(n5617) );
  XNOR2_X1 U7210 ( .A(n9794), .B(n8173), .ZN(n5618) );
  OR2_X1 U7211 ( .A1(n8218), .A2(n8187), .ZN(n5619) );
  XNOR2_X1 U7212 ( .A(n5618), .B(n5619), .ZN(n6636) );
  INV_X1 U7213 ( .A(n5618), .ZN(n5620) );
  NAND2_X1 U7214 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  XNOR2_X1 U7215 ( .A(n6479), .B(n8195), .ZN(n5622) );
  NOR2_X1 U7216 ( .A1(n6741), .A2(n8187), .ZN(n5623) );
  NAND2_X1 U7217 ( .A1(n5622), .A2(n5623), .ZN(n6733) );
  INV_X1 U7218 ( .A(n5622), .ZN(n6732) );
  INV_X1 U7219 ( .A(n5623), .ZN(n5624) );
  NAND2_X1 U7220 ( .A1(n6732), .A2(n5624), .ZN(n5625) );
  NAND2_X1 U7221 ( .A1(n6733), .A2(n5625), .ZN(n5630) );
  NAND3_X1 U7222 ( .A1(n5627), .A2(n6206), .A3(n5626), .ZN(n5641) );
  OR3_X2 U7223 ( .A1(n5632), .A2(n5748), .A3(n9772), .ZN(n8587) );
  INV_X1 U7224 ( .A(n6734), .ZN(n5629) );
  AOI211_X1 U7225 ( .C1(n5631), .C2(n5630), .A(n8587), .B(n5629), .ZN(n5646)
         );
  NOR2_X1 U7226 ( .A1(n8607), .A2(n8218), .ZN(n5645) );
  NAND2_X1 U7227 ( .A1(n9763), .A2(n8448), .ZN(n9739) );
  OR2_X1 U7228 ( .A1(n5632), .A2(n9739), .ZN(n5634) );
  INV_X1 U7229 ( .A(n5633), .ZN(n5640) );
  INV_X1 U7231 ( .A(n8583), .ZN(n8596) );
  OAI22_X1 U7232 ( .A1(n8596), .A2(n6509), .B1(n8608), .B2(n6820), .ZN(n5644)
         );
  INV_X1 U7233 ( .A(n5635), .ZN(n5638) );
  INV_X1 U7234 ( .A(n5722), .ZN(n5636) );
  NAND3_X1 U7235 ( .A1(n5638), .A2(n5637), .A3(n5636), .ZN(n5639) );
  AOI21_X1 U7236 ( .B1(n5641), .B2(n5640), .A(n5639), .ZN(n5642) );
  OR2_X2 U7237 ( .A1(n5642), .A2(P2_U3152), .ZN(n8606) );
  OAI22_X1 U7238 ( .A1(n8606), .A2(n6508), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5823), .ZN(n5643) );
  OR4_X1 U7239 ( .A1(n5646), .A2(n5645), .A3(n5644), .A4(n5643), .ZN(P2_U3215)
         );
  NAND2_X1 U7240 ( .A1(n5647), .A2(n5648), .ZN(n5650) );
  INV_X1 U7241 ( .A(n6805), .ZN(n5649) );
  AOI211_X1 U7242 ( .C1(n5651), .C2(n5650), .A(n8587), .B(n5649), .ZN(n5655)
         );
  NOR2_X1 U7243 ( .A1(n8607), .A2(n5082), .ZN(n5654) );
  OAI22_X1 U7244 ( .A1(n8596), .A2(n9780), .B1(n8608), .B2(n8221), .ZN(n5653)
         );
  OAI22_X1 U7245 ( .A1(n8606), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n4468), .ZN(n5652) );
  OR4_X1 U7246 ( .A1(n5655), .A2(n5654), .A3(n5653), .A4(n5652), .ZN(P2_U3220)
         );
  INV_X2 U7247 ( .A(n6150), .ZN(n8979) );
  NAND2_X1 U7248 ( .A1(n7725), .A2(P2_U3152), .ZN(n8233) );
  OAI222_X1 U7249 ( .A1(n8979), .A2(n5656), .B1(n8233), .B2(n5943), .C1(
        P2_U3152), .C2(n5764), .ZN(P2_U3357) );
  INV_X1 U7250 ( .A(n8233), .ZN(n7043) );
  OAI222_X1 U7251 ( .A1(n8979), .A2(n5657), .B1(n8980), .B2(n5988), .C1(
        P2_U3152), .C2(n5765), .ZN(P2_U3356) );
  OAI222_X1 U7252 ( .A1(n8979), .A2(n5658), .B1(n8980), .B2(n6087), .C1(
        P2_U3152), .C2(n5814), .ZN(P2_U3355) );
  OAI222_X1 U7253 ( .A1(n8979), .A2(n5659), .B1(n8980), .B2(n6052), .C1(
        P2_U3152), .C2(n5785), .ZN(P2_U3354) );
  NAND2_X2 U7254 ( .A1(n5942), .A2(P1_U3084), .ZN(n9493) );
  INV_X1 U7255 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7256 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5662), .ZN(n5660) );
  OAI222_X1 U7257 ( .A1(n9495), .A2(n5989), .B1(n9493), .B2(n5988), .C1(
        P1_U3084), .C2(n9591), .ZN(P1_U3351) );
  INV_X1 U7258 ( .A(n5861), .ZN(n6091) );
  OAI222_X1 U7259 ( .A1(n9495), .A2(n6088), .B1(n9493), .B2(n6087), .C1(
        P1_U3084), .C2(n6091), .ZN(P1_U3350) );
  AND2_X1 U7260 ( .A1(n6130), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5663) );
  INV_X1 U7261 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5669) );
  INV_X1 U7262 ( .A(n7400), .ZN(n5666) );
  NAND2_X1 U7263 ( .A1(n7272), .A2(P1_B_REG_SCAN_IN), .ZN(n5664) );
  MUX2_X1 U7264 ( .A(P1_B_REG_SCAN_IN), .B(n5664), .S(n7079), .Z(n5665) );
  AND2_X1 U7265 ( .A1(n7400), .A2(n7272), .ZN(n5667) );
  NAND2_X1 U7266 ( .A1(n6238), .A2(n9694), .ZN(n5668) );
  OAI21_X1 U7267 ( .B1(n9694), .B2(n5669), .A(n5668), .ZN(P1_U3441) );
  OAI222_X1 U7268 ( .A1(n8979), .A2(n5670), .B1(n8980), .B2(n6068), .C1(
        P2_U3152), .C2(n5803), .ZN(P2_U3353) );
  INV_X1 U7269 ( .A(n5830), .ZN(n5792) );
  OAI222_X1 U7270 ( .A1(n8979), .A2(n5671), .B1(n8980), .B2(n6119), .C1(
        P2_U3152), .C2(n5792), .ZN(P2_U3352) );
  OR2_X1 U7271 ( .A1(n5672), .A2(n9486), .ZN(n5673) );
  XNOR2_X1 U7272 ( .A(n5673), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9602) );
  OAI222_X1 U7273 ( .A1(n9495), .A2(n6053), .B1(n9493), .B2(n6052), .C1(
        P1_U3084), .C2(n6056), .ZN(P1_U3349) );
  NAND2_X1 U7274 ( .A1(n5672), .A2(n5674), .ZN(n5680) );
  NAND2_X1 U7275 ( .A1(n5680), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5675) );
  XNOR2_X1 U7276 ( .A(n5675), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6028) );
  INV_X1 U7277 ( .A(n6028), .ZN(n6123) );
  OAI222_X1 U7278 ( .A1(n9495), .A2(n6121), .B1(n9493), .B2(n6119), .C1(
        P1_U3084), .C2(n6123), .ZN(P1_U3347) );
  INV_X1 U7279 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7280 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5676) );
  OAI222_X1 U7281 ( .A1(n9495), .A2(n5945), .B1(n9493), .B2(n5943), .C1(
        P1_U3084), .C2(n5939), .ZN(P1_U3352) );
  INV_X1 U7282 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7283 ( .A1(n5672), .A2(n5677), .ZN(n5678) );
  NAND2_X1 U7284 ( .A1(n5678), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5679) );
  MUX2_X1 U7285 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5679), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5681) );
  INV_X1 U7286 ( .A(n5918), .ZN(n6070) );
  OAI222_X1 U7287 ( .A1(n9495), .A2(n6069), .B1(n9493), .B2(n6068), .C1(
        P1_U3084), .C2(n6070), .ZN(P1_U3348) );
  AND2_X1 U7288 ( .A1(n5672), .A2(n5682), .ZN(n5683) );
  INV_X1 U7289 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5685) );
  XNOR2_X1 U7290 ( .A(n5686), .B(n5685), .ZN(n6346) );
  OAI222_X1 U7291 ( .A1(n9495), .A2(n6288), .B1(n9493), .B2(n6287), .C1(
        P1_U3084), .C2(n6346), .ZN(P1_U3346) );
  INV_X1 U7292 ( .A(n6184), .ZN(n6191) );
  OAI222_X1 U7293 ( .A1(n8979), .A2(n5684), .B1(n8980), .B2(n6287), .C1(
        P2_U3152), .C2(n6191), .ZN(P2_U3351) );
  INV_X1 U7294 ( .A(n6642), .ZN(n5689) );
  NAND2_X1 U7295 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  NAND2_X1 U7296 ( .A1(n5687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5715) );
  XNOR2_X1 U7297 ( .A(n5715), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9628) );
  INV_X1 U7298 ( .A(n9495), .ZN(n9488) );
  AOI22_X1 U7299 ( .A1(n9628), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9488), .ZN(n5688) );
  OAI21_X1 U7300 ( .B1(n5689), .B2(n9493), .A(n5688), .ZN(P1_U3345) );
  INV_X1 U7301 ( .A(n6375), .ZN(n6382) );
  OAI222_X1 U7302 ( .A1(n8979), .A2(n5690), .B1(n8980), .B2(n5689), .C1(
        P2_U3152), .C2(n6382), .ZN(P2_U3350) );
  INV_X1 U7303 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5705) );
  NOR2_X1 U7304 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5691) );
  NAND2_X1 U7305 ( .A1(n5696), .A2(n5694), .ZN(n5698) );
  OR2_X1 U7306 ( .A1(n5696), .A2(n9486), .ZN(n5697) );
  INV_X2 U7307 ( .A(n7639), .ZN(n5707) );
  NAND2_X1 U7308 ( .A1(n7244), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7309 ( .A1(n7822), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U7310 ( .A1(n4305), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5701) );
  AND3_X1 U7311 ( .A1(n5703), .A2(n5702), .A3(n5701), .ZN(n7732) );
  INV_X1 U7312 ( .A(n7732), .ZN(n8119) );
  NAND2_X1 U7313 ( .A1(n8119), .A2(P1_U4006), .ZN(n5704) );
  OAI21_X1 U7314 ( .B1(P1_U4006), .B2(n5705), .A(n5704), .ZN(P1_U3586) );
  INV_X1 U7315 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U7316 ( .A1(n7346), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7317 ( .A1(n6114), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U7318 ( .A1(n5931), .A2(P1_U4006), .ZN(n5712) );
  OAI21_X1 U7319 ( .B1(P1_U4006), .B2(n9878), .A(n5712), .ZN(P1_U3555) );
  NAND2_X1 U7320 ( .A1(n8620), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5713) );
  OAI21_X1 U7321 ( .B1(n8858), .B2(n8620), .A(n5713), .ZN(P2_U3572) );
  INV_X1 U7322 ( .A(n6706), .ZN(n5719) );
  INV_X1 U7323 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7324 ( .A1(n5715), .A2(n5714), .ZN(n5716) );
  NAND2_X1 U7325 ( .A1(n5716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5717) );
  XNOR2_X1 U7326 ( .A(n5717), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9642) );
  AOI22_X1 U7327 ( .A1(n9642), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9488), .ZN(n5718) );
  OAI21_X1 U7328 ( .B1(n5719), .B2(n9493), .A(n5718), .ZN(P1_U3344) );
  INV_X1 U7329 ( .A(n6580), .ZN(n6388) );
  OAI222_X1 U7330 ( .A1(n8979), .A2(n5720), .B1(n8233), .B2(n5719), .C1(n6388), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI21_X1 U7331 ( .B1(n9754), .B2(n5721), .A(n5749), .ZN(n5724) );
  NAND2_X1 U7332 ( .A1(n5722), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8457) );
  NAND2_X1 U7333 ( .A1(n9754), .A2(n8457), .ZN(n5723) );
  NAND2_X1 U7334 ( .A1(n5724), .A2(n5723), .ZN(n8724) );
  NOR2_X1 U7335 ( .A1(n9729), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7336 ( .A(n5725), .ZN(n5731) );
  NAND2_X1 U7337 ( .A1(n5726), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5727) );
  MUX2_X1 U7338 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5727), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5728) );
  AND2_X1 U7339 ( .A1(n5728), .A2(n5576), .ZN(n9125) );
  AOI22_X1 U7340 ( .A1(n9125), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9488), .ZN(n5729) );
  OAI21_X1 U7341 ( .B1(n5731), .B2(n9493), .A(n5729), .ZN(P1_U3343) );
  INV_X1 U7342 ( .A(n6963), .ZN(n6588) );
  OAI222_X1 U7343 ( .A1(P2_U3152), .A2(n6588), .B1(n8980), .B2(n5731), .C1(
        n5730), .C2(n8979), .ZN(P2_U3348) );
  INV_X1 U7344 ( .A(n5732), .ZN(n5733) );
  INV_X1 U7345 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n5746) );
  NOR2_X1 U7346 ( .A1(n5734), .A2(P1_U3084), .ZN(n5742) );
  INV_X1 U7347 ( .A(n8117), .ZN(n5740) );
  NAND2_X1 U7348 ( .A1(n5742), .A2(n5740), .ZN(n9623) );
  INV_X1 U7349 ( .A(n5734), .ZN(n5737) );
  NAND4_X1 U7350 ( .A1(n5737), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .A4(n5973), .ZN(n5739) );
  OAI21_X1 U7351 ( .B1(n8117), .B2(P1_REG2_REG_0__SCAN_IN), .A(n5973), .ZN(
        n5738) );
  XOR2_X1 U7352 ( .A(P1_IR_REG_0__SCAN_IN), .B(n5738), .Z(n9583) );
  AOI21_X1 U7353 ( .B1(n9623), .B2(n5739), .A(n9583), .ZN(n5744) );
  OR2_X1 U7354 ( .A1(n5740), .A2(n5736), .ZN(n9585) );
  INV_X1 U7355 ( .A(n9585), .ZN(n5741) );
  INV_X1 U7356 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5905) );
  AND3_X1 U7357 ( .A1(n9686), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5905), .ZN(n5743) );
  AOI211_X1 U7358 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n5744), .B(
        n5743), .ZN(n5745) );
  OAI21_X1 U7359 ( .B1(n9671), .B2(n5746), .A(n5745), .ZN(P1_U3241) );
  OAI211_X1 U7360 ( .C1(n9754), .C2(n5748), .A(n8457), .B(n5747), .ZN(n5750)
         );
  NAND2_X1 U7361 ( .A1(n5750), .A2(n5749), .ZN(n5755) );
  NAND2_X1 U7362 ( .A1(n8620), .A2(n5755), .ZN(n5769) );
  NAND2_X1 U7363 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6810) );
  INV_X1 U7364 ( .A(n6810), .ZN(n5760) );
  INV_X1 U7365 ( .A(n5765), .ZN(n9513) );
  INV_X1 U7366 ( .A(n5764), .ZN(n9501) );
  NAND2_X1 U7367 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9499) );
  INV_X1 U7368 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5751) );
  INV_X1 U7369 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5752) );
  MUX2_X1 U7370 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5752), .S(n5765), .Z(n9510)
         );
  NOR2_X1 U7371 ( .A1(n9511), .A2(n9510), .ZN(n9509) );
  AOI21_X1 U7372 ( .B1(n9513), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9509), .ZN(
        n5806) );
  NAND2_X1 U7373 ( .A1(n5761), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5753) );
  OAI21_X1 U7374 ( .B1(n5761), .B2(P2_REG1_REG_3__SCAN_IN), .A(n5753), .ZN(
        n5805) );
  NOR2_X1 U7375 ( .A1(n5806), .A2(n5805), .ZN(n5804) );
  INV_X1 U7376 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5754) );
  MUX2_X1 U7377 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5754), .S(n5785), .Z(n5757)
         );
  INV_X1 U7378 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U7379 ( .A1(n5756), .A2(n5509), .ZN(n9732) );
  AOI211_X1 U7380 ( .C1(n5758), .C2(n5757), .A(n5774), .B(n9732), .ZN(n5759)
         );
  AOI211_X1 U7381 ( .C1(n9729), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n5760), .B(
        n5759), .ZN(n5773) );
  NAND2_X1 U7382 ( .A1(n5761), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5766) );
  MUX2_X1 U7383 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n5762), .S(n5761), .Z(n5810)
         );
  MUX2_X1 U7384 ( .A(n5763), .B(P2_REG2_REG_2__SCAN_IN), .S(n5765), .Z(n9516)
         );
  MUX2_X1 U7385 ( .A(n6215), .B(P2_REG2_REG_1__SCAN_IN), .S(n5764), .Z(n9504)
         );
  NAND3_X1 U7386 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9504), .ZN(n9503) );
  OAI21_X1 U7387 ( .B1(n5764), .B2(n6215), .A(n9503), .ZN(n9517) );
  NAND2_X1 U7388 ( .A1(n9516), .A2(n9517), .ZN(n9515) );
  OAI21_X1 U7389 ( .B1(n5765), .B2(n5763), .A(n9515), .ZN(n5811) );
  NAND2_X1 U7390 ( .A1(n5810), .A2(n5811), .ZN(n5809) );
  NAND2_X1 U7391 ( .A1(n5766), .A2(n5809), .ZN(n5771) );
  MUX2_X1 U7392 ( .A(n5767), .B(P2_REG2_REG_4__SCAN_IN), .S(n5785), .Z(n5770)
         );
  NOR2_X1 U7393 ( .A1(n5508), .A2(n5509), .ZN(n5768) );
  NAND2_X1 U7394 ( .A1(n5770), .A2(n5771), .ZN(n5784) );
  OAI211_X1 U7395 ( .C1(n5771), .C2(n5770), .A(n9728), .B(n5784), .ZN(n5772)
         );
  OAI211_X1 U7396 ( .C1(n9731), .C2(n5785), .A(n5773), .B(n5772), .ZN(P2_U3249) );
  NAND2_X1 U7397 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6629) );
  INV_X1 U7398 ( .A(n6629), .ZN(n5781) );
  INV_X1 U7399 ( .A(n5785), .ZN(n5775) );
  NAND2_X1 U7400 ( .A1(n5782), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5776) );
  OAI21_X1 U7401 ( .B1(n5782), .B2(P2_REG1_REG_5__SCAN_IN), .A(n5776), .ZN(
        n5794) );
  AOI21_X1 U7402 ( .B1(n5782), .B2(P2_REG1_REG_5__SCAN_IN), .A(n5793), .ZN(
        n5779) );
  NAND2_X1 U7403 ( .A1(n5830), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5777) );
  OAI21_X1 U7404 ( .B1(n5830), .B2(P2_REG1_REG_6__SCAN_IN), .A(n5777), .ZN(
        n5778) );
  NOR2_X1 U7405 ( .A1(n5779), .A2(n5778), .ZN(n5824) );
  AOI211_X1 U7406 ( .C1(n5779), .C2(n5778), .A(n5824), .B(n9732), .ZN(n5780)
         );
  AOI211_X1 U7407 ( .C1(n9729), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n5781), .B(
        n5780), .ZN(n5791) );
  NAND2_X1 U7408 ( .A1(n5782), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5786) );
  MUX2_X1 U7409 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n5783), .S(n5782), .Z(n5799)
         );
  OAI21_X1 U7410 ( .B1(n5785), .B2(n5767), .A(n5784), .ZN(n5800) );
  NAND2_X1 U7411 ( .A1(n5799), .A2(n5800), .ZN(n5798) );
  NAND2_X1 U7412 ( .A1(n5786), .A2(n5798), .ZN(n5789) );
  MUX2_X1 U7413 ( .A(n6402), .B(P2_REG2_REG_6__SCAN_IN), .S(n5830), .Z(n5787)
         );
  INV_X1 U7414 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U7415 ( .A1(n5788), .A2(n5789), .ZN(n5831) );
  OAI211_X1 U7416 ( .C1(n5789), .C2(n5788), .A(n9728), .B(n5831), .ZN(n5790)
         );
  OAI211_X1 U7417 ( .C1(n9731), .C2(n5792), .A(n5791), .B(n5790), .ZN(P2_U3251) );
  NAND2_X1 U7418 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n8217) );
  INV_X1 U7419 ( .A(n8217), .ZN(n5797) );
  AOI211_X1 U7420 ( .C1(n5795), .C2(n5794), .A(n5793), .B(n9732), .ZN(n5796)
         );
  AOI211_X1 U7421 ( .C1(n9729), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n5797), .B(
        n5796), .ZN(n5802) );
  OAI211_X1 U7422 ( .C1(n5800), .C2(n5799), .A(n9728), .B(n5798), .ZN(n5801)
         );
  OAI211_X1 U7423 ( .C1(n9731), .C2(n5803), .A(n5802), .B(n5801), .ZN(P2_U3250) );
  NOR2_X1 U7424 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4468), .ZN(n5808) );
  AOI211_X1 U7425 ( .C1(n5806), .C2(n5805), .A(n5804), .B(n9732), .ZN(n5807)
         );
  AOI211_X1 U7426 ( .C1(n9729), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n5808), .B(
        n5807), .ZN(n5813) );
  OAI211_X1 U7427 ( .C1(n5811), .C2(n5810), .A(n9728), .B(n5809), .ZN(n5812)
         );
  OAI211_X1 U7428 ( .C1(n9731), .C2(n5814), .A(n5813), .B(n5812), .ZN(P2_U3248) );
  INV_X1 U7429 ( .A(n6920), .ZN(n5821) );
  NAND2_X1 U7430 ( .A1(n5576), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5816) );
  MUX2_X1 U7431 ( .A(n5816), .B(P1_IR_REG_31__SCAN_IN), .S(n5815), .Z(n5819)
         );
  INV_X1 U7432 ( .A(n5817), .ZN(n5818) );
  INV_X1 U7433 ( .A(n9646), .ZN(n6333) );
  OAI222_X1 U7434 ( .A1(n9493), .A2(n5821), .B1(n6333), .B2(P1_U3084), .C1(
        n9865), .C2(n9495), .ZN(P1_U3342) );
  INV_X1 U7435 ( .A(n7054), .ZN(n6970) );
  OAI222_X1 U7436 ( .A1(P2_U3152), .A2(n6970), .B1(n8980), .B2(n5821), .C1(
        n5820), .C2(n8979), .ZN(P2_U3347) );
  NAND2_X1 U7437 ( .A1(n8620), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5822) );
  OAI21_X1 U7438 ( .B1(n8845), .B2(n8620), .A(n5822), .ZN(P2_U3575) );
  NOR2_X1 U7439 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5823), .ZN(n5829) );
  AOI21_X1 U7440 ( .B1(n5830), .B2(P2_REG1_REG_6__SCAN_IN), .A(n5824), .ZN(
        n5827) );
  INV_X1 U7441 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5825) );
  MUX2_X1 U7442 ( .A(n5825), .B(P2_REG1_REG_7__SCAN_IN), .S(n6184), .Z(n5826)
         );
  NOR2_X1 U7443 ( .A1(n5827), .A2(n5826), .ZN(n6183) );
  AOI211_X1 U7444 ( .C1(n5827), .C2(n5826), .A(n6183), .B(n9732), .ZN(n5828)
         );
  AOI211_X1 U7445 ( .C1(n9729), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n5829), .B(
        n5828), .ZN(n5836) );
  NAND2_X1 U7446 ( .A1(n5830), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7447 ( .A1(n5832), .A2(n5831), .ZN(n5834) );
  MUX2_X1 U7448 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6507), .S(n6184), .Z(n5833)
         );
  NAND2_X1 U7449 ( .A1(n5833), .A2(n5834), .ZN(n6190) );
  OAI211_X1 U7450 ( .C1(n5834), .C2(n5833), .A(n9728), .B(n6190), .ZN(n5835)
         );
  OAI211_X1 U7451 ( .C1(n9731), .C2(n6191), .A(n5836), .B(n5835), .ZN(P2_U3252) );
  INV_X1 U7452 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9972) );
  NOR2_X1 U7453 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9972), .ZN(n6170) );
  INV_X1 U7454 ( .A(n9591), .ZN(n5839) );
  INV_X1 U7455 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5837) );
  MUX2_X1 U7456 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n5837), .S(n5939), .Z(n9570)
         );
  NOR3_X1 U7457 ( .A1(n4528), .A2(n5905), .A3(n9570), .ZN(n9569) );
  AOI21_X1 U7458 ( .B1(n5940), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9569), .ZN(
        n9582) );
  INV_X1 U7459 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5838) );
  MUX2_X1 U7460 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n5838), .S(n9591), .Z(n9581)
         );
  NAND2_X1 U7461 ( .A1(n5861), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5840) );
  OAI21_X1 U7462 ( .B1(n5861), .B2(P1_REG1_REG_3__SCAN_IN), .A(n5840), .ZN(
        n5841) );
  NOR2_X1 U7463 ( .A1(n5842), .A2(n5841), .ZN(n5855) );
  AOI211_X1 U7464 ( .C1(n5842), .C2(n5841), .A(n5855), .B(n9579), .ZN(n5843)
         );
  AOI211_X1 U7465 ( .C1(n9685), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n6170), .B(
        n5843), .ZN(n5852) );
  INV_X1 U7466 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5845) );
  MUX2_X1 U7467 ( .A(n5845), .B(P1_REG2_REG_2__SCAN_IN), .S(n9591), .Z(n9589)
         );
  INV_X1 U7468 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5844) );
  NAND3_X1 U7469 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .A3(n9574), .ZN(n9573) );
  OAI21_X1 U7470 ( .B1(n5939), .B2(n5844), .A(n9573), .ZN(n9588) );
  NAND2_X1 U7471 ( .A1(n9589), .A2(n9588), .ZN(n9587) );
  OAI21_X1 U7472 ( .B1(n9591), .B2(n5845), .A(n9587), .ZN(n5850) );
  INV_X1 U7473 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5846) );
  INV_X1 U7474 ( .A(n5847), .ZN(n5849) );
  OAI211_X1 U7475 ( .C1(n5850), .C2(n5849), .A(n9676), .B(n5862), .ZN(n5851)
         );
  OAI211_X1 U7476 ( .C1(n9592), .C2(n6091), .A(n5852), .B(n5851), .ZN(P1_U3244) );
  NOR2_X1 U7477 ( .A1(n6028), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5853) );
  AOI21_X1 U7478 ( .B1(n6028), .B2(P1_REG1_REG_6__SCAN_IN), .A(n5853), .ZN(
        n5857) );
  NAND2_X1 U7479 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n5918), .ZN(n5854) );
  OAI21_X1 U7480 ( .B1(n5918), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5854), .ZN(
        n5915) );
  INV_X1 U7481 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6535) );
  AOI22_X1 U7482 ( .A1(n9602), .A2(P1_REG1_REG_4__SCAN_IN), .B1(n6535), .B2(
        n6056), .ZN(n9605) );
  AOI21_X1 U7483 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n5861), .A(n5855), .ZN(
        n9604) );
  NAND2_X1 U7484 ( .A1(n9605), .A2(n9604), .ZN(n9603) );
  OAI21_X1 U7485 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9602), .A(n9603), .ZN(
        n5916) );
  NOR2_X1 U7486 ( .A1(n5915), .A2(n5916), .ZN(n5914) );
  AOI21_X1 U7487 ( .B1(n5918), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5914), .ZN(
        n5856) );
  NAND2_X1 U7488 ( .A1(n5856), .A2(n5857), .ZN(n6027) );
  OAI21_X1 U7489 ( .B1(n5857), .B2(n5856), .A(n6027), .ZN(n5860) );
  AND2_X1 U7490 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6146) );
  INV_X1 U7491 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n5858) );
  NOR2_X1 U7492 ( .A1(n9671), .A2(n5858), .ZN(n5859) );
  AOI211_X1 U7493 ( .C1(n9686), .C2(n5860), .A(n6146), .B(n5859), .ZN(n5873)
         );
  NOR2_X1 U7494 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n5918), .ZN(n5867) );
  NAND2_X1 U7495 ( .A1(n5861), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5863) );
  INV_X1 U7496 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5864) );
  NOR2_X1 U7497 ( .A1(n9602), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5865) );
  INV_X1 U7498 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5866) );
  MUX2_X1 U7499 ( .A(n5866), .B(P1_REG2_REG_5__SCAN_IN), .S(n5918), .Z(n5912)
         );
  NOR2_X1 U7500 ( .A1(n5867), .A2(n5911), .ZN(n5871) );
  INV_X1 U7501 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5868) );
  MUX2_X1 U7502 ( .A(n5868), .B(P1_REG2_REG_6__SCAN_IN), .S(n6028), .Z(n5869)
         );
  INV_X1 U7503 ( .A(n5869), .ZN(n5870) );
  NAND2_X1 U7504 ( .A1(n5871), .A2(n5870), .ZN(n6020) );
  OAI211_X1 U7505 ( .C1(n5871), .C2(n5870), .A(n9676), .B(n6020), .ZN(n5872)
         );
  OAI211_X1 U7506 ( .C1(n9592), .C2(n6123), .A(n5873), .B(n5872), .ZN(P1_U3247) );
  NOR4_X1 U7507 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5882) );
  NOR4_X1 U7508 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5881) );
  NOR4_X1 U7509 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5877) );
  NOR4_X1 U7510 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5876) );
  NOR4_X1 U7511 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5875) );
  NOR4_X1 U7512 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5874) );
  NAND4_X1 U7513 ( .A1(n5877), .A2(n5876), .A3(n5875), .A4(n5874), .ZN(n5878)
         );
  NOR4_X1 U7514 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5879), .A4(n5878), .ZN(n5880) );
  NAND3_X1 U7515 ( .A1(n5882), .A2(n5881), .A3(n5880), .ZN(n5883) );
  NAND2_X1 U7516 ( .A1(n9690), .A2(n5883), .ZN(n6237) );
  INV_X1 U7517 ( .A(n6237), .ZN(n5884) );
  NOR2_X1 U7518 ( .A1(n6238), .A2(n5884), .ZN(n5891) );
  NAND2_X1 U7519 ( .A1(n5887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5889) );
  OR2_X1 U7520 ( .A1(n9696), .A2(n8097), .ZN(n5890) );
  INV_X1 U7521 ( .A(n6131), .ZN(n5893) );
  INV_X1 U7522 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9990) );
  AND2_X1 U7523 ( .A1(n7400), .A2(n7079), .ZN(n5892) );
  AOI21_X1 U7524 ( .B1(n9690), .B2(n9990), .A(n5892), .ZN(n5959) );
  NAND2_X1 U7525 ( .A1(n5959), .A2(n9694), .ZN(n9693) );
  INV_X1 U7526 ( .A(SI_0_), .ZN(n5896) );
  INV_X1 U7527 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5895) );
  OAI21_X1 U7528 ( .B1(n7725), .B2(n5896), .A(n5895), .ZN(n5898) );
  AND2_X1 U7529 ( .A1(n5898), .A2(n5897), .ZN(n9496) );
  AND2_X1 U7530 ( .A1(n5923), .A2(n5931), .ZN(n7840) );
  NOR2_X1 U7531 ( .A1(n5923), .A2(n5931), .ZN(n6159) );
  OR2_X1 U7532 ( .A1(n7840), .A2(n6159), .ZN(n8030) );
  NAND2_X1 U7533 ( .A1(n8109), .A2(n8097), .ZN(n6000) );
  OR2_X1 U7534 ( .A1(n6000), .A2(n5925), .ZN(n8108) );
  AND2_X1 U7535 ( .A1(n8108), .A2(n5963), .ZN(n5903) );
  NAND2_X1 U7536 ( .A1(n6114), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5901) );
  AND2_X1 U7537 ( .A1(n9372), .A2(n9120), .ZN(n5902) );
  AOI21_X1 U7538 ( .B1(n8030), .B2(n5903), .A(n5902), .ZN(n6286) );
  OAI21_X1 U7539 ( .B1(n5923), .B2(n5963), .A(n6286), .ZN(n5908) );
  NAND2_X1 U7540 ( .A1(n5908), .A2(n9561), .ZN(n5904) );
  OAI21_X1 U7541 ( .B1(n9561), .B2(n5905), .A(n5904), .ZN(P1_U3523) );
  NOR2_X1 U7542 ( .A1(n5959), .A2(n8107), .ZN(n5906) );
  INV_X1 U7543 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7544 ( .A1(n5908), .A2(n9719), .ZN(n5909) );
  OAI21_X1 U7545 ( .B1(n9719), .B2(n5910), .A(n5909), .ZN(P1_U3454) );
  AOI21_X1 U7546 ( .B1(n5913), .B2(n5912), .A(n5911), .ZN(n5921) );
  INV_X1 U7547 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6072) );
  NOR2_X1 U7548 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6072), .ZN(n6267) );
  AOI211_X1 U7549 ( .C1(n5916), .C2(n5915), .A(n5914), .B(n9579), .ZN(n5917)
         );
  AOI211_X1 U7550 ( .C1(n9685), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n6267), .B(
        n5917), .ZN(n5920) );
  NAND2_X1 U7551 ( .A1(n9678), .A2(n5918), .ZN(n5919) );
  OAI211_X1 U7552 ( .C1(n5921), .C2(n9637), .A(n5920), .B(n5919), .ZN(P1_U3246) );
  NAND2_X1 U7553 ( .A1(n5932), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5922) );
  OAI21_X1 U7554 ( .B1(n5923), .B2(n5938), .A(n5922), .ZN(n5924) );
  INV_X1 U7555 ( .A(n5924), .ZN(n5927) );
  INV_X1 U7556 ( .A(n5925), .ZN(n6232) );
  AND2_X2 U7557 ( .A1(n6232), .A2(n6132), .ZN(n6092) );
  INV_X1 U7558 ( .A(n7685), .ZN(n5928) );
  NAND2_X1 U7559 ( .A1(n5928), .A2(n6095), .ZN(n5937) );
  AND2_X4 U7560 ( .A1(n5930), .A2(n6001), .ZN(n9002) );
  NAND2_X1 U7561 ( .A1(n7684), .A2(n6092), .ZN(n5934) );
  NAND2_X1 U7562 ( .A1(n5932), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7563 ( .A1(n7687), .A2(n7685), .ZN(n7686) );
  NAND2_X1 U7564 ( .A1(n5937), .A2(n7686), .ZN(n5955) );
  INV_X1 U7565 ( .A(n5955), .ZN(n5953) );
  NAND2_X2 U7566 ( .A1(n5944), .A2(n5942), .ZN(n6067) );
  OR2_X1 U7567 ( .A1(n6067), .A2(n5943), .ZN(n5947) );
  NAND2_X2 U7568 ( .A1(n5944), .A2(n7725), .ZN(n6120) );
  OR2_X1 U7569 ( .A1(n4306), .A2(n5945), .ZN(n5946) );
  NAND2_X1 U7570 ( .A1(n5930), .A2(n6012), .ZN(n5950) );
  NAND2_X1 U7571 ( .A1(n9120), .A2(n6092), .ZN(n5949) );
  NAND2_X1 U7572 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  XNOR2_X1 U7573 ( .A(n5951), .B(n8482), .ZN(n5954) );
  INV_X1 U7574 ( .A(n5954), .ZN(n5952) );
  NAND2_X1 U7575 ( .A1(n5953), .A2(n5952), .ZN(n6038) );
  NAND2_X1 U7576 ( .A1(n5955), .A2(n5954), .ZN(n6039) );
  NAND2_X1 U7577 ( .A1(n6038), .A2(n6039), .ZN(n5958) );
  NAND2_X1 U7578 ( .A1(n9002), .A2(n9120), .ZN(n5957) );
  NAND2_X1 U7579 ( .A1(n6012), .A2(n6092), .ZN(n5956) );
  AND2_X1 U7580 ( .A1(n5957), .A2(n5956), .ZN(n6037) );
  XNOR2_X1 U7581 ( .A(n5958), .B(n6037), .ZN(n5977) );
  NAND3_X1 U7582 ( .A1(n6238), .A2(n5959), .A3(n6237), .ZN(n5965) );
  INV_X1 U7583 ( .A(n5968), .ZN(n5962) );
  AND2_X1 U7584 ( .A1(n9710), .A2(n8061), .ZN(n5961) );
  OR2_X1 U7585 ( .A1(n5963), .A2(n5899), .ZN(n6276) );
  NOR2_X1 U7586 ( .A1(n6276), .A2(n8107), .ZN(n5964) );
  AND2_X1 U7587 ( .A1(n5964), .A2(n5965), .ZN(n6135) );
  INV_X1 U7588 ( .A(n6135), .ZN(n5966) );
  NAND2_X1 U7589 ( .A1(n5965), .A2(n9710), .ZN(n6134) );
  NAND4_X1 U7590 ( .A1(n5966), .A2(n9694), .A3(n6131), .A4(n6134), .ZN(n9072)
         );
  NAND2_X1 U7591 ( .A1(n9694), .A2(n9178), .ZN(n5967) );
  OAI21_X2 U7592 ( .B1(n5968), .B2(n6276), .A(n9365), .ZN(n9084) );
  AOI22_X1 U7593 ( .A1(n9072), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9084), .B2(
        n6012), .ZN(n5976) );
  NOR2_X1 U7594 ( .A1(n5968), .A2(n8108), .ZN(n5974) );
  NAND2_X1 U7595 ( .A1(n7346), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7596 ( .A1(n7869), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7597 ( .A1(n6114), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7598 ( .A1(n7244), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5969) );
  NAND4_X2 U7599 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(n9118)
         );
  AOI22_X1 U7600 ( .A1(n9073), .A2(n9118), .B1(n9092), .B2(n5931), .ZN(n5975)
         );
  OAI211_X1 U7601 ( .C1(n5977), .C2(n9086), .A(n5976), .B(n5975), .ZN(P1_U3220) );
  INV_X1 U7602 ( .A(n7023), .ZN(n5983) );
  NOR2_X1 U7603 ( .A1(n5817), .A2(n9486), .ZN(n5978) );
  MUX2_X1 U7604 ( .A(n9486), .B(n5978), .S(P1_IR_REG_12__SCAN_IN), .Z(n5981)
         );
  INV_X1 U7605 ( .A(n5979), .ZN(n5980) );
  OAI222_X1 U7606 ( .A1(n9495), .A2(n5982), .B1(n9493), .B2(n5983), .C1(
        P1_U3084), .C2(n6349), .ZN(P1_U3341) );
  INV_X1 U7607 ( .A(n7222), .ZN(n7065) );
  OAI222_X1 U7608 ( .A1(n8979), .A2(n5984), .B1(n8980), .B2(n5983), .C1(
        P2_U3152), .C2(n7065), .ZN(P2_U3346) );
  INV_X1 U7609 ( .A(n7138), .ZN(n6035) );
  NAND2_X1 U7610 ( .A1(n5979), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7611 ( .A(n5985), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7313) );
  AOI22_X1 U7612 ( .A1(n7313), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9488), .ZN(n5986) );
  OAI21_X1 U7613 ( .B1(n6035), .B2(n9493), .A(n5986), .ZN(P1_U3340) );
  INV_X1 U7614 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6017) );
  AND2_X1 U7615 ( .A1(n5931), .A2(n7684), .ZN(n6157) );
  NAND2_X1 U7616 ( .A1(n6158), .A2(n6157), .ZN(n6156) );
  NAND2_X1 U7617 ( .A1(n9120), .A2(n6012), .ZN(n5987) );
  NAND2_X1 U7618 ( .A1(n6156), .A2(n5987), .ZN(n5993) );
  INV_X1 U7619 ( .A(n5993), .ZN(n5992) );
  OR2_X1 U7620 ( .A1(n6120), .A2(n5989), .ZN(n5990) );
  INV_X1 U7621 ( .A(n8033), .ZN(n5999) );
  NAND2_X1 U7622 ( .A1(n5992), .A2(n5999), .ZN(n6416) );
  NAND2_X1 U7623 ( .A1(n5993), .A2(n8033), .ZN(n5994) );
  NAND2_X1 U7624 ( .A1(n6416), .A2(n5994), .ZN(n6004) );
  INV_X1 U7625 ( .A(n6004), .ZN(n6283) );
  NAND2_X1 U7626 ( .A1(n5929), .A2(n9178), .ZN(n8016) );
  OR2_X1 U7627 ( .A1(n5929), .A2(n8097), .ZN(n5996) );
  NAND2_X1 U7628 ( .A1(n5900), .A2(n8104), .ZN(n5995) );
  INV_X1 U7629 ( .A(n6158), .ZN(n8032) );
  NAND2_X1 U7630 ( .A1(n8032), .A2(n6159), .ZN(n5998) );
  INV_X1 U7631 ( .A(n9120), .ZN(n7690) );
  NAND2_X1 U7632 ( .A1(n7690), .A2(n6012), .ZN(n5997) );
  XNOR2_X1 U7633 ( .A(n6408), .B(n5999), .ZN(n6011) );
  OR2_X1 U7634 ( .A1(n6000), .A2(n6232), .ZN(n6003) );
  OR2_X1 U7635 ( .A1(n6001), .A2(n8092), .ZN(n6002) );
  AND2_X1 U7636 ( .A1(n6003), .A2(n6002), .ZN(n7354) );
  NAND2_X1 U7637 ( .A1(n6004), .A2(n7158), .ZN(n6010) );
  NAND2_X1 U7638 ( .A1(n4305), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7639 ( .A1(n7244), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7640 ( .A1(n6114), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7641 ( .A1(n7346), .A2(n9972), .ZN(n6005) );
  AOI22_X1 U7642 ( .A1(n9380), .A2(n9120), .B1(n9372), .B2(n9117), .ZN(n6009)
         );
  OAI211_X1 U7643 ( .C1(n9374), .C2(n6011), .A(n6010), .B(n6009), .ZN(n6274)
         );
  INV_X1 U7644 ( .A(n6274), .ZN(n6015) );
  AND2_X1 U7645 ( .A1(n6161), .A2(n4307), .ZN(n6013) );
  NOR2_X1 U7646 ( .A1(n6432), .A2(n6013), .ZN(n6280) );
  AOI22_X1 U7647 ( .A1(n6280), .A2(n9437), .B1(n9465), .B2(n4307), .ZN(n6014)
         );
  OAI211_X1 U7648 ( .C1(n6283), .C2(n9535), .A(n6015), .B(n6014), .ZN(n6018)
         );
  NAND2_X1 U7649 ( .A1(n6018), .A2(n9719), .ZN(n6016) );
  OAI21_X1 U7650 ( .B1(n9719), .B2(n6017), .A(n6016), .ZN(P1_U3460) );
  NAND2_X1 U7651 ( .A1(n6018), .A2(n9561), .ZN(n6019) );
  OAI21_X1 U7652 ( .B1(n9561), .B2(n5838), .A(n6019), .ZN(P1_U3525) );
  INV_X1 U7653 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7654 ( .A1(n6028), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7655 ( .A1(n6021), .A2(n6020), .ZN(n6024) );
  INV_X1 U7656 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6022) );
  MUX2_X1 U7657 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6022), .S(n6346), .Z(n6023)
         );
  AOI21_X1 U7658 ( .B1(n6024), .B2(n6023), .A(n6345), .ZN(n6025) );
  OAI22_X1 U7659 ( .A1(n6025), .A2(n9637), .B1(n9592), .B2(n6346), .ZN(n6026)
         );
  INV_X1 U7660 ( .A(n6026), .ZN(n6033) );
  INV_X1 U7661 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6336) );
  MUX2_X1 U7662 ( .A(n6336), .B(P1_REG1_REG_7__SCAN_IN), .S(n6346), .Z(n6030)
         );
  OAI21_X1 U7663 ( .B1(n6028), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6027), .ZN(
        n6029) );
  NAND2_X1 U7664 ( .A1(n6030), .A2(n6029), .ZN(n6337) );
  OAI21_X1 U7665 ( .B1(n6030), .B2(n6029), .A(n6337), .ZN(n6031) );
  INV_X1 U7666 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6138) );
  NOR2_X1 U7667 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6138), .ZN(n6314) );
  AOI21_X1 U7668 ( .B1(n9686), .B2(n6031), .A(n6314), .ZN(n6032) );
  OAI211_X1 U7669 ( .C1(n9671), .C2(n6034), .A(n6033), .B(n6032), .ZN(P1_U3248) );
  INV_X1 U7670 ( .A(n7409), .ZN(n7402) );
  OAI222_X1 U7671 ( .A1(n8979), .A2(n6036), .B1(n8233), .B2(n6035), .C1(n7402), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  NAND2_X1 U7672 ( .A1(n6038), .A2(n6037), .ZN(n6040) );
  NAND2_X1 U7673 ( .A1(n6040), .A2(n6039), .ZN(n9067) );
  NAND2_X1 U7674 ( .A1(n4307), .A2(n5930), .ZN(n6042) );
  NAND2_X1 U7675 ( .A1(n9118), .A2(n6092), .ZN(n6041) );
  NAND2_X1 U7676 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  XNOR2_X1 U7677 ( .A(n6043), .B(n8482), .ZN(n6046) );
  NAND2_X1 U7678 ( .A1(n9002), .A2(n9118), .ZN(n6045) );
  NAND2_X1 U7679 ( .A1(n4307), .A2(n6092), .ZN(n6044) );
  AND2_X1 U7680 ( .A1(n6045), .A2(n6044), .ZN(n6047) );
  NAND2_X1 U7681 ( .A1(n6046), .A2(n6047), .ZN(n6051) );
  INV_X1 U7682 ( .A(n6046), .ZN(n6049) );
  INV_X1 U7683 ( .A(n6047), .ZN(n6048) );
  NAND2_X1 U7684 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  AND2_X1 U7685 ( .A1(n6051), .A2(n6050), .ZN(n9069) );
  NAND2_X1 U7686 ( .A1(n9067), .A2(n9069), .ZN(n9068) );
  NAND2_X1 U7687 ( .A1(n9068), .A2(n6051), .ZN(n6167) );
  OR2_X1 U7688 ( .A1(n6067), .A2(n6052), .ZN(n6055) );
  OR2_X1 U7689 ( .A1(n6120), .A2(n6053), .ZN(n6054) );
  NAND2_X1 U7690 ( .A1(n6526), .A2(n5930), .ZN(n6063) );
  NAND2_X1 U7691 ( .A1(n7244), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7692 ( .A1(n7869), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7693 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6073) );
  OAI21_X1 U7694 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n6073), .ZN(n6057) );
  INV_X1 U7695 ( .A(n6057), .ZN(n6464) );
  NAND2_X1 U7696 ( .A1(n7346), .A2(n6464), .ZN(n6059) );
  NAND2_X1 U7697 ( .A1(n6114), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7698 ( .A1(n9116), .A2(n6092), .ZN(n6062) );
  NAND2_X1 U7699 ( .A1(n6063), .A2(n6062), .ZN(n6064) );
  XNOR2_X1 U7700 ( .A(n6064), .B(n8482), .ZN(n6101) );
  NAND2_X1 U7701 ( .A1(n9002), .A2(n9116), .ZN(n6066) );
  NAND2_X1 U7702 ( .A1(n6526), .A2(n6092), .ZN(n6065) );
  AND2_X1 U7703 ( .A1(n6066), .A2(n6065), .ZN(n6100) );
  OR2_X1 U7704 ( .A1(n6101), .A2(n6100), .ZN(n6259) );
  NAND2_X1 U7705 ( .A1(n6488), .A2(n5930), .ZN(n6080) );
  NAND2_X1 U7706 ( .A1(n7244), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7707 ( .A1(n7869), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6077) );
  INV_X1 U7708 ( .A(n6073), .ZN(n6071) );
  NAND2_X1 U7709 ( .A1(n6071), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7710 ( .A1(n6073), .A2(n6072), .ZN(n6074) );
  AND2_X1 U7711 ( .A1(n6112), .A2(n6074), .ZN(n6424) );
  NAND2_X1 U7712 ( .A1(n7346), .A2(n6424), .ZN(n6076) );
  NAND2_X1 U7713 ( .A1(n6114), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7714 ( .A1(n9115), .A2(n6092), .ZN(n6079) );
  NAND2_X1 U7715 ( .A1(n9002), .A2(n9115), .ZN(n6083) );
  NAND2_X1 U7716 ( .A1(n6488), .A2(n6092), .ZN(n6082) );
  NAND2_X1 U7717 ( .A1(n6083), .A2(n6082), .ZN(n6261) );
  NAND2_X1 U7718 ( .A1(n6263), .A2(n6261), .ZN(n6084) );
  NAND2_X1 U7719 ( .A1(n6259), .A2(n6084), .ZN(n6086) );
  NOR2_X1 U7720 ( .A1(n6263), .A2(n6261), .ZN(n6102) );
  INV_X1 U7721 ( .A(n6102), .ZN(n6085) );
  NAND2_X1 U7722 ( .A1(n6086), .A2(n6085), .ZN(n6107) );
  OR2_X1 U7723 ( .A1(n6067), .A2(n6087), .ZN(n6090) );
  OR2_X1 U7724 ( .A1(n6120), .A2(n6088), .ZN(n6089) );
  OAI211_X1 U7725 ( .C1(n5944), .C2(n6091), .A(n6090), .B(n6089), .ZN(n6169)
         );
  NAND2_X1 U7726 ( .A1(n6169), .A2(n5930), .ZN(n6094) );
  NAND2_X1 U7727 ( .A1(n9117), .A2(n6092), .ZN(n6093) );
  NAND2_X1 U7728 ( .A1(n6094), .A2(n6093), .ZN(n6096) );
  XNOR2_X1 U7729 ( .A(n6096), .B(n8482), .ZN(n6105) );
  NAND2_X1 U7730 ( .A1(n9002), .A2(n9117), .ZN(n6098) );
  NAND2_X1 U7731 ( .A1(n6169), .A2(n6092), .ZN(n6097) );
  NAND2_X1 U7732 ( .A1(n6098), .A2(n6097), .ZN(n6103) );
  XNOR2_X1 U7733 ( .A(n6105), .B(n6103), .ZN(n6168) );
  NAND2_X1 U7734 ( .A1(n6167), .A2(n6099), .ZN(n6109) );
  AND2_X1 U7735 ( .A1(n6101), .A2(n6100), .ZN(n6257) );
  NOR2_X1 U7736 ( .A1(n6102), .A2(n6257), .ZN(n6106) );
  INV_X1 U7737 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7738 ( .A1(n6105), .A2(n6104), .ZN(n6197) );
  NAND2_X1 U7739 ( .A1(n6109), .A2(n6108), .ZN(n6292) );
  NAND2_X1 U7740 ( .A1(n7869), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7741 ( .A1(n7244), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6117) );
  INV_X1 U7742 ( .A(n6112), .ZN(n6110) );
  NAND2_X1 U7743 ( .A1(n6110), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6139) );
  INV_X1 U7744 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7745 ( .A1(n6112), .A2(n6111), .ZN(n6113) );
  AND2_X1 U7746 ( .A1(n6139), .A2(n6113), .ZN(n6501) );
  NAND2_X1 U7747 ( .A1(n7346), .A2(n6501), .ZN(n6116) );
  NAND2_X1 U7748 ( .A1(n6114), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6115) );
  NAND4_X1 U7749 ( .A1(n6118), .A2(n6117), .A3(n6116), .A4(n6115), .ZN(n9114)
         );
  NAND2_X1 U7750 ( .A1(n9002), .A2(n9114), .ZN(n6125) );
  OR2_X1 U7751 ( .A1(n6120), .A2(n6121), .ZN(n6122) );
  NAND2_X1 U7752 ( .A1(n6515), .A2(n8508), .ZN(n6124) );
  NAND2_X1 U7753 ( .A1(n6125), .A2(n6124), .ZN(n6291) );
  NAND2_X1 U7754 ( .A1(n9114), .A2(n8508), .ZN(n6127) );
  NAND2_X1 U7755 ( .A1(n6515), .A2(n5930), .ZN(n6126) );
  NAND2_X1 U7756 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  XNOR2_X1 U7757 ( .A(n6128), .B(n8482), .ZN(n6293) );
  XOR2_X1 U7758 ( .A(n6291), .B(n6293), .Z(n6129) );
  XNOR2_X1 U7759 ( .A(n6292), .B(n6129), .ZN(n6149) );
  AOI22_X1 U7760 ( .A1(n9092), .A2(n9115), .B1(n6515), .B2(n9084), .ZN(n6148)
         );
  AND3_X1 U7761 ( .A1(n6132), .A2(n6131), .A3(n6130), .ZN(n6133) );
  AOI21_X1 U7762 ( .B1(n6134), .B2(n6133), .A(P1_U3084), .ZN(n6136) );
  NAND2_X1 U7763 ( .A1(n7244), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7764 ( .A1(n7869), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6143) );
  INV_X1 U7765 ( .A(n6139), .ZN(n6137) );
  NAND2_X1 U7766 ( .A1(n6137), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7767 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  AND2_X1 U7768 ( .A1(n6306), .A2(n6140), .ZN(n6696) );
  NAND2_X1 U7769 ( .A1(n7346), .A2(n6696), .ZN(n6142) );
  NAND2_X1 U7770 ( .A1(n7822), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6141) );
  NAND4_X1 U7771 ( .A1(n6144), .A2(n6143), .A3(n6142), .A4(n6141), .ZN(n9113)
         );
  INV_X1 U7772 ( .A(n9113), .ZN(n6678) );
  NOR2_X1 U7773 ( .A1(n9095), .A2(n6678), .ZN(n6145) );
  AOI211_X1 U7774 ( .C1(n6501), .C2(n9099), .A(n6146), .B(n6145), .ZN(n6147)
         );
  OAI211_X1 U7775 ( .C1(n6149), .C2(n9086), .A(n6148), .B(n6147), .ZN(P1_U3237) );
  INV_X1 U7776 ( .A(n7338), .ZN(n6179) );
  AOI22_X1 U7777 ( .A1(n8667), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n6150), .ZN(n6151) );
  OAI21_X1 U7778 ( .B1(n6179), .B2(n8980), .A(n6151), .ZN(P2_U3343) );
  INV_X1 U7779 ( .A(n7233), .ZN(n6182) );
  OR2_X1 U7780 ( .A1(n5979), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7781 ( .A1(n6152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6224) );
  OR2_X1 U7782 ( .A1(n6224), .A2(n6153), .ZN(n6154) );
  NAND2_X1 U7783 ( .A1(n6224), .A2(n6153), .ZN(n6176) );
  OAI222_X1 U7784 ( .A1(n9493), .A2(n6182), .B1(n7311), .B2(P1_U3084), .C1(
        n6155), .C2(n9495), .ZN(P1_U3339) );
  OAI21_X1 U7785 ( .B1(n6158), .B2(n6157), .A(n6156), .ZN(n6233) );
  XNOR2_X1 U7786 ( .A(n8032), .B(n6159), .ZN(n6160) );
  AOI222_X1 U7787 ( .A1(n9355), .A2(n6160), .B1(n9118), .B2(n9372), .C1(n5931), 
        .C2(n9380), .ZN(n6231) );
  INV_X1 U7788 ( .A(n6161), .ZN(n6162) );
  AOI211_X1 U7789 ( .C1(n7684), .C2(n6012), .A(n9696), .B(n6162), .ZN(n6242)
         );
  AOI21_X1 U7790 ( .B1(n9465), .B2(n6012), .A(n6242), .ZN(n6163) );
  OAI211_X1 U7791 ( .C1(n9468), .C2(n6233), .A(n6231), .B(n6163), .ZN(n6165)
         );
  NAND2_X1 U7792 ( .A1(n6165), .A2(n9719), .ZN(n6164) );
  OAI21_X1 U7793 ( .B1(n9719), .B2(n4677), .A(n6164), .ZN(P1_U3457) );
  NAND2_X1 U7794 ( .A1(n6165), .A2(n9561), .ZN(n6166) );
  OAI21_X1 U7795 ( .B1(n9561), .B2(n5837), .A(n6166), .ZN(P1_U3524) );
  NAND2_X1 U7796 ( .A1(n6167), .A2(n6168), .ZN(n6198) );
  OAI21_X1 U7797 ( .B1(n6168), .B2(n6167), .A(n6198), .ZN(n6174) );
  AOI22_X1 U7798 ( .A1(n9073), .A2(n9116), .B1(n9092), .B2(n9118), .ZN(n6172)
         );
  AOI21_X1 U7799 ( .B1(n9084), .B2(n6169), .A(n6170), .ZN(n6171) );
  OAI211_X1 U7800 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9050), .A(n6172), .B(
        n6171), .ZN(n6173) );
  AOI21_X1 U7801 ( .B1(n6174), .B2(n9088), .A(n6173), .ZN(n6175) );
  INV_X1 U7802 ( .A(n6175), .ZN(P1_U3216) );
  NAND2_X1 U7803 ( .A1(n6176), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6178) );
  XNOR2_X1 U7804 ( .A(n6178), .B(n6177), .ZN(n9141) );
  OAI222_X1 U7805 ( .A1(n9495), .A2(n6180), .B1(n9493), .B2(n6179), .C1(
        P1_U3084), .C2(n9141), .ZN(P1_U3338) );
  INV_X1 U7806 ( .A(n7407), .ZN(n8646) );
  OAI222_X1 U7807 ( .A1(P2_U3152), .A2(n8646), .B1(n8233), .B2(n6182), .C1(
        n6181), .C2(n8979), .ZN(P2_U3344) );
  NAND2_X1 U7808 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6739) );
  INV_X1 U7809 ( .A(n6739), .ZN(n6189) );
  AOI21_X1 U7810 ( .B1(n6184), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6183), .ZN(
        n6187) );
  INV_X1 U7811 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6185) );
  MUX2_X1 U7812 ( .A(n6185), .B(P2_REG1_REG_8__SCAN_IN), .S(n6375), .Z(n6186)
         );
  AOI211_X1 U7813 ( .C1(n6187), .C2(n6186), .A(n6374), .B(n9732), .ZN(n6188)
         );
  AOI211_X1 U7814 ( .C1(n9729), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6189), .B(
        n6188), .ZN(n6195) );
  OAI21_X1 U7815 ( .B1(n6191), .B2(n6507), .A(n6190), .ZN(n6193) );
  MUX2_X1 U7816 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6566), .S(n6375), .Z(n6192)
         );
  NAND2_X1 U7817 ( .A1(n6192), .A2(n6193), .ZN(n6381) );
  OAI211_X1 U7818 ( .C1(n6193), .C2(n6192), .A(n9728), .B(n6381), .ZN(n6194)
         );
  OAI211_X1 U7819 ( .C1(n9731), .C2(n6382), .A(n6195), .B(n6194), .ZN(P2_U3253) );
  INV_X1 U7820 ( .A(n6259), .ZN(n6196) );
  NOR2_X1 U7821 ( .A1(n6196), .A2(n6257), .ZN(n6199) );
  NAND2_X1 U7822 ( .A1(n6198), .A2(n6197), .ZN(n6258) );
  XOR2_X1 U7823 ( .A(n6199), .B(n6258), .Z(n6204) );
  AOI22_X1 U7824 ( .A1(n9073), .A2(n9115), .B1(n9092), .B2(n9117), .ZN(n6203)
         );
  INV_X1 U7825 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6200) );
  NOR2_X1 U7826 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6200), .ZN(n9606) );
  INV_X1 U7827 ( .A(n6526), .ZN(n6467) );
  NOR2_X1 U7828 ( .A1(n9102), .A2(n6467), .ZN(n6201) );
  AOI211_X1 U7829 ( .C1(n6464), .C2(n9099), .A(n9606), .B(n6201), .ZN(n6202)
         );
  OAI211_X1 U7830 ( .C1(n6204), .C2(n9086), .A(n6203), .B(n6202), .ZN(P1_U3228) );
  NAND2_X1 U7831 ( .A1(n6206), .A2(n6369), .ZN(n6208) );
  INV_X1 U7832 ( .A(n9739), .ZN(n6209) );
  INV_X1 U7833 ( .A(n8305), .ZN(n6211) );
  AND2_X1 U7834 ( .A1(n8315), .A2(n8313), .ZN(n8251) );
  NOR2_X1 U7835 ( .A1(n8251), .A2(n6389), .ZN(n6210) );
  AOI211_X1 U7836 ( .C1(n6211), .C2(n8313), .A(n8857), .B(n6210), .ZN(n6214)
         );
  OR2_X1 U7837 ( .A1(n6771), .A2(n8859), .ZN(n6213) );
  OR2_X1 U7838 ( .A1(n5082), .A2(n8861), .ZN(n6212) );
  NAND2_X1 U7839 ( .A1(n6213), .A2(n6212), .ZN(n6253) );
  NOR2_X1 U7840 ( .A1(n6214), .A2(n6253), .ZN(n9768) );
  MUX2_X1 U7841 ( .A(n6215), .B(n9768), .S(n8826), .Z(n6222) );
  OR2_X1 U7842 ( .A1(n6216), .A2(n9744), .ZN(n6537) );
  AND2_X1 U7843 ( .A1(n7660), .A2(n6537), .ZN(n9749) );
  XNOR2_X1 U7844 ( .A(n8251), .B(n6217), .ZN(n9770) );
  OR2_X1 U7845 ( .A1(n6218), .A2(n7547), .ZN(n8831) );
  NAND3_X1 U7846 ( .A1(n6450), .A2(n9786), .A3(n6219), .ZN(n9767) );
  OAI22_X1 U7847 ( .A1(n8831), .A2(n9767), .B1(n6256), .B2(n9742), .ZN(n6220)
         );
  AOI21_X1 U7848 ( .B1(n8823), .B2(n9770), .A(n6220), .ZN(n6221) );
  OAI211_X1 U7849 ( .C1(n6205), .C2(n8869), .A(n6222), .B(n6221), .ZN(P2_U3295) );
  INV_X1 U7850 ( .A(n7593), .ZN(n6272) );
  OAI21_X1 U7851 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(P1_IR_REG_14__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7852 ( .A1(n6224), .A2(n6223), .ZN(n6246) );
  NAND2_X1 U7853 ( .A1(n6225), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6228) );
  INV_X1 U7854 ( .A(n6228), .ZN(n6226) );
  NAND2_X1 U7855 ( .A1(n6226), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7856 ( .A1(n6228), .A2(n6227), .ZN(n6484) );
  AOI22_X1 U7857 ( .A1(n9172), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9488), .ZN(n6230) );
  OAI21_X1 U7858 ( .B1(n6272), .B2(n9493), .A(n6230), .ZN(P1_U3336) );
  INV_X1 U7859 ( .A(n6231), .ZN(n6236) );
  NAND2_X1 U7860 ( .A1(n6232), .A2(n9178), .ZN(n6273) );
  AOI21_X1 U7861 ( .B1(n7354), .B2(n6273), .A(n6233), .ZN(n6235) );
  OAI22_X1 U7862 ( .A1(n9365), .A2(n4681), .B1(n7841), .B2(n6276), .ZN(n6234)
         );
  NOR3_X1 U7863 ( .A1(n6236), .A2(n6235), .A3(n6234), .ZN(n6244) );
  AND2_X1 U7864 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  INV_X2 U7865 ( .A(n9367), .ZN(n9319) );
  NOR2_X2 U7866 ( .A1(n6241), .A2(n9178), .ZN(n9370) );
  AOI22_X1 U7867 ( .A1(n6242), .A2(n9370), .B1(n9319), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6243) );
  OAI21_X1 U7868 ( .B1(n6244), .B2(n9319), .A(n6243), .ZN(P1_U3290) );
  INV_X1 U7869 ( .A(n8681), .ZN(n8676) );
  INV_X1 U7870 ( .A(n7455), .ZN(n6247) );
  OAI222_X1 U7871 ( .A1(P2_U3152), .A2(n8676), .B1(n8233), .B2(n6247), .C1(
        n9884), .C2(n8979), .ZN(P2_U3342) );
  XNOR2_X1 U7872 ( .A(n6246), .B(n6245), .ZN(n9158) );
  INV_X1 U7873 ( .A(n9158), .ZN(n9148) );
  OAI222_X1 U7874 ( .A1(n9495), .A2(n6248), .B1(P1_U3084), .B2(n9148), .C1(
        n6247), .C2(n9493), .ZN(P1_U3337) );
  NAND2_X1 U7875 ( .A1(n8620), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6249) );
  OAI21_X1 U7876 ( .B1(n8746), .B2(n8620), .A(n6249), .ZN(P2_U3581) );
  INV_X1 U7877 ( .A(n8606), .ZN(n8554) );
  NOR2_X1 U7878 ( .A1(n8554), .A2(P2_U3152), .ZN(n7678) );
  INV_X1 U7879 ( .A(n6888), .ZN(n8580) );
  INV_X1 U7880 ( .A(n8587), .ZN(n8604) );
  OAI21_X1 U7881 ( .B1(n6251), .B2(n6250), .A(n7672), .ZN(n6252) );
  AOI22_X1 U7882 ( .A1(n8580), .A2(n6253), .B1(n8604), .B2(n6252), .ZN(n6255)
         );
  OAI211_X1 U7883 ( .C1(n7678), .C2(n6256), .A(n6255), .B(n6254), .ZN(P2_U3224) );
  OR2_X1 U7884 ( .A1(n6258), .A2(n6257), .ZN(n6260) );
  NAND2_X1 U7885 ( .A1(n6260), .A2(n6259), .ZN(n6265) );
  INV_X1 U7886 ( .A(n6261), .ZN(n6262) );
  XNOR2_X1 U7887 ( .A(n6263), .B(n6262), .ZN(n6264) );
  XNOR2_X1 U7888 ( .A(n6265), .B(n6264), .ZN(n6270) );
  AOI22_X1 U7889 ( .A1(n9073), .A2(n9114), .B1(n9092), .B2(n9116), .ZN(n6269)
         );
  INV_X1 U7890 ( .A(n6488), .ZN(n9703) );
  NOR2_X1 U7891 ( .A1(n9102), .A2(n9703), .ZN(n6266) );
  AOI211_X1 U7892 ( .C1(n6424), .C2(n9099), .A(n6267), .B(n6266), .ZN(n6268)
         );
  OAI211_X1 U7893 ( .C1(n6270), .C2(n9086), .A(n6269), .B(n6268), .ZN(P1_U3225) );
  INV_X1 U7894 ( .A(n8697), .ZN(n8689) );
  OAI222_X1 U7895 ( .A1(P2_U3152), .A2(n8689), .B1(n8233), .B2(n6272), .C1(
        n6271), .C2(n8979), .ZN(P2_U3341) );
  MUX2_X1 U7896 ( .A(n6274), .B(P1_REG2_REG_2__SCAN_IN), .S(n9356), .Z(n6275)
         );
  INV_X1 U7897 ( .A(n6275), .ZN(n6282) );
  INV_X1 U7898 ( .A(n6276), .ZN(n6277) );
  INV_X1 U7899 ( .A(n4307), .ZN(n7839) );
  INV_X1 U7900 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6278) );
  OAI22_X1 U7901 ( .A1(n9364), .A2(n7839), .B1(n6278), .B2(n9365), .ZN(n6279)
         );
  AOI21_X1 U7902 ( .B1(n9322), .B2(n6280), .A(n6279), .ZN(n6281) );
  OAI211_X1 U7903 ( .C1(n6283), .C2(n7363), .A(n6282), .B(n6281), .ZN(P1_U3289) );
  OAI21_X1 U7904 ( .B1(n9322), .B2(n9183), .A(n7684), .ZN(n6285) );
  INV_X2 U7905 ( .A(n9365), .ZN(n9343) );
  AOI22_X1 U7906 ( .A1(n9356), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9343), .ZN(n6284) );
  OAI211_X1 U7907 ( .C1(n9356), .C2(n6286), .A(n6285), .B(n6284), .ZN(P1_U3291) );
  OR2_X1 U7908 ( .A1(n6287), .A2(n6067), .ZN(n6290) );
  OR2_X1 U7909 ( .A1(n6120), .A2(n6288), .ZN(n6289) );
  OAI211_X1 U7910 ( .C1(n5944), .C2(n6346), .A(n6290), .B(n6289), .ZN(n6697)
         );
  NAND2_X1 U7911 ( .A1(n9113), .A2(n8508), .ZN(n6295) );
  NAND2_X1 U7912 ( .A1(n6697), .A2(n5930), .ZN(n6294) );
  NAND2_X1 U7913 ( .A1(n6295), .A2(n6294), .ZN(n6296) );
  XNOR2_X1 U7914 ( .A(n6296), .B(n8482), .ZN(n6302) );
  INV_X1 U7915 ( .A(n6302), .ZN(n6300) );
  NAND2_X1 U7916 ( .A1(n9002), .A2(n9113), .ZN(n6298) );
  NAND2_X1 U7917 ( .A1(n6697), .A2(n8508), .ZN(n6297) );
  AND2_X1 U7918 ( .A1(n6298), .A2(n6297), .ZN(n6301) );
  INV_X1 U7919 ( .A(n6301), .ZN(n6299) );
  NAND2_X1 U7920 ( .A1(n6300), .A2(n6299), .ZN(n6650) );
  NAND2_X1 U7921 ( .A1(n6302), .A2(n6301), .ZN(n6648) );
  NAND2_X1 U7922 ( .A1(n6650), .A2(n6648), .ZN(n6303) );
  XNOR2_X1 U7923 ( .A(n6649), .B(n6303), .ZN(n6304) );
  NAND2_X1 U7924 ( .A1(n6304), .A2(n9088), .ZN(n6316) );
  NAND2_X1 U7925 ( .A1(n7244), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7926 ( .A1(n7869), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7927 ( .A1(n6306), .A2(n6305), .ZN(n6307) );
  AND2_X1 U7928 ( .A1(n6662), .A2(n6307), .ZN(n6690) );
  NAND2_X1 U7929 ( .A1(n7346), .A2(n6690), .ZN(n6309) );
  NAND2_X1 U7930 ( .A1(n7822), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6308) );
  NAND4_X1 U7931 ( .A1(n6311), .A2(n6310), .A3(n6309), .A4(n6308), .ZN(n9112)
         );
  INV_X1 U7932 ( .A(n9114), .ZN(n6606) );
  INV_X1 U7933 ( .A(n6696), .ZN(n6312) );
  OAI22_X1 U7934 ( .A1(n9051), .A2(n6606), .B1(n9050), .B2(n6312), .ZN(n6313)
         );
  AOI211_X1 U7935 ( .C1(n9073), .C2(n9112), .A(n6314), .B(n6313), .ZN(n6315)
         );
  OAI211_X1 U7936 ( .C1(n6677), .C2(n9102), .A(n6316), .B(n6315), .ZN(P1_U3211) );
  INV_X1 U7937 ( .A(n7242), .ZN(n6320) );
  NAND2_X1 U7938 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6322) );
  INV_X1 U7939 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8986) );
  INV_X1 U7940 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9033) );
  INV_X1 U7941 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9094) );
  INV_X1 U7942 ( .A(n7887), .ZN(n6327) );
  AND2_X1 U7943 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6326) );
  NAND2_X1 U7944 ( .A1(n6327), .A2(n6326), .ZN(n7889) );
  INV_X1 U7945 ( .A(n7889), .ZN(n8132) );
  NAND2_X1 U7946 ( .A1(n7822), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U7947 ( .A1(n4305), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U7948 ( .A1(n7244), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6328) );
  NAND3_X1 U7949 ( .A1(n6330), .A2(n6329), .A3(n6328), .ZN(n6331) );
  AOI21_X1 U7950 ( .B1(n8132), .B2(n7346), .A(n6331), .ZN(n9197) );
  NAND2_X1 U7951 ( .A1(n9119), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6332) );
  OAI21_X1 U7952 ( .B1(n9197), .B2(n9119), .A(n6332), .ZN(P1_U3584) );
  INV_X1 U7953 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9560) );
  AOI22_X1 U7954 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9646), .B1(n6333), .B2(
        n9560), .ZN(n9649) );
  NOR2_X1 U7955 ( .A1(n9125), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6334) );
  AOI21_X1 U7956 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9125), .A(n6334), .ZN(
        n9128) );
  INV_X1 U7957 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6335) );
  MUX2_X1 U7958 ( .A(n6335), .B(P1_REG1_REG_8__SCAN_IN), .S(n9628), .Z(n9617)
         );
  NAND2_X1 U7959 ( .A1(n6346), .A2(n6336), .ZN(n6338) );
  NAND2_X1 U7960 ( .A1(n6338), .A2(n6337), .ZN(n9616) );
  NOR2_X1 U7961 ( .A1(n9617), .A2(n9616), .ZN(n9615) );
  AOI21_X1 U7962 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9628), .A(n9615), .ZN(
        n9634) );
  NOR2_X1 U7963 ( .A1(n9642), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6339) );
  AOI21_X1 U7964 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9642), .A(n6339), .ZN(
        n9633) );
  NAND2_X1 U7965 ( .A1(n9634), .A2(n9633), .ZN(n9632) );
  OAI21_X1 U7966 ( .B1(n9642), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9632), .ZN(
        n9129) );
  NAND2_X1 U7967 ( .A1(n9128), .A2(n9129), .ZN(n9127) );
  OAI21_X1 U7968 ( .B1(n9125), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9127), .ZN(
        n9648) );
  NAND2_X1 U7969 ( .A1(n9649), .A2(n9648), .ZN(n9647) );
  OAI21_X1 U7970 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9646), .A(n9647), .ZN(
        n6342) );
  INV_X1 U7971 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6340) );
  MUX2_X1 U7972 ( .A(n6340), .B(P1_REG1_REG_12__SCAN_IN), .S(n6349), .Z(n6341)
         );
  NAND2_X1 U7973 ( .A1(n6341), .A2(n6342), .ZN(n6598) );
  OAI21_X1 U7974 ( .B1(n6342), .B2(n6341), .A(n6598), .ZN(n6355) );
  NAND2_X1 U7975 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7099) );
  NAND2_X1 U7976 ( .A1(n9685), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6343) );
  OAI211_X1 U7977 ( .C1(n9592), .C2(n6349), .A(n7099), .B(n6343), .ZN(n6354)
         );
  NOR2_X1 U7978 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n9646), .ZN(n6344) );
  AOI21_X1 U7979 ( .B1(n9646), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6344), .ZN(
        n9652) );
  NAND2_X1 U7980 ( .A1(n9642), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6347) );
  OAI21_X1 U7981 ( .B1(n9642), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6347), .ZN(
        n9639) );
  NOR2_X1 U7982 ( .A1(n9640), .A2(n9639), .ZN(n9638) );
  AOI21_X1 U7983 ( .B1(n9642), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9638), .ZN(
        n9123) );
  NAND2_X1 U7984 ( .A1(n9125), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6348) );
  OAI21_X1 U7985 ( .B1(n9125), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6348), .ZN(
        n9122) );
  NOR2_X1 U7986 ( .A1(n9123), .A2(n9122), .ZN(n9121) );
  NAND2_X1 U7987 ( .A1(n9652), .A2(n9651), .ZN(n9650) );
  OAI21_X1 U7988 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9646), .A(n9650), .ZN(
        n6352) );
  NAND2_X1 U7989 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7024), .ZN(n6350) );
  OAI21_X1 U7990 ( .B1(n7024), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6350), .ZN(
        n6351) );
  AOI211_X1 U7991 ( .C1(n6352), .C2(n6351), .A(n6592), .B(n9637), .ZN(n6353)
         );
  AOI211_X1 U7992 ( .C1(n9686), .C2(n6355), .A(n6354), .B(n6353), .ZN(n6356)
         );
  INV_X1 U7993 ( .A(n6356), .ZN(P1_U3253) );
  INV_X1 U7994 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6368) );
  INV_X1 U7995 ( .A(n8256), .ZN(n6358) );
  XNOR2_X1 U7996 ( .A(n6357), .B(n6358), .ZN(n9748) );
  NAND2_X1 U7997 ( .A1(n6359), .A2(n8219), .ZN(n6360) );
  NAND2_X1 U7998 ( .A1(n6360), .A2(n9786), .ZN(n6361) );
  NOR2_X1 U7999 ( .A1(n6403), .A2(n6361), .ZN(n9745) );
  XNOR2_X1 U8000 ( .A(n8256), .B(n6362), .ZN(n6363) );
  NAND2_X1 U8001 ( .A1(n6363), .A2(n8817), .ZN(n6365) );
  INV_X1 U8002 ( .A(n8861), .ZN(n7567) );
  AOI22_X1 U8003 ( .A1(n8636), .A2(n7567), .B1(n7566), .B2(n8638), .ZN(n6364)
         );
  NAND2_X1 U8004 ( .A1(n6365), .A2(n6364), .ZN(n9738) );
  AOI211_X1 U8005 ( .C1(n9772), .C2(n8219), .A(n9745), .B(n9738), .ZN(n6366)
         );
  OAI21_X1 U8006 ( .B1(n9790), .B2(n9748), .A(n6366), .ZN(n6371) );
  NAND2_X1 U8007 ( .A1(n6371), .A2(n9817), .ZN(n6367) );
  OAI21_X1 U8008 ( .B1(n9817), .B2(n6368), .A(n6367), .ZN(P2_U3466) );
  INV_X1 U8009 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8010 ( .A1(n6371), .A2(n9830), .ZN(n6372) );
  OAI21_X1 U8011 ( .B1(n9830), .B2(n6373), .A(n6372), .ZN(P2_U3525) );
  NAND2_X1 U8012 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6797) );
  INV_X1 U8013 ( .A(n6797), .ZN(n6380) );
  INV_X1 U8014 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6376) );
  MUX2_X1 U8015 ( .A(n6376), .B(P2_REG1_REG_9__SCAN_IN), .S(n6580), .Z(n6377)
         );
  AOI211_X1 U8016 ( .C1(n6378), .C2(n6377), .A(n6579), .B(n9732), .ZN(n6379)
         );
  AOI211_X1 U8017 ( .C1(n9729), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n6380), .B(
        n6379), .ZN(n6387) );
  OAI21_X1 U8018 ( .B1(n6382), .B2(n6566), .A(n6381), .ZN(n6385) );
  MUX2_X1 U8019 ( .A(n6831), .B(P2_REG2_REG_9__SCAN_IN), .S(n6580), .Z(n6383)
         );
  INV_X1 U8020 ( .A(n6383), .ZN(n6384) );
  NAND2_X1 U8021 ( .A1(n6384), .A2(n6385), .ZN(n6573) );
  OAI211_X1 U8022 ( .C1(n6385), .C2(n6384), .A(n9728), .B(n6573), .ZN(n6386)
         );
  OAI211_X1 U8023 ( .C1(n9731), .C2(n6388), .A(n6387), .B(n6386), .ZN(P2_U3254) );
  INV_X1 U8024 ( .A(n6389), .ZN(n6390) );
  INV_X1 U8025 ( .A(n6771), .ZN(n8641) );
  AND2_X1 U8026 ( .A1(n8641), .A2(n6770), .ZN(n8302) );
  NOR2_X1 U8027 ( .A1(n6390), .A2(n8302), .ZN(n8252) );
  INV_X1 U8028 ( .A(n8252), .ZN(n9764) );
  AOI22_X1 U8029 ( .A1(n9764), .A2(n8817), .B1(n7567), .B2(n6391), .ZN(n9766)
         );
  OAI22_X1 U8030 ( .A1(n9766), .A2(n9752), .B1(n6776), .B2(n9742), .ZN(n6392)
         );
  AOI21_X1 U8031 ( .B1(n9752), .B2(P2_REG2_REG_0__SCAN_IN), .A(n6392), .ZN(
        n6394) );
  OAI21_X1 U8032 ( .B1(n8864), .B2(n8828), .A(n9762), .ZN(n6393) );
  OAI211_X1 U8033 ( .C1(n8252), .C2(n8873), .A(n6394), .B(n6393), .ZN(P2_U3296) );
  NAND2_X1 U8034 ( .A1(n6396), .A2(n6395), .ZN(n6471) );
  INV_X1 U8035 ( .A(n6471), .ZN(n6398) );
  INV_X1 U8036 ( .A(n6396), .ZN(n6397) );
  AOI22_X1 U8037 ( .A1(n6398), .A2(n6470), .B1(n8258), .B2(n6397), .ZN(n9793)
         );
  OAI21_X1 U8038 ( .B1(n6400), .B2(n8258), .A(n6399), .ZN(n6401) );
  AOI222_X1 U8039 ( .A1(n8817), .A2(n6401), .B1(n8635), .B2(n7567), .C1(n8637), 
        .C2(n7566), .ZN(n9796) );
  MUX2_X1 U8040 ( .A(n6402), .B(n9796), .S(n8826), .Z(n6407) );
  NOR2_X1 U8041 ( .A1(n6403), .A2(n9794), .ZN(n6404) );
  OR2_X1 U8042 ( .A1(n6476), .A2(n6404), .ZN(n9795) );
  OAI22_X1 U8043 ( .A1(n9795), .A2(n8736), .B1(n6627), .B2(n9742), .ZN(n6405)
         );
  AOI21_X1 U8044 ( .B1(n8828), .B2(n6630), .A(n6405), .ZN(n6406) );
  OAI211_X1 U8045 ( .C1(n9793), .C2(n8873), .A(n6407), .B(n6406), .ZN(P2_U3290) );
  INV_X1 U8046 ( .A(n9118), .ZN(n6414) );
  NAND2_X1 U8047 ( .A1(n6414), .A2(n4307), .ZN(n6409) );
  NAND2_X1 U8048 ( .A1(n6456), .A2(n6169), .ZN(n6417) );
  INV_X1 U8049 ( .A(n6417), .ZN(n8065) );
  NAND2_X1 U8050 ( .A1(n6467), .A2(n9116), .ZN(n7917) );
  AND2_X1 U8051 ( .A1(n7917), .A2(n6457), .ZN(n8063) );
  INV_X1 U8052 ( .A(n9116), .ZN(n6419) );
  NAND2_X1 U8053 ( .A1(n6419), .A2(n6526), .ZN(n7914) );
  INV_X1 U8054 ( .A(n7914), .ZN(n6410) );
  INV_X1 U8055 ( .A(n9115), .ZN(n6455) );
  NAND2_X1 U8056 ( .A1(n6455), .A2(n6488), .ZN(n7918) );
  NAND2_X1 U8057 ( .A1(n9703), .A2(n9115), .ZN(n7920) );
  INV_X1 U8058 ( .A(n6607), .ZN(n8031) );
  XNOR2_X1 U8059 ( .A(n6493), .B(n8031), .ZN(n6411) );
  NAND2_X1 U8060 ( .A1(n6411), .A2(n9355), .ZN(n6413) );
  AOI22_X1 U8061 ( .A1(n9380), .A2(n9116), .B1(n9372), .B2(n9114), .ZN(n6412)
         );
  NAND2_X1 U8062 ( .A1(n6413), .A2(n6412), .ZN(n9705) );
  INV_X1 U8063 ( .A(n9705), .ZN(n6429) );
  NAND2_X1 U8064 ( .A1(n6414), .A2(n7839), .ZN(n6415) );
  NAND2_X1 U8065 ( .A1(n6416), .A2(n6415), .ZN(n6430) );
  NAND2_X1 U8066 ( .A1(n6430), .A2(n8028), .ZN(n6431) );
  NAND2_X1 U8067 ( .A1(n6456), .A2(n9695), .ZN(n6418) );
  NAND2_X1 U8068 ( .A1(n6431), .A2(n6418), .ZN(n6454) );
  NAND2_X1 U8069 ( .A1(n7914), .A2(n7917), .ZN(n8029) );
  NAND2_X1 U8070 ( .A1(n6454), .A2(n8029), .ZN(n6453) );
  NAND2_X1 U8071 ( .A1(n6419), .A2(n6467), .ZN(n6420) );
  NAND2_X1 U8072 ( .A1(n6453), .A2(n6420), .ZN(n6609) );
  INV_X1 U8073 ( .A(n6490), .ZN(n6421) );
  AOI21_X1 U8074 ( .B1(n6607), .B2(n6609), .A(n6421), .ZN(n9707) );
  INV_X1 U8075 ( .A(n9383), .ZN(n6704) );
  NAND2_X1 U8076 ( .A1(n6432), .A2(n9695), .ZN(n6463) );
  OR2_X1 U8077 ( .A1(n6463), .A2(n6526), .ZN(n6423) );
  INV_X1 U8078 ( .A(n6423), .ZN(n6462) );
  INV_X1 U8079 ( .A(n6499), .ZN(n6500) );
  OAI211_X1 U8080 ( .C1(n9703), .C2(n6462), .A(n6500), .B(n9437), .ZN(n9702)
         );
  INV_X1 U8081 ( .A(n9370), .ZN(n7256) );
  AOI22_X1 U8082 ( .A1(n9356), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6424), .B2(
        n9343), .ZN(n6426) );
  NAND2_X1 U8083 ( .A1(n9183), .A2(n6488), .ZN(n6425) );
  OAI211_X1 U8084 ( .C1(n9702), .C2(n7256), .A(n6426), .B(n6425), .ZN(n6427)
         );
  AOI21_X1 U8085 ( .B1(n9707), .B2(n6704), .A(n6427), .ZN(n6428) );
  OAI21_X1 U8086 ( .B1(n9319), .B2(n6429), .A(n6428), .ZN(P1_U3286) );
  OAI21_X1 U8087 ( .B1(n6430), .B2(n8028), .A(n6431), .ZN(n9700) );
  INV_X1 U8088 ( .A(n9322), .ZN(n9186) );
  OR2_X1 U8089 ( .A1(n6432), .A2(n9695), .ZN(n6433) );
  NAND2_X1 U8090 ( .A1(n6463), .A2(n6433), .ZN(n9697) );
  AOI22_X1 U8091 ( .A1(n9183), .A2(n6169), .B1(n9343), .B2(n9972), .ZN(n6434)
         );
  OAI21_X1 U8092 ( .B1(n9186), .B2(n9697), .A(n6434), .ZN(n6439) );
  XNOR2_X1 U8093 ( .A(n8064), .B(n8028), .ZN(n6437) );
  NAND2_X1 U8094 ( .A1(n9700), .A2(n7158), .ZN(n6436) );
  AOI22_X1 U8095 ( .A1(n9380), .A2(n9118), .B1(n9372), .B2(n9116), .ZN(n6435)
         );
  OAI211_X1 U8096 ( .C1(n9374), .C2(n6437), .A(n6436), .B(n6435), .ZN(n9698)
         );
  MUX2_X1 U8097 ( .A(n9698), .B(P1_REG2_REG_3__SCAN_IN), .S(n9319), .Z(n6438)
         );
  AOI211_X1 U8098 ( .C1(n7165), .C2(n9700), .A(n6439), .B(n6438), .ZN(n6440)
         );
  INV_X1 U8099 ( .A(n6440), .ZN(P1_U3288) );
  XNOR2_X1 U8100 ( .A(n6441), .B(n6443), .ZN(n9777) );
  NOR2_X1 U8101 ( .A1(n8826), .A2(n5763), .ZN(n6449) );
  NAND2_X1 U8102 ( .A1(n6444), .A2(n6443), .ZN(n6445) );
  NAND2_X1 U8103 ( .A1(n6442), .A2(n6445), .ZN(n6447) );
  OAI22_X1 U8104 ( .A1(n7676), .A2(n8859), .B1(n5100), .B2(n8861), .ZN(n6446)
         );
  AOI21_X1 U8105 ( .B1(n6447), .B2(n8817), .A(n6446), .ZN(n9775) );
  OAI22_X1 U8106 ( .A1(n9775), .A2(n9752), .B1(n7677), .B2(n9742), .ZN(n6448)
         );
  AOI211_X1 U8107 ( .C1(n8823), .C2(n9777), .A(n6449), .B(n6448), .ZN(n6452)
         );
  AOI21_X1 U8108 ( .B1(n9771), .B2(n6450), .A(n6539), .ZN(n9773) );
  AOI22_X1 U8109 ( .A1(n9773), .A2(n8864), .B1(n8828), .B2(n9771), .ZN(n6451)
         );
  NAND2_X1 U8110 ( .A1(n6452), .A2(n6451), .ZN(P2_U3294) );
  OAI21_X1 U8111 ( .B1(n6454), .B2(n8029), .A(n6453), .ZN(n6525) );
  OAI22_X1 U8112 ( .A1(n6456), .A2(n9331), .B1(n6455), .B2(n9329), .ZN(n6461)
         );
  NAND2_X1 U8113 ( .A1(n6458), .A2(n6457), .ZN(n7916) );
  XOR2_X1 U8114 ( .A(n8029), .B(n7916), .Z(n6459) );
  NOR2_X1 U8115 ( .A1(n6459), .A2(n9374), .ZN(n6460) );
  AOI211_X1 U8116 ( .C1(n7158), .C2(n6525), .A(n6461), .B(n6460), .ZN(n6529)
         );
  AOI21_X1 U8117 ( .B1(n6526), .B2(n6463), .A(n6462), .ZN(n6527) );
  NAND2_X1 U8118 ( .A1(n6527), .A2(n9322), .ZN(n6466) );
  AOI22_X1 U8119 ( .A1(n9356), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6464), .B2(
        n9343), .ZN(n6465) );
  OAI211_X1 U8120 ( .C1(n6467), .C2(n9364), .A(n6466), .B(n6465), .ZN(n6468)
         );
  AOI21_X1 U8121 ( .B1(n6525), .B2(n7165), .A(n6468), .ZN(n6469) );
  OAI21_X1 U8122 ( .B1(n6529), .B2(n9319), .A(n6469), .ZN(P1_U3287) );
  NAND3_X1 U8123 ( .A1(n6471), .A2(n8259), .A3(n6470), .ZN(n6472) );
  AND2_X1 U8124 ( .A1(n6473), .A2(n6472), .ZN(n6514) );
  XNOR2_X1 U8125 ( .A(n6474), .B(n8259), .ZN(n6475) );
  AOI222_X1 U8126 ( .A1(n8817), .A2(n6475), .B1(n8636), .B2(n7566), .C1(n8634), 
        .C2(n7567), .ZN(n6506) );
  INV_X1 U8127 ( .A(n6476), .ZN(n6478) );
  INV_X1 U8128 ( .A(n6567), .ZN(n6477) );
  AOI21_X1 U8129 ( .B1(n6479), .B2(n6478), .A(n6477), .ZN(n6511) );
  AOI22_X1 U8130 ( .A1(n6511), .A2(n9786), .B1(n9772), .B2(n6479), .ZN(n6480)
         );
  OAI211_X1 U8131 ( .C1(n9790), .C2(n6514), .A(n6506), .B(n6480), .ZN(n6482)
         );
  NAND2_X1 U8132 ( .A1(n6482), .A2(n9830), .ZN(n6481) );
  OAI21_X1 U8133 ( .B1(n9830), .B2(n5825), .A(n6481), .ZN(P2_U3527) );
  NAND2_X1 U8134 ( .A1(n6482), .A2(n9817), .ZN(n6483) );
  OAI21_X1 U8135 ( .B1(n9817), .B2(n5152), .A(n6483), .ZN(P2_U3472) );
  INV_X1 U8136 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6486) );
  INV_X1 U8137 ( .A(n7799), .ZN(n6487) );
  NAND2_X1 U8138 ( .A1(n6484), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6485) );
  XNOR2_X1 U8139 ( .A(n6485), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9677) );
  INV_X1 U8140 ( .A(n9677), .ZN(n9170) );
  OAI222_X1 U8141 ( .A1(n9495), .A2(n6486), .B1(n9493), .B2(n6487), .C1(
        P1_U3084), .C2(n9170), .ZN(P1_U3335) );
  INV_X1 U8142 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10031) );
  INV_X1 U8143 ( .A(n8707), .ZN(n8710) );
  OAI222_X1 U8144 ( .A1(n8979), .A2(n10031), .B1(n8233), .B2(n6487), .C1(
        P2_U3152), .C2(n8710), .ZN(P2_U3340) );
  NAND2_X1 U8145 ( .A1(n9115), .A2(n6488), .ZN(n6489) );
  AND2_X1 U8146 ( .A1(n6490), .A2(n6489), .ZN(n6492) );
  NAND2_X1 U8147 ( .A1(n6606), .A2(n6515), .ZN(n8067) );
  NAND2_X1 U8148 ( .A1(n6605), .A2(n9114), .ZN(n8070) );
  NAND2_X1 U8149 ( .A1(n8067), .A2(n8070), .ZN(n6494) );
  AND2_X1 U8150 ( .A1(n6494), .A2(n6489), .ZN(n6610) );
  NAND2_X1 U8151 ( .A1(n6490), .A2(n6610), .ZN(n6491) );
  OAI21_X1 U8152 ( .B1(n6492), .B2(n6494), .A(n6491), .ZN(n6498) );
  INV_X1 U8153 ( .A(n6498), .ZN(n6519) );
  NAND2_X1 U8154 ( .A1(n6493), .A2(n7918), .ZN(n6615) );
  NAND2_X1 U8155 ( .A1(n6615), .A2(n7920), .ZN(n7928) );
  INV_X1 U8156 ( .A(n6494), .ZN(n8034) );
  XNOR2_X1 U8157 ( .A(n7928), .B(n8034), .ZN(n6496) );
  AOI22_X1 U8158 ( .A1(n9380), .A2(n9115), .B1(n9372), .B2(n9113), .ZN(n6495)
         );
  OAI21_X1 U8159 ( .B1(n6496), .B2(n9374), .A(n6495), .ZN(n6497) );
  AOI21_X1 U8160 ( .B1(n6498), .B2(n7158), .A(n6497), .ZN(n6518) );
  MUX2_X1 U8161 ( .A(n6518), .B(n5868), .S(n9319), .Z(n6505) );
  AOI21_X1 U8162 ( .B1(n6515), .B2(n6500), .A(n6620), .ZN(n6516) );
  INV_X1 U8163 ( .A(n6501), .ZN(n6502) );
  OAI22_X1 U8164 ( .A1(n9364), .A2(n6605), .B1(n6502), .B2(n9365), .ZN(n6503)
         );
  AOI21_X1 U8165 ( .B1(n6516), .B2(n9322), .A(n6503), .ZN(n6504) );
  OAI211_X1 U8166 ( .C1(n6519), .C2(n7363), .A(n6505), .B(n6504), .ZN(P1_U3285) );
  INV_X2 U8167 ( .A(n9752), .ZN(n8826) );
  MUX2_X1 U8168 ( .A(n6507), .B(n6506), .S(n8826), .Z(n6513) );
  OAI22_X1 U8169 ( .A1(n8869), .A2(n6509), .B1(n9742), .B2(n6508), .ZN(n6510)
         );
  AOI21_X1 U8170 ( .B1(n6511), .B2(n8864), .A(n6510), .ZN(n6512) );
  OAI211_X1 U8171 ( .C1(n6514), .C2(n8873), .A(n6513), .B(n6512), .ZN(P2_U3289) );
  INV_X1 U8172 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6521) );
  AOI22_X1 U8173 ( .A1(n6516), .A2(n9437), .B1(n9465), .B2(n6515), .ZN(n6517)
         );
  OAI211_X1 U8174 ( .C1(n6519), .C2(n9535), .A(n6518), .B(n6517), .ZN(n6522)
         );
  NAND2_X1 U8175 ( .A1(n6522), .A2(n9561), .ZN(n6520) );
  OAI21_X1 U8176 ( .B1(n9561), .B2(n6521), .A(n6520), .ZN(P1_U3529) );
  INV_X1 U8177 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U8178 ( .A1(n6522), .A2(n9719), .ZN(n6523) );
  OAI21_X1 U8179 ( .B1(n9719), .B2(n6524), .A(n6523), .ZN(P1_U3472) );
  INV_X1 U8180 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6532) );
  INV_X1 U8181 ( .A(n6525), .ZN(n6530) );
  AOI22_X1 U8182 ( .A1(n6527), .A2(n9437), .B1(n9465), .B2(n6526), .ZN(n6528)
         );
  OAI211_X1 U8183 ( .C1(n6530), .C2(n9535), .A(n6529), .B(n6528), .ZN(n6533)
         );
  NAND2_X1 U8184 ( .A1(n6533), .A2(n9719), .ZN(n6531) );
  OAI21_X1 U8185 ( .B1(n9719), .B2(n6532), .A(n6531), .ZN(P1_U3466) );
  NAND2_X1 U8186 ( .A1(n6533), .A2(n9561), .ZN(n6534) );
  OAI21_X1 U8187 ( .B1(n9561), .B2(n6535), .A(n6534), .ZN(P1_U3527) );
  XNOR2_X1 U8188 ( .A(n8307), .B(n6536), .ZN(n9779) );
  INV_X1 U8189 ( .A(n6537), .ZN(n6538) );
  AND2_X1 U8190 ( .A1(n8826), .A2(n6538), .ZN(n7333) );
  INV_X1 U8191 ( .A(n7333), .ZN(n7670) );
  OAI22_X1 U8192 ( .A1(n8826), .A2(n5762), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9742), .ZN(n6541) );
  OAI21_X1 U8193 ( .B1(n6539), .B2(n9780), .A(n6554), .ZN(n9781) );
  NOR2_X1 U8194 ( .A1(n8736), .A2(n9781), .ZN(n6540) );
  AOI211_X1 U8195 ( .C1(n8828), .C2(n6542), .A(n6541), .B(n6540), .ZN(n6549)
         );
  AOI22_X1 U8196 ( .A1(n8640), .A2(n7566), .B1(n7567), .B2(n8638), .ZN(n6547)
         );
  INV_X1 U8197 ( .A(n6543), .ZN(n6545) );
  AND3_X1 U8198 ( .A1(n8254), .A2(n6442), .A3(n8316), .ZN(n6544) );
  OAI21_X1 U8199 ( .B1(n6545), .B2(n6544), .A(n8817), .ZN(n6546) );
  OAI211_X1 U8200 ( .C1(n9779), .C2(n7660), .A(n6547), .B(n6546), .ZN(n9782)
         );
  NAND2_X1 U8201 ( .A1(n9782), .A2(n8826), .ZN(n6548) );
  OAI211_X1 U8202 ( .C1(n9779), .C2(n7670), .A(n6549), .B(n6548), .ZN(P2_U3293) );
  XNOR2_X1 U8203 ( .A(n6550), .B(n4451), .ZN(n6552) );
  OAI22_X1 U8204 ( .A1(n6632), .A2(n8861), .B1(n5100), .B2(n8859), .ZN(n6551)
         );
  AOI21_X1 U8205 ( .B1(n6552), .B2(n8817), .A(n6551), .ZN(n9789) );
  XOR2_X1 U8206 ( .A(n8255), .B(n6553), .Z(n9791) );
  OR2_X1 U8207 ( .A1(n9791), .A2(n8873), .ZN(n6559) );
  XNOR2_X1 U8208 ( .A(n6554), .B(n6555), .ZN(n9787) );
  OAI22_X1 U8209 ( .A1(n8826), .A2(n5767), .B1(n6812), .B2(n9742), .ZN(n6557)
         );
  NOR2_X1 U8210 ( .A1(n8869), .A2(n6555), .ZN(n6556) );
  AOI211_X1 U8211 ( .C1(n8864), .C2(n9787), .A(n6557), .B(n6556), .ZN(n6558)
         );
  OAI211_X1 U8212 ( .C1(n9752), .C2(n9789), .A(n6559), .B(n6558), .ZN(P2_U3292) );
  NAND2_X1 U8213 ( .A1(n6561), .A2(n8332), .ZN(n6562) );
  NAND2_X1 U8214 ( .A1(n6560), .A2(n6562), .ZN(n9801) );
  AOI22_X1 U8215 ( .A1(n7566), .A2(n8635), .B1(n8633), .B2(n7567), .ZN(n6565)
         );
  XNOR2_X1 U8216 ( .A(n6821), .B(n8346), .ZN(n6563) );
  NAND2_X1 U8217 ( .A1(n6563), .A2(n8817), .ZN(n6564) );
  OAI211_X1 U8218 ( .C1(n9801), .C2(n7660), .A(n6565), .B(n6564), .ZN(n9804)
         );
  NAND2_X1 U8219 ( .A1(n9804), .A2(n8826), .ZN(n6572) );
  OAI22_X1 U8220 ( .A1(n8826), .A2(n6566), .B1(n6740), .B2(n9742), .ZN(n6570)
         );
  NAND2_X1 U8221 ( .A1(n6567), .A2(n9802), .ZN(n6568) );
  NAND2_X1 U8222 ( .A1(n6828), .A2(n6568), .ZN(n9803) );
  NOR2_X1 U8223 ( .A1(n9803), .A2(n8736), .ZN(n6569) );
  AOI211_X1 U8224 ( .C1(n8828), .C2(n9802), .A(n6570), .B(n6569), .ZN(n6571)
         );
  OAI211_X1 U8225 ( .C1(n9801), .C2(n7670), .A(n6572), .B(n6571), .ZN(P2_U3288) );
  NAND2_X1 U8226 ( .A1(n6580), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U8227 ( .A1(n6574), .A2(n6573), .ZN(n6577) );
  MUX2_X1 U8228 ( .A(n7662), .B(P2_REG2_REG_10__SCAN_IN), .S(n6963), .Z(n6575)
         );
  INV_X1 U8229 ( .A(n6575), .ZN(n6576) );
  NAND2_X1 U8230 ( .A1(n6576), .A2(n6577), .ZN(n6956) );
  OAI211_X1 U8231 ( .C1(n6577), .C2(n6576), .A(n9728), .B(n6956), .ZN(n6587)
         );
  INV_X1 U8232 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6578) );
  MUX2_X1 U8233 ( .A(n6578), .B(P2_REG1_REG_10__SCAN_IN), .S(n6963), .Z(n6582)
         );
  NOR2_X1 U8234 ( .A1(n6581), .A2(n6582), .ZN(n6962) );
  AOI21_X1 U8235 ( .B1(n6582), .B2(n6581), .A(n6962), .ZN(n6585) );
  INV_X1 U8236 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U8237 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7642) );
  OAI21_X1 U8238 ( .B1(n8724), .B2(n6583), .A(n7642), .ZN(n6584) );
  AOI21_X1 U8239 ( .B1(n9727), .B2(n6585), .A(n6584), .ZN(n6586) );
  OAI211_X1 U8240 ( .C1(n9731), .C2(n6588), .A(n6587), .B(n6586), .ZN(P2_U3255) );
  INV_X1 U8241 ( .A(n7803), .ZN(n6590) );
  OAI222_X1 U8242 ( .A1(n9495), .A2(n6589), .B1(n9493), .B2(n6590), .C1(n8097), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8243 ( .A1(n8979), .A2(n6591), .B1(n8980), .B2(n6590), .C1(
        P2_U3152), .C2(n9744), .ZN(P2_U3339) );
  INV_X1 U8244 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6604) );
  MUX2_X1 U8245 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n4536), .S(n7313), .Z(n6593)
         );
  INV_X1 U8246 ( .A(n6593), .ZN(n6594) );
  AOI211_X1 U8247 ( .C1(n6595), .C2(n6594), .A(n7306), .B(n9637), .ZN(n6596)
         );
  AOI21_X1 U8248 ( .B1(n9678), .B2(n7313), .A(n6596), .ZN(n6603) );
  INV_X1 U8249 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6597) );
  MUX2_X1 U8250 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6597), .S(n7313), .Z(n6600)
         );
  OAI21_X1 U8251 ( .B1(n7024), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6598), .ZN(
        n6599) );
  NAND2_X1 U8252 ( .A1(n6599), .A2(n6600), .ZN(n7312) );
  OAI21_X1 U8253 ( .B1(n6600), .B2(n6599), .A(n7312), .ZN(n6601) );
  AND2_X1 U8254 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7197) );
  AOI21_X1 U8255 ( .B1(n9686), .B2(n6601), .A(n7197), .ZN(n6602) );
  OAI211_X1 U8256 ( .C1(n9671), .C2(n6604), .A(n6603), .B(n6602), .ZN(P1_U3254) );
  INV_X1 U8257 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6623) );
  AND2_X1 U8258 ( .A1(n6606), .A2(n6605), .ZN(n6611) );
  OR2_X1 U8259 ( .A1(n6607), .A2(n6611), .ZN(n6608) );
  OR2_X1 U8260 ( .A1(n6609), .A2(n6608), .ZN(n6613) );
  OR2_X1 U8261 ( .A1(n6611), .A2(n6610), .ZN(n6612) );
  AND2_X1 U8262 ( .A1(n6613), .A2(n6612), .ZN(n6614) );
  NAND2_X1 U8263 ( .A1(n6678), .A2(n6697), .ZN(n7926) );
  NAND2_X1 U8264 ( .A1(n6677), .A2(n9113), .ZN(n7929) );
  NAND2_X1 U8265 ( .A1(n7926), .A2(n7929), .ZN(n8037) );
  OAI21_X1 U8266 ( .B1(n6614), .B2(n8037), .A(n6680), .ZN(n6703) );
  INV_X1 U8267 ( .A(n9468), .ZN(n9706) );
  AND2_X1 U8268 ( .A1(n8070), .A2(n7920), .ZN(n8062) );
  NAND2_X1 U8269 ( .A1(n6615), .A2(n8062), .ZN(n6616) );
  NAND2_X1 U8270 ( .A1(n6616), .A2(n8067), .ZN(n6674) );
  INV_X1 U8271 ( .A(n8037), .ZN(n6673) );
  XNOR2_X1 U8272 ( .A(n6674), .B(n6673), .ZN(n6617) );
  NAND2_X1 U8273 ( .A1(n6617), .A2(n9355), .ZN(n6619) );
  AOI22_X1 U8274 ( .A1(n9380), .A2(n9114), .B1(n9372), .B2(n9112), .ZN(n6618)
         );
  NAND2_X1 U8275 ( .A1(n6619), .A2(n6618), .ZN(n6700) );
  OAI211_X1 U8276 ( .C1(n6620), .C2(n6677), .A(n9437), .B(n6689), .ZN(n6699)
         );
  OAI21_X1 U8277 ( .B1(n6677), .B2(n9710), .A(n6699), .ZN(n6621) );
  AOI211_X1 U8278 ( .C1(n6703), .C2(n9706), .A(n6700), .B(n6621), .ZN(n6624)
         );
  OR2_X1 U8279 ( .A1(n6624), .A2(n9717), .ZN(n6622) );
  OAI21_X1 U8280 ( .B1(n9719), .B2(n6623), .A(n6622), .ZN(P1_U3475) );
  OR2_X1 U8281 ( .A1(n6624), .A2(n9724), .ZN(n6625) );
  OAI21_X1 U8282 ( .B1(n9561), .B2(n6336), .A(n6625), .ZN(P1_U3530) );
  OR2_X1 U8283 ( .A1(n8606), .A2(n6627), .ZN(n6628) );
  OAI211_X1 U8284 ( .C1(n8608), .C2(n6741), .A(n6629), .B(n6628), .ZN(n6634)
         );
  NAND2_X1 U8285 ( .A1(n8583), .A2(n6630), .ZN(n6631) );
  OAI21_X1 U8286 ( .B1(n8607), .B2(n6632), .A(n6631), .ZN(n6633) );
  NOR2_X1 U8287 ( .A1(n6634), .A2(n6633), .ZN(n6641) );
  NAND2_X1 U8288 ( .A1(n8601), .A2(n8637), .ZN(n6637) );
  OAI21_X1 U8289 ( .B1(n6638), .B2(n8587), .A(n6637), .ZN(n6639) );
  NAND3_X1 U8290 ( .A1(n6635), .A2(n4396), .A3(n6639), .ZN(n6640) );
  OAI211_X1 U8291 ( .C1(n6626), .C2(n8587), .A(n6641), .B(n6640), .ZN(P2_U3241) );
  NAND2_X1 U8292 ( .A1(n6642), .A2(n7896), .ZN(n6644) );
  AOI22_X1 U8293 ( .A1(n7804), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5941), .B2(
        n9628), .ZN(n6643) );
  NAND2_X1 U8294 ( .A1(n6644), .A2(n6643), .ZN(n6907) );
  NAND2_X1 U8295 ( .A1(n6907), .A2(n5930), .ZN(n6646) );
  NAND2_X1 U8296 ( .A1(n9112), .A2(n8508), .ZN(n6645) );
  NAND2_X1 U8297 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  XNOR2_X1 U8298 ( .A(n6647), .B(n6095), .ZN(n6661) );
  NAND2_X1 U8299 ( .A1(n6907), .A2(n8508), .ZN(n6652) );
  NAND2_X1 U8300 ( .A1(n9002), .A2(n9112), .ZN(n6651) );
  NAND2_X1 U8301 ( .A1(n6652), .A2(n6651), .ZN(n6654) );
  NAND2_X1 U8302 ( .A1(n6659), .A2(n6661), .ZN(n6658) );
  INV_X1 U8303 ( .A(n6658), .ZN(n6656) );
  NAND2_X1 U8304 ( .A1(n6656), .A2(n6657), .ZN(n6660) );
  AOI22_X1 U8305 ( .A1(n6661), .A2(n6660), .B1(n6713), .B2(n6659), .ZN(n6672)
         );
  AND2_X1 U8306 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9619) );
  INV_X1 U8307 ( .A(n6690), .ZN(n6668) );
  NAND2_X1 U8308 ( .A1(n7244), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U8309 ( .A1(n4305), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6666) );
  INV_X1 U8310 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U8311 ( .A1(n6662), .A2(n9896), .ZN(n6663) );
  AND2_X1 U8312 ( .A1(n6717), .A2(n6663), .ZN(n6788) );
  NAND2_X1 U8313 ( .A1(n7346), .A2(n6788), .ZN(n6665) );
  NAND2_X1 U8314 ( .A1(n7822), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6664) );
  NAND4_X1 U8315 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .ZN(n9111)
         );
  INV_X1 U8316 ( .A(n9111), .ZN(n6868) );
  OAI22_X1 U8317 ( .A1(n9050), .A2(n6668), .B1(n9095), .B2(n6868), .ZN(n6669)
         );
  AOI211_X1 U8318 ( .C1(n9092), .C2(n9113), .A(n9619), .B(n6669), .ZN(n6671)
         );
  NAND2_X1 U8319 ( .A1(n9084), .A2(n6907), .ZN(n6670) );
  OAI211_X1 U8320 ( .C1(n6672), .C2(n9086), .A(n6671), .B(n6670), .ZN(P1_U3219) );
  NAND2_X1 U8321 ( .A1(n6674), .A2(n6673), .ZN(n6675) );
  INV_X1 U8322 ( .A(n6907), .ZN(n6692) );
  NAND2_X1 U8323 ( .A1(n6692), .A2(n9112), .ZN(n7940) );
  INV_X1 U8324 ( .A(n9112), .ZN(n6676) );
  NAND2_X1 U8325 ( .A1(n6676), .A2(n6907), .ZN(n7933) );
  XNOR2_X1 U8326 ( .A(n6780), .B(n8036), .ZN(n6687) );
  OAI22_X1 U8327 ( .A1(n6678), .A2(n9331), .B1(n6868), .B2(n9329), .ZN(n6686)
         );
  NAND2_X1 U8328 ( .A1(n6678), .A2(n6677), .ZN(n6679) );
  NAND2_X1 U8329 ( .A1(n6682), .A2(n6681), .ZN(n6778) );
  NAND2_X1 U8330 ( .A1(n6683), .A2(n8036), .ZN(n6684) );
  NAND2_X1 U8331 ( .A1(n6778), .A2(n6684), .ZN(n6911) );
  NOR2_X1 U8332 ( .A1(n6911), .A2(n7354), .ZN(n6685) );
  AOI211_X1 U8333 ( .C1(n6687), .C2(n9355), .A(n6686), .B(n6685), .ZN(n6910)
         );
  INV_X1 U8334 ( .A(n6786), .ZN(n6688) );
  AOI21_X1 U8335 ( .B1(n6907), .B2(n6689), .A(n6688), .ZN(n6908) );
  AOI22_X1 U8336 ( .A1(n9356), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6690), .B2(
        n9343), .ZN(n6691) );
  OAI21_X1 U8337 ( .B1(n6692), .B2(n9364), .A(n6691), .ZN(n6694) );
  NOR2_X1 U8338 ( .A1(n6911), .A2(n7363), .ZN(n6693) );
  AOI211_X1 U8339 ( .C1(n6908), .C2(n9322), .A(n6694), .B(n6693), .ZN(n6695)
         );
  OAI21_X1 U8340 ( .B1(n6910), .B2(n9319), .A(n6695), .ZN(P1_U3283) );
  AOI22_X1 U8341 ( .A1(n9183), .A2(n6697), .B1(n6696), .B2(n9343), .ZN(n6698)
         );
  OAI21_X1 U8342 ( .B1(n6699), .B2(n7256), .A(n6698), .ZN(n6702) );
  MUX2_X1 U8343 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6700), .S(n9367), .Z(n6701)
         );
  AOI211_X1 U8344 ( .C1(n6704), .C2(n6703), .A(n6702), .B(n6701), .ZN(n6705)
         );
  INV_X1 U8345 ( .A(n6705), .ZN(P1_U3284) );
  NAND2_X1 U8346 ( .A1(n6706), .A2(n7896), .ZN(n6708) );
  AOI22_X1 U8347 ( .A1(n7804), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5941), .B2(
        n9642), .ZN(n6707) );
  NAND2_X1 U8348 ( .A1(n6708), .A2(n6707), .ZN(n6861) );
  INV_X1 U8349 ( .A(n6861), .ZN(n9711) );
  NAND2_X1 U8350 ( .A1(n6861), .A2(n5930), .ZN(n6710) );
  NAND2_X1 U8351 ( .A1(n9111), .A2(n8508), .ZN(n6709) );
  NAND2_X1 U8352 ( .A1(n6710), .A2(n6709), .ZN(n6711) );
  XNOR2_X1 U8353 ( .A(n6711), .B(n6095), .ZN(n6839) );
  AND2_X1 U8354 ( .A1(n9002), .A2(n9111), .ZN(n6712) );
  AOI21_X1 U8355 ( .B1(n6861), .B2(n8508), .A(n6712), .ZN(n6840) );
  XNOR2_X1 U8356 ( .A(n6839), .B(n6840), .ZN(n6714) );
  OAI21_X1 U8357 ( .B1(n6714), .B2(n6713), .A(n6843), .ZN(n6715) );
  NAND2_X1 U8358 ( .A1(n6715), .A2(n9088), .ZN(n6726) );
  AND2_X1 U8359 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9635) );
  INV_X1 U8360 ( .A(n6788), .ZN(n6723) );
  NAND2_X1 U8361 ( .A1(n7244), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U8362 ( .A1(n7869), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6721) );
  NAND2_X1 U8363 ( .A1(n6717), .A2(n6716), .ZN(n6718) );
  AND2_X1 U8364 ( .A1(n6851), .A2(n6718), .ZN(n6871) );
  NAND2_X1 U8365 ( .A1(n7346), .A2(n6871), .ZN(n6720) );
  NAND2_X1 U8366 ( .A1(n7822), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6719) );
  NAND4_X1 U8367 ( .A1(n6722), .A2(n6721), .A3(n6720), .A4(n6719), .ZN(n9110)
         );
  INV_X1 U8368 ( .A(n9110), .ZN(n6864) );
  OAI22_X1 U8369 ( .A1(n9050), .A2(n6723), .B1(n9095), .B2(n6864), .ZN(n6724)
         );
  AOI211_X1 U8370 ( .C1(n9092), .C2(n9112), .A(n9635), .B(n6724), .ZN(n6725)
         );
  OAI211_X1 U8371 ( .C1(n9711), .C2(n9102), .A(n6726), .B(n6725), .ZN(P1_U3229) );
  XNOR2_X1 U8372 ( .A(n9802), .B(n8195), .ZN(n6727) );
  NOR2_X1 U8373 ( .A1(n6820), .A2(n8187), .ZN(n6728) );
  NAND2_X1 U8374 ( .A1(n6727), .A2(n6728), .ZN(n6746) );
  INV_X1 U8375 ( .A(n6727), .ZN(n6793) );
  INV_X1 U8376 ( .A(n6728), .ZN(n6729) );
  NAND2_X1 U8377 ( .A1(n6793), .A2(n6729), .ZN(n6730) );
  AND2_X1 U8378 ( .A1(n6746), .A2(n6730), .ZN(n6735) );
  INV_X1 U8379 ( .A(n6735), .ZN(n6731) );
  AOI21_X1 U8380 ( .B1(n6734), .B2(n6731), .A(n8587), .ZN(n6738) );
  INV_X1 U8381 ( .A(n8601), .ZN(n8559) );
  NOR3_X1 U8382 ( .A1(n8559), .A2(n6732), .A3(n6741), .ZN(n6737) );
  NAND2_X1 U8383 ( .A1(n6736), .A2(n6735), .ZN(n6748) );
  OAI21_X1 U8384 ( .B1(n6738), .B2(n6737), .A(n6748), .ZN(n6745) );
  OAI21_X1 U8385 ( .B1(n8606), .B2(n6740), .A(n6739), .ZN(n6743) );
  OAI22_X1 U8386 ( .A1(n6741), .A2(n8607), .B1(n8608), .B2(n7655), .ZN(n6742)
         );
  AOI211_X1 U8387 ( .C1(n9802), .C2(n8583), .A(n6743), .B(n6742), .ZN(n6744)
         );
  NAND2_X1 U8388 ( .A1(n6745), .A2(n6744), .ZN(P2_U3223) );
  XNOR2_X1 U8389 ( .A(n6975), .B(n8173), .ZN(n6751) );
  NOR2_X1 U8390 ( .A1(n7655), .A2(n8187), .ZN(n6749) );
  XNOR2_X1 U8391 ( .A(n6751), .B(n6749), .ZN(n6803) );
  AND2_X1 U8392 ( .A1(n6803), .A2(n6746), .ZN(n6747) );
  NAND2_X1 U8393 ( .A1(n6748), .A2(n6747), .ZN(n6796) );
  INV_X1 U8394 ( .A(n6749), .ZN(n6750) );
  NAND2_X1 U8395 ( .A1(n6751), .A2(n6750), .ZN(n6752) );
  XNOR2_X1 U8396 ( .A(n5207), .B(n8195), .ZN(n6753) );
  NOR2_X1 U8397 ( .A1(n6819), .A2(n8187), .ZN(n6754) );
  NAND2_X1 U8398 ( .A1(n6753), .A2(n6754), .ZN(n6760) );
  INV_X1 U8399 ( .A(n6753), .ZN(n6759) );
  INV_X1 U8400 ( .A(n6754), .ZN(n6755) );
  NAND2_X1 U8401 ( .A1(n6759), .A2(n6755), .ZN(n6756) );
  NAND2_X1 U8402 ( .A1(n6760), .A2(n6756), .ZN(n7646) );
  XNOR2_X1 U8403 ( .A(n7007), .B(n8173), .ZN(n6882) );
  NOR2_X1 U8404 ( .A1(n7656), .A2(n8187), .ZN(n6883) );
  XNOR2_X1 U8405 ( .A(n6882), .B(n6883), .ZN(n6762) );
  INV_X1 U8406 ( .A(n6762), .ZN(n6758) );
  AOI21_X1 U8407 ( .B1(n6761), .B2(n6758), .A(n8587), .ZN(n6765) );
  NOR3_X1 U8408 ( .A1(n8559), .A2(n6759), .A3(n6819), .ZN(n6764) );
  NAND2_X1 U8409 ( .A1(n6763), .A2(n6762), .ZN(n6886) );
  OAI21_X1 U8410 ( .B1(n6765), .B2(n6764), .A(n6886), .ZN(n6769) );
  OAI22_X1 U8411 ( .A1(n8606), .A2(n6901), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5216), .ZN(n6767) );
  OAI22_X1 U8412 ( .A1(n7108), .A2(n8608), .B1(n8607), .B2(n6819), .ZN(n6766)
         );
  AOI211_X1 U8413 ( .C1(n7007), .C2(n8583), .A(n6767), .B(n6766), .ZN(n6768)
         );
  NAND2_X1 U8414 ( .A1(n6769), .A2(n6768), .ZN(P2_U3238) );
  OAI22_X1 U8415 ( .A1(n8559), .A2(n6771), .B1(n6770), .B2(n8587), .ZN(n6773)
         );
  NAND2_X1 U8416 ( .A1(n6773), .A2(n6772), .ZN(n6775) );
  INV_X1 U8417 ( .A(n8608), .ZN(n7681) );
  AOI22_X1 U8418 ( .A1(n7681), .A2(n6391), .B1(n9762), .B2(n8583), .ZN(n6774)
         );
  OAI211_X1 U8419 ( .C1(n7678), .C2(n6776), .A(n6775), .B(n6774), .ZN(P2_U3234) );
  NAND2_X1 U8420 ( .A1(n6907), .A2(n9112), .ZN(n6777) );
  OR2_X1 U8421 ( .A1(n6861), .A2(n6868), .ZN(n7939) );
  NAND2_X1 U8422 ( .A1(n6861), .A2(n6868), .ZN(n7934) );
  NAND2_X1 U8423 ( .A1(n7939), .A2(n7934), .ZN(n8038) );
  INV_X1 U8424 ( .A(n8038), .ZN(n6779) );
  XNOR2_X1 U8425 ( .A(n6863), .B(n6779), .ZN(n9714) );
  INV_X1 U8426 ( .A(n7933), .ZN(n7941) );
  XNOR2_X1 U8427 ( .A(n6943), .B(n8038), .ZN(n6781) );
  NAND2_X1 U8428 ( .A1(n6781), .A2(n9355), .ZN(n6783) );
  AOI22_X1 U8429 ( .A1(n9380), .A2(n9112), .B1(n9372), .B2(n9110), .ZN(n6782)
         );
  NAND2_X1 U8430 ( .A1(n6783), .A2(n6782), .ZN(n6784) );
  AOI21_X1 U8431 ( .B1(n9714), .B2(n7158), .A(n6784), .ZN(n9716) );
  NAND2_X1 U8432 ( .A1(n6786), .A2(n6861), .ZN(n6785) );
  NAND2_X1 U8433 ( .A1(n6785), .A2(n9437), .ZN(n6787) );
  OR2_X1 U8434 ( .A1(n6787), .A2(n6869), .ZN(n9709) );
  AOI22_X1 U8435 ( .A1(n9356), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6788), .B2(
        n9343), .ZN(n6790) );
  NAND2_X1 U8436 ( .A1(n9183), .A2(n6861), .ZN(n6789) );
  OAI211_X1 U8437 ( .C1(n9709), .C2(n7256), .A(n6790), .B(n6789), .ZN(n6791)
         );
  AOI21_X1 U8438 ( .B1(n9714), .B2(n7165), .A(n6791), .ZN(n6792) );
  OAI21_X1 U8439 ( .B1(n9716), .B2(n9319), .A(n6792), .ZN(P1_U3282) );
  INV_X1 U8440 ( .A(n6748), .ZN(n6795) );
  NOR3_X1 U8441 ( .A1(n8559), .A2(n6793), .A3(n6820), .ZN(n6794) );
  AOI21_X1 U8442 ( .B1(n6795), .B2(n8604), .A(n6794), .ZN(n6804) );
  NOR2_X1 U8443 ( .A1(n6796), .A2(n8587), .ZN(n6801) );
  AND2_X1 U8444 ( .A1(n8583), .A2(n6975), .ZN(n6800) );
  OAI21_X1 U8445 ( .B1(n8606), .B2(n6830), .A(n6797), .ZN(n6799) );
  OAI22_X1 U8446 ( .A1(n6820), .A2(n8607), .B1(n8608), .B2(n6819), .ZN(n6798)
         );
  NOR4_X1 U8447 ( .A1(n6801), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(n6802)
         );
  OAI21_X1 U8448 ( .B1(n6804), .B2(n6803), .A(n6802), .ZN(P2_U3233) );
  OAI21_X1 U8449 ( .B1(n6806), .B2(n6805), .A(n8229), .ZN(n6815) );
  INV_X1 U8450 ( .A(n6806), .ZN(n6808) );
  NAND3_X1 U8451 ( .A1(n8601), .A2(n6808), .A3(n6807), .ZN(n6809) );
  AOI21_X1 U8452 ( .B1(n6809), .B2(n8607), .A(n5100), .ZN(n6814) );
  AOI22_X1 U8453 ( .A1(n7681), .A2(n8637), .B1(n9785), .B2(n8583), .ZN(n6811)
         );
  OAI211_X1 U8454 ( .C1(n6812), .C2(n8606), .A(n6811), .B(n6810), .ZN(n6813)
         );
  AOI211_X1 U8455 ( .C1(n8604), .C2(n6815), .A(n6814), .B(n6813), .ZN(n6816)
         );
  INV_X1 U8456 ( .A(n6816), .ZN(P2_U3232) );
  INV_X1 U8457 ( .A(n7660), .ZN(n6826) );
  OAI21_X1 U8458 ( .B1(n6818), .B2(n8261), .A(n6817), .ZN(n6974) );
  OAI22_X1 U8459 ( .A1(n6820), .A2(n8859), .B1(n6819), .B2(n8861), .ZN(n6825)
         );
  OR2_X1 U8460 ( .A1(n6821), .A2(n8346), .ZN(n6822) );
  NAND2_X1 U8461 ( .A1(n6822), .A2(n8347), .ZN(n7652) );
  XNOR2_X1 U8462 ( .A(n7652), .B(n8261), .ZN(n6823) );
  NOR2_X1 U8463 ( .A1(n6823), .A2(n8857), .ZN(n6824) );
  AOI211_X1 U8464 ( .C1(n6826), .C2(n6974), .A(n6825), .B(n6824), .ZN(n6978)
         );
  INV_X1 U8465 ( .A(n7663), .ZN(n6827) );
  AOI21_X1 U8466 ( .B1(n6975), .B2(n6828), .A(n6827), .ZN(n6976) );
  INV_X1 U8467 ( .A(n6975), .ZN(n6829) );
  NOR2_X1 U8468 ( .A1(n8869), .A2(n6829), .ZN(n6833) );
  OAI22_X1 U8469 ( .A1(n8826), .A2(n6831), .B1(n6830), .B2(n9742), .ZN(n6832)
         );
  AOI211_X1 U8470 ( .C1(n6976), .C2(n8864), .A(n6833), .B(n6832), .ZN(n6835)
         );
  NAND2_X1 U8471 ( .A1(n6974), .A2(n7333), .ZN(n6834) );
  OAI211_X1 U8472 ( .C1(n6978), .C2(n9752), .A(n6835), .B(n6834), .ZN(P2_U3287) );
  INV_X1 U8473 ( .A(n6836), .ZN(n8206) );
  OAI222_X1 U8474 ( .A1(n9495), .A2(n7788), .B1(P1_U3084), .B2(n5899), .C1(
        n9493), .C2(n8206), .ZN(P1_U3333) );
  NAND2_X1 U8475 ( .A1(n5725), .A2(n7896), .ZN(n6838) );
  AOI22_X1 U8476 ( .A1(n7804), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5941), .B2(
        n9125), .ZN(n6837) );
  NAND2_X1 U8477 ( .A1(n6838), .A2(n6837), .ZN(n7068) );
  INV_X1 U8478 ( .A(n7068), .ZN(n6874) );
  INV_X1 U8479 ( .A(n6839), .ZN(n6841) );
  NAND2_X1 U8480 ( .A1(n6841), .A2(n6840), .ZN(n6842) );
  AND2_X1 U8481 ( .A1(n9002), .A2(n9110), .ZN(n6844) );
  AOI21_X1 U8482 ( .B1(n7068), .B2(n8508), .A(n6844), .ZN(n6916) );
  NAND2_X1 U8483 ( .A1(n7068), .A2(n5930), .ZN(n6846) );
  NAND2_X1 U8484 ( .A1(n9110), .A2(n8508), .ZN(n6845) );
  NAND2_X1 U8485 ( .A1(n6846), .A2(n6845), .ZN(n6847) );
  XNOR2_X1 U8486 ( .A(n6847), .B(n8482), .ZN(n6917) );
  XOR2_X1 U8487 ( .A(n6916), .B(n6917), .Z(n6848) );
  XNOR2_X1 U8488 ( .A(n6919), .B(n6848), .ZN(n6849) );
  NAND2_X1 U8489 ( .A1(n6849), .A2(n9088), .ZN(n6860) );
  NAND2_X1 U8490 ( .A1(n7869), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U8491 ( .A1(n7822), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6855) );
  INV_X1 U8492 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U8493 ( .A1(n6851), .A2(n6850), .ZN(n6852) );
  AND2_X1 U8494 ( .A1(n6928), .A2(n6852), .ZN(n6951) );
  NAND2_X1 U8495 ( .A1(n7346), .A2(n6951), .ZN(n6854) );
  NAND2_X1 U8496 ( .A1(n7244), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6853) );
  NAND4_X1 U8497 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n9109)
         );
  AND2_X1 U8498 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9126) );
  INV_X1 U8499 ( .A(n6871), .ZN(n6857) );
  OAI22_X1 U8500 ( .A1(n9051), .A2(n6868), .B1(n9050), .B2(n6857), .ZN(n6858)
         );
  AOI211_X1 U8501 ( .C1(n9073), .C2(n9109), .A(n9126), .B(n6858), .ZN(n6859)
         );
  OAI211_X1 U8502 ( .C1(n6874), .C2(n9102), .A(n6860), .B(n6859), .ZN(P1_U3215) );
  AND2_X1 U8503 ( .A1(n6861), .A2(n9111), .ZN(n6862) );
  OR2_X1 U8504 ( .A1(n7068), .A2(n6864), .ZN(n7938) );
  NAND2_X1 U8505 ( .A1(n7068), .A2(n6864), .ZN(n7937) );
  NAND2_X1 U8506 ( .A1(n7938), .A2(n7937), .ZN(n7015) );
  INV_X1 U8507 ( .A(n7015), .ZN(n8041) );
  XNOR2_X1 U8508 ( .A(n7022), .B(n8041), .ZN(n7070) );
  INV_X1 U8509 ( .A(n9109), .ZN(n7834) );
  INV_X1 U8510 ( .A(n7939), .ZN(n6865) );
  OAI21_X1 U8511 ( .B1(n6943), .B2(n6865), .A(n7934), .ZN(n6866) );
  XNOR2_X1 U8512 ( .A(n6866), .B(n7015), .ZN(n6867) );
  OAI222_X1 U8513 ( .A1(n9329), .A2(n7834), .B1(n9331), .B2(n6868), .C1(n6867), 
        .C2(n9374), .ZN(n7066) );
  INV_X1 U8514 ( .A(n6869), .ZN(n6870) );
  AND2_X1 U8515 ( .A1(n6869), .A2(n6874), .ZN(n6949) );
  AOI211_X1 U8516 ( .C1(n7068), .C2(n6870), .A(n9696), .B(n6949), .ZN(n7067)
         );
  NAND2_X1 U8517 ( .A1(n7067), .A2(n9370), .ZN(n6873) );
  AOI22_X1 U8518 ( .A1(n9356), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n6871), .B2(
        n9343), .ZN(n6872) );
  OAI211_X1 U8519 ( .C1(n6874), .C2(n9364), .A(n6873), .B(n6872), .ZN(n6875)
         );
  AOI21_X1 U8520 ( .B1(n7066), .B2(n9367), .A(n6875), .ZN(n6876) );
  OAI21_X1 U8521 ( .B1(n7070), .B2(n9383), .A(n6876), .ZN(P1_U3281) );
  INV_X1 U8522 ( .A(n7780), .ZN(n6939) );
  OAI222_X1 U8523 ( .A1(n8979), .A2(n6877), .B1(n8233), .B2(n6939), .C1(n8284), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  XNOR2_X1 U8524 ( .A(n7128), .B(n8173), .ZN(n6878) );
  OR2_X1 U8525 ( .A1(n7108), .A2(n8187), .ZN(n6879) );
  NAND2_X1 U8526 ( .A1(n6878), .A2(n6879), .ZN(n6983) );
  INV_X1 U8527 ( .A(n6878), .ZN(n6881) );
  INV_X1 U8528 ( .A(n6879), .ZN(n6880) );
  NAND2_X1 U8529 ( .A1(n6881), .A2(n6880), .ZN(n7366) );
  NAND2_X1 U8530 ( .A1(n6983), .A2(n7366), .ZN(n6887) );
  INV_X1 U8531 ( .A(n6882), .ZN(n6884) );
  NAND2_X1 U8532 ( .A1(n6884), .A2(n6883), .ZN(n6885) );
  XOR2_X1 U8533 ( .A(n6887), .B(n6984), .Z(n6892) );
  AOI22_X1 U8534 ( .A1(n7566), .A2(n8631), .B1(n8629), .B2(n7567), .ZN(n6995)
         );
  OAI22_X1 U8535 ( .A1(n6888), .A2(n6995), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7058), .ZN(n6890) );
  NOR2_X1 U8536 ( .A1(n8606), .A2(n7000), .ZN(n6889) );
  AOI211_X1 U8537 ( .C1(n7128), .C2(n8583), .A(n6890), .B(n6889), .ZN(n6891)
         );
  OAI21_X1 U8538 ( .B1(n6892), .B2(n8587), .A(n6891), .ZN(P2_U3226) );
  NAND2_X1 U8539 ( .A1(n6893), .A2(n6894), .ZN(n6895) );
  XNOR2_X1 U8540 ( .A(n6895), .B(n8264), .ZN(n7011) );
  XOR2_X1 U8541 ( .A(n6896), .B(n8264), .Z(n6897) );
  AOI222_X1 U8542 ( .A1(n8817), .A2(n6897), .B1(n8632), .B2(n7566), .C1(n8630), 
        .C2(n7567), .ZN(n7010) );
  OR2_X1 U8543 ( .A1(n7010), .A2(n9752), .ZN(n6906) );
  INV_X1 U8544 ( .A(n6898), .ZN(n7665) );
  INV_X1 U8545 ( .A(n6997), .ZN(n6899) );
  AOI21_X1 U8546 ( .B1(n7007), .B2(n7665), .A(n6899), .ZN(n7008) );
  NOR2_X1 U8547 ( .A1(n6900), .A2(n8869), .ZN(n6904) );
  OAI22_X1 U8548 ( .A1(n8826), .A2(n6902), .B1(n6901), .B2(n9742), .ZN(n6903)
         );
  AOI211_X1 U8549 ( .C1(n7008), .C2(n8864), .A(n6904), .B(n6903), .ZN(n6905)
         );
  OAI211_X1 U8550 ( .C1(n7011), .C2(n8873), .A(n6906), .B(n6905), .ZN(P2_U3285) );
  AOI22_X1 U8551 ( .A1(n6908), .A2(n9437), .B1(n9465), .B2(n6907), .ZN(n6909)
         );
  OAI211_X1 U8552 ( .C1(n9535), .C2(n6911), .A(n6910), .B(n6909), .ZN(n6913)
         );
  NAND2_X1 U8553 ( .A1(n6913), .A2(n9561), .ZN(n6912) );
  OAI21_X1 U8554 ( .B1(n9561), .B2(n6335), .A(n6912), .ZN(P1_U3531) );
  INV_X1 U8555 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U8556 ( .A1(n6913), .A2(n9719), .ZN(n6914) );
  OAI21_X1 U8557 ( .B1(n9719), .B2(n6915), .A(n6914), .ZN(P1_U3478) );
  AND2_X1 U8558 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  OAI22_X1 U8559 ( .A1(n6919), .A2(n6918), .B1(n6917), .B2(n6916), .ZN(n7090)
         );
  NAND2_X1 U8560 ( .A1(n6920), .A2(n7896), .ZN(n6922) );
  AOI22_X1 U8561 ( .A1(n7804), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5941), .B2(
        n9646), .ZN(n6921) );
  NAND2_X1 U8562 ( .A1(n7835), .A2(n5930), .ZN(n6924) );
  NAND2_X1 U8563 ( .A1(n9109), .A2(n8508), .ZN(n6923) );
  NAND2_X1 U8564 ( .A1(n6924), .A2(n6923), .ZN(n6925) );
  XNOR2_X1 U8565 ( .A(n6925), .B(n6095), .ZN(n7093) );
  AND2_X1 U8566 ( .A1(n9002), .A2(n9109), .ZN(n6926) );
  AOI21_X1 U8567 ( .B1(n7835), .B2(n8508), .A(n6926), .ZN(n7091) );
  XNOR2_X1 U8568 ( .A(n7093), .B(n7091), .ZN(n7089) );
  XNOR2_X1 U8569 ( .A(n7090), .B(n7089), .ZN(n6938) );
  AND2_X1 U8570 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9645) );
  INV_X1 U8571 ( .A(n6951), .ZN(n6934) );
  NAND2_X1 U8572 ( .A1(n7244), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U8573 ( .A1(n7869), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6932) );
  NAND2_X1 U8574 ( .A1(n6928), .A2(n6927), .ZN(n6929) );
  AND2_X1 U8575 ( .A1(n7029), .A2(n6929), .ZN(n7100) );
  NAND2_X1 U8576 ( .A1(n7346), .A2(n7100), .ZN(n6931) );
  NAND2_X1 U8577 ( .A1(n7822), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6930) );
  NAND4_X1 U8578 ( .A1(n6933), .A2(n6932), .A3(n6931), .A4(n6930), .ZN(n9108)
         );
  INV_X1 U8579 ( .A(n9108), .ZN(n7027) );
  OAI22_X1 U8580 ( .A1(n9050), .A2(n6934), .B1(n9095), .B2(n7027), .ZN(n6935)
         );
  AOI211_X1 U8581 ( .C1(n9092), .C2(n9110), .A(n9645), .B(n6935), .ZN(n6937)
         );
  NAND2_X1 U8582 ( .A1(n7835), .A2(n9084), .ZN(n6936) );
  OAI211_X1 U8583 ( .C1(n6938), .C2(n9086), .A(n6937), .B(n6936), .ZN(P1_U3234) );
  INV_X1 U8584 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7781) );
  OAI222_X1 U8585 ( .A1(n9495), .A2(n7781), .B1(P1_U3084), .B2(n8092), .C1(
        n9493), .C2(n6939), .ZN(P1_U3332) );
  NAND2_X1 U8586 ( .A1(n7022), .A2(n7015), .ZN(n6940) );
  OR2_X1 U8587 ( .A1(n7068), .A2(n9110), .ZN(n7018) );
  NAND2_X1 U8588 ( .A1(n6940), .A2(n7018), .ZN(n6942) );
  XNOR2_X1 U8589 ( .A(n7835), .B(n9109), .ZN(n8040) );
  INV_X1 U8590 ( .A(n8040), .ZN(n6941) );
  XNOR2_X1 U8591 ( .A(n6942), .B(n6941), .ZN(n9557) );
  NAND2_X1 U8592 ( .A1(n7938), .A2(n7939), .ZN(n7936) );
  NAND2_X1 U8593 ( .A1(n7937), .A2(n7934), .ZN(n7943) );
  NAND2_X1 U8594 ( .A1(n7943), .A2(n7938), .ZN(n7848) );
  NAND2_X1 U8595 ( .A1(n6945), .A2(n8040), .ZN(n7035) );
  OAI211_X1 U8596 ( .C1(n6945), .C2(n8040), .A(n7035), .B(n9355), .ZN(n6947)
         );
  AOI22_X1 U8597 ( .A1(n9380), .A2(n9110), .B1(n9372), .B2(n9108), .ZN(n6946)
         );
  NAND2_X1 U8598 ( .A1(n6947), .A2(n6946), .ZN(n6948) );
  AOI21_X1 U8599 ( .B1(n9557), .B2(n7158), .A(n6948), .ZN(n9559) );
  INV_X1 U8600 ( .A(n7835), .ZN(n9554) );
  OR2_X1 U8601 ( .A1(n6949), .A2(n9554), .ZN(n6950) );
  NAND2_X1 U8602 ( .A1(n7037), .A2(n6950), .ZN(n9555) );
  AOI22_X1 U8603 ( .A1(n9356), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n6951), .B2(
        n9343), .ZN(n6953) );
  NAND2_X1 U8604 ( .A1(n9183), .A2(n7835), .ZN(n6952) );
  OAI211_X1 U8605 ( .C1(n9555), .C2(n9186), .A(n6953), .B(n6952), .ZN(n6954)
         );
  AOI21_X1 U8606 ( .B1(n9557), .B2(n7165), .A(n6954), .ZN(n6955) );
  OAI21_X1 U8607 ( .B1(n9559), .B2(n9319), .A(n6955), .ZN(P1_U3280) );
  NAND2_X1 U8608 ( .A1(n6963), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U8609 ( .A1(n6957), .A2(n6956), .ZN(n6960) );
  MUX2_X1 U8610 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n6902), .S(n7054), .Z(n6958)
         );
  INV_X1 U8611 ( .A(n6958), .ZN(n6959) );
  NOR2_X1 U8612 ( .A1(n6960), .A2(n6959), .ZN(n7048) );
  AOI21_X1 U8613 ( .B1(n6960), .B2(n6959), .A(n7048), .ZN(n6973) );
  INV_X1 U8614 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6961) );
  MUX2_X1 U8615 ( .A(n6961), .B(P2_REG1_REG_11__SCAN_IN), .S(n7054), .Z(n6965)
         );
  AOI21_X1 U8616 ( .B1(n6965), .B2(n6964), .A(n7053), .ZN(n6966) );
  NAND2_X1 U8617 ( .A1(n9727), .A2(n6966), .ZN(n6969) );
  NOR2_X1 U8618 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5216), .ZN(n6967) );
  AOI21_X1 U8619 ( .B1(n9729), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6967), .ZN(
        n6968) );
  OAI211_X1 U8620 ( .C1(n9731), .C2(n6970), .A(n6969), .B(n6968), .ZN(n6971)
         );
  INV_X1 U8621 ( .A(n6971), .ZN(n6972) );
  OAI21_X1 U8622 ( .B1(n6973), .B2(n9730), .A(n6972), .ZN(P2_U3256) );
  INV_X1 U8623 ( .A(n6974), .ZN(n6979) );
  AOI22_X1 U8624 ( .A1(n6976), .A2(n9786), .B1(n9772), .B2(n6975), .ZN(n6977)
         );
  OAI211_X1 U8625 ( .C1(n6979), .C2(n9778), .A(n6978), .B(n6977), .ZN(n6981)
         );
  NAND2_X1 U8626 ( .A1(n6981), .A2(n9817), .ZN(n6980) );
  OAI21_X1 U8627 ( .B1(n9817), .B2(n5185), .A(n6980), .ZN(P2_U3478) );
  NAND2_X1 U8628 ( .A1(n6981), .A2(n9830), .ZN(n6982) );
  OAI21_X1 U8629 ( .B1(n9830), .B2(n6376), .A(n6982), .ZN(P2_U3529) );
  XNOR2_X1 U8630 ( .A(n8952), .B(n8173), .ZN(n7205) );
  NOR2_X1 U8631 ( .A1(n7211), .A2(n8187), .ZN(n7206) );
  XNOR2_X1 U8632 ( .A(n7205), .B(n7206), .ZN(n7376) );
  XNOR2_X1 U8633 ( .A(n7385), .B(n7376), .ZN(n6988) );
  OAI22_X1 U8634 ( .A1(n8606), .A2(n7119), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7227), .ZN(n6986) );
  OAI22_X1 U8635 ( .A1(n7108), .A2(n8607), .B1(n8608), .B2(n7261), .ZN(n6985)
         );
  AOI211_X1 U8636 ( .C1(n8952), .C2(n8583), .A(n6986), .B(n6985), .ZN(n6987)
         );
  OAI21_X1 U8637 ( .B1(n6988), .B2(n8587), .A(n6987), .ZN(P2_U3236) );
  NAND2_X1 U8638 ( .A1(n6893), .A2(n6989), .ZN(n6991) );
  AND2_X1 U8639 ( .A1(n6991), .A2(n6990), .ZN(n6992) );
  XOR2_X1 U8640 ( .A(n8266), .B(n6992), .Z(n7130) );
  NAND2_X1 U8641 ( .A1(n6993), .A2(n8338), .ZN(n6994) );
  XNOR2_X1 U8642 ( .A(n6994), .B(n8266), .ZN(n6996) );
  OAI21_X1 U8643 ( .B1(n6996), .B2(n8857), .A(n6995), .ZN(n7126) );
  AOI21_X1 U8644 ( .B1(n6997), .B2(n7128), .A(n9810), .ZN(n6998) );
  AND2_X1 U8645 ( .A1(n6998), .A2(n7116), .ZN(n7127) );
  INV_X1 U8646 ( .A(n8831), .ZN(n6999) );
  NAND2_X1 U8647 ( .A1(n7127), .A2(n6999), .ZN(n7003) );
  OAI22_X1 U8648 ( .A1(n8826), .A2(n7050), .B1(n7000), .B2(n9742), .ZN(n7001)
         );
  AOI21_X1 U8649 ( .B1(n7128), .B2(n8828), .A(n7001), .ZN(n7002) );
  NAND2_X1 U8650 ( .A1(n7003), .A2(n7002), .ZN(n7004) );
  AOI21_X1 U8651 ( .B1(n7126), .B2(n8826), .A(n7004), .ZN(n7005) );
  OAI21_X1 U8652 ( .B1(n7130), .B2(n8873), .A(n7005), .ZN(P2_U3284) );
  INV_X1 U8653 ( .A(n7768), .ZN(n7640) );
  OAI222_X1 U8654 ( .A1(n8979), .A2(n7006), .B1(n8233), .B2(n7640), .C1(
        P2_U3152), .C2(n5517), .ZN(P2_U3336) );
  AOI22_X1 U8655 ( .A1(n7008), .A2(n9786), .B1(n9772), .B2(n7007), .ZN(n7009)
         );
  OAI211_X1 U8656 ( .C1(n9790), .C2(n7011), .A(n7010), .B(n7009), .ZN(n7013)
         );
  NAND2_X1 U8657 ( .A1(n7013), .A2(n9830), .ZN(n7012) );
  OAI21_X1 U8658 ( .B1(n9830), .B2(n6961), .A(n7012), .ZN(P2_U3531) );
  NAND2_X1 U8659 ( .A1(n7013), .A2(n9817), .ZN(n7014) );
  OAI21_X1 U8660 ( .B1(n9817), .B2(n5214), .A(n7014), .ZN(P2_U3484) );
  NAND2_X1 U8661 ( .A1(n7835), .A2(n9109), .ZN(n7016) );
  AND2_X1 U8662 ( .A1(n7015), .A2(n7016), .ZN(n7021) );
  INV_X1 U8663 ( .A(n7016), .ZN(n7020) );
  OR2_X1 U8664 ( .A1(n7835), .A2(n9109), .ZN(n7017) );
  AND2_X1 U8665 ( .A1(n7018), .A2(n7017), .ZN(n7019) );
  NAND2_X1 U8666 ( .A1(n7023), .A2(n7896), .ZN(n7026) );
  AOI22_X1 U8667 ( .A1(n7804), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5941), .B2(
        n7024), .ZN(n7025) );
  OR2_X1 U8668 ( .A1(n9464), .A2(n7027), .ZN(n7950) );
  NAND2_X1 U8669 ( .A1(n9464), .A2(n7027), .ZN(n7949) );
  NAND2_X1 U8670 ( .A1(n7950), .A2(n7949), .ZN(n7136) );
  XNOR2_X1 U8671 ( .A(n7137), .B(n7136), .ZN(n9467) );
  NAND2_X1 U8672 ( .A1(n7244), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7034) );
  NAND2_X1 U8673 ( .A1(n7869), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8674 ( .A1(n7029), .A2(n7028), .ZN(n7030) );
  AND2_X1 U8675 ( .A1(n7149), .A2(n7030), .ZN(n7194) );
  NAND2_X1 U8676 ( .A1(n7346), .A2(n7194), .ZN(n7032) );
  NAND2_X1 U8677 ( .A1(n7822), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7031) );
  NAND4_X1 U8678 ( .A1(n7034), .A2(n7033), .A3(n7032), .A4(n7031), .ZN(n9107)
         );
  OR2_X1 U8679 ( .A1(n7835), .A2(n7834), .ZN(n7142) );
  INV_X1 U8680 ( .A(n7136), .ZN(n8042) );
  XNOR2_X1 U8681 ( .A(n7141), .B(n8042), .ZN(n7036) );
  OAI222_X1 U8682 ( .A1(n9331), .A2(n7834), .B1(n9329), .B2(n7237), .C1(n9374), 
        .C2(n7036), .ZN(n9462) );
  INV_X1 U8683 ( .A(n9464), .ZN(n7040) );
  AOI211_X1 U8684 ( .C1(n9464), .C2(n7037), .A(n9696), .B(n7160), .ZN(n9463)
         );
  NAND2_X1 U8685 ( .A1(n9463), .A2(n9370), .ZN(n7039) );
  AOI22_X1 U8686 ( .A1(n9356), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7100), .B2(
        n9343), .ZN(n7038) );
  OAI211_X1 U8687 ( .C1(n7040), .C2(n9364), .A(n7039), .B(n7038), .ZN(n7041)
         );
  AOI21_X1 U8688 ( .B1(n9462), .B2(n9367), .A(n7041), .ZN(n7042) );
  OAI21_X1 U8689 ( .B1(n9467), .B2(n9383), .A(n7042), .ZN(P1_U3279) );
  NAND2_X1 U8690 ( .A1(n7816), .A2(n7043), .ZN(n7044) );
  OAI211_X1 U8691 ( .C1(n9886), .C2(n8979), .A(n7044), .B(n8457), .ZN(P2_U3335) );
  NAND2_X1 U8692 ( .A1(n7816), .A2(n7045), .ZN(n7047) );
  NAND2_X1 U8693 ( .A1(n7046), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8112) );
  OAI211_X1 U8694 ( .C1(n7817), .C2(n9495), .A(n7047), .B(n8112), .ZN(P1_U3330) );
  NOR2_X1 U8695 ( .A1(n7054), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7049) );
  NOR2_X1 U8696 ( .A1(n7049), .A2(n7048), .ZN(n7052) );
  MUX2_X1 U8697 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7050), .S(n7222), .Z(n7051)
         );
  NAND2_X1 U8698 ( .A1(n7222), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7218) );
  OAI211_X1 U8699 ( .C1(n7222), .C2(P2_REG2_REG_12__SCAN_IN), .A(n7052), .B(
        n7218), .ZN(n7217) );
  OAI211_X1 U8700 ( .C1(n7052), .C2(n7051), .A(n7217), .B(n9728), .ZN(n7064)
         );
  MUX2_X1 U8701 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7055), .S(n7222), .Z(n7056)
         );
  OAI21_X1 U8702 ( .B1(n7057), .B2(n7056), .A(n7224), .ZN(n7062) );
  INV_X1 U8703 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7060) );
  OR2_X1 U8704 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7058), .ZN(n7059) );
  OAI21_X1 U8705 ( .B1(n8724), .B2(n7060), .A(n7059), .ZN(n7061) );
  AOI21_X1 U8706 ( .B1(n9727), .B2(n7062), .A(n7061), .ZN(n7063) );
  OAI211_X1 U8707 ( .C1(n9731), .C2(n7065), .A(n7064), .B(n7063), .ZN(P2_U3257) );
  INV_X1 U8708 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7072) );
  AOI211_X1 U8709 ( .C1(n9465), .C2(n7068), .A(n7067), .B(n7066), .ZN(n7069)
         );
  OAI21_X1 U8710 ( .B1(n9468), .B2(n7070), .A(n7069), .ZN(n7073) );
  NAND2_X1 U8711 ( .A1(n7073), .A2(n9561), .ZN(n7071) );
  OAI21_X1 U8712 ( .B1(n9561), .B2(n7072), .A(n7071), .ZN(P1_U3533) );
  INV_X1 U8713 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7075) );
  NAND2_X1 U8714 ( .A1(n7073), .A2(n9719), .ZN(n7074) );
  OAI21_X1 U8715 ( .B1(n9719), .B2(n7075), .A(n7074), .ZN(P1_U3484) );
  INV_X1 U8716 ( .A(n7861), .ZN(n7078) );
  OAI222_X1 U8717 ( .A1(P2_U3152), .A2(n7077), .B1(n8233), .B2(n7078), .C1(
        n7076), .C2(n8979), .ZN(P2_U3334) );
  OAI222_X1 U8718 ( .A1(n9495), .A2(n7862), .B1(P1_U3084), .B2(n7079), .C1(
        n9493), .C2(n7078), .ZN(P1_U3329) );
  NAND2_X1 U8719 ( .A1(n9464), .A2(n5930), .ZN(n7081) );
  NAND2_X1 U8720 ( .A1(n9108), .A2(n8508), .ZN(n7080) );
  NAND2_X1 U8721 ( .A1(n7081), .A2(n7080), .ZN(n7082) );
  XNOR2_X1 U8722 ( .A(n7082), .B(n8482), .ZN(n7084) );
  AND2_X1 U8723 ( .A1(n9002), .A2(n9108), .ZN(n7083) );
  AOI21_X1 U8724 ( .B1(n9464), .B2(n8508), .A(n7083), .ZN(n7085) );
  NAND2_X1 U8725 ( .A1(n7084), .A2(n7085), .ZN(n7181) );
  INV_X1 U8726 ( .A(n7084), .ZN(n7087) );
  INV_X1 U8727 ( .A(n7085), .ZN(n7086) );
  NAND2_X1 U8728 ( .A1(n7087), .A2(n7086), .ZN(n7088) );
  NAND2_X1 U8729 ( .A1(n7181), .A2(n7088), .ZN(n7098) );
  INV_X1 U8730 ( .A(n7091), .ZN(n7092) );
  NAND2_X1 U8731 ( .A1(n7093), .A2(n7092), .ZN(n7094) );
  INV_X1 U8732 ( .A(n7182), .ZN(n7097) );
  AOI21_X1 U8733 ( .B1(n7098), .B2(n7095), .A(n7097), .ZN(n7106) );
  INV_X1 U8734 ( .A(n7099), .ZN(n7103) );
  INV_X1 U8735 ( .A(n7100), .ZN(n7101) );
  OAI22_X1 U8736 ( .A1(n9050), .A2(n7101), .B1(n9095), .B2(n7237), .ZN(n7102)
         );
  AOI211_X1 U8737 ( .C1(n9092), .C2(n9109), .A(n7103), .B(n7102), .ZN(n7105)
         );
  NAND2_X1 U8738 ( .A1(n9464), .A2(n9084), .ZN(n7104) );
  OAI211_X1 U8739 ( .C1(n7106), .C2(n9086), .A(n7105), .B(n7104), .ZN(P1_U3222) );
  OAI21_X1 U8740 ( .B1(n8267), .B2(n7107), .A(n7170), .ZN(n7115) );
  OAI22_X1 U8741 ( .A1(n7108), .A2(n8859), .B1(n7261), .B2(n8861), .ZN(n7114)
         );
  AND2_X1 U8742 ( .A1(n7110), .A2(n7109), .ZN(n7112) );
  OAI21_X1 U8743 ( .B1(n7112), .B2(n8374), .A(n7111), .ZN(n8956) );
  NOR2_X1 U8744 ( .A1(n8956), .A2(n7660), .ZN(n7113) );
  AOI211_X1 U8745 ( .C1(n8817), .C2(n7115), .A(n7114), .B(n7113), .ZN(n8955)
         );
  AND2_X1 U8746 ( .A1(n7116), .A2(n8952), .ZN(n7117) );
  NOR2_X1 U8747 ( .A1(n7175), .A2(n7117), .ZN(n8953) );
  INV_X1 U8748 ( .A(n8952), .ZN(n7118) );
  NOR2_X1 U8749 ( .A1(n7118), .A2(n8869), .ZN(n7122) );
  OAI22_X1 U8750 ( .A1(n8826), .A2(n7120), .B1(n7119), .B2(n9742), .ZN(n7121)
         );
  AOI211_X1 U8751 ( .C1(n8953), .C2(n8864), .A(n7122), .B(n7121), .ZN(n7125)
         );
  INV_X1 U8752 ( .A(n8956), .ZN(n7123) );
  NAND2_X1 U8753 ( .A1(n7123), .A2(n7333), .ZN(n7124) );
  OAI211_X1 U8754 ( .C1(n8955), .C2(n9752), .A(n7125), .B(n7124), .ZN(P2_U3283) );
  INV_X1 U8755 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7132) );
  AOI211_X1 U8756 ( .C1(n9772), .C2(n7128), .A(n7127), .B(n7126), .ZN(n7129)
         );
  OAI21_X1 U8757 ( .B1(n9790), .B2(n7130), .A(n7129), .ZN(n7133) );
  NAND2_X1 U8758 ( .A1(n7133), .A2(n9817), .ZN(n7131) );
  OAI21_X1 U8759 ( .B1(n9817), .B2(n7132), .A(n7131), .ZN(P2_U3487) );
  NAND2_X1 U8760 ( .A1(n7133), .A2(n9830), .ZN(n7134) );
  OAI21_X1 U8761 ( .B1(n9830), .B2(n7055), .A(n7134), .ZN(P2_U3532) );
  AND2_X1 U8762 ( .A1(n9464), .A2(n9108), .ZN(n7135) );
  NAND2_X1 U8763 ( .A1(n7138), .A2(n7896), .ZN(n7140) );
  AOI22_X1 U8764 ( .A1(n7804), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5941), .B2(
        n7313), .ZN(n7139) );
  OR2_X1 U8765 ( .A1(n7236), .A2(n7237), .ZN(n7953) );
  NAND2_X1 U8766 ( .A1(n7236), .A2(n7237), .ZN(n7833) );
  NAND2_X1 U8767 ( .A1(n7953), .A2(n7833), .ZN(n8045) );
  XNOR2_X1 U8768 ( .A(n7239), .B(n8045), .ZN(n9551) );
  INV_X1 U8769 ( .A(n7142), .ZN(n7143) );
  NAND2_X1 U8770 ( .A1(n7949), .A2(n7143), .ZN(n7144) );
  AND2_X1 U8771 ( .A1(n7144), .A2(n7950), .ZN(n7954) );
  NAND2_X1 U8772 ( .A1(n7145), .A2(n8045), .ZN(n7146) );
  NAND2_X1 U8773 ( .A1(n4857), .A2(n7146), .ZN(n7147) );
  NAND2_X1 U8774 ( .A1(n7147), .A2(n9355), .ZN(n7156) );
  NAND2_X1 U8775 ( .A1(n7869), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7154) );
  NAND2_X1 U8776 ( .A1(n7822), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7153) );
  INV_X1 U8777 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7148) );
  NAND2_X1 U8778 ( .A1(n7149), .A2(n7148), .ZN(n7150) );
  AND2_X1 U8779 ( .A1(n7242), .A2(n7150), .ZN(n7436) );
  NAND2_X1 U8780 ( .A1(n7346), .A2(n7436), .ZN(n7152) );
  NAND2_X1 U8781 ( .A1(n7244), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7151) );
  NAND4_X1 U8782 ( .A1(n7154), .A2(n7153), .A3(n7152), .A4(n7151), .ZN(n9106)
         );
  AOI22_X1 U8783 ( .A1(n9372), .A2(n9106), .B1(n9380), .B2(n9108), .ZN(n7155)
         );
  NAND2_X1 U8784 ( .A1(n7156), .A2(n7155), .ZN(n7157) );
  AOI21_X1 U8785 ( .B1(n9551), .B2(n7158), .A(n7157), .ZN(n9553) );
  AOI21_X1 U8786 ( .B1(n4506), .B2(n7236), .A(n9696), .ZN(n7161) );
  NAND2_X1 U8787 ( .A1(n7161), .A2(n7251), .ZN(n9549) );
  AOI22_X1 U8788 ( .A1(n9356), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7194), .B2(
        n9343), .ZN(n7163) );
  NAND2_X1 U8789 ( .A1(n7236), .A2(n9183), .ZN(n7162) );
  OAI211_X1 U8790 ( .C1(n9549), .C2(n7256), .A(n7163), .B(n7162), .ZN(n7164)
         );
  AOI21_X1 U8791 ( .B1(n9551), .B2(n7165), .A(n7164), .ZN(n7166) );
  OAI21_X1 U8792 ( .B1(n9553), .B2(n9319), .A(n7166), .ZN(P1_U3278) );
  XNOR2_X1 U8793 ( .A(n7167), .B(n8268), .ZN(n9531) );
  INV_X1 U8794 ( .A(n9531), .ZN(n7180) );
  NAND2_X1 U8795 ( .A1(n7168), .A2(n8817), .ZN(n7173) );
  AOI21_X1 U8796 ( .B1(n7170), .B2(n7169), .A(n8268), .ZN(n7172) );
  AOI22_X1 U8797 ( .A1(n7567), .A2(n8627), .B1(n8629), .B2(n7566), .ZN(n7171)
         );
  OAI21_X1 U8798 ( .B1(n7173), .B2(n7172), .A(n7171), .ZN(n9530) );
  INV_X1 U8799 ( .A(n7174), .ZN(n7266) );
  OAI21_X1 U8800 ( .B1(n9527), .B2(n7175), .A(n7266), .ZN(n9528) );
  OAI22_X1 U8801 ( .A1(n8826), .A2(n8643), .B1(n7210), .B2(n9742), .ZN(n7176)
         );
  AOI21_X1 U8802 ( .B1(n7214), .B2(n8828), .A(n7176), .ZN(n7177) );
  OAI21_X1 U8803 ( .B1(n9528), .B2(n8736), .A(n7177), .ZN(n7178) );
  AOI21_X1 U8804 ( .B1(n9530), .B2(n8826), .A(n7178), .ZN(n7179) );
  OAI21_X1 U8805 ( .B1(n7180), .B2(n8873), .A(n7179), .ZN(P2_U3282) );
  NAND2_X1 U8806 ( .A1(n7236), .A2(n5930), .ZN(n7184) );
  NAND2_X1 U8807 ( .A1(n9107), .A2(n8508), .ZN(n7183) );
  NAND2_X1 U8808 ( .A1(n7184), .A2(n7183), .ZN(n7185) );
  XNOR2_X1 U8809 ( .A(n7185), .B(n8482), .ZN(n7190) );
  INV_X1 U8810 ( .A(n7190), .ZN(n7188) );
  AND2_X1 U8811 ( .A1(n9002), .A2(n9107), .ZN(n7186) );
  AOI21_X1 U8812 ( .B1(n7236), .B2(n8508), .A(n7186), .ZN(n7189) );
  INV_X1 U8813 ( .A(n7189), .ZN(n7187) );
  NAND2_X1 U8814 ( .A1(n7188), .A2(n7187), .ZN(n7428) );
  INV_X1 U8815 ( .A(n7428), .ZN(n7191) );
  AND2_X1 U8816 ( .A1(n7190), .A2(n7189), .ZN(n7422) );
  NOR2_X1 U8817 ( .A1(n7191), .A2(n7422), .ZN(n7192) );
  XNOR2_X1 U8818 ( .A(n7421), .B(n7192), .ZN(n7193) );
  NAND2_X1 U8819 ( .A1(n7193), .A2(n9088), .ZN(n7199) );
  INV_X1 U8820 ( .A(n7194), .ZN(n7195) );
  OAI22_X1 U8821 ( .A1(n9050), .A2(n7195), .B1(n9095), .B2(n7831), .ZN(n7196)
         );
  AOI211_X1 U8822 ( .C1(n9092), .C2(n9108), .A(n7197), .B(n7196), .ZN(n7198)
         );
  OAI211_X1 U8823 ( .C1(n7159), .C2(n9102), .A(n7199), .B(n7198), .ZN(P1_U3232) );
  XNOR2_X1 U8824 ( .A(n7214), .B(n8173), .ZN(n7200) );
  OR2_X1 U8825 ( .A1(n7261), .A2(n8187), .ZN(n7201) );
  NAND2_X1 U8826 ( .A1(n7200), .A2(n7201), .ZN(n7375) );
  INV_X1 U8827 ( .A(n7200), .ZN(n7203) );
  INV_X1 U8828 ( .A(n7201), .ZN(n7202) );
  NAND2_X1 U8829 ( .A1(n7203), .A2(n7202), .ZN(n7204) );
  NAND2_X1 U8830 ( .A1(n7375), .A2(n7204), .ZN(n7372) );
  NAND2_X1 U8831 ( .A1(n7385), .A2(n7376), .ZN(n7208) );
  INV_X1 U8832 ( .A(n7205), .ZN(n7207) );
  NAND2_X1 U8833 ( .A1(n7207), .A2(n7206), .ZN(n7370) );
  NAND2_X1 U8834 ( .A1(n7208), .A2(n7370), .ZN(n7209) );
  AOI21_X1 U8835 ( .B1(n7372), .B2(n7209), .A(n4366), .ZN(n7216) );
  NAND2_X1 U8836 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7414) );
  OAI21_X1 U8837 ( .B1(n8606), .B2(n7210), .A(n7414), .ZN(n7213) );
  OAI22_X1 U8838 ( .A1(n8382), .A2(n8608), .B1(n8607), .B2(n7211), .ZN(n7212)
         );
  AOI211_X1 U8839 ( .C1(n7214), .C2(n8583), .A(n7213), .B(n7212), .ZN(n7215)
         );
  OAI21_X1 U8840 ( .B1(n7216), .B2(n8587), .A(n7215), .ZN(P2_U3217) );
  NAND2_X1 U8841 ( .A1(n7218), .A2(n7217), .ZN(n7220) );
  AOI22_X1 U8842 ( .A1(n7409), .A2(n7120), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7402), .ZN(n7219) );
  NOR2_X1 U8843 ( .A1(n7220), .A2(n7219), .ZN(n7401) );
  AOI21_X1 U8844 ( .B1(n7220), .B2(n7219), .A(n7401), .ZN(n7221) );
  OR2_X1 U8845 ( .A1(n7221), .A2(n9730), .ZN(n7232) );
  OR2_X1 U8846 ( .A1(n7222), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7223) );
  NAND2_X1 U8847 ( .A1(n7224), .A2(n7223), .ZN(n7226) );
  AOI22_X1 U8848 ( .A1(n7409), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5254), .B2(
        n7402), .ZN(n7225) );
  NAND2_X1 U8849 ( .A1(n7225), .A2(n7226), .ZN(n7408) );
  OAI21_X1 U8850 ( .B1(n7226), .B2(n7225), .A(n7408), .ZN(n7230) );
  INV_X1 U8851 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7228) );
  OAI22_X1 U8852 ( .A1(n8724), .A2(n7228), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7227), .ZN(n7229) );
  AOI21_X1 U8853 ( .B1(n9727), .B2(n7230), .A(n7229), .ZN(n7231) );
  OAI211_X1 U8854 ( .C1(n9731), .C2(n7402), .A(n7232), .B(n7231), .ZN(P2_U3258) );
  NAND2_X1 U8855 ( .A1(n7233), .A2(n7896), .ZN(n7235) );
  AOI22_X1 U8856 ( .A1(n7804), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5941), .B2(
        n9659), .ZN(n7234) );
  XNOR2_X1 U8857 ( .A(n7832), .B(n7831), .ZN(n8046) );
  NOR2_X1 U8858 ( .A1(n7236), .A2(n9107), .ZN(n7238) );
  OAI22_X2 U8859 ( .A1(n7239), .A2(n7238), .B1(n7237), .B2(n7159), .ZN(n7337)
         );
  XOR2_X1 U8860 ( .A(n8046), .B(n7337), .Z(n9547) );
  INV_X1 U8861 ( .A(n9547), .ZN(n7259) );
  INV_X1 U8862 ( .A(n8046), .ZN(n7240) );
  XNOR2_X1 U8863 ( .A(n7342), .B(n7240), .ZN(n7241) );
  NAND2_X1 U8864 ( .A1(n7241), .A2(n9355), .ZN(n7250) );
  INV_X1 U8865 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U8866 ( .A1(n7242), .A2(n7492), .ZN(n7243) );
  AND2_X1 U8867 ( .A1(n7344), .A2(n7243), .ZN(n7355) );
  NAND2_X1 U8868 ( .A1(n7346), .A2(n7355), .ZN(n7248) );
  NAND2_X1 U8869 ( .A1(n7869), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7247) );
  NAND2_X1 U8870 ( .A1(n7822), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7246) );
  NAND2_X1 U8871 ( .A1(n7244), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7245) );
  NAND4_X1 U8872 ( .A1(n7248), .A2(n7247), .A3(n7246), .A4(n7245), .ZN(n9105)
         );
  AOI22_X1 U8873 ( .A1(n9380), .A2(n9107), .B1(n9372), .B2(n9105), .ZN(n7249)
         );
  NAND2_X1 U8874 ( .A1(n7250), .A2(n7249), .ZN(n9546) );
  INV_X1 U8875 ( .A(n7251), .ZN(n7253) );
  INV_X1 U8876 ( .A(n7357), .ZN(n7252) );
  OAI211_X1 U8877 ( .C1(n9544), .C2(n7253), .A(n7252), .B(n9437), .ZN(n9543)
         );
  AOI22_X1 U8878 ( .A1(n9356), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7436), .B2(
        n9343), .ZN(n7255) );
  NAND2_X1 U8879 ( .A1(n7832), .A2(n9183), .ZN(n7254) );
  OAI211_X1 U8880 ( .C1(n9543), .C2(n7256), .A(n7255), .B(n7254), .ZN(n7257)
         );
  AOI21_X1 U8881 ( .B1(n9546), .B2(n9367), .A(n7257), .ZN(n7258) );
  OAI21_X1 U8882 ( .B1(n7259), .B2(n9383), .A(n7258), .ZN(P1_U3277) );
  XNOR2_X1 U8883 ( .A(n7260), .B(n8376), .ZN(n7262) );
  OAI22_X1 U8884 ( .A1(n7509), .A2(n8861), .B1(n7261), .B2(n8859), .ZN(n7691)
         );
  AOI21_X1 U8885 ( .B1(n7262), .B2(n8817), .A(n7691), .ZN(n8950) );
  OAI21_X1 U8886 ( .B1(n7264), .B2(n8376), .A(n7263), .ZN(n8946) );
  INV_X1 U8887 ( .A(n7328), .ZN(n7265) );
  AOI21_X1 U8888 ( .B1(n8947), .B2(n7266), .A(n7265), .ZN(n8948) );
  NAND2_X1 U8889 ( .A1(n8948), .A2(n8864), .ZN(n7269) );
  INV_X1 U8890 ( .A(n7693), .ZN(n7267) );
  INV_X1 U8891 ( .A(n9742), .ZN(n8865) );
  AOI22_X1 U8892 ( .A1(n9752), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7267), .B2(
        n8865), .ZN(n7268) );
  OAI211_X1 U8893 ( .C1(n8383), .C2(n8869), .A(n7269), .B(n7268), .ZN(n7270)
         );
  AOI21_X1 U8894 ( .B1(n8946), .B2(n8823), .A(n7270), .ZN(n7271) );
  OAI21_X1 U8895 ( .B1(n9752), .B2(n8950), .A(n7271), .ZN(P2_U3281) );
  INV_X1 U8896 ( .A(n7756), .ZN(n7274) );
  OAI222_X1 U8897 ( .A1(n9495), .A2(n7757), .B1(n9493), .B2(n7274), .C1(n7272), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U8898 ( .A1(n8979), .A2(n7275), .B1(n8233), .B2(n7274), .C1(
        P2_U3152), .C2(n7273), .ZN(P2_U3333) );
  INV_X1 U8899 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U8900 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7276) );
  AOI21_X1 U8901 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7276), .ZN(n9838) );
  NOR2_X1 U8902 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7277) );
  AOI21_X1 U8903 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7277), .ZN(n9841) );
  NOR2_X1 U8904 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7278) );
  AOI21_X1 U8905 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7278), .ZN(n9844) );
  NOR2_X1 U8906 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7279) );
  AOI21_X1 U8907 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7279), .ZN(n9847) );
  NOR2_X1 U8908 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7280) );
  AOI21_X1 U8909 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7280), .ZN(n9850) );
  NOR2_X1 U8910 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7286) );
  XOR2_X1 U8911 ( .A(n9613), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10067) );
  NAND2_X1 U8912 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7284) );
  XOR2_X1 U8913 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10065) );
  NAND2_X1 U8914 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7282) );
  INV_X1 U8915 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9596) );
  XNOR2_X1 U8916 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9596), .ZN(n10063) );
  AOI21_X1 U8917 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9831) );
  INV_X1 U8918 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9835) );
  NAND3_X1 U8919 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9833) );
  OAI21_X1 U8920 ( .B1(n9831), .B2(n9835), .A(n9833), .ZN(n10062) );
  NAND2_X1 U8921 ( .A1(n10063), .A2(n10062), .ZN(n7281) );
  NAND2_X1 U8922 ( .A1(n7282), .A2(n7281), .ZN(n10064) );
  NAND2_X1 U8923 ( .A1(n10065), .A2(n10064), .ZN(n7283) );
  NAND2_X1 U8924 ( .A1(n7284), .A2(n7283), .ZN(n10066) );
  NOR2_X1 U8925 ( .A1(n10067), .A2(n10066), .ZN(n7285) );
  NOR2_X1 U8926 ( .A1(n7286), .A2(n7285), .ZN(n7287) );
  NOR2_X1 U8927 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7287), .ZN(n10051) );
  AND2_X1 U8928 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7287), .ZN(n10050) );
  NOR2_X1 U8929 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10050), .ZN(n7288) );
  NOR2_X1 U8930 ( .A1(n10051), .A2(n7288), .ZN(n7289) );
  NAND2_X1 U8931 ( .A1(n7289), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7291) );
  XOR2_X1 U8932 ( .A(n7289), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10049) );
  NAND2_X1 U8933 ( .A1(n10049), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7290) );
  NAND2_X1 U8934 ( .A1(n7291), .A2(n7290), .ZN(n7292) );
  NAND2_X1 U8935 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7292), .ZN(n7294) );
  XOR2_X1 U8936 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7292), .Z(n10061) );
  NAND2_X1 U8937 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10061), .ZN(n7293) );
  NAND2_X1 U8938 ( .A1(n7294), .A2(n7293), .ZN(n7295) );
  NAND2_X1 U8939 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7295), .ZN(n7297) );
  INV_X1 U8940 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9631) );
  XNOR2_X1 U8941 ( .A(n9631), .B(n7295), .ZN(n10060) );
  NAND2_X1 U8942 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10060), .ZN(n7296) );
  NAND2_X1 U8943 ( .A1(n7297), .A2(n7296), .ZN(n7298) );
  AND2_X1 U8944 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7298), .ZN(n7299) );
  INV_X1 U8945 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10059) );
  XNOR2_X1 U8946 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7298), .ZN(n10058) );
  NOR2_X1 U8947 ( .A1(n10059), .A2(n10058), .ZN(n10057) );
  NAND2_X1 U8948 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7300) );
  OAI21_X1 U8949 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7300), .ZN(n9858) );
  NAND2_X1 U8950 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7301) );
  OAI21_X1 U8951 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7301), .ZN(n9855) );
  NOR2_X1 U8952 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7302) );
  AOI21_X1 U8953 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7302), .ZN(n9852) );
  NAND2_X1 U8954 ( .A1(n9853), .A2(n9852), .ZN(n9851) );
  NAND2_X1 U8955 ( .A1(n9850), .A2(n9849), .ZN(n9848) );
  OAI21_X1 U8956 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9848), .ZN(n9846) );
  NAND2_X1 U8957 ( .A1(n9847), .A2(n9846), .ZN(n9845) );
  OAI21_X1 U8958 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9845), .ZN(n9843) );
  NAND2_X1 U8959 ( .A1(n9844), .A2(n9843), .ZN(n9842) );
  OAI21_X1 U8960 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9842), .ZN(n9840) );
  NAND2_X1 U8961 ( .A1(n9841), .A2(n9840), .ZN(n9839) );
  OAI21_X1 U8962 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9839), .ZN(n9837) );
  NAND2_X1 U8963 ( .A1(n9838), .A2(n9837), .ZN(n9836) );
  OAI21_X1 U8964 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9836), .ZN(n10054) );
  NOR2_X1 U8965 ( .A1(n10055), .A2(n10054), .ZN(n7303) );
  NAND2_X1 U8966 ( .A1(n10055), .A2(n10054), .ZN(n10053) );
  OAI21_X1 U8967 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7303), .A(n10053), .ZN(
        n7305) );
  XNOR2_X1 U8968 ( .A(n4903), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7304) );
  XNOR2_X1 U8969 ( .A(n7305), .B(n7304), .ZN(ADD_1071_U4) );
  NAND2_X1 U8970 ( .A1(n7307), .A2(n7311), .ZN(n7308) );
  INV_X1 U8971 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U8972 ( .A1(n7308), .A2(n9660), .ZN(n9134) );
  XNOR2_X1 U8973 ( .A(n9134), .B(n9141), .ZN(n7309) );
  INV_X1 U8974 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7356) );
  NOR2_X1 U8975 ( .A1(n7356), .A2(n7309), .ZN(n9135) );
  AOI211_X1 U8976 ( .C1(n7309), .C2(n7356), .A(n9135), .B(n9637), .ZN(n7310)
         );
  INV_X1 U8977 ( .A(n7310), .ZN(n7318) );
  AND2_X1 U8978 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3084), .ZN(n7316) );
  INV_X1 U8979 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9548) );
  AOI22_X1 U8980 ( .A1(n9659), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n9548), .B2(
        n7311), .ZN(n9665) );
  OAI21_X1 U8981 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7313), .A(n7312), .ZN(
        n9664) );
  NAND2_X1 U8982 ( .A1(n9665), .A2(n9664), .ZN(n9663) );
  INV_X1 U8983 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9542) );
  NOR2_X1 U8984 ( .A1(n9542), .A2(n7314), .ZN(n9142) );
  AOI211_X1 U8985 ( .C1(n7314), .C2(n9542), .A(n9142), .B(n9579), .ZN(n7315)
         );
  AOI211_X1 U8986 ( .C1(P1_ADDR_REG_15__SCAN_IN), .C2(n9685), .A(n7316), .B(
        n7315), .ZN(n7317) );
  OAI211_X1 U8987 ( .C1(n9592), .C2(n9141), .A(n7318), .B(n7317), .ZN(P1_U3256) );
  NAND2_X1 U8988 ( .A1(n7319), .A2(n7320), .ZN(n7321) );
  NAND2_X1 U8989 ( .A1(n7321), .A2(n8385), .ZN(n7508) );
  OAI21_X1 U8990 ( .B1(n8385), .B2(n7321), .A(n7508), .ZN(n7326) );
  OAI22_X1 U8991 ( .A1(n7565), .A2(n8861), .B1(n8382), .B2(n8859), .ZN(n7441)
         );
  NAND2_X1 U8992 ( .A1(n7322), .A2(n8385), .ZN(n7323) );
  NAND2_X1 U8993 ( .A1(n7324), .A2(n7323), .ZN(n8945) );
  NOR2_X1 U8994 ( .A1(n8945), .A2(n7660), .ZN(n7325) );
  AOI211_X1 U8995 ( .C1(n8817), .C2(n7326), .A(n7441), .B(n7325), .ZN(n8944)
         );
  INV_X1 U8996 ( .A(n7504), .ZN(n7327) );
  AOI21_X1 U8997 ( .B1(n8941), .B2(n7328), .A(n7327), .ZN(n8942) );
  NOR2_X1 U8998 ( .A1(n7329), .A2(n8869), .ZN(n7332) );
  OAI22_X1 U8999 ( .A1(n8826), .A2(n7330), .B1(n7443), .B2(n9742), .ZN(n7331)
         );
  AOI211_X1 U9000 ( .C1(n8942), .C2(n8864), .A(n7332), .B(n7331), .ZN(n7336)
         );
  INV_X1 U9001 ( .A(n8945), .ZN(n7334) );
  NAND2_X1 U9002 ( .A1(n7334), .A2(n7333), .ZN(n7335) );
  OAI211_X1 U9003 ( .C1(n8944), .C2(n9752), .A(n7336), .B(n7335), .ZN(P2_U3280) );
  NAND2_X1 U9004 ( .A1(n7338), .A2(n7896), .ZN(n7341) );
  INV_X1 U9005 ( .A(n9141), .ZN(n7339) );
  AOI22_X1 U9006 ( .A1(n7804), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5941), .B2(
        n7339), .ZN(n7340) );
  OR2_X1 U9007 ( .A1(n7496), .A2(n7467), .ZN(n7967) );
  NAND2_X1 U9008 ( .A1(n7496), .A2(n7467), .ZN(n7966) );
  NAND2_X1 U9009 ( .A1(n7967), .A2(n7966), .ZN(n8047) );
  XNOR2_X1 U9010 ( .A(n7454), .B(n8047), .ZN(n9536) );
  XNOR2_X1 U9011 ( .A(n7465), .B(n8047), .ZN(n7352) );
  NAND2_X1 U9012 ( .A1(n7869), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7350) );
  NAND2_X1 U9013 ( .A1(n7244), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7349) );
  NAND2_X1 U9014 ( .A1(n7344), .A2(n7343), .ZN(n7345) );
  AND2_X1 U9015 ( .A1(n7459), .A2(n7345), .ZN(n7533) );
  NAND2_X1 U9016 ( .A1(n7346), .A2(n7533), .ZN(n7348) );
  NAND2_X1 U9017 ( .A1(n7822), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7347) );
  NAND4_X1 U9018 ( .A1(n7350), .A2(n7349), .A3(n7348), .A4(n7347), .ZN(n9379)
         );
  OAI22_X1 U9019 ( .A1(n7831), .A2(n9331), .B1(n7610), .B2(n9329), .ZN(n7351)
         );
  AOI21_X1 U9020 ( .B1(n7352), .B2(n9355), .A(n7351), .ZN(n7353) );
  OAI21_X1 U9021 ( .B1(n9536), .B2(n7354), .A(n7353), .ZN(n9539) );
  NAND2_X1 U9022 ( .A1(n9539), .A2(n9367), .ZN(n7362) );
  INV_X1 U9023 ( .A(n7355), .ZN(n7493) );
  OAI22_X1 U9024 ( .A1(n9367), .A2(n7356), .B1(n7493), .B2(n9365), .ZN(n7360)
         );
  NAND2_X1 U9025 ( .A1(n7357), .A2(n9537), .ZN(n7469) );
  OR2_X1 U9026 ( .A1(n7357), .A2(n9537), .ZN(n7358) );
  NAND2_X1 U9027 ( .A1(n7469), .A2(n7358), .ZN(n9538) );
  NOR2_X1 U9028 ( .A1(n9538), .A2(n9186), .ZN(n7359) );
  AOI211_X1 U9029 ( .C1(n9183), .C2(n7496), .A(n7360), .B(n7359), .ZN(n7361)
         );
  OAI211_X1 U9030 ( .C1(n9536), .C2(n7363), .A(n7362), .B(n7361), .ZN(P1_U3276) );
  INV_X1 U9031 ( .A(n7743), .ZN(n7399) );
  OAI222_X1 U9032 ( .A1(P2_U3152), .A2(n7365), .B1(n8980), .B2(n7399), .C1(
        n7364), .C2(n8979), .ZN(P2_U3332) );
  INV_X1 U9033 ( .A(n7372), .ZN(n7368) );
  AND2_X1 U9034 ( .A1(n7370), .A2(n7366), .ZN(n7367) );
  AND2_X1 U9035 ( .A1(n7368), .A2(n7367), .ZN(n7369) );
  INV_X1 U9036 ( .A(n7375), .ZN(n7374) );
  INV_X1 U9037 ( .A(n7370), .ZN(n7371) );
  OR2_X1 U9038 ( .A1(n7374), .A2(n7373), .ZN(n7380) );
  AND2_X1 U9039 ( .A1(n7376), .A2(n7375), .ZN(n7383) );
  INV_X1 U9040 ( .A(n7383), .ZN(n7377) );
  XNOR2_X1 U9041 ( .A(n8947), .B(n8173), .ZN(n7381) );
  NAND2_X1 U9042 ( .A1(n7379), .A2(n7381), .ZN(n7445) );
  OR2_X1 U9043 ( .A1(n7381), .A2(n7380), .ZN(n7387) );
  INV_X1 U9044 ( .A(n7381), .ZN(n7382) );
  AND2_X1 U9045 ( .A1(n7383), .A2(n7382), .ZN(n7384) );
  XNOR2_X1 U9046 ( .A(n8941), .B(n8173), .ZN(n7391) );
  NOR2_X1 U9047 ( .A1(n7509), .A2(n8187), .ZN(n7389) );
  XNOR2_X1 U9048 ( .A(n7391), .B(n7389), .ZN(n7444) );
  NAND2_X1 U9049 ( .A1(n7388), .A2(n7444), .ZN(n7448) );
  INV_X1 U9050 ( .A(n7389), .ZN(n7390) );
  NAND2_X1 U9051 ( .A1(n7391), .A2(n7390), .ZN(n7392) );
  XNOR2_X1 U9052 ( .A(n5318), .B(n8195), .ZN(n7474) );
  NOR2_X1 U9053 ( .A1(n7565), .A2(n8187), .ZN(n7475) );
  XNOR2_X1 U9054 ( .A(n7474), .B(n7475), .ZN(n7476) );
  XNOR2_X1 U9055 ( .A(n7477), .B(n7476), .ZN(n7398) );
  INV_X1 U9056 ( .A(n7393), .ZN(n7503) );
  OAI22_X1 U9057 ( .A1(n8606), .A2(n7503), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5028), .ZN(n7396) );
  OAI22_X1 U9058 ( .A1(n7509), .A2(n8607), .B1(n8608), .B2(n7394), .ZN(n7395)
         );
  AOI211_X1 U9059 ( .C1(n5318), .C2(n8583), .A(n7396), .B(n7395), .ZN(n7397)
         );
  OAI21_X1 U9060 ( .B1(n7398), .B2(n8587), .A(n7397), .ZN(P2_U3230) );
  OAI222_X1 U9061 ( .A1(n9495), .A2(n7744), .B1(P1_U3084), .B2(n7400), .C1(
        n9493), .C2(n7399), .ZN(P1_U3327) );
  AOI21_X1 U9062 ( .B1(n7402), .B2(n7120), .A(n7401), .ZN(n7405) );
  NOR2_X1 U9063 ( .A1(n7407), .A2(n8643), .ZN(n7403) );
  AOI21_X1 U9064 ( .B1(n7407), .B2(n8643), .A(n7403), .ZN(n7404) );
  NOR2_X1 U9065 ( .A1(n7405), .A2(n7404), .ZN(n8642) );
  AOI21_X1 U9066 ( .B1(n7405), .B2(n7404), .A(n8642), .ZN(n7420) );
  NAND2_X1 U9067 ( .A1(n7407), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7406) );
  OAI21_X1 U9068 ( .B1(n7407), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7406), .ZN(
        n7412) );
  OAI21_X1 U9069 ( .B1(n7409), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7408), .ZN(
        n7410) );
  NAND2_X1 U9070 ( .A1(n7412), .A2(n7411), .ZN(n7413) );
  NAND2_X1 U9071 ( .A1(n8648), .A2(n7413), .ZN(n7417) );
  INV_X1 U9072 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7415) );
  OAI21_X1 U9073 ( .B1(n8724), .B2(n7415), .A(n7414), .ZN(n7416) );
  AOI21_X1 U9074 ( .B1(n9727), .B2(n7417), .A(n7416), .ZN(n7419) );
  OR2_X1 U9075 ( .A1(n9731), .A2(n8646), .ZN(n7418) );
  OAI211_X1 U9076 ( .C1(n7420), .C2(n9730), .A(n7419), .B(n7418), .ZN(P2_U3259) );
  NAND2_X1 U9077 ( .A1(n7431), .A2(n7428), .ZN(n7427) );
  NAND2_X1 U9078 ( .A1(n7832), .A2(n5930), .ZN(n7424) );
  NAND2_X1 U9079 ( .A1(n9106), .A2(n8508), .ZN(n7423) );
  NAND2_X1 U9080 ( .A1(n7424), .A2(n7423), .ZN(n7425) );
  XNOR2_X1 U9081 ( .A(n7425), .B(n8482), .ZN(n7429) );
  INV_X1 U9082 ( .A(n7429), .ZN(n7426) );
  AND2_X1 U9083 ( .A1(n7429), .A2(n7428), .ZN(n7430) );
  NAND2_X1 U9084 ( .A1(n7431), .A2(n7430), .ZN(n7485) );
  NAND2_X1 U9085 ( .A1(n7486), .A2(n7485), .ZN(n7434) );
  NAND2_X1 U9086 ( .A1(n7832), .A2(n8508), .ZN(n7433) );
  NAND2_X1 U9087 ( .A1(n9002), .A2(n9106), .ZN(n7432) );
  NAND2_X1 U9088 ( .A1(n7433), .A2(n7432), .ZN(n7484) );
  XNOR2_X1 U9089 ( .A(n7434), .B(n7484), .ZN(n7435) );
  NAND2_X1 U9090 ( .A1(n7435), .A2(n9088), .ZN(n7440) );
  AND2_X1 U9091 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9658) );
  INV_X1 U9092 ( .A(n7436), .ZN(n7437) );
  OAI22_X1 U9093 ( .A1(n9050), .A2(n7437), .B1(n9095), .B2(n7467), .ZN(n7438)
         );
  AOI211_X1 U9094 ( .C1(n9092), .C2(n9107), .A(n9658), .B(n7438), .ZN(n7439)
         );
  OAI211_X1 U9095 ( .C1(n9544), .C2(n9102), .A(n7440), .B(n7439), .ZN(P1_U3213) );
  AOI22_X1 U9096 ( .A1(n8580), .A2(n7441), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n7442) );
  OAI21_X1 U9097 ( .B1(n7443), .B2(n8606), .A(n7442), .ZN(n7450) );
  INV_X1 U9098 ( .A(n7444), .ZN(n7446) );
  NAND3_X1 U9099 ( .A1(n7698), .A2(n7446), .A3(n7445), .ZN(n7447) );
  AOI21_X1 U9100 ( .B1(n7448), .B2(n7447), .A(n8587), .ZN(n7449) );
  AOI211_X1 U9101 ( .C1(n8941), .C2(n8583), .A(n7450), .B(n7449), .ZN(n7451)
         );
  INV_X1 U9102 ( .A(n7451), .ZN(P2_U3228) );
  INV_X1 U9103 ( .A(n7733), .ZN(n7453) );
  OAI222_X1 U9104 ( .A1(n8979), .A2(n7452), .B1(n8233), .B2(n7453), .C1(n5509), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  OAI222_X1 U9105 ( .A1(n9495), .A2(n7734), .B1(P1_U3084), .B2(n8117), .C1(
        n7453), .C2(n9493), .ZN(P1_U3326) );
  NAND2_X1 U9106 ( .A1(n7455), .A2(n7896), .ZN(n7457) );
  AOI22_X1 U9107 ( .A1(n7804), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5941), .B2(
        n9158), .ZN(n7456) );
  NAND2_X1 U9108 ( .A1(n9459), .A2(n7610), .ZN(n8137) );
  NAND2_X1 U9109 ( .A1(n8135), .A2(n8137), .ZN(n8122) );
  XNOR2_X1 U9110 ( .A(n8123), .B(n8122), .ZN(n9461) );
  NAND2_X1 U9111 ( .A1(n4305), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7464) );
  INV_X1 U9112 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7458) );
  NAND2_X1 U9113 ( .A1(n7459), .A2(n7458), .ZN(n7460) );
  AND2_X1 U9114 ( .A1(n7808), .A2(n7460), .ZN(n7609) );
  NAND2_X1 U9115 ( .A1(n7346), .A2(n7609), .ZN(n7463) );
  NAND2_X1 U9116 ( .A1(n7244), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7462) );
  NAND2_X1 U9117 ( .A1(n7822), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7461) );
  NAND4_X1 U9118 ( .A1(n7464), .A2(n7463), .A3(n7462), .A4(n7461), .ZN(n9353)
         );
  XNOR2_X1 U9119 ( .A(n8136), .B(n8122), .ZN(n7466) );
  OAI222_X1 U9120 ( .A1(n9331), .A2(n7467), .B1(n9329), .B2(n8124), .C1(n7466), 
        .C2(n9374), .ZN(n9457) );
  INV_X1 U9121 ( .A(n9459), .ZN(n7539) );
  INV_X1 U9122 ( .A(n9363), .ZN(n7468) );
  AOI211_X1 U9123 ( .C1(n9459), .C2(n7469), .A(n9696), .B(n7468), .ZN(n9458)
         );
  NAND2_X1 U9124 ( .A1(n9458), .A2(n9370), .ZN(n7471) );
  AOI22_X1 U9125 ( .A1(n9356), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7533), .B2(
        n9343), .ZN(n7470) );
  OAI211_X1 U9126 ( .C1(n7539), .C2(n9364), .A(n7471), .B(n7470), .ZN(n7472)
         );
  AOI21_X1 U9127 ( .B1(n9457), .B2(n9367), .A(n7472), .ZN(n7473) );
  OAI21_X1 U9128 ( .B1(n9461), .B2(n9383), .A(n7473), .ZN(P1_U3275) );
  XNOR2_X1 U9129 ( .A(n7563), .B(n8173), .ZN(n7576) );
  NAND2_X1 U9130 ( .A1(n8624), .A2(n8250), .ZN(n7574) );
  XNOR2_X1 U9131 ( .A(n7576), .B(n7574), .ZN(n7572) );
  XNOR2_X1 U9132 ( .A(n7573), .B(n7572), .ZN(n7481) );
  NAND2_X1 U9133 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8702) );
  OAI21_X1 U9134 ( .B1(n8606), .B2(n7560), .A(n8702), .ZN(n7479) );
  OAI22_X1 U9135 ( .A1(n7565), .A2(n8607), .B1(n8608), .B2(n7633), .ZN(n7478)
         );
  AOI211_X1 U9136 ( .C1(n8932), .C2(n8583), .A(n7479), .B(n7478), .ZN(n7480)
         );
  OAI21_X1 U9137 ( .B1(n7481), .B2(n8587), .A(n7480), .ZN(P2_U3240) );
  NAND2_X1 U9138 ( .A1(n7496), .A2(n8508), .ZN(n7483) );
  NAND2_X1 U9139 ( .A1(n9002), .A2(n9105), .ZN(n7482) );
  NAND2_X1 U9140 ( .A1(n7483), .A2(n7482), .ZN(n7518) );
  NAND2_X1 U9141 ( .A1(n7496), .A2(n5930), .ZN(n7488) );
  NAND2_X1 U9142 ( .A1(n9105), .A2(n8508), .ZN(n7487) );
  NAND2_X1 U9143 ( .A1(n7488), .A2(n7487), .ZN(n7489) );
  XNOR2_X1 U9144 ( .A(n7489), .B(n6095), .ZN(n7490) );
  NAND2_X1 U9145 ( .A1(n7519), .A2(n7517), .ZN(n7491) );
  XOR2_X1 U9146 ( .A(n7518), .B(n7491), .Z(n7498) );
  OAI22_X1 U9147 ( .A1(n9051), .A2(n7831), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7492), .ZN(n7495) );
  OAI22_X1 U9148 ( .A1(n9050), .A2(n7493), .B1(n9095), .B2(n7610), .ZN(n7494)
         );
  AOI211_X1 U9149 ( .C1(n7496), .C2(n9084), .A(n7495), .B(n7494), .ZN(n7497)
         );
  OAI21_X1 U9150 ( .B1(n7498), .B2(n9086), .A(n7497), .ZN(P1_U3239) );
  INV_X1 U9151 ( .A(n7897), .ZN(n7638) );
  OAI222_X1 U9152 ( .A1(n7500), .A2(P2_U3152), .B1(n8233), .B2(n7638), .C1(
        n7499), .C2(n8979), .ZN(P2_U3329) );
  AOI21_X1 U9153 ( .B1(n8390), .B2(n7502), .A(n7501), .ZN(n8940) );
  INV_X1 U9154 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8677) );
  OAI22_X1 U9155 ( .A1(n8826), .A2(n8677), .B1(n7503), .B2(n9742), .ZN(n7515)
         );
  AOI211_X1 U9156 ( .C1(n5318), .C2(n7504), .A(n9810), .B(n7557), .ZN(n8938)
         );
  AND2_X1 U9157 ( .A1(n7506), .A2(n7505), .ZN(n7507) );
  NAND2_X1 U9158 ( .A1(n7507), .A2(n8817), .ZN(n7512) );
  AOI21_X1 U9159 ( .B1(n7508), .B2(n8387), .A(n8390), .ZN(n7511) );
  INV_X1 U9160 ( .A(n7509), .ZN(n8626) );
  AOI22_X1 U9161 ( .A1(n8626), .A2(n7566), .B1(n7567), .B2(n8624), .ZN(n7510)
         );
  OAI21_X1 U9162 ( .B1(n7512), .B2(n7511), .A(n7510), .ZN(n8937) );
  AOI21_X1 U9163 ( .B1(n8938), .B2(n9744), .A(n8937), .ZN(n7513) );
  NOR2_X1 U9164 ( .A1(n7513), .A2(n9752), .ZN(n7514) );
  AOI211_X1 U9165 ( .C1(n8828), .C2(n5318), .A(n7515), .B(n7514), .ZN(n7516)
         );
  OAI21_X1 U9166 ( .B1(n8940), .B2(n8873), .A(n7516), .ZN(P2_U3279) );
  INV_X1 U9167 ( .A(n7881), .ZN(n8232) );
  OAI222_X1 U9168 ( .A1(n9495), .A2(n7882), .B1(P1_U3084), .B2(n5736), .C1(
        n8232), .C2(n9493), .ZN(P1_U3325) );
  NAND2_X1 U9169 ( .A1(n9459), .A2(n5930), .ZN(n7521) );
  NAND2_X1 U9170 ( .A1(n9379), .A2(n8508), .ZN(n7520) );
  NAND2_X1 U9171 ( .A1(n7521), .A2(n7520), .ZN(n7522) );
  XNOR2_X1 U9172 ( .A(n7522), .B(n6095), .ZN(n7525) );
  NAND2_X1 U9173 ( .A1(n9459), .A2(n8508), .ZN(n7524) );
  NAND2_X1 U9174 ( .A1(n9002), .A2(n9379), .ZN(n7523) );
  NAND2_X1 U9175 ( .A1(n7524), .A2(n7523), .ZN(n7526) );
  NAND2_X1 U9176 ( .A1(n7525), .A2(n7526), .ZN(n7530) );
  INV_X1 U9177 ( .A(n7525), .ZN(n7528) );
  INV_X1 U9178 ( .A(n7526), .ZN(n7527) );
  NAND2_X1 U9179 ( .A1(n7528), .A2(n7527), .ZN(n7600) );
  NOR2_X1 U9180 ( .A1(n7601), .A2(n4821), .ZN(n7532) );
  AOI21_X1 U9181 ( .B1(n7530), .B2(n7600), .A(n7529), .ZN(n7531) );
  OAI21_X1 U9182 ( .B1(n7532), .B2(n7531), .A(n9088), .ZN(n7538) );
  NAND2_X1 U9183 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9147) );
  INV_X1 U9184 ( .A(n9147), .ZN(n7536) );
  INV_X1 U9185 ( .A(n7533), .ZN(n7534) );
  OAI22_X1 U9186 ( .A1(n9050), .A2(n7534), .B1(n9095), .B2(n8124), .ZN(n7535)
         );
  AOI211_X1 U9187 ( .C1(n9092), .C2(n9105), .A(n7536), .B(n7535), .ZN(n7537)
         );
  OAI211_X1 U9188 ( .C1(n7539), .C2(n9102), .A(n7538), .B(n7537), .ZN(P1_U3224) );
  XNOR2_X1 U9189 ( .A(n7540), .B(n8273), .ZN(n8925) );
  INV_X1 U9190 ( .A(n8925), .ZN(n7554) );
  AOI21_X1 U9191 ( .B1(n7558), .B2(n8927), .A(n9810), .ZN(n7541) );
  NAND2_X1 U9192 ( .A1(n7541), .A2(n7616), .ZN(n8928) );
  XNOR2_X1 U9193 ( .A(n7542), .B(n8273), .ZN(n7543) );
  NAND2_X1 U9194 ( .A1(n7543), .A2(n8817), .ZN(n8929) );
  OR2_X1 U9195 ( .A1(n8858), .A2(n8861), .ZN(n7545) );
  NAND2_X1 U9196 ( .A1(n8624), .A2(n7566), .ZN(n7544) );
  NAND2_X1 U9197 ( .A1(n7545), .A2(n7544), .ZN(n8926) );
  INV_X1 U9198 ( .A(n8926), .ZN(n7546) );
  OAI211_X1 U9199 ( .C1(n7547), .C2(n8928), .A(n8929), .B(n7546), .ZN(n7552)
         );
  INV_X1 U9200 ( .A(n7589), .ZN(n7548) );
  AOI22_X1 U9201 ( .A1(n9752), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n7548), .B2(
        n8865), .ZN(n7549) );
  OAI21_X1 U9202 ( .B1(n7550), .B2(n8869), .A(n7549), .ZN(n7551) );
  AOI21_X1 U9203 ( .B1(n7552), .B2(n8826), .A(n7551), .ZN(n7553) );
  OAI21_X1 U9204 ( .B1(n7554), .B2(n8873), .A(n7553), .ZN(P2_U3277) );
  AOI21_X1 U9205 ( .B1(n7556), .B2(n8272), .A(n7555), .ZN(n8936) );
  INV_X1 U9206 ( .A(n7558), .ZN(n7559) );
  AOI21_X1 U9207 ( .B1(n8932), .B2(n4553), .A(n7559), .ZN(n8933) );
  INV_X1 U9208 ( .A(n7560), .ZN(n7561) );
  AOI22_X1 U9209 ( .A1(n9752), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n7561), .B2(
        n8865), .ZN(n7562) );
  OAI21_X1 U9210 ( .B1(n7563), .B2(n8869), .A(n7562), .ZN(n7570) );
  XOR2_X1 U9211 ( .A(n8272), .B(n7564), .Z(n7568) );
  INV_X1 U9212 ( .A(n7565), .ZN(n8625) );
  AOI222_X1 U9213 ( .A1(n8817), .A2(n7568), .B1(n8623), .B2(n7567), .C1(n8625), 
        .C2(n7566), .ZN(n8935) );
  NOR2_X1 U9214 ( .A1(n8935), .A2(n9752), .ZN(n7569) );
  AOI211_X1 U9215 ( .C1(n8933), .C2(n8864), .A(n7570), .B(n7569), .ZN(n7571)
         );
  OAI21_X1 U9216 ( .B1(n8936), .B2(n8873), .A(n7571), .ZN(P2_U3278) );
  INV_X1 U9217 ( .A(n7574), .ZN(n7575) );
  NAND2_X1 U9218 ( .A1(n7576), .A2(n7575), .ZN(n7577) );
  XNOR2_X1 U9219 ( .A(n8927), .B(n8173), .ZN(n7578) );
  OR2_X1 U9220 ( .A1(n7633), .A2(n8187), .ZN(n7579) );
  NAND2_X1 U9221 ( .A1(n7578), .A2(n7579), .ZN(n7628) );
  INV_X1 U9222 ( .A(n7578), .ZN(n7581) );
  INV_X1 U9223 ( .A(n7579), .ZN(n7580) );
  NAND2_X1 U9224 ( .A1(n7581), .A2(n7580), .ZN(n7582) );
  NAND2_X1 U9225 ( .A1(n7628), .A2(n7582), .ZN(n7586) );
  INV_X1 U9226 ( .A(n7587), .ZN(n7584) );
  INV_X1 U9227 ( .A(n7586), .ZN(n7583) );
  NAND2_X1 U9228 ( .A1(n7584), .A2(n7583), .ZN(n7629) );
  INV_X1 U9229 ( .A(n7629), .ZN(n7585) );
  AOI21_X1 U9230 ( .B1(n7587), .B2(n7586), .A(n7585), .ZN(n7592) );
  NAND2_X1 U9231 ( .A1(n8580), .A2(n8926), .ZN(n7588) );
  NAND2_X1 U9232 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8722) );
  OAI211_X1 U9233 ( .C1(n8606), .C2(n7589), .A(n7588), .B(n8722), .ZN(n7590)
         );
  AOI21_X1 U9234 ( .B1(n8927), .B2(n8583), .A(n7590), .ZN(n7591) );
  OAI21_X1 U9235 ( .B1(n7592), .B2(n8587), .A(n7591), .ZN(P2_U3221) );
  NAND2_X1 U9236 ( .A1(n7593), .A2(n7896), .ZN(n7595) );
  AOI22_X1 U9237 ( .A1(n7804), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5941), .B2(
        n9172), .ZN(n7594) );
  NAND2_X1 U9238 ( .A1(n9453), .A2(n5930), .ZN(n7597) );
  NAND2_X1 U9239 ( .A1(n9353), .A2(n8508), .ZN(n7596) );
  NAND2_X1 U9240 ( .A1(n7597), .A2(n7596), .ZN(n7598) );
  XNOR2_X1 U9241 ( .A(n7598), .B(n6095), .ZN(n8467) );
  AND2_X1 U9242 ( .A1(n9002), .A2(n9353), .ZN(n7599) );
  AOI21_X1 U9243 ( .B1(n9453), .B2(n8508), .A(n7599), .ZN(n8468) );
  XNOR2_X1 U9244 ( .A(n8467), .B(n8468), .ZN(n7603) );
  OAI21_X1 U9245 ( .B1(n7603), .B2(n7602), .A(n8470), .ZN(n7604) );
  NAND2_X1 U9246 ( .A1(n7604), .A2(n9088), .ZN(n7614) );
  XNOR2_X1 U9247 ( .A(n7808), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U9248 ( .A1(n9344), .A2(n7346), .ZN(n7608) );
  NAND2_X1 U9249 ( .A1(n7869), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U9250 ( .A1(n7822), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7606) );
  NAND2_X1 U9251 ( .A1(n7244), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7605) );
  NAND4_X1 U9252 ( .A1(n7608), .A2(n7607), .A3(n7606), .A4(n7605), .ZN(n9371)
         );
  NOR2_X1 U9253 ( .A1(n9095), .A2(n9330), .ZN(n7612) );
  INV_X1 U9254 ( .A(n7609), .ZN(n9366) );
  OAI22_X1 U9255 ( .A1(n9051), .A2(n7610), .B1(n9050), .B2(n9366), .ZN(n7611)
         );
  AOI211_X1 U9256 ( .C1(P1_REG3_REG_17__SCAN_IN), .C2(P1_U3084), .A(n7612), 
        .B(n7611), .ZN(n7613) );
  OAI211_X1 U9257 ( .C1(n4517), .C2(n9102), .A(n7614), .B(n7613), .ZN(P1_U3226) );
  XNOR2_X1 U9258 ( .A(n7615), .B(n7620), .ZN(n8924) );
  AOI21_X1 U9259 ( .B1(n5344), .B2(n7616), .A(n4538), .ZN(n8921) );
  AOI22_X1 U9260 ( .A1(n9752), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n7630), .B2(
        n8865), .ZN(n7617) );
  OAI21_X1 U9261 ( .B1(n7618), .B2(n8869), .A(n7617), .ZN(n7626) );
  INV_X1 U9262 ( .A(n7619), .ZN(n7621) );
  INV_X1 U9263 ( .A(n7620), .ZN(n8275) );
  AOI21_X1 U9264 ( .B1(n7621), .B2(n8275), .A(n8857), .ZN(n7624) );
  OAI22_X1 U9265 ( .A1(n8844), .A2(n8861), .B1(n7633), .B2(n8859), .ZN(n7622)
         );
  AOI21_X1 U9266 ( .B1(n7624), .B2(n7623), .A(n7622), .ZN(n8923) );
  NOR2_X1 U9267 ( .A1(n8923), .A2(n9752), .ZN(n7625) );
  AOI211_X1 U9268 ( .C1(n8921), .C2(n8864), .A(n7626), .B(n7625), .ZN(n7627)
         );
  OAI21_X1 U9269 ( .B1(n8924), .B2(n8873), .A(n7627), .ZN(P2_U3276) );
  XNOR2_X1 U9270 ( .A(n5344), .B(n8195), .ZN(n8169) );
  NOR2_X1 U9271 ( .A1(n8858), .A2(n8187), .ZN(n8168) );
  XNOR2_X1 U9272 ( .A(n8169), .B(n8168), .ZN(n8171) );
  XNOR2_X1 U9273 ( .A(n8172), .B(n8171), .ZN(n7637) );
  INV_X1 U9274 ( .A(n7630), .ZN(n7632) );
  OAI22_X1 U9275 ( .A1(n8606), .A2(n7632), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7631), .ZN(n7635) );
  OAI22_X1 U9276 ( .A1(n8844), .A2(n8608), .B1(n8607), .B2(n7633), .ZN(n7634)
         );
  AOI211_X1 U9277 ( .C1(n5344), .C2(n8583), .A(n7635), .B(n7634), .ZN(n7636)
         );
  OAI21_X1 U9278 ( .B1(n7637), .B2(n8587), .A(n7636), .ZN(P2_U3235) );
  INV_X1 U9279 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7898) );
  OAI222_X1 U9280 ( .A1(n9495), .A2(n7898), .B1(n7639), .B2(P1_U3084), .C1(
        n9493), .C2(n7638), .ZN(P1_U3324) );
  OAI222_X1 U9281 ( .A1(n9495), .A2(n7769), .B1(n9493), .B2(n7640), .C1(n5929), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  INV_X1 U9282 ( .A(n8607), .ZN(n7641) );
  AOI22_X1 U9283 ( .A1(n7681), .A2(n8631), .B1(n7641), .B2(n8633), .ZN(n7643)
         );
  OAI211_X1 U9284 ( .C1(n7661), .C2(n8606), .A(n7643), .B(n7642), .ZN(n7648)
         );
  INV_X1 U9285 ( .A(n6761), .ZN(n7644) );
  AOI211_X1 U9286 ( .C1(n7646), .C2(n7645), .A(n8587), .B(n7644), .ZN(n7647)
         );
  AOI211_X1 U9287 ( .C1(n5207), .C2(n8583), .A(n7648), .B(n7647), .ZN(n7649)
         );
  INV_X1 U9288 ( .A(n7649), .ZN(P2_U3219) );
  OAI21_X1 U9289 ( .B1(n7650), .B2(n8262), .A(n6893), .ZN(n9807) );
  NAND2_X1 U9290 ( .A1(n7652), .A2(n7651), .ZN(n7653) );
  NAND2_X1 U9291 ( .A1(n7653), .A2(n8353), .ZN(n7654) );
  XOR2_X1 U9292 ( .A(n8262), .B(n7654), .Z(n7658) );
  OAI22_X1 U9293 ( .A1(n7656), .A2(n8861), .B1(n7655), .B2(n8859), .ZN(n7657)
         );
  AOI21_X1 U9294 ( .B1(n7658), .B2(n8817), .A(n7657), .ZN(n7659) );
  OAI21_X1 U9295 ( .B1(n9807), .B2(n7660), .A(n7659), .ZN(n9812) );
  NAND2_X1 U9296 ( .A1(n9812), .A2(n8826), .ZN(n7669) );
  OAI22_X1 U9297 ( .A1(n8826), .A2(n7662), .B1(n7661), .B2(n9742), .ZN(n7667)
         );
  NAND2_X1 U9298 ( .A1(n7663), .A2(n5207), .ZN(n7664) );
  NAND2_X1 U9299 ( .A1(n7665), .A2(n7664), .ZN(n9811) );
  NOR2_X1 U9300 ( .A1(n9811), .A2(n8736), .ZN(n7666) );
  AOI211_X1 U9301 ( .C1(n8828), .C2(n5207), .A(n7667), .B(n7666), .ZN(n7668)
         );
  OAI211_X1 U9302 ( .C1(n9807), .C2(n7670), .A(n7669), .B(n7668), .ZN(P2_U3286) );
  AOI22_X1 U9303 ( .A1(n8601), .A2(n6391), .B1(n8604), .B2(n5597), .ZN(n7675)
         );
  INV_X1 U9304 ( .A(n7672), .ZN(n7674) );
  NOR3_X1 U9305 ( .A1(n7675), .A2(n7674), .A3(n7673), .ZN(n7680) );
  OAI22_X1 U9306 ( .A1(n7678), .A2(n7677), .B1(n7676), .B2(n8607), .ZN(n7679)
         );
  NOR2_X1 U9307 ( .A1(n7680), .A2(n7679), .ZN(n7683) );
  AOI22_X1 U9308 ( .A1(n7681), .A2(n8639), .B1(n9771), .B2(n8583), .ZN(n7682)
         );
  OAI211_X1 U9309 ( .C1(n5647), .C2(n8587), .A(n7683), .B(n7682), .ZN(P2_U3239) );
  AOI22_X1 U9310 ( .A1(n9072), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9084), .B2(
        n7684), .ZN(n7689) );
  OAI21_X1 U9311 ( .B1(n7687), .B2(n7685), .A(n7686), .ZN(n9586) );
  NAND2_X1 U9312 ( .A1(n9586), .A2(n9088), .ZN(n7688) );
  OAI211_X1 U9313 ( .C1(n7690), .C2(n9095), .A(n7689), .B(n7688), .ZN(P1_U3230) );
  AND2_X1 U9314 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8651) );
  AOI21_X1 U9315 ( .B1(n8580), .B2(n7691), .A(n8651), .ZN(n7692) );
  OAI21_X1 U9316 ( .B1(n7693), .B2(n8606), .A(n7692), .ZN(n7694) );
  AOI21_X1 U9317 ( .B1(n8947), .B2(n8583), .A(n7694), .ZN(n7697) );
  NAND3_X1 U9318 ( .A1(n7695), .A2(n8601), .A3(n8627), .ZN(n7696) );
  OAI211_X1 U9319 ( .C1(n7698), .C2(n8587), .A(n7697), .B(n7696), .ZN(P2_U3243) );
  NAND2_X1 U9320 ( .A1(n7699), .A2(n8823), .ZN(n7708) );
  INV_X1 U9321 ( .A(n7700), .ZN(n7701) );
  NOR2_X1 U9322 ( .A1(n7701), .A2(n8869), .ZN(n7705) );
  OAI22_X1 U9323 ( .A1(n7703), .A2(n9742), .B1(n7702), .B2(n8826), .ZN(n7704)
         );
  AOI211_X1 U9324 ( .C1(n7706), .C2(n8864), .A(n7705), .B(n7704), .ZN(n7707)
         );
  OAI211_X1 U9325 ( .C1(n7709), .C2(n9752), .A(n7708), .B(n7707), .ZN(P2_U3267) );
  NOR2_X1 U9326 ( .A1(n7712), .A2(SI_29_), .ZN(n7710) );
  NAND2_X1 U9327 ( .A1(n7712), .A2(SI_29_), .ZN(n7713) );
  MUX2_X1 U9328 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7725), .Z(n7721) );
  NAND2_X1 U9329 ( .A1(n8978), .A2(n7896), .ZN(n7715) );
  INV_X1 U9330 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9494) );
  OR2_X1 U9331 ( .A1(n4306), .A2(n9494), .ZN(n7714) );
  NAND2_X1 U9332 ( .A1(n7244), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U9333 ( .A1(n7822), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U9334 ( .A1(n7869), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7716) );
  NAND3_X1 U9335 ( .A1(n7718), .A2(n7717), .A3(n7716), .ZN(n9103) );
  INV_X1 U9336 ( .A(n9103), .ZN(n7901) );
  OR2_X1 U9337 ( .A1(n9387), .A2(n7901), .ZN(n8014) );
  INV_X1 U9338 ( .A(n7719), .ZN(n7720) );
  NAND2_X1 U9339 ( .A1(n7720), .A2(SI_30_), .ZN(n7724) );
  NAND2_X1 U9340 ( .A1(n7722), .A2(n7721), .ZN(n7723) );
  NAND2_X1 U9341 ( .A1(n7724), .A2(n7723), .ZN(n7728) );
  MUX2_X1 U9342 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7725), .Z(n7726) );
  XNOR2_X1 U9343 ( .A(n7726), .B(SI_31_), .ZN(n7727) );
  NAND2_X1 U9344 ( .A1(n8973), .A2(n7896), .ZN(n7731) );
  INV_X1 U9345 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7729) );
  OR2_X1 U9346 ( .A1(n6120), .A2(n7729), .ZN(n7730) );
  NAND2_X1 U9347 ( .A1(n8114), .A2(n7732), .ZN(n8018) );
  NAND2_X1 U9348 ( .A1(n8014), .A2(n8018), .ZN(n8058) );
  INV_X1 U9349 ( .A(n8058), .ZN(n7904) );
  NAND2_X1 U9350 ( .A1(n7733), .A2(n7896), .ZN(n7736) );
  OR2_X1 U9351 ( .A1(n6120), .A2(n7734), .ZN(n7735) );
  XNOR2_X1 U9352 ( .A(n7887), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U9353 ( .A1(n9212), .A2(n7346), .ZN(n7742) );
  INV_X1 U9354 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U9355 ( .A1(n7822), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U9356 ( .A1(n7869), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7737) );
  OAI211_X1 U9357 ( .C1(n5700), .C2(n7739), .A(n7738), .B(n7737), .ZN(n7740)
         );
  INV_X1 U9358 ( .A(n7740), .ZN(n7741) );
  NAND2_X1 U9359 ( .A1(n7743), .A2(n7896), .ZN(n7746) );
  OR2_X1 U9360 ( .A1(n4306), .A2(n7744), .ZN(n7745) );
  NAND2_X1 U9361 ( .A1(n7761), .A2(n9094), .ZN(n7747) );
  NAND2_X1 U9362 ( .A1(n9222), .A2(n7346), .ZN(n7754) );
  INV_X1 U9363 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n7751) );
  NAND2_X1 U9364 ( .A1(n7244), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U9365 ( .A1(n4305), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7748) );
  OAI211_X1 U9366 ( .C1(n7751), .C2(n7750), .A(n7749), .B(n7748), .ZN(n7752)
         );
  INV_X1 U9367 ( .A(n7752), .ZN(n7753) );
  OR2_X1 U9368 ( .A1(n9406), .A2(n9209), .ZN(n7755) );
  NAND2_X1 U9369 ( .A1(n8155), .A2(n7755), .ZN(n7997) );
  NAND2_X1 U9370 ( .A1(n7756), .A2(n7896), .ZN(n7759) );
  OR2_X1 U9371 ( .A1(n6120), .A2(n7757), .ZN(n7758) );
  NAND2_X1 U9372 ( .A1(n7867), .A2(n9033), .ZN(n7760) );
  NAND2_X1 U9373 ( .A1(n7761), .A2(n7760), .ZN(n9234) );
  INV_X1 U9374 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U9375 ( .A1(n7869), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7763) );
  NAND2_X1 U9376 ( .A1(n7822), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7762) );
  OAI211_X1 U9377 ( .C1(n5700), .C2(n7764), .A(n7763), .B(n7762), .ZN(n7765)
         );
  INV_X1 U9378 ( .A(n7765), .ZN(n7766) );
  NOR2_X1 U9379 ( .A1(n7997), .A2(n4687), .ZN(n8086) );
  NAND2_X1 U9380 ( .A1(n7768), .A2(n7896), .ZN(n7771) );
  OR2_X1 U9381 ( .A1(n4306), .A2(n7769), .ZN(n7770) );
  INV_X1 U9382 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U9383 ( .A1(n7785), .A2(n7772), .ZN(n7773) );
  NAND2_X1 U9384 ( .A1(n7820), .A2(n7773), .ZN(n9061) );
  OR2_X1 U9385 ( .A1(n9061), .A2(n7868), .ZN(n7779) );
  INV_X1 U9386 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U9387 ( .A1(n7822), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U9388 ( .A1(n7869), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7774) );
  OAI211_X1 U9389 ( .C1(n5700), .C2(n7776), .A(n7775), .B(n7774), .ZN(n7777)
         );
  INV_X1 U9390 ( .A(n7777), .ZN(n7778) );
  NAND2_X1 U9391 ( .A1(n7779), .A2(n7778), .ZN(n9303) );
  NAND2_X1 U9392 ( .A1(n7780), .A2(n7896), .ZN(n7783) );
  OR2_X1 U9393 ( .A1(n6120), .A2(n7781), .ZN(n7782) );
  NAND2_X1 U9394 ( .A1(n7792), .A2(n9025), .ZN(n7784) );
  NAND2_X1 U9395 ( .A1(n7785), .A2(n7784), .ZN(n9294) );
  AOI22_X1 U9396 ( .A1(n7244), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n4305), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U9397 ( .A1(n7822), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7786) );
  OAI211_X1 U9398 ( .C1(n9294), .C2(n7868), .A(n7787), .B(n7786), .ZN(n9314)
         );
  INV_X1 U9399 ( .A(n9314), .ZN(n9049) );
  NAND2_X1 U9400 ( .A1(n6836), .A2(n7896), .ZN(n7790) );
  OR2_X1 U9401 ( .A1(n4306), .A2(n7788), .ZN(n7789) );
  INV_X1 U9402 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7795) );
  INV_X1 U9403 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U9404 ( .A1(n7809), .A2(n9048), .ZN(n7791) );
  NAND2_X1 U9405 ( .A1(n7792), .A2(n7791), .ZN(n9310) );
  OR2_X1 U9406 ( .A1(n9310), .A2(n7868), .ZN(n7794) );
  AOI22_X1 U9407 ( .A1(n7822), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n7869), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n7793) );
  OAI211_X1 U9408 ( .C1(n5700), .C2(n7795), .A(n7794), .B(n7793), .ZN(n9302)
         );
  INV_X1 U9409 ( .A(n9302), .ZN(n9328) );
  NAND2_X1 U9410 ( .A1(n9436), .A2(n9328), .ZN(n8025) );
  INV_X1 U9411 ( .A(n8025), .ZN(n7796) );
  NAND2_X1 U9412 ( .A1(n8024), .A2(n7796), .ZN(n7797) );
  NAND2_X1 U9413 ( .A1(n9432), .A2(n9049), .ZN(n8143) );
  NAND2_X1 U9414 ( .A1(n7797), .A2(n8143), .ZN(n7798) );
  OR2_X1 U9415 ( .A1(n8145), .A2(n7798), .ZN(n7985) );
  NAND2_X1 U9416 ( .A1(n7799), .A2(n7896), .ZN(n7801) );
  AOI22_X1 U9417 ( .A1(n7804), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9677), .B2(
        n5941), .ZN(n7800) );
  OR2_X1 U9418 ( .A1(n9448), .A2(n9330), .ZN(n8027) );
  NOR2_X1 U9419 ( .A1(n9453), .A2(n8124), .ZN(n9349) );
  INV_X1 U9420 ( .A(n9349), .ZN(n7802) );
  AND2_X1 U9421 ( .A1(n8027), .A2(n7802), .ZN(n7970) );
  NAND2_X1 U9422 ( .A1(n7803), .A2(n7896), .ZN(n7806) );
  AOI22_X1 U9423 ( .A1(n7804), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9178), .B2(
        n5941), .ZN(n7805) );
  INV_X1 U9424 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9173) );
  INV_X1 U9425 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7807) );
  INV_X1 U9426 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8994) );
  OAI21_X1 U9427 ( .B1(n7808), .B2(n7807), .A(n8994), .ZN(n7810) );
  AND2_X1 U9428 ( .A1(n7810), .A2(n7809), .ZN(n9334) );
  NAND2_X1 U9429 ( .A1(n9334), .A2(n7346), .ZN(n7814) );
  NAND2_X1 U9430 ( .A1(n7869), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7812) );
  NAND2_X1 U9431 ( .A1(n7822), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7811) );
  AND2_X1 U9432 ( .A1(n7812), .A2(n7811), .ZN(n7813) );
  OAI211_X1 U9433 ( .C1(n5700), .C2(n9173), .A(n7814), .B(n7813), .ZN(n9352)
         );
  INV_X1 U9434 ( .A(n9352), .ZN(n9082) );
  NAND2_X1 U9435 ( .A1(n9444), .A2(n9082), .ZN(n8140) );
  NAND2_X1 U9436 ( .A1(n9448), .A2(n9330), .ZN(n8139) );
  NAND2_X1 U9437 ( .A1(n8140), .A2(n8139), .ZN(n7976) );
  OR2_X1 U9438 ( .A1(n9444), .A2(n9082), .ZN(n8026) );
  AND2_X1 U9439 ( .A1(n8141), .A2(n8026), .ZN(n7978) );
  OAI211_X1 U9440 ( .C1(n7970), .C2(n7976), .A(n8024), .B(n7978), .ZN(n7815)
         );
  INV_X1 U9441 ( .A(n7815), .ZN(n7829) );
  NAND2_X1 U9442 ( .A1(n7816), .A2(n7896), .ZN(n7819) );
  OR2_X1 U9443 ( .A1(n6120), .A2(n7817), .ZN(n7818) );
  NAND2_X1 U9444 ( .A1(n7820), .A2(n8986), .ZN(n7821) );
  AND2_X1 U9445 ( .A1(n7865), .A2(n7821), .ZN(n9265) );
  NAND2_X1 U9446 ( .A1(n9265), .A2(n7346), .ZN(n7828) );
  INV_X1 U9447 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U9448 ( .A1(n7869), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U9449 ( .A1(n7822), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7823) );
  OAI211_X1 U9450 ( .C1(n5700), .C2(n7825), .A(n7824), .B(n7823), .ZN(n7826)
         );
  INV_X1 U9451 ( .A(n7826), .ZN(n7827) );
  OAI211_X1 U9452 ( .C1(n7985), .C2(n7829), .A(n8147), .B(n8144), .ZN(n8083)
         );
  INV_X1 U9453 ( .A(n8083), .ZN(n7878) );
  NOR2_X1 U9454 ( .A1(n7985), .A2(n4699), .ZN(n8079) );
  NAND2_X1 U9455 ( .A1(n9453), .A2(n8124), .ZN(n7971) );
  AND2_X1 U9456 ( .A1(n7971), .A2(n8137), .ZN(n7830) );
  NAND2_X1 U9457 ( .A1(n8139), .A2(n7830), .ZN(n7858) );
  NAND2_X1 U9458 ( .A1(n7832), .A2(n7831), .ZN(n7851) );
  AND2_X1 U9459 ( .A1(n7851), .A2(n7833), .ZN(n7854) );
  INV_X1 U9460 ( .A(n7854), .ZN(n7961) );
  NAND2_X1 U9461 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  NAND2_X1 U9462 ( .A1(n7949), .A2(n7836), .ZN(n7951) );
  NAND3_X1 U9463 ( .A1(n7848), .A2(n7933), .A3(n7926), .ZN(n7837) );
  OR3_X1 U9464 ( .A1(n7961), .A2(n7951), .A3(n7837), .ZN(n7838) );
  OR3_X1 U9465 ( .A1(n7858), .A2(n4706), .A3(n7838), .ZN(n8077) );
  INV_X1 U9466 ( .A(n6674), .ZN(n7847) );
  AOI21_X1 U9467 ( .B1(n7839), .B2(n9118), .A(n8092), .ZN(n7845) );
  INV_X1 U9468 ( .A(n7840), .ZN(n7843) );
  NAND2_X1 U9469 ( .A1(n7841), .A2(n9120), .ZN(n7842) );
  AND2_X1 U9470 ( .A1(n7843), .A2(n7842), .ZN(n7844) );
  NAND4_X1 U9471 ( .A1(n8062), .A2(n8063), .A3(n7845), .A4(n7844), .ZN(n7846)
         );
  INV_X1 U9472 ( .A(n7929), .ZN(n8072) );
  AOI21_X1 U9473 ( .B1(n7847), .B2(n7846), .A(n8072), .ZN(n7859) );
  INV_X1 U9474 ( .A(n7940), .ZN(n7935) );
  OAI21_X1 U9475 ( .B1(n7936), .B2(n7935), .A(n7848), .ZN(n7849) );
  OAI21_X1 U9476 ( .B1(n7951), .B2(n7849), .A(n7954), .ZN(n7853) );
  INV_X1 U9477 ( .A(n7953), .ZN(n7850) );
  NAND2_X1 U9478 ( .A1(n7851), .A2(n7850), .ZN(n7852) );
  NAND2_X1 U9479 ( .A1(n7852), .A2(n7960), .ZN(n7959) );
  AOI21_X1 U9480 ( .B1(n7854), .B2(n7853), .A(n7959), .ZN(n7855) );
  OAI211_X1 U9481 ( .C1(n7855), .C2(n4706), .A(n8135), .B(n7967), .ZN(n7856)
         );
  INV_X1 U9482 ( .A(n7856), .ZN(n7857) );
  OR2_X1 U9483 ( .A1(n7858), .A2(n7857), .ZN(n8075) );
  OAI21_X1 U9484 ( .B1(n8077), .B2(n7859), .A(n8075), .ZN(n7860) );
  NAND2_X1 U9485 ( .A1(n8079), .A2(n7860), .ZN(n7877) );
  NAND2_X1 U9486 ( .A1(n7861), .A2(n7896), .ZN(n7864) );
  OR2_X1 U9487 ( .A1(n6120), .A2(n7862), .ZN(n7863) );
  INV_X1 U9488 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U9489 ( .A1(n7865), .A2(n9041), .ZN(n7866) );
  NAND2_X1 U9490 ( .A1(n7867), .A2(n7866), .ZN(n9253) );
  OR2_X1 U9491 ( .A1(n9253), .A2(n7868), .ZN(n7875) );
  INV_X1 U9492 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U9493 ( .A1(n4305), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U9494 ( .A1(n7822), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7870) );
  OAI211_X1 U9495 ( .C1(n5700), .C2(n7872), .A(n7871), .B(n7870), .ZN(n7873)
         );
  INV_X1 U9496 ( .A(n7873), .ZN(n7874) );
  INV_X1 U9497 ( .A(n9273), .ZN(n9034) );
  NAND2_X1 U9498 ( .A1(n9418), .A2(n9034), .ZN(n8148) );
  NAND2_X1 U9499 ( .A1(n9421), .A2(n9249), .ZN(n7991) );
  NAND2_X1 U9500 ( .A1(n8148), .A2(n7991), .ZN(n7876) );
  AOI21_X1 U9501 ( .B1(n7878), .B2(n7877), .A(n7876), .ZN(n7880) );
  INV_X1 U9502 ( .A(n8149), .ZN(n7879) );
  NAND2_X1 U9503 ( .A1(n9411), .A2(n9250), .ZN(n8151) );
  OAI21_X1 U9504 ( .B1(n7880), .B2(n7879), .A(n8151), .ZN(n7895) );
  NAND2_X1 U9505 ( .A1(n7881), .A2(n7896), .ZN(n7884) );
  OR2_X1 U9506 ( .A1(n4306), .A2(n7882), .ZN(n7883) );
  INV_X1 U9507 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7886) );
  INV_X1 U9508 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7885) );
  OAI21_X1 U9509 ( .B1(n7887), .B2(n7886), .A(n7885), .ZN(n7888) );
  INV_X1 U9510 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U9511 ( .A1(n7822), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U9512 ( .A1(n4305), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7890) );
  OAI211_X1 U9513 ( .C1(n5700), .C2(n7892), .A(n7891), .B(n7890), .ZN(n7893)
         );
  NAND2_X1 U9514 ( .A1(n9396), .A2(n9208), .ZN(n8021) );
  NAND2_X1 U9515 ( .A1(n9403), .A2(n9096), .ZN(n8022) );
  NAND2_X1 U9516 ( .A1(n8021), .A2(n8022), .ZN(n7906) );
  AND2_X1 U9517 ( .A1(n9406), .A2(n9209), .ZN(n8154) );
  AND2_X1 U9518 ( .A1(n8155), .A2(n8154), .ZN(n7894) );
  OR2_X1 U9519 ( .A1(n7906), .A2(n7894), .ZN(n8084) );
  AOI21_X1 U9520 ( .B1(n8086), .B2(n7895), .A(n8084), .ZN(n7902) );
  NAND2_X1 U9521 ( .A1(n7897), .A2(n7896), .ZN(n7900) );
  OR2_X1 U9522 ( .A1(n6120), .A2(n7898), .ZN(n7899) );
  OR2_X1 U9523 ( .A1(n9392), .A2(n9197), .ZN(n8002) );
  NAND2_X1 U9524 ( .A1(n8002), .A2(n8158), .ZN(n8089) );
  NAND2_X1 U9525 ( .A1(n9387), .A2(n7901), .ZN(n8056) );
  NAND2_X1 U9526 ( .A1(n9392), .A2(n9197), .ZN(n8087) );
  OAI211_X1 U9527 ( .C1(n7902), .C2(n8089), .A(n8056), .B(n8087), .ZN(n7903)
         );
  AOI21_X1 U9528 ( .B1(n7904), .B2(n7903), .A(n8091), .ZN(n7905) );
  XNOR2_X1 U9529 ( .A(n7905), .B(n8097), .ZN(n8106) );
  NAND2_X1 U9530 ( .A1(n8002), .A2(n8087), .ZN(n8159) );
  INV_X1 U9531 ( .A(n8159), .ZN(n8055) );
  INV_X1 U9532 ( .A(n7906), .ZN(n8000) );
  INV_X1 U9533 ( .A(n8147), .ZN(n7907) );
  NAND2_X1 U9534 ( .A1(n8148), .A2(n7907), .ZN(n7908) );
  NAND3_X1 U9535 ( .A1(n8152), .A2(n8149), .A3(n7908), .ZN(n7913) );
  INV_X1 U9536 ( .A(n7991), .ZN(n7909) );
  NAND2_X1 U9537 ( .A1(n8149), .A2(n7909), .ZN(n7910) );
  AND2_X1 U9538 ( .A1(n7910), .A2(n8148), .ZN(n7911) );
  AND2_X1 U9539 ( .A1(n7911), .A2(n8151), .ZN(n8081) );
  INV_X1 U9540 ( .A(n8081), .ZN(n7912) );
  INV_X1 U9541 ( .A(n8016), .ZN(n8010) );
  MUX2_X1 U9542 ( .A(n7913), .B(n7912), .S(n8010), .Z(n7996) );
  NAND2_X1 U9543 ( .A1(n7918), .A2(n7914), .ZN(n8066) );
  INV_X1 U9544 ( .A(n8066), .ZN(n7915) );
  NAND2_X1 U9545 ( .A1(n7916), .A2(n7915), .ZN(n7923) );
  INV_X1 U9546 ( .A(n7917), .ZN(n7919) );
  NAND2_X1 U9547 ( .A1(n7919), .A2(n7918), .ZN(n7921) );
  NAND2_X1 U9548 ( .A1(n7921), .A2(n7920), .ZN(n8068) );
  NOR2_X1 U9549 ( .A1(n8068), .A2(n8016), .ZN(n7922) );
  NAND2_X1 U9550 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  NAND2_X1 U9551 ( .A1(n7924), .A2(n8034), .ZN(n7927) );
  NAND3_X1 U9552 ( .A1(n7927), .A2(n7929), .A3(n8070), .ZN(n7925) );
  NAND2_X1 U9553 ( .A1(n7925), .A2(n7926), .ZN(n7932) );
  OAI211_X1 U9554 ( .C1(n7928), .C2(n7927), .A(n8067), .B(n7926), .ZN(n7930)
         );
  NAND2_X1 U9555 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  MUX2_X1 U9556 ( .A(n7932), .B(n7931), .S(n8016), .Z(n7942) );
  OAI211_X1 U9557 ( .C1(n7942), .C2(n7941), .A(n7940), .B(n7939), .ZN(n7945)
         );
  INV_X1 U9558 ( .A(n7943), .ZN(n7944) );
  NAND2_X1 U9559 ( .A1(n7945), .A2(n7944), .ZN(n7946) );
  NAND2_X1 U9560 ( .A1(n7946), .A2(n7950), .ZN(n7947) );
  NAND2_X1 U9561 ( .A1(n7947), .A2(n8010), .ZN(n7948) );
  AND2_X1 U9562 ( .A1(n7951), .A2(n7950), .ZN(n7952) );
  NOR2_X1 U9563 ( .A1(n7961), .A2(n7952), .ZN(n7956) );
  AND3_X1 U9564 ( .A1(n7960), .A2(n7954), .A3(n7953), .ZN(n7955) );
  MUX2_X1 U9565 ( .A(n7956), .B(n7955), .S(n8016), .Z(n7957) );
  NAND2_X1 U9566 ( .A1(n7958), .A2(n7957), .ZN(n7965) );
  INV_X1 U9567 ( .A(n7959), .ZN(n7963) );
  NAND2_X1 U9568 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  MUX2_X1 U9569 ( .A(n7963), .B(n7962), .S(n8016), .Z(n7964) );
  INV_X1 U9570 ( .A(n8122), .ZN(n8049) );
  MUX2_X1 U9571 ( .A(n7967), .B(n7966), .S(n8010), .Z(n7968) );
  XNOR2_X1 U9572 ( .A(n9453), .B(n8124), .ZN(n9376) );
  INV_X1 U9573 ( .A(n9376), .ZN(n9360) );
  MUX2_X1 U9574 ( .A(n8135), .B(n8137), .S(n8016), .Z(n7969) );
  INV_X1 U9575 ( .A(n7970), .ZN(n7973) );
  NAND2_X1 U9576 ( .A1(n8139), .A2(n7971), .ZN(n7972) );
  MUX2_X1 U9577 ( .A(n7973), .B(n7972), .S(n8010), .Z(n7974) );
  INV_X1 U9578 ( .A(n7974), .ZN(n7975) );
  INV_X1 U9579 ( .A(n7976), .ZN(n7977) );
  NAND2_X1 U9580 ( .A1(n7980), .A2(n7977), .ZN(n7979) );
  NAND3_X1 U9581 ( .A1(n7980), .A2(n8027), .A3(n8026), .ZN(n7981) );
  AOI21_X1 U9582 ( .B1(n7982), .B2(n8144), .A(n8145), .ZN(n7990) );
  INV_X1 U9583 ( .A(n7983), .ZN(n7984) );
  NAND2_X1 U9584 ( .A1(n7984), .A2(n8024), .ZN(n7988) );
  INV_X1 U9585 ( .A(n7985), .ZN(n7987) );
  INV_X1 U9586 ( .A(n8144), .ZN(n7986) );
  AOI21_X1 U9587 ( .B1(n7988), .B2(n7987), .A(n7986), .ZN(n7989) );
  MUX2_X1 U9588 ( .A(n7990), .B(n7989), .S(n8016), .Z(n7993) );
  NAND2_X1 U9589 ( .A1(n8147), .A2(n7991), .ZN(n9260) );
  INV_X1 U9590 ( .A(n9260), .ZN(n9271) );
  NAND3_X1 U9591 ( .A1(n9271), .A2(n8149), .A3(n8148), .ZN(n7992) );
  NOR2_X1 U9592 ( .A1(n7993), .A2(n7992), .ZN(n7995) );
  XNOR2_X1 U9593 ( .A(n9406), .B(n9209), .ZN(n9218) );
  MUX2_X1 U9594 ( .A(n8152), .B(n8151), .S(n8016), .Z(n7994) );
  OAI211_X1 U9595 ( .C1(n7996), .C2(n7995), .A(n8153), .B(n7994), .ZN(n7999)
         );
  NAND2_X1 U9596 ( .A1(n7997), .A2(n8016), .ZN(n7998) );
  NAND2_X1 U9597 ( .A1(n7999), .A2(n7998), .ZN(n8006) );
  NAND2_X1 U9598 ( .A1(n8000), .A2(n8006), .ZN(n8001) );
  NAND2_X1 U9599 ( .A1(n8001), .A2(n8158), .ZN(n8004) );
  INV_X1 U9600 ( .A(n8002), .ZN(n8003) );
  AOI21_X1 U9601 ( .B1(n8055), .B2(n8004), .A(n8003), .ZN(n8012) );
  INV_X1 U9602 ( .A(n8154), .ZN(n9204) );
  NAND2_X1 U9603 ( .A1(n8022), .A2(n9204), .ZN(n8005) );
  OAI211_X1 U9604 ( .C1(n8006), .C2(n8005), .A(n8155), .B(n8158), .ZN(n8007)
         );
  NAND2_X1 U9605 ( .A1(n8007), .A2(n8021), .ZN(n8009) );
  INV_X1 U9606 ( .A(n8087), .ZN(n8008) );
  AOI21_X1 U9607 ( .B1(n8009), .B2(n8055), .A(n8008), .ZN(n8011) );
  NAND2_X1 U9608 ( .A1(n8119), .A2(n9103), .ZN(n8013) );
  NAND2_X1 U9609 ( .A1(n9387), .A2(n8013), .ZN(n8088) );
  NAND2_X1 U9610 ( .A1(n8014), .A2(n8119), .ZN(n8015) );
  NAND2_X1 U9611 ( .A1(n8015), .A2(n8114), .ZN(n8094) );
  INV_X1 U9612 ( .A(n8088), .ZN(n8017) );
  NAND3_X1 U9613 ( .A1(n8018), .A2(n8017), .A3(n8016), .ZN(n8019) );
  INV_X1 U9614 ( .A(n8091), .ZN(n8100) );
  AND2_X1 U9615 ( .A1(n8019), .A2(n8100), .ZN(n8020) );
  NAND2_X1 U9616 ( .A1(n8158), .A2(n8021), .ZN(n9188) );
  INV_X1 U9617 ( .A(n9188), .ZN(n9194) );
  NAND2_X1 U9618 ( .A1(n8152), .A2(n8151), .ZN(n9239) );
  OR2_X1 U9619 ( .A1(n9418), .A2(n9273), .ZN(n8129) );
  INV_X1 U9620 ( .A(n8129), .ZN(n8023) );
  AND2_X1 U9621 ( .A1(n9418), .A2(n9273), .ZN(n8130) );
  INV_X1 U9622 ( .A(n8145), .ZN(n9268) );
  NAND2_X1 U9623 ( .A1(n8024), .A2(n8143), .ZN(n9298) );
  NAND2_X1 U9624 ( .A1(n8141), .A2(n8025), .ZN(n9316) );
  NAND2_X1 U9625 ( .A1(n8027), .A2(n8139), .ZN(n9348) );
  INV_X1 U9626 ( .A(n9348), .ZN(n8050) );
  NOR4_X1 U9627 ( .A1(n8031), .A2(n8030), .A3(n8029), .A4(n8028), .ZN(n8035)
         );
  NAND4_X1 U9628 ( .A1(n8035), .A2(n8034), .A3(n8033), .A4(n8032), .ZN(n8039)
         );
  NOR4_X1 U9629 ( .A1(n8039), .A2(n8038), .A3(n6681), .A4(n8037), .ZN(n8043)
         );
  NAND4_X1 U9630 ( .A1(n8043), .A2(n8042), .A3(n8041), .A4(n8040), .ZN(n8044)
         );
  NOR4_X1 U9631 ( .A1(n8047), .A2(n8046), .A3(n8045), .A4(n8044), .ZN(n8048)
         );
  NAND4_X1 U9632 ( .A1(n8050), .A2(n8049), .A3(n8048), .A4(n9360), .ZN(n8051)
         );
  NOR4_X1 U9633 ( .A1(n9298), .A2(n9316), .A3(n4696), .A4(n8051), .ZN(n8052)
         );
  NAND4_X1 U9634 ( .A1(n9246), .A2(n9271), .A3(n9285), .A4(n8052), .ZN(n8053)
         );
  NOR4_X1 U9635 ( .A1(n9205), .A2(n9218), .A3(n9239), .A4(n8053), .ZN(n8054)
         );
  NAND4_X1 U9636 ( .A1(n8056), .A2(n8055), .A3(n9194), .A4(n8054), .ZN(n8057)
         );
  NOR3_X1 U9637 ( .A1(n8058), .A2(n8091), .A3(n8057), .ZN(n8059) );
  NOR2_X1 U9638 ( .A1(n8059), .A2(n5900), .ZN(n8096) );
  INV_X1 U9639 ( .A(n8096), .ZN(n8060) );
  OAI21_X1 U9640 ( .B1(n8101), .B2(n8061), .A(n8060), .ZN(n8099) );
  NAND3_X1 U9641 ( .A1(n8064), .A2(n8063), .A3(n8062), .ZN(n8074) );
  NOR2_X1 U9642 ( .A1(n8066), .A2(n8065), .ZN(n8069) );
  OAI21_X1 U9643 ( .B1(n8069), .B2(n8068), .A(n8067), .ZN(n8071) );
  NAND2_X1 U9644 ( .A1(n8071), .A2(n8070), .ZN(n8073) );
  AOI21_X1 U9645 ( .B1(n8074), .B2(n8073), .A(n8072), .ZN(n8076) );
  OAI21_X1 U9646 ( .B1(n8077), .B2(n8076), .A(n8075), .ZN(n8078) );
  NAND2_X1 U9647 ( .A1(n8079), .A2(n8078), .ZN(n8080) );
  NAND2_X1 U9648 ( .A1(n8080), .A2(n8149), .ZN(n8082) );
  OAI21_X1 U9649 ( .B1(n8083), .B2(n8082), .A(n8081), .ZN(n8085) );
  AOI21_X1 U9650 ( .B1(n8086), .B2(n8085), .A(n8084), .ZN(n8090) );
  OAI211_X1 U9651 ( .C1(n8090), .C2(n8089), .A(n8088), .B(n8087), .ZN(n8093)
         );
  AOI211_X1 U9652 ( .C1(n8094), .C2(n8093), .A(n8092), .B(n8091), .ZN(n8095)
         );
  NOR2_X1 U9653 ( .A1(n8096), .A2(n8095), .ZN(n8098) );
  MUX2_X1 U9654 ( .A(n8099), .B(n8098), .S(n8097), .Z(n8103) );
  AND4_X1 U9655 ( .A1(n8101), .A2(n5900), .A3(n8100), .A4(n5929), .ZN(n8102)
         );
  NOR2_X1 U9656 ( .A1(n8103), .A2(n8102), .ZN(n8105) );
  MUX2_X1 U9657 ( .A(n8106), .B(n8105), .S(n8104), .Z(n8113) );
  NOR4_X1 U9658 ( .A1(n8108), .A2(n8107), .A3(n5736), .A4(n8117), .ZN(n8111)
         );
  OAI21_X1 U9659 ( .B1(n8109), .B2(n8112), .A(P1_B_REG_SCAN_IN), .ZN(n8110) );
  OAI22_X1 U9660 ( .A1(n8113), .A2(n8112), .B1(n8111), .B2(n8110), .ZN(
        P1_U3240) );
  INV_X1 U9661 ( .A(n9448), .ZN(n9346) );
  INV_X1 U9662 ( .A(n9444), .ZN(n9337) );
  NAND2_X1 U9663 ( .A1(n9280), .A2(n9267), .ZN(n9262) );
  INV_X1 U9664 ( .A(n8131), .ZN(n9181) );
  NOR2_X1 U9665 ( .A1(n9387), .A2(n9181), .ZN(n8115) );
  XNOR2_X1 U9666 ( .A(n8115), .B(n8114), .ZN(n9384) );
  NAND2_X1 U9667 ( .A1(n9384), .A2(n9322), .ZN(n8121) );
  INV_X1 U9668 ( .A(P1_B_REG_SCAN_IN), .ZN(n8116) );
  NOR2_X1 U9669 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  NOR2_X1 U9670 ( .A1(n9329), .A2(n8118), .ZN(n8162) );
  NAND2_X1 U9671 ( .A1(n8162), .A2(n8119), .ZN(n9389) );
  NOR2_X1 U9672 ( .A1(n9319), .A2(n9389), .ZN(n9182) );
  AOI21_X1 U9673 ( .B1(n9356), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9182), .ZN(
        n8120) );
  OAI211_X1 U9674 ( .C1(n9386), .C2(n9364), .A(n8121), .B(n8120), .ZN(P1_U3261) );
  AOI22_X2 U9675 ( .A1(n8123), .A2(n8122), .B1(n9459), .B2(n9379), .ZN(n9361)
         );
  NOR2_X1 U9676 ( .A1(n9453), .A2(n9353), .ZN(n8125) );
  INV_X1 U9677 ( .A(n9436), .ZN(n9313) );
  AOI22_X1 U9678 ( .A1(n9292), .A2(n9298), .B1(n9314), .B2(n9432), .ZN(n9279)
         );
  NAND2_X1 U9679 ( .A1(n9426), .A2(n9303), .ZN(n8127) );
  OAI21_X1 U9680 ( .B1(n9421), .B2(n9287), .A(n9261), .ZN(n8128) );
  OAI21_X2 U9681 ( .B1(n9267), .B2(n9249), .A(n8128), .ZN(n9245) );
  INV_X1 U9682 ( .A(n9411), .ZN(n9237) );
  NAND2_X1 U9683 ( .A1(n9189), .A2(n9188), .ZN(n9187) );
  INV_X1 U9684 ( .A(n9396), .ZN(n9193) );
  AOI211_X1 U9685 ( .C1(n9190), .C2(n9392), .A(n8131), .B(n9696), .ZN(n9391)
         );
  INV_X1 U9686 ( .A(n9392), .ZN(n8134) );
  AOI22_X1 U9687 ( .A1(n8132), .A2(n9343), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9319), .ZN(n8133) );
  OAI21_X1 U9688 ( .B1(n8134), .B2(n9364), .A(n8133), .ZN(n8166) );
  NOR2_X1 U9689 ( .A1(n9348), .A2(n9349), .ZN(n8138) );
  NAND2_X1 U9690 ( .A1(n9350), .A2(n8139), .ZN(n9326) );
  INV_X1 U9691 ( .A(n8141), .ZN(n9299) );
  NOR2_X1 U9692 ( .A1(n9298), .A2(n9299), .ZN(n8142) );
  NAND2_X1 U9693 ( .A1(n9300), .A2(n8143), .ZN(n9286) );
  NAND2_X1 U9694 ( .A1(n9286), .A2(n8144), .ZN(n9269) );
  NOR2_X1 U9695 ( .A1(n9260), .A2(n8145), .ZN(n8146) );
  NAND2_X1 U9696 ( .A1(n9269), .A2(n8146), .ZN(n9270) );
  NAND2_X1 U9697 ( .A1(n9270), .A2(n8147), .ZN(n9247) );
  NAND2_X1 U9698 ( .A1(n9247), .A2(n8148), .ZN(n8150) );
  NAND2_X1 U9699 ( .A1(n8150), .A2(n8149), .ZN(n9238) );
  NOR2_X1 U9700 ( .A1(n9205), .A2(n8154), .ZN(n8157) );
  INV_X1 U9701 ( .A(n8155), .ZN(n8156) );
  AOI21_X1 U9702 ( .B1(n9225), .B2(n8157), .A(n8156), .ZN(n9195) );
  OAI21_X1 U9703 ( .B1(n9195), .B2(n9188), .A(n8158), .ZN(n8160) );
  XNOR2_X1 U9704 ( .A(n8160), .B(n8159), .ZN(n8161) );
  NAND2_X1 U9705 ( .A1(n8161), .A2(n9355), .ZN(n8164) );
  INV_X1 U9706 ( .A(n9208), .ZN(n9104) );
  NOR2_X1 U9707 ( .A1(n9394), .A2(n9319), .ZN(n8165) );
  OAI21_X1 U9708 ( .B1(n9395), .B2(n9383), .A(n8167), .ZN(P1_U3355) );
  NOR2_X1 U9709 ( .A1(n8845), .A2(n8187), .ZN(n8563) );
  NAND2_X1 U9710 ( .A1(n8621), .A2(n8250), .ZN(n8603) );
  XNOR2_X1 U9711 ( .A(n8842), .B(n8195), .ZN(n8177) );
  INV_X1 U9712 ( .A(n8177), .ZN(n8599) );
  NAND2_X1 U9713 ( .A1(n8169), .A2(n8168), .ZN(n8170) );
  XNOR2_X1 U9714 ( .A(n8916), .B(n8173), .ZN(n8174) );
  NOR2_X1 U9715 ( .A1(n8844), .A2(n8187), .ZN(n8175) );
  XNOR2_X1 U9716 ( .A(n8174), .B(n8175), .ZN(n8567) );
  INV_X1 U9717 ( .A(n8174), .ZN(n8176) );
  NAND2_X1 U9718 ( .A1(n8176), .A2(n8175), .ZN(n8597) );
  XNOR2_X1 U9719 ( .A(n4501), .B(n8195), .ZN(n8179) );
  XNOR2_X1 U9720 ( .A(n8898), .B(n8195), .ZN(n8181) );
  NOR2_X1 U9721 ( .A1(n8586), .A2(n8187), .ZN(n8588) );
  NAND2_X1 U9722 ( .A1(n8589), .A2(n8588), .ZN(n8184) );
  INV_X1 U9723 ( .A(n8180), .ZN(n8182) );
  NAND2_X1 U9724 ( .A1(n8182), .A2(n8181), .ZN(n8183) );
  XOR2_X1 U9725 ( .A(n8195), .B(n8894), .Z(n8577) );
  NAND2_X1 U9726 ( .A1(n8618), .A2(n8250), .ZN(n8576) );
  XNOR2_X1 U9727 ( .A(n8889), .B(n8195), .ZN(n8546) );
  NOR2_X1 U9728 ( .A1(n8761), .A2(n8187), .ZN(n8185) );
  NAND2_X1 U9729 ( .A1(n8546), .A2(n8185), .ZN(n8186) );
  OAI21_X1 U9730 ( .B1(n8546), .B2(n8185), .A(n8186), .ZN(n8209) );
  INV_X1 U9731 ( .A(n8186), .ZN(n8193) );
  XNOR2_X1 U9732 ( .A(n8883), .B(n8195), .ZN(n8188) );
  NOR2_X1 U9733 ( .A1(n8747), .A2(n8187), .ZN(n8189) );
  NAND2_X1 U9734 ( .A1(n8188), .A2(n8189), .ZN(n8194) );
  INV_X1 U9735 ( .A(n8188), .ZN(n8191) );
  INV_X1 U9736 ( .A(n8189), .ZN(n8190) );
  NAND2_X1 U9737 ( .A1(n8191), .A2(n8190), .ZN(n8192) );
  AND2_X1 U9738 ( .A1(n8194), .A2(n8192), .ZN(n8544) );
  NAND2_X1 U9739 ( .A1(n8549), .A2(n8194), .ZN(n8199) );
  NAND2_X1 U9740 ( .A1(n8615), .A2(n8250), .ZN(n8196) );
  XNOR2_X1 U9741 ( .A(n8196), .B(n8195), .ZN(n8197) );
  XNOR2_X1 U9742 ( .A(n8878), .B(n8197), .ZN(n8198) );
  XNOR2_X1 U9743 ( .A(n8199), .B(n8198), .ZN(n8205) );
  INV_X1 U9744 ( .A(n8741), .ZN(n8201) );
  OAI22_X1 U9745 ( .A1(n8201), .A2(n8606), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8200), .ZN(n8203) );
  OAI22_X1 U9746 ( .A1(n8747), .A2(n8607), .B1(n8746), .B2(n8608), .ZN(n8202)
         );
  AOI211_X1 U9747 ( .C1(n8878), .C2(n8583), .A(n8203), .B(n8202), .ZN(n8204)
         );
  OAI21_X1 U9748 ( .B1(n8205), .B2(n8587), .A(n8204), .ZN(P2_U3222) );
  OAI222_X1 U9749 ( .A1(n8979), .A2(n8207), .B1(n8233), .B2(n8206), .C1(n8282), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OR2_X1 U9750 ( .A1(n8747), .A2(n8861), .ZN(n8211) );
  OR2_X1 U9751 ( .A1(n8809), .A2(n8859), .ZN(n8210) );
  NAND2_X1 U9752 ( .A1(n8211), .A2(n8210), .ZN(n8774) );
  OAI22_X1 U9753 ( .A1(n8779), .A2(n8606), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8212), .ZN(n8213) );
  AOI21_X1 U9754 ( .B1(n8774), .B2(n8580), .A(n8213), .ZN(n8214) );
  OAI211_X1 U9755 ( .C1(n8781), .C2(n8596), .A(n8215), .B(n8214), .ZN(P2_U3242) );
  OR2_X1 U9756 ( .A1(n8606), .A2(n9741), .ZN(n8216) );
  OAI211_X1 U9757 ( .C1(n8608), .C2(n8218), .A(n8217), .B(n8216), .ZN(n8223)
         );
  NAND2_X1 U9758 ( .A1(n8583), .A2(n8219), .ZN(n8220) );
  OAI21_X1 U9759 ( .B1(n8607), .B2(n8221), .A(n8220), .ZN(n8222) );
  NOR2_X1 U9760 ( .A1(n8223), .A2(n8222), .ZN(n8231) );
  INV_X1 U9761 ( .A(n8224), .ZN(n8228) );
  NAND2_X1 U9762 ( .A1(n8601), .A2(n8638), .ZN(n8225) );
  OAI21_X1 U9763 ( .B1(n8226), .B2(n8587), .A(n8225), .ZN(n8227) );
  NAND3_X1 U9764 ( .A1(n8229), .A2(n8228), .A3(n8227), .ZN(n8230) );
  OAI211_X1 U9765 ( .C1(n6635), .C2(n8587), .A(n8231), .B(n8230), .ZN(P2_U3229) );
  OAI222_X1 U9766 ( .A1(n8979), .A2(n8234), .B1(n8233), .B2(n8232), .C1(n5508), 
        .C2(P2_U3152), .ZN(P2_U3330) );
  INV_X1 U9767 ( .A(n8241), .ZN(n8243) );
  INV_X1 U9768 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9989) );
  NOR2_X1 U9769 ( .A1(n5097), .A2(n9989), .ZN(n8236) );
  INV_X1 U9770 ( .A(n8731), .ZN(n9525) );
  AND2_X1 U9771 ( .A1(n8731), .A2(n8614), .ZN(n8288) );
  INV_X1 U9772 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U9773 ( .A1(n5086), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U9774 ( .A1(n8237), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8238) );
  OAI211_X1 U9775 ( .C1(n8240), .C2(n8725), .A(n8239), .B(n8238), .ZN(n8727)
         );
  OAI21_X1 U9776 ( .B1(n8243), .B2(n9525), .A(n8242), .ZN(n8247) );
  NOR2_X1 U9777 ( .A1(n5097), .A2(n5705), .ZN(n8244) );
  INV_X1 U9778 ( .A(n8614), .ZN(n8245) );
  NAND2_X1 U9779 ( .A1(n9525), .A2(n8245), .ZN(n8439) );
  NOR2_X1 U9780 ( .A1(n8246), .A2(n8727), .ZN(n8444) );
  AOI21_X1 U9781 ( .B1(n8247), .B2(n8287), .A(n8444), .ZN(n8248) );
  XNOR2_X1 U9782 ( .A(n8248), .B(n9744), .ZN(n8452) );
  NAND2_X1 U9783 ( .A1(n8250), .A2(n8249), .ZN(n8451) );
  NOR2_X1 U9784 ( .A1(n8444), .A2(n8288), .ZN(n8286) );
  NAND4_X1 U9785 ( .A1(n8253), .A2(n8448), .A3(n8252), .A4(n8251), .ZN(n8257)
         );
  NOR4_X1 U9786 ( .A1(n8257), .A2(n8256), .A3(n8255), .A4(n8254), .ZN(n8260)
         );
  NAND4_X1 U9787 ( .A1(n8260), .A2(n8259), .A3(n8332), .A4(n8258), .ZN(n8263)
         );
  NOR4_X1 U9788 ( .A1(n8264), .A2(n8263), .A3(n8262), .A4(n8261), .ZN(n8265)
         );
  NAND4_X1 U9789 ( .A1(n8268), .A2(n8267), .A3(n8266), .A4(n8265), .ZN(n8269)
         );
  NOR4_X1 U9790 ( .A1(n8270), .A2(n5317), .A3(n8376), .A4(n8269), .ZN(n8271)
         );
  NAND3_X1 U9791 ( .A1(n8273), .A2(n8272), .A3(n8271), .ZN(n8274) );
  NOR4_X1 U9792 ( .A1(n8843), .A2(n8855), .A3(n8275), .A4(n8274), .ZN(n8277)
         );
  INV_X1 U9793 ( .A(n8821), .ZN(n8276) );
  NAND4_X1 U9794 ( .A1(n4666), .A2(n4662), .A3(n8277), .A4(n8276), .ZN(n8278)
         );
  NOR4_X1 U9795 ( .A1(n8279), .A2(n8759), .A3(n8771), .A4(n8278), .ZN(n8280)
         );
  NAND4_X1 U9796 ( .A1(n8286), .A2(n8287), .A3(n8280), .A4(n4649), .ZN(n8281)
         );
  XOR2_X1 U9797 ( .A(n9744), .B(n8281), .Z(n8283) );
  AOI22_X1 U9798 ( .A1(n8283), .A2(n8284), .B1(n8450), .B2(n8282), .ZN(n8449)
         );
  NOR2_X1 U9799 ( .A1(n9744), .A2(n8284), .ZN(n8285) );
  INV_X1 U9800 ( .A(n8288), .ZN(n8440) );
  NAND2_X1 U9801 ( .A1(n8394), .A2(n8289), .ZN(n8292) );
  INV_X1 U9802 ( .A(n8290), .ZN(n8291) );
  MUX2_X1 U9803 ( .A(n8292), .B(n8291), .S(n8435), .Z(n8293) );
  INV_X1 U9804 ( .A(n8293), .ZN(n8393) );
  NAND2_X1 U9805 ( .A1(n4332), .A2(n8294), .ZN(n8341) );
  NAND2_X1 U9806 ( .A1(n8323), .A2(n8321), .ZN(n8296) );
  NAND2_X1 U9807 ( .A1(n8299), .A2(n8298), .ZN(n8295) );
  MUX2_X1 U9808 ( .A(n8296), .B(n8295), .S(n8435), .Z(n8325) );
  AND2_X1 U9809 ( .A1(n8298), .A2(n8297), .ZN(n8300) );
  OAI211_X1 U9810 ( .C1(n8325), .C2(n8300), .A(n8299), .B(n8327), .ZN(n8301)
         );
  NAND2_X1 U9811 ( .A1(n8301), .A2(n8442), .ZN(n8311) );
  INV_X1 U9812 ( .A(n8325), .ZN(n8309) );
  INV_X1 U9813 ( .A(n8302), .ZN(n8312) );
  AND2_X1 U9814 ( .A1(n8312), .A2(n8303), .ZN(n8304) );
  OAI211_X1 U9815 ( .C1(n8305), .C2(n8304), .A(n8317), .B(n8313), .ZN(n8306)
         );
  NAND3_X1 U9816 ( .A1(n8306), .A2(n8316), .A3(n8442), .ZN(n8308) );
  NAND3_X1 U9817 ( .A1(n8309), .A2(n8308), .A3(n8307), .ZN(n8310) );
  NAND2_X1 U9818 ( .A1(n9794), .A2(n8636), .ZN(n8322) );
  NAND2_X1 U9819 ( .A1(n8313), .A2(n8312), .ZN(n8314) );
  NAND3_X1 U9820 ( .A1(n8316), .A2(n8315), .A3(n8314), .ZN(n8318) );
  NAND3_X1 U9821 ( .A1(n8318), .A2(n8435), .A3(n8317), .ZN(n8319) );
  AND2_X1 U9822 ( .A1(n8321), .A2(n8320), .ZN(n8324) );
  OAI211_X1 U9823 ( .C1(n8325), .C2(n8324), .A(n8323), .B(n8322), .ZN(n8326)
         );
  NOR2_X1 U9824 ( .A1(n8327), .A2(n8442), .ZN(n8328) );
  NOR2_X1 U9825 ( .A1(n8329), .A2(n8328), .ZN(n8330) );
  NAND3_X1 U9826 ( .A1(n8350), .A2(n8332), .A3(n8331), .ZN(n8339) );
  INV_X1 U9827 ( .A(n8343), .ZN(n8334) );
  MUX2_X1 U9828 ( .A(n8334), .B(n8333), .S(n8442), .Z(n8336) );
  INV_X1 U9829 ( .A(n8337), .ZN(n8335) );
  OR2_X1 U9830 ( .A1(n8336), .A2(n8335), .ZN(n8355) );
  OAI211_X1 U9831 ( .C1(n8339), .C2(n8355), .A(n8338), .B(n8337), .ZN(n8340)
         );
  AND2_X1 U9832 ( .A1(n8343), .A2(n8342), .ZN(n8352) );
  INV_X1 U9833 ( .A(n8344), .ZN(n8345) );
  NOR2_X1 U9834 ( .A1(n8346), .A2(n8345), .ZN(n8349) );
  INV_X1 U9835 ( .A(n8347), .ZN(n8348) );
  AOI21_X1 U9836 ( .B1(n8350), .B2(n8349), .A(n8348), .ZN(n8351) );
  MUX2_X1 U9837 ( .A(n8352), .B(n8351), .S(n8435), .Z(n8354) );
  NAND2_X1 U9838 ( .A1(n8354), .A2(n8353), .ZN(n8357) );
  INV_X1 U9839 ( .A(n8355), .ZN(n8356) );
  NAND2_X1 U9840 ( .A1(n8357), .A2(n8356), .ZN(n8358) );
  AND2_X1 U9841 ( .A1(n8362), .A2(n4332), .ZN(n8361) );
  INV_X1 U9842 ( .A(n8359), .ZN(n8360) );
  INV_X1 U9843 ( .A(n8362), .ZN(n8363) );
  AOI21_X1 U9844 ( .B1(n8365), .B2(n8364), .A(n8363), .ZN(n8366) );
  MUX2_X1 U9845 ( .A(n8367), .B(n8366), .S(n8435), .Z(n8375) );
  INV_X1 U9846 ( .A(n8368), .ZN(n8369) );
  MUX2_X1 U9847 ( .A(n8370), .B(n8369), .S(n8442), .Z(n8371) );
  NOR2_X1 U9848 ( .A1(n8372), .A2(n8371), .ZN(n8373) );
  OAI21_X1 U9849 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8380) );
  MUX2_X1 U9850 ( .A(n8378), .B(n8377), .S(n8442), .Z(n8379) );
  NAND3_X1 U9851 ( .A1(n8380), .A2(n5497), .A3(n8379), .ZN(n8386) );
  MUX2_X1 U9852 ( .A(n8947), .B(n8627), .S(n8442), .Z(n8381) );
  OAI21_X1 U9853 ( .B1(n8383), .B2(n8382), .A(n8381), .ZN(n8384) );
  NAND3_X1 U9854 ( .A1(n8386), .A2(n8385), .A3(n8384), .ZN(n8391) );
  MUX2_X1 U9855 ( .A(n8388), .B(n8387), .S(n8442), .Z(n8389) );
  NAND3_X1 U9856 ( .A1(n8391), .A2(n8390), .A3(n8389), .ZN(n8392) );
  INV_X1 U9857 ( .A(n8407), .ZN(n8395) );
  OR2_X1 U9858 ( .A1(n8916), .A2(n8844), .ZN(n8406) );
  INV_X1 U9859 ( .A(n8411), .ZN(n8397) );
  AOI21_X1 U9860 ( .B1(n8398), .B2(n8397), .A(n8396), .ZN(n8399) );
  INV_X1 U9861 ( .A(n8400), .ZN(n8401) );
  AOI21_X1 U9862 ( .B1(n8403), .B2(n8402), .A(n8401), .ZN(n8409) );
  NAND2_X1 U9863 ( .A1(n8405), .A2(n8404), .ZN(n8408) );
  OAI211_X1 U9864 ( .C1(n8409), .C2(n8408), .A(n8407), .B(n8406), .ZN(n8410)
         );
  NAND2_X1 U9865 ( .A1(n8410), .A2(n4326), .ZN(n8412) );
  AOI21_X1 U9866 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8414) );
  NOR2_X1 U9867 ( .A1(n8821), .A2(n8414), .ZN(n8415) );
  AOI21_X1 U9868 ( .B1(n8418), .B2(n8416), .A(n8435), .ZN(n8417) );
  OAI21_X1 U9869 ( .B1(n8435), .B2(n8419), .A(n4666), .ZN(n8421) );
  NAND2_X1 U9870 ( .A1(n8772), .A2(n8435), .ZN(n8420) );
  OAI211_X1 U9871 ( .C1(n8422), .C2(n8421), .A(n8427), .B(n8420), .ZN(n8426)
         );
  AOI21_X1 U9872 ( .B1(n8425), .B2(n8423), .A(n8435), .ZN(n8424) );
  MUX2_X1 U9873 ( .A(n8429), .B(n8428), .S(n8435), .Z(n8430) );
  NAND2_X1 U9874 ( .A1(n8615), .A2(n8442), .ZN(n8432) );
  NAND2_X1 U9875 ( .A1(n8762), .A2(n8435), .ZN(n8431) );
  MUX2_X1 U9876 ( .A(n8432), .B(n8431), .S(n8878), .Z(n8433) );
  MUX2_X1 U9877 ( .A(n4325), .B(n8436), .S(n8435), .Z(n8437) );
  NAND4_X1 U9878 ( .A1(n8440), .A2(n8439), .A3(n8438), .A4(n8437), .ZN(n8446)
         );
  INV_X1 U9879 ( .A(n8441), .ZN(n8443) );
  MUX2_X1 U9880 ( .A(n8444), .B(n8443), .S(n8442), .Z(n8445) );
  NOR4_X1 U9881 ( .A1(n9754), .A2(n5509), .A3(n8453), .A4(n8859), .ZN(n8456)
         );
  OAI21_X1 U9882 ( .B1(n8457), .B2(n8454), .A(P2_B_REG_SCAN_IN), .ZN(n8455) );
  OAI22_X1 U9883 ( .A1(n8458), .A2(n8457), .B1(n8456), .B2(n8455), .ZN(
        P2_U3244) );
  NAND2_X1 U9884 ( .A1(n9403), .A2(n5930), .ZN(n8460) );
  NAND2_X1 U9885 ( .A1(n9226), .A2(n6092), .ZN(n8459) );
  NAND2_X1 U9886 ( .A1(n8460), .A2(n8459), .ZN(n8461) );
  XNOR2_X1 U9887 ( .A(n8461), .B(n8482), .ZN(n8463) );
  AND2_X1 U9888 ( .A1(n9226), .A2(n9002), .ZN(n8462) );
  AOI21_X1 U9889 ( .B1(n9403), .B2(n8508), .A(n8462), .ZN(n8464) );
  NAND2_X1 U9890 ( .A1(n8463), .A2(n8464), .ZN(n9014) );
  INV_X1 U9891 ( .A(n8463), .ZN(n8466) );
  INV_X1 U9892 ( .A(n8464), .ZN(n8465) );
  NAND2_X1 U9893 ( .A1(n8466), .A2(n8465), .ZN(n9001) );
  NAND2_X1 U9894 ( .A1(n9014), .A2(n9001), .ZN(n8538) );
  AOI22_X1 U9895 ( .A1(n9421), .A2(n8508), .B1(n9002), .B2(n9287), .ZN(n8984)
         );
  INV_X1 U9896 ( .A(n8467), .ZN(n8469) );
  NAND2_X1 U9897 ( .A1(n9448), .A2(n5930), .ZN(n8472) );
  NAND2_X1 U9898 ( .A1(n9371), .A2(n8508), .ZN(n8471) );
  NAND2_X1 U9899 ( .A1(n8472), .A2(n8471), .ZN(n8473) );
  XNOR2_X1 U9900 ( .A(n8473), .B(n8482), .ZN(n8477) );
  NAND2_X1 U9901 ( .A1(n8476), .A2(n8477), .ZN(n9077) );
  NAND2_X1 U9902 ( .A1(n9448), .A2(n6092), .ZN(n8475) );
  NAND2_X1 U9903 ( .A1(n9371), .A2(n9002), .ZN(n8474) );
  NAND2_X1 U9904 ( .A1(n8475), .A2(n8474), .ZN(n9080) );
  INV_X1 U9905 ( .A(n8476), .ZN(n8479) );
  INV_X1 U9906 ( .A(n8477), .ZN(n8478) );
  NAND2_X1 U9907 ( .A1(n9444), .A2(n5930), .ZN(n8481) );
  NAND2_X1 U9908 ( .A1(n9352), .A2(n8508), .ZN(n8480) );
  NAND2_X1 U9909 ( .A1(n8481), .A2(n8480), .ZN(n8483) );
  XNOR2_X1 U9910 ( .A(n8483), .B(n8482), .ZN(n8486) );
  AND2_X1 U9911 ( .A1(n9352), .A2(n9002), .ZN(n8484) );
  AOI21_X1 U9912 ( .B1(n9444), .B2(n8508), .A(n8484), .ZN(n8485) );
  XNOR2_X1 U9913 ( .A(n8486), .B(n8485), .ZN(n8992) );
  INV_X1 U9914 ( .A(n8485), .ZN(n8488) );
  INV_X1 U9915 ( .A(n8486), .ZN(n8487) );
  NAND2_X1 U9916 ( .A1(n9436), .A2(n5930), .ZN(n8490) );
  NAND2_X1 U9917 ( .A1(n9302), .A2(n8508), .ZN(n8489) );
  NAND2_X1 U9918 ( .A1(n8490), .A2(n8489), .ZN(n8491) );
  XNOR2_X1 U9919 ( .A(n8491), .B(n6095), .ZN(n8493) );
  AND2_X1 U9920 ( .A1(n9302), .A2(n9002), .ZN(n8492) );
  AOI21_X1 U9921 ( .B1(n9436), .B2(n8508), .A(n8492), .ZN(n8494) );
  XNOR2_X1 U9922 ( .A(n8493), .B(n8494), .ZN(n9047) );
  INV_X1 U9923 ( .A(n8493), .ZN(n8495) );
  NAND2_X1 U9924 ( .A1(n8495), .A2(n8494), .ZN(n9021) );
  NAND2_X1 U9925 ( .A1(n9432), .A2(n5930), .ZN(n8497) );
  NAND2_X1 U9926 ( .A1(n9314), .A2(n6092), .ZN(n8496) );
  NAND2_X1 U9927 ( .A1(n8497), .A2(n8496), .ZN(n8498) );
  XNOR2_X1 U9928 ( .A(n8498), .B(n6095), .ZN(n8504) );
  INV_X1 U9929 ( .A(n8504), .ZN(n8500) );
  AND2_X1 U9930 ( .A1(n9314), .A2(n9002), .ZN(n8499) );
  AOI21_X1 U9931 ( .B1(n9432), .B2(n8508), .A(n8499), .ZN(n8503) );
  NAND2_X1 U9932 ( .A1(n8500), .A2(n8503), .ZN(n8502) );
  AND2_X1 U9933 ( .A1(n9021), .A2(n8502), .ZN(n8501) );
  INV_X1 U9934 ( .A(n8502), .ZN(n8505) );
  XNOR2_X1 U9935 ( .A(n8504), .B(n8503), .ZN(n9024) );
  OR2_X1 U9936 ( .A1(n8505), .A2(n9024), .ZN(n8512) );
  AND2_X1 U9937 ( .A1(n9303), .A2(n9002), .ZN(n8506) );
  AOI21_X1 U9938 ( .B1(n9426), .B2(n6092), .A(n8506), .ZN(n8514) );
  AND2_X1 U9939 ( .A1(n8512), .A2(n8514), .ZN(n8507) );
  NAND2_X1 U9940 ( .A1(n8513), .A2(n8507), .ZN(n9056) );
  NAND2_X1 U9941 ( .A1(n9426), .A2(n5930), .ZN(n8510) );
  NAND2_X1 U9942 ( .A1(n9303), .A2(n8508), .ZN(n8509) );
  NAND2_X1 U9943 ( .A1(n8510), .A2(n8509), .ZN(n8511) );
  XNOR2_X1 U9944 ( .A(n8511), .B(n6095), .ZN(n9057) );
  NAND2_X1 U9945 ( .A1(n9421), .A2(n5930), .ZN(n8517) );
  NAND2_X1 U9946 ( .A1(n9287), .A2(n6092), .ZN(n8516) );
  NAND2_X1 U9947 ( .A1(n8517), .A2(n8516), .ZN(n8518) );
  XNOR2_X1 U9948 ( .A(n8518), .B(n6095), .ZN(n8519) );
  AOI22_X1 U9949 ( .A1(n9418), .A2(n6092), .B1(n9002), .B2(n9273), .ZN(n8523)
         );
  NAND2_X1 U9950 ( .A1(n9418), .A2(n5930), .ZN(n8521) );
  NAND2_X1 U9951 ( .A1(n9273), .A2(n8508), .ZN(n8520) );
  NAND2_X1 U9952 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  XNOR2_X1 U9953 ( .A(n8522), .B(n6095), .ZN(n8525) );
  XOR2_X1 U9954 ( .A(n8523), .B(n8525), .Z(n9040) );
  INV_X1 U9955 ( .A(n8523), .ZN(n8524) );
  NAND2_X1 U9956 ( .A1(n9411), .A2(n5930), .ZN(n8527) );
  NAND2_X1 U9957 ( .A1(n9227), .A2(n6092), .ZN(n8526) );
  NAND2_X1 U9958 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  XNOR2_X1 U9959 ( .A(n8528), .B(n6095), .ZN(n8529) );
  AOI22_X1 U9960 ( .A1(n9411), .A2(n6092), .B1(n9002), .B2(n9227), .ZN(n8530)
         );
  XNOR2_X1 U9961 ( .A(n8529), .B(n8530), .ZN(n9032) );
  INV_X1 U9962 ( .A(n8529), .ZN(n8531) );
  AOI22_X1 U9963 ( .A1(n9406), .A2(n6092), .B1(n9002), .B2(n9240), .ZN(n8534)
         );
  AOI22_X1 U9964 ( .A1(n9406), .A2(n5930), .B1(n6092), .B2(n9240), .ZN(n8532)
         );
  XNOR2_X1 U9965 ( .A(n8532), .B(n6095), .ZN(n8533) );
  XOR2_X1 U9966 ( .A(n8534), .B(n8533), .Z(n9090) );
  INV_X1 U9967 ( .A(n8533), .ZN(n8536) );
  INV_X1 U9968 ( .A(n8534), .ZN(n8535) );
  XOR2_X1 U9969 ( .A(n8538), .B(n9000), .Z(n8543) );
  AOI22_X1 U9970 ( .A1(n9240), .A2(n9092), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8540) );
  NAND2_X1 U9971 ( .A1(n9212), .A2(n9099), .ZN(n8539) );
  OAI211_X1 U9972 ( .C1(n9208), .C2(n9095), .A(n8540), .B(n8539), .ZN(n8541)
         );
  AOI21_X1 U9973 ( .B1(n9403), .B2(n9084), .A(n8541), .ZN(n8542) );
  OAI21_X1 U9974 ( .B1(n8543), .B2(n9086), .A(n8542), .ZN(P1_U3212) );
  NOR2_X1 U9975 ( .A1(n8545), .A2(n8544), .ZN(n8548) );
  INV_X1 U9976 ( .A(n8761), .ZN(n8617) );
  NAND3_X1 U9977 ( .A1(n8546), .A2(n8601), .A3(n8617), .ZN(n8547) );
  OAI21_X1 U9978 ( .B1(n8548), .B2(n8587), .A(n8547), .ZN(n8550) );
  NAND2_X1 U9979 ( .A1(n8550), .A2(n8549), .ZN(n8556) );
  NOR2_X1 U9980 ( .A1(n8551), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8553) );
  OAI22_X1 U9981 ( .A1(n8762), .A2(n8608), .B1(n8761), .B2(n8607), .ZN(n8552)
         );
  AOI211_X1 U9982 ( .C1(n8554), .C2(n8756), .A(n8553), .B(n8552), .ZN(n8555)
         );
  OAI211_X1 U9983 ( .C1(n4547), .C2(n8596), .A(n8556), .B(n8555), .ZN(P2_U3216) );
  OAI22_X1 U9984 ( .A1(n8586), .A2(n8861), .B1(n8860), .B2(n8859), .ZN(n8816)
         );
  AOI22_X1 U9985 ( .A1(n8816), .A2(n8580), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8557) );
  OAI21_X1 U9986 ( .B1(n8824), .B2(n8606), .A(n8557), .ZN(n8561) );
  NOR2_X1 U9987 ( .A1(n8558), .A2(n4340), .ZN(n8562) );
  NOR3_X1 U9988 ( .A1(n8562), .A2(n8845), .A3(n8559), .ZN(n8560) );
  AOI211_X1 U9989 ( .C1(n8905), .C2(n8583), .A(n8561), .B(n8560), .ZN(n8566)
         );
  INV_X1 U9990 ( .A(n8562), .ZN(n8564) );
  NAND2_X1 U9991 ( .A1(n8566), .A2(n8565), .ZN(P2_U3218) );
  XNOR2_X1 U9992 ( .A(n8568), .B(n8567), .ZN(n8574) );
  INV_X1 U9993 ( .A(n8866), .ZN(n8570) );
  OAI22_X1 U9994 ( .A1(n8606), .A2(n8570), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8569), .ZN(n8572) );
  OAI22_X1 U9995 ( .A1(n8858), .A2(n8607), .B1(n8608), .B2(n8860), .ZN(n8571)
         );
  AOI211_X1 U9996 ( .C1(n8916), .C2(n8583), .A(n8572), .B(n8571), .ZN(n8573)
         );
  OAI21_X1 U9997 ( .B1(n8574), .B2(n8587), .A(n8573), .ZN(P2_U3225) );
  XNOR2_X1 U9998 ( .A(n8577), .B(n8576), .ZN(n8578) );
  XNOR2_X1 U9999 ( .A(n8575), .B(n8578), .ZN(n8585) );
  INV_X1 U10000 ( .A(n8579), .ZN(n8787) );
  OAI22_X1 U10001 ( .A1(n8761), .A2(n8861), .B1(n8586), .B2(n8859), .ZN(n8790)
         );
  AOI22_X1 U10002 ( .A1(n8790), .A2(n8580), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8581) );
  OAI21_X1 U10003 ( .B1(n8787), .B2(n8606), .A(n8581), .ZN(n8582) );
  AOI21_X1 U10004 ( .B1(n8894), .B2(n8583), .A(n8582), .ZN(n8584) );
  OAI21_X1 U10005 ( .B1(n8585), .B2(n8587), .A(n8584), .ZN(P2_U3227) );
  INV_X1 U10006 ( .A(n8586), .ZN(n8619) );
  NAND2_X1 U10007 ( .A1(n8619), .A2(n8601), .ZN(n8591) );
  OR2_X1 U10008 ( .A1(n8588), .A2(n8587), .ZN(n8590) );
  MUX2_X1 U10009 ( .A(n8591), .B(n8590), .S(n8589), .Z(n8595) );
  NOR2_X1 U10010 ( .A1(n8606), .A2(n8802), .ZN(n8593) );
  OAI22_X1 U10011 ( .A1(n8809), .A2(n8608), .B1(n8607), .B2(n8845), .ZN(n8592)
         );
  AOI211_X1 U10012 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3152), .A(n8593), 
        .B(n8592), .ZN(n8594) );
  OAI211_X1 U10013 ( .C1(n8805), .C2(n8596), .A(n8595), .B(n8594), .ZN(
        P2_U3231) );
  NAND2_X1 U10014 ( .A1(n8598), .A2(n8597), .ZN(n8600) );
  XNOR2_X1 U10015 ( .A(n8600), .B(n8599), .ZN(n8602) );
  NAND3_X1 U10016 ( .A1(n8602), .A2(n8601), .A3(n8621), .ZN(n8613) );
  INV_X1 U10017 ( .A(n8602), .ZN(n8605) );
  NAND3_X1 U10018 ( .A1(n8605), .A2(n8604), .A3(n8603), .ZN(n8612) );
  OAI22_X1 U10019 ( .A1(n8606), .A2(n8839), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10029), .ZN(n8610) );
  OAI22_X1 U10020 ( .A1(n8845), .A2(n8608), .B1(n8607), .B2(n8844), .ZN(n8609)
         );
  AOI211_X1 U10021 ( .C1(n8910), .C2(n8583), .A(n8610), .B(n8609), .ZN(n8611)
         );
  NAND3_X1 U10022 ( .A1(n8613), .A2(n8612), .A3(n8611), .ZN(P2_U3237) );
  MUX2_X1 U10023 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8727), .S(P2_U3966), .Z(
        P2_U3583) );
  MUX2_X1 U10024 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8614), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10025 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8615), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U10026 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8616), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10027 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8617), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8618), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8619), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U10030 ( .A(n8621), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8620), .Z(
        P2_U3574) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8622), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8623), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10033 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8624), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8625), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10035 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8626), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8627), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8628), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10038 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8629), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10039 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8630), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8631), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8632), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8633), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8634), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10044 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8635), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10045 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8636), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10046 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8637), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10047 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8638), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10048 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8639), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10049 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8640), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6391), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U10051 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8641), .S(P2_U3966), .Z(
        P2_U3552) );
  AOI21_X1 U10052 ( .B1(n8646), .B2(n8643), .A(n8642), .ZN(n8668) );
  XNOR2_X1 U10053 ( .A(n8668), .B(n8667), .ZN(n8644) );
  NOR2_X1 U10054 ( .A1(n8644), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8669) );
  AOI21_X1 U10055 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8644), .A(n8669), .ZN(
        n8654) );
  NAND2_X1 U10056 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  NOR2_X1 U10057 ( .A1(n8649), .A2(n5291), .ZN(n8656) );
  AOI211_X1 U10058 ( .C1(n5291), .C2(n8649), .A(n8656), .B(n9732), .ZN(n8650)
         );
  AOI211_X1 U10059 ( .C1(n9729), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n8651), .B(
        n8650), .ZN(n8653) );
  INV_X1 U10060 ( .A(n9731), .ZN(n9514) );
  NAND2_X1 U10061 ( .A1(n9514), .A2(n8667), .ZN(n8652) );
  OAI211_X1 U10062 ( .C1(n8654), .C2(n9730), .A(n8653), .B(n8652), .ZN(
        P2_U3260) );
  INV_X1 U10063 ( .A(n8655), .ZN(n8657) );
  AOI21_X1 U10064 ( .B1(n8657), .B2(n8667), .A(n8656), .ZN(n8660) );
  XNOR2_X1 U10065 ( .A(n8681), .B(n8658), .ZN(n8659) );
  NAND2_X1 U10066 ( .A1(n8659), .A2(n8660), .ZN(n8682) );
  OAI21_X1 U10067 ( .B1(n8660), .B2(n8659), .A(n8682), .ZN(n8665) );
  NOR2_X1 U10068 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8661), .ZN(n8664) );
  INV_X1 U10069 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8662) );
  NOR2_X1 U10070 ( .A1(n8724), .A2(n8662), .ZN(n8663) );
  AOI211_X1 U10071 ( .C1(n9727), .C2(n8665), .A(n8664), .B(n8663), .ZN(n8675)
         );
  NAND2_X1 U10072 ( .A1(n8681), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8679) );
  INV_X1 U10073 ( .A(n8679), .ZN(n8666) );
  AOI21_X1 U10074 ( .B1(n7330), .B2(n8676), .A(n8666), .ZN(n8673) );
  INV_X1 U10075 ( .A(n8667), .ZN(n8671) );
  INV_X1 U10076 ( .A(n8668), .ZN(n8670) );
  AOI21_X1 U10077 ( .B1(n8671), .B2(n8670), .A(n8669), .ZN(n8672) );
  NAND2_X1 U10078 ( .A1(n8673), .A2(n8672), .ZN(n8678) );
  OAI211_X1 U10079 ( .C1(n8673), .C2(n8672), .A(n9728), .B(n8678), .ZN(n8674)
         );
  OAI211_X1 U10080 ( .C1(n9731), .C2(n8676), .A(n8675), .B(n8674), .ZN(
        P2_U3261) );
  XNOR2_X1 U10081 ( .A(n8697), .B(n8677), .ZN(n8693) );
  NAND2_X1 U10082 ( .A1(n8679), .A2(n8678), .ZN(n8694) );
  XOR2_X1 U10083 ( .A(n8693), .B(n8694), .Z(n8691) );
  INV_X1 U10084 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8680) );
  XNOR2_X1 U10085 ( .A(n8697), .B(n8680), .ZN(n8685) );
  OR2_X1 U10086 ( .A1(n8681), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8683) );
  OAI211_X1 U10087 ( .C1(n8685), .C2(n8684), .A(n9727), .B(n8699), .ZN(n8688)
         );
  NOR2_X1 U10088 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5028), .ZN(n8686) );
  AOI21_X1 U10089 ( .B1(n9729), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8686), .ZN(
        n8687) );
  OAI211_X1 U10090 ( .C1(n9731), .C2(n8689), .A(n8688), .B(n8687), .ZN(n8690)
         );
  AOI21_X1 U10091 ( .B1(n8691), .B2(n9728), .A(n8690), .ZN(n8692) );
  INV_X1 U10092 ( .A(n8692), .ZN(P2_U3262) );
  AOI22_X1 U10093 ( .A1(n8694), .A2(n8693), .B1(n8697), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8711) );
  XNOR2_X1 U10094 ( .A(n8711), .B(n8707), .ZN(n8695) );
  NAND2_X1 U10095 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8695), .ZN(n8712) );
  OAI211_X1 U10096 ( .C1(n8695), .C2(P2_REG2_REG_18__SCAN_IN), .A(n9728), .B(
        n8712), .ZN(n8706) );
  XNOR2_X1 U10097 ( .A(n8707), .B(n8696), .ZN(n8701) );
  NAND2_X1 U10098 ( .A1(n8697), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8698) );
  OAI21_X1 U10099 ( .B1(n8701), .B2(n8700), .A(n8708), .ZN(n8704) );
  OAI21_X1 U10100 ( .B1(n8724), .B2(n10055), .A(n8702), .ZN(n8703) );
  AOI21_X1 U10101 ( .B1(n9727), .B2(n8704), .A(n8703), .ZN(n8705) );
  OAI211_X1 U10102 ( .C1(n9731), .C2(n8710), .A(n8706), .B(n8705), .ZN(
        P2_U3263) );
  XNOR2_X1 U10103 ( .A(n8709), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8716) );
  OR2_X1 U10104 ( .A1(n8711), .A2(n8710), .ZN(n8713) );
  NAND2_X1 U10105 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  XNOR2_X1 U10106 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8714), .ZN(n8718) );
  NAND2_X1 U10107 ( .A1(n8718), .A2(n9728), .ZN(n8715) );
  OAI211_X1 U10108 ( .C1(n8716), .C2(n9732), .A(n8715), .B(n9731), .ZN(n8720)
         );
  INV_X1 U10109 ( .A(n8716), .ZN(n8717) );
  OAI22_X1 U10110 ( .A1(n8718), .A2(n9730), .B1(n8717), .B2(n9732), .ZN(n8719)
         );
  MUX2_X1 U10111 ( .A(n8720), .B(n8719), .S(n9744), .Z(n8721) );
  INV_X1 U10112 ( .A(n8721), .ZN(n8723) );
  OAI211_X1 U10113 ( .C1(n4902), .C2(n8724), .A(n8723), .B(n8722), .ZN(
        P2_U3264) );
  XNOR2_X1 U10114 ( .A(n8874), .B(n4320), .ZN(n8876) );
  NOR2_X1 U10115 ( .A1(n8826), .A2(n8725), .ZN(n8728) );
  NAND2_X1 U10116 ( .A1(n8727), .A2(n8726), .ZN(n9521) );
  NOR2_X1 U10117 ( .A1(n9752), .A2(n9521), .ZN(n8733) );
  AOI211_X1 U10118 ( .C1(n8874), .C2(n8828), .A(n8728), .B(n8733), .ZN(n8729)
         );
  OAI21_X1 U10119 ( .B1(n8876), .B2(n8736), .A(n8729), .ZN(P2_U3265) );
  OAI21_X1 U10120 ( .B1(n8731), .B2(n8730), .A(n4320), .ZN(n9522) );
  NOR2_X1 U10121 ( .A1(n8826), .A2(n8732), .ZN(n8734) );
  AOI211_X1 U10122 ( .C1(n9525), .C2(n8828), .A(n8734), .B(n8733), .ZN(n8735)
         );
  OAI21_X1 U10123 ( .B1(n8736), .B2(n9522), .A(n8735), .ZN(P2_U3266) );
  XNOR2_X1 U10124 ( .A(n8737), .B(n4649), .ZN(n8882) );
  INV_X1 U10125 ( .A(n8755), .ZN(n8740) );
  INV_X1 U10126 ( .A(n8738), .ZN(n8739) );
  AOI21_X1 U10127 ( .B1(n8878), .B2(n8740), .A(n8739), .ZN(n8879) );
  AOI22_X1 U10128 ( .A1(n8741), .A2(n8865), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9752), .ZN(n8742) );
  OAI21_X1 U10129 ( .B1(n8743), .B2(n8869), .A(n8742), .ZN(n8751) );
  AOI211_X1 U10130 ( .C1(n8745), .C2(n8744), .A(n8857), .B(n4327), .ZN(n8749)
         );
  OAI22_X1 U10131 ( .A1(n8747), .A2(n8859), .B1(n8746), .B2(n8861), .ZN(n8748)
         );
  NOR2_X1 U10132 ( .A1(n8749), .A2(n8748), .ZN(n8881) );
  NOR2_X1 U10133 ( .A1(n8881), .A2(n9752), .ZN(n8750) );
  AOI211_X1 U10134 ( .C1(n8864), .C2(n8879), .A(n8751), .B(n8750), .ZN(n8752)
         );
  OAI21_X1 U10135 ( .B1(n8882), .B2(n8873), .A(n8752), .ZN(P2_U3268) );
  XNOR2_X1 U10136 ( .A(n8753), .B(n8759), .ZN(n8887) );
  AOI21_X1 U10137 ( .B1(n8883), .B2(n8754), .A(n8755), .ZN(n8884) );
  AOI22_X1 U10138 ( .A1(n8756), .A2(n8865), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9752), .ZN(n8757) );
  OAI21_X1 U10139 ( .B1(n4547), .B2(n8869), .A(n8757), .ZN(n8767) );
  NOR2_X1 U10140 ( .A1(n8758), .A2(n8857), .ZN(n8765) );
  OAI21_X1 U10141 ( .B1(n8770), .B2(n8760), .A(n8759), .ZN(n8764) );
  OAI22_X1 U10142 ( .A1(n8762), .A2(n8861), .B1(n8761), .B2(n8859), .ZN(n8763)
         );
  AOI21_X1 U10143 ( .B1(n8765), .B2(n8764), .A(n8763), .ZN(n8886) );
  NOR2_X1 U10144 ( .A1(n8886), .A2(n9752), .ZN(n8766) );
  AOI211_X1 U10145 ( .C1(n8864), .C2(n8884), .A(n8767), .B(n8766), .ZN(n8768)
         );
  OAI21_X1 U10146 ( .B1(n8887), .B2(n8873), .A(n8768), .ZN(P2_U3269) );
  XOR2_X1 U10147 ( .A(n8771), .B(n8769), .Z(n8892) );
  OAI21_X1 U10148 ( .B1(n8788), .B2(n8772), .A(n8771), .ZN(n8773) );
  AOI21_X1 U10149 ( .B1(n4377), .B2(n8773), .A(n8857), .ZN(n8775) );
  NOR2_X1 U10150 ( .A1(n8775), .A2(n8774), .ZN(n8891) );
  INV_X1 U10151 ( .A(n8792), .ZN(n8777) );
  INV_X1 U10152 ( .A(n8754), .ZN(n8776) );
  AOI211_X1 U10153 ( .C1(n8889), .C2(n8777), .A(n9810), .B(n8776), .ZN(n8888)
         );
  NAND2_X1 U10154 ( .A1(n8888), .A2(n9744), .ZN(n8778) );
  OAI211_X1 U10155 ( .C1(n9742), .C2(n8779), .A(n8891), .B(n8778), .ZN(n8783)
         );
  OAI22_X1 U10156 ( .A1(n8781), .A2(n8869), .B1(n8826), .B2(n8780), .ZN(n8782)
         );
  AOI21_X1 U10157 ( .B1(n8783), .B2(n8826), .A(n8782), .ZN(n8784) );
  OAI21_X1 U10158 ( .B1(n8892), .B2(n8873), .A(n8784), .ZN(P2_U3270) );
  XNOR2_X1 U10159 ( .A(n8785), .B(n8789), .ZN(n8897) );
  OAI22_X1 U10160 ( .A1(n8787), .A2(n9742), .B1(n8786), .B2(n8826), .ZN(n8795)
         );
  AOI211_X1 U10161 ( .C1(n4316), .C2(n8789), .A(n8857), .B(n8788), .ZN(n8791)
         );
  NOR2_X1 U10162 ( .A1(n8791), .A2(n8790), .ZN(n8896) );
  AOI211_X1 U10163 ( .C1(n8894), .C2(n8799), .A(n9810), .B(n8792), .ZN(n8893)
         );
  NAND2_X1 U10164 ( .A1(n8893), .A2(n9744), .ZN(n8793) );
  AOI21_X1 U10165 ( .B1(n8896), .B2(n8793), .A(n9752), .ZN(n8794) );
  AOI211_X1 U10166 ( .C1(n8828), .C2(n8894), .A(n8795), .B(n8794), .ZN(n8796)
         );
  OAI21_X1 U10167 ( .B1(n8897), .B2(n8873), .A(n8796), .ZN(P2_U3271) );
  AOI21_X1 U10168 ( .B1(n4662), .B2(n8798), .A(n8797), .ZN(n8902) );
  INV_X1 U10169 ( .A(n8819), .ZN(n8801) );
  INV_X1 U10170 ( .A(n8799), .ZN(n8800) );
  AOI21_X1 U10171 ( .B1(n8898), .B2(n8801), .A(n8800), .ZN(n8899) );
  INV_X1 U10172 ( .A(n8802), .ZN(n8803) );
  AOI22_X1 U10173 ( .A1(n9752), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8803), .B2(
        n8865), .ZN(n8804) );
  OAI21_X1 U10174 ( .B1(n8805), .B2(n8869), .A(n8804), .ZN(n8813) );
  AOI211_X1 U10175 ( .C1(n8808), .C2(n8807), .A(n8857), .B(n8806), .ZN(n8811)
         );
  OAI22_X1 U10176 ( .A1(n8809), .A2(n8861), .B1(n8845), .B2(n8859), .ZN(n8810)
         );
  NOR2_X1 U10177 ( .A1(n8811), .A2(n8810), .ZN(n8901) );
  NOR2_X1 U10178 ( .A1(n8901), .A2(n9752), .ZN(n8812) );
  AOI211_X1 U10179 ( .C1(n8899), .C2(n8864), .A(n8813), .B(n8812), .ZN(n8814)
         );
  OAI21_X1 U10180 ( .B1(n8902), .B2(n8873), .A(n8814), .ZN(P2_U3272) );
  XNOR2_X1 U10181 ( .A(n8815), .B(n8821), .ZN(n8818) );
  AOI21_X1 U10182 ( .B1(n8818), .B2(n8817), .A(n8816), .ZN(n8908) );
  AND2_X1 U10183 ( .A1(n8905), .A2(n8836), .ZN(n8820) );
  OR3_X1 U10184 ( .A1(n8820), .A2(n8819), .A3(n9810), .ZN(n8907) );
  OR2_X1 U10185 ( .A1(n8822), .A2(n8821), .ZN(n8904) );
  NAND3_X1 U10186 ( .A1(n8904), .A2(n8903), .A3(n8823), .ZN(n8830) );
  OAI22_X1 U10187 ( .A1(n8826), .A2(n8825), .B1(n8824), .B2(n9742), .ZN(n8827)
         );
  AOI21_X1 U10188 ( .B1(n8905), .B2(n8828), .A(n8827), .ZN(n8829) );
  OAI211_X1 U10189 ( .C1(n8907), .C2(n8831), .A(n8830), .B(n8829), .ZN(n8832)
         );
  INV_X1 U10190 ( .A(n8832), .ZN(n8833) );
  OAI21_X1 U10191 ( .B1(n9752), .B2(n8908), .A(n8833), .ZN(P2_U3273) );
  XNOR2_X1 U10192 ( .A(n8835), .B(n8834), .ZN(n8914) );
  INV_X1 U10193 ( .A(n8862), .ZN(n8838) );
  INV_X1 U10194 ( .A(n8836), .ZN(n8837) );
  AOI21_X1 U10195 ( .B1(n8910), .B2(n8838), .A(n8837), .ZN(n8911) );
  INV_X1 U10196 ( .A(n8839), .ZN(n8840) );
  AOI22_X1 U10197 ( .A1(n9752), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8840), .B2(
        n8865), .ZN(n8841) );
  OAI21_X1 U10198 ( .B1(n8842), .B2(n8869), .A(n8841), .ZN(n8850) );
  AOI21_X1 U10199 ( .B1(n4345), .B2(n8843), .A(n8857), .ZN(n8848) );
  OAI22_X1 U10200 ( .A1(n8845), .A2(n8861), .B1(n8844), .B2(n8859), .ZN(n8846)
         );
  AOI21_X1 U10201 ( .B1(n8848), .B2(n8847), .A(n8846), .ZN(n8913) );
  NOR2_X1 U10202 ( .A1(n8913), .A2(n9752), .ZN(n8849) );
  AOI211_X1 U10203 ( .C1(n8911), .C2(n8864), .A(n8850), .B(n8849), .ZN(n8851)
         );
  OAI21_X1 U10204 ( .B1(n8914), .B2(n8873), .A(n8851), .ZN(P2_U3274) );
  XNOR2_X1 U10205 ( .A(n8852), .B(n8855), .ZN(n8920) );
  AOI21_X1 U10206 ( .B1(n8855), .B2(n8854), .A(n8853), .ZN(n8856) );
  OAI222_X1 U10207 ( .A1(n8861), .A2(n8860), .B1(n8859), .B2(n8858), .C1(n8857), .C2(n8856), .ZN(n8915) );
  AOI21_X1 U10208 ( .B1(n8916), .B2(n8863), .A(n8862), .ZN(n8917) );
  NAND2_X1 U10209 ( .A1(n8917), .A2(n8864), .ZN(n8868) );
  AOI22_X1 U10210 ( .A1(n9752), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8866), .B2(
        n8865), .ZN(n8867) );
  OAI211_X1 U10211 ( .C1(n8870), .C2(n8869), .A(n8868), .B(n8867), .ZN(n8871)
         );
  AOI21_X1 U10212 ( .B1(n8915), .B2(n8826), .A(n8871), .ZN(n8872) );
  OAI21_X1 U10213 ( .B1(n8920), .B2(n8873), .A(n8872), .ZN(P2_U3275) );
  NAND2_X1 U10214 ( .A1(n8874), .A2(n9772), .ZN(n8875) );
  OAI211_X1 U10215 ( .C1(n8876), .C2(n9810), .A(n9521), .B(n8875), .ZN(n8957)
         );
  MUX2_X1 U10216 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8957), .S(n9830), .Z(
        P2_U3551) );
  MUX2_X1 U10217 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8877), .S(n9830), .Z(
        P2_U3549) );
  AOI22_X1 U10218 ( .A1(n8879), .A2(n9786), .B1(n9772), .B2(n8878), .ZN(n8880)
         );
  OAI211_X1 U10219 ( .C1(n8882), .C2(n9790), .A(n8881), .B(n8880), .ZN(n8958)
         );
  MUX2_X1 U10220 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8958), .S(n9830), .Z(
        P2_U3548) );
  AOI22_X1 U10221 ( .A1(n8884), .A2(n9786), .B1(n9772), .B2(n8883), .ZN(n8885)
         );
  OAI211_X1 U10222 ( .C1(n8887), .C2(n9790), .A(n8886), .B(n8885), .ZN(n8959)
         );
  MUX2_X1 U10223 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8959), .S(n9830), .Z(
        P2_U3547) );
  AOI21_X1 U10224 ( .B1(n9772), .B2(n8889), .A(n8888), .ZN(n8890) );
  OAI211_X1 U10225 ( .C1(n8892), .C2(n9790), .A(n8891), .B(n8890), .ZN(n8960)
         );
  MUX2_X1 U10226 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8960), .S(n9830), .Z(
        P2_U3546) );
  AOI21_X1 U10227 ( .B1(n9772), .B2(n8894), .A(n8893), .ZN(n8895) );
  OAI211_X1 U10228 ( .C1(n8897), .C2(n9790), .A(n8896), .B(n8895), .ZN(n8961)
         );
  MUX2_X1 U10229 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8961), .S(n9830), .Z(
        P2_U3545) );
  AOI22_X1 U10230 ( .A1(n8899), .A2(n9786), .B1(n9772), .B2(n8898), .ZN(n8900)
         );
  OAI211_X1 U10231 ( .C1(n8902), .C2(n9790), .A(n8901), .B(n8900), .ZN(n8962)
         );
  MUX2_X1 U10232 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8962), .S(n9830), .Z(
        P2_U3544) );
  NAND3_X1 U10233 ( .A1(n8904), .A2(n8903), .A3(n9800), .ZN(n8909) );
  NAND2_X1 U10234 ( .A1(n8905), .A2(n9772), .ZN(n8906) );
  NAND4_X1 U10235 ( .A1(n8909), .A2(n8908), .A3(n8907), .A4(n8906), .ZN(n8963)
         );
  MUX2_X1 U10236 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8963), .S(n9830), .Z(
        P2_U3543) );
  AOI22_X1 U10237 ( .A1(n8911), .A2(n9786), .B1(n9772), .B2(n8910), .ZN(n8912)
         );
  OAI211_X1 U10238 ( .C1(n8914), .C2(n9790), .A(n8913), .B(n8912), .ZN(n8964)
         );
  MUX2_X1 U10239 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8964), .S(n9830), .Z(
        P2_U3542) );
  INV_X1 U10240 ( .A(n8915), .ZN(n8919) );
  AOI22_X1 U10241 ( .A1(n8917), .A2(n9786), .B1(n9772), .B2(n8916), .ZN(n8918)
         );
  OAI211_X1 U10242 ( .C1(n8920), .C2(n9790), .A(n8919), .B(n8918), .ZN(n8965)
         );
  MUX2_X1 U10243 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8965), .S(n9830), .Z(
        P2_U3541) );
  AOI22_X1 U10244 ( .A1(n8921), .A2(n9786), .B1(n9772), .B2(n5344), .ZN(n8922)
         );
  OAI211_X1 U10245 ( .C1(n8924), .C2(n9790), .A(n8923), .B(n8922), .ZN(n8966)
         );
  MUX2_X1 U10246 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8966), .S(n9830), .Z(
        P2_U3540) );
  NAND2_X1 U10247 ( .A1(n8925), .A2(n9800), .ZN(n8931) );
  AOI21_X1 U10248 ( .B1(n8927), .B2(n9772), .A(n8926), .ZN(n8930) );
  NAND4_X1 U10249 ( .A1(n8931), .A2(n8930), .A3(n8929), .A4(n8928), .ZN(n8967)
         );
  MUX2_X1 U10250 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8967), .S(n9830), .Z(
        P2_U3539) );
  AOI22_X1 U10251 ( .A1(n8933), .A2(n9786), .B1(n9772), .B2(n8932), .ZN(n8934)
         );
  OAI211_X1 U10252 ( .C1(n8936), .C2(n9790), .A(n8935), .B(n8934), .ZN(n8968)
         );
  MUX2_X1 U10253 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8968), .S(n9830), .Z(
        P2_U3538) );
  AOI211_X1 U10254 ( .C1(n9772), .C2(n5318), .A(n8938), .B(n8937), .ZN(n8939)
         );
  OAI21_X1 U10255 ( .B1(n8940), .B2(n9790), .A(n8939), .ZN(n8969) );
  MUX2_X1 U10256 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8969), .S(n9830), .Z(
        P2_U3537) );
  AOI22_X1 U10257 ( .A1(n8942), .A2(n9786), .B1(n9772), .B2(n8941), .ZN(n8943)
         );
  OAI211_X1 U10258 ( .C1(n9778), .C2(n8945), .A(n8944), .B(n8943), .ZN(n8970)
         );
  MUX2_X1 U10259 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8970), .S(n9830), .Z(
        P2_U3536) );
  INV_X1 U10260 ( .A(n8946), .ZN(n8951) );
  AOI22_X1 U10261 ( .A1(n8948), .A2(n9786), .B1(n9772), .B2(n8947), .ZN(n8949)
         );
  OAI211_X1 U10262 ( .C1(n8951), .C2(n9790), .A(n8950), .B(n8949), .ZN(n8971)
         );
  MUX2_X1 U10263 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8971), .S(n9830), .Z(
        P2_U3535) );
  AOI22_X1 U10264 ( .A1(n8953), .A2(n9786), .B1(n9772), .B2(n8952), .ZN(n8954)
         );
  OAI211_X1 U10265 ( .C1(n9778), .C2(n8956), .A(n8955), .B(n8954), .ZN(n8972)
         );
  MUX2_X1 U10266 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8972), .S(n9830), .Z(
        P2_U3533) );
  MUX2_X1 U10267 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8957), .S(n9817), .Z(
        P2_U3519) );
  MUX2_X1 U10268 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8958), .S(n9817), .Z(
        P2_U3516) );
  MUX2_X1 U10269 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8959), .S(n9817), .Z(
        P2_U3515) );
  MUX2_X1 U10270 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8960), .S(n9817), .Z(
        P2_U3514) );
  MUX2_X1 U10271 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8961), .S(n9817), .Z(
        P2_U3513) );
  MUX2_X1 U10272 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8962), .S(n9817), .Z(
        P2_U3512) );
  MUX2_X1 U10273 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8963), .S(n9817), .Z(
        P2_U3511) );
  MUX2_X1 U10274 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8964), .S(n9817), .Z(
        P2_U3510) );
  MUX2_X1 U10275 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8965), .S(n9817), .Z(
        P2_U3509) );
  MUX2_X1 U10276 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8966), .S(n9817), .Z(
        P2_U3508) );
  MUX2_X1 U10277 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8967), .S(n9817), .Z(
        P2_U3507) );
  MUX2_X1 U10278 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8968), .S(n9817), .Z(
        P2_U3505) );
  MUX2_X1 U10279 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8969), .S(n9817), .Z(
        P2_U3502) );
  MUX2_X1 U10280 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8970), .S(n9817), .Z(
        P2_U3499) );
  MUX2_X1 U10281 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8971), .S(n9817), .Z(
        P2_U3496) );
  MUX2_X1 U10282 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8972), .S(n9817), .Z(
        P2_U3490) );
  INV_X1 U10283 ( .A(n8973), .ZN(n9490) );
  NAND3_X1 U10284 ( .A1(n8974), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8975) );
  OAI22_X1 U10285 ( .A1(n4465), .A2(n8975), .B1(n5705), .B2(n8979), .ZN(n8976)
         );
  INV_X1 U10286 ( .A(n8976), .ZN(n8977) );
  OAI21_X1 U10287 ( .B1(n9490), .B2(n8980), .A(n8977), .ZN(P2_U3327) );
  INV_X1 U10288 ( .A(n8978), .ZN(n9492) );
  MUX2_X1 U10289 ( .A(n8981), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10290 ( .A1(n4794), .A2(n8983), .ZN(n8985) );
  XNOR2_X1 U10291 ( .A(n8985), .B(n8984), .ZN(n8991) );
  OAI22_X1 U10292 ( .A1(n9034), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8986), .ZN(n8989) );
  INV_X1 U10293 ( .A(n9265), .ZN(n8987) );
  OAI22_X1 U10294 ( .A1(n9051), .A2(n9026), .B1(n9050), .B2(n8987), .ZN(n8988)
         );
  AOI211_X1 U10295 ( .C1(n9421), .C2(n9084), .A(n8989), .B(n8988), .ZN(n8990)
         );
  OAI21_X1 U10296 ( .B1(n8991), .B2(n9086), .A(n8990), .ZN(P1_U3214) );
  XOR2_X1 U10297 ( .A(n8993), .B(n8992), .Z(n8999) );
  OAI22_X1 U10298 ( .A1(n9095), .A2(n9328), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8994), .ZN(n8997) );
  INV_X1 U10299 ( .A(n9334), .ZN(n8995) );
  OAI22_X1 U10300 ( .A1(n9051), .A2(n9330), .B1(n9050), .B2(n8995), .ZN(n8996)
         );
  AOI211_X1 U10301 ( .C1(n9444), .C2(n9084), .A(n8997), .B(n8996), .ZN(n8998)
         );
  OAI21_X1 U10302 ( .B1(n8999), .B2(n9086), .A(n8998), .ZN(P1_U3217) );
  NAND2_X1 U10303 ( .A1(n9396), .A2(n8508), .ZN(n9005) );
  INV_X1 U10304 ( .A(n9002), .ZN(n9003) );
  OR2_X1 U10305 ( .A1(n9208), .A2(n9003), .ZN(n9004) );
  NAND2_X1 U10306 ( .A1(n9005), .A2(n9004), .ZN(n9006) );
  XNOR2_X1 U10307 ( .A(n9006), .B(n8482), .ZN(n9010) );
  NOR2_X1 U10308 ( .A1(n9208), .A2(n9007), .ZN(n9008) );
  AOI21_X1 U10309 ( .B1(n9396), .B2(n5930), .A(n9008), .ZN(n9009) );
  XNOR2_X1 U10310 ( .A(n9010), .B(n9009), .ZN(n9015) );
  NAND4_X1 U10311 ( .A1(n9011), .A2(n9088), .A3(n9014), .A4(n9015), .ZN(n9020)
         );
  AOI22_X1 U10312 ( .A1(n9191), .A2(n9099), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n9013) );
  NAND2_X1 U10313 ( .A1(n9226), .A2(n9092), .ZN(n9012) );
  OAI211_X1 U10314 ( .C1(n9197), .C2(n9095), .A(n9013), .B(n9012), .ZN(n9017)
         );
  NOR3_X1 U10315 ( .A1(n9015), .A2(n9086), .A3(n9014), .ZN(n9016) );
  AOI211_X1 U10316 ( .C1(n9396), .C2(n9084), .A(n9017), .B(n9016), .ZN(n9018)
         );
  NAND3_X1 U10317 ( .A1(n9020), .A2(n9019), .A3(n9018), .ZN(P1_U3218) );
  NAND2_X1 U10318 ( .A1(n9022), .A2(n9021), .ZN(n9023) );
  XOR2_X1 U10319 ( .A(n9024), .B(n9023), .Z(n9030) );
  OAI22_X1 U10320 ( .A1(n9026), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9025), .ZN(n9028) );
  OAI22_X1 U10321 ( .A1(n9051), .A2(n9328), .B1(n9050), .B2(n9294), .ZN(n9027)
         );
  AOI211_X1 U10322 ( .C1(n9432), .C2(n9084), .A(n9028), .B(n9027), .ZN(n9029)
         );
  OAI21_X1 U10323 ( .B1(n9030), .B2(n9086), .A(n9029), .ZN(P1_U3221) );
  XOR2_X1 U10324 ( .A(n9032), .B(n9031), .Z(n9038) );
  OAI22_X1 U10325 ( .A1(n9034), .A2(n9051), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9033), .ZN(n9036) );
  OAI22_X1 U10326 ( .A1(n9209), .A2(n9095), .B1(n9050), .B2(n9234), .ZN(n9035)
         );
  AOI211_X1 U10327 ( .C1(n9411), .C2(n9084), .A(n9036), .B(n9035), .ZN(n9037)
         );
  OAI21_X1 U10328 ( .B1(n9038), .B2(n9086), .A(n9037), .ZN(P1_U3223) );
  XOR2_X1 U10329 ( .A(n9040), .B(n9039), .Z(n9045) );
  OAI22_X1 U10330 ( .A1(n9250), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9041), .ZN(n9043) );
  OAI22_X1 U10331 ( .A1(n9249), .A2(n9051), .B1(n9050), .B2(n9253), .ZN(n9042)
         );
  AOI211_X1 U10332 ( .C1(n9418), .C2(n9084), .A(n9043), .B(n9042), .ZN(n9044)
         );
  OAI21_X1 U10333 ( .B1(n9045), .B2(n9086), .A(n9044), .ZN(P1_U3227) );
  XOR2_X1 U10334 ( .A(n9046), .B(n9047), .Z(n9055) );
  OAI22_X1 U10335 ( .A1(n9095), .A2(n9049), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9048), .ZN(n9053) );
  OAI22_X1 U10336 ( .A1(n9051), .A2(n9082), .B1(n9050), .B2(n9310), .ZN(n9052)
         );
  AOI211_X1 U10337 ( .C1(n9436), .C2(n9084), .A(n9053), .B(n9052), .ZN(n9054)
         );
  OAI21_X1 U10338 ( .B1(n9055), .B2(n9086), .A(n9054), .ZN(P1_U3231) );
  AOI21_X1 U10339 ( .B1(n4322), .B2(n9056), .A(n9057), .ZN(n9060) );
  INV_X1 U10340 ( .A(n9057), .ZN(n9058) );
  OAI22_X1 U10341 ( .A1(n9060), .A2(n9059), .B1(n9058), .B2(n4322), .ZN(n9065)
         );
  AOI22_X1 U10342 ( .A1(n9073), .A2(n9287), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9063) );
  INV_X1 U10343 ( .A(n9061), .ZN(n9282) );
  AOI22_X1 U10344 ( .A1(n9092), .A2(n9314), .B1(n9282), .B2(n9099), .ZN(n9062)
         );
  OAI211_X1 U10345 ( .C1(n9284), .C2(n9102), .A(n9063), .B(n9062), .ZN(n9064)
         );
  AOI21_X1 U10346 ( .B1(n9065), .B2(n9088), .A(n9064), .ZN(n9066) );
  INV_X1 U10347 ( .A(n9066), .ZN(P1_U3233) );
  OAI21_X1 U10348 ( .B1(n9069), .B2(n9067), .A(n9068), .ZN(n9070) );
  NAND2_X1 U10349 ( .A1(n9070), .A2(n9088), .ZN(n9076) );
  AOI22_X1 U10350 ( .A1(n9072), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n9084), .B2(
        n4307), .ZN(n9075) );
  AOI22_X1 U10351 ( .A1(n9073), .A2(n9117), .B1(n9092), .B2(n9120), .ZN(n9074)
         );
  NAND3_X1 U10352 ( .A1(n9076), .A2(n9075), .A3(n9074), .ZN(P1_U3235) );
  NAND2_X1 U10353 ( .A1(n9078), .A2(n9077), .ZN(n9079) );
  XOR2_X1 U10354 ( .A(n9080), .B(n9079), .Z(n9087) );
  AOI22_X1 U10355 ( .A1(n9092), .A2(n9353), .B1(n9344), .B2(n9099), .ZN(n9081)
         );
  NAND2_X1 U10356 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9679) );
  OAI211_X1 U10357 ( .C1(n9082), .C2(n9095), .A(n9081), .B(n9679), .ZN(n9083)
         );
  AOI21_X1 U10358 ( .B1(n9448), .B2(n9084), .A(n9083), .ZN(n9085) );
  OAI21_X1 U10359 ( .B1(n9087), .B2(n9086), .A(n9085), .ZN(P1_U3236) );
  OAI211_X1 U10360 ( .C1(n9091), .C2(n9090), .A(n9089), .B(n9088), .ZN(n9101)
         );
  NAND2_X1 U10361 ( .A1(n9227), .A2(n9092), .ZN(n9093) );
  OAI21_X1 U10362 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9094), .A(n9093), .ZN(
        n9098) );
  NOR2_X1 U10363 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  AOI211_X1 U10364 ( .C1(n9222), .C2(n9099), .A(n9098), .B(n9097), .ZN(n9100)
         );
  OAI211_X1 U10365 ( .C1(n9224), .C2(n9102), .A(n9101), .B(n9100), .ZN(
        P1_U3238) );
  MUX2_X1 U10366 ( .A(n9103), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9119), .Z(
        P1_U3585) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9104), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10368 ( .A(n9226), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9119), .Z(
        P1_U3582) );
  MUX2_X1 U10369 ( .A(n9240), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9119), .Z(
        P1_U3581) );
  MUX2_X1 U10370 ( .A(n9227), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9119), .Z(
        P1_U3580) );
  MUX2_X1 U10371 ( .A(n9273), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9119), .Z(
        P1_U3579) );
  MUX2_X1 U10372 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9287), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9303), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10374 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9314), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10375 ( .A(n9302), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9119), .Z(
        P1_U3575) );
  MUX2_X1 U10376 ( .A(n9352), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9119), .Z(
        P1_U3574) );
  MUX2_X1 U10377 ( .A(n9371), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9119), .Z(
        P1_U3573) );
  MUX2_X1 U10378 ( .A(n9353), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9119), .Z(
        P1_U3572) );
  MUX2_X1 U10379 ( .A(n9379), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9119), .Z(
        P1_U3571) );
  MUX2_X1 U10380 ( .A(n9105), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9119), .Z(
        P1_U3570) );
  MUX2_X1 U10381 ( .A(n9106), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9119), .Z(
        P1_U3569) );
  MUX2_X1 U10382 ( .A(n9107), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9119), .Z(
        P1_U3568) );
  MUX2_X1 U10383 ( .A(n9108), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9119), .Z(
        P1_U3567) );
  MUX2_X1 U10384 ( .A(n9109), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9119), .Z(
        P1_U3566) );
  MUX2_X1 U10385 ( .A(n9110), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9119), .Z(
        P1_U3565) );
  MUX2_X1 U10386 ( .A(n9111), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9119), .Z(
        P1_U3564) );
  MUX2_X1 U10387 ( .A(n9112), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9119), .Z(
        P1_U3563) );
  MUX2_X1 U10388 ( .A(n9113), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9119), .Z(
        P1_U3562) );
  MUX2_X1 U10389 ( .A(n9114), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9119), .Z(
        P1_U3561) );
  MUX2_X1 U10390 ( .A(n9115), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9119), .Z(
        P1_U3560) );
  MUX2_X1 U10391 ( .A(n9116), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9119), .Z(
        P1_U3559) );
  MUX2_X1 U10392 ( .A(n9117), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9119), .Z(
        P1_U3558) );
  MUX2_X1 U10393 ( .A(n9118), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9119), .Z(
        P1_U3557) );
  MUX2_X1 U10394 ( .A(n9120), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9119), .Z(
        P1_U3556) );
  AOI211_X1 U10395 ( .C1(n9123), .C2(n9122), .A(n9121), .B(n9637), .ZN(n9124)
         );
  AOI21_X1 U10396 ( .B1(n9678), .B2(n9125), .A(n9124), .ZN(n9133) );
  AOI21_X1 U10397 ( .B1(n9685), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n9126), .ZN(
        n9132) );
  OAI21_X1 U10398 ( .B1(n9129), .B2(n9128), .A(n9127), .ZN(n9130) );
  NAND2_X1 U10399 ( .A1(n9130), .A2(n9686), .ZN(n9131) );
  NAND3_X1 U10400 ( .A1(n9133), .A2(n9132), .A3(n9131), .ZN(P1_U3251) );
  NOR2_X1 U10401 ( .A1(n9141), .A2(n9134), .ZN(n9136) );
  NAND2_X1 U10402 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9158), .ZN(n9137) );
  OAI21_X1 U10403 ( .B1(n9158), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9137), .ZN(
        n9138) );
  AOI211_X1 U10404 ( .C1(n9139), .C2(n9138), .A(n9157), .B(n9637), .ZN(n9151)
         );
  NOR2_X1 U10405 ( .A1(n9141), .A2(n9140), .ZN(n9143) );
  NOR2_X1 U10406 ( .A1(n9143), .A2(n9142), .ZN(n9145) );
  XNOR2_X1 U10407 ( .A(n9158), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9144) );
  NOR2_X1 U10408 ( .A1(n9145), .A2(n9144), .ZN(n9152) );
  AOI211_X1 U10409 ( .C1(n9145), .C2(n9144), .A(n9152), .B(n9579), .ZN(n9150)
         );
  NAND2_X1 U10410 ( .A1(n9685), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9146) );
  OAI211_X1 U10411 ( .C1(n9592), .C2(n9148), .A(n9147), .B(n9146), .ZN(n9149)
         );
  OR3_X1 U10412 ( .A1(n9151), .A2(n9150), .A3(n9149), .ZN(P1_U3257) );
  AND2_X1 U10413 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9156) );
  AOI21_X1 U10414 ( .B1(n9158), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9152), .ZN(
        n9154) );
  XNOR2_X1 U10415 ( .A(n9172), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9153) );
  NOR2_X1 U10416 ( .A1(n9154), .A2(n9153), .ZN(n9171) );
  AOI211_X1 U10417 ( .C1(n9154), .C2(n9153), .A(n9171), .B(n9579), .ZN(n9155)
         );
  AOI211_X1 U10418 ( .C1(P1_ADDR_REG_17__SCAN_IN), .C2(n9685), .A(n9156), .B(
        n9155), .ZN(n9164) );
  INV_X1 U10419 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9159) );
  MUX2_X1 U10420 ( .A(n9159), .B(P1_REG2_REG_17__SCAN_IN), .S(n9172), .Z(n9160) );
  AOI211_X1 U10421 ( .C1(n9161), .C2(n9160), .A(n9165), .B(n9637), .ZN(n9162)
         );
  AOI21_X1 U10422 ( .B1(n9678), .B2(n9172), .A(n9162), .ZN(n9163) );
  NAND2_X1 U10423 ( .A1(n9164), .A2(n9163), .ZN(P1_U3258) );
  OR2_X1 U10424 ( .A1(n9677), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U10425 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9677), .ZN(n9166) );
  NAND2_X1 U10426 ( .A1(n9167), .A2(n9166), .ZN(n9674) );
  NOR2_X1 U10427 ( .A1(n9673), .A2(n9674), .ZN(n9672) );
  AOI21_X1 U10428 ( .B1(n9677), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9672), .ZN(
        n9168) );
  XNOR2_X1 U10429 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9168), .ZN(n9176) );
  INV_X1 U10430 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9169) );
  AOI22_X1 U10431 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9677), .B1(n9170), .B2(
        n9169), .ZN(n9684) );
  AOI21_X1 U10432 ( .B1(n9172), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9171), .ZN(
        n9683) );
  NAND2_X1 U10433 ( .A1(n9684), .A2(n9683), .ZN(n9682) );
  OAI21_X1 U10434 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9677), .A(n9682), .ZN(
        n9174) );
  XOR2_X1 U10435 ( .A(n9174), .B(n9173), .Z(n9175) );
  AOI22_X1 U10436 ( .A1(n9176), .A2(n9676), .B1(n9686), .B2(n9175), .ZN(n9179)
         );
  INV_X1 U10437 ( .A(n9175), .ZN(n9177) );
  NAND2_X1 U10438 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n9180) );
  XNOR2_X1 U10439 ( .A(n9387), .B(n9181), .ZN(n9390) );
  AOI21_X1 U10440 ( .B1(n9319), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9182), .ZN(
        n9185) );
  NAND2_X1 U10441 ( .A1(n9387), .A2(n9183), .ZN(n9184) );
  OAI211_X1 U10442 ( .C1(n9390), .C2(n9186), .A(n9185), .B(n9184), .ZN(
        P1_U3262) );
  OAI21_X1 U10443 ( .B1(n9189), .B2(n9188), .A(n9187), .ZN(n9400) );
  AOI21_X1 U10444 ( .B1(n9396), .B2(n9210), .A(n4507), .ZN(n9397) );
  AOI22_X1 U10445 ( .A1(n9191), .A2(n9343), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9319), .ZN(n9192) );
  OAI21_X1 U10446 ( .B1(n9193), .B2(n9364), .A(n9192), .ZN(n9201) );
  XNOR2_X1 U10447 ( .A(n9195), .B(n9194), .ZN(n9199) );
  NAND2_X1 U10448 ( .A1(n9226), .A2(n9380), .ZN(n9196) );
  OAI21_X1 U10449 ( .B1(n9197), .B2(n9329), .A(n9196), .ZN(n9198) );
  AOI21_X1 U10450 ( .B1(n9199), .B2(n9355), .A(n9198), .ZN(n9399) );
  NOR2_X1 U10451 ( .A1(n9399), .A2(n9319), .ZN(n9200) );
  AOI211_X1 U10452 ( .C1(n9397), .C2(n9322), .A(n9201), .B(n9200), .ZN(n9202)
         );
  OAI21_X1 U10453 ( .B1(n9400), .B2(n9383), .A(n9202), .ZN(P1_U3263) );
  XOR2_X1 U10454 ( .A(n9205), .B(n9203), .Z(n9405) );
  XNOR2_X1 U10455 ( .A(n9206), .B(n9205), .ZN(n9207) );
  OAI222_X1 U10456 ( .A1(n9331), .A2(n9209), .B1(n9329), .B2(n9208), .C1(n9207), .C2(n9374), .ZN(n9401) );
  INV_X1 U10457 ( .A(n9220), .ZN(n9211) );
  AOI211_X1 U10458 ( .C1(n9403), .C2(n9211), .A(n9696), .B(n4508), .ZN(n9402)
         );
  NAND2_X1 U10459 ( .A1(n9402), .A2(n9370), .ZN(n9214) );
  AOI22_X1 U10460 ( .A1(n9212), .A2(n9343), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9319), .ZN(n9213) );
  OAI211_X1 U10461 ( .C1(n9215), .C2(n9364), .A(n9214), .B(n9213), .ZN(n9216)
         );
  AOI21_X1 U10462 ( .B1(n9401), .B2(n9367), .A(n9216), .ZN(n9217) );
  OAI21_X1 U10463 ( .B1(n9405), .B2(n9383), .A(n9217), .ZN(P1_U3264) );
  XNOR2_X1 U10464 ( .A(n9219), .B(n9218), .ZN(n9410) );
  INV_X1 U10465 ( .A(n9233), .ZN(n9221) );
  AOI21_X1 U10466 ( .B1(n9406), .B2(n9221), .A(n9220), .ZN(n9407) );
  AOI22_X1 U10467 ( .A1(n9222), .A2(n9343), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9319), .ZN(n9223) );
  OAI21_X1 U10468 ( .B1(n9224), .B2(n9364), .A(n9223), .ZN(n9230) );
  OAI21_X1 U10469 ( .B1(n4858), .B2(n8153), .A(n9225), .ZN(n9228) );
  AOI222_X1 U10470 ( .A1(n9355), .A2(n9228), .B1(n9227), .B2(n9380), .C1(n9226), .C2(n9372), .ZN(n9409) );
  NOR2_X1 U10471 ( .A1(n9409), .A2(n9356), .ZN(n9229) );
  AOI211_X1 U10472 ( .C1(n9322), .C2(n9407), .A(n9230), .B(n9229), .ZN(n9231)
         );
  OAI21_X1 U10473 ( .B1(n9410), .B2(n9383), .A(n9231), .ZN(P1_U3265) );
  XOR2_X1 U10474 ( .A(n9239), .B(n9232), .Z(n9415) );
  AOI21_X1 U10475 ( .B1(n9411), .B2(n9251), .A(n9233), .ZN(n9412) );
  INV_X1 U10476 ( .A(n9234), .ZN(n9235) );
  AOI22_X1 U10477 ( .A1(n9235), .A2(n9343), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9319), .ZN(n9236) );
  OAI21_X1 U10478 ( .B1(n9237), .B2(n9364), .A(n9236), .ZN(n9243) );
  XNOR2_X1 U10479 ( .A(n9238), .B(n9239), .ZN(n9241) );
  AOI222_X1 U10480 ( .A1(n9355), .A2(n9241), .B1(n9240), .B2(n9372), .C1(n9273), .C2(n9380), .ZN(n9414) );
  NOR2_X1 U10481 ( .A1(n9414), .A2(n9319), .ZN(n9242) );
  AOI211_X1 U10482 ( .C1(n9322), .C2(n9412), .A(n9243), .B(n9242), .ZN(n9244)
         );
  OAI21_X1 U10483 ( .B1(n9415), .B2(n9383), .A(n9244), .ZN(P1_U3266) );
  XOR2_X1 U10484 ( .A(n9246), .B(n9245), .Z(n9420) );
  XNOR2_X1 U10485 ( .A(n9247), .B(n9246), .ZN(n9248) );
  OAI222_X1 U10486 ( .A1(n9329), .A2(n9250), .B1(n9331), .B2(n9249), .C1(n9248), .C2(n9374), .ZN(n9416) );
  INV_X1 U10487 ( .A(n9418), .ZN(n9257) );
  INV_X1 U10488 ( .A(n9251), .ZN(n9252) );
  AOI211_X1 U10489 ( .C1(n9418), .C2(n9262), .A(n9696), .B(n9252), .ZN(n9417)
         );
  NAND2_X1 U10490 ( .A1(n9417), .A2(n9370), .ZN(n9256) );
  INV_X1 U10491 ( .A(n9253), .ZN(n9254) );
  AOI22_X1 U10492 ( .A1(n9254), .A2(n9343), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9319), .ZN(n9255) );
  OAI211_X1 U10493 ( .C1(n9257), .C2(n9364), .A(n9256), .B(n9255), .ZN(n9258)
         );
  AOI21_X1 U10494 ( .B1(n9416), .B2(n9367), .A(n9258), .ZN(n9259) );
  OAI21_X1 U10495 ( .B1(n9420), .B2(n9383), .A(n9259), .ZN(P1_U3267) );
  XNOR2_X1 U10496 ( .A(n9261), .B(n9260), .ZN(n9425) );
  INV_X1 U10497 ( .A(n9280), .ZN(n9264) );
  INV_X1 U10498 ( .A(n9262), .ZN(n9263) );
  AOI21_X1 U10499 ( .B1(n9421), .B2(n9264), .A(n9263), .ZN(n9422) );
  AOI22_X1 U10500 ( .A1(n9319), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9265), .B2(
        n9343), .ZN(n9266) );
  OAI21_X1 U10501 ( .B1(n9267), .B2(n9364), .A(n9266), .ZN(n9277) );
  AND2_X1 U10502 ( .A1(n9269), .A2(n9268), .ZN(n9272) );
  OAI211_X1 U10503 ( .C1(n9272), .C2(n9271), .A(n9270), .B(n9355), .ZN(n9275)
         );
  AOI22_X1 U10504 ( .A1(n9273), .A2(n9372), .B1(n9380), .B2(n9303), .ZN(n9274)
         );
  AND2_X1 U10505 ( .A1(n9275), .A2(n9274), .ZN(n9424) );
  NOR2_X1 U10506 ( .A1(n9424), .A2(n9319), .ZN(n9276) );
  AOI211_X1 U10507 ( .C1(n9422), .C2(n9322), .A(n9277), .B(n9276), .ZN(n9278)
         );
  OAI21_X1 U10508 ( .B1(n9425), .B2(n9383), .A(n9278), .ZN(P1_U3268) );
  XNOR2_X1 U10509 ( .A(n9279), .B(n9285), .ZN(n9430) );
  INV_X1 U10510 ( .A(n9293), .ZN(n9281) );
  AOI21_X1 U10511 ( .B1(n9426), .B2(n9281), .A(n9280), .ZN(n9427) );
  AOI22_X1 U10512 ( .A1(n9356), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9282), .B2(
        n9343), .ZN(n9283) );
  OAI21_X1 U10513 ( .B1(n9284), .B2(n9364), .A(n9283), .ZN(n9290) );
  XNOR2_X1 U10514 ( .A(n9286), .B(n9285), .ZN(n9288) );
  AOI222_X1 U10515 ( .A1(n9355), .A2(n9288), .B1(n9314), .B2(n9380), .C1(n9287), .C2(n9372), .ZN(n9429) );
  NOR2_X1 U10516 ( .A1(n9429), .A2(n9319), .ZN(n9289) );
  AOI211_X1 U10517 ( .C1(n9427), .C2(n9322), .A(n9290), .B(n9289), .ZN(n9291)
         );
  OAI21_X1 U10518 ( .B1(n9430), .B2(n9383), .A(n9291), .ZN(P1_U3269) );
  XNOR2_X1 U10519 ( .A(n9292), .B(n9298), .ZN(n9435) );
  AOI211_X1 U10520 ( .C1(n9432), .C2(n9309), .A(n9696), .B(n9293), .ZN(n9431)
         );
  INV_X1 U10521 ( .A(n9432), .ZN(n9297) );
  INV_X1 U10522 ( .A(n9294), .ZN(n9295) );
  AOI22_X1 U10523 ( .A1(n9356), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9295), .B2(
        n9343), .ZN(n9296) );
  OAI21_X1 U10524 ( .B1(n9297), .B2(n9364), .A(n9296), .ZN(n9306) );
  OAI21_X1 U10525 ( .B1(n4321), .B2(n9299), .A(n9298), .ZN(n9301) );
  NAND2_X1 U10526 ( .A1(n9301), .A2(n9300), .ZN(n9304) );
  AOI222_X1 U10527 ( .A1(n9355), .A2(n9304), .B1(n9303), .B2(n9372), .C1(n9302), .C2(n9380), .ZN(n9434) );
  NOR2_X1 U10528 ( .A1(n9434), .A2(n9356), .ZN(n9305) );
  AOI211_X1 U10529 ( .C1(n9431), .C2(n9370), .A(n9306), .B(n9305), .ZN(n9307)
         );
  OAI21_X1 U10530 ( .B1(n9435), .B2(n9383), .A(n9307), .ZN(P1_U3270) );
  XNOR2_X1 U10531 ( .A(n9308), .B(n9316), .ZN(n9441) );
  AOI21_X1 U10532 ( .B1(n9436), .B2(n9332), .A(n4512), .ZN(n9438) );
  INV_X1 U10533 ( .A(n9310), .ZN(n9311) );
  AOI22_X1 U10534 ( .A1(n9356), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9311), .B2(
        n9343), .ZN(n9312) );
  OAI21_X1 U10535 ( .B1(n9313), .B2(n9364), .A(n9312), .ZN(n9321) );
  AND2_X1 U10536 ( .A1(n9314), .A2(n9372), .ZN(n9318) );
  AOI211_X1 U10537 ( .C1(n9316), .C2(n9315), .A(n9374), .B(n4321), .ZN(n9317)
         );
  AOI211_X1 U10538 ( .C1(n9380), .C2(n9352), .A(n9318), .B(n9317), .ZN(n9440)
         );
  NOR2_X1 U10539 ( .A1(n9440), .A2(n9319), .ZN(n9320) );
  AOI211_X1 U10540 ( .C1(n9438), .C2(n9322), .A(n9321), .B(n9320), .ZN(n9323)
         );
  OAI21_X1 U10541 ( .B1(n9441), .B2(n9383), .A(n9323), .ZN(P1_U3271) );
  XNOR2_X1 U10542 ( .A(n9325), .B(n9324), .ZN(n9446) );
  XNOR2_X1 U10543 ( .A(n9326), .B(n4696), .ZN(n9327) );
  OAI222_X1 U10544 ( .A1(n9331), .A2(n9330), .B1(n9329), .B2(n9328), .C1(n9327), .C2(n9374), .ZN(n9442) );
  INV_X1 U10545 ( .A(n9341), .ZN(n9333) );
  AOI211_X1 U10546 ( .C1(n9444), .C2(n9333), .A(n9696), .B(n4513), .ZN(n9443)
         );
  NAND2_X1 U10547 ( .A1(n9443), .A2(n9370), .ZN(n9336) );
  AOI22_X1 U10548 ( .A1(n9356), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9334), .B2(
        n9343), .ZN(n9335) );
  OAI211_X1 U10549 ( .C1(n9337), .C2(n9364), .A(n9336), .B(n9335), .ZN(n9338)
         );
  AOI21_X1 U10550 ( .B1(n9442), .B2(n9367), .A(n9338), .ZN(n9339) );
  OAI21_X1 U10551 ( .B1(n9446), .B2(n9383), .A(n9339), .ZN(P1_U3272) );
  XNOR2_X1 U10552 ( .A(n9340), .B(n9348), .ZN(n9451) );
  INV_X1 U10553 ( .A(n9362), .ZN(n9342) );
  AOI211_X1 U10554 ( .C1(n9448), .C2(n9342), .A(n9696), .B(n9341), .ZN(n9447)
         );
  AOI22_X1 U10555 ( .A1(n9356), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9344), .B2(
        n9343), .ZN(n9345) );
  OAI21_X1 U10556 ( .B1(n9346), .B2(n9364), .A(n9345), .ZN(n9358) );
  INV_X1 U10557 ( .A(n9347), .ZN(n9373) );
  OAI21_X1 U10558 ( .B1(n9373), .B2(n9349), .A(n9348), .ZN(n9351) );
  NAND2_X1 U10559 ( .A1(n9351), .A2(n9350), .ZN(n9354) );
  AOI222_X1 U10560 ( .A1(n9355), .A2(n9354), .B1(n9353), .B2(n9380), .C1(n9352), .C2(n9372), .ZN(n9450) );
  NOR2_X1 U10561 ( .A1(n9450), .A2(n9356), .ZN(n9357) );
  AOI211_X1 U10562 ( .C1(n9447), .C2(n9370), .A(n9358), .B(n9357), .ZN(n9359)
         );
  OAI21_X1 U10563 ( .B1(n9451), .B2(n9383), .A(n9359), .ZN(P1_U3273) );
  XNOR2_X1 U10564 ( .A(n9361), .B(n9360), .ZN(n9456) );
  AOI211_X1 U10565 ( .C1(n9453), .C2(n9363), .A(n9696), .B(n9362), .ZN(n9452)
         );
  NOR2_X1 U10566 ( .A1(n4517), .A2(n9364), .ZN(n9369) );
  OAI22_X1 U10567 ( .A1(n9367), .A2(n9159), .B1(n9366), .B2(n9365), .ZN(n9368)
         );
  AOI211_X1 U10568 ( .C1(n9452), .C2(n9370), .A(n9369), .B(n9368), .ZN(n9382)
         );
  AND2_X1 U10569 ( .A1(n9372), .A2(n9371), .ZN(n9378) );
  AOI211_X1 U10570 ( .C1(n9376), .C2(n9375), .A(n9374), .B(n9373), .ZN(n9377)
         );
  AOI211_X1 U10571 ( .C1(n9380), .C2(n9379), .A(n9378), .B(n9377), .ZN(n9455)
         );
  OR2_X1 U10572 ( .A1(n9455), .A2(n9356), .ZN(n9381) );
  OAI211_X1 U10573 ( .C1(n9456), .C2(n9383), .A(n9382), .B(n9381), .ZN(
        P1_U3274) );
  NAND2_X1 U10574 ( .A1(n9384), .A2(n9437), .ZN(n9385) );
  OAI211_X1 U10575 ( .C1(n9386), .C2(n9710), .A(n9385), .B(n9389), .ZN(n9469)
         );
  MUX2_X1 U10576 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9469), .S(n9561), .Z(
        P1_U3554) );
  NAND2_X1 U10577 ( .A1(n9387), .A2(n9465), .ZN(n9388) );
  OAI211_X1 U10578 ( .C1(n9390), .C2(n9696), .A(n9389), .B(n9388), .ZN(n9470)
         );
  MUX2_X1 U10579 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9470), .S(n9561), .Z(
        P1_U3553) );
  MUX2_X1 U10580 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9471), .S(n9561), .Z(
        P1_U3552) );
  AOI22_X1 U10581 ( .A1(n9397), .A2(n9437), .B1(n9465), .B2(n9396), .ZN(n9398)
         );
  OAI211_X1 U10582 ( .C1(n9400), .C2(n9468), .A(n9399), .B(n9398), .ZN(n9472)
         );
  MUX2_X1 U10583 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9472), .S(n9561), .Z(
        P1_U3551) );
  AOI211_X1 U10584 ( .C1(n9465), .C2(n9403), .A(n9402), .B(n9401), .ZN(n9404)
         );
  OAI21_X1 U10585 ( .B1(n9405), .B2(n9468), .A(n9404), .ZN(n9473) );
  MUX2_X1 U10586 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9473), .S(n9561), .Z(
        P1_U3550) );
  AOI22_X1 U10587 ( .A1(n9407), .A2(n9437), .B1(n9465), .B2(n9406), .ZN(n9408)
         );
  OAI211_X1 U10588 ( .C1(n9410), .C2(n9468), .A(n9409), .B(n9408), .ZN(n9474)
         );
  MUX2_X1 U10589 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9474), .S(n9561), .Z(
        P1_U3549) );
  AOI22_X1 U10590 ( .A1(n9412), .A2(n9437), .B1(n9465), .B2(n9411), .ZN(n9413)
         );
  OAI211_X1 U10591 ( .C1(n9415), .C2(n9468), .A(n9414), .B(n9413), .ZN(n9475)
         );
  MUX2_X1 U10592 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9475), .S(n9561), .Z(
        P1_U3548) );
  AOI211_X1 U10593 ( .C1(n9465), .C2(n9418), .A(n9417), .B(n9416), .ZN(n9419)
         );
  OAI21_X1 U10594 ( .B1(n9420), .B2(n9468), .A(n9419), .ZN(n9476) );
  MUX2_X1 U10595 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9476), .S(n9561), .Z(
        P1_U3547) );
  AOI22_X1 U10596 ( .A1(n9422), .A2(n9437), .B1(n9465), .B2(n9421), .ZN(n9423)
         );
  OAI211_X1 U10597 ( .C1(n9425), .C2(n9468), .A(n9424), .B(n9423), .ZN(n9477)
         );
  MUX2_X1 U10598 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9477), .S(n9561), .Z(
        P1_U3546) );
  AOI22_X1 U10599 ( .A1(n9427), .A2(n9437), .B1(n9465), .B2(n9426), .ZN(n9428)
         );
  OAI211_X1 U10600 ( .C1(n9430), .C2(n9468), .A(n9429), .B(n9428), .ZN(n9478)
         );
  MUX2_X1 U10601 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9478), .S(n9561), .Z(
        P1_U3545) );
  AOI21_X1 U10602 ( .B1(n9465), .B2(n9432), .A(n9431), .ZN(n9433) );
  OAI211_X1 U10603 ( .C1(n9435), .C2(n9468), .A(n9434), .B(n9433), .ZN(n9479)
         );
  MUX2_X1 U10604 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9479), .S(n9561), .Z(
        P1_U3544) );
  AOI22_X1 U10605 ( .A1(n9438), .A2(n9437), .B1(n9465), .B2(n9436), .ZN(n9439)
         );
  OAI211_X1 U10606 ( .C1(n9441), .C2(n9468), .A(n9440), .B(n9439), .ZN(n9480)
         );
  MUX2_X1 U10607 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9480), .S(n9561), .Z(
        P1_U3543) );
  AOI211_X1 U10608 ( .C1(n9465), .C2(n9444), .A(n9443), .B(n9442), .ZN(n9445)
         );
  OAI21_X1 U10609 ( .B1(n9446), .B2(n9468), .A(n9445), .ZN(n9481) );
  MUX2_X1 U10610 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9481), .S(n9561), .Z(
        P1_U3542) );
  AOI21_X1 U10611 ( .B1(n9465), .B2(n9448), .A(n9447), .ZN(n9449) );
  OAI211_X1 U10612 ( .C1(n9451), .C2(n9468), .A(n9450), .B(n9449), .ZN(n9482)
         );
  MUX2_X1 U10613 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9482), .S(n9561), .Z(
        P1_U3541) );
  AOI21_X1 U10614 ( .B1(n9465), .B2(n9453), .A(n9452), .ZN(n9454) );
  OAI211_X1 U10615 ( .C1(n9456), .C2(n9468), .A(n9455), .B(n9454), .ZN(n9483)
         );
  MUX2_X1 U10616 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9483), .S(n9561), .Z(
        P1_U3540) );
  AOI211_X1 U10617 ( .C1(n9465), .C2(n9459), .A(n9458), .B(n9457), .ZN(n9460)
         );
  OAI21_X1 U10618 ( .B1(n9461), .B2(n9468), .A(n9460), .ZN(n9484) );
  MUX2_X1 U10619 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9484), .S(n9561), .Z(
        P1_U3539) );
  AOI211_X1 U10620 ( .C1(n9465), .C2(n9464), .A(n9463), .B(n9462), .ZN(n9466)
         );
  OAI21_X1 U10621 ( .B1(n9468), .B2(n9467), .A(n9466), .ZN(n9485) );
  MUX2_X1 U10622 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9485), .S(n9561), .Z(
        P1_U3535) );
  MUX2_X1 U10623 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9469), .S(n9719), .Z(
        P1_U3522) );
  MUX2_X1 U10624 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9470), .S(n9719), .Z(
        P1_U3521) );
  MUX2_X1 U10625 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9472), .S(n9719), .Z(
        P1_U3519) );
  MUX2_X1 U10626 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9473), .S(n9719), .Z(
        P1_U3518) );
  MUX2_X1 U10627 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9474), .S(n9719), .Z(
        P1_U3517) );
  MUX2_X1 U10628 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9475), .S(n9719), .Z(
        P1_U3516) );
  MUX2_X1 U10629 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9476), .S(n9719), .Z(
        P1_U3515) );
  MUX2_X1 U10630 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9477), .S(n9719), .Z(
        P1_U3514) );
  MUX2_X1 U10631 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9478), .S(n9719), .Z(
        P1_U3513) );
  MUX2_X1 U10632 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9479), .S(n9719), .Z(
        P1_U3512) );
  MUX2_X1 U10633 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9480), .S(n9719), .Z(
        P1_U3511) );
  MUX2_X1 U10634 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9481), .S(n9719), .Z(
        P1_U3510) );
  MUX2_X1 U10635 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9482), .S(n9719), .Z(
        P1_U3508) );
  MUX2_X1 U10636 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9483), .S(n9719), .Z(
        P1_U3505) );
  MUX2_X1 U10637 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9484), .S(n9719), .Z(
        P1_U3502) );
  MUX2_X1 U10638 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9485), .S(n9719), .Z(
        P1_U3490) );
  NOR4_X1 U10639 ( .A1(n5698), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9486), .ZN(n9487) );
  AOI21_X1 U10640 ( .B1(n9488), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9487), .ZN(
        n9489) );
  OAI21_X1 U10641 ( .B1(n9490), .B2(n9493), .A(n9489), .ZN(P1_U3322) );
  OAI222_X1 U10642 ( .A1(n9495), .A2(n9494), .B1(n9493), .B2(n9492), .C1(
        P1_U3084), .C2(n9491), .ZN(P1_U3323) );
  MUX2_X1 U10643 ( .A(n9496), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10644 ( .A1(n9729), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9508) );
  AOI211_X1 U10645 ( .C1(n9499), .C2(n9498), .A(n9497), .B(n9732), .ZN(n9500)
         );
  AOI21_X1 U10646 ( .B1(n9514), .B2(n9501), .A(n9500), .ZN(n9507) );
  INV_X1 U10647 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9502) );
  NOR2_X1 U10648 ( .A1(n9502), .A2(n5064), .ZN(n9505) );
  OAI211_X1 U10649 ( .C1(n9505), .C2(n9504), .A(n9728), .B(n9503), .ZN(n9506)
         );
  NAND3_X1 U10650 ( .A1(n9508), .A2(n9507), .A3(n9506), .ZN(P2_U3246) );
  AOI22_X1 U10651 ( .A1(n9729), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9520) );
  AOI211_X1 U10652 ( .C1(n9511), .C2(n9510), .A(n9509), .B(n9732), .ZN(n9512)
         );
  AOI21_X1 U10653 ( .B1(n9514), .B2(n9513), .A(n9512), .ZN(n9519) );
  OAI211_X1 U10654 ( .C1(n9517), .C2(n9516), .A(n9728), .B(n9515), .ZN(n9518)
         );
  NAND3_X1 U10655 ( .A1(n9520), .A2(n9519), .A3(n9518), .ZN(P2_U3247) );
  INV_X1 U10656 ( .A(n9521), .ZN(n9524) );
  NOR2_X1 U10657 ( .A1(n9522), .A2(n9810), .ZN(n9523) );
  INV_X1 U10658 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9526) );
  AOI22_X1 U10659 ( .A1(n9830), .A2(n9533), .B1(n9526), .B2(n9828), .ZN(
        P2_U3550) );
  OAI22_X1 U10660 ( .A1(n9528), .A2(n9810), .B1(n9527), .B2(n9808), .ZN(n9529)
         );
  AOI211_X1 U10661 ( .C1(n9531), .C2(n9800), .A(n9530), .B(n9529), .ZN(n9534)
         );
  AOI22_X1 U10662 ( .A1(n9830), .A2(n9534), .B1(n8645), .B2(n9828), .ZN(
        P2_U3534) );
  INV_X1 U10663 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9532) );
  AOI22_X1 U10664 ( .A1(n9817), .A2(n9533), .B1(n9532), .B2(n9816), .ZN(
        P2_U3518) );
  INV_X1 U10665 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U10666 ( .A1(n9817), .A2(n9534), .B1(n9971), .B2(n9816), .ZN(
        P2_U3493) );
  INV_X1 U10667 ( .A(n9535), .ZN(n9713) );
  INV_X1 U10668 ( .A(n9536), .ZN(n9541) );
  OAI22_X1 U10669 ( .A1(n9538), .A2(n9696), .B1(n9537), .B2(n9710), .ZN(n9540)
         );
  AOI211_X1 U10670 ( .C1(n9713), .C2(n9541), .A(n9540), .B(n9539), .ZN(n9563)
         );
  AOI22_X1 U10671 ( .A1(n9561), .A2(n9563), .B1(n9542), .B2(n9724), .ZN(
        P1_U3538) );
  OAI21_X1 U10672 ( .B1(n9544), .B2(n9710), .A(n9543), .ZN(n9545) );
  AOI211_X1 U10673 ( .C1(n9547), .C2(n9706), .A(n9546), .B(n9545), .ZN(n9565)
         );
  AOI22_X1 U10674 ( .A1(n9561), .A2(n9565), .B1(n9548), .B2(n9724), .ZN(
        P1_U3537) );
  OAI21_X1 U10675 ( .B1(n7159), .B2(n9710), .A(n9549), .ZN(n9550) );
  AOI21_X1 U10676 ( .B1(n9551), .B2(n9713), .A(n9550), .ZN(n9552) );
  AND2_X1 U10677 ( .A1(n9553), .A2(n9552), .ZN(n9567) );
  AOI22_X1 U10678 ( .A1(n9561), .A2(n9567), .B1(n6597), .B2(n9724), .ZN(
        P1_U3536) );
  OAI22_X1 U10679 ( .A1(n9555), .A2(n9696), .B1(n9554), .B2(n9710), .ZN(n9556)
         );
  AOI21_X1 U10680 ( .B1(n9557), .B2(n9713), .A(n9556), .ZN(n9558) );
  AND2_X1 U10681 ( .A1(n9559), .A2(n9558), .ZN(n9568) );
  AOI22_X1 U10682 ( .A1(n9561), .A2(n9568), .B1(n9560), .B2(n9724), .ZN(
        P1_U3534) );
  INV_X1 U10683 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9562) );
  AOI22_X1 U10684 ( .A1(n9719), .A2(n9563), .B1(n9562), .B2(n9717), .ZN(
        P1_U3499) );
  INV_X1 U10685 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9564) );
  AOI22_X1 U10686 ( .A1(n9719), .A2(n9565), .B1(n9564), .B2(n9717), .ZN(
        P1_U3496) );
  INV_X1 U10687 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9566) );
  AOI22_X1 U10688 ( .A1(n9719), .A2(n9567), .B1(n9566), .B2(n9717), .ZN(
        P1_U3493) );
  INV_X1 U10689 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U10690 ( .A1(n9719), .A2(n9568), .B1(n9889), .B2(n9717), .ZN(
        P1_U3487) );
  INV_X1 U10691 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10017) );
  XOR2_X1 U10692 ( .A(n10017), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U10693 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U10694 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9571) );
  AOI211_X1 U10695 ( .C1(n9571), .C2(n9570), .A(n9569), .B(n9579), .ZN(n9572)
         );
  AOI21_X1 U10696 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(P1_U3084), .A(n9572), 
        .ZN(n9578) );
  AOI22_X1 U10697 ( .A1(n9678), .A2(n5940), .B1(n9685), .B2(
        P1_ADDR_REG_1__SCAN_IN), .ZN(n9577) );
  AND2_X1 U10698 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9575) );
  OAI211_X1 U10699 ( .C1(n9575), .C2(n9574), .A(n9676), .B(n9573), .ZN(n9576)
         );
  NAND3_X1 U10700 ( .A1(n9578), .A2(n9577), .A3(n9576), .ZN(P1_U3242) );
  AOI211_X1 U10701 ( .C1(n9582), .C2(n9581), .A(n9580), .B(n9579), .ZN(n9594)
         );
  AOI21_X1 U10702 ( .B1(n9583), .B2(n9585), .A(n9119), .ZN(n9584) );
  OAI21_X1 U10703 ( .B1(n9586), .B2(n9585), .A(n9584), .ZN(n9611) );
  OAI211_X1 U10704 ( .C1(n9589), .C2(n9588), .A(n9676), .B(n9587), .ZN(n9590)
         );
  OAI211_X1 U10705 ( .C1(n9592), .C2(n9591), .A(n9611), .B(n9590), .ZN(n9593)
         );
  AOI211_X1 U10706 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(P1_U3084), .A(n9594), 
        .B(n9593), .ZN(n9595) );
  OAI21_X1 U10707 ( .B1(n9671), .B2(n9596), .A(n9595), .ZN(P1_U3243) );
  AOI21_X1 U10708 ( .B1(n9599), .B2(n9598), .A(n9597), .ZN(n9600) );
  INV_X1 U10709 ( .A(n9600), .ZN(n9601) );
  NAND2_X1 U10710 ( .A1(n9676), .A2(n9601), .ZN(n9610) );
  NAND2_X1 U10711 ( .A1(n9678), .A2(n9602), .ZN(n9609) );
  OAI21_X1 U10712 ( .B1(n9605), .B2(n9604), .A(n9603), .ZN(n9607) );
  AOI21_X1 U10713 ( .B1(n9686), .B2(n9607), .A(n9606), .ZN(n9608) );
  AND3_X1 U10714 ( .A1(n9610), .A2(n9609), .A3(n9608), .ZN(n9612) );
  OAI211_X1 U10715 ( .C1(n9613), .C2(n9671), .A(n9612), .B(n9611), .ZN(
        P1_U3245) );
  OAI21_X1 U10716 ( .B1(n5736), .B2(n9614), .A(n9628), .ZN(n9622) );
  AOI21_X1 U10717 ( .B1(n9617), .B2(n9616), .A(n9615), .ZN(n9618) );
  NAND2_X1 U10718 ( .A1(n9686), .A2(n9618), .ZN(n9621) );
  INV_X1 U10719 ( .A(n9619), .ZN(n9620) );
  OAI211_X1 U10720 ( .C1(n9623), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9624)
         );
  INV_X1 U10721 ( .A(n9624), .ZN(n9630) );
  INV_X1 U10722 ( .A(n9625), .ZN(n9626) );
  INV_X1 U10723 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10034) );
  NAND2_X1 U10724 ( .A1(n9626), .A2(n10034), .ZN(n9627) );
  OAI211_X1 U10725 ( .C1(n9628), .C2(n9627), .A(n9676), .B(n9640), .ZN(n9629)
         );
  OAI211_X1 U10726 ( .C1(n9631), .C2(n9671), .A(n9630), .B(n9629), .ZN(
        P1_U3249) );
  OAI21_X1 U10727 ( .B1(n9634), .B2(n9633), .A(n9632), .ZN(n9636) );
  AOI21_X1 U10728 ( .B1(n9636), .B2(n9686), .A(n9635), .ZN(n9644) );
  AOI211_X1 U10729 ( .C1(n9640), .C2(n9639), .A(n9638), .B(n9637), .ZN(n9641)
         );
  AOI21_X1 U10730 ( .B1(n9678), .B2(n9642), .A(n9641), .ZN(n9643) );
  OAI211_X1 U10731 ( .C1(n9671), .C2(n10059), .A(n9644), .B(n9643), .ZN(
        P1_U3250) );
  INV_X1 U10732 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9657) );
  AOI21_X1 U10733 ( .B1(n9678), .B2(n9646), .A(n9645), .ZN(n9656) );
  OAI21_X1 U10734 ( .B1(n9649), .B2(n9648), .A(n9647), .ZN(n9654) );
  OAI21_X1 U10735 ( .B1(n9652), .B2(n9651), .A(n9650), .ZN(n9653) );
  AOI22_X1 U10736 ( .A1(n9654), .A2(n9686), .B1(n9653), .B2(n9676), .ZN(n9655)
         );
  OAI211_X1 U10737 ( .C1(n9671), .C2(n9657), .A(n9656), .B(n9655), .ZN(
        P1_U3252) );
  INV_X1 U10738 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9670) );
  AOI21_X1 U10739 ( .B1(n9678), .B2(n9659), .A(n9658), .ZN(n9669) );
  OAI21_X1 U10740 ( .B1(n9662), .B2(n9661), .A(n9660), .ZN(n9667) );
  OAI21_X1 U10741 ( .B1(n9665), .B2(n9664), .A(n9663), .ZN(n9666) );
  AOI22_X1 U10742 ( .A1(n9667), .A2(n9676), .B1(n9686), .B2(n9666), .ZN(n9668)
         );
  OAI211_X1 U10743 ( .C1(n9671), .C2(n9670), .A(n9669), .B(n9668), .ZN(
        P1_U3255) );
  AOI21_X1 U10744 ( .B1(n9674), .B2(n9673), .A(n9672), .ZN(n9675) );
  NAND2_X1 U10745 ( .A1(n9676), .A2(n9675), .ZN(n9681) );
  NAND2_X1 U10746 ( .A1(n9678), .A2(n9677), .ZN(n9680) );
  AND3_X1 U10747 ( .A1(n9681), .A2(n9680), .A3(n9679), .ZN(n9689) );
  OAI21_X1 U10748 ( .B1(n9684), .B2(n9683), .A(n9682), .ZN(n9687) );
  AOI22_X1 U10749 ( .A1(n9687), .A2(n9686), .B1(n9685), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U10750 ( .A1(n9689), .A2(n9688), .ZN(P1_U3259) );
  INV_X1 U10751 ( .A(n9690), .ZN(n9691) );
  AND2_X1 U10752 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9860), .ZN(P1_U3292) );
  AND2_X1 U10753 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9860), .ZN(P1_U3293) );
  AND2_X1 U10754 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9860), .ZN(P1_U3294) );
  AND2_X1 U10755 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9860), .ZN(P1_U3295) );
  AND2_X1 U10756 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9860), .ZN(P1_U3296) );
  INV_X1 U10757 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10013) );
  NOR2_X1 U10758 ( .A1(n9692), .A2(n10013), .ZN(P1_U3297) );
  AND2_X1 U10759 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9860), .ZN(P1_U3298) );
  AND2_X1 U10760 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9860), .ZN(P1_U3299) );
  AND2_X1 U10761 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9860), .ZN(P1_U3300) );
  INV_X1 U10762 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9974) );
  NOR2_X1 U10763 ( .A1(n9692), .A2(n9974), .ZN(P1_U3301) );
  AND2_X1 U10764 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9860), .ZN(P1_U3302) );
  AND2_X1 U10765 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9860), .ZN(P1_U3303) );
  AND2_X1 U10766 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9860), .ZN(P1_U3304) );
  AND2_X1 U10767 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9860), .ZN(P1_U3305) );
  AND2_X1 U10768 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9860), .ZN(P1_U3306) );
  AND2_X1 U10769 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9860), .ZN(P1_U3307) );
  AND2_X1 U10770 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9860), .ZN(P1_U3308) );
  AND2_X1 U10771 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9860), .ZN(P1_U3310) );
  AND2_X1 U10772 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9860), .ZN(P1_U3311) );
  AND2_X1 U10773 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9860), .ZN(P1_U3312) );
  AND2_X1 U10774 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9860), .ZN(P1_U3313) );
  AND2_X1 U10775 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9860), .ZN(P1_U3314) );
  AND2_X1 U10776 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9860), .ZN(P1_U3315) );
  AND2_X1 U10777 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9860), .ZN(P1_U3316) );
  AND2_X1 U10778 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9860), .ZN(P1_U3317) );
  AND2_X1 U10779 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9860), .ZN(P1_U3318) );
  AND2_X1 U10780 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9860), .ZN(P1_U3319) );
  INV_X1 U10781 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10032) );
  NOR2_X1 U10782 ( .A1(n9692), .A2(n10032), .ZN(P1_U3320) );
  AND2_X1 U10783 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9860), .ZN(P1_U3321) );
  OAI21_X1 U10784 ( .B1(n9694), .B2(n9990), .A(n9693), .ZN(P1_U3440) );
  OAI22_X1 U10785 ( .A1(n9697), .A2(n9696), .B1(n9695), .B2(n9710), .ZN(n9699)
         );
  AOI211_X1 U10786 ( .C1(n9713), .C2(n9700), .A(n9699), .B(n9698), .ZN(n9721)
         );
  INV_X1 U10787 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9701) );
  AOI22_X1 U10788 ( .A1(n9719), .A2(n9721), .B1(n9701), .B2(n9717), .ZN(
        P1_U3463) );
  OAI21_X1 U10789 ( .B1(n9703), .B2(n9710), .A(n9702), .ZN(n9704) );
  AOI211_X1 U10790 ( .C1(n9707), .C2(n9706), .A(n9705), .B(n9704), .ZN(n9723)
         );
  INV_X1 U10791 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9708) );
  AOI22_X1 U10792 ( .A1(n9719), .A2(n9723), .B1(n9708), .B2(n9717), .ZN(
        P1_U3469) );
  OAI21_X1 U10793 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9712) );
  AOI21_X1 U10794 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(n9715) );
  AND2_X1 U10795 ( .A1(n9716), .A2(n9715), .ZN(n9726) );
  INV_X1 U10796 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9718) );
  AOI22_X1 U10797 ( .A1(n9719), .A2(n9726), .B1(n9718), .B2(n9717), .ZN(
        P1_U3481) );
  INV_X1 U10798 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9720) );
  AOI22_X1 U10799 ( .A1(n9561), .A2(n9721), .B1(n9720), .B2(n9724), .ZN(
        P1_U3526) );
  INV_X1 U10800 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9722) );
  AOI22_X1 U10801 ( .A1(n9561), .A2(n9723), .B1(n9722), .B2(n9724), .ZN(
        P1_U3528) );
  INV_X1 U10802 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9725) );
  AOI22_X1 U10803 ( .A1(n9561), .A2(n9726), .B1(n9725), .B2(n9724), .ZN(
        P1_U3532) );
  AOI22_X1 U10804 ( .A1(n9728), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n9727), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9737) );
  AOI22_X1 U10805 ( .A1(n9729), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9736) );
  NOR2_X1 U10806 ( .A1(n9730), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9734) );
  OAI21_X1 U10807 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n9732), .A(n9731), .ZN(
        n9733) );
  OAI21_X1 U10808 ( .B1(n9734), .B2(n9733), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9735) );
  OAI211_X1 U10809 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9737), .A(n9736), .B(
        n9735), .ZN(P2_U3245) );
  INV_X1 U10810 ( .A(n9738), .ZN(n9747) );
  OAI22_X1 U10811 ( .A1(n9742), .A2(n9741), .B1(n9740), .B2(n9739), .ZN(n9743)
         );
  AOI21_X1 U10812 ( .B1(n9745), .B2(n9744), .A(n9743), .ZN(n9746) );
  OAI211_X1 U10813 ( .C1(n9749), .C2(n9748), .A(n9747), .B(n9746), .ZN(n9750)
         );
  INV_X1 U10814 ( .A(n9750), .ZN(n9751) );
  AOI22_X1 U10815 ( .A1(n9752), .A2(n5783), .B1(n9751), .B2(n8826), .ZN(
        P2_U3291) );
  AND2_X1 U10816 ( .A1(n9758), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3297) );
  AND2_X1 U10817 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9758), .ZN(P2_U3298) );
  AND2_X1 U10818 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9758), .ZN(P2_U3299) );
  AND2_X1 U10819 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9758), .ZN(P2_U3300) );
  AND2_X1 U10820 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9758), .ZN(P2_U3301) );
  AND2_X1 U10821 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9758), .ZN(P2_U3302) );
  INV_X1 U10822 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9898) );
  NOR2_X1 U10823 ( .A1(n9755), .A2(n9898), .ZN(P2_U3303) );
  AND2_X1 U10824 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9758), .ZN(P2_U3304) );
  AND2_X1 U10825 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9758), .ZN(P2_U3305) );
  AND2_X1 U10826 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9758), .ZN(P2_U3306) );
  AND2_X1 U10827 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9758), .ZN(P2_U3307) );
  INV_X1 U10828 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9897) );
  NOR2_X1 U10829 ( .A1(n9755), .A2(n9897), .ZN(P2_U3308) );
  AND2_X1 U10830 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9758), .ZN(P2_U3309) );
  INV_X1 U10831 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10002) );
  NOR2_X1 U10832 ( .A1(n9755), .A2(n10002), .ZN(P2_U3310) );
  AND2_X1 U10833 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9758), .ZN(P2_U3311) );
  AND2_X1 U10834 ( .A1(n9758), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3312) );
  AND2_X1 U10835 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9758), .ZN(P2_U3313) );
  INV_X1 U10836 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9862) );
  NOR2_X1 U10837 ( .A1(n9755), .A2(n9862), .ZN(P2_U3314) );
  AND2_X1 U10838 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9758), .ZN(P2_U3315) );
  AND2_X1 U10839 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9758), .ZN(P2_U3316) );
  INV_X1 U10840 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10027) );
  NOR2_X1 U10841 ( .A1(n9755), .A2(n10027), .ZN(P2_U3317) );
  AND2_X1 U10842 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9758), .ZN(P2_U3318) );
  AND2_X1 U10843 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9758), .ZN(P2_U3319) );
  AND2_X1 U10844 ( .A1(n9758), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3320) );
  AND2_X1 U10845 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9758), .ZN(P2_U3321) );
  AND2_X1 U10846 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9758), .ZN(P2_U3322) );
  AND2_X1 U10847 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9758), .ZN(P2_U3323) );
  AND2_X1 U10848 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9758), .ZN(P2_U3324) );
  AND2_X1 U10849 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9758), .ZN(P2_U3325) );
  AND2_X1 U10850 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9758), .ZN(P2_U3326) );
  AOI22_X1 U10851 ( .A1(n9757), .A2(n9760), .B1(n9756), .B2(n9758), .ZN(
        P2_U3437) );
  AOI22_X1 U10852 ( .A1(n9761), .A2(n9760), .B1(n9759), .B2(n9758), .ZN(
        P2_U3438) );
  AOI22_X1 U10853 ( .A1(n9764), .A2(n9800), .B1(n9763), .B2(n9762), .ZN(n9765)
         );
  AND2_X1 U10854 ( .A1(n9766), .A2(n9765), .ZN(n9819) );
  AOI22_X1 U10855 ( .A1(n9817), .A2(n9819), .B1(n5063), .B2(n9816), .ZN(
        P2_U3451) );
  OAI211_X1 U10856 ( .C1(n6205), .C2(n9808), .A(n9768), .B(n9767), .ZN(n9769)
         );
  AOI21_X1 U10857 ( .B1(n9800), .B2(n9770), .A(n9769), .ZN(n9820) );
  AOI22_X1 U10858 ( .A1(n9817), .A2(n9820), .B1(n5050), .B2(n9816), .ZN(
        P2_U3454) );
  AOI22_X1 U10859 ( .A1(n9773), .A2(n9786), .B1(n9772), .B2(n9771), .ZN(n9774)
         );
  NAND2_X1 U10860 ( .A1(n9775), .A2(n9774), .ZN(n9776) );
  AOI21_X1 U10861 ( .B1(n9800), .B2(n9777), .A(n9776), .ZN(n9821) );
  AOI22_X1 U10862 ( .A1(n9817), .A2(n9821), .B1(n5073), .B2(n9816), .ZN(
        P2_U3457) );
  INV_X1 U10863 ( .A(n9778), .ZN(n9815) );
  INV_X1 U10864 ( .A(n9779), .ZN(n9784) );
  OAI22_X1 U10865 ( .A1(n9781), .A2(n9810), .B1(n9780), .B2(n9808), .ZN(n9783)
         );
  AOI211_X1 U10866 ( .C1(n9815), .C2(n9784), .A(n9783), .B(n9782), .ZN(n9823)
         );
  AOI22_X1 U10867 ( .A1(n9817), .A2(n9823), .B1(n5087), .B2(n9816), .ZN(
        P2_U3460) );
  AOI22_X1 U10868 ( .A1(n9787), .A2(n9786), .B1(n9772), .B2(n9785), .ZN(n9788)
         );
  OAI211_X1 U10869 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9788), .ZN(n9792)
         );
  INV_X1 U10870 ( .A(n9792), .ZN(n9824) );
  AOI22_X1 U10871 ( .A1(n9817), .A2(n9824), .B1(n5103), .B2(n9816), .ZN(
        P2_U3463) );
  INV_X1 U10872 ( .A(n9793), .ZN(n9799) );
  OAI22_X1 U10873 ( .A1(n9795), .A2(n9810), .B1(n9794), .B2(n9808), .ZN(n9798)
         );
  INV_X1 U10874 ( .A(n9796), .ZN(n9797) );
  AOI211_X1 U10875 ( .C1(n9800), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9826)
         );
  AOI22_X1 U10876 ( .A1(n9817), .A2(n9826), .B1(n5129), .B2(n9816), .ZN(
        P2_U3469) );
  INV_X1 U10877 ( .A(n9801), .ZN(n9806) );
  OAI22_X1 U10878 ( .A1(n9803), .A2(n9810), .B1(n4549), .B2(n9808), .ZN(n9805)
         );
  AOI211_X1 U10879 ( .C1(n9815), .C2(n9806), .A(n9805), .B(n9804), .ZN(n9827)
         );
  AOI22_X1 U10880 ( .A1(n9817), .A2(n9827), .B1(n5172), .B2(n9816), .ZN(
        P2_U3475) );
  INV_X1 U10881 ( .A(n9807), .ZN(n9814) );
  INV_X1 U10882 ( .A(n5207), .ZN(n9809) );
  OAI22_X1 U10883 ( .A1(n9811), .A2(n9810), .B1(n9809), .B2(n9808), .ZN(n9813)
         );
  AOI211_X1 U10884 ( .C1(n9815), .C2(n9814), .A(n9813), .B(n9812), .ZN(n9829)
         );
  AOI22_X1 U10885 ( .A1(n9817), .A2(n9829), .B1(n5202), .B2(n9816), .ZN(
        P2_U3481) );
  INV_X1 U10886 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9818) );
  AOI22_X1 U10887 ( .A1(n9830), .A2(n9819), .B1(n9818), .B2(n9828), .ZN(
        P2_U3520) );
  AOI22_X1 U10888 ( .A1(n9830), .A2(n9820), .B1(n5751), .B2(n9828), .ZN(
        P2_U3521) );
  AOI22_X1 U10889 ( .A1(n9830), .A2(n9821), .B1(n5752), .B2(n9828), .ZN(
        P2_U3522) );
  INV_X1 U10890 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U10891 ( .A1(n9830), .A2(n9823), .B1(n9822), .B2(n9828), .ZN(
        P2_U3523) );
  AOI22_X1 U10892 ( .A1(n9830), .A2(n9824), .B1(n5754), .B2(n9828), .ZN(
        P2_U3524) );
  INV_X1 U10893 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9825) );
  AOI22_X1 U10894 ( .A1(n9830), .A2(n9826), .B1(n9825), .B2(n9828), .ZN(
        P2_U3526) );
  AOI22_X1 U10895 ( .A1(n9830), .A2(n9827), .B1(n6185), .B2(n9828), .ZN(
        P2_U3528) );
  AOI22_X1 U10896 ( .A1(n9830), .A2(n9829), .B1(n6578), .B2(n9828), .ZN(
        P2_U3530) );
  INV_X1 U10897 ( .A(n9831), .ZN(n9832) );
  NAND2_X1 U10898 ( .A1(n9833), .A2(n9832), .ZN(n9834) );
  XOR2_X1 U10899 ( .A(n9835), .B(n9834), .Z(ADD_1071_U5) );
  XOR2_X1 U10900 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10901 ( .B1(n9838), .B2(n9837), .A(n9836), .ZN(ADD_1071_U56) );
  OAI21_X1 U10902 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(ADD_1071_U57) );
  OAI21_X1 U10903 ( .B1(n9844), .B2(n9843), .A(n9842), .ZN(ADD_1071_U58) );
  OAI21_X1 U10904 ( .B1(n9847), .B2(n9846), .A(n9845), .ZN(ADD_1071_U59) );
  OAI21_X1 U10905 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(ADD_1071_U60) );
  OAI21_X1 U10906 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(ADD_1071_U61) );
  AOI21_X1 U10907 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(ADD_1071_U62) );
  AOI21_X1 U10908 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(ADD_1071_U63) );
  NAND2_X1 U10909 ( .A1(n9860), .A2(P1_D_REG_14__SCAN_IN), .ZN(n10048) );
  AOI22_X1 U10910 ( .A1(n5866), .A2(keyinput80), .B1(keyinput67), .B2(n9862), 
        .ZN(n9861) );
  OAI221_X1 U10911 ( .B1(n5866), .B2(keyinput80), .C1(n9862), .C2(keyinput67), 
        .A(n9861), .ZN(n9871) );
  AOI22_X1 U10912 ( .A1(n5028), .A2(keyinput83), .B1(keyinput103), .B2(n9971), 
        .ZN(n9863) );
  OAI221_X1 U10913 ( .B1(n5028), .B2(keyinput83), .C1(n9971), .C2(keyinput103), 
        .A(n9863), .ZN(n9870) );
  AOI22_X1 U10914 ( .A1(n10034), .A2(keyinput101), .B1(n9865), .B2(keyinput81), 
        .ZN(n9864) );
  OAI221_X1 U10915 ( .B1(n10034), .B2(keyinput101), .C1(n9865), .C2(keyinput81), .A(n9864), .ZN(n9869) );
  XNOR2_X1 U10916 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput106), .ZN(n9867) );
  XNOR2_X1 U10917 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput73), .ZN(n9866) );
  NAND2_X1 U10918 ( .A1(n9867), .A2(n9866), .ZN(n9868) );
  NOR4_X1 U10919 ( .A1(n9871), .A2(n9870), .A3(n9869), .A4(n9868), .ZN(n9909)
         );
  INV_X1 U10920 ( .A(SI_2_), .ZN(n9987) );
  AOI22_X1 U10921 ( .A1(n9873), .A2(keyinput77), .B1(keyinput88), .B2(n9987), 
        .ZN(n9872) );
  OAI221_X1 U10922 ( .B1(n9873), .B2(keyinput77), .C1(n9987), .C2(keyinput88), 
        .A(n9872), .ZN(n9882) );
  INV_X1 U10923 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n10018) );
  AOI22_X1 U10924 ( .A1(n9875), .A2(keyinput105), .B1(keyinput86), .B2(n10018), 
        .ZN(n9874) );
  OAI221_X1 U10925 ( .B1(n9875), .B2(keyinput105), .C1(n10018), .C2(keyinput86), .A(n9874), .ZN(n9881) );
  INV_X1 U10926 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10014) );
  AOI22_X1 U10927 ( .A1(n6566), .A2(keyinput68), .B1(n10014), .B2(keyinput108), 
        .ZN(n9876) );
  OAI221_X1 U10928 ( .B1(n6566), .B2(keyinput68), .C1(n10014), .C2(keyinput108), .A(n9876), .ZN(n9880) );
  AOI22_X1 U10929 ( .A1(n5462), .A2(keyinput74), .B1(n9878), .B2(keyinput64), 
        .ZN(n9877) );
  OAI221_X1 U10930 ( .B1(n5462), .B2(keyinput74), .C1(n9878), .C2(keyinput64), 
        .A(n9877), .ZN(n9879) );
  NOR4_X1 U10931 ( .A1(n9882), .A2(n9881), .A3(n9880), .A4(n9879), .ZN(n9908)
         );
  INV_X1 U10932 ( .A(SI_4_), .ZN(n9993) );
  AOI22_X1 U10933 ( .A1(n9884), .A2(keyinput109), .B1(keyinput76), .B2(n9993), 
        .ZN(n9883) );
  OAI221_X1 U10934 ( .B1(n9884), .B2(keyinput109), .C1(n9993), .C2(keyinput76), 
        .A(n9883), .ZN(n9893) );
  AOI22_X1 U10935 ( .A1(n9886), .A2(keyinput92), .B1(n10013), .B2(keyinput120), 
        .ZN(n9885) );
  OAI221_X1 U10936 ( .B1(n9886), .B2(keyinput92), .C1(n10013), .C2(keyinput120), .A(n9885), .ZN(n9892) );
  AOI22_X1 U10937 ( .A1(n10002), .A2(keyinput122), .B1(keyinput95), .B2(n6578), 
        .ZN(n9887) );
  OAI221_X1 U10938 ( .B1(n10002), .B2(keyinput122), .C1(n6578), .C2(keyinput95), .A(n9887), .ZN(n9891) );
  AOI22_X1 U10939 ( .A1(n9889), .A2(keyinput114), .B1(n10031), .B2(keyinput126), .ZN(n9888) );
  OAI221_X1 U10940 ( .B1(n9889), .B2(keyinput114), .C1(n10031), .C2(
        keyinput126), .A(n9888), .ZN(n9890) );
  NOR4_X1 U10941 ( .A1(n9893), .A2(n9892), .A3(n9891), .A4(n9890), .ZN(n9907)
         );
  AOI22_X1 U10942 ( .A1(n10017), .A2(keyinput113), .B1(n5063), .B2(keyinput69), 
        .ZN(n9894) );
  OAI221_X1 U10943 ( .B1(n10017), .B2(keyinput113), .C1(n5063), .C2(keyinput69), .A(n9894), .ZN(n9905) );
  AOI22_X1 U10944 ( .A1(n9897), .A2(keyinput117), .B1(n9896), .B2(keyinput70), 
        .ZN(n9895) );
  OAI221_X1 U10945 ( .B1(n9897), .B2(keyinput117), .C1(n9896), .C2(keyinput70), 
        .A(n9895), .ZN(n9904) );
  XNOR2_X1 U10946 ( .A(n9898), .B(keyinput85), .ZN(n9903) );
  XNOR2_X1 U10947 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput102), .ZN(n9901) );
  XNOR2_X1 U10948 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput75), .ZN(n9900) );
  XNOR2_X1 U10949 ( .A(keyinput66), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n9899) );
  NAND3_X1 U10950 ( .A1(n9901), .A2(n9900), .A3(n9899), .ZN(n9902) );
  NOR4_X1 U10951 ( .A1(n9905), .A2(n9904), .A3(n9903), .A4(n9902), .ZN(n9906)
         );
  AND4_X1 U10952 ( .A1(n9909), .A2(n9908), .A3(n9907), .A4(n9906), .ZN(n10046)
         );
  OAI22_X1 U10953 ( .A1(P1_REG1_REG_25__SCAN_IN), .A2(keyinput79), .B1(
        P2_D_REG_16__SCAN_IN), .B2(keyinput123), .ZN(n9910) );
  AOI221_X1 U10954 ( .B1(P1_REG1_REG_25__SCAN_IN), .B2(keyinput79), .C1(
        keyinput123), .C2(P2_D_REG_16__SCAN_IN), .A(n9910), .ZN(n9917) );
  OAI22_X1 U10955 ( .A1(P2_D_REG_11__SCAN_IN), .A2(keyinput78), .B1(keyinput98), .B2(P2_ADDR_REG_11__SCAN_IN), .ZN(n9911) );
  AOI221_X1 U10956 ( .B1(P2_D_REG_11__SCAN_IN), .B2(keyinput78), .C1(
        P2_ADDR_REG_11__SCAN_IN), .C2(keyinput98), .A(n9911), .ZN(n9916) );
  OAI22_X1 U10957 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(keyinput115), .B1(
        P2_REG1_REG_1__SCAN_IN), .B2(keyinput111), .ZN(n9912) );
  AOI221_X1 U10958 ( .B1(P2_IR_REG_15__SCAN_IN), .B2(keyinput115), .C1(
        keyinput111), .C2(P2_REG1_REG_1__SCAN_IN), .A(n9912), .ZN(n9915) );
  OAI22_X1 U10959 ( .A1(P1_REG1_REG_21__SCAN_IN), .A2(keyinput93), .B1(
        keyinput119), .B2(P2_D_REG_31__SCAN_IN), .ZN(n9913) );
  AOI221_X1 U10960 ( .B1(P1_REG1_REG_21__SCAN_IN), .B2(keyinput93), .C1(
        P2_D_REG_31__SCAN_IN), .C2(keyinput119), .A(n9913), .ZN(n9914) );
  NAND4_X1 U10961 ( .A1(n9917), .A2(n9916), .A3(n9915), .A4(n9914), .ZN(n9945)
         );
  OAI22_X1 U10962 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput118), .B1(
        keyinput65), .B2(P2_IR_REG_25__SCAN_IN), .ZN(n9918) );
  AOI221_X1 U10963 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput118), .C1(
        P2_IR_REG_25__SCAN_IN), .C2(keyinput65), .A(n9918), .ZN(n9925) );
  OAI22_X1 U10964 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput124), .B1(keyinput91), .B2(P1_REG1_REG_16__SCAN_IN), .ZN(n9919) );
  AOI221_X1 U10965 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput124), .C1(
        P1_REG1_REG_16__SCAN_IN), .C2(keyinput91), .A(n9919), .ZN(n9924) );
  OAI22_X1 U10966 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(keyinput90), .B1(
        keyinput107), .B2(P2_ADDR_REG_12__SCAN_IN), .ZN(n9920) );
  AOI221_X1 U10967 ( .B1(P2_IR_REG_28__SCAN_IN), .B2(keyinput90), .C1(
        P2_ADDR_REG_12__SCAN_IN), .C2(keyinput107), .A(n9920), .ZN(n9923) );
  OAI22_X1 U10968 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(keyinput72), .B1(
        P2_REG2_REG_24__SCAN_IN), .B2(keyinput110), .ZN(n9921) );
  AOI221_X1 U10969 ( .B1(P1_DATAO_REG_5__SCAN_IN), .B2(keyinput72), .C1(
        keyinput110), .C2(P2_REG2_REG_24__SCAN_IN), .A(n9921), .ZN(n9922) );
  NAND4_X1 U10970 ( .A1(n9925), .A2(n9924), .A3(n9923), .A4(n9922), .ZN(n9944)
         );
  OAI22_X1 U10971 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(keyinput89), .B1(
        keyinput116), .B2(P2_ADDR_REG_4__SCAN_IN), .ZN(n9926) );
  AOI221_X1 U10972 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(keyinput89), .C1(
        P2_ADDR_REG_4__SCAN_IN), .C2(keyinput116), .A(n9926), .ZN(n9933) );
  OAI22_X1 U10973 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput104), .B1(
        P1_REG1_REG_24__SCAN_IN), .B2(keyinput127), .ZN(n9927) );
  AOI221_X1 U10974 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput104), .C1(
        keyinput127), .C2(P1_REG1_REG_24__SCAN_IN), .A(n9927), .ZN(n9932) );
  OAI22_X1 U10975 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput121), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput87), .ZN(n9928) );
  AOI221_X1 U10976 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput121), .C1(
        keyinput87), .C2(P2_REG3_REG_22__SCAN_IN), .A(n9928), .ZN(n9931) );
  OAI22_X1 U10977 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput125), .B1(
        keyinput94), .B2(P2_D_REG_8__SCAN_IN), .ZN(n9929) );
  AOI221_X1 U10978 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput125), .C1(
        P2_D_REG_8__SCAN_IN), .C2(keyinput94), .A(n9929), .ZN(n9930) );
  NAND4_X1 U10979 ( .A1(n9933), .A2(n9932), .A3(n9931), .A4(n9930), .ZN(n9943)
         );
  OAI22_X1 U10980 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput71), .B1(
        keyinput96), .B2(P1_REG3_REG_3__SCAN_IN), .ZN(n9934) );
  AOI221_X1 U10981 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput71), .C1(
        P1_REG3_REG_3__SCAN_IN), .C2(keyinput96), .A(n9934), .ZN(n9941) );
  OAI22_X1 U10982 ( .A1(P1_D_REG_22__SCAN_IN), .A2(keyinput99), .B1(
        P2_ADDR_REG_19__SCAN_IN), .B2(keyinput112), .ZN(n9935) );
  AOI221_X1 U10983 ( .B1(P1_D_REG_22__SCAN_IN), .B2(keyinput99), .C1(
        keyinput112), .C2(P2_ADDR_REG_19__SCAN_IN), .A(n9935), .ZN(n9940) );
  OAI22_X1 U10984 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput97), .B1(
        P2_REG2_REG_29__SCAN_IN), .B2(keyinput100), .ZN(n9936) );
  AOI221_X1 U10985 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput97), .C1(
        keyinput100), .C2(P2_REG2_REG_29__SCAN_IN), .A(n9936), .ZN(n9939) );
  OAI22_X1 U10986 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput82), .B1(
        keyinput84), .B2(P1_REG1_REG_31__SCAN_IN), .ZN(n9937) );
  AOI221_X1 U10987 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput82), .C1(
        P1_REG1_REG_31__SCAN_IN), .C2(keyinput84), .A(n9937), .ZN(n9938) );
  NAND4_X1 U10988 ( .A1(n9941), .A2(n9940), .A3(n9939), .A4(n9938), .ZN(n9942)
         );
  NOR4_X1 U10989 ( .A1(n9945), .A2(n9944), .A3(n9943), .A4(n9942), .ZN(n10045)
         );
  AOI22_X1 U10990 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput21), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput17), .ZN(n9946) );
  OAI221_X1 U10991 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput21), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput17), .A(n9946), .ZN(n9953) );
  AOI22_X1 U10992 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(keyinput31), .B1(
        P1_REG0_REG_11__SCAN_IN), .B2(keyinput50), .ZN(n9947) );
  OAI221_X1 U10993 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(keyinput31), .C1(
        P1_REG0_REG_11__SCAN_IN), .C2(keyinput50), .A(n9947), .ZN(n9952) );
  AOI22_X1 U10994 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(keyinput6), .B1(SI_21_), 
        .B2(keyinput13), .ZN(n9948) );
  OAI221_X1 U10995 ( .B1(P1_REG3_REG_9__SCAN_IN), .B2(keyinput6), .C1(SI_21_), 
        .C2(keyinput13), .A(n9948), .ZN(n9951) );
  AOI22_X1 U10996 ( .A1(SI_29_), .A2(keyinput10), .B1(P1_DATAO_REG_5__SCAN_IN), 
        .B2(keyinput8), .ZN(n9949) );
  OAI221_X1 U10997 ( .B1(SI_29_), .B2(keyinput10), .C1(P1_DATAO_REG_5__SCAN_IN), .C2(keyinput8), .A(n9949), .ZN(n9950) );
  NOR4_X1 U10998 ( .A1(n9953), .A2(n9952), .A3(n9951), .A4(n9950), .ZN(n9985)
         );
  AOI22_X1 U10999 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(keyinput9), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(keyinput0), .ZN(n9954) );
  OAI221_X1 U11000 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(keyinput9), .C1(
        P1_DATAO_REG_0__SCAN_IN), .C2(keyinput0), .A(n9954), .ZN(n9961) );
  AOI22_X1 U11001 ( .A1(P2_D_REG_16__SCAN_IN), .A2(keyinput59), .B1(
        P2_IR_REG_12__SCAN_IN), .B2(keyinput38), .ZN(n9955) );
  OAI221_X1 U11002 ( .B1(P2_D_REG_16__SCAN_IN), .B2(keyinput59), .C1(
        P2_IR_REG_12__SCAN_IN), .C2(keyinput38), .A(n9955), .ZN(n9960) );
  AOI22_X1 U11003 ( .A1(P2_REG1_REG_1__SCAN_IN), .A2(keyinput47), .B1(
        P1_REG1_REG_25__SCAN_IN), .B2(keyinput15), .ZN(n9956) );
  OAI221_X1 U11004 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(keyinput47), .C1(
        P1_REG1_REG_25__SCAN_IN), .C2(keyinput15), .A(n9956), .ZN(n9959) );
  AOI22_X1 U11005 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(keyinput34), .B1(
        P2_IR_REG_28__SCAN_IN), .B2(keyinput26), .ZN(n9957) );
  OAI221_X1 U11006 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(keyinput34), .C1(
        P2_IR_REG_28__SCAN_IN), .C2(keyinput26), .A(n9957), .ZN(n9958) );
  NOR4_X1 U11007 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n9984)
         );
  AOI22_X1 U11008 ( .A1(P2_D_REG_20__SCAN_IN), .A2(keyinput53), .B1(
        P1_REG1_REG_24__SCAN_IN), .B2(keyinput63), .ZN(n9962) );
  OAI221_X1 U11009 ( .B1(P2_D_REG_20__SCAN_IN), .B2(keyinput53), .C1(
        P1_REG1_REG_24__SCAN_IN), .C2(keyinput63), .A(n9962), .ZN(n9969) );
  AOI22_X1 U11010 ( .A1(P2_D_REG_14__SCAN_IN), .A2(keyinput3), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(keyinput45), .ZN(n9963) );
  OAI221_X1 U11011 ( .B1(P2_D_REG_14__SCAN_IN), .B2(keyinput3), .C1(
        P1_DATAO_REG_16__SCAN_IN), .C2(keyinput45), .A(n9963), .ZN(n9968) );
  AOI22_X1 U11012 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(keyinput43), .B1(
        P2_IR_REG_2__SCAN_IN), .B2(keyinput41), .ZN(n9964) );
  OAI221_X1 U11013 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(keyinput43), .C1(
        P2_IR_REG_2__SCAN_IN), .C2(keyinput41), .A(n9964), .ZN(n9967) );
  AOI22_X1 U11014 ( .A1(P1_REG1_REG_31__SCAN_IN), .A2(keyinput20), .B1(
        P2_D_REG_8__SCAN_IN), .B2(keyinput30), .ZN(n9965) );
  OAI221_X1 U11015 ( .B1(P1_REG1_REG_31__SCAN_IN), .B2(keyinput20), .C1(
        P2_D_REG_8__SCAN_IN), .C2(keyinput30), .A(n9965), .ZN(n9966) );
  NOR4_X1 U11016 ( .A1(n9969), .A2(n9968), .A3(n9967), .A4(n9966), .ZN(n9983)
         );
  AOI22_X1 U11017 ( .A1(n9972), .A2(keyinput32), .B1(keyinput39), .B2(n9971), 
        .ZN(n9970) );
  OAI221_X1 U11018 ( .B1(n9972), .B2(keyinput32), .C1(n9971), .C2(keyinput39), 
        .A(n9970), .ZN(n9981) );
  AOI22_X1 U11019 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(keyinput11), .B1(n9974), 
        .B2(keyinput35), .ZN(n9973) );
  OAI221_X1 U11020 ( .B1(P2_IR_REG_14__SCAN_IN), .B2(keyinput11), .C1(n9974), 
        .C2(keyinput35), .A(n9973), .ZN(n9980) );
  AOI22_X1 U11021 ( .A1(P2_D_REG_31__SCAN_IN), .A2(keyinput55), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(keyinput28), .ZN(n9975) );
  OAI221_X1 U11022 ( .B1(P2_D_REG_31__SCAN_IN), .B2(keyinput55), .C1(
        P1_DATAO_REG_23__SCAN_IN), .C2(keyinput28), .A(n9975), .ZN(n9979) );
  XOR2_X1 U11023 ( .A(n5063), .B(keyinput5), .Z(n9977) );
  XNOR2_X1 U11024 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput48), .ZN(n9976) );
  NAND2_X1 U11025 ( .A1(n9977), .A2(n9976), .ZN(n9978) );
  NOR4_X1 U11026 ( .A1(n9981), .A2(n9980), .A3(n9979), .A4(n9978), .ZN(n9982)
         );
  NAND4_X1 U11027 ( .A1(n9985), .A2(n9984), .A3(n9983), .A4(n9982), .ZN(n10044) );
  AOI22_X1 U11028 ( .A1(n4898), .A2(keyinput46), .B1(n9987), .B2(keyinput24), 
        .ZN(n9986) );
  OAI221_X1 U11029 ( .B1(n4898), .B2(keyinput46), .C1(n9987), .C2(keyinput24), 
        .A(n9986), .ZN(n9999) );
  AOI22_X1 U11030 ( .A1(n9990), .A2(keyinput33), .B1(keyinput18), .B2(n9989), 
        .ZN(n9988) );
  OAI221_X1 U11031 ( .B1(n9990), .B2(keyinput33), .C1(n9989), .C2(keyinput18), 
        .A(n9988), .ZN(n9998) );
  INV_X1 U11032 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9992) );
  AOI22_X1 U11033 ( .A1(n9993), .A2(keyinput12), .B1(keyinput29), .B2(n9992), 
        .ZN(n9991) );
  OAI221_X1 U11034 ( .B1(n9993), .B2(keyinput12), .C1(n9992), .C2(keyinput29), 
        .A(n9991), .ZN(n9997) );
  XNOR2_X1 U11035 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput42), .ZN(n9995) );
  XNOR2_X1 U11036 ( .A(keyinput2), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U11037 ( .A1(n9995), .A2(n9994), .ZN(n9996) );
  NOR4_X1 U11038 ( .A1(n9999), .A2(n9998), .A3(n9997), .A4(n9996), .ZN(n10042)
         );
  INV_X1 U11039 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10001) );
  AOI22_X1 U11040 ( .A1(n10002), .A2(keyinput58), .B1(keyinput52), .B2(n10001), 
        .ZN(n10000) );
  OAI221_X1 U11041 ( .B1(n10002), .B2(keyinput58), .C1(n10001), .C2(keyinput52), .A(n10000), .ZN(n10011) );
  INV_X1 U11042 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10004) );
  AOI22_X1 U11043 ( .A1(n7751), .A2(keyinput25), .B1(keyinput27), .B2(n10004), 
        .ZN(n10003) );
  OAI221_X1 U11044 ( .B1(n7751), .B2(keyinput25), .C1(n10004), .C2(keyinput27), 
        .A(n10003), .ZN(n10010) );
  XNOR2_X1 U11045 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput54), .ZN(n10008)
         );
  XNOR2_X1 U11046 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput57), .ZN(n10007) );
  XNOR2_X1 U11047 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput51), .ZN(n10006) );
  XNOR2_X1 U11048 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput7), .ZN(n10005)
         );
  NAND4_X1 U11049 ( .A1(n10008), .A2(n10007), .A3(n10006), .A4(n10005), .ZN(
        n10009) );
  NOR3_X1 U11050 ( .A1(n10011), .A2(n10010), .A3(n10009), .ZN(n10041) );
  AOI22_X1 U11051 ( .A1(n10014), .A2(keyinput44), .B1(n10013), .B2(keyinput56), 
        .ZN(n10012) );
  OAI221_X1 U11052 ( .B1(n10014), .B2(keyinput44), .C1(n10013), .C2(keyinput56), .A(n10012), .ZN(n10025) );
  AOI22_X1 U11053 ( .A1(n10017), .A2(keyinput49), .B1(n10016), .B2(keyinput40), 
        .ZN(n10015) );
  OAI221_X1 U11054 ( .B1(n10017), .B2(keyinput49), .C1(n10016), .C2(keyinput40), .A(n10015), .ZN(n10024) );
  XOR2_X1 U11055 ( .A(n5028), .B(keyinput19), .Z(n10022) );
  XOR2_X1 U11056 ( .A(n10018), .B(keyinput22), .Z(n10021) );
  XNOR2_X1 U11057 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput61), .ZN(n10020) );
  XNOR2_X1 U11058 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput1), .ZN(n10019) );
  NAND4_X1 U11059 ( .A1(n10022), .A2(n10021), .A3(n10020), .A4(n10019), .ZN(
        n10023) );
  NOR3_X1 U11060 ( .A1(n10025), .A2(n10024), .A3(n10023), .ZN(n10040) );
  AOI22_X1 U11061 ( .A1(n10027), .A2(keyinput14), .B1(keyinput4), .B2(n6566), 
        .ZN(n10026) );
  OAI221_X1 U11062 ( .B1(n10027), .B2(keyinput14), .C1(n6566), .C2(keyinput4), 
        .A(n10026), .ZN(n10038) );
  AOI22_X1 U11063 ( .A1(n10029), .A2(keyinput23), .B1(n5866), .B2(keyinput16), 
        .ZN(n10028) );
  OAI221_X1 U11064 ( .B1(n10029), .B2(keyinput23), .C1(n5866), .C2(keyinput16), 
        .A(n10028), .ZN(n10037) );
  AOI22_X1 U11065 ( .A1(n10032), .A2(keyinput60), .B1(keyinput62), .B2(n10031), 
        .ZN(n10030) );
  OAI221_X1 U11066 ( .B1(n10032), .B2(keyinput60), .C1(n10031), .C2(keyinput62), .A(n10030), .ZN(n10036) );
  AOI22_X1 U11067 ( .A1(n10034), .A2(keyinput37), .B1(keyinput36), .B2(n7702), 
        .ZN(n10033) );
  OAI221_X1 U11068 ( .B1(n10034), .B2(keyinput37), .C1(n7702), .C2(keyinput36), 
        .A(n10033), .ZN(n10035) );
  NOR4_X1 U11069 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10035), .ZN(
        n10039) );
  NAND4_X1 U11070 ( .A1(n10042), .A2(n10041), .A3(n10040), .A4(n10039), .ZN(
        n10043) );
  AOI211_X1 U11071 ( .C1(n10046), .C2(n10045), .A(n10044), .B(n10043), .ZN(
        n10047) );
  XNOR2_X1 U11072 ( .A(n10048), .B(n10047), .ZN(P1_U3309) );
  XOR2_X1 U11073 ( .A(n10049), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11074 ( .A1(n10051), .A2(n10050), .ZN(n10052) );
  XOR2_X1 U11075 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10052), .Z(ADD_1071_U51) );
  OAI21_X1 U11076 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(n10056) );
  XNOR2_X1 U11077 ( .A(n10056), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11078 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(ADD_1071_U47) );
  XOR2_X1 U11079 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10060), .Z(ADD_1071_U48) );
  XOR2_X1 U11080 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10061), .Z(ADD_1071_U49) );
  XOR2_X1 U11081 ( .A(n10063), .B(n10062), .Z(ADD_1071_U54) );
  XOR2_X1 U11082 ( .A(n10065), .B(n10064), .Z(ADD_1071_U53) );
  XNOR2_X1 U11083 ( .A(n10067), .B(n10066), .ZN(ADD_1071_U52) );
  CLKBUF_X3 U4888 ( .A(n4919), .Z(n5942) );
  AND4_X1 U4815 ( .A1(n5165), .A2(n5230), .A3(n5164), .A4(n4878), .ZN(n4880)
         );
  CLKBUF_X1 U4827 ( .A(n5614), .Z(n8195) );
  NAND2_X2 U6370 ( .A1(n5749), .A2(n7725), .ZN(n5147) );
  OR2_X1 U6530 ( .A1(n9754), .A2(n5640), .ZN(n9742) );
  CLKBUF_X1 U7230 ( .A(n9071), .Z(n4307) );
endmodule

